magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1260 -1260 137880 84568
<< dnwell >>
rect 1822 1724 134872 81473
<< nwell >>
rect 1738 81389 134956 81557
rect 1738 1808 1906 81389
rect 134788 1808 134956 81389
rect 1738 1640 134956 1808
<< metal1 >>
rect 1710 81361 134984 81585
rect 1790 80994 1854 81046
rect 134840 80994 134904 81046
rect 1790 80658 1854 80710
rect 134840 80658 134904 80710
rect 1790 80322 1854 80374
rect 134840 80322 134904 80374
rect 1790 79986 1854 80038
rect 134840 79986 134904 80038
rect 1790 79650 1854 79702
rect 134840 79650 134904 79702
rect 1790 79314 1854 79366
rect 134840 79314 134904 79366
rect 1790 78978 1854 79030
rect 134840 78978 134904 79030
rect 1790 78642 1854 78694
rect 134840 78642 134904 78694
rect 1790 78306 1854 78358
rect 134840 78306 134904 78358
rect 1790 77970 1854 78022
rect 134840 77970 134904 78022
rect 1790 77634 1854 77686
rect 134840 77634 134904 77686
rect 1790 77298 1854 77350
rect 134840 77298 134904 77350
rect 1790 76962 1854 77014
rect 134840 76962 134904 77014
rect 1790 76626 1854 76678
rect 134840 76626 134904 76678
rect 1790 76290 1854 76342
rect 134840 76290 134904 76342
rect 1790 75954 1854 76006
rect 134840 75954 134904 76006
rect 1790 75618 1854 75670
rect 134840 75618 134904 75670
rect 1790 75282 1854 75334
rect 134840 75282 134904 75334
rect 1790 74946 1854 74998
rect 134840 74946 134904 74998
rect 1790 74610 1854 74662
rect 134840 74610 134904 74662
rect 1790 74274 1854 74326
rect 134840 74274 134904 74326
rect 1790 73938 1854 73990
rect 134840 73938 134904 73990
rect 1790 73602 1854 73654
rect 134840 73602 134904 73654
rect 1790 73266 1854 73318
rect 134840 73266 134904 73318
rect 1790 72930 1854 72982
rect 134840 72930 134904 72982
rect 1790 72594 1854 72646
rect 134840 72594 134904 72646
rect 1790 72258 1854 72310
rect 134840 72258 134904 72310
rect 1790 71922 1854 71974
rect 134840 71922 134904 71974
rect 1790 71586 1854 71638
rect 134840 71586 134904 71638
rect 1790 71250 1854 71302
rect 134840 71250 134904 71302
rect 1790 70914 1854 70966
rect 134840 70914 134904 70966
rect 1790 70578 1854 70630
rect 134840 70578 134904 70630
rect 1790 70242 1854 70294
rect 134840 70242 134904 70294
rect 1790 69906 1854 69958
rect 134840 69906 134904 69958
rect 1790 69570 1854 69622
rect 134840 69570 134904 69622
rect 1790 69234 1854 69286
rect 134840 69234 134904 69286
rect 1790 68898 1854 68950
rect 134840 68898 134904 68950
rect 1790 68562 1854 68614
rect 134840 68562 134904 68614
rect 1790 68226 1854 68278
rect 134840 68226 134904 68278
rect 1790 67890 1854 67942
rect 134840 67890 134904 67942
rect 1790 67554 1854 67606
rect 134840 67554 134904 67606
rect 1790 67218 1854 67270
rect 134840 67218 134904 67270
rect 1790 66882 1854 66934
rect 134840 66882 134904 66934
rect 1790 66546 1854 66598
rect 134840 66546 134904 66598
rect 1790 66210 1854 66262
rect 134840 66210 134904 66262
rect 1790 65874 1854 65926
rect 134840 65874 134904 65926
rect 1790 65538 1854 65590
rect 134840 65538 134904 65590
rect 1790 65202 1854 65254
rect 134840 65202 134904 65254
rect 1790 64866 1854 64918
rect 134840 64866 134904 64918
rect 1790 64530 1854 64582
rect 134840 64530 134904 64582
rect 1790 64194 1854 64246
rect 134840 64194 134904 64246
rect 1790 63858 1854 63910
rect 134840 63858 134904 63910
rect 1790 63522 1854 63574
rect 134840 63522 134904 63574
rect 1790 63186 1854 63238
rect 134840 63186 134904 63238
rect 1790 62850 1854 62902
rect 134840 62850 134904 62902
rect 1790 62514 1854 62566
rect 134840 62514 134904 62566
rect 1790 62178 1854 62230
rect 134840 62178 134904 62230
rect 1790 61842 1854 61894
rect 134840 61842 134904 61894
rect 1790 61506 1854 61558
rect 134840 61506 134904 61558
rect 1790 61170 1854 61222
rect 134840 61170 134904 61222
rect 1790 60834 1854 60886
rect 134840 60834 134904 60886
rect 1790 60498 1854 60550
rect 134840 60498 134904 60550
rect 1790 60162 1854 60214
rect 134840 60162 134904 60214
rect 1790 59826 1854 59878
rect 134840 59826 134904 59878
rect 1790 59490 1854 59542
rect 134840 59490 134904 59542
rect 1790 59154 1854 59206
rect 134840 59154 134904 59206
rect 1790 58818 1854 58870
rect 134840 58818 134904 58870
rect 1790 58482 1854 58534
rect 134840 58482 134904 58534
rect 1790 58146 1854 58198
rect 134840 58146 134904 58198
rect 1790 57810 1854 57862
rect 134840 57810 134904 57862
rect 1790 57474 1854 57526
rect 134840 57474 134904 57526
rect 1790 57138 1854 57190
rect 134840 57138 134904 57190
rect 1790 56802 1854 56854
rect 134840 56802 134904 56854
rect 1790 56466 1854 56518
rect 134840 56466 134904 56518
rect 1790 56130 1854 56182
rect 134840 56130 134904 56182
rect 1790 55794 1854 55846
rect 134840 55794 134904 55846
rect 1790 55458 1854 55510
rect 134840 55458 134904 55510
rect 1790 55122 1854 55174
rect 134840 55122 134904 55174
rect 1790 54786 1854 54838
rect 134840 54786 134904 54838
rect 1790 54450 1854 54502
rect 134840 54450 134904 54502
rect 1790 54114 1854 54166
rect 134840 54114 134904 54166
rect 1790 53778 1854 53830
rect 134840 53778 134904 53830
rect 1790 53442 1854 53494
rect 134840 53442 134904 53494
rect 1790 53106 1854 53158
rect 134840 53106 134904 53158
rect 1790 52770 1854 52822
rect 134840 52770 134904 52822
rect 1790 52434 1854 52486
rect 134840 52434 134904 52486
rect 1790 52098 1854 52150
rect 134840 52098 134904 52150
rect 1790 51762 1854 51814
rect 134840 51762 134904 51814
rect 1790 51426 1854 51478
rect 134840 51426 134904 51478
rect 1790 51090 1854 51142
rect 134840 51090 134904 51142
rect 1790 50754 1854 50806
rect 134840 50754 134904 50806
rect 1790 50418 1854 50470
rect 134840 50418 134904 50470
rect 1790 50082 1854 50134
rect 134840 50082 134904 50134
rect 1790 49746 1854 49798
rect 134840 49746 134904 49798
rect 1790 49410 1854 49462
rect 134840 49410 134904 49462
rect 1790 49074 1854 49126
rect 134840 49074 134904 49126
rect 1790 48738 1854 48790
rect 134840 48738 134904 48790
rect 1790 48402 1854 48454
rect 134840 48402 134904 48454
rect 1790 48066 1854 48118
rect 134840 48066 134904 48118
rect 1790 47730 1854 47782
rect 134840 47730 134904 47782
rect 1790 47394 1854 47446
rect 134840 47394 134904 47446
rect 1790 47058 1854 47110
rect 134840 47058 134904 47110
rect 1790 46722 1854 46774
rect 134840 46722 134904 46774
rect 1790 46386 1854 46438
rect 134840 46386 134904 46438
rect 1790 46050 1854 46102
rect 134840 46050 134904 46102
rect 1790 45714 1854 45766
rect 134840 45714 134904 45766
rect 1790 45378 1854 45430
rect 134840 45378 134904 45430
rect 1790 45042 1854 45094
rect 134840 45042 134904 45094
rect 1790 44706 1854 44758
rect 134840 44706 134904 44758
rect 1790 44370 1854 44422
rect 134840 44370 134904 44422
rect 1790 44034 1854 44086
rect 134840 44034 134904 44086
rect 1790 43698 1854 43750
rect 134840 43698 134904 43750
rect 1790 43362 1854 43414
rect 134840 43362 134904 43414
rect 1790 43026 1854 43078
rect 134840 43026 134904 43078
rect 1790 42690 1854 42742
rect 134840 42690 134904 42742
rect 1790 42354 1854 42406
rect 134840 42354 134904 42406
rect 1790 42018 1854 42070
rect 134840 42018 134904 42070
rect 1790 41682 1854 41734
rect 134840 41682 134904 41734
rect 1790 41346 1854 41398
rect 134840 41346 134904 41398
rect 1790 41010 1854 41062
rect 134840 41010 134904 41062
rect 1790 40674 1854 40726
rect 134840 40674 134904 40726
rect 1790 40338 1854 40390
rect 134840 40338 134904 40390
rect 1790 40002 1854 40054
rect 134840 40002 134904 40054
rect 1790 39666 1854 39718
rect 134840 39666 134904 39718
rect 1790 39330 1854 39382
rect 134840 39330 134904 39382
rect 1790 38994 1854 39046
rect 134840 38994 134904 39046
rect 1790 38658 1854 38710
rect 134840 38658 134904 38710
rect 1790 38322 1854 38374
rect 134840 38322 134904 38374
rect 1790 37986 1854 38038
rect 134840 37986 134904 38038
rect 1790 37650 1854 37702
rect 134840 37650 134904 37702
rect 1790 37314 1854 37366
rect 134840 37314 134904 37366
rect 1790 36978 1854 37030
rect 134840 36978 134904 37030
rect 1790 36642 1854 36694
rect 1790 36306 1854 36358
rect 1790 35970 1854 36022
rect 1790 35634 1854 35686
rect 1790 35298 1854 35350
rect 1790 34962 1854 35014
rect 1790 34626 1854 34678
rect 1790 34290 1854 34342
rect 1790 33954 1854 34006
rect 1790 33618 1854 33670
rect 1790 33282 1854 33334
rect 1790 32946 1854 32998
rect 1790 32610 1854 32662
rect 1790 32274 1854 32326
rect 1790 31938 1854 31990
rect 1790 31602 1854 31654
rect 1790 31266 1854 31318
rect 1790 30930 1854 30982
rect 1790 30594 1854 30646
rect 1790 30258 1854 30310
rect 1790 29922 1854 29974
rect 1790 29586 1854 29638
rect 1790 29250 1854 29302
rect 1790 28914 1854 28966
rect 1790 28578 1854 28630
rect 1790 28242 1854 28294
rect 1790 27906 1854 27958
rect 1790 27570 1854 27622
rect 1790 27234 1854 27286
rect 1790 26898 1854 26950
rect 1790 26562 1854 26614
rect 1790 26226 1854 26278
rect 1790 25890 1854 25942
rect 1790 25554 1854 25606
rect 1790 25218 1854 25270
rect 1790 24882 1854 24934
rect 1790 24546 1854 24598
rect 1790 24210 1854 24262
rect 1790 23874 1854 23926
rect 14881 23796 14909 28381
rect 14961 23796 14989 29939
rect 15041 23796 15069 31209
rect 15121 23796 15149 32767
rect 15201 23796 15229 34037
rect 15281 23796 15309 35595
rect 15361 23796 15389 36865
rect 134840 36642 134904 36694
rect 134840 36306 134904 36358
rect 134840 35970 134904 36022
rect 134840 35634 134904 35686
rect 134840 35298 134904 35350
rect 134840 34962 134904 35014
rect 134840 34626 134904 34678
rect 134840 34290 134904 34342
rect 134840 33954 134904 34006
rect 134840 33618 134904 33670
rect 134840 33282 134904 33334
rect 134840 32946 134904 32998
rect 134840 32610 134904 32662
rect 134840 32274 134904 32326
rect 134840 31938 134904 31990
rect 134840 31602 134904 31654
rect 134840 31266 134904 31318
rect 134840 30930 134904 30982
rect 134840 30594 134904 30646
rect 134840 30258 134904 30310
rect 134840 29922 134904 29974
rect 134840 29586 134904 29638
rect 134840 29250 134904 29302
rect 134840 28914 134904 28966
rect 134840 28578 134904 28630
rect 134840 28242 134904 28294
rect 134840 27906 134904 27958
rect 134840 27570 134904 27622
rect 134840 27234 134904 27286
rect 134840 26898 134904 26950
rect 134840 26562 134904 26614
rect 134840 26226 134904 26278
rect 134840 25890 134904 25942
rect 134840 25554 134904 25606
rect 134840 25218 134904 25270
rect 134840 24882 134904 24934
rect 134840 24546 134904 24598
rect 134840 24210 134904 24262
rect 134840 23874 134904 23926
rect 1790 23538 1854 23590
rect 1790 23202 1854 23254
rect 1790 22866 1854 22918
rect 1790 22530 1854 22582
rect 1790 22194 1854 22246
rect 1790 21858 1854 21910
rect 1790 21522 1854 21574
rect 1790 21186 1854 21238
rect 1790 20850 1854 20902
rect 1790 20514 1854 20566
rect 1790 20178 1854 20230
rect 1790 19842 1854 19894
rect 1790 19506 1854 19558
rect 1790 19170 1854 19222
rect 1790 18834 1854 18886
rect 1790 18498 1854 18550
rect 1790 18162 1854 18214
rect 1790 17826 1854 17878
rect 1790 17490 1854 17542
rect 1790 17154 1854 17206
rect 1790 16818 1854 16870
rect 1790 16482 1854 16534
rect 1790 16146 1854 16198
rect 1790 15810 1854 15862
rect 1790 15474 1854 15526
rect 1790 15138 1854 15190
rect 1790 14802 1854 14854
rect 1790 14466 1854 14518
rect 1790 14130 1854 14182
rect 1790 13794 1854 13846
rect 1790 13458 1854 13510
rect 1790 13122 1854 13174
rect 1790 12786 1854 12838
rect 1790 12450 1854 12502
rect 1790 12114 1854 12166
rect 1790 11778 1854 11830
rect 1790 11442 1854 11494
rect 1790 11106 1854 11158
rect 1790 10770 1854 10822
rect 121521 10727 121549 23796
rect 121601 11997 121629 23796
rect 121681 13555 121709 23796
rect 121761 14825 121789 23796
rect 121841 16383 121869 23796
rect 121921 17653 121949 23796
rect 122001 19211 122029 23796
rect 134840 23538 134904 23590
rect 134840 23202 134904 23254
rect 134840 22866 134904 22918
rect 134840 22530 134904 22582
rect 134840 22194 134904 22246
rect 134840 21858 134904 21910
rect 134840 21522 134904 21574
rect 134840 21186 134904 21238
rect 134840 20850 134904 20902
rect 134840 20514 134904 20566
rect 134840 20178 134904 20230
rect 134840 19842 134904 19894
rect 134840 19506 134904 19558
rect 134840 19170 134904 19222
rect 134840 18834 134904 18886
rect 134840 18498 134904 18550
rect 134840 18162 134904 18214
rect 134840 17826 134904 17878
rect 134840 17490 134904 17542
rect 134840 17154 134904 17206
rect 134840 16818 134904 16870
rect 134840 16482 134904 16534
rect 134840 16146 134904 16198
rect 134840 15810 134904 15862
rect 134840 15474 134904 15526
rect 134840 15138 134904 15190
rect 134840 14802 134904 14854
rect 134840 14466 134904 14518
rect 134840 14130 134904 14182
rect 134840 13794 134904 13846
rect 134840 13458 134904 13510
rect 134840 13122 134904 13174
rect 134840 12786 134904 12838
rect 134840 12450 134904 12502
rect 134840 12114 134904 12166
rect 134840 11778 134904 11830
rect 134840 11442 134904 11494
rect 134840 11106 134904 11158
rect 134840 10770 134904 10822
rect 1790 10434 1854 10486
rect 134840 10434 134904 10486
rect 1790 10098 1854 10150
rect 134840 10098 134904 10150
rect 1790 9762 1854 9814
rect 134840 9762 134904 9814
rect 1790 9426 1854 9478
rect 134840 9426 134904 9478
rect 1790 9090 1854 9142
rect 134840 9090 134904 9142
rect 1790 8754 1854 8806
rect 134840 8754 134904 8806
rect 1790 8418 1854 8470
rect 134840 8418 134904 8470
rect 1790 8082 1854 8134
rect 134840 8082 134904 8134
rect 1790 7746 1854 7798
rect 134840 7746 134904 7798
rect 1790 7410 1854 7462
rect 134840 7410 134904 7462
rect 1790 7074 1854 7126
rect 134840 7074 134904 7126
rect 1790 6738 1854 6790
rect 134840 6738 134904 6790
rect 1790 6402 1854 6454
rect 134840 6402 134904 6454
rect 1790 6066 1854 6118
rect 134840 6066 134904 6118
rect 1790 5730 1854 5782
rect 134840 5730 134904 5782
rect 1790 5394 1854 5446
rect 134840 5394 134904 5446
rect 1790 5058 1854 5110
rect 134840 5058 134904 5110
rect 1790 4722 1854 4774
rect 134840 4722 134904 4774
rect 1790 4386 1854 4438
rect 134840 4386 134904 4438
rect 1790 4050 1854 4102
rect 134840 4050 134904 4102
rect 1790 3714 1854 3766
rect 134840 3714 134904 3766
rect 1790 3378 1854 3430
rect 134840 3378 134904 3430
rect 1790 3042 1854 3094
rect 134840 3042 134904 3094
rect 1790 2706 1854 2758
rect 134840 2706 134904 2758
rect 1790 2370 1854 2422
rect 134840 2370 134904 2422
rect 1790 2034 1854 2086
rect 134840 2034 134904 2086
rect 1710 1612 134984 1836
<< metal2 >>
rect 1710 1612 1934 81585
rect 2130 81449 2186 81497
rect 3810 81449 3866 81497
rect 5490 81449 5546 81497
rect 7170 81449 7226 81497
rect 8850 81449 8906 81497
rect 10530 81449 10586 81497
rect 12210 81449 12266 81497
rect 13890 81449 13946 81497
rect 15570 81449 15626 81497
rect 17250 81449 17306 81497
rect 18930 81449 18986 81497
rect 20610 81449 20666 81497
rect 22290 81449 22346 81497
rect 23970 81449 24026 81497
rect 25650 81449 25706 81497
rect 27330 81449 27386 81497
rect 29010 81449 29066 81497
rect 30690 81449 30746 81497
rect 32370 81449 32426 81497
rect 34050 81449 34106 81497
rect 35730 81449 35786 81497
rect 37410 81449 37466 81497
rect 39090 81449 39146 81497
rect 40770 81449 40826 81497
rect 42450 81449 42506 81497
rect 44130 81449 44186 81497
rect 45810 81449 45866 81497
rect 47490 81449 47546 81497
rect 49170 81449 49226 81497
rect 50850 81449 50906 81497
rect 52530 81449 52586 81497
rect 54210 81449 54266 81497
rect 55890 81449 55946 81497
rect 57570 81449 57626 81497
rect 59250 81449 59306 81497
rect 60930 81449 60986 81497
rect 62610 81449 62666 81497
rect 64290 81449 64346 81497
rect 65970 81449 66026 81497
rect 67650 81449 67706 81497
rect 69330 81449 69386 81497
rect 71010 81449 71066 81497
rect 72690 81449 72746 81497
rect 74370 81449 74426 81497
rect 76050 81449 76106 81497
rect 77730 81449 77786 81497
rect 79410 81449 79466 81497
rect 81090 81449 81146 81497
rect 82770 81449 82826 81497
rect 84450 81449 84506 81497
rect 86130 81449 86186 81497
rect 87810 81449 87866 81497
rect 89490 81449 89546 81497
rect 91170 81449 91226 81497
rect 92850 81449 92906 81497
rect 94530 81449 94586 81497
rect 96210 81449 96266 81497
rect 97890 81449 97946 81497
rect 99570 81449 99626 81497
rect 101250 81449 101306 81497
rect 102930 81449 102986 81497
rect 104610 81449 104666 81497
rect 106290 81449 106346 81497
rect 107970 81449 108026 81497
rect 109650 81449 109706 81497
rect 111330 81449 111386 81497
rect 113010 81449 113066 81497
rect 114690 81449 114746 81497
rect 116370 81449 116426 81497
rect 118050 81449 118106 81497
rect 119730 81449 119786 81497
rect 121410 81449 121466 81497
rect 123090 81449 123146 81497
rect 124770 81449 124826 81497
rect 126450 81449 126506 81497
rect 128130 81449 128186 81497
rect 129810 81449 129866 81497
rect 131490 81449 131546 81497
rect 133170 81449 133226 81497
rect 122202 79111 122230 80493
rect 122202 79083 122300 79111
rect 28618 76995 28674 77043
rect 31114 76995 31170 77043
rect 33610 76995 33666 77043
rect 36106 76995 36162 77043
rect 38602 76995 38658 77043
rect 41098 76995 41154 77043
rect 43594 76995 43650 77043
rect 46090 76995 46146 77043
rect 48586 76995 48642 77043
rect 51082 76995 51138 77043
rect 53578 76995 53634 77043
rect 56074 76995 56130 77043
rect 58570 76995 58626 77043
rect 61066 76995 61122 77043
rect 63562 76995 63618 77043
rect 66058 76995 66114 77043
rect 68554 76995 68610 77043
rect 71050 76995 71106 77043
rect 73546 76995 73602 77043
rect 76042 76995 76098 77043
rect 78538 76995 78594 77043
rect 81034 76995 81090 77043
rect 83530 76995 83586 77043
rect 86026 76995 86082 77043
rect 88522 76995 88578 77043
rect 91018 76995 91074 77043
rect 93514 76995 93570 77043
rect 96010 76995 96066 77043
rect 98506 76995 98562 77043
rect 101002 76995 101058 77043
rect 103498 76995 103554 77043
rect 105994 76995 106050 77043
rect 110061 74892 110117 74915
rect 110075 71182 110103 74855
rect 110199 71182 110227 73441
rect 114060 70705 114088 72027
rect 15347 36841 15403 36889
rect 15267 35571 15323 35619
rect 15187 34013 15243 34061
rect 15107 32743 15163 32791
rect 15027 31185 15083 31233
rect 14947 29915 15003 29963
rect 14867 28357 14923 28405
rect 14764 8341 14792 28054
rect 22822 18225 22850 19547
rect 122202 19538 122230 79083
rect 121987 19187 122043 19235
rect 26525 15397 26553 19070
rect 121907 17629 121963 17677
rect 121827 16359 121883 16407
rect 121747 14801 121803 14849
rect 26649 9457 26677 12569
rect 26773 9457 26801 13983
rect 121667 13531 121723 13579
rect 28618 13209 28674 13257
rect 31114 13209 31170 13257
rect 33610 13209 33666 13257
rect 36106 13209 36162 13257
rect 38602 13209 38658 13257
rect 41098 13209 41154 13257
rect 43594 13209 43650 13257
rect 46090 13209 46146 13257
rect 48586 13209 48642 13257
rect 51082 13209 51138 13257
rect 53578 13209 53634 13257
rect 56074 13209 56130 13257
rect 58570 13209 58626 13257
rect 61066 13209 61122 13257
rect 63562 13209 63618 13257
rect 66058 13209 66114 13257
rect 68554 13209 68610 13257
rect 71050 13209 71106 13257
rect 73546 13209 73602 13257
rect 76042 13209 76098 13257
rect 78538 13209 78594 13257
rect 81034 13209 81090 13257
rect 83530 13209 83586 13257
rect 86026 13209 86082 13257
rect 88522 13209 88578 13257
rect 91018 13209 91074 13257
rect 93514 13209 93570 13257
rect 96010 13209 96066 13257
rect 98506 13209 98562 13257
rect 101002 13209 101058 13257
rect 103498 13209 103554 13257
rect 105994 13209 106050 13257
rect 121587 11973 121643 12021
rect 121507 10703 121563 10751
rect 14694 8313 14792 8341
rect 14764 2704 14792 8313
rect 2130 1700 2186 1748
rect 3810 1700 3866 1748
rect 5490 1700 5546 1748
rect 7170 1700 7226 1748
rect 8850 1700 8906 1748
rect 10530 1700 10586 1748
rect 12210 1700 12266 1748
rect 13890 1700 13946 1748
rect 15570 1700 15626 1748
rect 17250 1700 17306 1748
rect 18930 1700 18986 1748
rect 20610 1700 20666 1748
rect 22290 1700 22346 1748
rect 23970 1700 24026 1748
rect 25650 1700 25706 1748
rect 27330 1700 27386 1748
rect 29010 1700 29066 1748
rect 30690 1700 30746 1748
rect 32370 1700 32426 1748
rect 34050 1700 34106 1748
rect 35730 1700 35786 1748
rect 37410 1700 37466 1748
rect 39090 1700 39146 1748
rect 40770 1700 40826 1748
rect 42450 1700 42506 1748
rect 44130 1700 44186 1748
rect 45810 1700 45866 1748
rect 47490 1700 47546 1748
rect 49170 1700 49226 1748
rect 50850 1700 50906 1748
rect 52530 1700 52586 1748
rect 54210 1700 54266 1748
rect 55890 1700 55946 1748
rect 57570 1700 57626 1748
rect 59250 1700 59306 1748
rect 60930 1700 60986 1748
rect 62610 1700 62666 1748
rect 64290 1700 64346 1748
rect 65970 1700 66026 1748
rect 67650 1700 67706 1748
rect 69330 1700 69386 1748
rect 71010 1700 71066 1748
rect 72690 1700 72746 1748
rect 74370 1700 74426 1748
rect 76050 1700 76106 1748
rect 77730 1700 77786 1748
rect 79410 1700 79466 1748
rect 81090 1700 81146 1748
rect 82770 1700 82826 1748
rect 84450 1700 84506 1748
rect 86130 1700 86186 1748
rect 87810 1700 87866 1748
rect 89490 1700 89546 1748
rect 91170 1700 91226 1748
rect 92850 1700 92906 1748
rect 94530 1700 94586 1748
rect 96210 1700 96266 1748
rect 97890 1700 97946 1748
rect 99570 1700 99626 1748
rect 101250 1700 101306 1748
rect 102930 1700 102986 1748
rect 104610 1700 104666 1748
rect 106290 1700 106346 1748
rect 107970 1700 108026 1748
rect 109650 1700 109706 1748
rect 111330 1700 111386 1748
rect 113010 1700 113066 1748
rect 114690 1700 114746 1748
rect 116370 1700 116426 1748
rect 118050 1700 118106 1748
rect 119730 1700 119786 1748
rect 121410 1700 121466 1748
rect 123090 1700 123146 1748
rect 124770 1700 124826 1748
rect 126450 1700 126506 1748
rect 128130 1700 128186 1748
rect 129810 1700 129866 1748
rect 131490 1700 131546 1748
rect 133170 1700 133226 1748
rect 134760 1612 134984 81585
<< metal3 >>
rect 272 82688 136348 83036
rect 952 82008 135668 82356
rect 2040 81328 2252 81540
rect 3672 81328 4020 81540
rect 5440 81328 5652 81540
rect 7072 81328 7284 81540
rect 8704 81328 9052 81540
rect 10472 81328 10684 81540
rect 12104 81328 12316 81540
rect 13736 81328 14084 81540
rect 15504 81328 15716 81540
rect 17136 81328 17348 81540
rect 18904 81328 19116 81540
rect 20536 81328 20748 81540
rect 22168 81328 22380 81540
rect 23936 81328 24148 81540
rect 25568 81328 25780 81540
rect 27200 81328 27412 81540
rect 28968 81328 29180 81540
rect 30600 81328 30812 81540
rect 32232 81328 32580 81540
rect 34000 81328 34212 81540
rect 35632 81328 35844 81540
rect 37264 81328 37612 81540
rect 39032 81328 39244 81540
rect 40664 81328 40876 81540
rect 42296 81328 42644 81540
rect 44064 81328 44276 81540
rect 45696 81328 45908 81540
rect 47464 81328 47676 81540
rect 49096 81328 49308 81540
rect 50728 81328 50940 81540
rect 52496 81328 52708 81540
rect 54128 81328 54340 81540
rect 55760 81328 55972 81540
rect 57528 81328 57740 81540
rect 59160 81328 59372 81540
rect 60792 81328 61140 81540
rect 62560 81328 62772 81540
rect 64192 81328 64404 81540
rect 65824 81328 66172 81540
rect 67592 81328 67804 81540
rect 69224 81328 69436 81540
rect 70856 81328 71204 81540
rect 72624 81328 72836 81540
rect 74256 81328 74468 81540
rect 76024 81328 76236 81540
rect 77656 81328 77868 81540
rect 79288 81328 79500 81540
rect 81056 81464 81404 81540
rect 81056 81328 81268 81464
rect 82688 81328 82900 81540
rect 84320 81328 84532 81540
rect 86088 81328 86300 81540
rect 87720 81328 87932 81540
rect 89352 81328 89700 81540
rect 91120 81328 91332 81540
rect 92752 81328 92964 81540
rect 94384 81328 94732 81540
rect 96152 81328 96364 81540
rect 97784 81328 97996 81540
rect 99416 81328 99764 81540
rect 101184 81328 101396 81540
rect 102816 81328 103028 81540
rect 104584 81328 104796 81540
rect 106216 81328 106428 81540
rect 107848 81328 108060 81540
rect 109616 81328 109828 81540
rect 111248 81328 111460 81540
rect 112880 81328 113092 81540
rect 114648 81328 114860 81540
rect 116280 81328 116492 81540
rect 117912 81328 118260 81540
rect 119544 81464 119892 81540
rect 119680 81328 119892 81464
rect 121312 81328 121524 81540
rect 122944 81328 123292 81540
rect 124712 81328 124924 81540
rect 126344 81328 126556 81540
rect 127976 81328 128324 81540
rect 129744 81328 129956 81540
rect 131376 81328 131588 81540
rect 133144 81328 133356 81540
rect 1768 81056 2116 81132
rect 1768 80920 1980 81056
rect 134776 80996 134988 81132
rect 134776 80920 135396 80996
rect 118048 80724 118396 80860
rect 119272 80724 119484 80860
rect 117950 80648 122340 80724
rect 118796 80463 122216 80523
rect 118456 80104 118804 80316
rect 119680 80104 119892 80316
rect 122264 79696 122476 79908
rect 133960 79832 136076 79908
rect 133960 79696 134172 79832
rect 1224 79424 1980 79500
rect 1768 79288 1980 79424
rect 118048 79364 118396 79500
rect 119272 79364 119484 79500
rect 134776 79424 135396 79500
rect 118048 79288 119484 79364
rect 133824 79228 134036 79364
rect 134823 79291 134921 79424
rect 130696 79016 130908 79228
rect 133824 79152 136620 79228
rect 115328 78608 117988 78684
rect 115328 78472 115540 78608
rect 116416 78472 116628 78608
rect 122264 78472 123020 78548
rect 122264 78336 122476 78472
rect 133960 78412 134172 78548
rect 133960 78336 134852 78412
rect 1768 77596 1980 77732
rect 1224 77520 1980 77596
rect 134776 77656 135396 77732
rect 134776 77520 134988 77656
rect 115328 77248 118124 77324
rect 28560 76840 28772 77188
rect 28968 77087 29044 77188
rect 28851 76989 29044 77087
rect 28968 76976 29044 76989
rect 31008 76840 31220 77188
rect 31280 76976 31492 77188
rect 33456 77068 33668 77188
rect 33864 77087 34076 77188
rect 33456 76916 33687 77068
rect 33843 76989 34076 77087
rect 34000 76976 34076 76989
rect 33456 76840 33804 76916
rect 36040 76840 36252 77188
rect 36448 77087 36524 77188
rect 36339 76989 36524 77087
rect 36448 76976 36524 76989
rect 38488 76840 38700 77188
rect 38896 77087 38972 77188
rect 38835 77052 38972 77087
rect 41072 77068 41148 77188
rect 41344 77087 41556 77188
rect 38835 76989 39108 77052
rect 38896 76976 39108 76989
rect 41072 76916 41175 77068
rect 41331 76989 41556 77087
rect 41344 76976 41556 76989
rect 41072 76840 41284 76916
rect 43520 76840 43732 77188
rect 43928 77087 44004 77188
rect 43827 76989 44004 77087
rect 43928 76976 44004 76989
rect 45968 76840 46180 77188
rect 46376 77087 46452 77188
rect 46323 77052 46452 77087
rect 48552 77068 48628 77188
rect 48824 77087 49036 77188
rect 46323 76989 46588 77052
rect 46376 76976 46588 76989
rect 48552 76916 48663 77068
rect 48819 76989 49036 77087
rect 48960 76976 49036 76989
rect 48552 76840 48764 76916
rect 51000 76840 51212 77188
rect 51408 77087 51484 77188
rect 51315 76989 51484 77087
rect 51408 76976 51484 76989
rect 53448 76840 53660 77188
rect 53856 77087 53932 77188
rect 53811 76989 53932 77087
rect 53856 76976 53932 76989
rect 56032 76840 56244 77188
rect 56304 76976 56516 77188
rect 58480 76840 58692 77188
rect 58888 77087 58964 77188
rect 58803 76989 58964 77087
rect 58888 76976 58964 76989
rect 60928 77068 61140 77188
rect 61336 77150 61548 77188
rect 61299 77112 61548 77150
rect 60928 76916 61143 77068
rect 61299 76989 61397 77112
rect 60928 76840 61276 76916
rect 63512 76840 63724 77188
rect 63920 77087 63996 77188
rect 63795 76989 63996 77087
rect 63920 76976 63996 76989
rect 65960 76840 66172 77188
rect 66368 77087 66444 77188
rect 66291 77052 66444 77087
rect 68408 77068 68620 77188
rect 68816 77150 69028 77188
rect 68787 77112 69028 77150
rect 66291 76989 66580 77052
rect 66368 76976 66580 76989
rect 68408 76916 68631 77068
rect 68787 76989 68885 77112
rect 68408 76840 68756 76916
rect 70992 76840 71204 77188
rect 71400 77087 71476 77188
rect 71283 76989 71476 77087
rect 71400 76976 71476 76989
rect 73440 76840 73652 77188
rect 73848 77087 73924 77188
rect 73779 76989 73924 77087
rect 73848 76976 73924 76989
rect 75888 77068 76100 77188
rect 76296 77087 76508 77188
rect 75888 76916 76119 77068
rect 76275 76989 76508 77087
rect 76432 76976 76508 76989
rect 75888 76840 76236 76916
rect 78472 76840 78684 77188
rect 78880 77087 78956 77188
rect 78771 76989 78956 77087
rect 78880 76976 78956 76989
rect 80920 76840 81132 77188
rect 81328 77087 81404 77188
rect 81267 77052 81404 77087
rect 83504 77068 83580 77188
rect 83776 77087 83988 77188
rect 81267 76989 81540 77052
rect 81328 76976 81540 76989
rect 83504 76916 83607 77068
rect 83763 76989 83988 77087
rect 83912 76976 83988 76989
rect 83504 76840 83716 76916
rect 85952 76840 86164 77188
rect 86360 77087 86436 77188
rect 86259 76989 86436 77087
rect 86360 76976 86436 76989
rect 88400 76840 88612 77188
rect 88808 77087 88884 77188
rect 88755 77052 88884 77087
rect 90984 77068 91060 77188
rect 91256 77087 91468 77188
rect 88755 76989 89020 77052
rect 88808 76976 89020 76989
rect 90984 76916 91095 77068
rect 91251 76989 91468 77087
rect 91392 76976 91468 76989
rect 90984 76840 91196 76916
rect 93432 76840 93644 77188
rect 93840 77087 93916 77188
rect 93747 76989 93916 77087
rect 93840 76976 93916 76989
rect 95880 76840 96092 77188
rect 96288 77087 96364 77188
rect 96243 76989 96364 77087
rect 96288 76976 96364 76989
rect 98464 76840 98676 77188
rect 98872 77087 98948 77188
rect 98739 76989 98948 77087
rect 98872 76976 98948 76989
rect 100912 76840 101124 77188
rect 101320 77087 101396 77188
rect 101235 76989 101396 77087
rect 101320 76976 101396 76989
rect 103360 77068 103572 77188
rect 103768 77150 103980 77188
rect 103731 77112 103980 77150
rect 103360 76916 103575 77068
rect 103731 76989 103829 77112
rect 103360 76840 103708 76916
rect 105944 76840 106156 77188
rect 106352 77087 106428 77188
rect 115328 77112 115540 77248
rect 116416 77112 116628 77248
rect 106227 76989 106428 77087
rect 106352 76976 106428 76989
rect 122264 76840 122476 77052
rect 28832 76568 29044 76780
rect 31280 76704 36524 76780
rect 31280 76568 31492 76704
rect 33728 76568 34076 76704
rect 36312 76644 36524 76704
rect 36312 76568 38700 76644
rect 38760 76568 38972 76780
rect 41208 76644 41556 76780
rect 41208 76568 43732 76644
rect 43792 76568 44004 76780
rect 46240 76568 46452 76780
rect 48688 76704 51484 76780
rect 48688 76568 49036 76704
rect 51272 76568 51484 76704
rect 53720 76644 53932 76780
rect 56304 76704 61412 76780
rect 53720 76568 56244 76644
rect 56304 76568 56516 76704
rect 58752 76568 58964 76704
rect 61200 76568 61412 76704
rect 63784 76568 63996 76780
rect 66232 76568 66444 76780
rect 68680 76568 68892 76780
rect 71264 76644 71476 76780
rect 71166 76568 71476 76644
rect 73712 76704 76508 76780
rect 73712 76568 73924 76704
rect 76160 76644 76508 76704
rect 78744 76644 78956 76780
rect 81192 76644 81404 76780
rect 76160 76568 78684 76644
rect 78744 76568 81404 76644
rect 83640 76644 83988 76780
rect 86224 76644 86436 76780
rect 88672 76644 88884 76780
rect 83640 76568 86436 76644
rect 88574 76568 88884 76644
rect 91120 76644 91468 76780
rect 91120 76568 93644 76644
rect 93704 76568 93916 76780
rect 96152 76644 96364 76780
rect 98736 76704 103844 76780
rect 96152 76568 98676 76644
rect 98736 76568 98948 76704
rect 101184 76568 101396 76704
rect 103632 76568 103844 76704
rect 106216 76568 106428 76780
rect 1224 76024 1980 76100
rect 1768 75888 1980 76024
rect 134776 76024 135396 76100
rect 28832 75888 31492 75964
rect 28832 75752 29044 75888
rect 31280 75752 31492 75888
rect 33728 75752 33940 75964
rect 36312 75752 36524 75964
rect 38662 75888 38972 75964
rect 38760 75828 38972 75888
rect 41208 75828 41420 75964
rect 43694 75888 49036 75964
rect 38760 75752 41420 75828
rect 43792 75752 44004 75888
rect 46240 75752 46452 75888
rect 48688 75752 49036 75888
rect 51272 75828 51484 75964
rect 53720 75828 53932 75964
rect 51272 75752 53932 75828
rect 56168 75752 56516 75964
rect 58752 75828 58964 75964
rect 61200 75888 66444 75964
rect 58752 75752 59508 75828
rect 61200 75752 61412 75888
rect 63648 75752 63996 75888
rect 66232 75828 66444 75888
rect 68680 75888 71204 75964
rect 71264 75888 73924 75964
rect 68680 75828 68892 75888
rect 66232 75752 68892 75828
rect 71264 75752 71476 75888
rect 73712 75752 73924 75888
rect 76160 75752 76372 75964
rect 78646 75888 78956 75964
rect 78744 75752 78956 75888
rect 81192 75828 81404 75964
rect 83640 75828 83852 75964
rect 81192 75752 83852 75828
rect 86224 75888 88612 75964
rect 88672 75888 91468 75964
rect 93606 75888 93916 75964
rect 86224 75752 86436 75888
rect 88672 75752 88884 75888
rect 91120 75752 91468 75888
rect 93704 75828 93916 75888
rect 96152 75828 96364 75964
rect 93704 75752 96364 75828
rect 98600 75752 98948 75964
rect 101184 75752 101396 75964
rect 103632 75888 106428 75964
rect 103632 75752 103844 75888
rect 106080 75752 106428 75888
rect 115328 75692 115540 75964
rect 116416 75692 116628 75964
rect 134776 75888 134988 76024
rect 115328 75616 116628 75692
rect 122264 75480 122476 75692
rect 28832 75072 29044 75284
rect 31416 75072 31628 75284
rect 33864 75072 34076 75284
rect 36312 75072 36524 75284
rect 38896 75072 39108 75284
rect 41344 75072 41556 75284
rect 43792 75148 44004 75284
rect 43792 75072 44140 75148
rect 46376 75072 46588 75284
rect 48824 75072 49036 75284
rect 51272 75148 51484 75284
rect 51272 75072 51620 75148
rect 53856 75072 54068 75284
rect 56304 75072 56516 75284
rect 58752 75072 59100 75284
rect 61336 75072 61548 75284
rect 63784 75072 63996 75284
rect 66232 75072 66580 75284
rect 68816 75072 69028 75284
rect 71264 75072 71476 75284
rect 73848 75072 74060 75284
rect 76296 75072 76508 75284
rect 78744 75072 78956 75284
rect 81328 75072 81540 75284
rect 83776 75072 83988 75284
rect 86224 75148 86436 75284
rect 86224 75072 86572 75148
rect 88808 75072 89020 75284
rect 91256 75072 91468 75284
rect 93704 75072 93916 75284
rect 96288 75072 96500 75284
rect 98736 75072 98948 75284
rect 101184 75072 101532 75284
rect 103768 75072 103980 75284
rect 106216 75072 106428 75284
rect 28921 75055 29019 75072
rect 31417 75055 31515 75072
rect 33913 75055 34011 75072
rect 36409 75055 36507 75072
rect 38905 75055 39003 75072
rect 41401 75055 41499 75072
rect 43897 75055 43995 75072
rect 46393 75055 46491 75072
rect 48889 75055 48987 75072
rect 51385 75055 51483 75072
rect 53881 75055 53979 75072
rect 56377 75055 56475 75072
rect 58873 75055 58971 75072
rect 61369 75055 61467 75072
rect 63865 75055 63963 75072
rect 66361 75055 66459 75072
rect 68857 75055 68955 75072
rect 71353 75055 71451 75072
rect 73849 75055 73947 75072
rect 76345 75055 76443 75072
rect 78841 75055 78939 75072
rect 81337 75055 81435 75072
rect 83833 75055 83931 75072
rect 86329 75055 86427 75072
rect 88825 75055 88923 75072
rect 91321 75055 91419 75072
rect 93817 75055 93915 75072
rect 96313 75055 96411 75072
rect 98809 75055 98907 75072
rect 101305 75055 101403 75072
rect 103801 75055 103899 75072
rect 106297 75055 106395 75072
rect 110056 74888 110122 74919
rect 110089 74825 122300 74885
rect 1768 74196 1980 74468
rect 115328 74392 116628 74468
rect 115328 74256 115540 74392
rect 116416 74256 116628 74392
rect 1224 74120 1980 74196
rect 122264 73984 122476 74332
rect 132600 74060 132812 74332
rect 133280 74196 133492 74332
rect 134776 74196 134988 74468
rect 133280 74120 135396 74196
rect 133280 74060 133492 74120
rect 132600 73984 133492 74060
rect 110213 73411 122300 73471
rect 28968 73108 29316 73244
rect 30328 73108 30540 73244
rect 31552 73168 32988 73244
rect 31552 73108 31764 73168
rect 28968 73032 31764 73108
rect 32776 73108 32988 73168
rect 34000 73168 35436 73244
rect 34000 73108 34212 73168
rect 32776 73032 34212 73108
rect 35224 73108 35436 73168
rect 36448 73168 39244 73244
rect 36448 73108 36796 73168
rect 35224 73032 36796 73108
rect 37808 73032 38020 73168
rect 39032 73108 39244 73168
rect 40256 73168 41692 73244
rect 40256 73108 40468 73168
rect 39032 73032 40468 73108
rect 41480 73108 41692 73168
rect 42704 73168 45500 73244
rect 42704 73108 43052 73168
rect 41480 73032 43052 73108
rect 44064 73032 44276 73168
rect 45288 73108 45500 73168
rect 46512 73168 47948 73244
rect 46512 73108 46724 73168
rect 45288 73032 46724 73108
rect 47736 73108 47948 73168
rect 48960 73168 51756 73244
rect 48960 73108 49172 73168
rect 47736 73032 49172 73108
rect 50184 73032 50532 73168
rect 51544 73108 51756 73168
rect 52768 73168 54204 73244
rect 52768 73108 52980 73168
rect 51544 73032 52980 73108
rect 53992 73108 54204 73168
rect 55216 73168 56380 73244
rect 55216 73108 55428 73168
rect 56440 73108 56652 73244
rect 57664 73168 60460 73244
rect 57664 73108 58012 73168
rect 53992 73032 58012 73108
rect 59024 73032 59236 73168
rect 60248 73108 60460 73168
rect 61472 73168 62908 73244
rect 61472 73108 61684 73168
rect 60248 73032 61684 73108
rect 62696 73108 62908 73168
rect 63920 73168 66716 73244
rect 63920 73108 64268 73168
rect 62696 73032 64268 73108
rect 65280 73032 65492 73168
rect 66504 73108 66716 73168
rect 67728 73168 69164 73244
rect 67728 73108 67940 73168
rect 66504 73032 67940 73108
rect 68952 73108 69164 73168
rect 70176 73168 71748 73244
rect 70176 73108 70388 73168
rect 68952 73032 70388 73108
rect 71400 73108 71748 73168
rect 72760 73108 72972 73244
rect 73984 73168 75420 73244
rect 73984 73108 74196 73168
rect 71400 73032 74196 73108
rect 75208 73108 75420 73168
rect 76432 73168 77868 73244
rect 76432 73108 76644 73168
rect 75208 73032 76644 73108
rect 77656 73108 77868 73168
rect 78880 73168 81676 73244
rect 78880 73108 79228 73168
rect 77656 73032 79228 73108
rect 80240 73032 80452 73168
rect 81464 73108 81676 73168
rect 82688 73168 84124 73244
rect 82688 73108 82900 73168
rect 81464 73032 82900 73108
rect 83912 73108 84124 73168
rect 85136 73168 87932 73244
rect 85136 73108 85484 73168
rect 83912 73032 85484 73108
rect 86496 73032 86708 73168
rect 87720 73108 87932 73168
rect 88944 73168 90380 73244
rect 88944 73108 89156 73168
rect 87720 73032 89156 73108
rect 90168 73108 90380 73168
rect 91392 73168 93780 73244
rect 91392 73108 91604 73168
rect 90168 73032 91604 73108
rect 92616 73108 92964 73168
rect 93976 73108 94188 73244
rect 95200 73168 96636 73244
rect 95200 73108 95412 73168
rect 92616 73032 95412 73108
rect 96424 73108 96636 73168
rect 97648 73168 99084 73244
rect 97648 73108 97860 73168
rect 96424 73032 97860 73108
rect 98872 73108 99084 73168
rect 100096 73108 100444 73244
rect 101456 73168 102892 73244
rect 101456 73108 101668 73168
rect 98872 73032 101668 73108
rect 102680 73108 102892 73168
rect 103904 73168 105340 73244
rect 103904 73108 104116 73168
rect 102680 73032 104116 73108
rect 105128 73108 105340 73168
rect 106352 73168 107924 73244
rect 106352 73108 106700 73168
rect 105128 73032 106700 73108
rect 107712 73108 107924 73168
rect 107712 73032 109692 73108
rect 115328 73032 116628 73108
rect 115328 72972 115540 73032
rect 115328 72896 115948 72972
rect 116416 72896 116628 73032
rect 1224 72624 1980 72700
rect 122264 72624 122476 72836
rect 132600 72760 136076 72836
rect 132600 72624 132812 72760
rect 133280 72624 133492 72760
rect 1768 72488 1980 72624
rect 134776 72564 134988 72700
rect 134776 72488 135396 72564
rect 115272 72296 115332 72356
rect 122132 72296 134125 72356
rect 114074 71997 122300 72057
rect 28560 71400 28772 71612
rect 29512 71476 29724 71612
rect 29784 71476 30132 71612
rect 29512 71400 30132 71476
rect 30736 71536 31356 71612
rect 30736 71400 30948 71536
rect 31144 71400 31356 71536
rect 31960 71476 32172 71612
rect 32368 71476 32580 71612
rect 31960 71400 32580 71476
rect 33184 71536 33804 71612
rect 33184 71400 33396 71536
rect 33592 71400 33804 71536
rect 34408 71476 34620 71612
rect 34816 71476 35028 71612
rect 34408 71400 35028 71476
rect 35632 71476 35980 71612
rect 36040 71476 36252 71612
rect 35632 71400 36252 71476
rect 36992 71536 37612 71612
rect 36992 71400 37204 71536
rect 37264 71400 37612 71536
rect 38216 71476 38428 71612
rect 38624 71476 38836 71612
rect 38216 71400 38836 71476
rect 39440 71536 40060 71612
rect 39440 71400 39652 71536
rect 39848 71400 40060 71536
rect 40664 71476 40876 71612
rect 41072 71476 41284 71612
rect 40664 71400 41284 71476
rect 41888 71536 42508 71612
rect 41888 71400 42236 71536
rect 42296 71400 42508 71536
rect 43248 71536 43868 71612
rect 43248 71400 43460 71536
rect 43520 71400 43868 71536
rect 44472 71476 44684 71612
rect 44880 71536 46316 71612
rect 44880 71476 45092 71536
rect 44472 71400 45092 71476
rect 45696 71400 45908 71536
rect 46104 71400 46316 71536
rect 46920 71476 47132 71612
rect 47328 71476 47540 71612
rect 46920 71400 47540 71476
rect 48144 71536 48764 71612
rect 48144 71400 48356 71536
rect 48552 71400 48764 71536
rect 49368 71536 49988 71612
rect 49368 71400 49716 71536
rect 49776 71400 49988 71536
rect 50728 71476 50940 71612
rect 51000 71476 51348 71612
rect 50728 71400 51348 71476
rect 51952 71536 52572 71612
rect 51952 71400 52164 71536
rect 52360 71400 52572 71536
rect 53176 71476 53388 71612
rect 53584 71476 53796 71612
rect 53176 71400 53796 71476
rect 54400 71536 55020 71612
rect 54400 71400 54612 71536
rect 54808 71400 55020 71536
rect 55624 71476 55836 71612
rect 56032 71476 56244 71612
rect 55624 71400 56244 71476
rect 56848 71536 57468 71612
rect 56848 71400 57196 71536
rect 57256 71400 57468 71536
rect 58208 71536 58828 71612
rect 58208 71400 58420 71536
rect 58480 71400 58828 71536
rect 59432 71476 59644 71612
rect 59840 71476 60052 71612
rect 59432 71400 60052 71476
rect 60656 71536 61276 71612
rect 60656 71400 60868 71536
rect 61064 71400 61276 71536
rect 61880 71476 62092 71612
rect 62288 71476 62500 71612
rect 61880 71400 62500 71476
rect 63104 71536 63724 71612
rect 63104 71400 63452 71536
rect 63512 71400 63724 71536
rect 64464 71536 65084 71612
rect 64464 71400 64676 71536
rect 64736 71400 65084 71536
rect 65688 71476 65900 71612
rect 66096 71476 66308 71612
rect 65688 71400 66308 71476
rect 66912 71536 67532 71612
rect 66912 71400 67124 71536
rect 67320 71400 67532 71536
rect 68136 71476 68348 71612
rect 68544 71476 68756 71612
rect 68136 71400 68756 71476
rect 69360 71536 69980 71612
rect 69360 71400 69572 71536
rect 69768 71400 69980 71536
rect 70584 71476 70932 71612
rect 70992 71476 71204 71612
rect 70584 71400 71204 71476
rect 71944 71476 72156 71612
rect 72216 71476 72564 71612
rect 71944 71400 72564 71476
rect 73168 71536 73788 71612
rect 73168 71400 73380 71536
rect 73576 71400 73788 71536
rect 74392 71476 74604 71612
rect 74800 71476 75012 71612
rect 74392 71400 75012 71476
rect 75616 71536 76236 71612
rect 75616 71400 75828 71536
rect 76024 71400 76236 71536
rect 76840 71476 77052 71612
rect 77248 71476 77460 71612
rect 76840 71400 77460 71476
rect 78064 71400 78412 71612
rect 78472 71400 78684 71612
rect 79424 71536 80044 71612
rect 79424 71400 79636 71536
rect 79696 71400 80044 71536
rect 80648 71476 80860 71612
rect 81056 71476 81268 71612
rect 80648 71400 81268 71476
rect 81872 71536 82492 71612
rect 81872 71400 82084 71536
rect 82280 71400 82492 71536
rect 83096 71476 83308 71612
rect 83504 71476 83716 71612
rect 83096 71400 83716 71476
rect 84320 71536 84940 71612
rect 84320 71400 84668 71536
rect 84728 71400 84940 71536
rect 85680 71536 86300 71612
rect 85680 71400 85892 71536
rect 85952 71400 86300 71536
rect 86904 71476 87116 71612
rect 87312 71476 87524 71612
rect 86904 71400 87524 71476
rect 88128 71536 88748 71612
rect 88128 71400 88340 71536
rect 88536 71400 88748 71536
rect 89352 71476 89564 71612
rect 89760 71476 89972 71612
rect 89352 71400 89972 71476
rect 90576 71536 91196 71612
rect 90576 71400 90788 71536
rect 90984 71400 91196 71536
rect 91800 71476 92148 71612
rect 92208 71476 92420 71612
rect 91800 71400 92420 71476
rect 93160 71476 93372 71612
rect 93432 71476 93780 71612
rect 93160 71400 93780 71476
rect 94384 71536 95004 71612
rect 94384 71400 94596 71536
rect 94792 71400 95004 71536
rect 95608 71476 95820 71612
rect 96016 71476 96228 71612
rect 95608 71400 96228 71476
rect 96832 71536 97452 71612
rect 96832 71400 97044 71536
rect 97240 71400 97452 71536
rect 98056 71476 98268 71612
rect 98464 71476 98676 71612
rect 98056 71400 98676 71476
rect 99280 71536 99900 71612
rect 99280 71400 99628 71536
rect 99688 71400 99900 71536
rect 100640 71536 101260 71612
rect 100640 71400 100852 71536
rect 100912 71400 101260 71536
rect 101864 71476 102076 71612
rect 102272 71476 102484 71612
rect 101864 71400 102484 71476
rect 103088 71536 103708 71612
rect 103088 71400 103300 71536
rect 103496 71400 103708 71536
rect 104312 71476 104524 71612
rect 104720 71476 104932 71612
rect 104312 71400 104932 71476
rect 105536 71536 106156 71612
rect 105536 71400 105884 71536
rect 105944 71400 106156 71536
rect 106896 71536 107516 71612
rect 106896 71400 107108 71536
rect 107168 71400 107516 71536
rect 108120 71476 108332 71612
rect 108528 71476 108740 71612
rect 108120 71400 108740 71476
rect 98192 71340 98268 71400
rect 98192 71264 98676 71340
rect 122264 71264 122476 71476
rect 132600 71340 132812 71476
rect 133280 71340 133492 71476
rect 132600 71264 134852 71340
rect 1224 70992 1980 71068
rect 1768 70856 1980 70992
rect 28152 70992 28636 71068
rect 27064 70796 27276 70932
rect 28152 70856 28364 70992
rect 28696 70932 28908 71068
rect 29376 70992 29860 71068
rect 29920 70992 30812 71068
rect 29376 70932 29588 70992
rect 29920 70932 30132 70992
rect 28696 70856 30132 70932
rect 30600 70932 30812 70992
rect 31144 70932 31492 71068
rect 31824 70932 32036 71068
rect 30600 70856 32036 70932
rect 32504 70932 32716 71068
rect 33048 70932 33260 71068
rect 33728 70992 34620 71068
rect 33728 70932 33940 70992
rect 32504 70856 33940 70932
rect 34272 70856 34620 70992
rect 34952 70932 35164 71068
rect 35632 70932 35844 71068
rect 34952 70856 35844 70932
rect 36176 70992 37068 71068
rect 36176 70856 36388 70992
rect 36856 70856 37068 70992
rect 37400 70932 37748 71068
rect 38080 70992 38972 71068
rect 38080 70932 38292 70992
rect 37400 70856 38292 70932
rect 38760 70932 38972 70992
rect 39304 70932 39516 71068
rect 39984 70992 40740 71068
rect 39984 70932 40196 70992
rect 38760 70856 40196 70932
rect 40528 70856 40740 70992
rect 41208 70932 41420 71068
rect 41752 70932 42100 71068
rect 41208 70856 42100 70932
rect 42432 70992 43324 71068
rect 42432 70856 42644 70992
rect 43112 70932 43324 70992
rect 43656 70932 43868 71068
rect 44336 70992 45228 71068
rect 44336 70932 44548 70992
rect 44880 70932 45228 70992
rect 43112 70856 44548 70932
rect 44646 70856 45228 70932
rect 45560 70856 45772 71068
rect 46240 70992 47676 71068
rect 46240 70856 46452 70992
rect 46784 70856 46996 70992
rect 47464 70932 47676 70992
rect 48008 70992 49580 71068
rect 48008 70932 48356 70992
rect 47464 70856 48356 70932
rect 48688 70856 48900 70992
rect 49368 70932 49580 70992
rect 49912 70932 50124 71068
rect 50592 70932 50804 71068
rect 49368 70856 50804 70932
rect 51136 70992 52028 71068
rect 51136 70856 51348 70992
rect 51816 70932 52028 70992
rect 52360 70992 53252 71068
rect 53350 70992 53932 71068
rect 52360 70932 52708 70992
rect 51816 70856 52708 70932
rect 53040 70856 53252 70992
rect 53720 70932 53932 70992
rect 54264 70932 54476 71068
rect 53720 70856 54476 70932
rect 54944 70992 56108 71068
rect 54944 70856 55156 70992
rect 55488 70932 55836 70992
rect 56168 70932 56380 71068
rect 56848 70992 58284 71068
rect 56848 70932 57060 70992
rect 55488 70856 57060 70932
rect 57392 70856 57604 70992
rect 58072 70932 58284 70992
rect 58616 70932 58964 71068
rect 59296 70932 59508 71068
rect 58072 70856 59508 70932
rect 59976 70932 60188 71068
rect 60520 70932 60732 71068
rect 61200 70992 61956 71068
rect 61200 70932 61412 70992
rect 59976 70856 61412 70932
rect 61744 70856 61956 70992
rect 62424 70932 62636 71068
rect 62968 70932 63316 71068
rect 62424 70856 63316 70932
rect 63648 70992 64540 71068
rect 63648 70856 63860 70992
rect 64328 70932 64540 70992
rect 64872 70932 65084 71068
rect 65552 70992 66988 71068
rect 65552 70932 65764 70992
rect 64328 70856 65764 70932
rect 66096 70856 66444 70992
rect 66776 70856 66988 70992
rect 67456 70992 68212 71068
rect 67456 70856 67668 70992
rect 68000 70856 68212 70992
rect 68680 70932 68892 71068
rect 69224 70932 69572 71068
rect 69904 70992 70796 71068
rect 69904 70932 70116 70992
rect 68680 70856 70116 70932
rect 70584 70932 70796 70992
rect 71128 70932 71340 71068
rect 71808 70992 72292 71068
rect 72352 70992 73244 71068
rect 71808 70932 72020 70992
rect 72352 70932 72564 70992
rect 70584 70856 72020 70932
rect 72118 70856 72564 70932
rect 73032 70932 73244 70992
rect 73576 70932 73924 71068
rect 74256 70932 74468 71068
rect 73032 70856 74468 70932
rect 74936 70932 75148 71068
rect 75480 70932 75692 71068
rect 74936 70856 75692 70932
rect 76160 70992 77052 71068
rect 76160 70856 76372 70992
rect 76704 70856 77052 70992
rect 77384 70932 77596 71068
rect 78064 70992 78548 71068
rect 78608 70992 79500 71068
rect 78064 70932 78276 70992
rect 78608 70932 78820 70992
rect 77384 70856 78820 70932
rect 79288 70856 79500 70992
rect 79832 70932 80180 71068
rect 80512 70992 81404 71068
rect 80512 70932 80724 70992
rect 79832 70856 80724 70932
rect 81192 70932 81404 70992
rect 81736 70932 81948 71068
rect 81192 70856 81948 70932
rect 82416 70992 83172 71068
rect 82416 70856 82628 70992
rect 82960 70856 83172 70992
rect 83640 70932 83852 71068
rect 84184 70932 84532 71068
rect 84630 70992 85756 71068
rect 84864 70932 85076 70992
rect 83640 70856 85076 70932
rect 85544 70932 85756 70992
rect 86088 70932 86300 71068
rect 86768 70992 88204 71068
rect 86768 70932 86980 70992
rect 85544 70856 86980 70932
rect 87312 70856 87660 70992
rect 87992 70856 88204 70992
rect 88672 70992 89428 71068
rect 88672 70856 88884 70992
rect 89216 70856 89428 70992
rect 89896 70932 90108 71068
rect 90440 70932 90788 71068
rect 89896 70856 90788 70932
rect 91120 70992 92012 71068
rect 91120 70856 91332 70992
rect 91800 70932 92012 70992
rect 92344 70932 92556 71068
rect 93024 70992 94460 71068
rect 93024 70932 93236 70992
rect 93568 70932 93780 70992
rect 91800 70856 93236 70932
rect 93334 70856 93780 70932
rect 94248 70932 94460 70992
rect 94792 70932 95140 71068
rect 95472 70992 96364 71068
rect 95472 70932 95684 70992
rect 94248 70856 95684 70932
rect 96152 70932 96364 70992
rect 96696 70932 96908 71068
rect 96152 70856 96908 70932
rect 97376 70992 98268 71068
rect 97376 70856 97588 70992
rect 97920 70932 98268 70992
rect 98600 70932 98812 71068
rect 99280 70992 100988 71068
rect 99280 70932 99492 70992
rect 97920 70856 99492 70932
rect 99824 70856 100036 70992
rect 100504 70932 100716 70992
rect 101048 70932 101396 71068
rect 101728 70932 101940 71068
rect 100504 70856 101940 70932
rect 102408 70932 102620 71068
rect 102952 70932 103164 71068
rect 102408 70856 103164 70932
rect 103632 70992 104388 71068
rect 103632 70856 103844 70992
rect 104176 70856 104388 70992
rect 104856 70932 105068 71068
rect 105400 70932 105748 71068
rect 104856 70856 105748 70932
rect 106080 70992 106972 71068
rect 106080 70856 106292 70992
rect 106760 70932 106972 70992
rect 107304 70932 107516 71068
rect 107984 70992 110780 71068
rect 107984 70932 108196 70992
rect 106760 70856 108196 70932
rect 108528 70856 108876 70992
rect 134776 70932 134988 71068
rect 27064 70720 29044 70796
rect 27064 70660 27276 70720
rect 27064 70584 27412 70660
rect 27336 70524 27412 70584
rect 109616 70584 109828 70932
rect 134776 70856 135396 70932
rect 109616 70524 109692 70584
rect 27336 70312 27684 70524
rect 109344 70448 109692 70524
rect 110704 70524 110916 70660
rect 113424 70524 113636 70660
rect 114240 70584 115404 70660
rect 114240 70524 114452 70584
rect 110704 70448 114452 70524
rect 109344 70312 109556 70448
rect 27336 70252 27412 70312
rect 109480 70252 109556 70312
rect 20808 69904 21020 70116
rect 21216 70040 21972 70116
rect 21216 69904 21428 70040
rect 21624 69904 21972 70040
rect 22032 69904 22244 70116
rect 22440 69904 22652 70116
rect 27336 70040 27684 70252
rect 27608 69980 27684 70040
rect 20944 69844 21020 69904
rect 21624 69844 21700 69904
rect 20808 69496 21020 69844
rect 21352 69768 21700 69844
rect 27336 69768 27684 69980
rect 109344 70040 109556 70252
rect 109344 69980 109420 70040
rect 109344 69768 109556 69980
rect 114240 69904 114452 70116
rect 114648 69904 114860 70116
rect 115056 69980 115268 70116
rect 115056 69904 115404 69980
rect 115464 69904 115676 70116
rect 115872 69904 116084 70116
rect 132600 69904 133492 69980
rect 115872 69844 115948 69904
rect 21352 69708 21428 69768
rect 27472 69708 27548 69768
rect 109344 69708 109420 69768
rect 21216 69632 21972 69708
rect 21216 69496 21428 69632
rect 21624 69496 21972 69632
rect 22032 69496 22244 69708
rect 22440 69496 22652 69708
rect 27336 69496 27684 69708
rect 109344 69496 109556 69708
rect 114240 69496 114452 69708
rect 114648 69496 114860 69708
rect 115056 69496 115268 69708
rect 115366 69632 115676 69708
rect 115464 69496 115676 69632
rect 115872 69496 116084 69844
rect 132600 69768 132812 69904
rect 133280 69844 133492 69904
rect 133182 69768 133492 69844
rect 27472 69436 27548 69496
rect 109480 69436 109556 69496
rect 1768 69300 1980 69436
rect 1224 69224 1980 69300
rect 1768 69088 1980 69224
rect 20808 69088 21020 69300
rect 21216 69088 21428 69300
rect 21624 69088 21972 69300
rect 22032 69088 22244 69300
rect 22440 69088 22652 69300
rect 27336 69224 27684 69436
rect 109344 69224 109556 69436
rect 134776 69360 135396 69436
rect 27472 69164 27548 69224
rect 109480 69164 109556 69224
rect 20808 69028 20884 69088
rect 20808 68816 21020 69028
rect 27336 68952 27684 69164
rect 109344 68952 109556 69164
rect 114240 69088 114452 69300
rect 114648 69088 114860 69300
rect 115056 69088 115268 69300
rect 115464 69088 115676 69300
rect 115872 69088 116084 69300
rect 134776 69088 134988 69360
rect 115464 69028 115540 69088
rect 115192 68952 115540 69028
rect 115872 69028 115948 69088
rect 27472 68892 27548 68952
rect 109344 68892 109420 68952
rect 115192 68892 115268 68952
rect 21216 68680 21428 68892
rect 21624 68756 21972 68892
rect 21488 68680 21972 68756
rect 22032 68680 22244 68892
rect 22440 68680 22652 68892
rect 21216 68620 21292 68680
rect 21488 68620 21564 68680
rect 20808 68272 21020 68620
rect 21216 68544 21564 68620
rect 21624 68620 21700 68680
rect 21216 68272 21428 68544
rect 21624 68272 21972 68620
rect 22032 68272 22244 68484
rect 22440 68272 22652 68484
rect 27336 68408 27684 68892
rect 109344 68408 109556 68892
rect 114240 68756 114452 68892
rect 114240 68680 114588 68756
rect 114648 68680 114860 68892
rect 115056 68816 115676 68892
rect 115872 68816 116084 69028
rect 115056 68680 115268 68816
rect 114512 68620 114588 68680
rect 115192 68620 115268 68680
rect 114512 68544 115268 68620
rect 27472 68348 27548 68408
rect 109480 68348 109556 68408
rect 20944 68212 21020 68272
rect 22168 68212 22244 68272
rect 22576 68212 22652 68272
rect 20808 68000 21020 68212
rect 21216 67864 21428 68076
rect 21624 67864 21972 68076
rect 21216 67804 21292 67864
rect 21896 67804 21972 67864
rect 1768 67532 1980 67668
rect 20808 67592 21020 67804
rect 21216 67592 21428 67804
rect 21624 67592 21972 67804
rect 22032 67864 22244 68212
rect 22440 67864 22652 68212
rect 22032 67804 22108 67864
rect 22440 67804 22516 67864
rect 1224 67456 1980 67532
rect 22032 67456 22244 67804
rect 22168 67396 22244 67456
rect 20808 67184 21020 67396
rect 21216 67260 21428 67396
rect 21216 67184 21564 67260
rect 21216 67124 21428 67184
rect 21624 67124 21972 67396
rect 22032 67184 22244 67396
rect 22440 67456 22652 67804
rect 27336 67728 27684 68348
rect 109344 67728 109556 68348
rect 114240 68272 114452 68484
rect 114648 68272 114860 68484
rect 115056 68272 115268 68544
rect 115464 68680 115676 68816
rect 115464 68620 115540 68680
rect 115464 68348 115676 68620
rect 115366 68272 115676 68348
rect 115872 68272 116084 68620
rect 132600 68484 132812 68620
rect 133280 68544 134852 68620
rect 133280 68484 133492 68544
rect 132600 68408 133492 68484
rect 114240 68212 114316 68272
rect 114648 68212 114724 68272
rect 116008 68212 116084 68272
rect 114240 67864 114452 68212
rect 114648 67864 114860 68212
rect 115056 68000 115404 68076
rect 115056 67864 115268 68000
rect 115464 67940 115676 68076
rect 115872 68000 116084 68212
rect 114376 67804 114452 67864
rect 114784 67804 114860 67864
rect 115192 67804 115268 67864
rect 115328 67864 115676 67940
rect 115328 67804 115404 67864
rect 27336 67668 27412 67728
rect 27336 67592 27684 67668
rect 109344 67592 109556 67668
rect 22440 67396 22516 67456
rect 27462 67396 27560 67592
rect 109344 67396 109448 67592
rect 114240 67456 114452 67804
rect 114648 67456 114860 67804
rect 115056 67728 115404 67804
rect 115056 67668 115268 67728
rect 115464 67668 115676 67804
rect 115056 67592 115676 67668
rect 115872 67592 116084 67804
rect 134776 67592 135396 67668
rect 134776 67456 134988 67592
rect 114240 67396 114316 67456
rect 114648 67396 114724 67456
rect 22440 67184 22652 67396
rect 27336 67184 27684 67396
rect 109344 67184 109556 67396
rect 114240 67184 114452 67396
rect 114648 67184 114860 67396
rect 27472 67124 27548 67184
rect 109480 67124 109556 67184
rect 21216 67048 21972 67124
rect 21352 66988 21428 67048
rect 20808 66776 21020 66988
rect 21216 66776 21428 66988
rect 21526 66912 21972 66988
rect 21624 66776 21972 66912
rect 22032 66776 22244 66988
rect 22440 66776 22652 66988
rect 27336 66912 27684 67124
rect 109344 66912 109556 67124
rect 115056 67048 115268 67396
rect 115464 67124 115676 67396
rect 115872 67184 116084 67396
rect 132600 67184 133492 67260
rect 115192 66988 115268 67048
rect 115328 67048 115676 67124
rect 132600 67124 132812 67184
rect 132600 67048 133220 67124
rect 115328 66988 115404 67048
rect 27336 66852 27412 66912
rect 109344 66852 109420 66912
rect 27336 66640 27684 66852
rect 109344 66640 109556 66852
rect 114240 66776 114452 66988
rect 114648 66776 114860 66988
rect 115056 66912 115404 66988
rect 115056 66852 115268 66912
rect 115464 66852 115676 66988
rect 115056 66776 115676 66852
rect 115872 66776 116084 66988
rect 132600 66912 132812 67048
rect 133280 66912 133492 67184
rect 27472 66580 27548 66640
rect 109344 66580 109420 66640
rect 20808 66368 21020 66580
rect 21216 66504 21972 66580
rect 21216 66444 21428 66504
rect 21216 66368 21564 66444
rect 21624 66368 21972 66504
rect 22032 66368 22244 66580
rect 22440 66368 22652 66580
rect 27336 66368 27684 66580
rect 109344 66368 109556 66580
rect 114240 66368 114452 66580
rect 114648 66368 114860 66580
rect 115056 66504 115676 66580
rect 115056 66444 115268 66504
rect 115056 66368 115404 66444
rect 115464 66368 115676 66504
rect 115872 66368 116084 66580
rect 27608 66308 27684 66368
rect 109480 66308 109556 66368
rect 1224 65960 1980 66036
rect 20808 65960 21020 66172
rect 21216 65960 21428 66172
rect 21526 66096 21972 66172
rect 21624 65960 21972 66096
rect 22032 65960 22244 66172
rect 22440 65960 22652 66172
rect 27336 66096 27684 66308
rect 109344 66096 109556 66308
rect 27608 66036 27684 66096
rect 109480 66036 109556 66096
rect 1768 65824 1980 65960
rect 27336 65824 27684 66036
rect 27608 65764 27684 65824
rect 20808 65552 21020 65764
rect 21216 65552 21428 65764
rect 21624 65628 21972 65764
rect 21526 65552 21972 65628
rect 22032 65552 22244 65764
rect 22440 65552 22652 65764
rect 27336 65552 27684 65764
rect 27608 65492 27684 65552
rect 20808 65144 21020 65356
rect 21216 65280 21564 65356
rect 21216 65220 21428 65280
rect 21624 65220 21972 65356
rect 21216 65144 21972 65220
rect 22032 65144 22244 65356
rect 22440 65144 22652 65356
rect 27336 65280 27684 65492
rect 109344 65824 109556 66036
rect 114240 65960 114452 66172
rect 114648 65960 114860 66172
rect 115056 65960 115268 66172
rect 115366 66096 115676 66172
rect 115464 65960 115676 66096
rect 115872 65960 116084 66172
rect 134776 65900 134988 66036
rect 134776 65824 135396 65900
rect 109344 65764 109420 65824
rect 134776 65764 134852 65824
rect 109344 65552 109556 65764
rect 114240 65552 114452 65764
rect 114648 65552 114860 65764
rect 115056 65688 115676 65764
rect 115056 65628 115268 65688
rect 115056 65552 115404 65628
rect 115464 65552 115676 65688
rect 115872 65552 116084 65764
rect 132600 65688 134852 65764
rect 132600 65552 132812 65688
rect 133280 65552 133492 65688
rect 109344 65492 109420 65552
rect 109344 65280 109556 65492
rect 27472 65220 27548 65280
rect 109480 65220 109556 65280
rect 20944 65084 21020 65144
rect 20808 65008 22108 65084
rect 27336 65008 27684 65220
rect 109344 65008 109556 65220
rect 114240 65144 114452 65356
rect 114648 65144 114860 65356
rect 115056 65144 115268 65356
rect 115366 65280 115676 65356
rect 115464 65144 115676 65280
rect 115872 65144 116084 65356
rect 20808 64736 21020 65008
rect 27608 64948 27684 65008
rect 109480 64948 109556 65008
rect 115872 65084 115948 65144
rect 21216 64736 21428 64948
rect 21624 64812 21972 64948
rect 21488 64736 21972 64812
rect 22032 64736 22244 64948
rect 22440 64736 22652 64948
rect 20808 64676 20884 64736
rect 21216 64676 21292 64736
rect 21488 64676 21564 64736
rect 1768 64132 1980 64404
rect 1224 64056 1980 64132
rect 20808 64328 21020 64676
rect 21216 64600 21564 64676
rect 21216 64404 21428 64600
rect 21624 64404 21972 64676
rect 21216 64328 21972 64404
rect 22032 64328 22244 64540
rect 22440 64328 22652 64540
rect 27336 64464 27684 64948
rect 109344 64464 109556 64948
rect 114240 64736 114452 64948
rect 114648 64736 114860 64948
rect 115056 64736 115268 64948
rect 115464 64736 115676 64948
rect 115600 64676 115676 64736
rect 115056 64600 115676 64676
rect 109344 64404 109420 64464
rect 20808 64268 20884 64328
rect 22032 64268 22108 64328
rect 22440 64268 22516 64328
rect 20808 64056 21020 64268
rect 21216 63996 21428 64132
rect 21216 63920 21564 63996
rect 21624 63920 21972 64132
rect 22032 63920 22244 64268
rect 21352 63860 21428 63920
rect 20808 63648 21020 63860
rect 21216 63648 21428 63860
rect 21488 63860 21564 63920
rect 21896 63860 21972 63920
rect 22168 63860 22244 63920
rect 21488 63784 21972 63860
rect 21624 63648 21972 63784
rect 22032 63512 22244 63860
rect 22440 63920 22652 64268
rect 22440 63860 22516 63920
rect 22440 63512 22652 63860
rect 27336 63784 27684 64404
rect 109344 63996 109556 64404
rect 114240 64328 114452 64540
rect 114376 64268 114452 64328
rect 109246 63920 109556 63996
rect 109344 63784 109556 63920
rect 114240 63920 114452 64268
rect 114648 64328 114860 64540
rect 115056 64404 115268 64600
rect 115056 64328 115404 64404
rect 115464 64328 115676 64600
rect 115872 64736 116084 65084
rect 115872 64676 115948 64736
rect 115872 64328 116084 64676
rect 134640 64464 136076 64540
rect 134640 64404 134716 64464
rect 114648 64268 114724 64328
rect 116008 64268 116084 64328
rect 114648 63920 114860 64268
rect 115056 63996 115268 64132
rect 115366 64056 115676 64132
rect 115872 64056 116084 64268
rect 132600 64268 132812 64404
rect 133280 64328 134716 64404
rect 133280 64268 133492 64328
rect 132600 64192 133492 64268
rect 134776 64132 134988 64404
rect 134776 64056 135396 64132
rect 115056 63920 115404 63996
rect 114240 63860 114316 63920
rect 114648 63860 114724 63920
rect 115056 63860 115132 63920
rect 115328 63860 115404 63920
rect 115464 63920 115676 64056
rect 115464 63860 115540 63920
rect 22032 63452 22108 63512
rect 22576 63452 22652 63512
rect 20808 63240 21020 63452
rect 21216 63316 21428 63452
rect 21624 63316 21972 63452
rect 21216 63240 21972 63316
rect 22032 63240 22244 63452
rect 22440 63240 22652 63452
rect 27336 63240 27684 63588
rect 109208 63512 109556 63588
rect 114240 63512 114452 63860
rect 114648 63512 114860 63860
rect 115056 63648 115268 63860
rect 115328 63784 115676 63860
rect 115464 63648 115676 63784
rect 115872 63648 116084 63860
rect 109344 63240 109556 63512
rect 114376 63452 114452 63512
rect 114784 63452 114860 63512
rect 114240 63240 114452 63452
rect 114648 63240 114860 63452
rect 21216 63180 21428 63240
rect 21216 63104 21564 63180
rect 21624 63104 21972 63240
rect 27608 63180 27684 63240
rect 109480 63180 109556 63240
rect 21352 63044 21428 63104
rect 20808 62832 21020 63044
rect 21216 62832 21428 63044
rect 21488 63044 21564 63104
rect 21488 62968 21972 63044
rect 21624 62832 21972 62968
rect 22032 62832 22244 63044
rect 22440 62832 22652 63044
rect 27336 62968 27684 63180
rect 109344 62968 109556 63180
rect 115056 63104 115268 63452
rect 115464 63104 115676 63452
rect 115872 63240 116084 63452
rect 115056 63044 115132 63104
rect 115464 63044 115540 63104
rect 27608 62908 27684 62968
rect 109480 62908 109556 62968
rect 1224 62560 1980 62636
rect 1768 62424 1980 62560
rect 20808 62424 21020 62636
rect 21216 62424 21428 62636
rect 21624 62424 21972 62636
rect 22032 62424 22244 62636
rect 22440 62424 22652 62636
rect 27336 62424 27684 62908
rect 109344 62424 109556 62908
rect 114240 62832 114452 63044
rect 114648 62832 114860 63044
rect 115056 62832 115268 63044
rect 115464 62832 115676 63044
rect 115872 62832 116084 63044
rect 132600 62772 132812 62908
rect 133280 62772 133492 62908
rect 132600 62696 134852 62772
rect 134776 62636 134852 62696
rect 114240 62424 114452 62636
rect 114648 62424 114860 62636
rect 115056 62424 115268 62636
rect 115464 62424 115676 62636
rect 115872 62424 116084 62636
rect 134776 62500 134988 62636
rect 134776 62424 135396 62500
rect 27472 62364 27548 62424
rect 109344 62364 109420 62424
rect 115464 62364 115540 62424
rect 20808 62016 21020 62228
rect 21216 62016 21428 62228
rect 21624 62016 21972 62228
rect 22032 62016 22244 62228
rect 22440 62016 22652 62228
rect 27336 62152 27684 62364
rect 109344 62152 109556 62364
rect 115192 62288 115540 62364
rect 115192 62228 115268 62288
rect 27336 62092 27412 62152
rect 109344 62092 109420 62152
rect 21624 61956 21700 62016
rect 21352 61880 21700 61956
rect 27336 61880 27684 62092
rect 109344 61880 109556 62092
rect 114240 62016 114452 62228
rect 114648 62016 114860 62228
rect 115056 62152 115676 62228
rect 115056 62016 115268 62152
rect 115464 62016 115676 62152
rect 115872 62016 116084 62228
rect 134050 62059 134200 62123
rect 21352 61820 21428 61880
rect 27608 61820 27684 61880
rect 109480 61820 109556 61880
rect 20808 61608 21020 61820
rect 21216 61744 21972 61820
rect 21216 61608 21428 61744
rect 21624 61608 21972 61744
rect 22032 61608 22244 61820
rect 22440 61608 22652 61820
rect 27336 61608 27684 61820
rect 109344 61608 109556 61820
rect 114240 61608 114452 61820
rect 114648 61608 114860 61820
rect 115056 61608 115268 61820
rect 115464 61608 115676 61820
rect 115872 61608 116084 61820
rect 27472 61548 27548 61608
rect 109344 61548 109420 61608
rect 20808 61200 21020 61412
rect 21216 61200 21428 61412
rect 21624 61200 21972 61412
rect 22032 61200 22244 61412
rect 22440 61200 22652 61412
rect 27336 61336 27684 61548
rect 27608 61276 27684 61336
rect 20944 61140 21020 61200
rect 21624 61140 21700 61200
rect 1224 60928 1980 61004
rect 1768 60792 1980 60928
rect 20808 60792 21020 61140
rect 21352 61064 21700 61140
rect 27336 61064 27684 61276
rect 109344 61336 109556 61548
rect 132600 61412 132812 61548
rect 133280 61412 133492 61548
rect 109344 61276 109420 61336
rect 109344 61064 109556 61276
rect 114240 61200 114452 61412
rect 114648 61200 114860 61412
rect 115056 61336 115676 61412
rect 115056 61276 115268 61336
rect 115056 61200 115404 61276
rect 115464 61200 115676 61336
rect 115872 61200 116084 61412
rect 132600 61336 133492 61412
rect 115872 61140 115948 61200
rect 21352 61004 21428 61064
rect 27472 61004 27548 61064
rect 109344 61004 109420 61064
rect 21216 60928 21972 61004
rect 21216 60868 21428 60928
rect 21216 60792 21564 60868
rect 21624 60792 21972 60928
rect 22032 60792 22244 61004
rect 22440 60792 22652 61004
rect 20808 60732 20884 60792
rect 21352 60732 21428 60792
rect 20808 60384 21020 60732
rect 21216 60384 21428 60732
rect 21488 60732 21564 60792
rect 21488 60656 21972 60732
rect 21624 60384 21972 60656
rect 22032 60384 22244 60596
rect 22440 60384 22652 60596
rect 27336 60520 27684 61004
rect 109344 60520 109556 61004
rect 114240 60792 114452 61004
rect 114648 60792 114860 61004
rect 115056 60792 115268 61004
rect 115366 60928 115676 61004
rect 115464 60792 115676 60928
rect 115872 60792 116084 61140
rect 134776 60868 134988 61004
rect 134776 60792 135396 60868
rect 115056 60732 115132 60792
rect 115464 60732 115540 60792
rect 116008 60732 116084 60792
rect 27472 60460 27548 60520
rect 109344 60460 109420 60520
rect 20808 60324 20884 60384
rect 20808 60112 21020 60324
rect 27336 60248 27684 60460
rect 109344 60248 109556 60460
rect 114240 60384 114452 60596
rect 114648 60384 114860 60596
rect 115056 60384 115268 60732
rect 115464 60460 115676 60732
rect 115366 60384 115676 60460
rect 115872 60384 116084 60732
rect 115872 60324 115948 60384
rect 27472 60188 27548 60248
rect 109344 60188 109420 60248
rect 21216 59976 21428 60188
rect 21624 59976 21972 60188
rect 22032 59976 22244 60188
rect 22440 59976 22652 60188
rect 21216 59916 21292 59976
rect 21624 59916 21700 59976
rect 22032 59916 22108 59976
rect 22440 59916 22516 59976
rect 20808 59704 21020 59916
rect 21216 59840 21972 59916
rect 21216 59704 21428 59840
rect 21624 59704 21972 59840
rect 22032 59568 22244 59916
rect 22440 59568 22652 59916
rect 27336 59840 27684 60188
rect 109344 59840 109556 60188
rect 114240 59976 114452 60188
rect 114376 59916 114452 59976
rect 22168 59508 22244 59568
rect 22576 59508 22652 59568
rect 20808 59296 21020 59508
rect 1224 59160 1980 59236
rect 1768 59024 1980 59160
rect 21216 59160 21428 59508
rect 21624 59160 21972 59508
rect 22032 59296 22244 59508
rect 22440 59296 22652 59508
rect 27336 59296 27684 59644
rect 109344 59296 109556 59644
rect 114240 59568 114452 59916
rect 114648 59976 114860 60188
rect 115056 60112 115404 60188
rect 115056 60052 115268 60112
rect 115464 60052 115676 60188
rect 115872 60112 116084 60324
rect 115056 59976 115676 60052
rect 114648 59916 114724 59976
rect 115192 59916 115268 59976
rect 114648 59568 114860 59916
rect 115056 59704 115268 59916
rect 115464 59916 115540 59976
rect 115464 59704 115676 59916
rect 115872 59704 116084 59916
rect 114240 59508 114316 59568
rect 114648 59508 114724 59568
rect 114240 59296 114452 59508
rect 114648 59296 114860 59508
rect 115056 59372 115268 59508
rect 115464 59372 115676 59508
rect 115056 59296 115676 59372
rect 115872 59296 116084 59508
rect 27472 59236 27548 59296
rect 109344 59236 109420 59296
rect 21216 59100 21292 59160
rect 21896 59100 21972 59160
rect 20808 58888 21020 59100
rect 21216 58888 21428 59100
rect 21624 58888 21972 59100
rect 22032 58888 22244 59100
rect 22440 58888 22652 59100
rect 27336 59024 27684 59236
rect 109344 59024 109556 59236
rect 115056 59160 115268 59296
rect 115464 59160 115676 59296
rect 115192 59100 115268 59160
rect 115600 59100 115676 59160
rect 134776 59160 135396 59236
rect 27336 58964 27412 59024
rect 109344 58964 109420 59024
rect 21624 58828 21700 58888
rect 21352 58752 21700 58828
rect 21352 58692 21428 58752
rect 20808 58480 21020 58692
rect 21216 58616 21972 58692
rect 21216 58480 21428 58616
rect 21624 58480 21972 58616
rect 22032 58480 22244 58692
rect 22440 58480 22652 58692
rect 27336 58480 27684 58964
rect 109344 58480 109556 58964
rect 114240 58888 114452 59100
rect 114648 58888 114860 59100
rect 115056 58888 115268 59100
rect 115464 58888 115676 59100
rect 115872 58888 116084 59100
rect 134776 59024 134988 59160
rect 114240 58480 114452 58692
rect 114648 58480 114860 58692
rect 115056 58480 115268 58692
rect 115464 58556 115676 58692
rect 115366 58480 115676 58556
rect 115872 58480 116084 58692
rect 27472 58420 27548 58480
rect 109480 58420 109556 58480
rect 20808 58072 21020 58284
rect 21216 58072 21428 58284
rect 21624 58148 21972 58284
rect 21526 58072 21972 58148
rect 22032 58072 22244 58284
rect 22440 58072 22652 58284
rect 27336 58208 27684 58420
rect 109344 58208 109556 58420
rect 27336 58148 27412 58208
rect 109344 58148 109420 58208
rect 27336 57936 27684 58148
rect 109344 57936 109556 58148
rect 114240 58072 114452 58284
rect 114648 58072 114860 58284
rect 115056 58208 115404 58284
rect 115056 58072 115268 58208
rect 115464 58148 115676 58284
rect 115366 58072 115676 58148
rect 115872 58072 116084 58284
rect 27472 57876 27548 57936
rect 109344 57876 109420 57936
rect 20808 57664 21020 57876
rect 21216 57800 21564 57876
rect 21216 57740 21428 57800
rect 21624 57740 21972 57876
rect 21216 57664 21972 57740
rect 22032 57664 22244 57876
rect 22440 57664 22652 57876
rect 27336 57664 27684 57876
rect 109344 57664 109556 57876
rect 114240 57664 114452 57876
rect 114648 57664 114860 57876
rect 115056 57800 115404 57876
rect 115056 57740 115268 57800
rect 115464 57740 115676 57876
rect 115056 57664 115676 57740
rect 115872 57664 116084 57876
rect 21624 57604 21700 57664
rect 27608 57604 27684 57664
rect 109480 57604 109556 57664
rect 1224 57528 1980 57604
rect 1768 57392 1980 57528
rect 21488 57528 21700 57604
rect 21488 57468 21564 57528
rect 20808 57256 21020 57468
rect 21216 57392 21564 57468
rect 21216 57256 21428 57392
rect 21624 57256 21972 57468
rect 22032 57256 22244 57468
rect 22440 57256 22652 57468
rect 27336 57392 27684 57604
rect 109344 57392 109556 57604
rect 134776 57528 135396 57604
rect 27472 57332 27548 57392
rect 109480 57332 109556 57392
rect 20944 57196 21020 57256
rect 20808 56848 21020 57196
rect 27336 57120 27684 57332
rect 109344 57120 109556 57332
rect 114240 57256 114452 57468
rect 114648 57256 114860 57468
rect 115056 57256 115268 57468
rect 115464 57256 115676 57468
rect 115872 57256 116084 57468
rect 134776 57392 134988 57528
rect 116008 57196 116084 57256
rect 27336 57060 27412 57120
rect 109344 57060 109420 57120
rect 20944 56788 21020 56848
rect 20808 56440 21020 56788
rect 21216 56848 21428 57060
rect 21624 56848 21972 57060
rect 22032 56848 22244 57060
rect 22440 56848 22652 57060
rect 27336 56848 27684 57060
rect 109344 56848 109556 57060
rect 114240 56848 114452 57060
rect 114648 56848 114860 57060
rect 115056 56924 115268 57060
rect 115464 56924 115676 57060
rect 115056 56848 115676 56924
rect 115872 56848 116084 57196
rect 21216 56788 21292 56848
rect 21896 56788 21972 56848
rect 21216 56516 21428 56788
rect 21624 56516 21972 56788
rect 27462 56652 27560 56848
rect 109344 56652 109448 56848
rect 115192 56788 115268 56848
rect 115600 56788 115676 56848
rect 116008 56788 116084 56848
rect 21216 56440 21972 56516
rect 22032 56440 22244 56652
rect 22440 56440 22652 56652
rect 27336 56576 27684 56652
rect 109344 56576 109556 56652
rect 27472 56516 27548 56576
rect 109344 56516 109420 56576
rect 20808 56380 20884 56440
rect 20808 56168 21020 56380
rect 27336 56304 27684 56516
rect 109344 56304 109556 56516
rect 114240 56440 114452 56652
rect 114648 56440 114860 56652
rect 115056 56440 115268 56788
rect 115464 56440 115676 56788
rect 115872 56440 116084 56788
rect 116008 56380 116084 56440
rect 27608 56244 27684 56304
rect 109480 56244 109556 56304
rect 21216 56032 21428 56244
rect 21624 56032 21972 56244
rect 21216 55972 21292 56032
rect 21896 55972 21972 56032
rect 1224 55896 1980 55972
rect 1768 55760 1980 55896
rect 20808 55760 21020 55972
rect 21216 55760 21428 55972
rect 21624 55836 21972 55972
rect 21526 55760 21972 55836
rect 22032 56032 22244 56244
rect 22440 56032 22652 56244
rect 22032 55972 22108 56032
rect 22440 55972 22516 56032
rect 22032 55624 22244 55972
rect 22440 55624 22652 55972
rect 27336 55896 27684 56244
rect 109344 55896 109556 56244
rect 114240 56032 114452 56244
rect 114648 56032 114860 56244
rect 115056 56032 115268 56244
rect 115464 56108 115676 56244
rect 115872 56168 116084 56380
rect 115366 56032 115676 56108
rect 114376 55972 114452 56032
rect 114784 55972 114860 56032
rect 115192 55972 115268 56032
rect 22032 55564 22108 55624
rect 22440 55564 22516 55624
rect 20808 55352 21020 55564
rect 21216 55488 21564 55564
rect 21216 55428 21428 55488
rect 21624 55428 21972 55564
rect 21216 55352 21972 55428
rect 21216 55216 21428 55352
rect 21624 55216 21972 55352
rect 22032 55216 22244 55564
rect 22440 55216 22652 55564
rect 21216 55156 21292 55216
rect 21624 55156 21700 55216
rect 22032 55156 22108 55216
rect 22440 55156 22516 55216
rect 20808 54944 21020 55156
rect 21216 54944 21428 55156
rect 21624 54944 21972 55156
rect 22032 54944 22244 55156
rect 22440 54944 22652 55156
rect 27336 55080 27684 55700
rect 109344 55080 109556 55700
rect 114240 55624 114452 55972
rect 114376 55564 114452 55624
rect 27608 55020 27684 55080
rect 109480 55020 109556 55080
rect 20808 54536 21020 54748
rect 21216 54536 21428 54748
rect 21624 54612 21972 54748
rect 21526 54536 21972 54612
rect 22032 54536 22244 54748
rect 22440 54536 22652 54748
rect 27336 54536 27684 55020
rect 27608 54476 27684 54536
rect 1224 54128 1980 54204
rect 20808 54128 21020 54340
rect 21216 54264 21564 54340
rect 21216 54204 21428 54264
rect 21624 54204 21972 54340
rect 21216 54128 21972 54204
rect 22032 54128 22244 54340
rect 22440 54128 22652 54340
rect 27336 54264 27684 54476
rect 109344 54536 109556 55020
rect 114240 55216 114452 55564
rect 114648 55624 114860 55972
rect 115056 55896 115676 55972
rect 115056 55836 115268 55896
rect 115056 55760 115404 55836
rect 115464 55760 115676 55896
rect 115872 55760 116084 55972
rect 134776 55896 135396 55972
rect 134776 55760 134988 55896
rect 114648 55564 114724 55624
rect 114648 55216 114860 55564
rect 115056 55216 115268 55564
rect 115366 55488 115676 55564
rect 115464 55216 115676 55488
rect 115872 55352 116084 55564
rect 114240 55156 114316 55216
rect 114648 55156 114724 55216
rect 115056 55156 115132 55216
rect 115600 55156 115676 55216
rect 114240 54944 114452 55156
rect 114648 54944 114860 55156
rect 115056 54944 115268 55156
rect 115464 55020 115676 55156
rect 115366 54944 115676 55020
rect 115872 54944 116084 55156
rect 114240 54536 114452 54748
rect 114648 54536 114860 54748
rect 115056 54672 115404 54748
rect 115056 54612 115268 54672
rect 115464 54612 115676 54748
rect 115056 54536 115676 54612
rect 115872 54536 116084 54748
rect 109344 54476 109420 54536
rect 109344 54264 109556 54476
rect 27608 54204 27684 54264
rect 109480 54204 109556 54264
rect 1768 53992 1980 54128
rect 27336 53992 27684 54204
rect 109344 53992 109556 54204
rect 114240 54128 114452 54340
rect 114648 54128 114860 54340
rect 115056 54128 115268 54340
rect 115464 54204 115676 54340
rect 115366 54128 115676 54204
rect 115872 54128 116084 54340
rect 134776 54068 134988 54204
rect 134776 53992 135396 54068
rect 27336 53932 27412 53992
rect 109344 53932 109420 53992
rect 20808 53720 21020 53932
rect 21216 53856 21972 53932
rect 21216 53720 21428 53856
rect 21624 53720 21972 53856
rect 22032 53720 22244 53932
rect 22440 53720 22652 53932
rect 27336 53720 27684 53932
rect 109344 53720 109556 53932
rect 114240 53720 114452 53932
rect 114648 53720 114860 53932
rect 115056 53856 115404 53932
rect 115056 53796 115268 53856
rect 115464 53796 115676 53932
rect 115056 53720 115676 53796
rect 115872 53720 116084 53932
rect 27336 53660 27412 53720
rect 109344 53660 109420 53720
rect 115464 53660 115540 53720
rect 20808 53312 21020 53524
rect 21216 53448 21972 53524
rect 21216 53388 21428 53448
rect 21216 53312 21564 53388
rect 21624 53312 21972 53448
rect 22032 53312 22244 53524
rect 22440 53312 22652 53524
rect 27336 53448 27684 53660
rect 109344 53448 109556 53660
rect 115192 53584 115540 53660
rect 115192 53524 115268 53584
rect 27336 53388 27412 53448
rect 109480 53388 109556 53448
rect 20944 53252 21020 53312
rect 20808 52904 21020 53252
rect 27336 53176 27684 53388
rect 109344 53176 109556 53388
rect 114240 53312 114452 53524
rect 114648 53312 114860 53524
rect 115056 53448 115676 53524
rect 115056 53312 115268 53448
rect 115464 53312 115676 53448
rect 115872 53312 116084 53524
rect 116008 53252 116084 53312
rect 27608 53116 27684 53176
rect 109480 53116 109556 53176
rect 21216 52904 21428 53116
rect 21526 53040 21972 53116
rect 21624 52904 21972 53040
rect 22032 52904 22244 53116
rect 22440 52904 22652 53116
rect 27336 52904 27684 53116
rect 109344 52904 109556 53116
rect 114240 52904 114452 53116
rect 114648 52904 114860 53116
rect 115056 52904 115268 53116
rect 115464 52904 115676 53116
rect 115872 52904 116084 53252
rect 27336 52844 27412 52904
rect 109480 52844 109556 52904
rect 1224 52496 1980 52572
rect 20808 52496 21020 52708
rect 21216 52496 21428 52708
rect 21624 52496 21972 52708
rect 22032 52496 22244 52708
rect 22440 52496 22652 52708
rect 27336 52632 27684 52844
rect 27608 52572 27684 52632
rect 1768 52360 1980 52496
rect 20944 52436 21020 52496
rect 21624 52436 21700 52496
rect 20808 52224 21020 52436
rect 21352 52360 21700 52436
rect 27336 52360 27684 52572
rect 109344 52632 109556 52844
rect 109344 52572 109420 52632
rect 109344 52360 109556 52572
rect 114240 52496 114452 52708
rect 114648 52496 114860 52708
rect 115056 52572 115268 52708
rect 115464 52572 115676 52708
rect 115056 52496 115676 52572
rect 115872 52496 116084 52708
rect 115192 52436 115268 52496
rect 115872 52436 115948 52496
rect 134776 52436 134988 52572
rect 115192 52360 115540 52436
rect 21352 52300 21428 52360
rect 27472 52300 27548 52360
rect 109480 52300 109556 52360
rect 115464 52300 115540 52360
rect 21216 52224 21972 52300
rect 21216 52164 21428 52224
rect 21216 52088 21564 52164
rect 21624 52088 21972 52224
rect 22032 52088 22244 52300
rect 22440 52088 22652 52300
rect 21352 52028 21428 52088
rect 20808 51680 21020 52028
rect 21216 51680 21428 52028
rect 21488 52028 21564 52088
rect 21488 51952 21972 52028
rect 21624 51680 21972 51952
rect 22032 51680 22244 51892
rect 22440 51680 22652 51892
rect 27336 51816 27684 52300
rect 27608 51756 27684 51816
rect 20808 51620 20884 51680
rect 22032 51620 22108 51680
rect 22576 51620 22652 51680
rect 20808 51408 21020 51620
rect 21216 51272 21428 51484
rect 21624 51348 21972 51484
rect 21488 51272 21972 51348
rect 22032 51272 22244 51620
rect 22440 51272 22652 51620
rect 21216 51212 21292 51272
rect 21488 51212 21564 51272
rect 20808 51000 21020 51212
rect 21216 51136 21564 51212
rect 21624 51212 21700 51272
rect 22032 51212 22108 51272
rect 22440 51212 22516 51272
rect 21216 51000 21428 51136
rect 21624 51000 21972 51212
rect 22032 51000 22244 51212
rect 22440 51000 22652 51212
rect 27336 51136 27684 51756
rect 27608 51076 27684 51136
rect 1224 50864 1980 50940
rect 1768 50728 1980 50864
rect 20808 50592 21020 50804
rect 21216 50592 21428 50804
rect 21624 50592 21972 50804
rect 22032 50592 22244 50804
rect 22440 50592 22652 50804
rect 27336 50592 27684 51076
rect 109344 51816 109556 52300
rect 114240 52088 114452 52300
rect 114648 52088 114860 52300
rect 115056 52088 115268 52300
rect 115464 52088 115676 52300
rect 115872 52224 116084 52436
rect 134776 52360 135396 52436
rect 115056 52028 115132 52088
rect 109344 51756 109420 51816
rect 109344 51136 109556 51756
rect 114240 51680 114452 51892
rect 114648 51680 114860 51892
rect 115056 51680 115268 52028
rect 115464 51680 115676 52028
rect 115872 51680 116084 52028
rect 114376 51620 114452 51680
rect 114784 51620 114860 51680
rect 115464 51620 115540 51680
rect 114240 51272 114452 51620
rect 114648 51272 114860 51620
rect 115192 51544 115540 51620
rect 115872 51620 115948 51680
rect 115192 51484 115268 51544
rect 115056 51408 115676 51484
rect 115872 51408 116084 51620
rect 115056 51272 115268 51408
rect 114240 51212 114316 51272
rect 114784 51212 114860 51272
rect 115192 51212 115268 51272
rect 109344 51076 109420 51136
rect 109344 50592 109556 51076
rect 114240 51000 114452 51212
rect 114648 51000 114860 51212
rect 115056 51000 115268 51212
rect 115464 51272 115676 51408
rect 115464 51212 115540 51272
rect 115464 51000 115676 51212
rect 115872 51000 116084 51212
rect 134776 50804 134988 50940
rect 114240 50592 114452 50804
rect 114648 50592 114860 50804
rect 115056 50592 115268 50804
rect 115464 50592 115676 50804
rect 115872 50592 116084 50804
rect 134776 50728 135396 50804
rect 27472 50532 27548 50592
rect 109344 50532 109420 50592
rect 115464 50532 115540 50592
rect 20808 50184 21020 50396
rect 21216 50184 21428 50396
rect 21624 50260 21972 50396
rect 21526 50184 21972 50260
rect 22032 50184 22244 50396
rect 22440 50184 22652 50396
rect 27336 50320 27684 50532
rect 109344 50320 109556 50532
rect 115192 50456 115540 50532
rect 115192 50396 115268 50456
rect 27336 50260 27412 50320
rect 109344 50260 109420 50320
rect 27336 50048 27684 50260
rect 109344 50048 109556 50260
rect 114240 50184 114452 50396
rect 114648 50184 114860 50396
rect 115056 50320 115676 50396
rect 115056 50184 115268 50320
rect 115464 50184 115676 50320
rect 115872 50184 116084 50396
rect 27608 49988 27684 50048
rect 109480 49988 109556 50048
rect 20808 49776 21020 49988
rect 21216 49912 21564 49988
rect 21216 49852 21428 49912
rect 21624 49852 21972 49988
rect 21216 49776 21972 49852
rect 22032 49776 22244 49988
rect 22440 49776 22652 49988
rect 27336 49776 27684 49988
rect 109344 49776 109556 49988
rect 114240 49776 114452 49988
rect 114648 49776 114860 49988
rect 115056 49776 115268 49988
rect 115464 49852 115676 49988
rect 115366 49776 115676 49852
rect 115872 49776 116084 49988
rect 27472 49716 27548 49776
rect 109480 49716 109556 49776
rect 20808 49368 21020 49580
rect 21216 49368 21428 49580
rect 21624 49368 21972 49580
rect 22032 49368 22244 49580
rect 22440 49368 22652 49580
rect 27336 49504 27684 49716
rect 109344 49504 109556 49716
rect 27336 49444 27412 49504
rect 109344 49444 109420 49504
rect 27336 49232 27684 49444
rect 109344 49232 109556 49444
rect 114240 49368 114452 49580
rect 114648 49368 114860 49580
rect 115056 49504 115404 49580
rect 115056 49444 115268 49504
rect 115464 49444 115676 49580
rect 115056 49368 115676 49444
rect 115872 49368 116084 49580
rect 115464 49308 115540 49368
rect 115192 49232 115540 49308
rect 27472 49172 27548 49232
rect 109344 49172 109420 49232
rect 115192 49172 115268 49232
rect 1768 49036 1980 49172
rect 1224 48960 1980 49036
rect 20808 48960 21020 49172
rect 21216 48960 21428 49172
rect 21624 49036 21972 49172
rect 21526 48960 21972 49036
rect 22032 48960 22244 49172
rect 22440 48960 22652 49172
rect 27336 48960 27684 49172
rect 109344 48960 109556 49172
rect 114240 48960 114452 49172
rect 114648 48960 114860 49172
rect 115056 49096 115676 49172
rect 115056 48960 115268 49096
rect 115464 48960 115676 49096
rect 115872 48960 116084 49172
rect 134776 49036 134988 49172
rect 134776 48960 135396 49036
rect 27336 48900 27412 48960
rect 109480 48900 109556 48960
rect 20808 48552 21020 48764
rect 21216 48688 21564 48764
rect 21216 48628 21428 48688
rect 21624 48628 21972 48764
rect 21216 48552 21972 48628
rect 22032 48552 22244 48764
rect 22440 48552 22652 48764
rect 27336 48688 27684 48900
rect 109344 48688 109556 48900
rect 27472 48628 27548 48688
rect 109480 48628 109556 48688
rect 20808 48492 20884 48552
rect 20808 48280 21020 48492
rect 27336 48416 27684 48628
rect 109344 48416 109556 48628
rect 114240 48552 114452 48764
rect 114648 48552 114860 48764
rect 115056 48552 115268 48764
rect 115464 48552 115676 48764
rect 115872 48552 116084 48764
rect 115872 48492 115948 48552
rect 27336 48356 27412 48416
rect 109344 48356 109420 48416
rect 21216 48144 21428 48356
rect 21624 48144 21972 48356
rect 22032 48144 22244 48356
rect 22440 48144 22652 48356
rect 21216 48084 21292 48144
rect 21896 48084 21972 48144
rect 20808 47736 21020 48084
rect 21216 47948 21428 48084
rect 21624 47948 21972 48084
rect 21216 47872 21972 47948
rect 21216 47812 21428 47872
rect 21216 47736 21564 47812
rect 21624 47736 21972 47872
rect 22032 47736 22244 47948
rect 20944 47676 21020 47736
rect 22168 47676 22244 47736
rect 1224 47464 1980 47540
rect 20808 47464 21020 47676
rect 1768 47328 1980 47464
rect 21216 47328 21428 47540
rect 21526 47464 21972 47540
rect 21624 47328 21972 47464
rect 22032 47328 22244 47676
rect 22440 47736 22652 47948
rect 27336 47872 27684 48356
rect 109344 47872 109556 48356
rect 114240 48144 114452 48356
rect 114648 48144 114860 48356
rect 115056 48280 115404 48356
rect 115056 48220 115268 48280
rect 115464 48220 115676 48356
rect 115872 48280 116084 48492
rect 115056 48144 115676 48220
rect 115192 48084 115268 48144
rect 27472 47812 27548 47872
rect 109344 47812 109420 47872
rect 22440 47676 22516 47736
rect 22440 47328 22652 47676
rect 21216 47268 21292 47328
rect 21624 47268 21700 47328
rect 22032 47268 22108 47328
rect 22576 47268 22652 47328
rect 20808 47056 21020 47268
rect 21216 47056 21428 47268
rect 21624 47056 21972 47268
rect 22032 46920 22244 47268
rect 22168 46860 22244 46920
rect 20808 46648 21020 46860
rect 21216 46724 21428 46860
rect 21624 46724 21972 46860
rect 21216 46648 21972 46724
rect 22032 46648 22244 46860
rect 22440 46920 22652 47268
rect 27336 47192 27684 47812
rect 109344 47192 109556 47812
rect 114240 47736 114452 47948
rect 114648 47736 114860 47948
rect 115056 47736 115268 48084
rect 115366 48008 115676 48084
rect 115464 47736 115676 48008
rect 115872 47736 116084 48084
rect 114240 47676 114316 47736
rect 114648 47676 114724 47736
rect 116008 47676 116084 47736
rect 114240 47328 114452 47676
rect 114648 47328 114860 47676
rect 115056 47328 115268 47540
rect 114376 47268 114452 47328
rect 114784 47268 114860 47328
rect 115192 47268 115268 47328
rect 115464 47328 115676 47540
rect 115872 47464 116084 47676
rect 134776 47464 135396 47540
rect 134776 47328 134988 47464
rect 115464 47268 115540 47328
rect 22440 46860 22516 46920
rect 22440 46648 22652 46860
rect 27336 46648 27684 46996
rect 109344 46648 109556 46996
rect 114240 46920 114452 47268
rect 114648 46920 114860 47268
rect 115056 47192 115676 47268
rect 115056 47132 115268 47192
rect 115056 47056 115404 47132
rect 115464 47056 115676 47192
rect 115872 47056 116084 47268
rect 114240 46860 114316 46920
rect 114648 46860 114724 46920
rect 114240 46648 114452 46860
rect 114648 46648 114860 46860
rect 21216 46512 21428 46648
rect 21624 46512 21972 46648
rect 21352 46452 21428 46512
rect 21896 46452 21972 46512
rect 27336 46588 27412 46648
rect 109480 46588 109556 46648
rect 20808 46240 21020 46452
rect 21216 46240 21428 46452
rect 21624 46240 21972 46452
rect 22032 46240 22244 46452
rect 22440 46240 22652 46452
rect 27336 46376 27684 46588
rect 109344 46376 109556 46588
rect 115056 46512 115268 46860
rect 115366 46784 115676 46860
rect 115464 46512 115676 46784
rect 115872 46648 116084 46860
rect 115056 46452 115132 46512
rect 115600 46452 115676 46512
rect 27608 46316 27684 46376
rect 109480 46316 109556 46376
rect 27336 46240 27684 46316
rect 109344 46240 109556 46316
rect 114240 46240 114452 46452
rect 114648 46240 114860 46452
rect 115056 46240 115268 46452
rect 115464 46316 115676 46452
rect 115366 46240 115676 46316
rect 115872 46240 116084 46452
rect 27462 46044 27560 46240
rect 109344 46044 109448 46240
rect 1768 45636 1980 45908
rect 20808 45832 21020 46044
rect 21216 45832 21428 46044
rect 21624 45832 21972 46044
rect 22032 45832 22244 46044
rect 22440 45832 22652 46044
rect 27336 45832 27684 46044
rect 109344 45832 109556 46044
rect 114240 45832 114452 46044
rect 114648 45908 114860 46044
rect 115056 45968 115404 46044
rect 114648 45832 114996 45908
rect 115056 45832 115268 45968
rect 115464 45832 115676 46044
rect 115872 45832 116084 46044
rect 21624 45772 21700 45832
rect 27608 45772 27684 45832
rect 109480 45772 109556 45832
rect 21352 45696 21700 45772
rect 21352 45636 21428 45696
rect 1224 45560 1980 45636
rect 20808 45424 21020 45636
rect 21216 45560 21972 45636
rect 21216 45424 21428 45560
rect 21624 45424 21972 45560
rect 22032 45500 22244 45636
rect 22032 45424 22380 45500
rect 22440 45424 22652 45636
rect 27336 45560 27684 45772
rect 109344 45560 109556 45772
rect 114920 45772 114996 45832
rect 115872 45772 115948 45832
rect 114920 45696 115948 45772
rect 134776 45772 134988 45908
rect 134776 45696 135396 45772
rect 27472 45500 27548 45560
rect 109480 45500 109556 45560
rect 114240 45500 114452 45636
rect 25878 45424 27684 45500
rect 22304 45364 22380 45424
rect 22304 45288 22924 45364
rect 22848 45228 22924 45288
rect 24208 45288 26052 45364
rect 27336 45288 27684 45424
rect 109344 45288 109556 45500
rect 113734 45424 114452 45500
rect 114648 45424 114860 45636
rect 115056 45424 115268 45636
rect 115464 45500 115676 45636
rect 115366 45424 115676 45500
rect 115872 45424 116084 45636
rect 134776 45560 134988 45696
rect 114648 45364 114724 45424
rect 24208 45228 24284 45288
rect 25976 45228 26052 45288
rect 27472 45228 27548 45288
rect 109480 45228 109556 45288
rect 112200 45288 113500 45364
rect 112200 45228 112276 45288
rect 113424 45228 113500 45288
rect 114104 45288 114724 45364
rect 114104 45228 114180 45288
rect 20808 45016 21020 45228
rect 21216 45016 21428 45228
rect 21624 45092 21972 45228
rect 21526 45016 21972 45092
rect 22032 45016 22244 45228
rect 22440 45016 22652 45228
rect 22848 45092 23060 45228
rect 23256 45152 24284 45228
rect 24344 45152 25916 45228
rect 22848 45016 23196 45092
rect 23256 45016 23604 45152
rect 24344 45016 24556 45152
rect 25976 45016 26188 45228
rect 27336 45016 27684 45228
rect 109344 45016 109556 45228
rect 110704 45152 112276 45228
rect 110704 45016 110916 45152
rect 112336 45092 112548 45228
rect 113424 45152 113772 45228
rect 113832 45152 114180 45228
rect 112336 45016 113364 45092
rect 113424 45016 113636 45152
rect 113832 45016 114044 45152
rect 114240 45016 114452 45228
rect 114648 45016 114860 45228
rect 115056 45152 115404 45228
rect 115056 45092 115268 45152
rect 115464 45092 115676 45228
rect 115056 45016 115676 45092
rect 115872 45016 116084 45228
rect 23120 44956 23196 45016
rect 24344 44956 24420 45016
rect 27472 44956 27548 45016
rect 109344 44956 109420 45016
rect 113288 44956 113364 45016
rect 113832 44956 113908 45016
rect 115464 44956 115540 45016
rect 23120 44880 24420 44956
rect 20808 44608 21020 44820
rect 21216 44744 21564 44820
rect 21216 44684 21428 44744
rect 21624 44684 21972 44820
rect 21216 44608 21972 44684
rect 22032 44608 22244 44820
rect 22440 44744 23332 44820
rect 27336 44744 27684 44956
rect 109344 44744 109556 44956
rect 113288 44880 113908 44956
rect 115192 44880 115540 44956
rect 115192 44820 115268 44880
rect 22440 44608 22652 44744
rect 27472 44684 27548 44744
rect 109344 44684 109420 44744
rect 20808 44548 20884 44608
rect 21352 44548 21428 44608
rect 20808 44200 21020 44548
rect 21352 44472 21700 44548
rect 27336 44472 27684 44684
rect 109344 44608 112412 44684
rect 114240 44608 114452 44820
rect 114648 44608 114860 44820
rect 115056 44744 115676 44820
rect 115056 44608 115268 44744
rect 115464 44608 115676 44744
rect 115872 44608 116084 44820
rect 109344 44472 109556 44608
rect 21624 44412 21700 44472
rect 27608 44412 27684 44472
rect 109480 44412 109556 44472
rect 115872 44548 115948 44608
rect 21216 44200 21428 44412
rect 21624 44200 21972 44412
rect 22032 44200 22244 44412
rect 22440 44200 22652 44412
rect 20808 44140 20884 44200
rect 21352 44140 21428 44200
rect 21760 44140 21836 44200
rect 1224 44064 1980 44140
rect 1768 43928 1980 44064
rect 20808 43792 21020 44140
rect 21216 43792 21428 44140
rect 21624 43792 21972 44140
rect 22032 43792 22244 44004
rect 22440 43792 22652 44004
rect 27336 43928 27684 44412
rect 27608 43868 27684 43928
rect 20808 43732 20884 43792
rect 20808 43520 21020 43732
rect 27336 43656 27684 43868
rect 109344 43928 109556 44412
rect 114240 44200 114452 44412
rect 114648 44200 114860 44412
rect 115056 44336 115676 44412
rect 115056 44276 115268 44336
rect 115056 44200 115404 44276
rect 115464 44200 115676 44336
rect 115872 44200 116084 44548
rect 115328 44140 115404 44200
rect 115872 44140 115948 44200
rect 109344 43868 109420 43928
rect 109344 43656 109556 43868
rect 114240 43792 114452 44004
rect 114648 43792 114860 44004
rect 115056 43868 115268 44140
rect 115328 44064 115676 44140
rect 115464 43868 115676 44064
rect 115056 43792 115676 43868
rect 115872 43792 116084 44140
rect 134776 44004 134988 44140
rect 134776 43928 135396 44004
rect 115192 43732 115268 43792
rect 115872 43732 115948 43792
rect 115192 43656 115540 43732
rect 27472 43596 27548 43656
rect 109344 43596 109420 43656
rect 115464 43596 115540 43656
rect 21216 43460 21428 43596
rect 21216 43384 21564 43460
rect 21624 43384 21972 43596
rect 22032 43384 22244 43596
rect 21488 43324 21564 43384
rect 21896 43324 21972 43384
rect 22168 43324 22244 43384
rect 20808 43112 21020 43324
rect 21216 43188 21428 43324
rect 21488 43248 21972 43324
rect 21216 43112 21564 43188
rect 21624 43112 21972 43248
rect 22032 42976 22244 43324
rect 22440 43384 22652 43596
rect 22440 43324 22516 43384
rect 22440 42976 22652 43324
rect 27336 43248 27684 43596
rect 109344 43248 109556 43596
rect 114240 43384 114452 43596
rect 114648 43384 114860 43596
rect 115056 43384 115268 43596
rect 115464 43384 115676 43596
rect 115872 43520 116084 43732
rect 114240 43324 114316 43384
rect 114648 43324 114724 43384
rect 115056 43324 115132 43384
rect 115464 43324 115540 43384
rect 22168 42916 22244 42976
rect 22576 42916 22652 42976
rect 20808 42704 21020 42916
rect 21216 42644 21428 42916
rect 21624 42644 21972 42916
rect 22032 42704 22244 42916
rect 22440 42704 22652 42916
rect 27336 42704 27684 43052
rect 109344 42704 109556 43052
rect 114240 42976 114452 43324
rect 114648 42976 114860 43324
rect 115056 43112 115268 43324
rect 115464 43112 115676 43324
rect 115872 43112 116084 43324
rect 114240 42916 114316 42976
rect 114784 42916 114860 42976
rect 114240 42704 114452 42916
rect 114648 42704 114860 42916
rect 21216 42568 21972 42644
rect 27336 42644 27412 42704
rect 109344 42644 109420 42704
rect 115056 42644 115268 42916
rect 21624 42508 21700 42568
rect 1224 42432 1980 42508
rect 1768 42296 1980 42432
rect 20808 42296 21020 42508
rect 21216 42432 21972 42508
rect 21216 42296 21428 42432
rect 21624 42296 21972 42432
rect 22032 42296 22244 42508
rect 22440 42296 22652 42508
rect 27336 42432 27684 42644
rect 109344 42432 109556 42644
rect 115056 42568 115404 42644
rect 115056 42508 115132 42568
rect 115328 42508 115404 42568
rect 115464 42568 115676 42916
rect 115872 42704 116084 42916
rect 115464 42508 115540 42568
rect 27472 42372 27548 42432
rect 109344 42372 109420 42432
rect 20808 41888 21020 42100
rect 21216 41888 21428 42100
rect 21624 41888 21972 42100
rect 22032 41888 22244 42100
rect 22440 41888 22652 42100
rect 27336 41888 27684 42372
rect 27608 41828 27684 41888
rect 20808 41480 21020 41692
rect 21216 41480 21428 41692
rect 21624 41480 21972 41692
rect 22032 41480 22244 41692
rect 22440 41480 22652 41692
rect 27336 41616 27684 41828
rect 27608 41556 27684 41616
rect 21624 41420 21700 41480
rect 21352 41344 21700 41420
rect 27336 41344 27684 41556
rect 109344 41888 109556 42372
rect 114240 42296 114452 42508
rect 114648 42296 114860 42508
rect 115056 42296 115268 42508
rect 115328 42432 115676 42508
rect 115464 42296 115676 42432
rect 115872 42296 116084 42508
rect 134776 42372 134988 42508
rect 134776 42296 135396 42372
rect 114240 41888 114452 42100
rect 114648 41888 114860 42100
rect 115056 41888 115268 42100
rect 115464 41964 115676 42100
rect 115366 41888 115676 41964
rect 115872 41888 116084 42100
rect 109344 41828 109420 41888
rect 109344 41616 109556 41828
rect 109344 41556 109420 41616
rect 109344 41344 109556 41556
rect 114240 41480 114452 41692
rect 114648 41480 114860 41692
rect 115056 41616 115404 41692
rect 115056 41556 115268 41616
rect 115464 41556 115676 41692
rect 115056 41480 115676 41556
rect 115872 41480 116084 41692
rect 21352 41284 21428 41344
rect 27608 41284 27684 41344
rect 109480 41284 109556 41344
rect 20808 41072 21020 41284
rect 21216 41208 21972 41284
rect 21216 41072 21428 41208
rect 21624 41072 21972 41208
rect 22032 41072 22244 41284
rect 22440 41072 22652 41284
rect 27336 41072 27684 41284
rect 109344 41072 109556 41284
rect 114240 41072 114452 41284
rect 114648 41072 114860 41284
rect 115056 41072 115268 41284
rect 115464 41148 115676 41284
rect 115366 41072 115676 41148
rect 115872 41072 116084 41284
rect 27472 41012 27548 41072
rect 109480 41012 109556 41072
rect 1224 40800 1980 40876
rect 1768 40528 1980 40800
rect 20808 40664 21020 40876
rect 21216 40664 21428 40876
rect 21624 40664 21972 40876
rect 22032 40664 22244 40876
rect 22440 40664 22652 40876
rect 27336 40800 27684 41012
rect 109344 40800 109556 41012
rect 27336 40740 27412 40800
rect 109344 40740 109420 40800
rect 20808 40604 20884 40664
rect 20808 40256 21020 40604
rect 27336 40528 27684 40740
rect 109344 40528 109556 40740
rect 114240 40664 114452 40876
rect 114648 40664 114860 40876
rect 115056 40800 115404 40876
rect 115056 40664 115268 40800
rect 115464 40740 115676 40876
rect 115366 40664 115676 40740
rect 115872 40664 116084 40876
rect 134776 40800 135396 40876
rect 115872 40604 115948 40664
rect 27472 40468 27548 40528
rect 109344 40468 109420 40528
rect 21216 40256 21428 40468
rect 21624 40332 21972 40468
rect 21488 40256 21972 40332
rect 22032 40256 22244 40468
rect 22440 40256 22652 40468
rect 20808 40196 20884 40256
rect 21216 40196 21292 40256
rect 21488 40196 21564 40256
rect 20808 39848 21020 40196
rect 21216 40120 21564 40196
rect 21216 39924 21428 40120
rect 21624 39924 21972 40196
rect 21216 39848 21972 39924
rect 22032 39848 22244 40060
rect 22440 39848 22652 40060
rect 27336 39984 27684 40468
rect 109344 39984 109556 40468
rect 114240 40256 114452 40468
rect 114648 40256 114860 40468
rect 115056 40392 115404 40468
rect 115056 40332 115268 40392
rect 115464 40332 115676 40468
rect 115056 40256 115676 40332
rect 115872 40256 116084 40604
rect 134776 40528 134988 40800
rect 115192 40196 115268 40256
rect 115872 40196 115948 40256
rect 27608 39924 27684 39984
rect 20808 39788 20884 39848
rect 20808 39576 21020 39788
rect 27336 39712 27684 39924
rect 27608 39652 27684 39712
rect 21216 39440 21428 39652
rect 21624 39516 21972 39652
rect 21488 39440 21972 39516
rect 21216 39380 21292 39440
rect 21488 39380 21564 39440
rect 21896 39380 21972 39440
rect 20808 39168 21020 39380
rect 21216 39304 21564 39380
rect 21216 39168 21428 39304
rect 21624 39244 21972 39380
rect 21526 39168 21972 39244
rect 22032 39440 22244 39652
rect 22440 39440 22652 39652
rect 22032 39380 22108 39440
rect 22576 39380 22652 39440
rect 21352 39108 21428 39168
rect 1224 39032 1980 39108
rect 21352 39032 21700 39108
rect 1768 38896 1980 39032
rect 21624 38972 21700 39032
rect 22032 39032 22244 39380
rect 22440 39032 22652 39380
rect 27336 39304 27684 39652
rect 109344 39712 109556 39924
rect 114240 39848 114452 40060
rect 114648 39848 114860 40060
rect 115056 39848 115268 40196
rect 115366 40120 115676 40196
rect 115464 39848 115676 40120
rect 115872 39848 116084 40196
rect 115872 39788 115948 39848
rect 109344 39652 109420 39712
rect 109344 39304 109556 39652
rect 114240 39440 114452 39652
rect 114648 39440 114860 39652
rect 115056 39440 115268 39652
rect 115464 39516 115676 39652
rect 115872 39576 116084 39788
rect 114376 39380 114452 39440
rect 114784 39380 114860 39440
rect 115192 39380 115268 39440
rect 115328 39440 115676 39516
rect 115328 39380 115404 39440
rect 115600 39380 115676 39440
rect 22032 38972 22108 39032
rect 22440 38972 22516 39032
rect 20808 38760 21020 38972
rect 21216 38896 21564 38972
rect 21216 38624 21428 38896
rect 21624 38624 21972 38972
rect 21896 38564 21972 38624
rect 20808 38352 21020 38564
rect 21216 38352 21428 38564
rect 21624 38352 21972 38564
rect 22032 38624 22244 38972
rect 22440 38624 22652 38972
rect 22032 38564 22108 38624
rect 22576 38564 22652 38624
rect 22032 38352 22244 38564
rect 22440 38352 22652 38564
rect 27336 38488 27684 39108
rect 109344 38488 109556 39108
rect 114240 39032 114452 39380
rect 114648 39032 114860 39380
rect 115056 39304 115404 39380
rect 115056 39168 115268 39304
rect 115464 39168 115676 39380
rect 115872 39168 116084 39380
rect 134776 39032 135396 39108
rect 114240 38972 114316 39032
rect 114648 38972 114724 39032
rect 114240 38624 114452 38972
rect 114648 38624 114860 38972
rect 115056 38624 115268 38972
rect 114240 38564 114316 38624
rect 114784 38564 114860 38624
rect 115192 38564 115268 38624
rect 115464 38624 115676 38972
rect 115872 38760 116084 38972
rect 134776 38896 134988 39032
rect 115464 38564 115540 38624
rect 27472 38428 27548 38488
rect 109344 38428 109420 38488
rect 21624 38292 21700 38352
rect 21352 38216 21700 38292
rect 21352 38156 21428 38216
rect 20808 37944 21020 38156
rect 21216 38080 21972 38156
rect 21216 37944 21428 38080
rect 21624 37944 21972 38080
rect 22032 37944 22244 38156
rect 22440 37944 22652 38156
rect 27336 37944 27684 38428
rect 109344 37944 109556 38428
rect 114240 38352 114452 38564
rect 114648 38352 114860 38564
rect 115056 38488 115676 38564
rect 115056 38428 115268 38488
rect 115056 38352 115404 38428
rect 115464 38352 115676 38488
rect 115872 38352 116084 38564
rect 114240 37944 114452 38156
rect 114648 37944 114860 38156
rect 115056 37944 115268 38156
rect 115366 38080 115676 38156
rect 115464 37944 115676 38080
rect 115872 37944 116084 38156
rect 27336 37884 27412 37944
rect 109480 37884 109556 37944
rect 14008 37536 14220 37748
rect 20808 37536 21020 37748
rect 21216 37536 21428 37748
rect 21624 37536 21972 37748
rect 22032 37536 22244 37748
rect 22440 37536 22652 37748
rect 27336 37672 27684 37884
rect 27608 37612 27684 37672
rect 1768 37340 1980 37476
rect 27336 37400 27684 37612
rect 109344 37672 109556 37884
rect 109344 37612 109420 37672
rect 109344 37400 109556 37612
rect 114240 37536 114452 37748
rect 114648 37536 114860 37748
rect 115056 37536 115268 37748
rect 115464 37536 115676 37748
rect 115872 37536 116084 37748
rect 115464 37476 115540 37536
rect 115192 37400 115540 37476
rect 134776 37400 135396 37476
rect 27336 37340 27412 37400
rect 109344 37340 109420 37400
rect 115192 37340 115268 37400
rect 1224 37264 1980 37340
rect 20808 37128 21020 37340
rect 21216 37128 21428 37340
rect 21624 37204 21972 37340
rect 21526 37128 21972 37204
rect 22032 37128 22244 37340
rect 22440 37128 22652 37340
rect 27336 37128 27684 37340
rect 27608 37068 27684 37128
rect 0 36856 13812 36932
rect 13600 36720 13812 36856
rect 14641 36835 15375 36895
rect 20808 36720 21020 36932
rect 21216 36856 21564 36932
rect 21216 36796 21428 36856
rect 21624 36796 21972 36932
rect 21216 36720 21972 36796
rect 22032 36720 22244 36932
rect 22440 36720 22652 36932
rect 27336 36856 27684 37068
rect 109344 37128 109556 37340
rect 114240 37128 114452 37340
rect 114648 37128 114860 37340
rect 115056 37264 115676 37340
rect 115056 37128 115268 37264
rect 115464 37128 115676 37264
rect 115872 37128 116084 37340
rect 134776 37264 134988 37400
rect 109344 37068 109420 37128
rect 109344 36856 109556 37068
rect 27608 36796 27684 36856
rect 109480 36796 109556 36856
rect 20808 36660 20884 36720
rect 14008 36252 14220 36388
rect 20808 36312 21020 36660
rect 27336 36584 27684 36796
rect 109344 36584 109556 36796
rect 114240 36720 114452 36932
rect 114648 36720 114860 36932
rect 115056 36720 115268 36932
rect 115464 36720 115676 36932
rect 115872 36720 116084 36932
rect 116008 36660 116084 36720
rect 27336 36524 27412 36584
rect 109480 36524 109556 36584
rect 21216 36388 21428 36524
rect 21216 36312 21564 36388
rect 21624 36312 21972 36524
rect 22032 36312 22244 36524
rect 22440 36312 22652 36524
rect 27336 36312 27684 36524
rect 109344 36312 109556 36524
rect 114240 36312 114452 36524
rect 114648 36312 114860 36524
rect 115056 36312 115268 36524
rect 115464 36388 115676 36524
rect 115366 36312 115676 36388
rect 115872 36312 116084 36660
rect 27472 36252 27548 36312
rect 109344 36252 109420 36312
rect 14008 36176 14318 36252
rect 0 35904 2116 35980
rect 2040 35844 2116 35904
rect 20808 35904 21020 36116
rect 21216 35980 21428 36116
rect 21526 36040 21972 36116
rect 21216 35904 21564 35980
rect 21624 35904 21972 36040
rect 22032 35904 22244 36116
rect 22440 35904 22652 36116
rect 27336 36040 27684 36252
rect 109344 36040 109556 36252
rect 27472 35980 27548 36040
rect 109480 35980 109556 36040
rect 20808 35844 20884 35904
rect 21624 35844 21700 35904
rect 2040 35768 13812 35844
rect 1773 35708 1871 35709
rect 1224 35632 1980 35708
rect 1768 35496 1980 35632
rect 13600 35496 13812 35768
rect 20808 35632 21020 35844
rect 21352 35768 21700 35844
rect 27336 35768 27684 35980
rect 109344 35768 109556 35980
rect 114240 35904 114452 36116
rect 114648 35904 114860 36116
rect 115056 36040 115404 36116
rect 115056 35980 115268 36040
rect 115464 35980 115676 36116
rect 115056 35904 115676 35980
rect 115872 35904 116084 36116
rect 116008 35844 116084 35904
rect 21352 35708 21428 35768
rect 27608 35708 27684 35768
rect 109480 35708 109556 35768
rect 14641 35565 15295 35625
rect 21216 35572 21428 35708
rect 21526 35632 21972 35708
rect 21216 35496 21564 35572
rect 21624 35496 21972 35632
rect 22032 35496 22244 35708
rect 22440 35496 22652 35708
rect 27336 35496 27684 35708
rect 109344 35496 109556 35708
rect 114240 35496 114452 35708
rect 21216 35436 21292 35496
rect 21488 35436 21564 35496
rect 22032 35436 22108 35496
rect 22576 35436 22652 35496
rect 20808 35224 21020 35436
rect 21216 35224 21428 35436
rect 21488 35360 21972 35436
rect 21624 35224 21972 35360
rect 22032 35088 22244 35436
rect 22440 35088 22652 35436
rect 27462 35300 27560 35496
rect 109344 35300 109448 35496
rect 114376 35436 114452 35496
rect 27336 35224 27684 35300
rect 27608 35164 27684 35224
rect 22032 35028 22108 35088
rect 22576 35028 22652 35088
rect 14008 34680 14220 34892
rect 20808 34816 21020 35028
rect 21216 34816 21972 34892
rect 21216 34680 21428 34816
rect 21624 34680 21972 34816
rect 22032 34680 22244 35028
rect 22440 34680 22652 35028
rect 21352 34620 21428 34680
rect 21760 34620 21836 34680
rect 22168 34620 22244 34680
rect 22576 34620 22652 34680
rect 20808 34408 21020 34620
rect 21216 34408 21428 34620
rect 21624 34408 21972 34620
rect 22032 34408 22244 34620
rect 22440 34408 22652 34620
rect 27336 34544 27684 35164
rect 109344 35224 109556 35300
rect 109344 35164 109420 35224
rect 109344 34544 109556 35164
rect 114240 35088 114452 35436
rect 114648 35496 114860 35708
rect 115056 35496 115268 35708
rect 115464 35496 115676 35708
rect 115872 35632 116084 35844
rect 134776 35572 134988 35844
rect 134776 35496 135396 35572
rect 114648 35436 114724 35496
rect 115056 35436 115132 35496
rect 115464 35436 115540 35496
rect 114648 35088 114860 35436
rect 115056 35360 115676 35436
rect 115056 35224 115268 35360
rect 115464 35224 115676 35360
rect 115872 35224 116084 35436
rect 114240 35028 114316 35088
rect 114784 35028 114860 35088
rect 114240 34680 114452 35028
rect 114648 34680 114860 35028
rect 114240 34620 114316 34680
rect 114784 34620 114860 34680
rect 27608 34484 27684 34544
rect 1224 34029 1844 34076
rect 1224 34000 1871 34029
rect 1773 33931 1871 34000
rect 13600 33940 13812 34076
rect 14641 34007 15215 34067
rect 20808 34000 21020 34212
rect 21216 34000 21428 34212
rect 21624 34000 21972 34212
rect 22032 34000 22244 34212
rect 22440 34000 22652 34212
rect 27336 34000 27684 34484
rect 109344 34000 109556 34484
rect 114240 34408 114452 34620
rect 114648 34408 114860 34620
rect 115056 34680 115268 34892
rect 115464 34680 115676 34892
rect 115872 34816 116084 35028
rect 115056 34620 115132 34680
rect 115600 34620 115676 34680
rect 115056 34408 115268 34620
rect 115464 34408 115676 34620
rect 115872 34408 116084 34620
rect 114240 34000 114452 34212
rect 114648 34000 114860 34212
rect 115056 34076 115268 34212
rect 115056 34000 115404 34076
rect 115464 34000 115676 34212
rect 115872 34000 116084 34212
rect 21624 33940 21700 34000
rect 2040 33864 13812 33940
rect 21352 33864 21700 33940
rect 27336 33940 27412 34000
rect 109344 33940 109420 34000
rect 134776 33940 134988 34076
rect 2040 33804 2116 33864
rect 21352 33804 21428 33864
rect 0 33728 2116 33804
rect 20808 33592 21020 33804
rect 21216 33728 21972 33804
rect 21216 33592 21428 33728
rect 21624 33592 21972 33728
rect 22032 33592 22244 33804
rect 22440 33592 22652 33804
rect 27336 33728 27684 33940
rect 109344 33728 109556 33940
rect 134776 33864 135396 33940
rect 27472 33668 27548 33728
rect 109480 33668 109556 33728
rect 14008 33456 14356 33532
rect 27336 33456 27684 33668
rect 109344 33456 109556 33668
rect 114240 33592 114452 33804
rect 114648 33592 114860 33804
rect 115056 33592 115268 33804
rect 115366 33728 115676 33804
rect 115464 33592 115676 33728
rect 115872 33592 116084 33804
rect 14008 33320 14220 33456
rect 27608 33396 27684 33456
rect 109480 33396 109556 33456
rect 20808 33184 21020 33396
rect 21216 33184 21428 33396
rect 21624 33184 21972 33396
rect 22032 33184 22244 33396
rect 22440 33184 22652 33396
rect 27336 33184 27684 33396
rect 109344 33184 109556 33396
rect 114240 33184 114452 33396
rect 114648 33184 114860 33396
rect 115056 33184 115268 33396
rect 115464 33184 115676 33396
rect 115872 33184 116084 33396
rect 27472 33124 27548 33184
rect 109344 33124 109420 33184
rect 115464 33124 115540 33184
rect 13600 32852 13812 32988
rect 0 32776 13812 32852
rect 14641 32737 15135 32797
rect 20808 32776 21020 32988
rect 21216 32776 21428 32988
rect 21624 32776 21972 32988
rect 22032 32776 22244 32988
rect 22440 32776 22652 32988
rect 27336 32912 27684 33124
rect 109344 32912 109556 33124
rect 115192 33048 115540 33124
rect 115192 32988 115268 33048
rect 27336 32852 27412 32912
rect 109344 32852 109420 32912
rect 21624 32716 21700 32776
rect 21352 32640 21700 32716
rect 27336 32640 27684 32852
rect 109344 32640 109556 32852
rect 114240 32776 114452 32988
rect 114648 32776 114860 32988
rect 115056 32912 115676 32988
rect 115056 32776 115268 32912
rect 115464 32776 115676 32912
rect 115872 32776 116084 32988
rect 21352 32580 21428 32640
rect 27608 32580 27684 32640
rect 109480 32580 109556 32640
rect 1224 32368 1980 32444
rect 20808 32368 21020 32580
rect 21216 32504 21972 32580
rect 21216 32368 21428 32504
rect 21624 32368 21972 32504
rect 22032 32368 22244 32580
rect 22440 32368 22652 32580
rect 27336 32368 27684 32580
rect 109344 32368 109556 32580
rect 114240 32368 114452 32580
rect 114648 32368 114860 32580
rect 115056 32368 115268 32580
rect 115464 32444 115676 32580
rect 115366 32368 115676 32444
rect 115872 32368 116084 32580
rect 1768 32232 1980 32368
rect 27472 32308 27548 32368
rect 109480 32308 109556 32368
rect 14008 31824 14220 32172
rect 20808 31960 21020 32172
rect 21216 31960 21428 32172
rect 21624 31960 21972 32172
rect 22032 31960 22244 32172
rect 22440 31960 22652 32172
rect 27336 32096 27684 32308
rect 109344 32096 109556 32308
rect 134776 32308 134988 32444
rect 134776 32232 135396 32308
rect 27336 32036 27412 32096
rect 109344 32036 109420 32096
rect 20944 31900 21020 31960
rect 20808 31688 21020 31900
rect 27336 31824 27684 32036
rect 109344 31824 109556 32036
rect 114240 31960 114452 32172
rect 114648 31960 114860 32172
rect 115056 32096 115404 32172
rect 115056 32036 115268 32096
rect 115464 32036 115676 32172
rect 115056 31960 115676 32036
rect 115872 31960 116084 32172
rect 115464 31900 115540 31960
rect 115192 31824 115540 31900
rect 115872 31900 115948 31960
rect 27472 31764 27548 31824
rect 109344 31764 109420 31824
rect 115192 31764 115268 31824
rect 21216 31688 21972 31764
rect 21216 31628 21428 31688
rect 21216 31552 21564 31628
rect 21624 31552 21972 31688
rect 22032 31552 22244 31764
rect 22440 31552 22652 31764
rect 21216 31492 21292 31552
rect 21488 31492 21564 31552
rect 13600 31084 13812 31220
rect 14641 31179 15055 31239
rect 0 31008 13812 31084
rect 20808 31144 21020 31492
rect 21216 31144 21428 31492
rect 21488 31416 21972 31492
rect 21624 31144 21972 31416
rect 22032 31144 22244 31356
rect 22440 31144 22652 31356
rect 27336 31280 27684 31764
rect 109344 31280 109556 31764
rect 114240 31552 114452 31764
rect 114648 31552 114860 31764
rect 115056 31688 115676 31764
rect 115872 31688 116084 31900
rect 115056 31628 115268 31688
rect 115056 31552 115404 31628
rect 115464 31552 115676 31688
rect 115192 31492 115268 31552
rect 27608 31220 27684 31280
rect 20808 31084 20884 31144
rect 22032 31084 22108 31144
rect 22440 31084 22516 31144
rect 20808 30872 21020 31084
rect 21216 30736 21428 30948
rect 21624 30812 21972 30948
rect 21488 30736 21972 30812
rect 22032 30736 22244 31084
rect 22440 30736 22652 31084
rect 21216 30676 21292 30736
rect 21488 30676 21564 30736
rect 22168 30676 22244 30736
rect 22576 30676 22652 30736
rect 1768 30540 1980 30676
rect 1224 30464 1980 30540
rect 14008 30464 14220 30676
rect 20808 30464 21020 30676
rect 21216 30600 21564 30676
rect 21216 30540 21428 30600
rect 21624 30540 21972 30676
rect 21216 30464 21972 30540
rect 21352 30404 21428 30464
rect 21352 30328 21700 30404
rect 22032 30328 22244 30676
rect 22440 30328 22652 30676
rect 27336 30600 27684 31220
rect 109344 30600 109556 31220
rect 114240 31144 114452 31356
rect 114648 31144 114860 31356
rect 115056 31144 115268 31492
rect 115328 31492 115404 31552
rect 115328 31416 115676 31492
rect 115464 31144 115676 31416
rect 115872 31144 116084 31492
rect 114376 31084 114452 31144
rect 114784 31084 114860 31144
rect 114240 30736 114452 31084
rect 114648 30736 114860 31084
rect 115872 31084 115948 31144
rect 115056 30812 115268 30948
rect 115056 30736 115404 30812
rect 115464 30736 115676 30948
rect 115872 30872 116084 31084
rect 114240 30676 114316 30736
rect 114648 30676 114724 30736
rect 115192 30676 115268 30736
rect 21624 30268 21700 30328
rect 22168 30268 22244 30328
rect 22576 30268 22652 30328
rect 13600 29996 13812 30132
rect 20808 30056 21020 30268
rect 0 29920 13812 29996
rect 14641 29909 14975 29969
rect 21216 29920 21428 30268
rect 21352 29860 21428 29920
rect 20808 29648 21020 29860
rect 21216 29648 21428 29860
rect 21624 29920 21972 30268
rect 22032 30056 22244 30268
rect 22440 30056 22652 30268
rect 27336 30056 27684 30404
rect 109344 30056 109556 30404
rect 114240 30328 114452 30676
rect 114648 30328 114860 30676
rect 115056 30464 115268 30676
rect 115328 30676 115404 30736
rect 115600 30676 115676 30736
rect 115328 30600 115676 30676
rect 115464 30464 115676 30600
rect 115872 30464 116084 30676
rect 134776 30540 134988 30676
rect 134776 30464 135396 30540
rect 114240 30268 114316 30328
rect 114784 30268 114860 30328
rect 114240 30056 114452 30268
rect 114648 30056 114860 30268
rect 27472 29996 27548 30056
rect 109480 29996 109556 30056
rect 21624 29860 21700 29920
rect 21624 29724 21972 29860
rect 21526 29648 21972 29724
rect 22032 29648 22244 29860
rect 22440 29648 22652 29860
rect 27336 29784 27684 29996
rect 109344 29784 109556 29996
rect 115056 29920 115268 30268
rect 115192 29860 115268 29920
rect 27336 29724 27412 29784
rect 109344 29724 109420 29784
rect 21896 29588 21972 29648
rect 22440 29588 22516 29648
rect 21896 29512 22516 29588
rect 27336 29512 27684 29724
rect 109344 29512 109556 29724
rect 114240 29648 114452 29860
rect 114648 29648 114860 29860
rect 115056 29724 115268 29860
rect 115464 29920 115676 30268
rect 115872 30056 116084 30268
rect 115464 29860 115540 29920
rect 115056 29648 115404 29724
rect 115464 29648 115676 29860
rect 115872 29648 116084 29860
rect 27336 29452 27412 29512
rect 109480 29452 109556 29512
rect 14008 29180 14220 29316
rect 20808 29240 21020 29452
rect 21216 29376 21564 29452
rect 21216 29240 21428 29376
rect 21624 29240 21972 29452
rect 22032 29240 22244 29452
rect 22440 29240 22652 29452
rect 27336 29240 27684 29452
rect 109344 29240 109556 29452
rect 114240 29240 114452 29452
rect 114648 29240 114860 29452
rect 115056 29240 115268 29452
rect 115366 29376 115676 29452
rect 115464 29316 115676 29376
rect 115366 29240 115676 29316
rect 115872 29240 116084 29452
rect 27472 29180 27548 29240
rect 109480 29180 109556 29240
rect 14008 29104 17892 29180
rect 1224 28968 1980 29044
rect 1768 28832 1980 28968
rect 20808 28832 21020 29044
rect 21216 28832 21428 29044
rect 21624 28832 21972 29044
rect 22032 28832 22244 29044
rect 22440 28832 22652 29044
rect 27336 28968 27684 29180
rect 109344 28968 109556 29180
rect 27608 28908 27684 28968
rect 109480 28908 109556 28968
rect 27336 28696 27684 28908
rect 109344 28696 109556 28908
rect 114240 28832 114452 29044
rect 114648 28832 114860 29044
rect 115056 28968 115404 29044
rect 115056 28832 115268 28968
rect 115464 28832 115676 29044
rect 115872 28832 116084 29044
rect 134776 28968 135396 29044
rect 134776 28832 134988 28968
rect 115464 28772 115540 28832
rect 115192 28696 115540 28772
rect 27472 28636 27548 28696
rect 109344 28636 109420 28696
rect 115192 28636 115268 28696
rect 20808 28424 21020 28636
rect 21216 28424 21428 28636
rect 21624 28500 21972 28636
rect 21526 28424 21972 28500
rect 22032 28424 22244 28636
rect 22440 28424 22652 28636
rect 27336 28424 27684 28636
rect 109344 28424 109556 28636
rect 114240 28424 114452 28636
rect 114648 28424 114860 28636
rect 115056 28560 115676 28636
rect 115056 28424 115268 28560
rect 115464 28424 115676 28560
rect 115872 28424 116084 28636
rect 13600 28228 13812 28364
rect 14641 28351 14895 28411
rect 27608 28364 27684 28424
rect 109480 28364 109556 28424
rect 0 28152 13812 28228
rect 20808 28092 21020 28228
rect 14694 28017 14778 28091
rect 18942 28016 21020 28092
rect 21216 28152 21564 28228
rect 21216 28092 21428 28152
rect 21624 28092 21972 28228
rect 21216 28016 21972 28092
rect 22032 28016 22244 28228
rect 22440 28016 22652 28228
rect 27336 28152 27684 28364
rect 109344 28152 109556 28364
rect 27472 28092 27548 28152
rect 109480 28092 109556 28152
rect 20808 27956 20884 28016
rect 14008 27684 14220 27820
rect 14008 27608 15988 27684
rect 20808 27608 21020 27956
rect 27336 27880 27684 28092
rect 109344 27880 109556 28092
rect 114240 28016 114452 28228
rect 114648 28016 114860 28228
rect 115056 28016 115268 28228
rect 115464 28016 115676 28228
rect 115872 28016 116084 28228
rect 115464 27956 115540 28016
rect 116008 27956 116084 28016
rect 27472 27820 27548 27880
rect 109480 27820 109556 27880
rect 115192 27880 115540 27956
rect 115192 27820 115268 27880
rect 20944 27548 21020 27608
rect 1768 27276 1980 27412
rect 1224 27200 1980 27276
rect 17408 27200 17620 27548
rect 17816 27472 18436 27548
rect 17816 27200 18028 27472
rect 18224 27200 18436 27472
rect 18632 27336 18980 27412
rect 18632 27200 18844 27336
rect 19040 27276 19252 27412
rect 19040 27200 20748 27276
rect 20808 27200 21020 27548
rect 21216 27608 21428 27820
rect 21624 27608 21972 27820
rect 22032 27608 22244 27820
rect 22440 27608 22652 27820
rect 21216 27548 21292 27608
rect 21624 27548 21700 27608
rect 21216 27200 21428 27548
rect 21624 27276 21972 27548
rect 21526 27200 21972 27276
rect 22032 27200 22244 27412
rect 20808 27140 20884 27200
rect 22168 27140 22244 27200
rect 20808 26928 21020 27140
rect 21216 26928 21564 27004
rect 21216 26868 21428 26928
rect 18496 26792 19116 26868
rect 20710 26792 21428 26868
rect 21624 26792 21972 27004
rect 22032 26792 22244 27140
rect 22440 27200 22652 27412
rect 27336 27336 27684 27820
rect 109344 27336 109556 27820
rect 114240 27608 114452 27820
rect 114648 27608 114860 27820
rect 115056 27744 115676 27820
rect 115056 27684 115268 27744
rect 115056 27608 115404 27684
rect 115464 27608 115676 27744
rect 115872 27608 116084 27956
rect 115192 27548 115268 27608
rect 27472 27276 27548 27336
rect 109480 27276 109556 27336
rect 22440 27140 22516 27200
rect 22440 26792 22652 27140
rect 18496 26732 18572 26792
rect 19040 26732 19116 26792
rect 21216 26732 21292 26792
rect 21760 26732 21836 26792
rect 22168 26732 22244 26792
rect 22576 26732 22652 26792
rect 17408 26596 17620 26732
rect 17816 26596 18028 26732
rect 18224 26656 18572 26732
rect 18224 26596 18436 26656
rect 17408 26520 17756 26596
rect 17816 26520 18436 26596
rect 17952 26460 18028 26520
rect 17952 26384 18300 26460
rect 18632 26384 18844 26732
rect 19040 26384 19252 26732
rect 20808 26520 21020 26732
rect 21216 26520 21428 26732
rect 21624 26520 21972 26732
rect 22032 26384 22244 26732
rect 22440 26384 22652 26732
rect 27336 26656 27684 27276
rect 109344 26656 109556 27276
rect 114240 27200 114452 27412
rect 114648 27200 114860 27412
rect 115056 27200 115268 27548
rect 115328 27548 115404 27608
rect 115872 27548 115948 27608
rect 115328 27472 115676 27548
rect 115464 27276 115676 27472
rect 115464 27200 115812 27276
rect 115872 27200 116084 27548
rect 117912 27472 118668 27548
rect 117912 27412 117988 27472
rect 117640 27336 117988 27412
rect 117640 27200 117852 27336
rect 118048 27200 118260 27412
rect 118456 27276 118668 27472
rect 118864 27276 119076 27548
rect 118456 27200 119076 27276
rect 119272 27200 119484 27548
rect 134776 27276 134988 27412
rect 134776 27200 135396 27276
rect 114240 27140 114316 27200
rect 114648 27140 114724 27200
rect 116008 27140 116084 27200
rect 114240 26792 114452 27140
rect 114648 26792 114860 27140
rect 115056 26792 115268 27004
rect 115464 26868 115676 27004
rect 115872 26928 116084 27140
rect 114376 26732 114452 26792
rect 114784 26732 114860 26792
rect 115192 26732 115268 26792
rect 115328 26792 115676 26868
rect 115774 26792 117716 26868
rect 115328 26732 115404 26792
rect 18632 26324 18708 26384
rect 22032 26324 22108 26384
rect 22440 26324 22516 26384
rect 17718 26248 18708 26324
rect 20808 26112 21020 26324
rect 3128 25976 4156 26052
rect 3128 25840 3340 25976
rect 3944 25916 4156 25976
rect 18496 25976 19116 26052
rect 21216 25976 21428 26324
rect 21624 26052 21972 26324
rect 22032 26112 22244 26324
rect 22440 26112 22652 26324
rect 27336 26112 27684 26460
rect 109344 26112 109556 26460
rect 114240 26384 114452 26732
rect 114376 26324 114452 26384
rect 114240 26112 114452 26324
rect 114648 26384 114860 26732
rect 115056 26656 115404 26732
rect 115464 26732 115540 26792
rect 115056 26520 115268 26656
rect 115464 26520 115676 26732
rect 115872 26520 116084 26732
rect 117640 26384 117852 26732
rect 118048 26384 118260 26732
rect 118456 26656 118804 26732
rect 118456 26596 118668 26656
rect 118864 26596 119076 26732
rect 118456 26520 119076 26596
rect 119272 26520 119484 26732
rect 114648 26324 114724 26384
rect 114648 26112 114860 26324
rect 27472 26052 27548 26112
rect 109480 26052 109556 26112
rect 18496 25916 18572 25976
rect 19040 25916 19116 25976
rect 21352 25916 21428 25976
rect 21488 25976 21972 26052
rect 21488 25916 21564 25976
rect 3846 25840 4156 25916
rect 17408 25704 17620 25916
rect 17816 25780 18028 25916
rect 18224 25840 18572 25916
rect 18224 25780 18436 25840
rect 17816 25704 18436 25780
rect 18632 25704 18844 25916
rect 19040 25704 19252 25916
rect 20808 25704 21020 25916
rect 21216 25840 21564 25916
rect 21216 25780 21428 25840
rect 21624 25780 21972 25916
rect 21216 25704 21972 25780
rect 22032 25704 22244 25916
rect 22440 25704 22652 25916
rect 27336 25840 27684 26052
rect 109344 25840 109556 26052
rect 115056 25976 115268 26324
rect 115464 25976 115676 26324
rect 115872 26112 116084 26324
rect 115056 25916 115132 25976
rect 115600 25916 115676 25976
rect 118320 25976 119348 26052
rect 118320 25916 118396 25976
rect 119272 25916 119348 25976
rect 27608 25780 27684 25840
rect 109480 25780 109556 25840
rect 21624 25644 21700 25704
rect 1224 25568 1980 25644
rect 1768 25432 1980 25568
rect 21488 25568 21700 25644
rect 21488 25508 21564 25568
rect 2494 25301 2644 25365
rect 20808 25296 21020 25508
rect 21216 25432 21564 25508
rect 21216 25296 21428 25432
rect 21624 25372 21972 25508
rect 21526 25296 21972 25372
rect 22032 25296 22244 25508
rect 22440 25296 22652 25508
rect 27336 25296 27684 25780
rect 109344 25296 109556 25780
rect 114240 25704 114452 25916
rect 114648 25704 114860 25916
rect 115056 25704 115268 25916
rect 115464 25704 115676 25916
rect 115872 25704 116084 25916
rect 117640 25704 117852 25916
rect 118048 25840 118396 25916
rect 118048 25704 118260 25840
rect 118456 25780 118668 25916
rect 118864 25780 119076 25916
rect 118456 25704 119076 25780
rect 119272 25780 119484 25916
rect 119272 25704 120844 25780
rect 134776 25508 134988 25644
rect 114240 25296 114452 25508
rect 114648 25296 114860 25508
rect 115056 25372 115268 25508
rect 115464 25372 115676 25508
rect 115056 25296 115676 25372
rect 115872 25296 116084 25508
rect 134776 25432 135396 25508
rect 27336 25236 27412 25296
rect 109344 25236 109420 25296
rect 17272 25160 17892 25236
rect 17272 25100 17348 25160
rect 17816 25100 17892 25160
rect 15912 24964 16124 25100
rect 16320 25024 17348 25100
rect 15912 24888 16260 24964
rect 16320 24888 16532 25024
rect 17408 24964 17620 25100
rect 17816 24964 18028 25100
rect 18224 24964 18436 25100
rect 17408 24888 17756 24964
rect 17816 24888 18436 24964
rect 18632 24888 18844 25100
rect 19040 24888 19252 25100
rect 20808 24888 21020 25100
rect 21216 25024 21564 25100
rect 21216 24888 21428 25024
rect 21624 24888 21972 25100
rect 22032 24888 22244 25100
rect 22440 24888 22652 25100
rect 27336 25024 27684 25236
rect 109344 25024 109556 25236
rect 119136 25160 120436 25236
rect 119136 25100 119212 25160
rect 120360 25100 120436 25160
rect 27472 24964 27548 25024
rect 109480 24964 109556 25024
rect 16184 24828 16260 24888
rect 17408 24828 17484 24888
rect 16184 24752 17484 24828
rect 27336 24752 27684 24964
rect 109344 24752 109556 24964
rect 114240 24888 114452 25100
rect 114648 24888 114860 25100
rect 115056 24888 115268 25100
rect 115464 24888 115676 25100
rect 115872 24888 116084 25100
rect 117640 24888 117852 25100
rect 118048 24888 118260 25100
rect 118456 24964 118668 25100
rect 118864 25024 119212 25100
rect 118864 24964 119076 25024
rect 118456 24888 119076 24964
rect 119272 24888 119484 25100
rect 120360 24888 120572 25100
rect 120768 24888 120980 25100
rect 27608 24692 27684 24752
rect 109480 24692 109556 24752
rect 3128 24556 3340 24692
rect 3944 24556 4156 24692
rect 2350 24480 4156 24556
rect 20808 24480 21020 24692
rect 21216 24616 21972 24692
rect 21216 24480 21428 24616
rect 21624 24480 21972 24616
rect 22032 24480 22244 24692
rect 22440 24480 22652 24692
rect 27336 24480 27684 24692
rect 27608 24420 27684 24480
rect 20808 24072 21020 24284
rect 21216 24072 21428 24284
rect 21624 24148 21972 24284
rect 21526 24072 21972 24148
rect 22032 24072 22244 24284
rect 22440 24072 22652 24284
rect 27336 24208 27684 24420
rect 109344 24480 109556 24692
rect 114240 24480 114452 24692
rect 114648 24480 114860 24692
rect 115056 24480 115268 24692
rect 115464 24480 115676 24692
rect 115872 24480 116084 24692
rect 109344 24420 109420 24480
rect 115464 24420 115540 24480
rect 109344 24208 109556 24420
rect 115192 24344 115540 24420
rect 115192 24284 115268 24344
rect 27336 24148 27412 24208
rect 109344 24148 109420 24208
rect 20944 24012 21020 24072
rect 1224 23936 2388 24012
rect 1768 23800 1980 23936
rect 20808 23664 21020 24012
rect 21352 23936 21700 24012
rect 27336 23936 27684 24148
rect 109344 23936 109556 24148
rect 114240 24072 114452 24284
rect 114648 24072 114860 24284
rect 115056 24208 115676 24284
rect 115056 24072 115268 24208
rect 115464 24072 115676 24208
rect 115872 24072 116084 24284
rect 21352 23876 21428 23936
rect 21624 23876 21700 23936
rect 27608 23876 27684 23936
rect 109480 23876 109556 23936
rect 115872 24012 115948 24072
rect 21216 23800 21564 23876
rect 21216 23740 21428 23800
rect 21216 23664 21564 23740
rect 21624 23664 21972 23876
rect 22032 23664 22244 23876
rect 22440 23664 22652 23876
rect 20808 23604 20884 23664
rect 21488 23604 21564 23664
rect 18496 23528 19116 23604
rect 18496 23468 18572 23528
rect 19040 23468 19116 23528
rect 3264 23392 4020 23468
rect 17718 23392 18028 23468
rect 3264 23332 3340 23392
rect 3944 23332 4020 23392
rect 17816 23332 18028 23392
rect 18224 23392 18572 23468
rect 3128 23256 3884 23332
rect 3128 23196 3340 23256
rect 544 23120 3884 23196
rect 3944 23120 4156 23332
rect 17816 23256 18164 23332
rect 18224 23256 18436 23392
rect 18632 23256 18844 23468
rect 19040 23256 19252 23468
rect 20808 23256 21020 23604
rect 21216 23256 21428 23604
rect 21488 23528 21972 23604
rect 21624 23256 21972 23528
rect 22032 23256 22244 23468
rect 22440 23256 22652 23468
rect 27336 23392 27684 23876
rect 109344 23392 109556 23876
rect 114240 23664 114452 23876
rect 114648 23664 114860 23876
rect 115056 23664 115268 23876
rect 115464 23664 115676 23876
rect 115872 23664 116084 24012
rect 134776 23876 134988 24012
rect 134776 23800 135396 23876
rect 115056 23604 115132 23664
rect 115600 23604 115676 23664
rect 116008 23604 116084 23664
rect 109344 23332 109420 23392
rect 18088 23196 18164 23256
rect 18632 23196 18708 23256
rect 20944 23196 21020 23256
rect 18088 23120 18708 23196
rect 20808 22984 21020 23196
rect 27336 23120 27684 23332
rect 109344 23120 109556 23332
rect 114240 23256 114452 23468
rect 114648 23256 114860 23468
rect 115056 23256 115268 23604
rect 115464 23256 115676 23604
rect 115872 23256 116084 23604
rect 117640 23256 117852 23468
rect 118048 23256 118260 23468
rect 118456 23256 118668 23468
rect 118864 23256 119076 23468
rect 115464 23196 115540 23256
rect 115192 23120 115540 23196
rect 115872 23196 115948 23256
rect 27472 23060 27548 23120
rect 109344 23060 109420 23120
rect 115192 23060 115268 23120
rect 21216 22984 21564 23060
rect 21216 22924 21428 22984
rect 21624 22924 21972 23060
rect 17680 22848 18300 22924
rect 21216 22848 21972 22924
rect 22032 22848 22244 23060
rect 17680 22788 17756 22848
rect 18224 22788 18300 22848
rect 21352 22788 21428 22848
rect 22168 22788 22244 22848
rect 16592 22516 16804 22788
rect 17000 22712 17756 22788
rect 16592 22440 16940 22516
rect 17000 22440 17212 22712
rect 17816 22516 18028 22788
rect 17816 22440 18164 22516
rect 18224 22440 18436 22788
rect 18632 22440 18844 22788
rect 19040 22440 19252 22788
rect 20808 22576 21020 22788
rect 21216 22576 21428 22788
rect 21526 22712 21972 22788
rect 21624 22576 21972 22712
rect 22032 22440 22244 22788
rect 22440 22848 22652 23060
rect 22440 22788 22516 22848
rect 22440 22440 22652 22788
rect 27336 22712 27684 23060
rect 109344 22712 109556 23060
rect 114240 22848 114452 23060
rect 114648 22848 114860 23060
rect 115056 22984 115676 23060
rect 115872 22984 116084 23196
rect 118358 22984 118940 23060
rect 115056 22924 115268 22984
rect 115056 22848 115404 22924
rect 115464 22848 115676 22984
rect 118728 22848 119756 22924
rect 114240 22788 114316 22848
rect 114648 22788 114724 22848
rect 115056 22788 115132 22848
rect 115328 22788 115404 22848
rect 118728 22788 118804 22848
rect 119680 22788 119756 22848
rect 16864 22380 16940 22440
rect 17816 22380 17892 22440
rect 1224 22304 1980 22380
rect 16864 22304 17892 22380
rect 18088 22380 18164 22440
rect 18632 22380 18708 22440
rect 22032 22380 22108 22440
rect 22576 22380 22652 22440
rect 18088 22304 18708 22380
rect 1768 22244 1980 22304
rect 1768 22168 3204 22244
rect 20808 22168 21020 22380
rect 21216 22032 21428 22380
rect 21624 22108 21972 22380
rect 21488 22032 21972 22108
rect 22032 22032 22244 22380
rect 22440 22032 22652 22380
rect 21216 21972 21292 22032
rect 21488 21972 21564 22032
rect 22032 21972 22108 22032
rect 22576 21972 22652 22032
rect 3128 21700 3340 21836
rect 3944 21700 4156 21836
rect 20808 21760 21020 21972
rect 21216 21896 21564 21972
rect 21216 21760 21428 21896
rect 21624 21836 21972 21972
rect 21526 21760 21972 21836
rect 22032 21760 22244 21972
rect 22440 21760 22652 21972
rect 27336 21896 27684 22516
rect 109344 21896 109556 22516
rect 114240 22440 114452 22788
rect 114648 22440 114860 22788
rect 115056 22576 115268 22788
rect 115328 22712 115676 22788
rect 115464 22576 115676 22712
rect 115872 22576 116084 22788
rect 117640 22516 117852 22788
rect 118048 22712 118396 22788
rect 118456 22712 118804 22788
rect 117640 22440 117988 22516
rect 118048 22440 118260 22712
rect 118456 22440 118668 22712
rect 118864 22516 119076 22788
rect 118864 22440 119620 22516
rect 119680 22440 120028 22788
rect 120088 22440 120300 22788
rect 114376 22380 114452 22440
rect 114784 22380 114860 22440
rect 117912 22380 117988 22440
rect 118456 22380 118532 22440
rect 114240 22032 114452 22380
rect 114648 22032 114860 22380
rect 115056 22032 115268 22380
rect 115464 22108 115676 22380
rect 115872 22168 116084 22380
rect 117912 22304 118532 22380
rect 119544 22380 119620 22440
rect 120088 22380 120164 22440
rect 119544 22304 120164 22380
rect 134776 22244 134988 22380
rect 118358 22168 118940 22244
rect 134776 22168 135396 22244
rect 114240 21972 114316 22032
rect 114648 21972 114724 22032
rect 115192 21972 115268 22032
rect 115328 22032 115676 22108
rect 115328 21972 115404 22032
rect 27472 21836 27548 21896
rect 109344 21836 109420 21896
rect 3128 21624 4156 21700
rect 20808 21352 21020 21564
rect 21216 21488 21564 21564
rect 21216 21352 21428 21488
rect 21624 21352 21972 21564
rect 22032 21352 22244 21564
rect 22440 21352 22652 21564
rect 27336 21352 27684 21836
rect 27608 21292 27684 21352
rect 18088 21216 18708 21292
rect 18088 21156 18164 21216
rect 18632 21156 18708 21216
rect 17816 21080 18164 21156
rect 17816 20944 18028 21080
rect 18224 21020 18436 21156
rect 18224 20944 18572 21020
rect 18632 20944 18844 21156
rect 19040 20944 19252 21156
rect 20808 20944 21020 21156
rect 21216 20944 21428 21156
rect 21624 20944 21972 21156
rect 22032 20944 22244 21156
rect 22440 20944 22652 21156
rect 27336 21080 27684 21292
rect 109344 21352 109556 21836
rect 114240 21760 114452 21972
rect 114648 21760 114860 21972
rect 115056 21896 115404 21972
rect 115056 21836 115268 21896
rect 115464 21836 115676 21972
rect 115056 21760 115676 21836
rect 115872 21760 116084 21972
rect 114240 21352 114452 21564
rect 114648 21352 114860 21564
rect 115056 21352 115268 21564
rect 115464 21352 115676 21564
rect 115872 21428 116084 21564
rect 115872 21352 118124 21428
rect 109344 21292 109420 21352
rect 109344 21080 109556 21292
rect 117912 21216 118532 21292
rect 117912 21156 117988 21216
rect 27336 21020 27412 21080
rect 109344 21020 109420 21080
rect 18496 20884 18572 20944
rect 19040 20884 19116 20944
rect 18496 20808 19116 20884
rect 27336 20808 27684 21020
rect 109344 20808 109556 21020
rect 114240 20944 114452 21156
rect 114648 20944 114860 21156
rect 115056 21080 115676 21156
rect 115056 21020 115268 21080
rect 115056 20944 115404 21020
rect 115464 20944 115676 21080
rect 115872 20944 116084 21156
rect 117640 21080 117988 21156
rect 118048 21080 118396 21156
rect 117640 21020 117852 21080
rect 117640 20944 117988 21020
rect 118048 20944 118260 21080
rect 118456 20944 118668 21156
rect 118864 20944 119076 21156
rect 117912 20884 117988 20944
rect 118456 20884 118532 20944
rect 117912 20808 118532 20884
rect 27336 20748 27412 20808
rect 109344 20748 109420 20808
rect 1224 20536 1980 20612
rect 20808 20536 21020 20748
rect 21216 20672 21972 20748
rect 21216 20536 21428 20672
rect 21624 20536 21972 20672
rect 22032 20536 22244 20748
rect 22440 20536 22652 20748
rect 27336 20536 27684 20748
rect 109344 20536 109556 20748
rect 114240 20536 114452 20748
rect 114648 20536 114860 20748
rect 115056 20536 115268 20748
rect 115366 20672 115676 20748
rect 115464 20536 115676 20672
rect 115872 20536 116084 20748
rect 134776 20536 135396 20612
rect 1768 20400 1980 20536
rect 27472 20476 27548 20536
rect 109480 20476 109556 20536
rect 3128 20400 3748 20476
rect 3846 20400 4156 20476
rect 3128 20340 3340 20400
rect 3944 20340 4156 20400
rect 17680 20400 18300 20476
rect 17680 20340 17756 20400
rect 18224 20340 18300 20400
rect 3128 20264 4156 20340
rect 16592 20204 16804 20340
rect 17000 20264 17756 20340
rect 16592 20128 16940 20204
rect 17000 20128 17212 20264
rect 17816 20128 18028 20340
rect 18224 20128 18436 20340
rect 18632 20128 18844 20340
rect 19040 20128 19252 20340
rect 20808 20204 21020 20340
rect 20808 20128 21156 20204
rect 21216 20128 21428 20340
rect 21624 20128 21972 20340
rect 22032 20128 22244 20340
rect 22440 20128 22652 20340
rect 27336 20264 27684 20476
rect 109344 20264 109556 20476
rect 118728 20400 119756 20476
rect 134776 20400 134988 20536
rect 118728 20340 118804 20400
rect 119680 20340 119756 20400
rect 27608 20204 27684 20264
rect 109480 20204 109556 20264
rect 16864 20068 16940 20128
rect 17816 20068 17892 20128
rect 16864 19992 17892 20068
rect 27336 19992 27684 20204
rect 109344 20068 109556 20204
rect 114240 20128 114452 20340
rect 114648 20128 114860 20340
rect 115056 20128 115268 20340
rect 115464 20128 115676 20340
rect 115872 20128 116084 20340
rect 117640 20128 117852 20340
rect 118048 20204 118260 20340
rect 118456 20264 118804 20340
rect 118048 20128 118396 20204
rect 118456 20128 118668 20264
rect 118864 20204 119076 20340
rect 118864 20128 119620 20204
rect 119680 20128 120028 20340
rect 120088 20204 120300 20340
rect 120088 20128 122884 20204
rect 118320 20068 118396 20128
rect 118864 20068 118940 20128
rect 109344 19992 109692 20068
rect 118320 19992 118940 20068
rect 119544 20068 119620 20128
rect 120088 20068 120164 20128
rect 119544 19992 120164 20068
rect 27472 19932 27548 19992
rect 109344 19932 109420 19992
rect 27336 19796 27684 19932
rect 22440 19660 22652 19796
rect 23256 19660 23604 19796
rect 25976 19660 26188 19796
rect 27064 19720 29044 19796
rect 109344 19720 109556 19932
rect 22440 19584 27004 19660
rect 27064 19584 27276 19720
rect 109616 19584 109828 19796
rect 122808 19720 123020 19932
rect 122216 19501 122300 19575
rect 26966 19312 28908 19388
rect 28152 19252 28364 19312
rect 28696 19252 28908 19312
rect 29376 19312 30812 19388
rect 29376 19252 29588 19312
rect 28152 19176 28636 19252
rect 28696 19176 29588 19252
rect 29920 19176 30132 19312
rect 30600 19252 30812 19312
rect 31144 19312 32716 19388
rect 31144 19252 31492 19312
rect 30600 19176 31492 19252
rect 31824 19176 32036 19312
rect 32504 19252 32716 19312
rect 33048 19252 33260 19388
rect 32504 19176 33260 19252
rect 33728 19312 34620 19388
rect 33728 19176 33940 19312
rect 34272 19252 34620 19312
rect 34952 19252 35164 19388
rect 35632 19312 37748 19388
rect 35632 19252 35844 19312
rect 34272 19176 35844 19252
rect 36176 19176 36388 19312
rect 36856 19252 37068 19312
rect 37400 19252 37748 19312
rect 38080 19252 38292 19388
rect 36856 19176 37340 19252
rect 37400 19176 38292 19252
rect 38760 19252 38972 19388
rect 39304 19252 39516 19388
rect 38760 19176 39516 19252
rect 39984 19312 40740 19388
rect 39984 19176 40196 19312
rect 40528 19176 40740 19312
rect 41208 19252 41420 19388
rect 41752 19252 42100 19388
rect 41208 19176 42100 19252
rect 42432 19312 43324 19388
rect 42432 19176 42644 19312
rect 43112 19176 43324 19312
rect 43656 19252 43868 19388
rect 44336 19312 45228 19388
rect 44336 19252 44548 19312
rect 43422 19176 44548 19252
rect 44880 19252 45228 19312
rect 45560 19252 45772 19388
rect 46240 19312 46996 19388
rect 46240 19252 46452 19312
rect 44880 19176 46452 19252
rect 46784 19176 46996 19312
rect 47464 19252 47676 19388
rect 48008 19252 48356 19388
rect 48688 19312 49580 19388
rect 48688 19252 48900 19312
rect 47464 19176 48900 19252
rect 49368 19252 49580 19312
rect 49912 19252 50124 19388
rect 50592 19312 52028 19388
rect 50592 19252 50804 19312
rect 49368 19176 50804 19252
rect 51136 19176 51348 19312
rect 51816 19252 52028 19312
rect 52360 19252 52708 19388
rect 53040 19252 53252 19388
rect 51816 19176 53252 19252
rect 53720 19252 53932 19388
rect 54264 19252 54476 19388
rect 53720 19176 54476 19252
rect 54944 19312 55836 19388
rect 54944 19176 55156 19312
rect 55488 19176 55836 19312
rect 56168 19252 56380 19388
rect 56848 19312 58284 19388
rect 56848 19252 57060 19312
rect 56168 19176 57060 19252
rect 57392 19176 57604 19312
rect 58072 19252 58284 19312
rect 58616 19312 59508 19388
rect 58616 19252 58964 19312
rect 58072 19176 58964 19252
rect 59296 19176 59508 19312
rect 59976 19252 60188 19388
rect 60520 19252 60732 19388
rect 61200 19312 61956 19388
rect 61200 19252 61412 19312
rect 59976 19176 60732 19252
rect 60830 19176 61412 19252
rect 61744 19176 61956 19312
rect 62424 19252 62636 19388
rect 62968 19312 64540 19388
rect 62968 19252 63316 19312
rect 62424 19176 63316 19252
rect 63648 19176 63860 19312
rect 64328 19252 64540 19312
rect 64872 19252 65084 19388
rect 65552 19312 66444 19388
rect 65552 19252 65764 19312
rect 64328 19176 65764 19252
rect 66096 19176 66444 19312
rect 66776 19176 66988 19388
rect 67456 19312 68892 19388
rect 67456 19176 67668 19312
rect 68000 19176 68212 19312
rect 68680 19252 68892 19312
rect 69224 19252 69572 19388
rect 69904 19312 71340 19388
rect 69904 19252 70116 19312
rect 68680 19176 70116 19252
rect 70584 19252 70796 19312
rect 71128 19252 71340 19312
rect 71808 19252 72020 19388
rect 70584 19176 71068 19252
rect 71128 19176 72020 19252
rect 72352 19312 73244 19388
rect 72352 19176 72564 19312
rect 73032 19252 73244 19312
rect 73576 19252 73924 19388
rect 74256 19312 75148 19388
rect 74256 19252 74468 19312
rect 73032 19176 74468 19252
rect 74936 19252 75148 19312
rect 75480 19252 75692 19388
rect 74936 19176 75692 19252
rect 76160 19312 77596 19388
rect 76160 19176 76372 19312
rect 76704 19176 77052 19312
rect 77384 19252 77596 19312
rect 78064 19312 80724 19388
rect 78064 19252 78276 19312
rect 77384 19176 78276 19252
rect 78608 19176 78820 19312
rect 79288 19252 79500 19312
rect 79288 19176 79772 19252
rect 79832 19176 80180 19312
rect 80512 19176 80724 19312
rect 81192 19252 81404 19388
rect 81736 19252 81948 19388
rect 82416 19312 83852 19388
rect 82416 19252 82628 19312
rect 81192 19176 82628 19252
rect 82960 19176 83172 19312
rect 83640 19252 83852 19312
rect 84184 19252 84532 19388
rect 83640 19176 84532 19252
rect 84864 19312 85756 19388
rect 84864 19176 85076 19312
rect 85544 19252 85756 19312
rect 86088 19252 86300 19388
rect 86768 19252 86980 19388
rect 85544 19176 86980 19252
rect 87312 19312 88204 19388
rect 87312 19176 87660 19312
rect 87992 19176 88204 19312
rect 88672 19312 89428 19388
rect 88672 19252 88884 19312
rect 88302 19176 88884 19252
rect 89216 19176 89428 19312
rect 89896 19252 90108 19388
rect 90440 19252 90788 19388
rect 91120 19312 92012 19388
rect 91120 19252 91332 19312
rect 89896 19176 91332 19252
rect 91800 19176 92012 19312
rect 92344 19252 92556 19388
rect 93024 19312 94460 19388
rect 94558 19312 95140 19388
rect 93024 19252 93236 19312
rect 92344 19176 93508 19252
rect 93568 19176 93780 19312
rect 94248 19252 94460 19312
rect 94792 19252 95140 19312
rect 95472 19252 95684 19388
rect 94248 19176 95684 19252
rect 96152 19252 96364 19388
rect 96696 19252 96908 19388
rect 97376 19312 98268 19388
rect 97376 19252 97588 19312
rect 96152 19176 97588 19252
rect 97920 19176 98268 19312
rect 98600 19252 98812 19388
rect 99280 19312 100716 19388
rect 99280 19252 99492 19312
rect 98600 19176 99492 19252
rect 99824 19176 100036 19312
rect 100504 19252 100716 19312
rect 101048 19252 101396 19388
rect 101728 19252 101940 19388
rect 100504 19176 101940 19252
rect 102408 19252 102620 19388
rect 102952 19252 103164 19388
rect 103632 19312 104388 19388
rect 103632 19252 103844 19312
rect 102408 19176 103844 19252
rect 104176 19176 104388 19312
rect 104856 19252 105068 19388
rect 105400 19252 105748 19388
rect 106080 19312 106972 19388
rect 106080 19252 106292 19312
rect 104856 19176 105748 19252
rect 105846 19176 106292 19252
rect 106760 19252 106972 19312
rect 107304 19252 107516 19388
rect 107984 19312 108876 19388
rect 107984 19252 108196 19312
rect 106760 19176 107244 19252
rect 107304 19176 108196 19252
rect 108528 19176 108876 19312
rect 123216 19312 136620 19388
rect 122015 19181 122353 19241
rect 123216 19176 123428 19312
rect 3128 19040 4156 19116
rect 1768 18844 1980 18980
rect 3128 18844 3340 19040
rect 1224 18768 3340 18844
rect 3944 18768 4156 19040
rect 14552 19040 16668 19116
rect 14552 18768 14764 19040
rect 134776 18904 135396 18980
rect 28152 18632 28500 18844
rect 28560 18632 28772 18844
rect 29512 18708 29724 18844
rect 29784 18708 30132 18844
rect 29512 18632 30132 18708
rect 30736 18768 31356 18844
rect 30736 18632 30948 18768
rect 31144 18632 31356 18768
rect 31960 18708 32172 18844
rect 32368 18708 32580 18844
rect 31960 18632 32580 18708
rect 33184 18768 33804 18844
rect 33184 18632 33396 18768
rect 33592 18632 33804 18768
rect 34408 18708 34620 18844
rect 34816 18708 35028 18844
rect 34408 18632 35028 18708
rect 35632 18768 36252 18844
rect 35632 18632 35980 18768
rect 36040 18632 36252 18768
rect 36992 18768 37612 18844
rect 36992 18632 37204 18768
rect 37264 18632 37612 18768
rect 38216 18708 38428 18844
rect 38624 18708 38836 18844
rect 38216 18632 38836 18708
rect 39440 18768 40060 18844
rect 39440 18632 39652 18768
rect 39848 18632 40060 18768
rect 40664 18708 40876 18844
rect 41072 18708 41284 18844
rect 40664 18632 41284 18708
rect 41888 18768 42508 18844
rect 41888 18632 42236 18768
rect 42296 18632 42508 18768
rect 43248 18768 43868 18844
rect 43248 18632 43460 18768
rect 43520 18632 43868 18768
rect 44472 18708 44684 18844
rect 44880 18708 45092 18844
rect 44472 18632 45092 18708
rect 45696 18768 46316 18844
rect 45696 18632 45908 18768
rect 46104 18632 46316 18768
rect 46920 18708 47132 18844
rect 47328 18708 47540 18844
rect 46920 18632 47540 18708
rect 48144 18768 48764 18844
rect 48144 18632 48356 18768
rect 48552 18632 48764 18768
rect 49368 18708 49716 18844
rect 49776 18708 49988 18844
rect 49368 18632 49988 18708
rect 50728 18708 50940 18844
rect 51000 18708 51348 18844
rect 50728 18632 51348 18708
rect 51952 18768 52572 18844
rect 51952 18632 52164 18768
rect 52360 18632 52572 18768
rect 53176 18708 53388 18844
rect 53584 18708 53796 18844
rect 53176 18632 53796 18708
rect 54400 18768 55020 18844
rect 54400 18632 54612 18768
rect 54808 18632 55020 18768
rect 55624 18708 55836 18844
rect 56032 18708 56244 18844
rect 55624 18632 56244 18708
rect 56848 18768 57468 18844
rect 56848 18632 57196 18768
rect 57256 18632 57468 18768
rect 58208 18768 58828 18844
rect 58208 18632 58420 18768
rect 58480 18632 58828 18768
rect 59432 18708 59644 18844
rect 59840 18708 60052 18844
rect 59432 18632 60052 18708
rect 60656 18768 61276 18844
rect 60656 18632 60868 18768
rect 61064 18632 61276 18768
rect 61880 18708 62092 18844
rect 62288 18708 62500 18844
rect 61880 18632 62500 18708
rect 63104 18708 63452 18844
rect 63512 18708 63724 18844
rect 63104 18632 63724 18708
rect 64464 18768 65084 18844
rect 64464 18632 64676 18768
rect 64736 18632 65084 18768
rect 65688 18708 65900 18844
rect 66096 18768 67532 18844
rect 66096 18708 66308 18768
rect 65688 18632 66308 18708
rect 66912 18632 67124 18768
rect 67320 18632 67532 18768
rect 68136 18708 68348 18844
rect 68544 18708 68756 18844
rect 68136 18632 68756 18708
rect 69360 18768 69980 18844
rect 69360 18632 69572 18768
rect 69768 18632 69980 18768
rect 70584 18708 70932 18844
rect 70992 18708 71204 18844
rect 70584 18632 71204 18708
rect 71944 18708 72156 18844
rect 72216 18708 72564 18844
rect 71944 18632 72564 18708
rect 73168 18768 73788 18844
rect 73168 18632 73380 18768
rect 73576 18632 73788 18768
rect 74392 18708 74604 18844
rect 74800 18708 75012 18844
rect 74392 18632 75012 18708
rect 75616 18768 76236 18844
rect 75616 18632 75828 18768
rect 76024 18632 76236 18768
rect 76840 18708 77052 18844
rect 77248 18708 77460 18844
rect 76840 18632 77460 18708
rect 78064 18768 78684 18844
rect 78064 18632 78412 18768
rect 78472 18632 78684 18768
rect 79424 18768 80044 18844
rect 79424 18632 79636 18768
rect 79696 18632 80044 18768
rect 80648 18708 80860 18844
rect 81056 18708 81268 18844
rect 80648 18632 81268 18708
rect 81872 18768 82492 18844
rect 81872 18632 82084 18768
rect 82280 18632 82492 18768
rect 83096 18708 83308 18844
rect 83504 18708 83716 18844
rect 83096 18632 83716 18708
rect 84320 18708 84668 18844
rect 84728 18708 84940 18844
rect 84320 18632 84940 18708
rect 85680 18768 86300 18844
rect 85680 18632 85892 18768
rect 85952 18632 86300 18768
rect 86904 18708 87116 18844
rect 87312 18708 87524 18844
rect 86904 18632 87524 18708
rect 88128 18768 88748 18844
rect 88128 18632 88340 18768
rect 88536 18632 88748 18768
rect 89352 18708 89564 18844
rect 89760 18708 89972 18844
rect 89352 18632 89972 18708
rect 90576 18768 91196 18844
rect 90576 18632 90788 18768
rect 90984 18632 91196 18768
rect 91800 18708 92148 18844
rect 92208 18708 92420 18844
rect 91800 18632 92420 18708
rect 93160 18708 93372 18844
rect 93432 18708 93780 18844
rect 93160 18632 93780 18708
rect 94384 18768 95004 18844
rect 94384 18632 94596 18768
rect 94792 18632 95004 18768
rect 95608 18708 95820 18844
rect 96016 18708 96228 18844
rect 95608 18632 96228 18708
rect 96832 18768 97452 18844
rect 96832 18632 97044 18768
rect 97240 18632 97452 18768
rect 98056 18708 98268 18844
rect 98464 18708 98676 18844
rect 98056 18632 98676 18708
rect 99280 18708 99628 18844
rect 99688 18708 99900 18844
rect 99280 18632 99900 18708
rect 100640 18768 101260 18844
rect 100640 18632 100852 18768
rect 100912 18632 101260 18768
rect 101864 18708 102076 18844
rect 102272 18708 102484 18844
rect 101864 18632 102484 18708
rect 103088 18768 103708 18844
rect 103088 18632 103300 18768
rect 103496 18632 103708 18768
rect 104312 18708 104524 18844
rect 104720 18708 104932 18844
rect 104312 18632 104932 18708
rect 105536 18768 106156 18844
rect 105536 18632 105884 18768
rect 105944 18632 106156 18768
rect 106896 18768 107516 18844
rect 106896 18632 107108 18768
rect 107168 18632 107516 18768
rect 108120 18768 108604 18844
rect 134776 18768 134988 18904
rect 108120 18632 108332 18768
rect 119990 18496 123020 18572
rect 122808 18360 123020 18496
rect 14694 18195 22836 18255
rect 2569 17896 28439 17956
rect 121935 17623 122353 17683
rect 123216 17680 136620 17756
rect 3128 17484 3340 17620
rect 3710 17544 4156 17620
rect 3944 17484 4156 17544
rect 3128 17408 4156 17484
rect 14552 17544 17076 17620
rect 14552 17408 14764 17544
rect 123216 17408 123428 17680
rect 1768 17076 1980 17348
rect 20128 17272 21564 17348
rect 20128 17136 20340 17272
rect 21216 17136 21564 17272
rect 134776 17212 134988 17348
rect 28968 17136 30540 17212
rect 1224 17000 1980 17076
rect 28968 17000 29316 17136
rect 30328 17076 30540 17136
rect 31552 17136 32988 17212
rect 31552 17076 31764 17136
rect 30328 17000 31764 17076
rect 32776 17076 32988 17136
rect 34000 17136 35436 17212
rect 34000 17076 34212 17136
rect 32776 17000 34212 17076
rect 35224 17076 35436 17136
rect 36448 17076 36796 17212
rect 37808 17136 39244 17212
rect 37808 17076 38020 17136
rect 35224 17000 38020 17076
rect 39032 17076 39244 17136
rect 40256 17136 41692 17212
rect 40256 17076 40468 17136
rect 39032 17000 40468 17076
rect 41480 17076 41692 17136
rect 42704 17076 43052 17212
rect 44064 17136 45500 17212
rect 44064 17076 44276 17136
rect 41480 17000 44276 17076
rect 45288 17076 45500 17136
rect 46512 17136 47948 17212
rect 46512 17076 46724 17136
rect 45288 17000 46724 17076
rect 47736 17076 47948 17136
rect 48960 17136 50532 17212
rect 48960 17076 49172 17136
rect 47736 17000 49172 17076
rect 50184 17076 50532 17136
rect 51544 17076 51756 17212
rect 52768 17136 54204 17212
rect 52768 17076 52980 17136
rect 50184 17000 52980 17076
rect 53992 17076 54204 17136
rect 55216 17136 56652 17212
rect 55216 17076 55428 17136
rect 53992 17000 55428 17076
rect 56440 17076 56652 17136
rect 57664 17136 60460 17212
rect 57664 17076 58012 17136
rect 56440 17000 58012 17076
rect 59024 17000 59236 17136
rect 60248 17076 60460 17136
rect 61472 17136 62908 17212
rect 61472 17076 61684 17136
rect 60248 17000 61684 17076
rect 62696 17076 62908 17136
rect 63920 17076 64268 17212
rect 65280 17136 66716 17212
rect 65280 17076 65492 17136
rect 62696 17000 65492 17076
rect 66504 17076 66716 17136
rect 67728 17136 69164 17212
rect 67728 17076 67940 17136
rect 66504 17000 67940 17076
rect 68952 17076 69164 17136
rect 70176 17136 71748 17212
rect 70176 17076 70388 17136
rect 68952 17000 70388 17076
rect 71400 17076 71748 17136
rect 72760 17076 72972 17212
rect 73984 17136 75420 17212
rect 73984 17076 74196 17136
rect 71400 17000 74196 17076
rect 75208 17076 75420 17136
rect 76432 17136 77868 17212
rect 76432 17076 76644 17136
rect 75208 17000 76644 17076
rect 77656 17076 77868 17136
rect 78880 17136 81676 17212
rect 78880 17076 79228 17136
rect 77656 17000 79228 17076
rect 80240 17000 80452 17136
rect 81464 17076 81676 17136
rect 82688 17136 84124 17212
rect 82688 17076 82900 17136
rect 81464 17000 82900 17076
rect 83912 17076 84124 17136
rect 85136 17136 87932 17212
rect 85136 17076 85484 17136
rect 86496 17076 86708 17136
rect 83912 17000 85484 17076
rect 86398 17000 86708 17076
rect 87720 17076 87932 17136
rect 88944 17136 90380 17212
rect 88944 17076 89156 17136
rect 87720 17000 89156 17076
rect 90168 17076 90380 17136
rect 91392 17136 92964 17212
rect 91392 17076 91604 17136
rect 90168 17000 91604 17076
rect 92616 17076 92964 17136
rect 93976 17076 94188 17212
rect 95200 17136 96636 17212
rect 95200 17076 95412 17136
rect 92616 17000 95412 17076
rect 96424 17076 96636 17136
rect 97648 17136 99084 17212
rect 97648 17076 97860 17136
rect 96424 17000 97860 17076
rect 98872 17076 99084 17136
rect 100096 17136 102892 17212
rect 100096 17076 100444 17136
rect 98872 17000 100444 17076
rect 101456 17000 101668 17136
rect 102680 17076 102892 17136
rect 103904 17136 105340 17212
rect 103904 17076 104116 17136
rect 102680 17000 104116 17076
rect 105128 17076 105340 17136
rect 106352 17136 107924 17212
rect 106352 17076 106700 17136
rect 105128 17000 106700 17076
rect 107712 17000 107924 17136
rect 134776 17136 135396 17212
rect 122808 16864 123020 17076
rect 134776 17000 134988 17136
rect 121855 16353 122353 16413
rect 123216 16396 123428 16532
rect 123216 16320 136620 16396
rect 3128 16184 4156 16260
rect 3128 16048 3340 16184
rect 3944 16048 4156 16184
rect 14552 16048 14764 16260
rect 20128 15912 21564 15988
rect 20128 15776 20340 15912
rect 21216 15852 21564 15912
rect 21216 15776 22516 15852
rect 1224 15504 3204 15580
rect 122808 15504 123020 15716
rect 1768 15368 1980 15504
rect 134776 15444 134988 15580
rect 14694 15367 26539 15427
rect 134776 15368 135396 15444
rect 28921 15172 29019 15197
rect 31417 15172 31515 15197
rect 33913 15172 34011 15197
rect 36409 15172 36507 15197
rect 38905 15172 39003 15197
rect 41401 15172 41499 15197
rect 43897 15172 43995 15197
rect 46393 15172 46491 15197
rect 48889 15172 48987 15197
rect 51385 15172 51483 15197
rect 53881 15172 53979 15197
rect 56377 15172 56475 15197
rect 58873 15172 58971 15197
rect 61369 15172 61467 15197
rect 63865 15172 63963 15197
rect 66361 15172 66459 15197
rect 68857 15172 68955 15197
rect 71353 15172 71451 15197
rect 73849 15172 73947 15197
rect 76345 15172 76443 15197
rect 78841 15172 78939 15197
rect 81337 15172 81435 15197
rect 83833 15172 83931 15197
rect 86329 15172 86427 15197
rect 88825 15172 88923 15197
rect 91321 15172 91419 15197
rect 93817 15172 93915 15197
rect 96313 15172 96411 15197
rect 98809 15172 98907 15197
rect 101305 15172 101403 15197
rect 103801 15172 103899 15197
rect 106297 15172 106395 15197
rect 28832 15096 29142 15172
rect 31416 15096 31764 15172
rect 33864 15096 34174 15172
rect 36312 15096 36622 15172
rect 38896 15096 39244 15172
rect 41344 15096 41692 15172
rect 43792 15096 44102 15172
rect 46376 15096 46724 15172
rect 48824 15096 49134 15172
rect 51272 15096 51582 15172
rect 53856 15096 54204 15172
rect 56304 15096 56614 15172
rect 58752 15096 59236 15172
rect 61336 15096 61684 15172
rect 63784 15096 64094 15172
rect 66232 15096 66716 15172
rect 68816 15096 69164 15172
rect 71264 15096 71574 15172
rect 73848 15096 74196 15172
rect 76296 15096 76606 15172
rect 78744 15096 79054 15172
rect 81328 15096 81676 15172
rect 83776 15096 84086 15172
rect 86224 15096 86534 15172
rect 88808 15096 89156 15172
rect 91256 15096 91566 15172
rect 93704 15096 94014 15172
rect 96288 15096 96636 15172
rect 98736 15096 99046 15172
rect 101184 15096 101668 15172
rect 103768 15096 104116 15172
rect 106216 15096 106526 15172
rect 121775 14795 122353 14855
rect 123216 14824 136620 14900
rect 544 14688 3340 14764
rect 3128 14628 3340 14688
rect 3944 14628 4156 14764
rect 3128 14552 4156 14628
rect 14552 14552 14764 14764
rect 123216 14688 123428 14824
rect 20128 14356 20340 14628
rect 21216 14356 21564 14628
rect 20128 14280 21564 14356
rect 28832 14280 29044 14492
rect 31280 14280 31492 14492
rect 33728 14356 33940 14492
rect 33630 14280 33940 14356
rect 36312 14280 36524 14492
rect 38760 14356 38972 14492
rect 38760 14280 41148 14356
rect 41208 14280 41420 14492
rect 43792 14280 44004 14492
rect 46240 14280 46452 14492
rect 48688 14280 49036 14492
rect 51272 14280 51484 14492
rect 53720 14356 53932 14492
rect 56168 14356 56516 14492
rect 58382 14416 58964 14492
rect 58752 14356 58964 14416
rect 61200 14356 61412 14492
rect 53720 14280 56516 14356
rect 58654 14280 58964 14356
rect 61102 14280 61412 14356
rect 63648 14280 63996 14492
rect 66232 14280 66444 14492
rect 68680 14280 68892 14492
rect 71264 14280 71476 14492
rect 73712 14280 73924 14492
rect 76160 14356 76372 14492
rect 76062 14280 76372 14356
rect 78744 14280 78956 14492
rect 81192 14280 81404 14492
rect 83640 14280 83852 14492
rect 86224 14356 86436 14492
rect 86126 14280 86436 14356
rect 88672 14280 88884 14492
rect 91120 14280 91468 14492
rect 93704 14280 93916 14492
rect 96152 14356 96364 14492
rect 98600 14416 101396 14492
rect 98600 14356 98948 14416
rect 96152 14280 98948 14356
rect 101184 14280 101396 14416
rect 103632 14416 106428 14492
rect 103632 14356 103844 14416
rect 103534 14280 103844 14356
rect 106080 14280 106428 14416
rect 14694 13953 26787 14013
rect 122808 14008 123020 14356
rect 1224 13872 1980 13948
rect 134776 13872 135396 13948
rect 1768 13812 1980 13872
rect 1768 13736 3204 13812
rect 134823 13771 134921 13872
rect 28832 13600 29044 13676
rect 28851 13487 29044 13600
rect 28968 13464 29044 13487
rect 31280 13600 33668 13676
rect 33728 13600 34076 13676
rect 36312 13600 36524 13676
rect 38760 13600 38972 13676
rect 41110 13600 41556 13676
rect 43792 13600 44004 13676
rect 46240 13600 49036 13676
rect 51272 13600 51484 13676
rect 53720 13600 53932 13676
rect 31280 13464 31492 13600
rect 33843 13487 34076 13600
rect 36339 13487 36524 13600
rect 38835 13487 38972 13600
rect 41331 13487 41556 13600
rect 43827 13487 44004 13600
rect 46323 13487 46452 13600
rect 48819 13487 49036 13600
rect 51315 13487 51484 13600
rect 53811 13487 53932 13600
rect 34000 13464 34076 13487
rect 36448 13464 36524 13487
rect 38896 13464 38972 13487
rect 41344 13464 41556 13487
rect 43928 13464 44004 13487
rect 46376 13464 46452 13487
rect 48960 13464 49036 13487
rect 51408 13464 51484 13487
rect 53856 13464 53932 13487
rect 56304 13600 58692 13676
rect 58752 13600 61140 13676
rect 61200 13600 63724 13676
rect 63784 13600 63996 13676
rect 66232 13600 66444 13676
rect 68680 13600 68892 13676
rect 71264 13600 71476 13676
rect 73712 13600 76100 13676
rect 76160 13600 76508 13676
rect 78744 13600 78956 13676
rect 81192 13600 81404 13676
rect 83640 13600 86164 13676
rect 86224 13600 86436 13676
rect 88672 13600 88884 13676
rect 91120 13600 91468 13676
rect 93704 13600 93916 13676
rect 96152 13600 96364 13676
rect 98736 13600 98948 13676
rect 101184 13600 103572 13676
rect 103632 13600 103844 13676
rect 106216 13600 106428 13676
rect 56304 13464 56516 13600
rect 58803 13487 58964 13600
rect 61299 13487 61397 13600
rect 63795 13487 63996 13600
rect 66291 13487 66444 13600
rect 68787 13487 68885 13600
rect 71283 13487 71476 13600
rect 73779 13487 73924 13600
rect 76275 13487 76508 13600
rect 78771 13487 78956 13600
rect 81267 13487 81404 13600
rect 83763 13487 83988 13600
rect 86259 13487 86436 13600
rect 88755 13487 88884 13600
rect 91251 13487 91468 13600
rect 93747 13487 93916 13600
rect 96243 13487 96364 13600
rect 98739 13487 98948 13600
rect 101235 13487 101396 13600
rect 103731 13487 103829 13600
rect 106227 13487 106428 13600
rect 123216 13600 136620 13676
rect 121695 13525 122353 13585
rect 58888 13464 58964 13487
rect 63920 13464 63996 13487
rect 66368 13464 66444 13487
rect 71400 13464 71476 13487
rect 73848 13464 73924 13487
rect 76432 13464 76508 13487
rect 78880 13464 78956 13487
rect 81328 13464 81404 13487
rect 83912 13464 83988 13487
rect 86360 13464 86436 13487
rect 88808 13464 88884 13487
rect 91392 13464 91468 13487
rect 93840 13464 93916 13487
rect 96288 13464 96364 13487
rect 98872 13464 98948 13487
rect 101320 13464 101396 13487
rect 106352 13464 106428 13487
rect 123216 13464 123428 13600
rect 3128 13268 3340 13404
rect 3944 13268 4156 13404
rect 3128 13192 4156 13268
rect 14552 13192 14764 13404
rect 28560 13132 28772 13404
rect 28968 13263 29180 13268
rect 28851 13192 29180 13263
rect 28851 13165 29044 13192
rect 20128 13056 21564 13132
rect 28288 13056 28772 13132
rect 28968 13132 29044 13165
rect 31008 13132 31220 13404
rect 33456 13328 33804 13404
rect 28968 13056 29142 13132
rect 30736 13056 31220 13132
rect 31280 13192 31628 13268
rect 31280 13056 31492 13192
rect 33456 13184 33687 13328
rect 34000 13263 34212 13268
rect 33843 13192 34212 13263
rect 33456 13056 33668 13184
rect 33843 13165 34076 13192
rect 33864 13056 34076 13165
rect 36040 13056 36252 13404
rect 36448 13263 36660 13268
rect 36339 13192 36660 13263
rect 36339 13165 36524 13192
rect 36448 13132 36524 13165
rect 36448 13056 36622 13132
rect 38488 13056 38700 13404
rect 41072 13328 41284 13404
rect 38896 13263 39108 13268
rect 38835 13192 39108 13263
rect 38835 13165 38972 13192
rect 38896 13132 38972 13165
rect 41072 13184 41175 13328
rect 41344 13263 41556 13268
rect 38896 13056 39070 13132
rect 41072 13056 41148 13184
rect 41331 13165 41556 13263
rect 41344 13056 41556 13165
rect 43520 13056 43732 13404
rect 43928 13263 44140 13268
rect 43827 13192 44140 13263
rect 43827 13165 44004 13192
rect 43928 13132 44004 13165
rect 43928 13056 44102 13132
rect 45968 13056 46180 13404
rect 48552 13328 48764 13404
rect 46376 13263 46588 13268
rect 46323 13192 46588 13263
rect 46323 13165 46452 13192
rect 46376 13132 46452 13165
rect 48552 13184 48663 13328
rect 48960 13263 49172 13268
rect 48819 13192 49172 13263
rect 48552 13132 48628 13184
rect 48819 13165 49036 13192
rect 46376 13056 46550 13132
rect 48280 13056 48628 13132
rect 48824 13056 49036 13165
rect 51000 13056 51212 13404
rect 51408 13263 51620 13268
rect 51315 13192 51620 13263
rect 51315 13165 51484 13192
rect 51408 13132 51484 13165
rect 51408 13056 51582 13132
rect 53448 13056 53660 13404
rect 53856 13263 54068 13268
rect 53811 13192 54068 13263
rect 53811 13165 53932 13192
rect 53856 13132 53932 13165
rect 53856 13056 54030 13132
rect 56032 13056 56244 13404
rect 56304 13192 56652 13268
rect 56304 13056 56516 13192
rect 58480 13056 58692 13404
rect 60928 13328 61276 13404
rect 58888 13263 59100 13268
rect 58803 13192 59100 13263
rect 58803 13165 58964 13192
rect 58888 13132 58964 13165
rect 60928 13184 61143 13328
rect 58888 13056 59062 13132
rect 60928 13056 61140 13184
rect 61299 13132 61397 13263
rect 61299 13094 61548 13132
rect 61336 13056 61548 13094
rect 63512 13056 63724 13404
rect 63920 13263 64132 13268
rect 63795 13192 64132 13263
rect 63795 13165 63996 13192
rect 63920 13132 63996 13165
rect 63920 13056 64094 13132
rect 65960 13056 66172 13404
rect 68408 13328 68756 13404
rect 66368 13263 66580 13268
rect 66291 13192 66580 13263
rect 66291 13165 66444 13192
rect 66368 13132 66444 13165
rect 68408 13184 68631 13328
rect 68408 13132 68620 13184
rect 66368 13056 66542 13132
rect 68272 13056 68620 13132
rect 68787 13132 68885 13263
rect 68787 13094 69028 13132
rect 68816 13056 69028 13094
rect 70992 13056 71204 13404
rect 71400 13263 71612 13268
rect 71283 13192 71612 13263
rect 71283 13165 71476 13192
rect 71400 13132 71476 13165
rect 71400 13056 71574 13132
rect 73440 13056 73652 13404
rect 75888 13328 76236 13404
rect 73848 13263 74060 13268
rect 73779 13192 74060 13263
rect 73779 13165 73924 13192
rect 73848 13132 73924 13165
rect 75888 13184 76119 13328
rect 76432 13263 76644 13268
rect 76275 13192 76644 13263
rect 73848 13056 74022 13132
rect 75888 13056 76100 13184
rect 76275 13165 76508 13192
rect 76296 13056 76508 13165
rect 78472 13056 78684 13404
rect 78880 13263 79092 13268
rect 78771 13192 79092 13263
rect 78771 13165 78956 13192
rect 78880 13132 78956 13165
rect 78880 13056 79054 13132
rect 80920 13056 81132 13404
rect 83504 13328 83716 13404
rect 81328 13263 81540 13268
rect 81267 13192 81540 13263
rect 81267 13165 81404 13192
rect 81328 13132 81404 13165
rect 83504 13184 83607 13328
rect 83912 13263 84124 13268
rect 83763 13192 84124 13263
rect 81328 13056 81502 13132
rect 83504 13056 83580 13184
rect 83763 13165 83988 13192
rect 83776 13056 83988 13165
rect 85952 13056 86164 13404
rect 86360 13263 86572 13268
rect 86259 13192 86572 13263
rect 86259 13165 86436 13192
rect 86360 13132 86436 13165
rect 86360 13056 86534 13132
rect 88400 13056 88612 13404
rect 90984 13328 91196 13404
rect 88808 13263 89020 13268
rect 88755 13192 89020 13263
rect 88755 13165 88884 13192
rect 88808 13132 88884 13165
rect 90984 13184 91095 13328
rect 91392 13263 91604 13268
rect 91251 13192 91604 13263
rect 88808 13056 88982 13132
rect 90984 13056 91060 13184
rect 91251 13165 91468 13192
rect 91256 13056 91468 13165
rect 93432 13056 93644 13404
rect 93840 13263 94052 13268
rect 93747 13192 94052 13263
rect 93747 13165 93916 13192
rect 93840 13132 93916 13165
rect 93840 13056 94014 13132
rect 95880 13056 96092 13404
rect 96288 13263 96500 13268
rect 96243 13192 96500 13263
rect 96243 13165 96364 13192
rect 96288 13132 96364 13165
rect 96288 13056 96462 13132
rect 98464 13056 98676 13404
rect 98872 13263 99084 13268
rect 98739 13192 99084 13263
rect 98739 13165 98948 13192
rect 98872 13132 98948 13165
rect 98872 13056 99046 13132
rect 100912 13056 101124 13404
rect 103360 13328 103708 13404
rect 101320 13263 101532 13268
rect 101235 13192 101532 13263
rect 101235 13165 101396 13192
rect 101320 13132 101396 13165
rect 103360 13184 103575 13328
rect 101320 13056 101494 13132
rect 103360 13056 103572 13184
rect 103731 13132 103829 13263
rect 103731 13094 103980 13132
rect 103768 13056 103980 13094
rect 105944 13056 106156 13404
rect 106352 13263 106564 13268
rect 106227 13192 106564 13263
rect 106227 13165 106428 13192
rect 106352 13132 106428 13165
rect 106352 13056 106526 13132
rect 20128 12920 20340 13056
rect 21216 12920 21564 13056
rect 122808 12648 123020 12860
rect 14694 12539 26663 12599
rect 28696 12512 29180 12588
rect 31144 12512 31492 12588
rect 1224 12240 1980 12316
rect 28696 12240 28908 12512
rect 31144 12316 31356 12512
rect 33728 12316 33940 12588
rect 31144 12240 31492 12316
rect 33456 12240 33940 12316
rect 36176 12512 36660 12588
rect 38624 12512 39108 12588
rect 41208 12512 41556 12588
rect 43656 12512 44140 12588
rect 46104 12512 46588 12588
rect 36176 12240 36388 12512
rect 38624 12240 38836 12512
rect 41208 12316 41420 12512
rect 43656 12316 43868 12512
rect 41208 12240 41556 12316
rect 43422 12240 43868 12316
rect 46104 12316 46316 12512
rect 46104 12240 46588 12316
rect 48688 12240 48900 12588
rect 51136 12512 51620 12588
rect 53584 12512 54068 12588
rect 56168 12512 56516 12588
rect 58616 12512 59100 12588
rect 51136 12240 51348 12512
rect 53584 12316 53796 12512
rect 56168 12316 56380 12512
rect 58616 12316 58828 12512
rect 53584 12240 54068 12316
rect 56168 12240 56516 12316
rect 58616 12240 59100 12316
rect 61064 12240 61412 12588
rect 63648 12512 64132 12588
rect 66096 12512 66580 12588
rect 63648 12240 63860 12512
rect 66096 12240 66308 12512
rect 68544 12240 68892 12588
rect 71128 12512 71612 12588
rect 73576 12512 74060 12588
rect 71128 12316 71340 12512
rect 73576 12316 73788 12512
rect 71128 12240 71612 12316
rect 73342 12240 73788 12316
rect 76160 12240 76372 12588
rect 78608 12512 79092 12588
rect 81056 12512 81540 12588
rect 78608 12240 78820 12512
rect 81056 12240 81268 12512
rect 83640 12316 83852 12588
rect 86088 12512 86572 12588
rect 88536 12512 89020 12588
rect 86088 12316 86300 12512
rect 88536 12316 88748 12512
rect 83640 12240 84124 12316
rect 86088 12240 86572 12316
rect 88536 12240 89020 12316
rect 91120 12240 91332 12588
rect 93568 12512 94052 12588
rect 96016 12512 96500 12588
rect 98600 12512 99084 12588
rect 101048 12512 101532 12588
rect 93568 12240 93780 12512
rect 96016 12240 96228 12512
rect 98600 12316 98812 12512
rect 101048 12316 101260 12512
rect 98600 12240 99084 12316
rect 101048 12240 101532 12316
rect 103496 12240 103844 12588
rect 106080 12512 106564 12588
rect 106080 12240 106292 12512
rect 134776 12240 135396 12316
rect 1768 11968 1980 12240
rect 14552 11696 14764 12044
rect 28696 11968 29044 12044
rect 28696 11832 28908 11968
rect 31144 11832 31356 12044
rect 33592 11968 34076 12044
rect 36176 11968 36524 12044
rect 38624 11968 38972 12044
rect 41072 11968 44004 12044
rect 46104 11968 46452 12044
rect 48688 11968 49036 12044
rect 51136 11968 51484 12044
rect 53584 11968 53932 12044
rect 33592 11832 33940 11968
rect 36176 11908 36388 11968
rect 38624 11908 38836 11968
rect 36176 11832 38836 11908
rect 41072 11832 41420 11968
rect 43656 11832 43868 11968
rect 46104 11832 46316 11968
rect 48688 11832 48900 11968
rect 51136 11832 51348 11968
rect 53584 11908 53796 11968
rect 53584 11832 53932 11908
rect 56168 11832 56380 12044
rect 58616 11968 58964 12044
rect 58616 11832 58828 11968
rect 61064 11832 61276 12044
rect 63648 11968 63996 12044
rect 66096 11968 66444 12044
rect 63648 11908 63860 11968
rect 66096 11908 66308 11968
rect 63648 11832 66308 11908
rect 68544 11832 68892 12044
rect 71128 11968 71476 12044
rect 73576 11968 73924 12044
rect 76024 11968 76508 12044
rect 78608 11968 78956 12044
rect 81056 11968 81404 12044
rect 83504 11968 83988 12044
rect 86088 11968 86436 12044
rect 88536 11968 88884 12044
rect 91120 11968 91468 12044
rect 93568 11968 93916 12044
rect 96016 11968 96364 12044
rect 98600 11968 98948 12044
rect 101048 11968 101396 12044
rect 71128 11832 71340 11968
rect 73576 11832 73788 11968
rect 76024 11832 76372 11968
rect 78608 11908 78820 11968
rect 81056 11908 81268 11968
rect 83504 11908 83852 11968
rect 78608 11832 83852 11908
rect 86088 11832 86300 11968
rect 88536 11908 88748 11968
rect 88536 11832 88884 11908
rect 91120 11832 91332 11968
rect 93568 11832 93780 11968
rect 96016 11832 96228 11968
rect 98600 11832 98812 11968
rect 101048 11832 101260 11968
rect 103496 11832 103708 12044
rect 106080 11968 106428 12044
rect 106080 11832 106292 11968
rect 121615 11967 122353 12027
rect 123216 11832 123428 12044
rect 134776 11968 134988 12240
rect 20128 11696 21564 11772
rect 20128 11560 20340 11696
rect 21216 11560 21564 11696
rect 28832 11560 29044 11772
rect 31280 11560 31492 11772
rect 33494 11696 33940 11772
rect 36214 11696 36524 11772
rect 38662 11696 38972 11772
rect 33728 11560 33940 11696
rect 28832 11500 28908 11560
rect 31280 11500 31356 11560
rect 33864 11500 33940 11560
rect 36312 11560 36524 11696
rect 38760 11560 38972 11696
rect 41208 11560 41556 11772
rect 43792 11560 44004 11772
rect 46240 11696 46550 11772
rect 46240 11560 46452 11696
rect 48688 11560 49036 11772
rect 51272 11560 51484 11772
rect 53720 11696 54030 11772
rect 53720 11560 53932 11696
rect 56168 11560 56516 11772
rect 58752 11696 59062 11772
rect 58752 11560 58964 11696
rect 61200 11560 61412 11772
rect 63686 11696 63996 11772
rect 63784 11560 63996 11696
rect 66232 11560 66444 11772
rect 68582 11696 68892 11772
rect 68680 11560 68892 11696
rect 71264 11696 71574 11772
rect 71264 11560 71476 11696
rect 73712 11560 73924 11772
rect 76160 11560 76372 11772
rect 78646 11696 78956 11772
rect 81094 11696 81404 11772
rect 78744 11560 78956 11696
rect 81192 11560 81404 11696
rect 83640 11696 84086 11772
rect 86224 11696 86534 11772
rect 88672 11696 88982 11772
rect 83640 11560 83988 11696
rect 86224 11560 86436 11696
rect 88672 11560 88884 11696
rect 91120 11560 91468 11772
rect 93704 11560 93916 11772
rect 96054 11696 96364 11772
rect 96152 11560 96364 11696
rect 98600 11696 99046 11772
rect 101184 11696 101494 11772
rect 98600 11560 98948 11696
rect 101184 11560 101396 11696
rect 103632 11560 103844 11772
rect 106118 11696 106428 11772
rect 106216 11560 106428 11696
rect 36312 11500 36388 11560
rect 38760 11500 38836 11560
rect 28696 11364 28908 11500
rect 28190 11288 28908 11364
rect 31144 11288 31356 11500
rect 33592 11288 33940 11500
rect 36176 11288 36388 11500
rect 38624 11288 38836 11500
rect 41208 11500 41284 11560
rect 43792 11500 43868 11560
rect 46240 11500 46316 11560
rect 48824 11500 48900 11560
rect 51272 11500 51348 11560
rect 53720 11500 53796 11560
rect 41208 11288 41420 11500
rect 43384 11424 43868 11500
rect 43656 11288 43868 11424
rect 46104 11288 46316 11500
rect 48688 11288 48900 11500
rect 51136 11288 51348 11500
rect 53584 11288 53796 11500
rect 56168 11500 56244 11560
rect 58752 11500 58828 11560
rect 61200 11500 61276 11560
rect 63784 11500 63860 11560
rect 66232 11500 66308 11560
rect 68680 11500 68756 11560
rect 71264 11500 71340 11560
rect 73712 11500 73788 11560
rect 76160 11500 76236 11560
rect 78744 11500 78820 11560
rect 81192 11500 81268 11560
rect 56168 11288 56380 11500
rect 58616 11288 58828 11500
rect 61064 11288 61412 11500
rect 63648 11288 63860 11500
rect 66096 11288 66308 11500
rect 68544 11288 68892 11500
rect 71128 11288 71340 11500
rect 73304 11424 73788 11500
rect 73576 11288 73788 11424
rect 76024 11288 76372 11500
rect 78608 11288 78820 11500
rect 81056 11288 81268 11500
rect 83640 11500 83716 11560
rect 86224 11500 86300 11560
rect 88672 11500 88748 11560
rect 91256 11500 91332 11560
rect 93704 11500 93780 11560
rect 96152 11500 96228 11560
rect 83640 11288 83852 11500
rect 86088 11288 86300 11500
rect 88536 11288 88748 11500
rect 91120 11288 91332 11500
rect 93568 11288 93780 11500
rect 96016 11288 96228 11500
rect 98600 11500 98676 11560
rect 101184 11500 101260 11560
rect 103632 11500 103708 11560
rect 106216 11500 106292 11560
rect 98600 11288 98812 11500
rect 101048 11288 101260 11500
rect 103496 11288 103844 11500
rect 106080 11364 106292 11500
rect 106080 11288 108468 11364
rect 122808 11288 123020 11500
rect 28598 11016 31356 11092
rect 33728 11016 36388 11092
rect 38624 11016 38836 11092
rect 41208 11016 41420 11092
rect 43656 11016 46452 11092
rect 48688 11016 53932 11092
rect 56168 11016 56380 11092
rect 58616 11016 58828 11092
rect 61064 11016 61412 11092
rect 63648 11016 63860 11092
rect 66096 11016 73788 11092
rect 76160 11016 78820 11092
rect 81056 11016 81268 11092
rect 83640 11016 83852 11092
rect 86088 11016 96364 11092
rect 98600 11016 98812 11092
rect 101048 11016 101260 11092
rect 103496 11016 103844 11092
rect 106080 11016 108332 11092
rect 28746 10985 28844 11016
rect 31242 10985 31340 11016
rect 33738 10985 33836 11016
rect 36234 10985 36332 11016
rect 38730 10985 38828 11016
rect 41226 10985 41324 11016
rect 43722 10985 43820 11016
rect 46218 10985 46316 11016
rect 48714 10985 48812 11016
rect 51210 10985 51308 11016
rect 53706 10985 53804 11016
rect 56202 10985 56300 11016
rect 58698 10985 58796 11016
rect 61194 10985 61292 11016
rect 63690 10985 63788 11016
rect 66186 10985 66284 11016
rect 68682 10985 68780 11016
rect 71178 10985 71276 11016
rect 73674 10985 73772 11016
rect 76170 10985 76268 11016
rect 78666 10985 78764 11016
rect 81162 10985 81260 11016
rect 83658 10985 83756 11016
rect 86154 10985 86252 11016
rect 88650 10985 88748 11016
rect 91146 10985 91244 11016
rect 93642 10985 93740 11016
rect 96138 10985 96236 11016
rect 98634 10985 98732 11016
rect 101130 10985 101228 11016
rect 103626 10985 103724 11016
rect 106122 10985 106220 11016
rect 121535 10697 122353 10757
rect 123216 10744 123428 10956
rect 27064 10608 28636 10684
rect 1224 10472 1980 10548
rect 1768 10336 1980 10472
rect 2448 10412 2796 10548
rect 2040 10336 2796 10412
rect 14552 10336 14764 10548
rect 27064 10472 27276 10608
rect 108256 10472 108468 10684
rect 134776 10412 134988 10548
rect 134776 10336 135396 10412
rect 2040 10276 2116 10336
rect 544 10200 2116 10276
rect 0 9928 2932 10004
rect 2720 9792 2932 9928
rect 122808 9792 123020 10004
rect 27064 9520 28228 9596
rect 27064 9384 27276 9520
rect 108256 9384 108468 9596
rect 2448 8976 2796 9188
rect 14552 9052 14764 9188
rect 14552 8976 16396 9052
rect 2448 8916 2524 8976
rect 1768 8840 2524 8916
rect 1768 8780 1980 8840
rect 1224 8704 1980 8780
rect 134776 8780 134988 8916
rect 134776 8704 135396 8780
rect 0 8296 6060 8372
rect 2720 8100 2932 8236
rect 5848 8160 6060 8296
rect 0 8024 2932 8100
rect 544 7616 2796 7692
rect 2448 7480 2796 7616
rect 14552 7480 14764 7692
rect 1224 7208 1980 7284
rect 1768 6936 1980 7208
rect 134776 7148 134988 7284
rect 134776 7072 135396 7148
rect 134776 6936 134988 7072
rect 1224 5440 1980 5516
rect 1768 5304 1980 5440
rect 134776 5380 134988 5516
rect 134776 5304 135396 5380
rect 1224 3808 1980 3884
rect 1768 3672 1980 3808
rect 16320 3808 17756 3884
rect 16320 3672 16532 3808
rect 17544 3748 17756 3808
rect 18632 3748 18844 3884
rect 19856 3808 21292 3884
rect 19856 3748 20068 3808
rect 20944 3748 21292 3808
rect 22168 3748 22380 3884
rect 23392 3808 25916 3884
rect 23392 3748 23604 3808
rect 17544 3672 20340 3748
rect 20944 3672 23604 3748
rect 24480 3672 24692 3808
rect 25704 3748 25916 3808
rect 26792 3748 27140 3884
rect 28016 3808 29452 3884
rect 28016 3748 28228 3808
rect 25704 3672 28228 3748
rect 29240 3748 29452 3808
rect 30328 3748 30540 3884
rect 31552 3808 34076 3884
rect 31552 3748 31764 3808
rect 29240 3672 31764 3748
rect 32640 3672 32852 3808
rect 33864 3748 34076 3808
rect 34952 3808 37612 3884
rect 34952 3748 35300 3808
rect 33864 3672 35300 3748
rect 36176 3672 36388 3808
rect 37400 3748 37612 3808
rect 38488 3748 38700 3884
rect 39712 3808 41148 3884
rect 39712 3748 39924 3808
rect 37400 3672 39924 3748
rect 40800 3748 41148 3808
rect 42024 3748 42236 3884
rect 43248 3808 45772 3884
rect 43248 3748 43460 3808
rect 40800 3672 43460 3748
rect 44336 3672 44548 3808
rect 45560 3748 45772 3808
rect 46648 3748 46996 3884
rect 47872 3808 49308 3884
rect 47872 3748 48084 3808
rect 45560 3672 48084 3748
rect 49096 3748 49308 3808
rect 50184 3748 50396 3884
rect 51408 3808 53932 3884
rect 51408 3748 51620 3808
rect 49096 3672 51620 3748
rect 52496 3672 52708 3808
rect 53720 3748 53932 3808
rect 54808 3748 55156 3884
rect 56032 3808 57468 3884
rect 56032 3748 56244 3808
rect 53720 3672 56244 3748
rect 57256 3748 57468 3808
rect 58344 3748 58556 3884
rect 59568 3748 59780 3884
rect 57256 3672 59780 3748
rect 134776 3748 134988 3884
rect 134776 3672 135396 3748
rect 15912 2856 16124 3068
rect 17136 2856 17348 3068
rect 18224 2856 18436 3068
rect 19584 3009 19660 3068
rect 20672 3009 20884 3068
rect 21896 3009 21972 3068
rect 19487 2932 19660 3009
rect 20655 2932 20884 3009
rect 21823 2932 21972 3009
rect 19448 2856 19660 2932
rect 20536 2856 20884 2932
rect 21760 2856 21972 2932
rect 22984 2856 23196 3068
rect 24208 3009 24284 3068
rect 24159 2932 24284 3009
rect 24072 2856 24284 2932
rect 25296 2856 25508 3068
rect 26520 3009 26596 3068
rect 27744 3009 27820 3068
rect 28832 3009 29044 3068
rect 30056 3009 30132 3068
rect 26495 2932 26596 3009
rect 27663 2932 27820 3009
rect 28831 2932 29044 3009
rect 29999 2932 30132 3009
rect 26384 2856 26596 2932
rect 27608 2856 27820 2932
rect 28696 2856 29044 2932
rect 29920 2856 30132 2932
rect 31144 2856 31356 3068
rect 32368 3009 32444 3068
rect 33592 3009 33668 3068
rect 34680 3009 34892 3068
rect 35904 3009 35980 3068
rect 32335 2932 32444 3009
rect 33503 2932 33668 3009
rect 34671 2932 34892 3009
rect 35839 2932 35980 3009
rect 32232 2856 32444 2932
rect 33456 2856 33668 2932
rect 34544 2856 34892 2932
rect 35768 2856 35980 2932
rect 36992 2856 37204 3068
rect 38216 3009 38292 3068
rect 39440 3009 39516 3068
rect 40528 3009 40740 3068
rect 41752 3009 41828 3068
rect 38175 2932 38292 3009
rect 39343 2932 39516 3009
rect 40511 2932 40740 3009
rect 41679 2932 41828 3009
rect 38080 2856 38292 2932
rect 39304 2856 39516 2932
rect 40392 2856 40740 2932
rect 41616 2856 41828 2932
rect 42840 2856 43052 3068
rect 44064 3009 44140 3068
rect 44015 2932 44140 3009
rect 43928 2856 44140 2932
rect 45152 2856 45364 3068
rect 46376 3009 46452 3068
rect 47600 3009 47676 3068
rect 48688 3009 48900 3068
rect 49912 3009 49988 3068
rect 46351 2932 46452 3009
rect 47519 2932 47676 3009
rect 48687 2932 48900 3009
rect 49855 2932 49988 3009
rect 46240 2856 46452 2932
rect 47464 2856 47676 2932
rect 48552 2856 48900 2932
rect 49776 2856 49988 2932
rect 51000 2856 51212 3068
rect 52224 3009 52300 3068
rect 53448 3009 53524 3068
rect 54536 3009 54748 3068
rect 55760 3009 55836 3068
rect 52191 2932 52300 3009
rect 53359 2932 53524 3009
rect 54527 2932 54748 3009
rect 55695 2932 55836 3009
rect 52088 2856 52300 2932
rect 53312 2856 53524 2932
rect 54400 2856 54748 2932
rect 55624 2856 55836 2932
rect 56848 2856 57060 3068
rect 58072 3009 58148 3068
rect 59296 3009 59372 3068
rect 58031 2932 58148 3009
rect 59199 2932 59372 3009
rect 57936 2856 58148 2932
rect 59160 2856 59372 2932
rect 14778 2674 17030 2734
rect 16320 2448 17756 2524
rect 16320 2312 16532 2448
rect 17544 2388 17756 2448
rect 18632 2388 18844 2524
rect 19856 2448 22380 2524
rect 19856 2388 20068 2448
rect 17544 2312 20068 2388
rect 20944 2312 21292 2448
rect 22168 2388 22380 2448
rect 23392 2448 25916 2524
rect 23392 2388 23604 2448
rect 22168 2312 23604 2388
rect 24480 2312 24692 2448
rect 25704 2388 25916 2448
rect 26792 2388 27140 2524
rect 28016 2448 29452 2524
rect 28016 2388 28228 2448
rect 25704 2312 28228 2388
rect 29240 2388 29452 2448
rect 30328 2388 30540 2524
rect 31552 2448 34076 2524
rect 31552 2388 31764 2448
rect 29240 2312 31764 2388
rect 32640 2312 32852 2448
rect 33864 2388 34076 2448
rect 34952 2388 35300 2524
rect 36176 2448 37612 2524
rect 36176 2388 36388 2448
rect 33864 2312 36388 2388
rect 37400 2388 37612 2448
rect 38488 2388 38700 2524
rect 39712 2448 42236 2524
rect 39712 2388 39924 2448
rect 37400 2312 39924 2388
rect 40800 2312 41148 2448
rect 42024 2388 42236 2448
rect 43248 2448 45772 2524
rect 43248 2388 43460 2448
rect 42024 2312 43460 2388
rect 44336 2312 44548 2448
rect 45560 2388 45772 2448
rect 46648 2388 46996 2524
rect 47872 2448 49308 2524
rect 47872 2388 48084 2448
rect 45560 2312 48084 2388
rect 49096 2388 49308 2448
rect 50184 2388 50396 2524
rect 51408 2448 53932 2524
rect 51408 2388 51620 2448
rect 49096 2312 51620 2388
rect 52496 2312 52708 2448
rect 53720 2388 53932 2448
rect 54808 2448 57468 2524
rect 54808 2388 55156 2448
rect 53720 2312 55156 2388
rect 56032 2312 56244 2448
rect 57256 2388 57468 2448
rect 58344 2388 58556 2524
rect 59568 2388 59780 2524
rect 57256 2312 59780 2388
rect 1768 1980 1980 2116
rect 134776 2040 135396 2116
rect 1768 1904 2116 1980
rect 134776 1904 134988 2040
rect 2040 1844 2116 1904
rect 2040 1632 2252 1844
rect 3672 1632 4020 1844
rect 5440 1632 5652 1844
rect 7072 1632 7284 1844
rect 8704 1632 9052 1844
rect 10472 1632 10684 1844
rect 12104 1632 12316 1844
rect 13736 1632 14084 1844
rect 15504 1632 15716 1844
rect 17136 1708 17348 1844
rect 17136 1632 17484 1708
rect 18904 1632 19116 1844
rect 20302 1768 20748 1844
rect 20536 1708 20748 1768
rect 20536 1632 20884 1708
rect 22168 1632 22380 1844
rect 23936 1632 24148 1844
rect 25568 1632 25780 1844
rect 27200 1632 27412 1844
rect 28968 1632 29180 1844
rect 30600 1708 30812 1844
rect 32232 1708 32580 1844
rect 30464 1632 30812 1708
rect 32096 1632 32580 1708
rect 34000 1632 34212 1844
rect 35632 1632 35844 1844
rect 37264 1632 37612 1844
rect 39032 1632 39244 1844
rect 40664 1632 40876 1844
rect 42296 1632 42644 1844
rect 44064 1632 44276 1844
rect 45696 1632 45908 1844
rect 47464 1708 47676 1844
rect 47328 1632 47676 1708
rect 49096 1632 49308 1844
rect 50728 1632 50940 1844
rect 52496 1632 52708 1844
rect 54128 1632 54340 1844
rect 55760 1708 55972 1844
rect 55488 1632 55972 1708
rect 57528 1632 57740 1844
rect 59160 1708 59372 1844
rect 59160 1632 59508 1708
rect 60792 1632 61140 1844
rect 62560 1632 62772 1844
rect 64192 1632 64404 1844
rect 65824 1632 66172 1844
rect 67592 1632 67804 1844
rect 69224 1632 69436 1844
rect 70856 1632 71204 1844
rect 72624 1632 72836 1844
rect 74256 1632 74468 1844
rect 76024 1632 76236 1844
rect 77656 1632 77868 1844
rect 79288 1632 79500 1844
rect 81056 1632 81268 1844
rect 82688 1632 82900 1844
rect 84320 1632 84532 1844
rect 86088 1632 86300 1844
rect 87720 1632 87932 1844
rect 89352 1632 89700 1844
rect 91120 1632 91332 1844
rect 92752 1632 92964 1844
rect 94384 1632 94732 1844
rect 96152 1632 96364 1844
rect 97784 1632 97996 1844
rect 99416 1632 99764 1844
rect 101184 1632 101396 1844
rect 102816 1632 103028 1844
rect 104584 1632 104796 1844
rect 106216 1632 106428 1844
rect 107848 1632 108060 1844
rect 109616 1632 109828 1844
rect 111248 1632 111460 1844
rect 112880 1632 113092 1844
rect 114648 1632 114860 1844
rect 116280 1632 116492 1844
rect 117912 1632 118260 1844
rect 119680 1632 119892 1844
rect 121312 1632 121524 1844
rect 122944 1632 123292 1844
rect 124712 1632 124924 1844
rect 126344 1632 126556 1844
rect 127976 1632 128324 1844
rect 129744 1632 129956 1844
rect 131376 1632 131588 1844
rect 133144 1632 133356 1844
rect 952 952 135668 1300
rect 272 272 136348 620
<< metal4 >>
rect 272 272 620 83036
rect 952 952 1300 82356
rect 2176 81502 2252 82084
rect 3944 81502 4020 82084
rect 5440 81502 5516 82084
rect 7208 81502 7284 82084
rect 8704 81502 8780 82084
rect 10472 81502 10548 82084
rect 12104 81502 12180 82084
rect 14008 81502 14084 82084
rect 15640 81502 15716 82084
rect 17136 81502 17212 82084
rect 18904 81502 18980 82084
rect 20672 81502 20748 82084
rect 22168 81502 22244 82084
rect 23936 81502 24012 82084
rect 25704 81502 25780 82084
rect 27200 81502 27276 82084
rect 2040 81094 2116 81404
rect 28696 77150 28772 83308
rect 28968 81502 29044 82084
rect 30600 81502 30676 82084
rect 31008 77150 31084 83308
rect 32368 81502 32444 82084
rect 33456 77150 33532 83308
rect 34136 81502 34212 82084
rect 35632 81502 35708 82084
rect 36176 77150 36252 83308
rect 37536 81502 37612 82084
rect 38488 77150 38564 83308
rect 39168 81502 39244 82084
rect 40664 81502 40740 82084
rect 41072 77150 41148 83308
rect 42432 81502 42508 82084
rect 43520 77150 43596 83308
rect 44200 81502 44276 82084
rect 45696 81502 45772 82084
rect 46104 77150 46180 83308
rect 47464 81502 47540 82084
rect 48552 77150 48628 83308
rect 49232 81502 49308 82084
rect 50728 81502 50804 82084
rect 51136 77150 51212 83308
rect 52632 81502 52708 82084
rect 53584 77150 53660 83308
rect 54128 81502 54204 82084
rect 55896 81502 55972 82084
rect 56168 77150 56244 83308
rect 57664 81502 57740 82084
rect 58480 77150 58556 83308
rect 59160 81502 59236 82084
rect 60792 81502 60868 82084
rect 60928 77150 61004 83308
rect 62696 81502 62772 82084
rect 63648 77150 63724 83308
rect 64192 81502 64268 82084
rect 65824 81502 65900 82084
rect 66096 77150 66172 83308
rect 67592 81502 67668 82084
rect 68544 77150 68620 83308
rect 69224 81502 69300 82084
rect 70856 81502 70932 82084
rect 70992 77150 71068 83308
rect 72624 81502 72700 82084
rect 73576 77150 73652 83308
rect 74392 81502 74468 82084
rect 75888 77150 75964 83308
rect 76160 81502 76236 82084
rect 77656 81502 77732 82084
rect 78608 77150 78684 83308
rect 79424 81502 79500 82084
rect 81056 77150 81132 83308
rect 81328 81502 81404 82084
rect 82688 81502 82764 82084
rect 83504 77150 83580 83308
rect 84456 81502 84532 82084
rect 85952 77150 86028 83308
rect 86224 81502 86300 82084
rect 87720 81502 87796 82084
rect 88400 77150 88476 83308
rect 89352 81502 89428 82084
rect 90984 77150 91060 83308
rect 91120 81502 91196 82084
rect 92888 81502 92964 82084
rect 93568 77150 93644 83308
rect 94384 81502 94460 82084
rect 96016 77150 96092 83308
rect 96288 81502 96364 82084
rect 97920 81502 97996 82084
rect 98464 77150 98540 83308
rect 99688 81502 99764 82084
rect 101048 77150 101124 83308
rect 101320 81502 101396 82084
rect 102952 81502 103028 82084
rect 103360 77150 103436 83308
rect 104584 81502 104660 82084
rect 106080 77150 106156 83308
rect 106352 81502 106428 82084
rect 107848 81502 107924 82084
rect 109616 81502 109692 82084
rect 111384 81502 111460 82084
rect 112880 81502 112956 82084
rect 114648 81502 114724 82084
rect 116416 81502 116492 82084
rect 117912 81502 117988 82084
rect 118048 80822 118124 82764
rect 117912 78646 117988 80724
rect 118184 79424 118260 81366
rect 118456 80278 118532 83308
rect 119544 81502 119620 82084
rect 119680 80278 119756 83308
rect 121448 81502 121524 82084
rect 123216 81502 123292 82084
rect 124712 81502 124788 82084
rect 126344 81502 126420 82084
rect 128112 81502 128188 82084
rect 129880 81502 129956 82084
rect 122264 79832 122340 80686
rect 28968 76780 29044 77014
rect 28832 76704 29044 76780
rect 28832 75208 28908 76704
rect 28968 75926 29044 76644
rect 31280 75926 31356 76644
rect 31416 75208 31492 77014
rect 33728 75926 33804 76644
rect 34000 75208 34076 77014
rect 36312 75926 36388 76644
rect 36448 75208 36524 77014
rect 38624 75888 38700 76606
rect 38896 75926 38972 76644
rect 39032 75208 39108 77014
rect 41344 75926 41420 76644
rect 41480 75208 41556 77014
rect 43928 76780 44004 77014
rect 43792 76704 44004 76780
rect 43656 75888 43732 76606
rect 43792 75208 43868 76704
rect 43928 75926 44004 76644
rect 46376 75926 46452 76644
rect 46512 75208 46588 77014
rect 48688 75926 48764 76644
rect 48960 75208 49036 77014
rect 51408 76780 51484 77014
rect 51272 76704 51484 76780
rect 51272 75208 51348 76704
rect 51408 75926 51484 76644
rect 53720 75926 53796 76644
rect 53856 75208 53932 77014
rect 56168 75888 56244 76606
rect 56304 75926 56380 76644
rect 56440 75208 56516 77014
rect 58752 75926 58828 76644
rect 58888 75208 58964 77014
rect 61336 75926 61412 76644
rect 28968 73168 29044 75110
rect 31552 73168 31628 75110
rect 34000 73168 34076 75110
rect 36448 73168 36524 75110
rect 39032 73168 39108 75110
rect 41480 73168 41556 75110
rect 44064 73168 44140 75110
rect 46512 73168 46588 75110
rect 48960 73168 49036 75110
rect 51544 73168 51620 75110
rect 53992 73168 54068 75110
rect 56304 73206 56380 75148
rect 59024 73168 59100 75110
rect 28560 71030 28636 71476
rect 28696 70992 28772 71438
rect 28968 70758 29044 73108
rect 59432 71536 59508 75790
rect 61472 75208 61548 77150
rect 63784 75926 63860 76644
rect 63920 75208 63996 77014
rect 66368 75926 66444 76644
rect 66504 75208 66580 77014
rect 68816 75926 68892 76644
rect 68952 75208 69028 77150
rect 71400 76780 71476 77014
rect 71264 76704 71476 76780
rect 71128 75926 71204 76644
rect 71264 75208 71340 76704
rect 71400 75926 71476 76644
rect 73712 75926 73788 76644
rect 73848 75208 73924 77014
rect 76160 75926 76236 76644
rect 76432 75208 76508 77014
rect 78608 75888 78684 76606
rect 78744 75926 78820 76644
rect 78880 75208 78956 77014
rect 81328 75926 81404 76644
rect 81464 75208 81540 77014
rect 83776 75926 83852 76644
rect 83912 75208 83988 77014
rect 86360 76780 86436 77014
rect 86224 76704 86436 76780
rect 86224 75208 86300 76704
rect 86360 75926 86436 76644
rect 88536 75926 88612 76644
rect 88808 75926 88884 76644
rect 88944 75208 89020 77014
rect 91256 75208 91332 77150
rect 93840 76780 93916 77014
rect 93704 76704 93916 76780
rect 91392 75926 91468 76644
rect 93568 75888 93644 76606
rect 93704 75208 93780 76704
rect 93840 75926 93916 76644
rect 96152 75926 96228 76644
rect 96288 75208 96364 77014
rect 98600 75888 98676 76606
rect 98736 75926 98812 76644
rect 98872 75208 98948 77014
rect 101184 75926 101260 76644
rect 101320 75208 101396 77014
rect 103768 75926 103844 76644
rect 103904 75208 103980 77150
rect 106216 75926 106292 76644
rect 106352 75208 106428 77014
rect 61472 73168 61548 75110
rect 63920 73168 63996 75110
rect 66504 73168 66580 75110
rect 68952 73168 69028 75110
rect 71400 73168 71476 75110
rect 73984 73168 74060 75110
rect 76432 73168 76508 75110
rect 78880 73168 78956 75110
rect 81464 73168 81540 75110
rect 83912 73168 83988 75110
rect 86496 73168 86572 75110
rect 88944 73168 89020 75110
rect 91392 73168 91468 75110
rect 93704 73206 93780 75148
rect 96424 73168 96500 75110
rect 98872 73168 98948 75110
rect 101456 73168 101532 75110
rect 103904 73168 103980 75110
rect 106352 73168 106428 75110
rect 115328 74392 115404 77150
rect 116552 75888 116628 78510
rect 118048 77286 118124 79364
rect 29784 71030 29860 71476
rect 31280 70992 31356 71438
rect 31960 71030 32036 71476
rect 32504 70992 32580 71438
rect 33728 70992 33804 71438
rect 34408 71030 34484 71476
rect 34952 70992 35028 71438
rect 35768 71030 35844 71476
rect 36176 70992 36252 71438
rect 36992 71030 37068 71476
rect 37536 70992 37612 71438
rect 38216 71030 38292 71476
rect 39984 70992 40060 71438
rect 40664 71030 40740 71476
rect 41208 70992 41284 71438
rect 41888 71030 41964 71476
rect 42432 70992 42508 71438
rect 43248 71030 43324 71476
rect 44608 70856 44684 71438
rect 45696 71030 45772 71476
rect 46240 70992 46316 71438
rect 46920 71030 46996 71476
rect 48688 70992 48764 71438
rect 49912 70992 49988 71438
rect 50728 71030 50804 71476
rect 51272 70992 51348 71438
rect 52496 70992 52572 71438
rect 53176 71030 53252 71476
rect 53312 70992 53388 71438
rect 54400 71030 54476 71476
rect 54944 70992 55020 71438
rect 56032 71030 56108 71476
rect 57392 70992 57468 71438
rect 58616 70992 58692 71438
rect 59432 71030 59508 71476
rect 59976 70992 60052 71438
rect 61200 70992 61276 71438
rect 61880 71030 61956 71476
rect 62424 70992 62500 71438
rect 63104 71030 63180 71476
rect 63648 70992 63724 71438
rect 65008 70992 65084 71438
rect 66096 70992 66172 71438
rect 66912 71030 66988 71476
rect 67456 70992 67532 71438
rect 68136 71030 68212 71476
rect 68680 70992 68756 71438
rect 69904 70992 69980 71438
rect 70584 71030 70660 71476
rect 72080 70856 72156 71438
rect 72216 71030 72292 71476
rect 73712 70992 73788 71438
rect 74392 71030 74468 71476
rect 74936 70992 75012 71438
rect 75616 71030 75692 71476
rect 76160 70992 76236 71438
rect 76840 71030 76916 71476
rect 77384 70992 77460 71438
rect 78200 71030 78276 71476
rect 78472 71030 78548 71476
rect 79424 71030 79500 71476
rect 79968 70992 80044 71438
rect 80648 71030 80724 71476
rect 81872 71030 81948 71476
rect 82416 70992 82492 71438
rect 83096 71030 83172 71476
rect 83640 70992 83716 71438
rect 84592 70992 84668 71438
rect 86088 70992 86164 71438
rect 86904 71030 86980 71476
rect 88128 71030 88204 71476
rect 88672 70992 88748 71438
rect 89352 71030 89428 71476
rect 89896 70992 89972 71438
rect 90712 71030 90788 71476
rect 91120 70992 91196 71438
rect 92344 70992 92420 71438
rect 93296 70856 93372 71438
rect 94928 70992 95004 71438
rect 95608 71030 95684 71476
rect 96832 71030 96908 71476
rect 97376 70992 97452 71438
rect 98600 70992 98676 71302
rect 99824 70992 99900 71438
rect 100912 71030 100988 71476
rect 101864 71030 101940 71476
rect 102408 70992 102484 71438
rect 103088 71030 103164 71476
rect 103632 70992 103708 71438
rect 104312 71030 104388 71476
rect 104856 70992 104932 71438
rect 105536 71030 105612 71476
rect 106080 70992 106156 71438
rect 107304 70992 107380 71438
rect 108528 70992 108604 71438
rect 109616 70856 109692 73070
rect 110704 70584 110780 71030
rect 115328 70622 115404 74332
rect 115464 73032 115540 75654
rect 122264 75616 122340 78374
rect 122400 76976 122476 79734
rect 122944 78510 123020 81404
rect 130832 79190 130908 83308
rect 131376 81502 131452 82084
rect 133144 81502 133220 82084
rect 134776 77656 134852 78374
rect 114240 70040 114316 70486
rect 115872 70040 115948 72934
rect 122264 72798 122340 75556
rect 122400 74294 122476 76916
rect 122400 71400 122476 74022
rect 22168 69670 22244 69980
rect 22440 69670 22516 69980
rect 114376 69632 114452 69942
rect 114648 69670 114724 69980
rect 115328 69632 115404 69942
rect 115464 69670 115540 69980
rect 20808 69224 20884 69534
rect 21352 69224 21428 69534
rect 21624 69262 21700 69572
rect 22168 69262 22244 69572
rect 22440 69224 22516 69534
rect 114240 69262 114316 69572
rect 114648 69224 114724 69534
rect 115056 69262 115132 69572
rect 115600 69262 115676 69572
rect 116008 69262 116084 69572
rect 21760 68854 21836 69164
rect 20808 68544 20884 68854
rect 22032 68816 22108 69126
rect 22440 68816 22516 69126
rect 114376 68816 114452 69126
rect 114784 68816 114860 69126
rect 115192 68854 115268 69164
rect 22032 68408 22108 68718
rect 22440 68446 22516 68756
rect 114376 68408 114452 68718
rect 114648 68446 114724 68756
rect 116008 68582 116084 68892
rect 21896 68038 21972 68348
rect 20808 67728 20884 68038
rect 27472 67902 27548 68212
rect 20808 67358 20884 67668
rect 21216 67358 21292 67668
rect 21624 67358 21700 67668
rect 27336 67592 27412 67902
rect 109480 67864 109556 68174
rect 115328 68038 115404 68348
rect 109344 67358 109420 67804
rect 115872 67728 115948 68038
rect 20808 66950 20884 67260
rect 21488 66912 21564 67222
rect 22032 66950 22108 67260
rect 22440 66950 22516 67260
rect 109480 67086 109556 67396
rect 115600 67358 115676 67668
rect 116008 67358 116084 67668
rect 114376 66950 114452 67260
rect 114648 66912 114724 67222
rect 115872 66950 115948 67260
rect 133144 67086 133220 69844
rect 20808 66504 20884 66814
rect 21624 66504 21700 66814
rect 22032 66542 22108 66852
rect 22440 66504 22516 66814
rect 114376 66542 114452 66852
rect 114784 66542 114860 66852
rect 115600 66542 115676 66852
rect 115872 66504 115948 66814
rect 20944 66134 21020 66444
rect 21352 66096 21428 66406
rect 21488 66096 21564 66406
rect 22168 66096 22244 66406
rect 22576 66134 22652 66444
rect 114240 66096 114316 66406
rect 114648 66096 114724 66406
rect 115056 66096 115132 66406
rect 115328 66096 115404 66406
rect 116008 66096 116084 66406
rect 20808 65726 20884 66036
rect 21760 65688 21836 65998
rect 22032 65726 22108 66036
rect 22576 65688 22652 65998
rect 114376 65726 114452 66036
rect 114648 65688 114724 65998
rect 115600 65688 115676 65998
rect 116008 65688 116084 65998
rect 20944 65280 21020 65590
rect 21352 65318 21428 65628
rect 21488 65318 21564 65628
rect 22032 65280 22108 65590
rect 22440 65318 22516 65628
rect 114376 65280 114452 65590
rect 114648 65318 114724 65628
rect 115192 65280 115268 65590
rect 115328 65280 115404 65590
rect 115872 65280 115948 65590
rect 21896 64872 21972 65182
rect 22032 64464 22108 65046
rect 22168 64910 22244 65220
rect 22440 64872 22516 65182
rect 22168 64464 22244 64774
rect 22576 64502 22652 64812
rect 27608 64736 27684 65046
rect 114240 64872 114316 65182
rect 114648 64872 114724 65182
rect 115056 64910 115132 65220
rect 115464 64872 115540 65182
rect 21760 64094 21836 64404
rect 27336 64230 27412 64540
rect 109344 64328 109420 64774
rect 114376 64502 114452 64812
rect 114648 64464 114724 64774
rect 132600 64366 132676 66988
rect 20808 63784 20884 64094
rect 27608 63920 27684 64230
rect 20808 63376 20884 63686
rect 21896 63376 21972 63686
rect 27472 63550 27548 63860
rect 109208 63550 109284 63996
rect 109480 63920 109556 64230
rect 115328 64056 115404 64366
rect 109344 63550 109420 63860
rect 116008 63784 116084 64094
rect 115464 63414 115540 63724
rect 115872 63414 115948 63724
rect 20808 63006 20884 63316
rect 22032 62968 22108 63278
rect 22576 62968 22652 63278
rect 114240 63006 114316 63316
rect 114784 62968 114860 63278
rect 116008 63006 116084 63316
rect 20808 62560 20884 62870
rect 21760 62560 21836 62870
rect 22032 62598 22108 62908
rect 22440 62598 22516 62908
rect 20808 62152 20884 62462
rect 21216 62152 21292 62462
rect 21624 62190 21700 62500
rect 22032 62152 22108 62462
rect 22576 62190 22652 62500
rect 109344 62288 109420 62598
rect 114240 62560 114316 62870
rect 114648 62560 114724 62870
rect 115056 62560 115132 62870
rect 115464 62598 115540 62908
rect 115872 62598 115948 62908
rect 114376 62190 114452 62500
rect 114784 62190 114860 62500
rect 115192 62190 115268 62500
rect 115872 62152 115948 62462
rect 20944 61782 21020 62092
rect 21352 61782 21428 62092
rect 22168 61744 22244 62054
rect 22440 61744 22516 62054
rect 114240 61744 114316 62054
rect 114648 61782 114724 62092
rect 115464 61744 115540 62054
rect 116008 61744 116084 62054
rect 20944 61336 21020 61646
rect 21760 61336 21836 61646
rect 22032 61374 22108 61684
rect 22440 61374 22516 61684
rect 114240 61336 114316 61646
rect 114648 61336 114724 61646
rect 115056 61336 115132 61646
rect 115600 61336 115676 61646
rect 115872 61374 115948 61684
rect 133416 61472 133492 64230
rect 134095 62091 134155 72326
rect 134776 70992 134852 71302
rect 134776 68582 134852 69164
rect 21352 60966 21428 61276
rect 22168 60966 22244 61276
rect 22440 60928 22516 61238
rect 22168 60520 22244 60830
rect 22576 60558 22652 60868
rect 109480 60830 109556 61140
rect 114240 60966 114316 61276
rect 114648 60966 114724 61276
rect 115328 60928 115404 61238
rect 114240 60558 114316 60868
rect 114648 60558 114724 60868
rect 20808 59878 20884 60188
rect 21896 60112 21972 60422
rect 22032 60112 22108 60422
rect 22440 60112 22516 60422
rect 114376 60150 114452 60460
rect 114648 60112 114724 60422
rect 115192 60150 115268 60460
rect 115328 60150 115404 60460
rect 20808 59432 20884 59742
rect 21760 59432 21836 59742
rect 27336 59606 27412 59916
rect 116008 59878 116084 60188
rect 109480 59568 109556 59878
rect 115464 59432 115540 59742
rect 116008 59432 116084 59742
rect 20808 59024 20884 59334
rect 22032 59024 22108 59334
rect 22440 59024 22516 59334
rect 114376 59062 114452 59372
rect 114784 59062 114860 59372
rect 115872 59062 115948 59372
rect 20808 58654 20884 58964
rect 21216 58616 21292 58926
rect 22168 58654 22244 58964
rect 22440 58654 22516 58964
rect 20808 58208 20884 58518
rect 21352 58208 21428 58518
rect 21760 58208 21836 58518
rect 22168 58208 22244 58518
rect 22440 58208 22516 58518
rect 27608 58344 27684 58654
rect 109480 58344 109556 58654
rect 114376 58616 114452 58926
rect 114784 58616 114860 58926
rect 115464 58654 115540 58964
rect 115872 58616 115948 58926
rect 114240 58208 114316 58518
rect 114784 58246 114860 58556
rect 115056 58208 115132 58518
rect 115328 58246 115404 58556
rect 116008 58208 116084 58518
rect 20944 57838 21020 58148
rect 21488 57838 21564 58148
rect 22032 57800 22108 58110
rect 22440 57800 22516 58110
rect 114376 57838 114452 58148
rect 114784 57800 114860 58110
rect 115192 57838 115268 58148
rect 115328 57838 115404 58148
rect 115872 57838 115948 58148
rect 20808 57392 20884 57702
rect 22168 57392 22244 57702
rect 22576 57430 22652 57740
rect 114240 57430 114316 57740
rect 114648 57430 114724 57740
rect 115600 57430 115676 57740
rect 116008 57392 116084 57702
rect 21216 57022 21292 57332
rect 21760 56984 21836 57294
rect 22032 57022 22108 57332
rect 22440 57022 22516 57332
rect 114240 56984 114316 57294
rect 114648 56984 114724 57294
rect 115192 57022 115268 57332
rect 115600 56984 115676 57294
rect 22032 56576 22108 56886
rect 22440 56576 22516 56886
rect 114240 56614 114316 56924
rect 114784 56576 114860 56886
rect 21352 56206 21428 56516
rect 21624 56206 21700 56516
rect 20944 55896 21020 56206
rect 22168 56168 22244 56478
rect 22440 56168 22516 56478
rect 114240 56168 114316 56478
rect 114648 56206 114724 56516
rect 115056 56206 115132 56516
rect 20808 55526 20884 55836
rect 21488 55526 21564 55836
rect 27472 55488 27548 55934
rect 109344 55624 109420 56070
rect 115192 56032 115404 56108
rect 115192 55934 115268 56032
rect 109480 55624 109556 55934
rect 116008 55896 116084 56206
rect 20944 55118 21020 55428
rect 27608 55216 27684 55526
rect 109480 55216 109556 55526
rect 115328 55488 115404 55798
rect 116008 55526 116084 55836
rect 116008 55080 116084 55390
rect 20808 54672 20884 54982
rect 21624 54710 21700 55020
rect 22032 54710 22108 55020
rect 22440 54672 22516 54982
rect 114376 54710 114452 55020
rect 114784 54710 114860 55020
rect 115192 54672 115268 54982
rect 115328 54710 115404 55020
rect 115872 54672 115948 54982
rect 20944 54302 21020 54612
rect 21352 54302 21428 54612
rect 21488 54302 21564 54612
rect 22168 54302 22244 54612
rect 22576 54264 22652 54574
rect 114240 54302 114316 54612
rect 114784 54264 114860 54574
rect 115464 54302 115540 54612
rect 116008 54302 116084 54612
rect 20808 53856 20884 54166
rect 21760 53856 21836 54166
rect 22168 53856 22244 54166
rect 22440 53894 22516 54204
rect 114376 53894 114452 54204
rect 114784 53894 114860 54204
rect 115192 53894 115268 54204
rect 115328 53894 115404 54204
rect 116008 53856 116084 54166
rect 20808 53448 20884 53758
rect 21624 53486 21700 53796
rect 22032 53448 22108 53758
rect 22440 53448 22516 53758
rect 114376 53448 114452 53758
rect 114784 53448 114860 53758
rect 115872 53486 115948 53796
rect 21352 53040 21428 53350
rect 21488 53040 21564 53350
rect 22168 53078 22244 53388
rect 22440 53040 22516 53350
rect 114240 53078 114316 53388
rect 114648 53040 114724 53350
rect 115464 53040 115540 53350
rect 20944 52632 21020 52942
rect 21216 52670 21292 52980
rect 21760 52632 21836 52942
rect 22168 52632 22244 52942
rect 22576 52670 22652 52980
rect 114240 52632 114316 52942
rect 114784 52670 114860 52980
rect 115192 52670 115268 52980
rect 115600 52670 115676 52980
rect 115872 52670 115948 52980
rect 22168 52262 22244 52572
rect 20808 51952 20884 52262
rect 22440 52224 22516 52534
rect 22168 51816 22244 52126
rect 22576 51854 22652 52164
rect 27472 52088 27548 52398
rect 114376 52224 114452 52534
rect 114784 52224 114860 52534
rect 115192 52224 115268 52534
rect 114240 51854 114316 52164
rect 114648 51854 114724 52164
rect 116008 51952 116084 52262
rect 21760 51446 21836 51756
rect 115192 51446 115268 51756
rect 20808 51136 20884 51446
rect 20808 50728 20884 51038
rect 21352 50728 21428 51038
rect 21896 50766 21972 51076
rect 22168 50728 22244 51038
rect 22576 50766 22652 51076
rect 27336 51000 27412 51310
rect 115872 51136 115948 51446
rect 114240 50766 114316 51076
rect 114648 50766 114724 51076
rect 115056 50766 115132 51076
rect 115464 50728 115540 51038
rect 116008 50728 116084 51038
rect 20808 50320 20884 50630
rect 21896 50320 21972 50630
rect 22032 50358 22108 50668
rect 22440 50320 22516 50630
rect 114376 50320 114452 50630
rect 114784 50358 114860 50668
rect 115872 50358 115948 50668
rect 20944 49912 21020 50222
rect 21216 49912 21292 50222
rect 21488 49950 21564 50260
rect 22168 49950 22244 50260
rect 22576 49912 22652 50222
rect 114240 49950 114316 50260
rect 114784 49912 114860 50222
rect 115600 49912 115676 50222
rect 115872 49912 115948 50222
rect 20808 49542 20884 49852
rect 21760 49504 21836 49814
rect 22168 49504 22244 49814
rect 22440 49542 22516 49852
rect 114240 49504 114316 49814
rect 114648 49504 114724 49814
rect 115192 49542 115268 49852
rect 115328 49542 115404 49852
rect 115872 49542 115948 49852
rect 20944 49134 21020 49444
rect 21216 49096 21292 49406
rect 21624 49134 21700 49444
rect 22032 49096 22108 49406
rect 22440 49096 22516 49406
rect 114376 49134 114452 49444
rect 114648 49134 114724 49444
rect 115872 49096 115948 49406
rect 20808 48688 20884 48998
rect 21352 48726 21428 49036
rect 21488 48726 21564 49036
rect 22168 48726 22244 49036
rect 22576 48726 22652 49036
rect 114240 48688 114316 48998
rect 114648 48726 114724 49036
rect 115600 48726 115676 49036
rect 116008 48688 116084 48998
rect 20808 48008 20884 48318
rect 21760 48280 21836 48590
rect 22168 48280 22244 48590
rect 22440 48318 22516 48628
rect 114376 48318 114452 48628
rect 114648 48280 114724 48590
rect 115056 48280 115132 48590
rect 115464 48318 115540 48628
rect 22168 47910 22244 48220
rect 22440 47910 22516 48220
rect 114240 47910 114316 48220
rect 114784 47872 114860 48182
rect 115328 48008 115404 48318
rect 115872 48008 115948 48318
rect 20808 47230 20884 47540
rect 21488 47464 21564 47774
rect 115056 47502 115132 47812
rect 20944 46784 21020 47094
rect 21352 46822 21428 47132
rect 21760 46784 21836 47094
rect 27336 46958 27412 47268
rect 115872 47230 115948 47540
rect 109344 46920 109420 47230
rect 20808 46376 20884 46686
rect 22168 46376 22244 46686
rect 22576 46414 22652 46724
rect 27336 46550 27412 46860
rect 109480 46550 109556 46860
rect 115328 46784 115404 47094
rect 115872 46784 115948 47094
rect 114240 46414 114316 46724
rect 114648 46414 114724 46724
rect 116008 46414 116084 46724
rect 20944 46006 21020 46316
rect 21216 45968 21292 46278
rect 22032 46006 22108 46316
rect 22576 46006 22652 46316
rect 114376 45968 114452 46278
rect 114784 45968 114860 46278
rect 115192 45968 115268 46278
rect 115328 46006 115404 46316
rect 115464 45968 115540 46278
rect 115872 45968 115948 46278
rect 20944 45560 21020 45870
rect 21352 45598 21428 45908
rect 22032 45560 22108 45870
rect 22440 45598 22516 45908
rect 114376 45560 114452 45870
rect 114648 45598 114724 45908
rect 115464 45598 115540 45908
rect 116008 45598 116084 45908
rect 20808 45152 20884 45462
rect 21760 45190 21836 45500
rect 22032 45190 22108 45500
rect 22440 45152 22516 45462
rect 25840 45190 25916 45500
rect 113696 45190 113772 45500
rect 114376 45190 114452 45500
rect 114784 45190 114860 45500
rect 115192 45190 115268 45500
rect 115328 45190 115404 45500
rect 115872 45190 115948 45500
rect 20944 44782 21020 45092
rect 21216 44782 21292 45092
rect 21488 44782 21564 45092
rect 22032 44782 22108 45092
rect 22576 44782 22652 45092
rect 23256 44782 23332 45092
rect 21352 44336 21428 44646
rect 22168 44374 22244 44684
rect 112336 44646 112412 45092
rect 114376 44744 114452 45054
rect 114648 44782 114724 45092
rect 115872 44782 115948 45092
rect 22440 44336 22516 44646
rect 114240 44374 114316 44684
rect 114648 44336 114724 44646
rect 115464 44336 115540 44646
rect 22168 43928 22244 44238
rect 22576 43928 22652 44238
rect 114376 43966 114452 44276
rect 114784 43966 114860 44276
rect 21760 43558 21836 43868
rect 20808 43248 20884 43558
rect 22032 43520 22108 43830
rect 22440 43520 22516 43830
rect 21488 43384 21700 43460
rect 27472 43384 27548 43694
rect 109344 43384 109420 43694
rect 114376 43520 114452 43830
rect 114784 43520 114860 43830
rect 115192 43520 115268 43830
rect 20808 42878 20884 43188
rect 21216 42878 21292 43188
rect 21488 43150 21564 43384
rect 27608 42976 27684 43286
rect 109344 43014 109420 43324
rect 116008 43286 116084 43596
rect 20808 42432 20884 42742
rect 22168 42470 22244 42780
rect 22440 42470 22516 42780
rect 109344 42568 109420 42878
rect 115056 42840 115132 43150
rect 116008 42840 116084 43150
rect 114240 42470 114316 42780
rect 114784 42432 114860 42742
rect 115872 42432 115948 42742
rect 20944 42062 21020 42372
rect 21760 42024 21836 42334
rect 22168 42024 22244 42334
rect 22576 42062 22652 42372
rect 114240 42062 114316 42372
rect 114648 42062 114724 42372
rect 115056 42062 115132 42372
rect 116008 42024 116084 42334
rect 20808 41616 20884 41926
rect 21216 41616 21292 41926
rect 21624 41654 21700 41964
rect 22032 41654 22108 41964
rect 22440 41616 22516 41926
rect 114376 41616 114452 41926
rect 114784 41654 114860 41964
rect 115192 41654 115268 41964
rect 115328 41654 115404 41964
rect 115872 41654 115948 41964
rect 20808 41246 20884 41556
rect 21352 41246 21428 41556
rect 22032 41208 22108 41518
rect 22576 41208 22652 41518
rect 114376 41208 114452 41518
rect 114784 41208 114860 41518
rect 115600 41208 115676 41518
rect 116008 41246 116084 41556
rect 20808 40800 20884 41110
rect 21760 40800 21836 41110
rect 22032 40838 22108 41148
rect 22440 40800 22516 41110
rect 114376 40838 114452 41148
rect 114648 40800 114724 41110
rect 115192 40838 115268 41148
rect 115328 40838 115404 41148
rect 115464 40838 115540 41148
rect 116008 40800 116084 41110
rect 21216 40392 21292 40702
rect 21624 40430 21700 40740
rect 22032 40392 22108 40702
rect 22576 40430 22652 40740
rect 22168 39984 22244 40294
rect 22440 39984 22516 40294
rect 27472 40256 27548 40566
rect 109480 40294 109556 40604
rect 114376 40392 114452 40702
rect 114648 40430 114724 40740
rect 115328 40430 115404 40740
rect 20808 39304 20884 39614
rect 21760 39576 21836 39886
rect 22032 39614 22108 39924
rect 22576 39614 22652 39924
rect 109344 39848 109420 40294
rect 114240 40022 114316 40332
rect 114648 40022 114724 40332
rect 115192 40196 115268 40294
rect 115192 40120 115404 40196
rect 114240 39576 114316 39886
rect 114648 39576 114724 39886
rect 115192 39614 115268 39924
rect 20808 38896 20884 39206
rect 21488 38934 21564 39244
rect 27472 39070 27548 39380
rect 109480 39070 109556 39380
rect 115872 39342 115948 39652
rect 115464 38896 115540 39206
rect 116008 38934 116084 39244
rect 20808 38526 20884 38836
rect 116008 38488 116084 38798
rect 20808 38080 20884 38390
rect 21352 38118 21428 38428
rect 22032 38080 22108 38390
rect 22440 38118 22516 38428
rect 20944 37710 21020 38020
rect 21760 37672 21836 37982
rect 22168 37710 22244 38020
rect 22440 37672 22516 37982
rect 27336 37846 27412 38156
rect 109480 37808 109556 38118
rect 114376 38080 114452 38390
rect 114648 38118 114724 38428
rect 115192 38080 115268 38390
rect 115328 38080 115404 38390
rect 115872 38080 115948 38390
rect 114240 37710 114316 38020
rect 114648 37672 114724 37982
rect 115056 37710 115132 38020
rect 115464 37672 115540 37982
rect 116008 37672 116084 37982
rect 14144 34854 14220 37612
rect 20808 37264 20884 37574
rect 21216 37264 21292 37574
rect 21624 37302 21700 37612
rect 22032 37264 22108 37574
rect 22576 37302 22652 37612
rect 114376 37302 114452 37612
rect 114784 37302 114860 37612
rect 115872 37302 115948 37612
rect 20808 36894 20884 37204
rect 21352 36894 21428 37204
rect 21488 36894 21564 37204
rect 22168 36894 22244 37204
rect 22576 36856 22652 37166
rect 114240 36894 114316 37204
rect 114784 36856 114860 37166
rect 115600 36856 115676 37166
rect 115872 36856 115948 37166
rect 21760 36448 21836 36758
rect 22032 36486 22108 36796
rect 22440 36486 22516 36796
rect 114240 36448 114316 36758
rect 114648 36448 114724 36758
rect 115192 36486 115268 36796
rect 115464 36486 115540 36796
rect 14008 32134 14084 34756
rect 14280 33494 14356 36252
rect 20944 36040 21020 36350
rect 21488 36040 21564 36350
rect 21624 36078 21700 36388
rect 22032 36040 22108 36350
rect 22440 36040 22516 36350
rect 114376 36078 114452 36388
rect 114784 36078 114860 36388
rect 115192 36078 115268 36388
rect 115328 36078 115404 36388
rect 116008 36040 116084 36350
rect 20808 35398 20884 35708
rect 21488 35632 21564 35942
rect 22168 35670 22244 35980
rect 22440 35632 22516 35942
rect 114240 35632 114316 35942
rect 114648 35670 114724 35980
rect 115464 35632 115540 35942
rect 21390 35496 21700 35572
rect 115872 35398 115948 35708
rect 20944 34990 21020 35300
rect 20808 34544 20884 34854
rect 21896 34816 21972 35262
rect 27472 34990 27548 35300
rect 109344 34718 109420 35028
rect 115464 34854 115540 35300
rect 115872 34990 115948 35300
rect 20808 34174 20884 34484
rect 21216 34174 21292 34484
rect 22032 34174 22108 34484
rect 22440 34174 22516 34484
rect 109480 34408 109556 34718
rect 116008 34544 116084 34854
rect 20808 33728 20884 34038
rect 21352 33766 21428 34076
rect 22032 33728 22108 34038
rect 22440 33766 22516 34076
rect 109480 33864 109556 34174
rect 114240 34136 114316 34446
rect 114648 34136 114724 34446
rect 115192 34174 115268 34484
rect 115600 34136 115676 34446
rect 116008 34136 116084 34446
rect 114240 33766 114316 34076
rect 114784 33728 114860 34038
rect 115328 33728 115404 34038
rect 115600 33728 115676 34038
rect 116008 33766 116084 34076
rect 14144 32036 14220 33396
rect 20808 33320 20884 33630
rect 21352 33320 21428 33630
rect 21760 33320 21836 33630
rect 22168 33320 22244 33630
rect 22440 33320 22516 33630
rect 114240 33320 114316 33630
rect 114648 33358 114724 33668
rect 115056 33320 115132 33630
rect 115600 33358 115676 33668
rect 116008 33320 116084 33630
rect 20808 32912 20884 33222
rect 21624 32950 21700 33260
rect 22032 32950 22108 33260
rect 22440 32912 22516 33222
rect 114376 32950 114452 33260
rect 114784 32950 114860 33260
rect 115192 32950 115268 33260
rect 115872 32950 115948 33260
rect 20944 32542 21020 32852
rect 21216 32504 21292 32814
rect 22032 32504 22108 32814
rect 22576 32504 22652 32814
rect 114376 32504 114452 32814
rect 114784 32504 114860 32814
rect 115600 32504 115676 32814
rect 115872 32504 115948 32814
rect 20944 32096 21020 32406
rect 21760 32096 21836 32406
rect 22032 32134 22108 32444
rect 22440 32096 22516 32406
rect 114240 32096 114316 32406
rect 114648 32096 114724 32406
rect 115192 32134 115268 32444
rect 115328 32134 115404 32444
rect 115872 32134 115948 32444
rect 14008 31960 14220 32036
rect 14008 30638 14084 31960
rect 14008 27782 14084 30540
rect 14144 29240 14220 31862
rect 20944 31416 21020 31726
rect 21216 31688 21292 31998
rect 21624 31688 21700 31998
rect 22032 31688 22108 31998
rect 22576 31726 22652 32036
rect 109480 31590 109556 31900
rect 114376 31726 114452 32036
rect 114784 31726 114860 32036
rect 22168 31280 22244 31590
rect 22440 31280 22516 31590
rect 20808 30600 20884 30910
rect 21760 30872 21836 31182
rect 109344 31144 109420 31590
rect 114240 31280 114316 31590
rect 114648 31280 114724 31590
rect 115872 31454 115948 31764
rect 27336 30736 27412 31046
rect 115464 30910 115540 31220
rect 115872 30638 115948 30948
rect 20808 30192 20884 30502
rect 21352 30230 21428 30540
rect 27472 30328 27548 30638
rect 109344 30328 109420 30638
rect 20944 29784 21020 30094
rect 22168 29784 22244 30094
rect 22576 29784 22652 30094
rect 109344 29958 109420 30268
rect 115464 30192 115540 30502
rect 116008 30230 116084 30540
rect 114240 29784 114316 30094
rect 114648 29784 114724 30094
rect 115872 29822 115948 30132
rect 20808 29414 20884 29724
rect 21488 29414 21564 29724
rect 21760 29376 21836 29686
rect 22032 29376 22108 29686
rect 22440 29414 22516 29724
rect 114240 29414 114316 29724
rect 114648 29414 114724 29724
rect 115328 29376 115404 29686
rect 115464 29414 115540 29724
rect 115872 29376 115948 29686
rect 2312 23974 2388 24556
rect 2539 17926 2599 25333
rect 3808 23294 3884 25916
rect 15912 25024 15988 27646
rect 17816 27472 17892 29142
rect 20808 28968 20884 29278
rect 21760 28968 21836 29278
rect 22168 29006 22244 29316
rect 22576 29006 22652 29316
rect 114240 28968 114316 29278
rect 114648 28968 114724 29278
rect 115056 28968 115132 29278
rect 115328 29006 115404 29316
rect 116008 29006 116084 29316
rect 20944 28598 21020 28908
rect 21216 28560 21292 28870
rect 21624 28598 21700 28908
rect 22032 28560 22108 28870
rect 22576 28598 22652 28908
rect 114376 28598 114452 28908
rect 114784 28598 114860 28908
rect 115192 28598 115268 28908
rect 115872 28560 115948 28870
rect 20944 28152 21020 28462
rect 21352 28190 21428 28500
rect 21488 28190 21564 28500
rect 22168 28190 22244 28500
rect 22440 28190 22516 28500
rect 114376 28152 114452 28462
rect 114784 28152 114860 28462
rect 115600 28152 115676 28462
rect 115872 28152 115948 28462
rect 18904 27374 18980 28092
rect 21760 27782 21836 28092
rect 22032 27782 22108 28092
rect 22440 27744 22516 28054
rect 114376 27782 114452 28092
rect 114784 27782 114860 28092
rect 115192 27782 115268 28092
rect 22032 27336 22108 27646
rect 22576 27374 22652 27684
rect 114376 27374 114452 27684
rect 114784 27374 114860 27684
rect 17408 26656 17484 27238
rect 18360 26694 18436 27276
rect 18632 26694 18708 27276
rect 19040 26694 19116 27276
rect 20672 26792 20748 27238
rect 20808 26694 20884 27004
rect 21352 26966 21428 27276
rect 21488 26966 21564 27276
rect 115600 26928 115676 27238
rect 115736 26792 115812 27238
rect 17544 25840 17620 26558
rect 17680 26248 17756 26558
rect 18224 25840 18300 26422
rect 18632 25840 18708 26422
rect 20808 26248 20884 26558
rect 21216 26248 21292 26558
rect 21896 26286 21972 26596
rect 27336 26384 27412 26694
rect 109344 26422 109420 26732
rect 115872 26694 115948 27004
rect 117640 26830 117716 27276
rect 117776 26656 117852 27238
rect 118184 26694 118260 27276
rect 118728 27200 118940 27276
rect 118728 26694 118804 27200
rect 119272 26694 119348 27276
rect 20808 25840 20884 26150
rect 22168 25878 22244 26188
rect 22576 25878 22652 26188
rect 27472 25976 27548 26286
rect 109344 25976 109420 26286
rect 115464 26248 115540 26558
rect 115872 26248 115948 26558
rect 114240 25878 114316 26188
rect 114648 25878 114724 26188
rect 116008 25878 116084 26188
rect 117640 25840 117716 26422
rect 118184 25840 118260 26422
rect 119000 25878 119076 26596
rect 119272 25840 119348 26558
rect 17408 25062 17484 25780
rect 18224 25024 18300 25742
rect 18768 25024 18844 25742
rect 19176 25062 19252 25780
rect 20808 25470 20884 25780
rect 22168 25432 22244 25742
rect 22576 25470 22652 25780
rect 114240 25432 114316 25742
rect 114784 25470 114860 25780
rect 115056 25432 115132 25742
rect 115600 25432 115676 25742
rect 116008 25432 116084 25742
rect 20808 25062 20884 25372
rect 21352 25062 21428 25372
rect 21488 25062 21564 25372
rect 21760 25024 21836 25334
rect 22168 25062 22244 25372
rect 22440 25024 22516 25334
rect 114240 25062 114316 25372
rect 114648 25062 114724 25372
rect 115192 25024 115268 25334
rect 115464 25062 115540 25372
rect 115872 25024 115948 25334
rect 117640 25062 117716 25780
rect 118184 25062 118260 25780
rect 119000 25062 119076 25780
rect 119408 25024 119484 25742
rect 120768 25024 120844 25742
rect 17680 23392 17756 24926
rect 18224 23392 18300 24926
rect 20808 24616 20884 24926
rect 21896 24654 21972 24964
rect 22168 24616 22244 24926
rect 22576 24654 22652 24964
rect 114240 24616 114316 24926
rect 114648 24616 114724 24926
rect 115056 24654 115132 24964
rect 115464 24616 115540 24926
rect 116008 24654 116084 24964
rect 20944 24246 21020 24556
rect 21624 24246 21700 24556
rect 22032 24246 22108 24556
rect 22440 24208 22516 24518
rect 114376 24208 114452 24518
rect 114784 24246 114860 24556
rect 115872 24208 115948 24518
rect 21216 23800 21292 24110
rect 21488 23838 21564 24148
rect 22032 23800 22108 24110
rect 22440 23838 22516 24148
rect 22168 23392 22244 23702
rect 22440 23430 22516 23740
rect 27608 23702 27684 24012
rect 114240 23838 114316 24148
rect 114784 23800 114860 24110
rect 115192 23800 115268 24110
rect 115600 23800 115676 24110
rect 3128 21760 3204 22206
rect 3672 17544 3748 20438
rect 3808 20400 3884 23158
rect 18224 22750 18300 23332
rect 18632 22750 18708 23332
rect 19040 22712 19116 23294
rect 20944 22712 21020 23022
rect 21352 22984 21428 23294
rect 21488 22712 21564 23022
rect 21624 22984 21700 23294
rect 22032 23022 22108 23332
rect 22576 23022 22652 23332
rect 27472 23256 27548 23702
rect 114240 23392 114316 23702
rect 114784 23430 114860 23740
rect 117640 23430 117716 24964
rect 118184 23392 118260 24926
rect 27336 22886 27412 23196
rect 109344 22848 109420 23158
rect 114376 22984 114452 23294
rect 114784 22984 114860 23294
rect 18360 21118 18436 22516
rect 18632 21118 18708 22516
rect 20808 22304 20884 22614
rect 21624 22342 21700 22652
rect 27472 22478 27548 22788
rect 109480 22478 109556 22788
rect 116008 22750 116084 23060
rect 117640 22750 117716 23332
rect 118048 22750 118124 23332
rect 118320 22750 118396 23060
rect 118592 22750 118668 23332
rect 118864 22712 118940 23022
rect 119000 22712 119076 23294
rect 20944 21934 21020 22244
rect 27336 22032 27412 22342
rect 109344 22070 109420 22380
rect 115056 22304 115132 22614
rect 115872 22342 115948 22652
rect 115872 21896 115948 22206
rect 20944 21526 21020 21836
rect 21352 21526 21428 21836
rect 21488 21526 21564 21836
rect 21760 21526 21836 21836
rect 22168 21526 22244 21836
rect 22440 21488 22516 21798
rect 20944 21080 21020 21390
rect 21624 21080 21700 21390
rect 22168 21080 22244 21390
rect 22440 21118 22516 21428
rect 109344 21254 109420 21564
rect 114240 21488 114316 21798
rect 114648 21526 114724 21836
rect 115056 21488 115132 21798
rect 115600 21526 115676 21836
rect 116008 21488 116084 21798
rect 114240 21080 114316 21390
rect 114648 21080 114724 21390
rect 115600 21080 115676 21390
rect 115872 21118 115948 21428
rect 118048 21080 118124 21390
rect 118320 21118 118396 22244
rect 118456 21254 118532 22516
rect 118864 22206 118940 22516
rect 17816 20302 17892 21020
rect 18360 20264 18436 20982
rect 18632 20264 18708 20982
rect 19176 20302 19252 21020
rect 20808 20672 20884 20982
rect 21352 20710 21428 21020
rect 21760 20672 21836 20982
rect 22032 20672 22108 20982
rect 22440 20672 22516 20982
rect 114240 20710 114316 21020
rect 114648 20710 114724 21020
rect 115192 20672 115268 20982
rect 115328 20672 115404 20982
rect 116008 20710 116084 21020
rect 20944 20302 21020 20612
rect 21352 20264 21428 20574
rect 21760 20264 21836 20574
rect 22168 20302 22244 20612
rect 22440 20264 22516 20574
rect 114240 20302 114316 20612
rect 114648 20302 114724 20612
rect 115056 20302 115132 20612
rect 115464 20264 115540 20574
rect 116008 20264 116084 20574
rect 117640 20264 117716 20982
rect 118184 20302 118260 21020
rect 118592 20302 118668 21020
rect 119000 20302 119076 21020
rect 16592 19078 16668 20204
rect 3128 15542 3204 16124
rect 14552 14726 14628 17484
rect 14688 16184 14764 18806
rect 17000 17582 17076 20204
rect 21080 17348 21156 20166
rect 22440 19720 22516 20166
rect 21080 17272 21292 17348
rect 3128 13328 3204 13774
rect 14552 11968 14628 14590
rect 14688 13366 14764 16124
rect 14552 9150 14628 11772
rect 14688 10510 14764 13268
rect 20264 11734 20340 14356
rect 21216 13056 21292 15814
rect 21352 14552 21428 17174
rect 22440 15814 22516 19660
rect 26928 19312 27004 19622
rect 28288 18768 28364 19214
rect 28560 18768 28636 19214
rect 28968 17136 29044 19758
rect 109616 19720 109692 20030
rect 29512 18768 29588 19214
rect 30736 18768 30812 19214
rect 32504 18806 32580 19252
rect 33184 18768 33260 19214
rect 33728 18806 33804 19252
rect 34544 18768 34620 19214
rect 35632 18768 35708 19214
rect 37264 18768 37340 19214
rect 38216 18768 38292 19214
rect 38760 18806 38836 19252
rect 39440 18768 39516 19214
rect 39984 18806 40060 19252
rect 40664 18768 40740 19214
rect 41208 18806 41284 19252
rect 42024 18768 42100 19214
rect 42432 18806 42508 19252
rect 43248 18768 43324 19214
rect 43384 18806 43460 19252
rect 44472 18768 44548 19214
rect 45696 18768 45772 19214
rect 46920 18768 46996 19214
rect 47464 18806 47540 19252
rect 48144 18768 48220 19214
rect 49912 18806 49988 19252
rect 51272 18806 51348 19252
rect 51952 18768 52028 19214
rect 53176 18768 53252 19214
rect 53720 18806 53796 19252
rect 54400 18768 54476 19214
rect 54944 18806 55020 19252
rect 55624 18768 55700 19214
rect 56168 18806 56244 19252
rect 57392 18806 57468 19252
rect 58208 18768 58284 19214
rect 59432 18768 59508 19214
rect 59976 18806 60052 19252
rect 60656 18768 60732 19214
rect 60792 18806 60868 19252
rect 61880 18768 61956 19214
rect 62424 18806 62500 19252
rect 63104 18768 63180 19214
rect 64464 18768 64540 19214
rect 66232 18806 66308 19252
rect 66912 18768 66988 19214
rect 67456 18806 67532 19252
rect 68680 18806 68756 19252
rect 69360 18768 69436 19214
rect 70992 18768 71068 19214
rect 71944 18768 72020 19214
rect 72352 18806 72428 19252
rect 73168 18768 73244 19214
rect 74936 18806 75012 19252
rect 75616 18768 75692 19214
rect 76160 18806 76236 19252
rect 77384 18806 77460 19252
rect 78064 18768 78140 19214
rect 79696 18768 79772 19214
rect 80648 18768 80724 19214
rect 81192 18806 81268 19252
rect 81872 18768 81948 19214
rect 83640 18806 83716 19252
rect 84320 18768 84396 19214
rect 84864 18806 84940 19252
rect 86088 18806 86164 19252
rect 86904 18768 86980 19214
rect 87312 18806 87388 19252
rect 88128 18768 88204 19214
rect 88264 18806 88340 19252
rect 89352 18768 89428 19214
rect 89896 18806 89972 19252
rect 90712 18768 90788 19214
rect 91800 18768 91876 19214
rect 92344 18806 92420 19252
rect 93432 18768 93508 19214
rect 94520 18806 94596 19388
rect 95608 18768 95684 19214
rect 96152 18806 96228 19252
rect 96832 18768 96908 19214
rect 98192 18768 98268 19214
rect 98600 18806 98676 19252
rect 99824 18806 99900 19252
rect 101184 18806 101260 19252
rect 101864 18768 101940 19214
rect 102408 18806 102484 19252
rect 103088 18768 103164 19214
rect 104312 18768 104388 19214
rect 104856 18806 104932 19252
rect 105536 18768 105612 19214
rect 105808 18806 105884 19252
rect 107168 18768 107244 19214
rect 107304 18806 107380 19252
rect 108528 18806 108604 19252
rect 28968 15134 29044 17076
rect 28832 13600 28908 14318
rect 14688 7654 14764 10412
rect 28152 9558 28228 11364
rect 16320 3808 16396 9014
rect 2040 1224 2116 1670
rect 3808 1224 3884 1670
rect 5576 1224 5652 1670
rect 7072 1224 7148 1670
rect 8704 1224 8780 1670
rect 10472 1224 10548 1670
rect 12104 1224 12180 1670
rect 14008 1224 14084 1670
rect 15504 1224 15580 1670
rect 16048 0 16124 2894
rect 17136 0 17212 2894
rect 17408 1224 17484 1670
rect 18224 0 18300 2894
rect 19040 1224 19116 1670
rect 19584 0 19660 2894
rect 20264 1768 20340 3710
rect 20536 0 20612 2894
rect 20808 1224 20884 1670
rect 21760 0 21836 2894
rect 22168 1224 22244 1670
rect 23120 0 23196 2894
rect 23936 1224 24012 1670
rect 24208 0 24284 2894
rect 25432 0 25508 2894
rect 25704 1224 25780 1670
rect 26520 0 26596 2894
rect 27336 1224 27412 1670
rect 27608 0 27684 2894
rect 28288 0 28364 13094
rect 28560 10646 28636 11092
rect 28696 11016 28772 11870
rect 28832 11696 28908 12278
rect 28968 12006 29044 13540
rect 29104 13230 29180 15172
rect 31416 13600 31492 14318
rect 29104 12550 29180 13132
rect 28696 0 28772 2894
rect 28968 1224 29044 1670
rect 30056 0 30132 2894
rect 30464 1224 30540 1670
rect 30736 0 30812 13094
rect 31280 12006 31356 13540
rect 31552 13230 31628 15172
rect 31688 15134 31764 17076
rect 34000 15134 34076 17076
rect 33592 13638 33668 14356
rect 33864 13600 33940 14318
rect 31416 12550 31492 13132
rect 31144 11016 31220 11870
rect 31416 11696 31492 12278
rect 33456 11696 33532 12278
rect 31280 0 31356 2894
rect 32096 1224 32172 1670
rect 32368 0 32444 2894
rect 33456 0 33532 2894
rect 33592 0 33668 13094
rect 33864 12550 33940 13132
rect 34000 12006 34076 13540
rect 34136 13230 34212 15172
rect 36448 15134 36524 17076
rect 36448 13600 36524 14318
rect 33864 11016 33940 11870
rect 34000 1224 34076 1670
rect 34544 0 34620 2894
rect 35768 1224 35844 1670
rect 35904 0 35980 2894
rect 36040 0 36116 13094
rect 36176 11696 36252 12278
rect 36448 12006 36524 13540
rect 36584 13230 36660 15172
rect 38896 13600 38972 14318
rect 36584 12550 36660 13132
rect 36312 11016 36388 11870
rect 36992 0 37068 2894
rect 37400 1224 37476 1670
rect 38080 0 38156 2894
rect 38488 0 38564 13094
rect 38624 11696 38700 12278
rect 38896 12006 38972 13540
rect 39032 13230 39108 15172
rect 39168 15134 39244 17076
rect 41072 13600 41148 14318
rect 41208 13600 41284 14318
rect 39032 12550 39108 13132
rect 38760 11016 38836 11870
rect 39168 1224 39244 1670
rect 39440 0 39516 2894
rect 39712 544 39788 2350
rect 40664 0 40740 2894
rect 40800 1224 40876 1670
rect 41072 0 41148 13094
rect 41344 12006 41420 13540
rect 41480 13230 41556 15172
rect 41616 15134 41692 17076
rect 43928 17000 44140 17076
rect 43928 15134 44004 17000
rect 43792 13600 43868 14318
rect 41480 12550 41556 13132
rect 41344 11016 41420 11870
rect 41480 11696 41556 12278
rect 43384 11462 43460 12316
rect 41752 0 41828 2894
rect 42432 1224 42508 1670
rect 42840 0 42916 2894
rect 43520 0 43596 13094
rect 43928 12006 44004 13540
rect 44064 13230 44140 15172
rect 46240 13600 46316 14318
rect 44064 12550 44140 13132
rect 43792 11016 43868 11870
rect 43928 0 44004 2894
rect 44200 1224 44276 1670
rect 45288 0 45364 2894
rect 45696 1224 45772 1670
rect 45968 0 46044 13094
rect 46376 12006 46452 13540
rect 46512 13230 46588 15172
rect 46648 15134 46724 17076
rect 48960 15134 49036 17076
rect 51408 17000 51620 17076
rect 48824 13600 48900 14318
rect 46512 12550 46588 13132
rect 46240 11016 46316 11870
rect 46512 11696 46588 12278
rect 46376 0 46452 2894
rect 47328 1224 47404 1670
rect 47600 0 47676 2894
rect 48280 0 48356 13094
rect 48824 12550 48900 13132
rect 48688 11016 48764 11870
rect 48824 11696 48900 12278
rect 48960 12006 49036 13540
rect 49096 13230 49172 15172
rect 51408 15134 51484 17000
rect 51408 13600 51484 14318
rect 48688 0 48764 2894
rect 49096 1224 49172 1670
rect 49776 0 49852 2894
rect 50728 1224 50804 1670
rect 51000 0 51076 13094
rect 51136 11016 51212 11870
rect 51272 11696 51348 12278
rect 51408 12006 51484 13540
rect 51544 13230 51620 15172
rect 53856 13600 53932 14318
rect 51544 12550 51620 13132
rect 51136 0 51212 2894
rect 52224 0 52300 2894
rect 52496 1224 52572 1670
rect 53312 0 53388 2894
rect 53584 0 53660 13094
rect 53856 12006 53932 13540
rect 53992 13230 54068 15172
rect 54128 15134 54204 17076
rect 56440 15134 56516 17076
rect 56440 13600 56516 14318
rect 53992 12550 54068 13132
rect 53856 11016 53932 11870
rect 53992 11696 54068 12278
rect 54128 1224 54204 1670
rect 54400 0 54476 2894
rect 55488 1224 55564 1670
rect 55760 0 55836 2894
rect 56032 0 56108 13094
rect 56304 12006 56380 13540
rect 56576 13230 56652 15172
rect 58344 14416 58420 18670
rect 119952 18496 120028 20166
rect 122808 19856 122884 20166
rect 58616 13638 58692 14356
rect 58888 13600 58964 14318
rect 56440 12550 56516 13132
rect 56304 11016 56380 11870
rect 56440 11696 56516 12278
rect 56984 0 57060 2894
rect 57528 1224 57604 1670
rect 58072 0 58148 2894
rect 58480 0 58556 13094
rect 58888 12006 58964 13540
rect 59024 13230 59100 15172
rect 59160 15134 59236 17076
rect 61064 13638 61140 14356
rect 59024 12550 59100 13132
rect 58752 11016 58828 11870
rect 59024 11696 59100 12278
rect 59160 0 59236 2894
rect 59432 1224 59508 1670
rect 60792 1224 60868 1670
rect 60928 0 61004 13094
rect 61200 12006 61276 13676
rect 61336 13600 61412 14318
rect 61336 12550 61412 13132
rect 61472 13094 61548 15172
rect 61608 15134 61684 17076
rect 63920 15134 63996 17076
rect 63648 13638 63724 14356
rect 63784 13600 63860 14318
rect 61200 11016 61276 11870
rect 61336 11696 61412 12278
rect 62560 1224 62636 1670
rect 63512 0 63588 13094
rect 63648 11696 63724 12278
rect 63920 12006 63996 13540
rect 64056 13230 64132 15172
rect 66232 13600 66308 14318
rect 64056 12550 64132 13132
rect 63784 11016 63860 11870
rect 64328 1224 64404 1670
rect 65824 1224 65900 1670
rect 65960 0 66036 13094
rect 66096 11016 66172 11870
rect 66232 11696 66308 12278
rect 66368 12006 66444 13540
rect 66504 13230 66580 15172
rect 66640 15134 66716 17076
rect 66504 12550 66580 13132
rect 67592 1224 67668 1670
rect 68272 0 68348 13094
rect 68544 11696 68620 12278
rect 68680 12006 68756 13676
rect 68816 13600 68892 14318
rect 68816 12550 68892 13132
rect 68952 13094 69028 15172
rect 69088 15134 69164 17076
rect 71400 15134 71476 17076
rect 71264 13600 71340 14318
rect 68816 11016 68892 11870
rect 69224 1224 69300 1670
rect 70856 1224 70932 1670
rect 70992 0 71068 13094
rect 71400 12006 71476 13540
rect 71536 13230 71612 15172
rect 73848 13600 73924 14318
rect 71536 12550 71612 13132
rect 71264 11016 71340 11870
rect 71536 11696 71612 12278
rect 73304 11462 73380 12316
rect 72760 1224 72836 1670
rect 73440 0 73516 13094
rect 73848 12006 73924 13540
rect 73984 13230 74060 15172
rect 74120 15134 74196 17076
rect 76432 15134 76508 17076
rect 76024 13638 76100 14356
rect 76296 13600 76372 14318
rect 73984 12550 74060 13132
rect 73712 11016 73788 11870
rect 74256 1224 74332 1670
rect 75888 0 75964 13094
rect 76296 12550 76372 13132
rect 76160 11696 76236 12278
rect 76432 12006 76508 13540
rect 76568 13230 76644 15172
rect 78880 15134 78956 17076
rect 78880 13600 78956 14318
rect 76296 11016 76372 11870
rect 76160 1224 76236 1670
rect 77656 1224 77732 1670
rect 78472 0 78548 13094
rect 78608 11696 78684 12278
rect 78880 12006 78956 13540
rect 79016 13230 79092 15172
rect 81328 13600 81404 14318
rect 79016 12550 79092 13132
rect 78744 11016 78820 11870
rect 79288 1224 79364 1670
rect 80920 0 80996 13094
rect 81056 11696 81132 12278
rect 81328 12006 81404 13540
rect 81464 13230 81540 15172
rect 81600 15134 81676 17076
rect 83912 15134 83988 17076
rect 83640 13600 83716 14318
rect 81464 12550 81540 13132
rect 81192 11016 81268 11870
rect 81056 1224 81132 1670
rect 82824 1224 82900 1670
rect 83504 0 83580 13094
rect 83776 12550 83852 13132
rect 83912 12006 83988 13540
rect 84048 13230 84124 15172
rect 86360 15134 86436 17076
rect 86088 13638 86164 14356
rect 86224 13600 86300 14318
rect 83776 11016 83852 11870
rect 84048 11696 84124 12278
rect 84320 1224 84396 1670
rect 85952 0 86028 13094
rect 86360 12006 86436 13540
rect 86496 13230 86572 15172
rect 88672 13600 88748 14318
rect 86496 12550 86572 13132
rect 86224 11016 86300 11870
rect 86496 11696 86572 12278
rect 86224 1224 86300 1670
rect 87720 1224 87796 1670
rect 88536 0 88612 13094
rect 88808 12006 88884 13540
rect 88944 13230 89020 15172
rect 89080 15134 89156 17076
rect 91392 15134 91468 17076
rect 93840 17000 94052 17076
rect 91256 13600 91332 14318
rect 88944 12550 89020 13132
rect 88808 11016 88884 11870
rect 88944 11696 89020 12278
rect 89352 1224 89428 1670
rect 90984 0 91060 13094
rect 91256 12550 91332 13132
rect 91120 11016 91196 11870
rect 91256 11696 91332 12278
rect 91392 12006 91468 13540
rect 91528 13230 91604 15172
rect 93840 15134 93916 17000
rect 93840 13600 93916 14318
rect 91256 1224 91332 1670
rect 92752 1224 92828 1670
rect 93432 0 93508 13094
rect 93568 11016 93644 11870
rect 93704 11462 93780 12316
rect 93840 12006 93916 13540
rect 93976 13230 94052 15172
rect 96288 13600 96364 14318
rect 93976 12550 94052 13132
rect 94384 1224 94460 1670
rect 95880 0 95956 13094
rect 96016 11696 96092 12278
rect 96288 12006 96364 13540
rect 96424 13230 96500 15172
rect 96560 15134 96636 17076
rect 98872 15134 98948 17076
rect 98872 13600 98948 14318
rect 96424 12550 96500 13132
rect 96152 11016 96228 11870
rect 96152 1224 96228 1670
rect 97784 1224 97860 1670
rect 98464 0 98540 13094
rect 98872 12006 98948 13540
rect 99008 13230 99084 15172
rect 101320 13600 101396 14318
rect 99008 12550 99084 13132
rect 98736 11016 98812 11870
rect 99008 11696 99084 12278
rect 99552 1224 99628 1670
rect 100912 0 100988 13094
rect 101320 12006 101396 13540
rect 101456 13230 101532 15172
rect 101592 15134 101668 17076
rect 103496 13638 103572 14356
rect 101456 12550 101532 13132
rect 101184 11016 101260 11870
rect 101456 11696 101532 12278
rect 101320 1224 101396 1670
rect 102816 1224 102892 1670
rect 103360 0 103436 13094
rect 103632 12006 103708 13676
rect 103768 13600 103844 14318
rect 103768 12550 103844 13132
rect 103904 13094 103980 15172
rect 104040 15134 104116 17076
rect 106352 15134 106428 17076
rect 122808 17038 122884 19796
rect 106352 13600 106428 14318
rect 103632 11016 103708 11870
rect 103768 11696 103844 12278
rect 104584 1224 104660 1670
rect 105944 0 106020 13094
rect 106080 11696 106156 12278
rect 106352 12006 106428 13540
rect 106488 13230 106564 15172
rect 122808 14280 122884 16902
rect 122944 15640 123020 18398
rect 106488 12550 106564 13132
rect 106216 11016 106292 11870
rect 122808 11462 122884 14084
rect 122944 12822 123020 15580
rect 108256 10608 108332 11054
rect 108392 9520 108468 11326
rect 122944 9928 123020 12686
rect 106216 1224 106292 1670
rect 107848 1224 107924 1670
rect 109752 1224 109828 1670
rect 111248 1224 111324 1670
rect 113016 1224 113092 1670
rect 114784 1224 114860 1670
rect 116280 1224 116356 1670
rect 118048 1224 118124 1670
rect 119816 1224 119892 1670
rect 121312 1224 121388 1670
rect 123080 1224 123156 1670
rect 123216 0 123292 11870
rect 123352 0 123428 10782
rect 124712 1224 124788 1670
rect 126344 1224 126420 1670
rect 127976 1224 128052 1670
rect 129744 1224 129820 1670
rect 131512 1224 131588 1670
rect 133144 1224 133220 1670
rect 135320 952 135668 82356
rect 136000 272 136348 83036
use sky130_sram_2kbyte_1rw1r_32x512_8_col_addr_dff  sky130_sram_2kbyte_1rw1r_32x512_8_col_addr_dff_1
timestamp 1626065694
transform -1 0 119964 0 -1 80801
box -36 -49 2372 1467
use sky130_sram_2kbyte_1rw1r_32x512_8_col_addr_dff  sky130_sram_2kbyte_1rw1r_32x512_8_col_addr_dff_0
timestamp 1626065694
transform 1 0 15862 0 1 2396
box -36 -49 2372 1467
use sky130_sram_2kbyte_1rw1r_32x512_8_data_dff  sky130_sram_2kbyte_1rw1r_32x512_8_data_dff_0
timestamp 1626065694
transform 1 0 22870 0 1 2396
box -36 -49 37412 1467
use sky130_sram_2kbyte_1rw1r_32x512_8_row_addr_dff  sky130_sram_2kbyte_1rw1r_32x512_8_row_addr_dff_1
timestamp 1626065694
transform 1 0 13526 0 1 27746
box -36 -49 1204 9951
use sky130_sram_2kbyte_1rw1r_32x512_8_row_addr_dff  sky130_sram_2kbyte_1rw1r_32x512_8_row_addr_dff_0
timestamp 1626065694
transform -1 0 123468 0 -1 19846
box -36 -49 1204 9951
use sky130_sram_2kbyte_1rw1r_32x512_8_wmask_dff  sky130_sram_2kbyte_1rw1r_32x512_8_wmask_dff_0
timestamp 1626065694
transform 1 0 18198 0 1 2396
box -36 -49 4708 1467
use sky130_sram_2kbyte_1rw1r_32x512_8_control_logic_r  sky130_sram_2kbyte_1rw1r_32x512_8_control_logic_r_0
timestamp 1626065694
transform -1 0 134082 0 -1 79804
box -75 -49 11782 18431
use sky130_sram_2kbyte_1rw1r_32x512_8_control_logic_rw  sky130_sram_2kbyte_1rw1r_32x512_8_control_logic_rw_0
timestamp 1626065694
transform 1 0 2612 0 1 7620
box -75 -49 12082 18431
use sky130_sram_2kbyte_1rw1r_32x512_8_cr_3  sky130_sram_2kbyte_1rw1r_32x512_8_cr_3_0
timestamp 1626065694
transform 1 0 14862 0 1 9422
box 2083 -6379 5297 4372
use sky130_sram_2kbyte_1rw1r_32x512_8_cr_5  sky130_sram_2kbyte_1rw1r_32x512_8_cr_5_0
timestamp 1626065694
transform 1 0 14862 0 1 9422
box 101765 67036 104019 70732
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_3
timestamp 1626065694
transform 1 0 122183 0 1 80456
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_2
timestamp 1626065694
transform 1 0 14745 0 1 28017
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_1
timestamp 1626065694
transform 1 0 14745 0 1 2667
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_32  sky130_sram_2kbyte_1rw1r_32x512_8_contact_32_0
timestamp 1626065694
transform 1 0 122183 0 1 19501
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_71
timestamp 1626065694
transform 1 0 135592 0 1 82149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_70
timestamp 1626065694
transform 1 0 135456 0 1 82149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_69
timestamp 1626065694
transform 1 0 135320 0 1 82285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_68
timestamp 1626065694
transform 1 0 135320 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_67
timestamp 1626065694
transform 1 0 135592 0 1 82285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_66
timestamp 1626065694
transform 1 0 135456 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_65
timestamp 1626065694
transform 1 0 135320 0 1 82149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_64
timestamp 1626065694
transform 1 0 135592 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_63
timestamp 1626065694
transform 1 0 135456 0 1 82285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_62
timestamp 1626065694
transform 1 0 136136 0 1 82693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_61
timestamp 1626065694
transform 1 0 136136 0 1 82965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_60
timestamp 1626065694
transform 1 0 136272 0 1 82829
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_59
timestamp 1626065694
transform 1 0 136272 0 1 82693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_58
timestamp 1626065694
transform 1 0 136000 0 1 82965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_57
timestamp 1626065694
transform 1 0 136136 0 1 82829
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_56
timestamp 1626065694
transform 1 0 136272 0 1 82965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_55
timestamp 1626065694
transform 1 0 136000 0 1 82693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_54
timestamp 1626065694
transform 1 0 136000 0 1 82829
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_53
timestamp 1626065694
transform 1 0 1088 0 1 82149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_52
timestamp 1626065694
transform 1 0 272 0 1 82693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_51
timestamp 1626065694
transform 1 0 952 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_50
timestamp 1626065694
transform 1 0 1088 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_49
timestamp 1626065694
transform 1 0 408 0 1 82965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_48
timestamp 1626065694
transform 1 0 544 0 1 82693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_47
timestamp 1626065694
transform 1 0 408 0 1 82693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_46
timestamp 1626065694
transform 1 0 1224 0 1 82285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_45
timestamp 1626065694
transform 1 0 544 0 1 82965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_44
timestamp 1626065694
transform 1 0 272 0 1 82965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_43
timestamp 1626065694
transform 1 0 952 0 1 82285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_42
timestamp 1626065694
transform 1 0 952 0 1 82149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_41
timestamp 1626065694
transform 1 0 1224 0 1 82149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_40
timestamp 1626065694
transform 1 0 1088 0 1 82285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_39
timestamp 1626065694
transform 1 0 544 0 1 82829
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_38
timestamp 1626065694
transform 1 0 272 0 1 82829
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_37
timestamp 1626065694
transform 1 0 1224 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_36
timestamp 1626065694
transform 1 0 408 0 1 82829
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_35
timestamp 1626065694
transform 1 0 272 0 1 549
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_34
timestamp 1626065694
transform 1 0 272 0 1 413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_33
timestamp 1626065694
transform 1 0 952 0 1 957
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_32
timestamp 1626065694
transform 1 0 1224 0 1 957
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_31
timestamp 1626065694
transform 1 0 544 0 1 413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_30
timestamp 1626065694
transform 1 0 1224 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_29
timestamp 1626065694
transform 1 0 1088 0 1 957
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_28
timestamp 1626065694
transform 1 0 272 0 1 277
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_27
timestamp 1626065694
transform 1 0 408 0 1 549
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_26
timestamp 1626065694
transform 1 0 1088 0 1 1093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_25
timestamp 1626065694
transform 1 0 1088 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_24
timestamp 1626065694
transform 1 0 952 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_23
timestamp 1626065694
transform 1 0 952 0 1 1093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_22
timestamp 1626065694
transform 1 0 1224 0 1 1093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_21
timestamp 1626065694
transform 1 0 544 0 1 549
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_20
timestamp 1626065694
transform 1 0 408 0 1 413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_19
timestamp 1626065694
transform 1 0 544 0 1 277
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_18
timestamp 1626065694
transform 1 0 408 0 1 277
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_17
timestamp 1626065694
transform 1 0 136136 0 1 413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_16
timestamp 1626065694
transform 1 0 136136 0 1 277
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_15
timestamp 1626065694
transform 1 0 135320 0 1 1093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_14
timestamp 1626065694
transform 1 0 135592 0 1 957
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_13
timestamp 1626065694
transform 1 0 136000 0 1 549
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_12
timestamp 1626065694
transform 1 0 135456 0 1 1093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_11
timestamp 1626065694
transform 1 0 136272 0 1 549
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_10
timestamp 1626065694
transform 1 0 136000 0 1 277
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_9
timestamp 1626065694
transform 1 0 136272 0 1 277
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_8
timestamp 1626065694
transform 1 0 135456 0 1 957
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_7
timestamp 1626065694
transform 1 0 135320 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_6
timestamp 1626065694
transform 1 0 135592 0 1 1093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_5
timestamp 1626065694
transform 1 0 135456 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_4
timestamp 1626065694
transform 1 0 135320 0 1 957
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_3
timestamp 1626065694
transform 1 0 135592 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_2
timestamp 1626065694
transform 1 0 136136 0 1 549
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_1
timestamp 1626065694
transform 1 0 136272 0 1 413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_39  sky130_sram_2kbyte_1rw1r_32x512_8_contact_39_0
timestamp 1626065694
transform 1 0 136000 0 1 413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_38  sky130_sram_2kbyte_1rw1r_32x512_8_contact_38_3
timestamp 1626065694
transform 1 0 134776 0 1 81377
box 0 0 192 192
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_38  sky130_sram_2kbyte_1rw1r_32x512_8_contact_38_2
timestamp 1626065694
transform 1 0 1726 0 1 81377
box 0 0 192 192
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_38  sky130_sram_2kbyte_1rw1r_32x512_8_contact_38_1
timestamp 1626065694
transform 1 0 1726 0 1 1628
box 0 0 192 192
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_38  sky130_sram_2kbyte_1rw1r_32x512_8_contact_38_0
timestamp 1626065694
transform 1 0 134776 0 1 1628
box 0 0 192 192
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_420
timestamp 1626065694
transform 1 0 133165 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_419
timestamp 1626065694
transform 1 0 134839 0 1 80983
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_418
timestamp 1626065694
transform 1 0 129805 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_417
timestamp 1626065694
transform 1 0 131485 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_416
timestamp 1626065694
transform 1 0 128125 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_415
timestamp 1626065694
transform 1 0 130742 0 1 79098
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_414
timestamp 1626065694
transform 1 0 134839 0 1 79303
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_413
timestamp 1626065694
transform 1 0 133879 0 1 79203
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_412
timestamp 1626065694
transform 1 0 126445 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_411
timestamp 1626065694
transform 1 0 119761 0 1 80200
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_410
timestamp 1626065694
transform 1 0 119725 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_409
timestamp 1626065694
transform 1 0 121405 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_408
timestamp 1626065694
transform 1 0 123085 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_407
timestamp 1626065694
transform 1 0 124765 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_406
timestamp 1626065694
transform 1 0 122267 0 1 73404
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_405
timestamp 1626065694
transform 1 0 122267 0 1 74818
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_404
timestamp 1626065694
transform 1 0 134839 0 1 77623
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_403
timestamp 1626065694
transform 1 0 134839 0 1 74263
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_402
timestamp 1626065694
transform 1 0 134839 0 1 75943
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_401
timestamp 1626065694
transform 1 0 111325 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_400
timestamp 1626065694
transform 1 0 113005 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_399
timestamp 1626065694
transform 1 0 114685 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_398
timestamp 1626065694
transform 1 0 116365 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_397
timestamp 1626065694
transform 1 0 118045 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_396
timestamp 1626065694
transform 1 0 118593 0 1 80200
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_395
timestamp 1626065694
transform 1 0 106285 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_394
timestamp 1626065694
transform 1 0 107965 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_393
timestamp 1626065694
transform 1 0 109645 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_392
timestamp 1626065694
transform 1 0 102925 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_391
timestamp 1626065694
transform 1 0 104605 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_390
timestamp 1626065694
transform 1 0 110180 0 1 73404
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_389
timestamp 1626065694
transform 1 0 110056 0 1 74818
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_388
timestamp 1626065694
transform 1 0 103493 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_387
timestamp 1626065694
transform 1 0 105989 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_386
timestamp 1626065694
transform 1 0 114041 0 1 71990
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_385
timestamp 1626065694
transform 1 0 134839 0 1 69223
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_384
timestamp 1626065694
transform 1 0 134839 0 1 70903
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_383
timestamp 1626065694
transform 1 0 134839 0 1 72583
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_382
timestamp 1626065694
transform 1 0 134839 0 1 67543
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_381
timestamp 1626065694
transform 1 0 122267 0 1 71990
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_380
timestamp 1626065694
transform 1 0 134839 0 1 64183
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_379
timestamp 1626065694
transform 1 0 134839 0 1 65863
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_378
timestamp 1626065694
transform 1 0 134839 0 1 62503
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_377
timestamp 1626065694
transform 1 0 94525 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_376
timestamp 1626065694
transform 1 0 96205 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_375
timestamp 1626065694
transform 1 0 97885 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_374
timestamp 1626065694
transform 1 0 99565 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_373
timestamp 1626065694
transform 1 0 101245 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_372
timestamp 1626065694
transform 1 0 87805 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_371
timestamp 1626065694
transform 1 0 89485 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_370
timestamp 1626065694
transform 1 0 91165 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_369
timestamp 1626065694
transform 1 0 92845 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_368
timestamp 1626065694
transform 1 0 86125 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_367
timestamp 1626065694
transform 1 0 86021 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_366
timestamp 1626065694
transform 1 0 88517 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_365
timestamp 1626065694
transform 1 0 91013 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_364
timestamp 1626065694
transform 1 0 93509 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_363
timestamp 1626065694
transform 1 0 98501 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_362
timestamp 1626065694
transform 1 0 100997 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_361
timestamp 1626065694
transform 1 0 96005 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_360
timestamp 1626065694
transform 1 0 77725 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_359
timestamp 1626065694
transform 1 0 79405 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_358
timestamp 1626065694
transform 1 0 81085 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_357
timestamp 1626065694
transform 1 0 82765 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_356
timestamp 1626065694
transform 1 0 84445 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_355
timestamp 1626065694
transform 1 0 69325 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_354
timestamp 1626065694
transform 1 0 71005 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_353
timestamp 1626065694
transform 1 0 72685 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_352
timestamp 1626065694
transform 1 0 74365 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_351
timestamp 1626065694
transform 1 0 76045 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_350
timestamp 1626065694
transform 1 0 73541 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_349
timestamp 1626065694
transform 1 0 76037 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_348
timestamp 1626065694
transform 1 0 68549 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_347
timestamp 1626065694
transform 1 0 71045 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_346
timestamp 1626065694
transform 1 0 81029 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_345
timestamp 1626065694
transform 1 0 83525 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_344
timestamp 1626065694
transform 1 0 78533 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_343
timestamp 1626065694
transform 1 0 134839 0 1 57463
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_342
timestamp 1626065694
transform 1 0 134839 0 1 59143
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_341
timestamp 1626065694
transform 1 0 134839 0 1 60823
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_340
timestamp 1626065694
transform 1 0 134092 0 1 62054
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_339
timestamp 1626065694
transform 1 0 134839 0 1 52423
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_338
timestamp 1626065694
transform 1 0 134839 0 1 54103
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_337
timestamp 1626065694
transform 1 0 134839 0 1 55783
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_336
timestamp 1626065694
transform 1 0 134839 0 1 50743
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_335
timestamp 1626065694
transform 1 0 134839 0 1 49063
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_334
timestamp 1626065694
transform 1 0 134839 0 1 47383
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_333
timestamp 1626065694
transform 1 0 134839 0 1 44023
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_332
timestamp 1626065694
transform 1 0 134839 0 1 45703
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_331
timestamp 1626065694
transform 1 0 134839 0 1 42343
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_330
timestamp 1626065694
transform 1 0 60925 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_329
timestamp 1626065694
transform 1 0 62605 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_328
timestamp 1626065694
transform 1 0 64285 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_327
timestamp 1626065694
transform 1 0 65965 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_326
timestamp 1626065694
transform 1 0 67645 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_325
timestamp 1626065694
transform 1 0 59245 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_324
timestamp 1626065694
transform 1 0 52525 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_323
timestamp 1626065694
transform 1 0 54205 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_322
timestamp 1626065694
transform 1 0 55885 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_321
timestamp 1626065694
transform 1 0 57565 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_320
timestamp 1626065694
transform 1 0 53573 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_319
timestamp 1626065694
transform 1 0 56069 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_318
timestamp 1626065694
transform 1 0 58565 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_317
timestamp 1626065694
transform 1 0 61061 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_316
timestamp 1626065694
transform 1 0 63557 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_315
timestamp 1626065694
transform 1 0 66053 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_314
timestamp 1626065694
transform 1 0 47485 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_313
timestamp 1626065694
transform 1 0 49165 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_312
timestamp 1626065694
transform 1 0 50845 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_311
timestamp 1626065694
transform 1 0 44125 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_310
timestamp 1626065694
transform 1 0 45805 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_309
timestamp 1626065694
transform 1 0 37405 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_308
timestamp 1626065694
transform 1 0 39085 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_307
timestamp 1626065694
transform 1 0 40765 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_306
timestamp 1626065694
transform 1 0 42445 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_305
timestamp 1626065694
transform 1 0 35725 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_304
timestamp 1626065694
transform 1 0 36101 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_303
timestamp 1626065694
transform 1 0 38597 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_302
timestamp 1626065694
transform 1 0 41093 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_301
timestamp 1626065694
transform 1 0 43589 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_300
timestamp 1626065694
transform 1 0 46085 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_299
timestamp 1626065694
transform 1 0 48581 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_298
timestamp 1626065694
transform 1 0 51077 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_297
timestamp 1626065694
transform 1 0 17245 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_296
timestamp 1626065694
transform 1 0 27325 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_295
timestamp 1626065694
transform 1 0 29005 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_294
timestamp 1626065694
transform 1 0 30685 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_293
timestamp 1626065694
transform 1 0 32365 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_292
timestamp 1626065694
transform 1 0 34045 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_291
timestamp 1626065694
transform 1 0 25645 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_290
timestamp 1626065694
transform 1 0 18925 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_289
timestamp 1626065694
transform 1 0 20605 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_288
timestamp 1626065694
transform 1 0 22285 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_287
timestamp 1626065694
transform 1 0 23965 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_286
timestamp 1626065694
transform 1 0 33605 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_285
timestamp 1626065694
transform 1 0 28613 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_284
timestamp 1626065694
transform 1 0 31109 0 1 76982
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_283
timestamp 1626065694
transform 1 0 8845 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_282
timestamp 1626065694
transform 1 0 10525 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_281
timestamp 1626065694
transform 1 0 12205 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_280
timestamp 1626065694
transform 1 0 13885 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_279
timestamp 1626065694
transform 1 0 15565 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_278
timestamp 1626065694
transform 1 0 5485 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_277
timestamp 1626065694
transform 1 0 7165 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_276
timestamp 1626065694
transform 1 0 3805 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_275
timestamp 1626065694
transform 1 0 1789 0 1 80983
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_274
timestamp 1626065694
transform 1 0 2125 0 1 81436
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_273
timestamp 1626065694
transform 1 0 1789 0 1 79303
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_272
timestamp 1626065694
transform 1 0 1789 0 1 74263
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_271
timestamp 1626065694
transform 1 0 1789 0 1 75943
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_270
timestamp 1626065694
transform 1 0 1789 0 1 77623
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_269
timestamp 1626065694
transform 1 0 1789 0 1 70903
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_268
timestamp 1626065694
transform 1 0 1789 0 1 72583
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_267
timestamp 1626065694
transform 1 0 1789 0 1 69223
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_266
timestamp 1626065694
transform 1 0 1789 0 1 67543
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_265
timestamp 1626065694
transform 1 0 1789 0 1 64183
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_264
timestamp 1626065694
transform 1 0 1789 0 1 65863
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_263
timestamp 1626065694
transform 1 0 1789 0 1 62503
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_262
timestamp 1626065694
transform 1 0 1789 0 1 57463
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_261
timestamp 1626065694
transform 1 0 1789 0 1 59143
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_260
timestamp 1626065694
transform 1 0 1789 0 1 60823
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_259
timestamp 1626065694
transform 1 0 1789 0 1 54103
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_258
timestamp 1626065694
transform 1 0 1789 0 1 55783
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_257
timestamp 1626065694
transform 1 0 1789 0 1 52423
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_256
timestamp 1626065694
transform 1 0 1789 0 1 50743
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_255
timestamp 1626065694
transform 1 0 1789 0 1 49063
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_254
timestamp 1626065694
transform 1 0 1789 0 1 47383
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_253
timestamp 1626065694
transform 1 0 1789 0 1 42343
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_252
timestamp 1626065694
transform 1 0 1789 0 1 44023
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_251
timestamp 1626065694
transform 1 0 1789 0 1 45703
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_250
timestamp 1626065694
transform 1 0 13663 0 1 36757
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_249
timestamp 1626065694
transform 1 0 14608 0 1 36828
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_248
timestamp 1626065694
transform 1 0 15342 0 1 36828
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_247
timestamp 1626065694
transform 1 0 1789 0 1 37303
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_246
timestamp 1626065694
transform 1 0 1789 0 1 38983
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_245
timestamp 1626065694
transform 1 0 1789 0 1 40663
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_244
timestamp 1626065694
transform 1 0 1789 0 1 33943
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_243
timestamp 1626065694
transform 1 0 1789 0 1 35623
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_242
timestamp 1626065694
transform 1 0 1789 0 1 32263
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_241
timestamp 1626065694
transform 1 0 13663 0 1 32801
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_240
timestamp 1626065694
transform 1 0 13663 0 1 33929
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_239
timestamp 1626065694
transform 1 0 15102 0 1 32730
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_238
timestamp 1626065694
transform 1 0 14608 0 1 34000
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_237
timestamp 1626065694
transform 1 0 15262 0 1 35558
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_236
timestamp 1626065694
transform 1 0 15182 0 1 34000
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_235
timestamp 1626065694
transform 1 0 14608 0 1 32730
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_234
timestamp 1626065694
transform 1 0 14608 0 1 35558
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_233
timestamp 1626065694
transform 1 0 13663 0 1 35629
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_232
timestamp 1626065694
transform 1 0 14942 0 1 29902
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_231
timestamp 1626065694
transform 1 0 14608 0 1 31172
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_230
timestamp 1626065694
transform 1 0 15022 0 1 31172
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_229
timestamp 1626065694
transform 1 0 14608 0 1 28344
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_228
timestamp 1626065694
transform 1 0 13663 0 1 28273
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_227
timestamp 1626065694
transform 1 0 13663 0 1 29973
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_226
timestamp 1626065694
transform 1 0 14862 0 1 28344
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_225
timestamp 1626065694
transform 1 0 14608 0 1 29902
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_224
timestamp 1626065694
transform 1 0 13663 0 1 31101
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_223
timestamp 1626065694
transform 1 0 1789 0 1 30583
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_222
timestamp 1626065694
transform 1 0 1789 0 1 27223
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_221
timestamp 1626065694
transform 1 0 1789 0 1 28903
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_220
timestamp 1626065694
transform 1 0 1789 0 1 23863
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_219
timestamp 1626065694
transform 1 0 1789 0 1 25543
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_218
timestamp 1626065694
transform 1 0 2536 0 1 25296
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_217
timestamp 1626065694
transform 1 0 1789 0 1 22183
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_216
timestamp 1626065694
transform 1 0 17245 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_215
timestamp 1626065694
transform 1 0 22803 0 1 18188
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_214
timestamp 1626065694
transform 1 0 33605 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_213
timestamp 1626065694
transform 1 0 26506 0 1 15360
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_212
timestamp 1626065694
transform 1 0 26630 0 1 12532
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_211
timestamp 1626065694
transform 1 0 26754 0 1 13946
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_210
timestamp 1626065694
transform 1 0 28613 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_209
timestamp 1626065694
transform 1 0 31109 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_208
timestamp 1626065694
transform 1 0 14661 0 1 18188
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_207
timestamp 1626065694
transform 1 0 1789 0 1 17143
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_206
timestamp 1626065694
transform 1 0 1789 0 1 18823
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_205
timestamp 1626065694
transform 1 0 1789 0 1 20503
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_204
timestamp 1626065694
transform 1 0 1789 0 1 13783
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_203
timestamp 1626065694
transform 1 0 1789 0 1 12103
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_202
timestamp 1626065694
transform 1 0 1789 0 1 15463
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_201
timestamp 1626065694
transform 1 0 14661 0 1 12532
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_200
timestamp 1626065694
transform 1 0 14661 0 1 13946
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_199
timestamp 1626065694
transform 1 0 14661 0 1 15360
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_198
timestamp 1626065694
transform 1 0 1789 0 1 5383
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_197
timestamp 1626065694
transform 1 0 1789 0 1 7063
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_196
timestamp 1626065694
transform 1 0 1789 0 1 8743
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_195
timestamp 1626065694
transform 1 0 2749 0 1 8147
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_194
timestamp 1626065694
transform 1 0 2749 0 1 9847
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_193
timestamp 1626065694
transform 1 0 5970 0 1 8252
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_192
timestamp 1626065694
transform 1 0 1789 0 1 10423
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_191
timestamp 1626065694
transform 1 0 1789 0 1 3703
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_190
timestamp 1626065694
transform 1 0 1789 0 1 2023
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_189
timestamp 1626065694
transform 1 0 2125 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_188
timestamp 1626065694
transform 1 0 3805 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_187
timestamp 1626065694
transform 1 0 7165 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_186
timestamp 1626065694
transform 1 0 5485 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_185
timestamp 1626065694
transform 1 0 13885 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_184
timestamp 1626065694
transform 1 0 15565 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_183
timestamp 1626065694
transform 1 0 10525 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_182
timestamp 1626065694
transform 1 0 15999 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_181
timestamp 1626065694
transform 1 0 17167 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_180
timestamp 1626065694
transform 1 0 12205 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_179
timestamp 1626065694
transform 1 0 8845 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_178
timestamp 1626065694
transform 1 0 18335 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_177
timestamp 1626065694
transform 1 0 19503 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_176
timestamp 1626065694
transform 1 0 20671 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_175
timestamp 1626065694
transform 1 0 21839 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_174
timestamp 1626065694
transform 1 0 18925 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_173
timestamp 1626065694
transform 1 0 22285 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_172
timestamp 1626065694
transform 1 0 23965 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_171
timestamp 1626065694
transform 1 0 25645 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_170
timestamp 1626065694
transform 1 0 23007 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_169
timestamp 1626065694
transform 1 0 24175 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_168
timestamp 1626065694
transform 1 0 25343 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_167
timestamp 1626065694
transform 1 0 20605 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_166
timestamp 1626065694
transform 1 0 29005 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_165
timestamp 1626065694
transform 1 0 34045 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_164
timestamp 1626065694
transform 1 0 30685 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_163
timestamp 1626065694
transform 1 0 26511 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_162
timestamp 1626065694
transform 1 0 27679 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_161
timestamp 1626065694
transform 1 0 28847 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_160
timestamp 1626065694
transform 1 0 30015 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_159
timestamp 1626065694
transform 1 0 31183 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_158
timestamp 1626065694
transform 1 0 32351 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_157
timestamp 1626065694
transform 1 0 33519 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_156
timestamp 1626065694
transform 1 0 32365 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_155
timestamp 1626065694
transform 1 0 27325 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_154
timestamp 1626065694
transform 1 0 53573 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_153
timestamp 1626065694
transform 1 0 56069 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_152
timestamp 1626065694
transform 1 0 58565 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_151
timestamp 1626065694
transform 1 0 61061 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_150
timestamp 1626065694
transform 1 0 63557 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_149
timestamp 1626065694
transform 1 0 66053 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_148
timestamp 1626065694
transform 1 0 36101 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_147
timestamp 1626065694
transform 1 0 38597 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_146
timestamp 1626065694
transform 1 0 41093 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_145
timestamp 1626065694
transform 1 0 43589 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_144
timestamp 1626065694
transform 1 0 46085 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_143
timestamp 1626065694
transform 1 0 48581 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_142
timestamp 1626065694
transform 1 0 51077 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_141
timestamp 1626065694
transform 1 0 37023 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_140
timestamp 1626065694
transform 1 0 40765 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_139
timestamp 1626065694
transform 1 0 42445 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_138
timestamp 1626065694
transform 1 0 38191 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_137
timestamp 1626065694
transform 1 0 34687 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_136
timestamp 1626065694
transform 1 0 39359 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_135
timestamp 1626065694
transform 1 0 40527 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_134
timestamp 1626065694
transform 1 0 41695 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_133
timestamp 1626065694
transform 1 0 35855 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_132
timestamp 1626065694
transform 1 0 35725 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_131
timestamp 1626065694
transform 1 0 37405 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_130
timestamp 1626065694
transform 1 0 39085 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_129
timestamp 1626065694
transform 1 0 44125 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_128
timestamp 1626065694
transform 1 0 44031 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_127
timestamp 1626065694
transform 1 0 49165 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_126
timestamp 1626065694
transform 1 0 45199 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_125
timestamp 1626065694
transform 1 0 42863 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_124
timestamp 1626065694
transform 1 0 50845 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_123
timestamp 1626065694
transform 1 0 51039 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_122
timestamp 1626065694
transform 1 0 46367 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_121
timestamp 1626065694
transform 1 0 47535 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_120
timestamp 1626065694
transform 1 0 45805 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_119
timestamp 1626065694
transform 1 0 48703 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_118
timestamp 1626065694
transform 1 0 49871 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_117
timestamp 1626065694
transform 1 0 47485 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_116
timestamp 1626065694
transform 1 0 53375 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_115
timestamp 1626065694
transform 1 0 54543 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_114
timestamp 1626065694
transform 1 0 55711 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_113
timestamp 1626065694
transform 1 0 56879 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_112
timestamp 1626065694
transform 1 0 58047 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_111
timestamp 1626065694
transform 1 0 59215 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_110
timestamp 1626065694
transform 1 0 52525 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_109
timestamp 1626065694
transform 1 0 54205 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_108
timestamp 1626065694
transform 1 0 52207 0 1 2923
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_107
timestamp 1626065694
transform 1 0 57565 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_106
timestamp 1626065694
transform 1 0 55885 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_105
timestamp 1626065694
transform 1 0 59245 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_104
timestamp 1626065694
transform 1 0 67645 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_103
timestamp 1626065694
transform 1 0 62605 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_102
timestamp 1626065694
transform 1 0 64285 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_101
timestamp 1626065694
transform 1 0 60925 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_100
timestamp 1626065694
transform 1 0 65965 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_99
timestamp 1626065694
transform 1 0 134839 0 1 37303
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_98
timestamp 1626065694
transform 1 0 134839 0 1 38983
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_97
timestamp 1626065694
transform 1 0 134839 0 1 40663
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_96
timestamp 1626065694
transform 1 0 134839 0 1 32263
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_95
timestamp 1626065694
transform 1 0 134839 0 1 33943
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_94
timestamp 1626065694
transform 1 0 134839 0 1 35623
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_93
timestamp 1626065694
transform 1 0 134839 0 1 28903
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_92
timestamp 1626065694
transform 1 0 134839 0 1 30583
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_91
timestamp 1626065694
transform 1 0 134839 0 1 27223
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_90
timestamp 1626065694
transform 1 0 134839 0 1 25543
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_89
timestamp 1626065694
transform 1 0 134839 0 1 22183
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_88
timestamp 1626065694
transform 1 0 134839 0 1 23863
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_87
timestamp 1626065694
transform 1 0 86021 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_86
timestamp 1626065694
transform 1 0 88517 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_85
timestamp 1626065694
transform 1 0 91013 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_84
timestamp 1626065694
transform 1 0 93509 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_83
timestamp 1626065694
transform 1 0 96005 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_82
timestamp 1626065694
transform 1 0 98501 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_81
timestamp 1626065694
transform 1 0 100997 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_80
timestamp 1626065694
transform 1 0 68549 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_79
timestamp 1626065694
transform 1 0 71045 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_78
timestamp 1626065694
transform 1 0 73541 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_77
timestamp 1626065694
transform 1 0 76037 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_76
timestamp 1626065694
transform 1 0 78533 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_75
timestamp 1626065694
transform 1 0 81029 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_74
timestamp 1626065694
transform 1 0 83525 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_73
timestamp 1626065694
transform 1 0 69325 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_72
timestamp 1626065694
transform 1 0 71005 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_71
timestamp 1626065694
transform 1 0 72685 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_70
timestamp 1626065694
transform 1 0 76045 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_69
timestamp 1626065694
transform 1 0 74365 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_68
timestamp 1626065694
transform 1 0 79405 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_67
timestamp 1626065694
transform 1 0 82765 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_66
timestamp 1626065694
transform 1 0 81085 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_65
timestamp 1626065694
transform 1 0 84445 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_64
timestamp 1626065694
transform 1 0 77725 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_63
timestamp 1626065694
transform 1 0 92845 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_62
timestamp 1626065694
transform 1 0 87805 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_61
timestamp 1626065694
transform 1 0 91165 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_60
timestamp 1626065694
transform 1 0 89485 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_59
timestamp 1626065694
transform 1 0 86125 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_58
timestamp 1626065694
transform 1 0 99565 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_57
timestamp 1626065694
transform 1 0 97885 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_56
timestamp 1626065694
transform 1 0 101245 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_55
timestamp 1626065694
transform 1 0 96205 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_54
timestamp 1626065694
transform 1 0 94525 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_53
timestamp 1626065694
transform 1 0 134839 0 1 17143
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_52
timestamp 1626065694
transform 1 0 134839 0 1 18823
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_51
timestamp 1626065694
transform 1 0 134839 0 1 20503
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_50
timestamp 1626065694
transform 1 0 123265 0 1 19245
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_49
timestamp 1626065694
transform 1 0 123265 0 1 17545
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_48
timestamp 1626065694
transform 1 0 123265 0 1 16417
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_47
timestamp 1626065694
transform 1 0 122320 0 1 19174
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_46
timestamp 1626065694
transform 1 0 121982 0 1 19174
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_45
timestamp 1626065694
transform 1 0 122320 0 1 17616
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_44
timestamp 1626065694
transform 1 0 121902 0 1 17616
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_43
timestamp 1626065694
transform 1 0 122320 0 1 16346
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_42
timestamp 1626065694
transform 1 0 121822 0 1 16346
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_41
timestamp 1626065694
transform 1 0 122320 0 1 11960
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_40
timestamp 1626065694
transform 1 0 121582 0 1 11960
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_39
timestamp 1626065694
transform 1 0 122320 0 1 10690
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_38
timestamp 1626065694
transform 1 0 121502 0 1 10690
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_37
timestamp 1626065694
transform 1 0 121742 0 1 14788
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_36
timestamp 1626065694
transform 1 0 122320 0 1 13518
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_35
timestamp 1626065694
transform 1 0 121662 0 1 13518
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_34
timestamp 1626065694
transform 1 0 123265 0 1 14717
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_33
timestamp 1626065694
transform 1 0 123265 0 1 13589
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_32
timestamp 1626065694
transform 1 0 123265 0 1 11889
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_31
timestamp 1626065694
transform 1 0 123265 0 1 10761
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_30
timestamp 1626065694
transform 1 0 122320 0 1 14788
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_29
timestamp 1626065694
transform 1 0 134839 0 1 15463
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_28
timestamp 1626065694
transform 1 0 134839 0 1 12103
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_27
timestamp 1626065694
transform 1 0 134839 0 1 13783
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_26
timestamp 1626065694
transform 1 0 103493 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_25
timestamp 1626065694
transform 1 0 105989 0 1 13196
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_24
timestamp 1626065694
transform 1 0 109645 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_23
timestamp 1626065694
transform 1 0 106285 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_22
timestamp 1626065694
transform 1 0 104605 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_21
timestamp 1626065694
transform 1 0 107965 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_20
timestamp 1626065694
transform 1 0 102925 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_19
timestamp 1626065694
transform 1 0 116365 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_18
timestamp 1626065694
transform 1 0 118045 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_17
timestamp 1626065694
transform 1 0 113005 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_16
timestamp 1626065694
transform 1 0 111325 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_15
timestamp 1626065694
transform 1 0 114685 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_14
timestamp 1626065694
transform 1 0 134839 0 1 5383
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_13
timestamp 1626065694
transform 1 0 134839 0 1 7063
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_12
timestamp 1626065694
transform 1 0 134839 0 1 8743
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_11
timestamp 1626065694
transform 1 0 134839 0 1 10423
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_10
timestamp 1626065694
transform 1 0 126445 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_9
timestamp 1626065694
transform 1 0 119725 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_8
timestamp 1626065694
transform 1 0 121405 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_7
timestamp 1626065694
transform 1 0 123085 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_6
timestamp 1626065694
transform 1 0 124765 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_5
timestamp 1626065694
transform 1 0 134839 0 1 3703
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_4
timestamp 1626065694
transform 1 0 128125 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_3
timestamp 1626065694
transform 1 0 129805 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_2
timestamp 1626065694
transform 1 0 131485 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1626065694
transform 1 0 133165 0 1 1687
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1626065694
transform 1 0 134839 0 1 2023
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_cr_4  sky130_sram_2kbyte_1rw1r_32x512_8_cr_4_0
timestamp 1626065694
transform 1 0 14862 0 1 9422
box 4376 -6402 91393 1462
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_707
timestamp 1626065694
transform 1 0 133166 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_706
timestamp 1626065694
transform 1 0 134840 0 1 80652
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_705
timestamp 1626065694
transform 1 0 134840 0 1 80988
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_704
timestamp 1626065694
transform 1 0 131486 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_703
timestamp 1626065694
transform 1 0 128126 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_702
timestamp 1626065694
transform 1 0 129806 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_701
timestamp 1626065694
transform 1 0 134840 0 1 79308
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_700
timestamp 1626065694
transform 1 0 134840 0 1 79644
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_699
timestamp 1626065694
transform 1 0 134840 0 1 79980
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_698
timestamp 1626065694
transform 1 0 134840 0 1 80316
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_697
timestamp 1626065694
transform 1 0 134840 0 1 77964
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_696
timestamp 1626065694
transform 1 0 134840 0 1 78300
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_695
timestamp 1626065694
transform 1 0 134840 0 1 78636
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_694
timestamp 1626065694
transform 1 0 134840 0 1 78972
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_693
timestamp 1626065694
transform 1 0 119726 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_692
timestamp 1626065694
transform 1 0 121406 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_691
timestamp 1626065694
transform 1 0 123086 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_690
timestamp 1626065694
transform 1 0 124766 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_689
timestamp 1626065694
transform 1 0 126446 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_688
timestamp 1626065694
transform 1 0 134840 0 1 77292
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_687
timestamp 1626065694
transform 1 0 134840 0 1 77628
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_686
timestamp 1626065694
transform 1 0 134840 0 1 72924
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_685
timestamp 1626065694
transform 1 0 134840 0 1 73260
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_684
timestamp 1626065694
transform 1 0 134840 0 1 73596
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_683
timestamp 1626065694
transform 1 0 134840 0 1 73932
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_682
timestamp 1626065694
transform 1 0 134840 0 1 74268
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_681
timestamp 1626065694
transform 1 0 134840 0 1 74604
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_680
timestamp 1626065694
transform 1 0 134840 0 1 74940
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_679
timestamp 1626065694
transform 1 0 134840 0 1 75276
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_678
timestamp 1626065694
transform 1 0 134840 0 1 75612
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_677
timestamp 1626065694
transform 1 0 134840 0 1 75948
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_676
timestamp 1626065694
transform 1 0 134840 0 1 76284
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_675
timestamp 1626065694
transform 1 0 134840 0 1 76620
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_674
timestamp 1626065694
transform 1 0 134840 0 1 76956
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_673
timestamp 1626065694
transform 1 0 111326 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_672
timestamp 1626065694
transform 1 0 113006 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_671
timestamp 1626065694
transform 1 0 114686 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_670
timestamp 1626065694
transform 1 0 116366 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_669
timestamp 1626065694
transform 1 0 118046 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_668
timestamp 1626065694
transform 1 0 107966 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_667
timestamp 1626065694
transform 1 0 109646 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_666
timestamp 1626065694
transform 1 0 102926 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_665
timestamp 1626065694
transform 1 0 104606 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_664
timestamp 1626065694
transform 1 0 106286 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_663
timestamp 1626065694
transform 1 0 105990 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_662
timestamp 1626065694
transform 1 0 103494 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_661
timestamp 1626065694
transform 1 0 134840 0 1 68220
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_660
timestamp 1626065694
transform 1 0 134840 0 1 68556
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_659
timestamp 1626065694
transform 1 0 134840 0 1 68892
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_658
timestamp 1626065694
transform 1 0 134840 0 1 69228
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_657
timestamp 1626065694
transform 1 0 134840 0 1 69564
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_656
timestamp 1626065694
transform 1 0 134840 0 1 69900
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_655
timestamp 1626065694
transform 1 0 134840 0 1 70236
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_654
timestamp 1626065694
transform 1 0 134840 0 1 70572
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_653
timestamp 1626065694
transform 1 0 134840 0 1 70908
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_652
timestamp 1626065694
transform 1 0 134840 0 1 71244
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_651
timestamp 1626065694
transform 1 0 134840 0 1 71580
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_650
timestamp 1626065694
transform 1 0 134840 0 1 71916
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_649
timestamp 1626065694
transform 1 0 134840 0 1 72252
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_648
timestamp 1626065694
transform 1 0 134840 0 1 72588
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_647
timestamp 1626065694
transform 1 0 134840 0 1 67548
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_646
timestamp 1626065694
transform 1 0 134840 0 1 67884
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_645
timestamp 1626065694
transform 1 0 134840 0 1 63852
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_644
timestamp 1626065694
transform 1 0 134840 0 1 64188
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_643
timestamp 1626065694
transform 1 0 134840 0 1 64524
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_642
timestamp 1626065694
transform 1 0 134840 0 1 64860
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_641
timestamp 1626065694
transform 1 0 134840 0 1 65196
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_640
timestamp 1626065694
transform 1 0 134840 0 1 65532
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_639
timestamp 1626065694
transform 1 0 134840 0 1 65868
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_638
timestamp 1626065694
transform 1 0 134840 0 1 66204
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_637
timestamp 1626065694
transform 1 0 134840 0 1 66540
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_636
timestamp 1626065694
transform 1 0 134840 0 1 66876
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_635
timestamp 1626065694
transform 1 0 134840 0 1 67212
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_634
timestamp 1626065694
transform 1 0 134840 0 1 62508
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_633
timestamp 1626065694
transform 1 0 134840 0 1 62844
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_632
timestamp 1626065694
transform 1 0 134840 0 1 63180
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_631
timestamp 1626065694
transform 1 0 134840 0 1 63516
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_630
timestamp 1626065694
transform 1 0 94526 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_629
timestamp 1626065694
transform 1 0 96206 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_628
timestamp 1626065694
transform 1 0 97886 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_627
timestamp 1626065694
transform 1 0 99566 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_626
timestamp 1626065694
transform 1 0 101246 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_625
timestamp 1626065694
transform 1 0 87806 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_624
timestamp 1626065694
transform 1 0 89486 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_623
timestamp 1626065694
transform 1 0 91166 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_622
timestamp 1626065694
transform 1 0 92846 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_621
timestamp 1626065694
transform 1 0 86126 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_620
timestamp 1626065694
transform 1 0 86022 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_619
timestamp 1626065694
transform 1 0 88518 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_618
timestamp 1626065694
transform 1 0 91014 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_617
timestamp 1626065694
transform 1 0 93510 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_616
timestamp 1626065694
transform 1 0 98502 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_615
timestamp 1626065694
transform 1 0 100998 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_614
timestamp 1626065694
transform 1 0 96006 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_613
timestamp 1626065694
transform 1 0 77726 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_612
timestamp 1626065694
transform 1 0 79406 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_611
timestamp 1626065694
transform 1 0 81086 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_610
timestamp 1626065694
transform 1 0 82766 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_609
timestamp 1626065694
transform 1 0 84446 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_608
timestamp 1626065694
transform 1 0 69326 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_607
timestamp 1626065694
transform 1 0 71006 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_606
timestamp 1626065694
transform 1 0 72686 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_605
timestamp 1626065694
transform 1 0 74366 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_604
timestamp 1626065694
transform 1 0 76046 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_603
timestamp 1626065694
transform 1 0 73542 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_602
timestamp 1626065694
transform 1 0 76038 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_601
timestamp 1626065694
transform 1 0 68550 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_600
timestamp 1626065694
transform 1 0 71046 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_599
timestamp 1626065694
transform 1 0 83526 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_598
timestamp 1626065694
transform 1 0 78534 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_597
timestamp 1626065694
transform 1 0 81030 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_596
timestamp 1626065694
transform 1 0 134840 0 1 57132
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_595
timestamp 1626065694
transform 1 0 134840 0 1 57468
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_594
timestamp 1626065694
transform 1 0 134840 0 1 57804
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_593
timestamp 1626065694
transform 1 0 134840 0 1 58140
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_592
timestamp 1626065694
transform 1 0 134840 0 1 58476
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_591
timestamp 1626065694
transform 1 0 134840 0 1 58812
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_590
timestamp 1626065694
transform 1 0 134840 0 1 59148
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_589
timestamp 1626065694
transform 1 0 134840 0 1 59484
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_588
timestamp 1626065694
transform 1 0 134840 0 1 59820
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_587
timestamp 1626065694
transform 1 0 134840 0 1 60156
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_586
timestamp 1626065694
transform 1 0 134840 0 1 60492
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_585
timestamp 1626065694
transform 1 0 134840 0 1 60828
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_584
timestamp 1626065694
transform 1 0 134840 0 1 61164
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_583
timestamp 1626065694
transform 1 0 134840 0 1 61500
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_582
timestamp 1626065694
transform 1 0 134840 0 1 61836
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_581
timestamp 1626065694
transform 1 0 134840 0 1 62172
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_580
timestamp 1626065694
transform 1 0 134840 0 1 52428
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_579
timestamp 1626065694
transform 1 0 134840 0 1 52764
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_578
timestamp 1626065694
transform 1 0 134840 0 1 53100
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_577
timestamp 1626065694
transform 1 0 134840 0 1 53436
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_576
timestamp 1626065694
transform 1 0 134840 0 1 53772
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_575
timestamp 1626065694
transform 1 0 134840 0 1 54108
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_574
timestamp 1626065694
transform 1 0 134840 0 1 54444
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_573
timestamp 1626065694
transform 1 0 134840 0 1 54780
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_572
timestamp 1626065694
transform 1 0 134840 0 1 55116
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_571
timestamp 1626065694
transform 1 0 134840 0 1 55452
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_570
timestamp 1626065694
transform 1 0 134840 0 1 55788
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_569
timestamp 1626065694
transform 1 0 134840 0 1 56124
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_568
timestamp 1626065694
transform 1 0 134840 0 1 56460
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_567
timestamp 1626065694
transform 1 0 134840 0 1 56796
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_566
timestamp 1626065694
transform 1 0 134840 0 1 52092
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_565
timestamp 1626065694
transform 1 0 134840 0 1 48732
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_564
timestamp 1626065694
transform 1 0 134840 0 1 50412
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_563
timestamp 1626065694
transform 1 0 134840 0 1 50748
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_562
timestamp 1626065694
transform 1 0 134840 0 1 49068
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_561
timestamp 1626065694
transform 1 0 134840 0 1 50076
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_560
timestamp 1626065694
transform 1 0 134840 0 1 51084
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_559
timestamp 1626065694
transform 1 0 134840 0 1 51420
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_558
timestamp 1626065694
transform 1 0 134840 0 1 48060
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_557
timestamp 1626065694
transform 1 0 134840 0 1 51756
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_556
timestamp 1626065694
transform 1 0 134840 0 1 47388
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_555
timestamp 1626065694
transform 1 0 134840 0 1 49404
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_554
timestamp 1626065694
transform 1 0 134840 0 1 49740
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_553
timestamp 1626065694
transform 1 0 134840 0 1 48396
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_552
timestamp 1626065694
transform 1 0 134840 0 1 47052
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_551
timestamp 1626065694
transform 1 0 134840 0 1 47724
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_550
timestamp 1626065694
transform 1 0 134840 0 1 44028
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_549
timestamp 1626065694
transform 1 0 134840 0 1 45372
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_548
timestamp 1626065694
transform 1 0 134840 0 1 46044
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_547
timestamp 1626065694
transform 1 0 134840 0 1 46380
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_546
timestamp 1626065694
transform 1 0 134840 0 1 45708
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_545
timestamp 1626065694
transform 1 0 134840 0 1 41676
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_544
timestamp 1626065694
transform 1 0 134840 0 1 45036
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_543
timestamp 1626065694
transform 1 0 134840 0 1 42012
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_542
timestamp 1626065694
transform 1 0 134840 0 1 42348
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_541
timestamp 1626065694
transform 1 0 134840 0 1 42684
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_540
timestamp 1626065694
transform 1 0 134840 0 1 46716
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_539
timestamp 1626065694
transform 1 0 134840 0 1 43020
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_538
timestamp 1626065694
transform 1 0 134840 0 1 43356
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_537
timestamp 1626065694
transform 1 0 134840 0 1 43692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_536
timestamp 1626065694
transform 1 0 134840 0 1 44364
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_535
timestamp 1626065694
transform 1 0 134840 0 1 44700
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_534
timestamp 1626065694
transform 1 0 60926 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_533
timestamp 1626065694
transform 1 0 62606 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_532
timestamp 1626065694
transform 1 0 64286 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_531
timestamp 1626065694
transform 1 0 65966 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_530
timestamp 1626065694
transform 1 0 67646 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_529
timestamp 1626065694
transform 1 0 59246 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_528
timestamp 1626065694
transform 1 0 52526 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_527
timestamp 1626065694
transform 1 0 54206 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_526
timestamp 1626065694
transform 1 0 55886 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_525
timestamp 1626065694
transform 1 0 57566 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_524
timestamp 1626065694
transform 1 0 53574 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_523
timestamp 1626065694
transform 1 0 56070 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_522
timestamp 1626065694
transform 1 0 58566 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_521
timestamp 1626065694
transform 1 0 61062 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_520
timestamp 1626065694
transform 1 0 63558 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_519
timestamp 1626065694
transform 1 0 66054 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_518
timestamp 1626065694
transform 1 0 47486 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_517
timestamp 1626065694
transform 1 0 49166 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_516
timestamp 1626065694
transform 1 0 50846 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_515
timestamp 1626065694
transform 1 0 44126 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_514
timestamp 1626065694
transform 1 0 45806 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_513
timestamp 1626065694
transform 1 0 37406 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_512
timestamp 1626065694
transform 1 0 39086 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_511
timestamp 1626065694
transform 1 0 40766 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_510
timestamp 1626065694
transform 1 0 42446 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_509
timestamp 1626065694
transform 1 0 35726 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_508
timestamp 1626065694
transform 1 0 38598 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_507
timestamp 1626065694
transform 1 0 41094 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_506
timestamp 1626065694
transform 1 0 36102 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_505
timestamp 1626065694
transform 1 0 43590 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_504
timestamp 1626065694
transform 1 0 46086 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_503
timestamp 1626065694
transform 1 0 48582 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_502
timestamp 1626065694
transform 1 0 51078 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_501
timestamp 1626065694
transform 1 0 17246 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_500
timestamp 1626065694
transform 1 0 27326 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_499
timestamp 1626065694
transform 1 0 29006 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_498
timestamp 1626065694
transform 1 0 30686 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_497
timestamp 1626065694
transform 1 0 32366 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_496
timestamp 1626065694
transform 1 0 34046 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_495
timestamp 1626065694
transform 1 0 25646 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_494
timestamp 1626065694
transform 1 0 18926 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_493
timestamp 1626065694
transform 1 0 20606 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_492
timestamp 1626065694
transform 1 0 22286 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_491
timestamp 1626065694
transform 1 0 23966 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_490
timestamp 1626065694
transform 1 0 33606 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_489
timestamp 1626065694
transform 1 0 28614 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_488
timestamp 1626065694
transform 1 0 31110 0 1 76987
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_487
timestamp 1626065694
transform 1 0 8846 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_486
timestamp 1626065694
transform 1 0 10526 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_485
timestamp 1626065694
transform 1 0 12206 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_484
timestamp 1626065694
transform 1 0 13886 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_483
timestamp 1626065694
transform 1 0 15566 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_482
timestamp 1626065694
transform 1 0 5486 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_481
timestamp 1626065694
transform 1 0 7166 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_480
timestamp 1626065694
transform 1 0 3806 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_479
timestamp 1626065694
transform 1 0 1790 0 1 80652
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_478
timestamp 1626065694
transform 1 0 1790 0 1 80988
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_477
timestamp 1626065694
transform 1 0 2126 0 1 81441
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_476
timestamp 1626065694
transform 1 0 1790 0 1 78972
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_475
timestamp 1626065694
transform 1 0 1790 0 1 79308
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_474
timestamp 1626065694
transform 1 0 1790 0 1 79644
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_473
timestamp 1626065694
transform 1 0 1790 0 1 79980
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_472
timestamp 1626065694
transform 1 0 1790 0 1 80316
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_471
timestamp 1626065694
transform 1 0 1790 0 1 77964
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_470
timestamp 1626065694
transform 1 0 1790 0 1 78300
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_469
timestamp 1626065694
transform 1 0 1790 0 1 78636
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_468
timestamp 1626065694
transform 1 0 1790 0 1 73260
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_467
timestamp 1626065694
transform 1 0 1790 0 1 73596
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_466
timestamp 1626065694
transform 1 0 1790 0 1 73932
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_465
timestamp 1626065694
transform 1 0 1790 0 1 74268
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_464
timestamp 1626065694
transform 1 0 1790 0 1 74604
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_463
timestamp 1626065694
transform 1 0 1790 0 1 74940
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_462
timestamp 1626065694
transform 1 0 1790 0 1 75276
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_461
timestamp 1626065694
transform 1 0 1790 0 1 75612
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_460
timestamp 1626065694
transform 1 0 1790 0 1 76956
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_459
timestamp 1626065694
transform 1 0 1790 0 1 75948
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_458
timestamp 1626065694
transform 1 0 1790 0 1 76284
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_457
timestamp 1626065694
transform 1 0 1790 0 1 76620
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_456
timestamp 1626065694
transform 1 0 1790 0 1 77628
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_455
timestamp 1626065694
transform 1 0 1790 0 1 77292
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_454
timestamp 1626065694
transform 1 0 1790 0 1 72924
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_453
timestamp 1626065694
transform 1 0 1790 0 1 69564
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_452
timestamp 1626065694
transform 1 0 1790 0 1 69900
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_451
timestamp 1626065694
transform 1 0 1790 0 1 69228
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_450
timestamp 1626065694
transform 1 0 1790 0 1 70236
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_449
timestamp 1626065694
transform 1 0 1790 0 1 70572
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_448
timestamp 1626065694
transform 1 0 1790 0 1 70908
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_447
timestamp 1626065694
transform 1 0 1790 0 1 71244
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_446
timestamp 1626065694
transform 1 0 1790 0 1 71580
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_445
timestamp 1626065694
transform 1 0 1790 0 1 71916
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_444
timestamp 1626065694
transform 1 0 1790 0 1 72252
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_443
timestamp 1626065694
transform 1 0 1790 0 1 72588
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_442
timestamp 1626065694
transform 1 0 1790 0 1 68556
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_441
timestamp 1626065694
transform 1 0 1790 0 1 68892
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_440
timestamp 1626065694
transform 1 0 1790 0 1 67548
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_439
timestamp 1626065694
transform 1 0 1790 0 1 67884
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_438
timestamp 1626065694
transform 1 0 1790 0 1 68220
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_437
timestamp 1626065694
transform 1 0 1790 0 1 63516
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_436
timestamp 1626065694
transform 1 0 1790 0 1 63852
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_435
timestamp 1626065694
transform 1 0 1790 0 1 64188
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_434
timestamp 1626065694
transform 1 0 1790 0 1 64524
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_433
timestamp 1626065694
transform 1 0 1790 0 1 64860
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_432
timestamp 1626065694
transform 1 0 1790 0 1 65196
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_431
timestamp 1626065694
transform 1 0 1790 0 1 65532
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_430
timestamp 1626065694
transform 1 0 1790 0 1 65868
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_429
timestamp 1626065694
transform 1 0 1790 0 1 66204
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_428
timestamp 1626065694
transform 1 0 1790 0 1 66540
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_427
timestamp 1626065694
transform 1 0 1790 0 1 66876
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_426
timestamp 1626065694
transform 1 0 1790 0 1 67212
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_425
timestamp 1626065694
transform 1 0 1790 0 1 62508
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_424
timestamp 1626065694
transform 1 0 1790 0 1 62844
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_423
timestamp 1626065694
transform 1 0 1790 0 1 63180
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_422
timestamp 1626065694
transform 1 0 1790 0 1 57132
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_421
timestamp 1626065694
transform 1 0 1790 0 1 57468
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_420
timestamp 1626065694
transform 1 0 1790 0 1 57804
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_419
timestamp 1626065694
transform 1 0 1790 0 1 58140
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_418
timestamp 1626065694
transform 1 0 1790 0 1 58476
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_417
timestamp 1626065694
transform 1 0 1790 0 1 58812
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_416
timestamp 1626065694
transform 1 0 1790 0 1 59148
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_415
timestamp 1626065694
transform 1 0 1790 0 1 59484
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_414
timestamp 1626065694
transform 1 0 1790 0 1 59820
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_413
timestamp 1626065694
transform 1 0 1790 0 1 60156
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_412
timestamp 1626065694
transform 1 0 1790 0 1 60492
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_411
timestamp 1626065694
transform 1 0 1790 0 1 60828
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_410
timestamp 1626065694
transform 1 0 1790 0 1 61164
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_409
timestamp 1626065694
transform 1 0 1790 0 1 61500
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_408
timestamp 1626065694
transform 1 0 1790 0 1 61836
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_407
timestamp 1626065694
transform 1 0 1790 0 1 62172
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_406
timestamp 1626065694
transform 1 0 1790 0 1 56796
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_405
timestamp 1626065694
transform 1 0 1790 0 1 54108
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_404
timestamp 1626065694
transform 1 0 1790 0 1 54444
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_403
timestamp 1626065694
transform 1 0 1790 0 1 54780
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_402
timestamp 1626065694
transform 1 0 1790 0 1 55116
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_401
timestamp 1626065694
transform 1 0 1790 0 1 55452
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_400
timestamp 1626065694
transform 1 0 1790 0 1 55788
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_399
timestamp 1626065694
transform 1 0 1790 0 1 56124
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_398
timestamp 1626065694
transform 1 0 1790 0 1 56460
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_397
timestamp 1626065694
transform 1 0 1790 0 1 52764
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_396
timestamp 1626065694
transform 1 0 1790 0 1 52428
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_395
timestamp 1626065694
transform 1 0 1790 0 1 52092
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_394
timestamp 1626065694
transform 1 0 1790 0 1 53100
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_393
timestamp 1626065694
transform 1 0 1790 0 1 53436
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_392
timestamp 1626065694
transform 1 0 1790 0 1 53772
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_391
timestamp 1626065694
transform 1 0 1790 0 1 49740
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_390
timestamp 1626065694
transform 1 0 1790 0 1 50748
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_389
timestamp 1626065694
transform 1 0 1790 0 1 49068
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_388
timestamp 1626065694
transform 1 0 1790 0 1 51084
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_387
timestamp 1626065694
transform 1 0 1790 0 1 51756
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_386
timestamp 1626065694
transform 1 0 1790 0 1 47052
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_385
timestamp 1626065694
transform 1 0 1790 0 1 47388
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_384
timestamp 1626065694
transform 1 0 1790 0 1 51420
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_383
timestamp 1626065694
transform 1 0 1790 0 1 49404
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_382
timestamp 1626065694
transform 1 0 1790 0 1 48732
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_381
timestamp 1626065694
transform 1 0 1790 0 1 50076
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_380
timestamp 1626065694
transform 1 0 1790 0 1 50412
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_379
timestamp 1626065694
transform 1 0 1790 0 1 47724
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_378
timestamp 1626065694
transform 1 0 1790 0 1 48060
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_377
timestamp 1626065694
transform 1 0 1790 0 1 48396
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_376
timestamp 1626065694
transform 1 0 1790 0 1 41676
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_375
timestamp 1626065694
transform 1 0 1790 0 1 46044
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_374
timestamp 1626065694
transform 1 0 1790 0 1 46380
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_373
timestamp 1626065694
transform 1 0 1790 0 1 42012
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_372
timestamp 1626065694
transform 1 0 1790 0 1 46716
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_371
timestamp 1626065694
transform 1 0 1790 0 1 42348
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_370
timestamp 1626065694
transform 1 0 1790 0 1 42684
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_369
timestamp 1626065694
transform 1 0 1790 0 1 43020
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_368
timestamp 1626065694
transform 1 0 1790 0 1 43356
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_367
timestamp 1626065694
transform 1 0 1790 0 1 43692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_366
timestamp 1626065694
transform 1 0 1790 0 1 44028
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_365
timestamp 1626065694
transform 1 0 1790 0 1 44364
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_364
timestamp 1626065694
transform 1 0 1790 0 1 44700
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_363
timestamp 1626065694
transform 1 0 1790 0 1 45036
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_362
timestamp 1626065694
transform 1 0 1790 0 1 45372
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_361
timestamp 1626065694
transform 1 0 1790 0 1 45708
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_360
timestamp 1626065694
transform 1 0 1790 0 1 31260
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_359
timestamp 1626065694
transform 1 0 15343 0 1 36833
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_358
timestamp 1626065694
transform 1 0 1790 0 1 37308
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_357
timestamp 1626065694
transform 1 0 1790 0 1 37644
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_356
timestamp 1626065694
transform 1 0 1790 0 1 37980
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_355
timestamp 1626065694
transform 1 0 1790 0 1 38316
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_354
timestamp 1626065694
transform 1 0 1790 0 1 38652
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_353
timestamp 1626065694
transform 1 0 1790 0 1 38988
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_352
timestamp 1626065694
transform 1 0 1790 0 1 39324
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_351
timestamp 1626065694
transform 1 0 1790 0 1 39660
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_350
timestamp 1626065694
transform 1 0 1790 0 1 39996
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_349
timestamp 1626065694
transform 1 0 1790 0 1 40332
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_348
timestamp 1626065694
transform 1 0 1790 0 1 40668
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_347
timestamp 1626065694
transform 1 0 1790 0 1 41004
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_346
timestamp 1626065694
transform 1 0 1790 0 1 41340
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_345
timestamp 1626065694
transform 1 0 1790 0 1 36972
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_344
timestamp 1626065694
transform 1 0 1790 0 1 36636
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_343
timestamp 1626065694
transform 1 0 1790 0 1 32604
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_342
timestamp 1626065694
transform 1 0 1790 0 1 32940
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_341
timestamp 1626065694
transform 1 0 1790 0 1 33276
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_340
timestamp 1626065694
transform 1 0 1790 0 1 33612
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_339
timestamp 1626065694
transform 1 0 1790 0 1 33948
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_338
timestamp 1626065694
transform 1 0 1790 0 1 34284
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_337
timestamp 1626065694
transform 1 0 1790 0 1 34620
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_336
timestamp 1626065694
transform 1 0 1790 0 1 31932
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_335
timestamp 1626065694
transform 1 0 1790 0 1 31596
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_334
timestamp 1626065694
transform 1 0 1790 0 1 34956
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_333
timestamp 1626065694
transform 1 0 1790 0 1 35292
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_332
timestamp 1626065694
transform 1 0 1790 0 1 35628
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_331
timestamp 1626065694
transform 1 0 1790 0 1 35964
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_330
timestamp 1626065694
transform 1 0 1790 0 1 36300
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_329
timestamp 1626065694
transform 1 0 1790 0 1 32268
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_328
timestamp 1626065694
transform 1 0 15183 0 1 34005
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_327
timestamp 1626065694
transform 1 0 15263 0 1 35563
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_326
timestamp 1626065694
transform 1 0 15103 0 1 32735
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_325
timestamp 1626065694
transform 1 0 15023 0 1 31177
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_324
timestamp 1626065694
transform 1 0 14863 0 1 28349
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_323
timestamp 1626065694
transform 1 0 14943 0 1 29907
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_322
timestamp 1626065694
transform 1 0 1790 0 1 26220
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_321
timestamp 1626065694
transform 1 0 1790 0 1 26556
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_320
timestamp 1626065694
transform 1 0 1790 0 1 26892
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_319
timestamp 1626065694
transform 1 0 1790 0 1 27228
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_318
timestamp 1626065694
transform 1 0 1790 0 1 27564
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_317
timestamp 1626065694
transform 1 0 1790 0 1 27900
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_316
timestamp 1626065694
transform 1 0 1790 0 1 28236
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_315
timestamp 1626065694
transform 1 0 1790 0 1 28572
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_314
timestamp 1626065694
transform 1 0 1790 0 1 28908
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_313
timestamp 1626065694
transform 1 0 1790 0 1 30252
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_312
timestamp 1626065694
transform 1 0 1790 0 1 29244
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_311
timestamp 1626065694
transform 1 0 1790 0 1 30588
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_310
timestamp 1626065694
transform 1 0 1790 0 1 30924
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_309
timestamp 1626065694
transform 1 0 1790 0 1 29580
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_308
timestamp 1626065694
transform 1 0 1790 0 1 29916
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_307
timestamp 1626065694
transform 1 0 1790 0 1 21516
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_306
timestamp 1626065694
transform 1 0 1790 0 1 22860
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_305
timestamp 1626065694
transform 1 0 1790 0 1 21852
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_304
timestamp 1626065694
transform 1 0 1790 0 1 23196
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_303
timestamp 1626065694
transform 1 0 1790 0 1 23532
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_302
timestamp 1626065694
transform 1 0 1790 0 1 23868
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_301
timestamp 1626065694
transform 1 0 1790 0 1 25212
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_300
timestamp 1626065694
transform 1 0 1790 0 1 25548
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_299
timestamp 1626065694
transform 1 0 1790 0 1 25884
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_298
timestamp 1626065694
transform 1 0 1790 0 1 22188
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_297
timestamp 1626065694
transform 1 0 1790 0 1 24540
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_296
timestamp 1626065694
transform 1 0 1790 0 1 24876
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_295
timestamp 1626065694
transform 1 0 1790 0 1 21180
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_294
timestamp 1626065694
transform 1 0 1790 0 1 24204
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_293
timestamp 1626065694
transform 1 0 1790 0 1 22524
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_292
timestamp 1626065694
transform 1 0 17246 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_291
timestamp 1626065694
transform 1 0 28614 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_290
timestamp 1626065694
transform 1 0 31110 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_289
timestamp 1626065694
transform 1 0 33606 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_288
timestamp 1626065694
transform 1 0 1790 0 1 17148
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_287
timestamp 1626065694
transform 1 0 1790 0 1 17484
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_286
timestamp 1626065694
transform 1 0 1790 0 1 17820
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_285
timestamp 1626065694
transform 1 0 1790 0 1 18156
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_284
timestamp 1626065694
transform 1 0 1790 0 1 18492
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_283
timestamp 1626065694
transform 1 0 1790 0 1 18828
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_282
timestamp 1626065694
transform 1 0 1790 0 1 19164
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_281
timestamp 1626065694
transform 1 0 1790 0 1 19500
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_280
timestamp 1626065694
transform 1 0 1790 0 1 19836
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_279
timestamp 1626065694
transform 1 0 1790 0 1 20172
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_278
timestamp 1626065694
transform 1 0 1790 0 1 20508
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_277
timestamp 1626065694
transform 1 0 1790 0 1 20844
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_276
timestamp 1626065694
transform 1 0 1790 0 1 16140
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_275
timestamp 1626065694
transform 1 0 1790 0 1 16476
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_274
timestamp 1626065694
transform 1 0 1790 0 1 16812
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_273
timestamp 1626065694
transform 1 0 1790 0 1 15804
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_272
timestamp 1626065694
transform 1 0 1790 0 1 11436
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_271
timestamp 1626065694
transform 1 0 1790 0 1 11772
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_270
timestamp 1626065694
transform 1 0 1790 0 1 13788
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_269
timestamp 1626065694
transform 1 0 1790 0 1 12108
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_268
timestamp 1626065694
transform 1 0 1790 0 1 12444
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_267
timestamp 1626065694
transform 1 0 1790 0 1 12780
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_266
timestamp 1626065694
transform 1 0 1790 0 1 14124
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_265
timestamp 1626065694
transform 1 0 1790 0 1 14460
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_264
timestamp 1626065694
transform 1 0 1790 0 1 10764
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_263
timestamp 1626065694
transform 1 0 1790 0 1 11100
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_262
timestamp 1626065694
transform 1 0 1790 0 1 14796
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_261
timestamp 1626065694
transform 1 0 1790 0 1 15132
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_260
timestamp 1626065694
transform 1 0 1790 0 1 15468
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_259
timestamp 1626065694
transform 1 0 1790 0 1 13116
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_258
timestamp 1626065694
transform 1 0 1790 0 1 13452
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_257
timestamp 1626065694
transform 1 0 1790 0 1 5388
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_256
timestamp 1626065694
transform 1 0 1790 0 1 5724
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_255
timestamp 1626065694
transform 1 0 1790 0 1 6060
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_254
timestamp 1626065694
transform 1 0 1790 0 1 6396
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_253
timestamp 1626065694
transform 1 0 1790 0 1 6732
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_252
timestamp 1626065694
transform 1 0 1790 0 1 7068
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_251
timestamp 1626065694
transform 1 0 1790 0 1 7404
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_250
timestamp 1626065694
transform 1 0 1790 0 1 7740
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_249
timestamp 1626065694
transform 1 0 1790 0 1 8076
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_248
timestamp 1626065694
transform 1 0 1790 0 1 8412
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_247
timestamp 1626065694
transform 1 0 1790 0 1 8748
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_246
timestamp 1626065694
transform 1 0 1790 0 1 9084
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_245
timestamp 1626065694
transform 1 0 1790 0 1 9420
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_244
timestamp 1626065694
transform 1 0 1790 0 1 9756
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_243
timestamp 1626065694
transform 1 0 1790 0 1 10092
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_242
timestamp 1626065694
transform 1 0 1790 0 1 10428
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_241
timestamp 1626065694
transform 1 0 1790 0 1 4380
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_240
timestamp 1626065694
transform 1 0 1790 0 1 4716
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_239
timestamp 1626065694
transform 1 0 1790 0 1 5052
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_238
timestamp 1626065694
transform 1 0 1790 0 1 3036
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_237
timestamp 1626065694
transform 1 0 1790 0 1 3372
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_236
timestamp 1626065694
transform 1 0 1790 0 1 3708
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_235
timestamp 1626065694
transform 1 0 1790 0 1 4044
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_234
timestamp 1626065694
transform 1 0 1790 0 1 2028
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_233
timestamp 1626065694
transform 1 0 1790 0 1 2364
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_232
timestamp 1626065694
transform 1 0 1790 0 1 2700
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_231
timestamp 1626065694
transform 1 0 2126 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_230
timestamp 1626065694
transform 1 0 3806 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_229
timestamp 1626065694
transform 1 0 7166 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_228
timestamp 1626065694
transform 1 0 5486 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_227
timestamp 1626065694
transform 1 0 13886 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_226
timestamp 1626065694
transform 1 0 15566 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_225
timestamp 1626065694
transform 1 0 10526 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_224
timestamp 1626065694
transform 1 0 12206 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_223
timestamp 1626065694
transform 1 0 8846 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_222
timestamp 1626065694
transform 1 0 18926 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_221
timestamp 1626065694
transform 1 0 22286 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_220
timestamp 1626065694
transform 1 0 23966 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_219
timestamp 1626065694
transform 1 0 25646 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_218
timestamp 1626065694
transform 1 0 20606 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_217
timestamp 1626065694
transform 1 0 29006 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_216
timestamp 1626065694
transform 1 0 34046 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_215
timestamp 1626065694
transform 1 0 30686 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_214
timestamp 1626065694
transform 1 0 27326 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_213
timestamp 1626065694
transform 1 0 32366 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_212
timestamp 1626065694
transform 1 0 53574 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_211
timestamp 1626065694
transform 1 0 56070 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_210
timestamp 1626065694
transform 1 0 58566 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_209
timestamp 1626065694
transform 1 0 61062 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_208
timestamp 1626065694
transform 1 0 63558 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_207
timestamp 1626065694
transform 1 0 66054 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_206
timestamp 1626065694
transform 1 0 36102 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_205
timestamp 1626065694
transform 1 0 38598 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_204
timestamp 1626065694
transform 1 0 41094 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_203
timestamp 1626065694
transform 1 0 43590 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_202
timestamp 1626065694
transform 1 0 46086 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_201
timestamp 1626065694
transform 1 0 48582 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_200
timestamp 1626065694
transform 1 0 51078 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_199
timestamp 1626065694
transform 1 0 40766 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_198
timestamp 1626065694
transform 1 0 42446 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_197
timestamp 1626065694
transform 1 0 35726 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_196
timestamp 1626065694
transform 1 0 37406 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_195
timestamp 1626065694
transform 1 0 39086 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_194
timestamp 1626065694
transform 1 0 49166 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_193
timestamp 1626065694
transform 1 0 50846 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_192
timestamp 1626065694
transform 1 0 45806 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_191
timestamp 1626065694
transform 1 0 47486 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_190
timestamp 1626065694
transform 1 0 44126 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_189
timestamp 1626065694
transform 1 0 52526 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_188
timestamp 1626065694
transform 1 0 59246 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_187
timestamp 1626065694
transform 1 0 54206 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_186
timestamp 1626065694
transform 1 0 57566 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_185
timestamp 1626065694
transform 1 0 55886 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_184
timestamp 1626065694
transform 1 0 60926 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_183
timestamp 1626065694
transform 1 0 62606 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_182
timestamp 1626065694
transform 1 0 64286 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_181
timestamp 1626065694
transform 1 0 67646 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_180
timestamp 1626065694
transform 1 0 65966 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_179
timestamp 1626065694
transform 1 0 134840 0 1 31260
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_178
timestamp 1626065694
transform 1 0 134840 0 1 36636
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_177
timestamp 1626065694
transform 1 0 134840 0 1 36972
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_176
timestamp 1626065694
transform 1 0 134840 0 1 37308
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_175
timestamp 1626065694
transform 1 0 134840 0 1 37644
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_174
timestamp 1626065694
transform 1 0 134840 0 1 37980
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_173
timestamp 1626065694
transform 1 0 134840 0 1 38316
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_172
timestamp 1626065694
transform 1 0 134840 0 1 38652
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_171
timestamp 1626065694
transform 1 0 134840 0 1 38988
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_170
timestamp 1626065694
transform 1 0 134840 0 1 39324
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_169
timestamp 1626065694
transform 1 0 134840 0 1 39660
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_168
timestamp 1626065694
transform 1 0 134840 0 1 39996
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_167
timestamp 1626065694
transform 1 0 134840 0 1 40332
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_166
timestamp 1626065694
transform 1 0 134840 0 1 40668
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_165
timestamp 1626065694
transform 1 0 134840 0 1 41004
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_164
timestamp 1626065694
transform 1 0 134840 0 1 41340
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_163
timestamp 1626065694
transform 1 0 134840 0 1 31932
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_162
timestamp 1626065694
transform 1 0 134840 0 1 32268
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_161
timestamp 1626065694
transform 1 0 134840 0 1 32604
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_160
timestamp 1626065694
transform 1 0 134840 0 1 32940
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_159
timestamp 1626065694
transform 1 0 134840 0 1 33276
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_158
timestamp 1626065694
transform 1 0 134840 0 1 33612
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_157
timestamp 1626065694
transform 1 0 134840 0 1 33948
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_156
timestamp 1626065694
transform 1 0 134840 0 1 34284
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_155
timestamp 1626065694
transform 1 0 134840 0 1 34620
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_154
timestamp 1626065694
transform 1 0 134840 0 1 34956
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_153
timestamp 1626065694
transform 1 0 134840 0 1 35292
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_152
timestamp 1626065694
transform 1 0 134840 0 1 35628
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_151
timestamp 1626065694
transform 1 0 134840 0 1 35964
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_150
timestamp 1626065694
transform 1 0 134840 0 1 36300
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_149
timestamp 1626065694
transform 1 0 134840 0 1 31596
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_148
timestamp 1626065694
transform 1 0 134840 0 1 27564
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_147
timestamp 1626065694
transform 1 0 134840 0 1 27900
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_146
timestamp 1626065694
transform 1 0 134840 0 1 28236
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_145
timestamp 1626065694
transform 1 0 134840 0 1 28572
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_144
timestamp 1626065694
transform 1 0 134840 0 1 28908
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_143
timestamp 1626065694
transform 1 0 134840 0 1 29244
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_142
timestamp 1626065694
transform 1 0 134840 0 1 29580
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_141
timestamp 1626065694
transform 1 0 134840 0 1 29916
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_140
timestamp 1626065694
transform 1 0 134840 0 1 30252
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_139
timestamp 1626065694
transform 1 0 134840 0 1 30588
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_138
timestamp 1626065694
transform 1 0 134840 0 1 30924
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_137
timestamp 1626065694
transform 1 0 134840 0 1 26220
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_136
timestamp 1626065694
transform 1 0 134840 0 1 26556
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_135
timestamp 1626065694
transform 1 0 134840 0 1 26892
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_134
timestamp 1626065694
transform 1 0 134840 0 1 27228
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_133
timestamp 1626065694
transform 1 0 134840 0 1 21516
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_132
timestamp 1626065694
transform 1 0 134840 0 1 21852
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_131
timestamp 1626065694
transform 1 0 134840 0 1 22860
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_130
timestamp 1626065694
transform 1 0 134840 0 1 22188
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_129
timestamp 1626065694
transform 1 0 134840 0 1 23196
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_128
timestamp 1626065694
transform 1 0 134840 0 1 25212
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_127
timestamp 1626065694
transform 1 0 134840 0 1 25548
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_126
timestamp 1626065694
transform 1 0 134840 0 1 25884
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_125
timestamp 1626065694
transform 1 0 134840 0 1 23532
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_124
timestamp 1626065694
transform 1 0 134840 0 1 23868
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_123
timestamp 1626065694
transform 1 0 134840 0 1 24204
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_122
timestamp 1626065694
transform 1 0 134840 0 1 24540
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_121
timestamp 1626065694
transform 1 0 134840 0 1 24876
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_120
timestamp 1626065694
transform 1 0 134840 0 1 22524
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_119
timestamp 1626065694
transform 1 0 134840 0 1 21180
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_118
timestamp 1626065694
transform 1 0 86022 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_117
timestamp 1626065694
transform 1 0 88518 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_116
timestamp 1626065694
transform 1 0 91014 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_115
timestamp 1626065694
transform 1 0 93510 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_114
timestamp 1626065694
transform 1 0 96006 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_113
timestamp 1626065694
transform 1 0 98502 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_112
timestamp 1626065694
transform 1 0 100998 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_111
timestamp 1626065694
transform 1 0 68550 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_110
timestamp 1626065694
transform 1 0 71046 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_109
timestamp 1626065694
transform 1 0 73542 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_108
timestamp 1626065694
transform 1 0 76038 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_107
timestamp 1626065694
transform 1 0 78534 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_106
timestamp 1626065694
transform 1 0 81030 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_105
timestamp 1626065694
transform 1 0 83526 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_104
timestamp 1626065694
transform 1 0 69326 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_103
timestamp 1626065694
transform 1 0 71006 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_102
timestamp 1626065694
transform 1 0 72686 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_101
timestamp 1626065694
transform 1 0 76046 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_100
timestamp 1626065694
transform 1 0 74366 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_99
timestamp 1626065694
transform 1 0 82766 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_98
timestamp 1626065694
transform 1 0 81086 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_97
timestamp 1626065694
transform 1 0 84446 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_96
timestamp 1626065694
transform 1 0 77726 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_95
timestamp 1626065694
transform 1 0 79406 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_94
timestamp 1626065694
transform 1 0 87806 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_93
timestamp 1626065694
transform 1 0 91166 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_92
timestamp 1626065694
transform 1 0 89486 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_91
timestamp 1626065694
transform 1 0 92846 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_90
timestamp 1626065694
transform 1 0 86126 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_89
timestamp 1626065694
transform 1 0 99566 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_88
timestamp 1626065694
transform 1 0 97886 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_87
timestamp 1626065694
transform 1 0 96206 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_86
timestamp 1626065694
transform 1 0 101246 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_85
timestamp 1626065694
transform 1 0 94526 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_84
timestamp 1626065694
transform 1 0 134840 0 1 15804
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_83
timestamp 1626065694
transform 1 0 134840 0 1 16140
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_82
timestamp 1626065694
transform 1 0 134840 0 1 16476
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_81
timestamp 1626065694
transform 1 0 134840 0 1 16812
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_80
timestamp 1626065694
transform 1 0 134840 0 1 17148
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_79
timestamp 1626065694
transform 1 0 134840 0 1 17484
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_78
timestamp 1626065694
transform 1 0 134840 0 1 17820
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_77
timestamp 1626065694
transform 1 0 134840 0 1 18156
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_76
timestamp 1626065694
transform 1 0 134840 0 1 18492
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_75
timestamp 1626065694
transform 1 0 134840 0 1 18828
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_74
timestamp 1626065694
transform 1 0 134840 0 1 19164
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_73
timestamp 1626065694
transform 1 0 134840 0 1 19500
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_72
timestamp 1626065694
transform 1 0 134840 0 1 19836
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_71
timestamp 1626065694
transform 1 0 134840 0 1 20172
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_70
timestamp 1626065694
transform 1 0 134840 0 1 20508
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_69
timestamp 1626065694
transform 1 0 134840 0 1 20844
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_68
timestamp 1626065694
transform 1 0 121983 0 1 19179
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_67
timestamp 1626065694
transform 1 0 121903 0 1 17621
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_66
timestamp 1626065694
transform 1 0 121823 0 1 16351
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_65
timestamp 1626065694
transform 1 0 121583 0 1 11965
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_64
timestamp 1626065694
transform 1 0 121503 0 1 10695
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_63
timestamp 1626065694
transform 1 0 121663 0 1 13523
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_62
timestamp 1626065694
transform 1 0 121743 0 1 14793
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_61
timestamp 1626065694
transform 1 0 134840 0 1 15132
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_60
timestamp 1626065694
transform 1 0 134840 0 1 15468
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_59
timestamp 1626065694
transform 1 0 134840 0 1 10764
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_58
timestamp 1626065694
transform 1 0 134840 0 1 11100
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_57
timestamp 1626065694
transform 1 0 134840 0 1 11436
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_56
timestamp 1626065694
transform 1 0 134840 0 1 11772
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_55
timestamp 1626065694
transform 1 0 134840 0 1 12108
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_54
timestamp 1626065694
transform 1 0 134840 0 1 12444
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_53
timestamp 1626065694
transform 1 0 134840 0 1 12780
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_52
timestamp 1626065694
transform 1 0 134840 0 1 13116
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_51
timestamp 1626065694
transform 1 0 134840 0 1 13452
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_50
timestamp 1626065694
transform 1 0 134840 0 1 13788
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_49
timestamp 1626065694
transform 1 0 134840 0 1 14124
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_48
timestamp 1626065694
transform 1 0 134840 0 1 14460
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_47
timestamp 1626065694
transform 1 0 134840 0 1 14796
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_46
timestamp 1626065694
transform 1 0 103494 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_45
timestamp 1626065694
transform 1 0 105990 0 1 13201
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_44
timestamp 1626065694
transform 1 0 109646 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_43
timestamp 1626065694
transform 1 0 106286 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_42
timestamp 1626065694
transform 1 0 104606 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_41
timestamp 1626065694
transform 1 0 107966 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_40
timestamp 1626065694
transform 1 0 102926 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_39
timestamp 1626065694
transform 1 0 116366 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_38
timestamp 1626065694
transform 1 0 118046 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_37
timestamp 1626065694
transform 1 0 113006 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_36
timestamp 1626065694
transform 1 0 111326 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_35
timestamp 1626065694
transform 1 0 114686 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_34
timestamp 1626065694
transform 1 0 134840 0 1 5388
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_33
timestamp 1626065694
transform 1 0 134840 0 1 5724
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_32
timestamp 1626065694
transform 1 0 134840 0 1 6060
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_31
timestamp 1626065694
transform 1 0 134840 0 1 6396
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_30
timestamp 1626065694
transform 1 0 134840 0 1 6732
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_29
timestamp 1626065694
transform 1 0 134840 0 1 7068
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_28
timestamp 1626065694
transform 1 0 134840 0 1 7404
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_27
timestamp 1626065694
transform 1 0 134840 0 1 7740
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_26
timestamp 1626065694
transform 1 0 134840 0 1 8076
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_25
timestamp 1626065694
transform 1 0 134840 0 1 8412
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_24
timestamp 1626065694
transform 1 0 134840 0 1 8748
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_23
timestamp 1626065694
transform 1 0 134840 0 1 9084
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_22
timestamp 1626065694
transform 1 0 134840 0 1 9420
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_21
timestamp 1626065694
transform 1 0 134840 0 1 9756
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_20
timestamp 1626065694
transform 1 0 134840 0 1 10092
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_19
timestamp 1626065694
transform 1 0 134840 0 1 10428
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_18
timestamp 1626065694
transform 1 0 119726 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_17
timestamp 1626065694
transform 1 0 121406 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_16
timestamp 1626065694
transform 1 0 123086 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_15
timestamp 1626065694
transform 1 0 124766 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_14
timestamp 1626065694
transform 1 0 126446 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_13
timestamp 1626065694
transform 1 0 134840 0 1 4380
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_12
timestamp 1626065694
transform 1 0 134840 0 1 4716
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_11
timestamp 1626065694
transform 1 0 134840 0 1 5052
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_10
timestamp 1626065694
transform 1 0 134840 0 1 3708
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_9
timestamp 1626065694
transform 1 0 134840 0 1 3372
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_8
timestamp 1626065694
transform 1 0 134840 0 1 4044
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_7
timestamp 1626065694
transform 1 0 134840 0 1 3036
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_6
timestamp 1626065694
transform 1 0 128126 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_5
timestamp 1626065694
transform 1 0 129806 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_4
timestamp 1626065694
transform 1 0 131486 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_3
timestamp 1626065694
transform 1 0 133166 0 1 1692
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1626065694
transform 1 0 134840 0 1 2028
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1626065694
transform 1 0 134840 0 1 2364
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1626065694
transform 1 0 134840 0 1 2700
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1259
timestamp 1626065694
transform 1 0 127793 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1258
timestamp 1626065694
transform 1 0 132161 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1257
timestamp 1626065694
transform 1 0 132497 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1256
timestamp 1626065694
transform 1 0 132833 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1255
timestamp 1626065694
transform 1 0 133169 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1254
timestamp 1626065694
transform 1 0 133505 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1253
timestamp 1626065694
transform 1 0 133841 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1252
timestamp 1626065694
transform 1 0 134177 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1251
timestamp 1626065694
transform 1 0 134843 0 1 80651
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1250
timestamp 1626065694
transform 1 0 134843 0 1 80987
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1249
timestamp 1626065694
transform 1 0 130145 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1248
timestamp 1626065694
transform 1 0 130481 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1247
timestamp 1626065694
transform 1 0 130817 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1246
timestamp 1626065694
transform 1 0 131153 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1245
timestamp 1626065694
transform 1 0 131489 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1244
timestamp 1626065694
transform 1 0 131825 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1243
timestamp 1626065694
transform 1 0 128129 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1242
timestamp 1626065694
transform 1 0 128465 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1241
timestamp 1626065694
transform 1 0 128801 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1240
timestamp 1626065694
transform 1 0 129137 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1239
timestamp 1626065694
transform 1 0 129473 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1238
timestamp 1626065694
transform 1 0 129809 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1237
timestamp 1626065694
transform 1 0 134843 0 1 79307
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1236
timestamp 1626065694
transform 1 0 134843 0 1 79643
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1235
timestamp 1626065694
transform 1 0 134843 0 1 79979
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1234
timestamp 1626065694
transform 1 0 134843 0 1 80315
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1233
timestamp 1626065694
transform 1 0 134843 0 1 77963
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1232
timestamp 1626065694
transform 1 0 134843 0 1 78299
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1231
timestamp 1626065694
transform 1 0 134843 0 1 78635
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1230
timestamp 1626065694
transform 1 0 134843 0 1 78971
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1229
timestamp 1626065694
transform 1 0 126785 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1228
timestamp 1626065694
transform 1 0 127121 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1227
timestamp 1626065694
transform 1 0 127457 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1226
timestamp 1626065694
transform 1 0 119393 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1225
timestamp 1626065694
transform 1 0 119729 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1224
timestamp 1626065694
transform 1 0 120065 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1223
timestamp 1626065694
transform 1 0 120401 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1222
timestamp 1626065694
transform 1 0 120737 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1221
timestamp 1626065694
transform 1 0 121073 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1220
timestamp 1626065694
transform 1 0 121409 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1219
timestamp 1626065694
transform 1 0 121745 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1218
timestamp 1626065694
transform 1 0 122081 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1217
timestamp 1626065694
transform 1 0 122417 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1216
timestamp 1626065694
transform 1 0 122753 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1215
timestamp 1626065694
transform 1 0 123089 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1214
timestamp 1626065694
transform 1 0 123425 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1213
timestamp 1626065694
transform 1 0 123761 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1212
timestamp 1626065694
transform 1 0 124097 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1211
timestamp 1626065694
transform 1 0 124433 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1210
timestamp 1626065694
transform 1 0 124769 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1209
timestamp 1626065694
transform 1 0 125105 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1208
timestamp 1626065694
transform 1 0 125441 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1207
timestamp 1626065694
transform 1 0 125777 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1206
timestamp 1626065694
transform 1 0 126113 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1205
timestamp 1626065694
transform 1 0 126449 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1204
timestamp 1626065694
transform 1 0 134843 0 1 77627
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1203
timestamp 1626065694
transform 1 0 134843 0 1 72923
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1202
timestamp 1626065694
transform 1 0 134843 0 1 73259
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1201
timestamp 1626065694
transform 1 0 134843 0 1 73595
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1200
timestamp 1626065694
transform 1 0 134843 0 1 73931
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1199
timestamp 1626065694
transform 1 0 134843 0 1 74267
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1198
timestamp 1626065694
transform 1 0 134843 0 1 74603
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1197
timestamp 1626065694
transform 1 0 134843 0 1 74939
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1196
timestamp 1626065694
transform 1 0 134843 0 1 75275
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1195
timestamp 1626065694
transform 1 0 134843 0 1 75611
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1194
timestamp 1626065694
transform 1 0 134843 0 1 75947
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1193
timestamp 1626065694
transform 1 0 134843 0 1 76283
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1192
timestamp 1626065694
transform 1 0 134843 0 1 76619
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1191
timestamp 1626065694
transform 1 0 134843 0 1 76955
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1190
timestamp 1626065694
transform 1 0 134843 0 1 77291
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1189
timestamp 1626065694
transform 1 0 110993 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1188
timestamp 1626065694
transform 1 0 111329 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1187
timestamp 1626065694
transform 1 0 111665 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1186
timestamp 1626065694
transform 1 0 112001 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1185
timestamp 1626065694
transform 1 0 112337 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1184
timestamp 1626065694
transform 1 0 112673 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1183
timestamp 1626065694
transform 1 0 113009 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1182
timestamp 1626065694
transform 1 0 113345 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1181
timestamp 1626065694
transform 1 0 113681 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1180
timestamp 1626065694
transform 1 0 114017 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1179
timestamp 1626065694
transform 1 0 114353 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1178
timestamp 1626065694
transform 1 0 114689 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1177
timestamp 1626065694
transform 1 0 115025 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1176
timestamp 1626065694
transform 1 0 115361 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1175
timestamp 1626065694
transform 1 0 115697 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1174
timestamp 1626065694
transform 1 0 116033 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1173
timestamp 1626065694
transform 1 0 116369 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1172
timestamp 1626065694
transform 1 0 116705 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1171
timestamp 1626065694
transform 1 0 117041 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1170
timestamp 1626065694
transform 1 0 117377 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1169
timestamp 1626065694
transform 1 0 117713 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1168
timestamp 1626065694
transform 1 0 118049 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1167
timestamp 1626065694
transform 1 0 118385 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1166
timestamp 1626065694
transform 1 0 118721 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1165
timestamp 1626065694
transform 1 0 119057 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1164
timestamp 1626065694
transform 1 0 106625 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1163
timestamp 1626065694
transform 1 0 106961 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1162
timestamp 1626065694
transform 1 0 107297 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1161
timestamp 1626065694
transform 1 0 107633 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1160
timestamp 1626065694
transform 1 0 107969 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1159
timestamp 1626065694
transform 1 0 108305 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1158
timestamp 1626065694
transform 1 0 108641 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1157
timestamp 1626065694
transform 1 0 108977 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1156
timestamp 1626065694
transform 1 0 109313 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1155
timestamp 1626065694
transform 1 0 109649 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1154
timestamp 1626065694
transform 1 0 109985 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1153
timestamp 1626065694
transform 1 0 110321 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1152
timestamp 1626065694
transform 1 0 110657 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1151
timestamp 1626065694
transform 1 0 103265 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1150
timestamp 1626065694
transform 1 0 103601 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1149
timestamp 1626065694
transform 1 0 103937 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1148
timestamp 1626065694
transform 1 0 104273 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1147
timestamp 1626065694
transform 1 0 104609 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1146
timestamp 1626065694
transform 1 0 104945 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1145
timestamp 1626065694
transform 1 0 105281 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1144
timestamp 1626065694
transform 1 0 105617 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1143
timestamp 1626065694
transform 1 0 105953 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1142
timestamp 1626065694
transform 1 0 106289 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1141
timestamp 1626065694
transform 1 0 102593 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1140
timestamp 1626065694
transform 1 0 102929 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1139
timestamp 1626065694
transform 1 0 134843 0 1 68219
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1138
timestamp 1626065694
transform 1 0 134843 0 1 68555
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1137
timestamp 1626065694
transform 1 0 134843 0 1 68891
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1136
timestamp 1626065694
transform 1 0 134843 0 1 69227
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1135
timestamp 1626065694
transform 1 0 134843 0 1 69563
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1134
timestamp 1626065694
transform 1 0 134843 0 1 69899
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1133
timestamp 1626065694
transform 1 0 134843 0 1 70235
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1132
timestamp 1626065694
transform 1 0 134843 0 1 70571
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1131
timestamp 1626065694
transform 1 0 134843 0 1 70907
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1130
timestamp 1626065694
transform 1 0 134843 0 1 71243
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1129
timestamp 1626065694
transform 1 0 134843 0 1 71579
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1128
timestamp 1626065694
transform 1 0 134843 0 1 71915
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1127
timestamp 1626065694
transform 1 0 134843 0 1 72251
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1126
timestamp 1626065694
transform 1 0 134843 0 1 72587
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1125
timestamp 1626065694
transform 1 0 134843 0 1 67547
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1124
timestamp 1626065694
transform 1 0 134843 0 1 67883
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1123
timestamp 1626065694
transform 1 0 134843 0 1 63851
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1122
timestamp 1626065694
transform 1 0 134843 0 1 64187
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1121
timestamp 1626065694
transform 1 0 134843 0 1 64523
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1120
timestamp 1626065694
transform 1 0 134843 0 1 64859
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1119
timestamp 1626065694
transform 1 0 134843 0 1 65195
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1118
timestamp 1626065694
transform 1 0 134843 0 1 65531
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1117
timestamp 1626065694
transform 1 0 134843 0 1 65867
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1116
timestamp 1626065694
transform 1 0 134843 0 1 66203
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1115
timestamp 1626065694
transform 1 0 134843 0 1 66539
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1114
timestamp 1626065694
transform 1 0 134843 0 1 66875
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1113
timestamp 1626065694
transform 1 0 134843 0 1 67211
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1112
timestamp 1626065694
transform 1 0 134843 0 1 62507
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1111
timestamp 1626065694
transform 1 0 134843 0 1 62843
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1110
timestamp 1626065694
transform 1 0 134843 0 1 63179
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1109
timestamp 1626065694
transform 1 0 134843 0 1 63515
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1108
timestamp 1626065694
transform 1 0 93857 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1107
timestamp 1626065694
transform 1 0 94193 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1106
timestamp 1626065694
transform 1 0 94529 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1105
timestamp 1626065694
transform 1 0 94865 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1104
timestamp 1626065694
transform 1 0 95201 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1103
timestamp 1626065694
transform 1 0 95537 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1102
timestamp 1626065694
transform 1 0 95873 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1101
timestamp 1626065694
transform 1 0 96209 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1100
timestamp 1626065694
transform 1 0 96545 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1099
timestamp 1626065694
transform 1 0 96881 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1098
timestamp 1626065694
transform 1 0 97217 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1097
timestamp 1626065694
transform 1 0 97553 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1096
timestamp 1626065694
transform 1 0 97889 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1095
timestamp 1626065694
transform 1 0 98225 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1094
timestamp 1626065694
transform 1 0 98561 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1093
timestamp 1626065694
transform 1 0 98897 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1092
timestamp 1626065694
transform 1 0 99233 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1091
timestamp 1626065694
transform 1 0 99569 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1090
timestamp 1626065694
transform 1 0 99905 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1089
timestamp 1626065694
transform 1 0 100241 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1088
timestamp 1626065694
transform 1 0 100577 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1087
timestamp 1626065694
transform 1 0 100913 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1086
timestamp 1626065694
transform 1 0 101249 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1085
timestamp 1626065694
transform 1 0 101585 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1084
timestamp 1626065694
transform 1 0 101921 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1083
timestamp 1626065694
transform 1 0 102257 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1082
timestamp 1626065694
transform 1 0 86465 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1081
timestamp 1626065694
transform 1 0 86801 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1080
timestamp 1626065694
transform 1 0 87137 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1079
timestamp 1626065694
transform 1 0 87473 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1078
timestamp 1626065694
transform 1 0 87809 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1077
timestamp 1626065694
transform 1 0 88145 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1076
timestamp 1626065694
transform 1 0 88481 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1075
timestamp 1626065694
transform 1 0 88817 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1074
timestamp 1626065694
transform 1 0 89153 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1073
timestamp 1626065694
transform 1 0 89489 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1072
timestamp 1626065694
transform 1 0 89825 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1071
timestamp 1626065694
transform 1 0 90161 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1070
timestamp 1626065694
transform 1 0 90497 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1069
timestamp 1626065694
transform 1 0 90833 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1068
timestamp 1626065694
transform 1 0 91169 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1067
timestamp 1626065694
transform 1 0 91505 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1066
timestamp 1626065694
transform 1 0 91841 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1065
timestamp 1626065694
transform 1 0 92177 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1064
timestamp 1626065694
transform 1 0 92513 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1063
timestamp 1626065694
transform 1 0 92849 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1062
timestamp 1626065694
transform 1 0 93185 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1061
timestamp 1626065694
transform 1 0 93521 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1060
timestamp 1626065694
transform 1 0 85457 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1059
timestamp 1626065694
transform 1 0 85793 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1058
timestamp 1626065694
transform 1 0 86129 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1057
timestamp 1626065694
transform 1 0 77057 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1056
timestamp 1626065694
transform 1 0 77393 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1055
timestamp 1626065694
transform 1 0 77729 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1054
timestamp 1626065694
transform 1 0 78065 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1053
timestamp 1626065694
transform 1 0 78401 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1052
timestamp 1626065694
transform 1 0 78737 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1051
timestamp 1626065694
transform 1 0 79073 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1050
timestamp 1626065694
transform 1 0 79409 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1049
timestamp 1626065694
transform 1 0 79745 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1048
timestamp 1626065694
transform 1 0 80081 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1047
timestamp 1626065694
transform 1 0 80417 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1046
timestamp 1626065694
transform 1 0 80753 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1045
timestamp 1626065694
transform 1 0 81089 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1044
timestamp 1626065694
transform 1 0 81425 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1043
timestamp 1626065694
transform 1 0 81761 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1042
timestamp 1626065694
transform 1 0 82097 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1041
timestamp 1626065694
transform 1 0 82433 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1040
timestamp 1626065694
transform 1 0 82769 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1039
timestamp 1626065694
transform 1 0 83105 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1038
timestamp 1626065694
transform 1 0 83441 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1037
timestamp 1626065694
transform 1 0 83777 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1036
timestamp 1626065694
transform 1 0 84113 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1035
timestamp 1626065694
transform 1 0 84449 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1034
timestamp 1626065694
transform 1 0 84785 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1033
timestamp 1626065694
transform 1 0 85121 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1032
timestamp 1626065694
transform 1 0 76385 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1031
timestamp 1626065694
transform 1 0 76721 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1030
timestamp 1626065694
transform 1 0 68993 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1029
timestamp 1626065694
transform 1 0 69329 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1028
timestamp 1626065694
transform 1 0 69665 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1027
timestamp 1626065694
transform 1 0 70001 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1026
timestamp 1626065694
transform 1 0 70337 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1025
timestamp 1626065694
transform 1 0 70673 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1024
timestamp 1626065694
transform 1 0 71009 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1023
timestamp 1626065694
transform 1 0 71345 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1022
timestamp 1626065694
transform 1 0 71681 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1021
timestamp 1626065694
transform 1 0 72017 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1020
timestamp 1626065694
transform 1 0 72353 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1019
timestamp 1626065694
transform 1 0 72689 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1018
timestamp 1626065694
transform 1 0 73025 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1017
timestamp 1626065694
transform 1 0 68321 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1016
timestamp 1626065694
transform 1 0 68657 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1015
timestamp 1626065694
transform 1 0 73361 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1014
timestamp 1626065694
transform 1 0 73697 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1013
timestamp 1626065694
transform 1 0 74033 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1012
timestamp 1626065694
transform 1 0 74369 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1011
timestamp 1626065694
transform 1 0 74705 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1010
timestamp 1626065694
transform 1 0 75041 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1009
timestamp 1626065694
transform 1 0 75377 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1008
timestamp 1626065694
transform 1 0 75713 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1007
timestamp 1626065694
transform 1 0 76049 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1006
timestamp 1626065694
transform 1 0 134843 0 1 57131
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1005
timestamp 1626065694
transform 1 0 134843 0 1 57467
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1004
timestamp 1626065694
transform 1 0 134843 0 1 57803
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1003
timestamp 1626065694
transform 1 0 134843 0 1 58139
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1002
timestamp 1626065694
transform 1 0 134843 0 1 58475
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1001
timestamp 1626065694
transform 1 0 134843 0 1 58811
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1000
timestamp 1626065694
transform 1 0 134843 0 1 59147
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_999
timestamp 1626065694
transform 1 0 134843 0 1 59483
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_998
timestamp 1626065694
transform 1 0 134843 0 1 59819
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_997
timestamp 1626065694
transform 1 0 134843 0 1 60155
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_996
timestamp 1626065694
transform 1 0 134843 0 1 60491
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_995
timestamp 1626065694
transform 1 0 134843 0 1 60827
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_994
timestamp 1626065694
transform 1 0 134843 0 1 61163
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_993
timestamp 1626065694
transform 1 0 134843 0 1 61499
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_992
timestamp 1626065694
transform 1 0 134843 0 1 61835
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_991
timestamp 1626065694
transform 1 0 134843 0 1 62171
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_990
timestamp 1626065694
transform 1 0 134843 0 1 52763
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_989
timestamp 1626065694
transform 1 0 134843 0 1 53099
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_988
timestamp 1626065694
transform 1 0 134843 0 1 53435
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_987
timestamp 1626065694
transform 1 0 134843 0 1 53771
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_986
timestamp 1626065694
transform 1 0 134843 0 1 54107
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_985
timestamp 1626065694
transform 1 0 134843 0 1 54443
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_984
timestamp 1626065694
transform 1 0 134843 0 1 54779
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_983
timestamp 1626065694
transform 1 0 134843 0 1 55115
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_982
timestamp 1626065694
transform 1 0 134843 0 1 55451
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_981
timestamp 1626065694
transform 1 0 134843 0 1 55787
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_980
timestamp 1626065694
transform 1 0 134843 0 1 56123
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_979
timestamp 1626065694
transform 1 0 134843 0 1 56459
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_978
timestamp 1626065694
transform 1 0 134843 0 1 52091
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_977
timestamp 1626065694
transform 1 0 134843 0 1 56795
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_976
timestamp 1626065694
transform 1 0 134843 0 1 52427
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_975
timestamp 1626065694
transform 1 0 134843 0 1 48731
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_974
timestamp 1626065694
transform 1 0 134843 0 1 50075
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_973
timestamp 1626065694
transform 1 0 134843 0 1 49067
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_972
timestamp 1626065694
transform 1 0 134843 0 1 50411
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_971
timestamp 1626065694
transform 1 0 134843 0 1 50747
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_970
timestamp 1626065694
transform 1 0 134843 0 1 51083
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_969
timestamp 1626065694
transform 1 0 134843 0 1 51419
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_968
timestamp 1626065694
transform 1 0 134843 0 1 48059
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_967
timestamp 1626065694
transform 1 0 134843 0 1 51755
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_966
timestamp 1626065694
transform 1 0 134843 0 1 47387
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_965
timestamp 1626065694
transform 1 0 134843 0 1 47723
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_964
timestamp 1626065694
transform 1 0 134843 0 1 48395
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_963
timestamp 1626065694
transform 1 0 134843 0 1 49403
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_962
timestamp 1626065694
transform 1 0 134843 0 1 49739
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_961
timestamp 1626065694
transform 1 0 134843 0 1 47051
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_960
timestamp 1626065694
transform 1 0 134843 0 1 45707
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_959
timestamp 1626065694
transform 1 0 134843 0 1 46379
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_958
timestamp 1626065694
transform 1 0 134843 0 1 41675
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_957
timestamp 1626065694
transform 1 0 134843 0 1 42011
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_956
timestamp 1626065694
transform 1 0 134843 0 1 45035
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_955
timestamp 1626065694
transform 1 0 134843 0 1 45371
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_954
timestamp 1626065694
transform 1 0 134843 0 1 42347
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_953
timestamp 1626065694
transform 1 0 134843 0 1 42683
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_952
timestamp 1626065694
transform 1 0 134843 0 1 46715
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_951
timestamp 1626065694
transform 1 0 134843 0 1 44699
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_950
timestamp 1626065694
transform 1 0 134843 0 1 44363
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_949
timestamp 1626065694
transform 1 0 134843 0 1 43019
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_948
timestamp 1626065694
transform 1 0 134843 0 1 43355
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_947
timestamp 1626065694
transform 1 0 134843 0 1 43691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_946
timestamp 1626065694
transform 1 0 134843 0 1 46043
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_945
timestamp 1626065694
transform 1 0 134843 0 1 44027
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_944
timestamp 1626065694
transform 1 0 59921 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_943
timestamp 1626065694
transform 1 0 60257 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_942
timestamp 1626065694
transform 1 0 60593 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_941
timestamp 1626065694
transform 1 0 60929 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_940
timestamp 1626065694
transform 1 0 61265 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_939
timestamp 1626065694
transform 1 0 61601 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_938
timestamp 1626065694
transform 1 0 61937 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_937
timestamp 1626065694
transform 1 0 62273 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_936
timestamp 1626065694
transform 1 0 62609 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_935
timestamp 1626065694
transform 1 0 62945 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_934
timestamp 1626065694
transform 1 0 63281 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_933
timestamp 1626065694
transform 1 0 63617 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_932
timestamp 1626065694
transform 1 0 63953 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_931
timestamp 1626065694
transform 1 0 64289 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_930
timestamp 1626065694
transform 1 0 64625 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_929
timestamp 1626065694
transform 1 0 64961 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_928
timestamp 1626065694
transform 1 0 65297 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_927
timestamp 1626065694
transform 1 0 65633 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_926
timestamp 1626065694
transform 1 0 65969 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_925
timestamp 1626065694
transform 1 0 66305 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_924
timestamp 1626065694
transform 1 0 66641 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_923
timestamp 1626065694
transform 1 0 66977 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_922
timestamp 1626065694
transform 1 0 67313 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_921
timestamp 1626065694
transform 1 0 67649 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_920
timestamp 1626065694
transform 1 0 67985 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_919
timestamp 1626065694
transform 1 0 58577 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_918
timestamp 1626065694
transform 1 0 58913 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_917
timestamp 1626065694
transform 1 0 59249 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_916
timestamp 1626065694
transform 1 0 59585 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_915
timestamp 1626065694
transform 1 0 51521 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_914
timestamp 1626065694
transform 1 0 51857 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_913
timestamp 1626065694
transform 1 0 52193 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_912
timestamp 1626065694
transform 1 0 52529 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_911
timestamp 1626065694
transform 1 0 52865 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_910
timestamp 1626065694
transform 1 0 53201 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_909
timestamp 1626065694
transform 1 0 53537 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_908
timestamp 1626065694
transform 1 0 53873 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_907
timestamp 1626065694
transform 1 0 54209 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_906
timestamp 1626065694
transform 1 0 54545 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_905
timestamp 1626065694
transform 1 0 54881 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_904
timestamp 1626065694
transform 1 0 55217 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_903
timestamp 1626065694
transform 1 0 55553 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_902
timestamp 1626065694
transform 1 0 55889 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_901
timestamp 1626065694
transform 1 0 56225 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_900
timestamp 1626065694
transform 1 0 56561 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_899
timestamp 1626065694
transform 1 0 56897 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_898
timestamp 1626065694
transform 1 0 57233 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_897
timestamp 1626065694
transform 1 0 57569 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_896
timestamp 1626065694
transform 1 0 57905 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_895
timestamp 1626065694
transform 1 0 58241 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_894
timestamp 1626065694
transform 1 0 42785 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_893
timestamp 1626065694
transform 1 0 46817 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_892
timestamp 1626065694
transform 1 0 47153 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_891
timestamp 1626065694
transform 1 0 47489 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_890
timestamp 1626065694
transform 1 0 47825 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_889
timestamp 1626065694
transform 1 0 48161 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_888
timestamp 1626065694
transform 1 0 48497 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_887
timestamp 1626065694
transform 1 0 48833 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_886
timestamp 1626065694
transform 1 0 49169 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_885
timestamp 1626065694
transform 1 0 49505 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_884
timestamp 1626065694
transform 1 0 49841 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_883
timestamp 1626065694
transform 1 0 50177 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_882
timestamp 1626065694
transform 1 0 50513 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_881
timestamp 1626065694
transform 1 0 50849 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_880
timestamp 1626065694
transform 1 0 51185 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_879
timestamp 1626065694
transform 1 0 43121 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_878
timestamp 1626065694
transform 1 0 43457 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_877
timestamp 1626065694
transform 1 0 43793 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_876
timestamp 1626065694
transform 1 0 44129 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_875
timestamp 1626065694
transform 1 0 44465 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_874
timestamp 1626065694
transform 1 0 44801 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_873
timestamp 1626065694
transform 1 0 45137 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_872
timestamp 1626065694
transform 1 0 45473 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_871
timestamp 1626065694
transform 1 0 45809 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_870
timestamp 1626065694
transform 1 0 46145 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_869
timestamp 1626065694
transform 1 0 46481 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_868
timestamp 1626065694
transform 1 0 37745 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_867
timestamp 1626065694
transform 1 0 38081 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_866
timestamp 1626065694
transform 1 0 38417 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_865
timestamp 1626065694
transform 1 0 38753 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_864
timestamp 1626065694
transform 1 0 39089 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_863
timestamp 1626065694
transform 1 0 39425 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_862
timestamp 1626065694
transform 1 0 39761 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_861
timestamp 1626065694
transform 1 0 40097 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_860
timestamp 1626065694
transform 1 0 40433 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_859
timestamp 1626065694
transform 1 0 40769 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_858
timestamp 1626065694
transform 1 0 41105 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_857
timestamp 1626065694
transform 1 0 41441 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_856
timestamp 1626065694
transform 1 0 41777 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_855
timestamp 1626065694
transform 1 0 42113 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_854
timestamp 1626065694
transform 1 0 42449 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_853
timestamp 1626065694
transform 1 0 34385 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_852
timestamp 1626065694
transform 1 0 34721 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_851
timestamp 1626065694
transform 1 0 35057 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_850
timestamp 1626065694
transform 1 0 35393 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_849
timestamp 1626065694
transform 1 0 35729 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_848
timestamp 1626065694
transform 1 0 36065 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_847
timestamp 1626065694
transform 1 0 36401 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_846
timestamp 1626065694
transform 1 0 36737 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_845
timestamp 1626065694
transform 1 0 37073 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_844
timestamp 1626065694
transform 1 0 37409 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_843
timestamp 1626065694
transform 1 0 17249 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_842
timestamp 1626065694
transform 1 0 25985 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_841
timestamp 1626065694
transform 1 0 26321 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_840
timestamp 1626065694
transform 1 0 26657 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_839
timestamp 1626065694
transform 1 0 26993 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_838
timestamp 1626065694
transform 1 0 27329 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_837
timestamp 1626065694
transform 1 0 27665 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_836
timestamp 1626065694
transform 1 0 28001 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_835
timestamp 1626065694
transform 1 0 28337 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_834
timestamp 1626065694
transform 1 0 28673 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_833
timestamp 1626065694
transform 1 0 29009 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_832
timestamp 1626065694
transform 1 0 29345 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_831
timestamp 1626065694
transform 1 0 29681 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_830
timestamp 1626065694
transform 1 0 30017 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_829
timestamp 1626065694
transform 1 0 30353 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_828
timestamp 1626065694
transform 1 0 30689 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_827
timestamp 1626065694
transform 1 0 31025 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_826
timestamp 1626065694
transform 1 0 31361 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_825
timestamp 1626065694
transform 1 0 31697 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_824
timestamp 1626065694
transform 1 0 32033 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_823
timestamp 1626065694
transform 1 0 32369 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_822
timestamp 1626065694
transform 1 0 32705 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_821
timestamp 1626065694
transform 1 0 33041 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_820
timestamp 1626065694
transform 1 0 33377 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_819
timestamp 1626065694
transform 1 0 33713 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_818
timestamp 1626065694
transform 1 0 34049 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_817
timestamp 1626065694
transform 1 0 25313 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_816
timestamp 1626065694
transform 1 0 25649 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_815
timestamp 1626065694
transform 1 0 17585 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_814
timestamp 1626065694
transform 1 0 17921 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_813
timestamp 1626065694
transform 1 0 18257 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_812
timestamp 1626065694
transform 1 0 18593 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_811
timestamp 1626065694
transform 1 0 18929 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_810
timestamp 1626065694
transform 1 0 19265 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_809
timestamp 1626065694
transform 1 0 19601 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_808
timestamp 1626065694
transform 1 0 19937 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_807
timestamp 1626065694
transform 1 0 20273 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_806
timestamp 1626065694
transform 1 0 20609 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_805
timestamp 1626065694
transform 1 0 20945 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_804
timestamp 1626065694
transform 1 0 21281 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_803
timestamp 1626065694
transform 1 0 21617 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_802
timestamp 1626065694
transform 1 0 21953 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_801
timestamp 1626065694
transform 1 0 22289 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_800
timestamp 1626065694
transform 1 0 22625 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_799
timestamp 1626065694
transform 1 0 22961 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_798
timestamp 1626065694
transform 1 0 23297 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_797
timestamp 1626065694
transform 1 0 23633 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_796
timestamp 1626065694
transform 1 0 23969 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_795
timestamp 1626065694
transform 1 0 24305 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_794
timestamp 1626065694
transform 1 0 24641 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_793
timestamp 1626065694
transform 1 0 24977 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_792
timestamp 1626065694
transform 1 0 9185 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_791
timestamp 1626065694
transform 1 0 9521 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_790
timestamp 1626065694
transform 1 0 9857 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_789
timestamp 1626065694
transform 1 0 10193 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_788
timestamp 1626065694
transform 1 0 10529 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_787
timestamp 1626065694
transform 1 0 10865 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_786
timestamp 1626065694
transform 1 0 11201 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_785
timestamp 1626065694
transform 1 0 11537 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_784
timestamp 1626065694
transform 1 0 11873 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_783
timestamp 1626065694
transform 1 0 12209 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_782
timestamp 1626065694
transform 1 0 12545 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_781
timestamp 1626065694
transform 1 0 12881 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_780
timestamp 1626065694
transform 1 0 13217 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_779
timestamp 1626065694
transform 1 0 13553 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_778
timestamp 1626065694
transform 1 0 13889 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_777
timestamp 1626065694
transform 1 0 14225 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_776
timestamp 1626065694
transform 1 0 14561 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_775
timestamp 1626065694
transform 1 0 14897 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_774
timestamp 1626065694
transform 1 0 15233 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_773
timestamp 1626065694
transform 1 0 15569 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_772
timestamp 1626065694
transform 1 0 15905 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_771
timestamp 1626065694
transform 1 0 16241 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_770
timestamp 1626065694
transform 1 0 16577 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_769
timestamp 1626065694
transform 1 0 16913 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_768
timestamp 1626065694
transform 1 0 8849 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_767
timestamp 1626065694
transform 1 0 4481 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_766
timestamp 1626065694
transform 1 0 4817 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_765
timestamp 1626065694
transform 1 0 5153 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_764
timestamp 1626065694
transform 1 0 5489 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_763
timestamp 1626065694
transform 1 0 5825 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_762
timestamp 1626065694
transform 1 0 6161 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_761
timestamp 1626065694
transform 1 0 6497 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_760
timestamp 1626065694
transform 1 0 6833 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_759
timestamp 1626065694
transform 1 0 7169 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_758
timestamp 1626065694
transform 1 0 7505 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_757
timestamp 1626065694
transform 1 0 7841 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_756
timestamp 1626065694
transform 1 0 8177 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_755
timestamp 1626065694
transform 1 0 8513 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_754
timestamp 1626065694
transform 1 0 3809 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_753
timestamp 1626065694
transform 1 0 4145 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_752
timestamp 1626065694
transform 1 0 1793 0 1 80651
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_751
timestamp 1626065694
transform 1 0 1793 0 1 80987
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_750
timestamp 1626065694
transform 1 0 2129 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_749
timestamp 1626065694
transform 1 0 2465 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_748
timestamp 1626065694
transform 1 0 2801 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_747
timestamp 1626065694
transform 1 0 3137 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_746
timestamp 1626065694
transform 1 0 3473 0 1 81440
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_745
timestamp 1626065694
transform 1 0 1793 0 1 78971
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_744
timestamp 1626065694
transform 1 0 1793 0 1 79307
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_743
timestamp 1626065694
transform 1 0 1793 0 1 79643
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_742
timestamp 1626065694
transform 1 0 1793 0 1 79979
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_741
timestamp 1626065694
transform 1 0 1793 0 1 80315
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_740
timestamp 1626065694
transform 1 0 1793 0 1 77963
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_739
timestamp 1626065694
transform 1 0 1793 0 1 78299
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_738
timestamp 1626065694
transform 1 0 1793 0 1 78635
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_737
timestamp 1626065694
transform 1 0 1793 0 1 73259
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_736
timestamp 1626065694
transform 1 0 1793 0 1 73595
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_735
timestamp 1626065694
transform 1 0 1793 0 1 73931
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_734
timestamp 1626065694
transform 1 0 1793 0 1 74267
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_733
timestamp 1626065694
transform 1 0 1793 0 1 74603
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_732
timestamp 1626065694
transform 1 0 1793 0 1 74939
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_731
timestamp 1626065694
transform 1 0 1793 0 1 75275
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_730
timestamp 1626065694
transform 1 0 1793 0 1 75611
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_729
timestamp 1626065694
transform 1 0 1793 0 1 76955
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_728
timestamp 1626065694
transform 1 0 1793 0 1 75947
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_727
timestamp 1626065694
transform 1 0 1793 0 1 76283
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_726
timestamp 1626065694
transform 1 0 1793 0 1 76619
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_725
timestamp 1626065694
transform 1 0 1793 0 1 77627
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_724
timestamp 1626065694
transform 1 0 1793 0 1 77291
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_723
timestamp 1626065694
transform 1 0 1793 0 1 72923
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_722
timestamp 1626065694
transform 1 0 1793 0 1 69563
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_721
timestamp 1626065694
transform 1 0 1793 0 1 69899
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_720
timestamp 1626065694
transform 1 0 1793 0 1 70235
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_719
timestamp 1626065694
transform 1 0 1793 0 1 70571
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_718
timestamp 1626065694
transform 1 0 1793 0 1 70907
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_717
timestamp 1626065694
transform 1 0 1793 0 1 71243
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_716
timestamp 1626065694
transform 1 0 1793 0 1 71579
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_715
timestamp 1626065694
transform 1 0 1793 0 1 71915
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_714
timestamp 1626065694
transform 1 0 1793 0 1 72251
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_713
timestamp 1626065694
transform 1 0 1793 0 1 72587
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_712
timestamp 1626065694
transform 1 0 1793 0 1 68555
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_711
timestamp 1626065694
transform 1 0 1793 0 1 68891
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_710
timestamp 1626065694
transform 1 0 1793 0 1 69227
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_709
timestamp 1626065694
transform 1 0 1793 0 1 67547
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_708
timestamp 1626065694
transform 1 0 1793 0 1 67883
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_707
timestamp 1626065694
transform 1 0 1793 0 1 68219
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_706
timestamp 1626065694
transform 1 0 1793 0 1 63515
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_705
timestamp 1626065694
transform 1 0 1793 0 1 63851
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_704
timestamp 1626065694
transform 1 0 1793 0 1 64187
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_703
timestamp 1626065694
transform 1 0 1793 0 1 64523
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_702
timestamp 1626065694
transform 1 0 1793 0 1 64859
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_701
timestamp 1626065694
transform 1 0 1793 0 1 65195
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_700
timestamp 1626065694
transform 1 0 1793 0 1 65531
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_699
timestamp 1626065694
transform 1 0 1793 0 1 65867
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_698
timestamp 1626065694
transform 1 0 1793 0 1 66203
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_697
timestamp 1626065694
transform 1 0 1793 0 1 66539
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_696
timestamp 1626065694
transform 1 0 1793 0 1 66875
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_695
timestamp 1626065694
transform 1 0 1793 0 1 67211
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_694
timestamp 1626065694
transform 1 0 1793 0 1 62507
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_693
timestamp 1626065694
transform 1 0 1793 0 1 62843
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_692
timestamp 1626065694
transform 1 0 1793 0 1 63179
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_691
timestamp 1626065694
transform 1 0 1793 0 1 57131
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_690
timestamp 1626065694
transform 1 0 1793 0 1 57467
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_689
timestamp 1626065694
transform 1 0 1793 0 1 57803
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_688
timestamp 1626065694
transform 1 0 1793 0 1 58139
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_687
timestamp 1626065694
transform 1 0 1793 0 1 58475
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_686
timestamp 1626065694
transform 1 0 1793 0 1 58811
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_685
timestamp 1626065694
transform 1 0 1793 0 1 59147
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_684
timestamp 1626065694
transform 1 0 1793 0 1 59483
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_683
timestamp 1626065694
transform 1 0 1793 0 1 59819
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_682
timestamp 1626065694
transform 1 0 1793 0 1 60155
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_681
timestamp 1626065694
transform 1 0 1793 0 1 60491
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_680
timestamp 1626065694
transform 1 0 1793 0 1 60827
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_679
timestamp 1626065694
transform 1 0 1793 0 1 61163
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_678
timestamp 1626065694
transform 1 0 1793 0 1 61499
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_677
timestamp 1626065694
transform 1 0 1793 0 1 61835
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_676
timestamp 1626065694
transform 1 0 1793 0 1 62171
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_675
timestamp 1626065694
transform 1 0 1793 0 1 56795
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_674
timestamp 1626065694
transform 1 0 1793 0 1 54107
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_673
timestamp 1626065694
transform 1 0 1793 0 1 54443
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_672
timestamp 1626065694
transform 1 0 1793 0 1 54779
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_671
timestamp 1626065694
transform 1 0 1793 0 1 55115
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_670
timestamp 1626065694
transform 1 0 1793 0 1 55451
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_669
timestamp 1626065694
transform 1 0 1793 0 1 55787
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_668
timestamp 1626065694
transform 1 0 1793 0 1 56123
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_667
timestamp 1626065694
transform 1 0 1793 0 1 56459
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_666
timestamp 1626065694
transform 1 0 1793 0 1 52427
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_665
timestamp 1626065694
transform 1 0 1793 0 1 52763
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_664
timestamp 1626065694
transform 1 0 1793 0 1 52091
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_663
timestamp 1626065694
transform 1 0 1793 0 1 53099
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_662
timestamp 1626065694
transform 1 0 1793 0 1 53435
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_661
timestamp 1626065694
transform 1 0 1793 0 1 53771
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_660
timestamp 1626065694
transform 1 0 1793 0 1 49739
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_659
timestamp 1626065694
transform 1 0 1793 0 1 50075
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_658
timestamp 1626065694
transform 1 0 1793 0 1 50747
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_657
timestamp 1626065694
transform 1 0 1793 0 1 51083
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_656
timestamp 1626065694
transform 1 0 1793 0 1 47051
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_655
timestamp 1626065694
transform 1 0 1793 0 1 47387
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_654
timestamp 1626065694
transform 1 0 1793 0 1 51419
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_653
timestamp 1626065694
transform 1 0 1793 0 1 49403
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_652
timestamp 1626065694
transform 1 0 1793 0 1 48731
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_651
timestamp 1626065694
transform 1 0 1793 0 1 47723
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_650
timestamp 1626065694
transform 1 0 1793 0 1 50411
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_649
timestamp 1626065694
transform 1 0 1793 0 1 49067
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_648
timestamp 1626065694
transform 1 0 1793 0 1 51755
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_647
timestamp 1626065694
transform 1 0 1793 0 1 48059
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_646
timestamp 1626065694
transform 1 0 1793 0 1 48395
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_645
timestamp 1626065694
transform 1 0 1793 0 1 42011
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_644
timestamp 1626065694
transform 1 0 1793 0 1 46043
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_643
timestamp 1626065694
transform 1 0 1793 0 1 46379
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_642
timestamp 1626065694
transform 1 0 1793 0 1 46715
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_641
timestamp 1626065694
transform 1 0 1793 0 1 42347
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_640
timestamp 1626065694
transform 1 0 1793 0 1 42683
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_639
timestamp 1626065694
transform 1 0 1793 0 1 43019
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_638
timestamp 1626065694
transform 1 0 1793 0 1 43355
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_637
timestamp 1626065694
transform 1 0 1793 0 1 43691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_636
timestamp 1626065694
transform 1 0 1793 0 1 44027
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_635
timestamp 1626065694
transform 1 0 1793 0 1 44363
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_634
timestamp 1626065694
transform 1 0 1793 0 1 44699
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_633
timestamp 1626065694
transform 1 0 1793 0 1 45035
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_632
timestamp 1626065694
transform 1 0 1793 0 1 45371
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_631
timestamp 1626065694
transform 1 0 1793 0 1 45707
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_630
timestamp 1626065694
transform 1 0 1793 0 1 41675
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_629
timestamp 1626065694
transform 1 0 1793 0 1 31259
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_628
timestamp 1626065694
transform 1 0 1793 0 1 36971
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_627
timestamp 1626065694
transform 1 0 1793 0 1 37643
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_626
timestamp 1626065694
transform 1 0 1793 0 1 37979
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_625
timestamp 1626065694
transform 1 0 1793 0 1 38315
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_624
timestamp 1626065694
transform 1 0 1793 0 1 38651
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_623
timestamp 1626065694
transform 1 0 1793 0 1 38987
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_622
timestamp 1626065694
transform 1 0 1793 0 1 39323
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_621
timestamp 1626065694
transform 1 0 1793 0 1 39659
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_620
timestamp 1626065694
transform 1 0 1793 0 1 39995
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_619
timestamp 1626065694
transform 1 0 1793 0 1 40331
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_618
timestamp 1626065694
transform 1 0 1793 0 1 40667
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_617
timestamp 1626065694
transform 1 0 1793 0 1 41003
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_616
timestamp 1626065694
transform 1 0 1793 0 1 41339
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_615
timestamp 1626065694
transform 1 0 1793 0 1 37307
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_614
timestamp 1626065694
transform 1 0 1793 0 1 36635
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_613
timestamp 1626065694
transform 1 0 1793 0 1 32267
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_612
timestamp 1626065694
transform 1 0 1793 0 1 32603
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_611
timestamp 1626065694
transform 1 0 1793 0 1 32939
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_610
timestamp 1626065694
transform 1 0 1793 0 1 33275
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_609
timestamp 1626065694
transform 1 0 1793 0 1 33611
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_608
timestamp 1626065694
transform 1 0 1793 0 1 33947
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_607
timestamp 1626065694
transform 1 0 1793 0 1 34283
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_606
timestamp 1626065694
transform 1 0 1793 0 1 34619
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_605
timestamp 1626065694
transform 1 0 1793 0 1 31595
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_604
timestamp 1626065694
transform 1 0 1793 0 1 34955
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_603
timestamp 1626065694
transform 1 0 1793 0 1 35291
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_602
timestamp 1626065694
transform 1 0 1793 0 1 35627
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_601
timestamp 1626065694
transform 1 0 1793 0 1 35963
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_600
timestamp 1626065694
transform 1 0 1793 0 1 36299
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_599
timestamp 1626065694
transform 1 0 1793 0 1 31931
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_598
timestamp 1626065694
transform 1 0 1793 0 1 26555
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_597
timestamp 1626065694
transform 1 0 1793 0 1 26891
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_596
timestamp 1626065694
transform 1 0 1793 0 1 27227
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_595
timestamp 1626065694
transform 1 0 1793 0 1 27563
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_594
timestamp 1626065694
transform 1 0 1793 0 1 27899
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_593
timestamp 1626065694
transform 1 0 1793 0 1 28235
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_592
timestamp 1626065694
transform 1 0 1793 0 1 28571
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_591
timestamp 1626065694
transform 1 0 1793 0 1 28907
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_590
timestamp 1626065694
transform 1 0 1793 0 1 30251
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_589
timestamp 1626065694
transform 1 0 1793 0 1 29243
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_588
timestamp 1626065694
transform 1 0 1793 0 1 29579
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_587
timestamp 1626065694
transform 1 0 1793 0 1 30587
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_586
timestamp 1626065694
transform 1 0 1793 0 1 30923
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_585
timestamp 1626065694
transform 1 0 1793 0 1 29915
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_584
timestamp 1626065694
transform 1 0 1793 0 1 26219
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_583
timestamp 1626065694
transform 1 0 1793 0 1 22859
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_582
timestamp 1626065694
transform 1 0 1793 0 1 21851
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_581
timestamp 1626065694
transform 1 0 1793 0 1 25211
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_580
timestamp 1626065694
transform 1 0 1793 0 1 23195
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_579
timestamp 1626065694
transform 1 0 1793 0 1 23531
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_578
timestamp 1626065694
transform 1 0 1793 0 1 23867
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_577
timestamp 1626065694
transform 1 0 1793 0 1 25547
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_576
timestamp 1626065694
transform 1 0 1793 0 1 25883
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_575
timestamp 1626065694
transform 1 0 1793 0 1 24539
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_574
timestamp 1626065694
transform 1 0 1793 0 1 22187
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_573
timestamp 1626065694
transform 1 0 1793 0 1 24875
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_572
timestamp 1626065694
transform 1 0 1793 0 1 21179
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_571
timestamp 1626065694
transform 1 0 1793 0 1 24203
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_570
timestamp 1626065694
transform 1 0 1793 0 1 22523
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_569
timestamp 1626065694
transform 1 0 1793 0 1 21515
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_568
timestamp 1626065694
transform 1 0 17249 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_567
timestamp 1626065694
transform 1 0 1793 0 1 17483
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_566
timestamp 1626065694
transform 1 0 1793 0 1 17819
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_565
timestamp 1626065694
transform 1 0 1793 0 1 18155
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_564
timestamp 1626065694
transform 1 0 1793 0 1 18491
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_563
timestamp 1626065694
transform 1 0 1793 0 1 18827
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_562
timestamp 1626065694
transform 1 0 1793 0 1 19163
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_561
timestamp 1626065694
transform 1 0 1793 0 1 19499
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_560
timestamp 1626065694
transform 1 0 1793 0 1 19835
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_559
timestamp 1626065694
transform 1 0 1793 0 1 20171
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_558
timestamp 1626065694
transform 1 0 1793 0 1 20507
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_557
timestamp 1626065694
transform 1 0 1793 0 1 20843
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_556
timestamp 1626065694
transform 1 0 1793 0 1 16139
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_555
timestamp 1626065694
transform 1 0 1793 0 1 16475
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_554
timestamp 1626065694
transform 1 0 1793 0 1 16811
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_553
timestamp 1626065694
transform 1 0 1793 0 1 17147
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_552
timestamp 1626065694
transform 1 0 1793 0 1 15803
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_551
timestamp 1626065694
transform 1 0 1793 0 1 13787
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_550
timestamp 1626065694
transform 1 0 1793 0 1 11771
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_549
timestamp 1626065694
transform 1 0 1793 0 1 11435
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_548
timestamp 1626065694
transform 1 0 1793 0 1 12107
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_547
timestamp 1626065694
transform 1 0 1793 0 1 14123
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_546
timestamp 1626065694
transform 1 0 1793 0 1 12443
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_545
timestamp 1626065694
transform 1 0 1793 0 1 12779
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_544
timestamp 1626065694
transform 1 0 1793 0 1 13115
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_543
timestamp 1626065694
transform 1 0 1793 0 1 14459
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_542
timestamp 1626065694
transform 1 0 1793 0 1 10763
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_541
timestamp 1626065694
transform 1 0 1793 0 1 14795
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_540
timestamp 1626065694
transform 1 0 1793 0 1 11099
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_539
timestamp 1626065694
transform 1 0 1793 0 1 15131
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_538
timestamp 1626065694
transform 1 0 1793 0 1 15467
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_537
timestamp 1626065694
transform 1 0 1793 0 1 13451
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_536
timestamp 1626065694
transform 1 0 1793 0 1 5387
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_535
timestamp 1626065694
transform 1 0 1793 0 1 5723
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_534
timestamp 1626065694
transform 1 0 1793 0 1 6059
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_533
timestamp 1626065694
transform 1 0 1793 0 1 6395
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_532
timestamp 1626065694
transform 1 0 1793 0 1 6731
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_531
timestamp 1626065694
transform 1 0 1793 0 1 7067
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_530
timestamp 1626065694
transform 1 0 1793 0 1 7403
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_529
timestamp 1626065694
transform 1 0 1793 0 1 7739
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_528
timestamp 1626065694
transform 1 0 1793 0 1 8075
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_527
timestamp 1626065694
transform 1 0 1793 0 1 8411
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_526
timestamp 1626065694
transform 1 0 1793 0 1 8747
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_525
timestamp 1626065694
transform 1 0 1793 0 1 9083
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_524
timestamp 1626065694
transform 1 0 1793 0 1 9419
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_523
timestamp 1626065694
transform 1 0 1793 0 1 9755
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_522
timestamp 1626065694
transform 1 0 1793 0 1 10091
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_521
timestamp 1626065694
transform 1 0 1793 0 1 10427
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_520
timestamp 1626065694
transform 1 0 4481 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_519
timestamp 1626065694
transform 1 0 1793 0 1 4379
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_518
timestamp 1626065694
transform 1 0 1793 0 1 4715
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_517
timestamp 1626065694
transform 1 0 1793 0 1 5051
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_516
timestamp 1626065694
transform 1 0 1793 0 1 3035
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_515
timestamp 1626065694
transform 1 0 1793 0 1 3371
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_514
timestamp 1626065694
transform 1 0 1793 0 1 3707
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_513
timestamp 1626065694
transform 1 0 1793 0 1 4043
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_512
timestamp 1626065694
transform 1 0 1793 0 1 2027
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_511
timestamp 1626065694
transform 1 0 1793 0 1 2363
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_510
timestamp 1626065694
transform 1 0 1793 0 1 2699
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_509
timestamp 1626065694
transform 1 0 2129 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_508
timestamp 1626065694
transform 1 0 2465 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_507
timestamp 1626065694
transform 1 0 2801 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_506
timestamp 1626065694
transform 1 0 3137 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_505
timestamp 1626065694
transform 1 0 3473 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_504
timestamp 1626065694
transform 1 0 3809 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_503
timestamp 1626065694
transform 1 0 4145 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_502
timestamp 1626065694
transform 1 0 7505 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_501
timestamp 1626065694
transform 1 0 8177 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_500
timestamp 1626065694
transform 1 0 5825 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_499
timestamp 1626065694
transform 1 0 6161 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_498
timestamp 1626065694
transform 1 0 6497 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_497
timestamp 1626065694
transform 1 0 6833 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_496
timestamp 1626065694
transform 1 0 5489 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_495
timestamp 1626065694
transform 1 0 8513 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_494
timestamp 1626065694
transform 1 0 7169 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_493
timestamp 1626065694
transform 1 0 4817 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_492
timestamp 1626065694
transform 1 0 7841 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_491
timestamp 1626065694
transform 1 0 5153 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_490
timestamp 1626065694
transform 1 0 13889 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_489
timestamp 1626065694
transform 1 0 14225 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_488
timestamp 1626065694
transform 1 0 14561 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_487
timestamp 1626065694
transform 1 0 14897 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_486
timestamp 1626065694
transform 1 0 15233 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_485
timestamp 1626065694
transform 1 0 15569 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_484
timestamp 1626065694
transform 1 0 15905 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_483
timestamp 1626065694
transform 1 0 16241 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_482
timestamp 1626065694
transform 1 0 16577 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_481
timestamp 1626065694
transform 1 0 16913 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_480
timestamp 1626065694
transform 1 0 10529 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_479
timestamp 1626065694
transform 1 0 10865 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_478
timestamp 1626065694
transform 1 0 11201 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_477
timestamp 1626065694
transform 1 0 11537 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_476
timestamp 1626065694
transform 1 0 9857 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_475
timestamp 1626065694
transform 1 0 9185 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_474
timestamp 1626065694
transform 1 0 11873 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_473
timestamp 1626065694
transform 1 0 12209 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_472
timestamp 1626065694
transform 1 0 12545 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_471
timestamp 1626065694
transform 1 0 12881 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_470
timestamp 1626065694
transform 1 0 13217 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_469
timestamp 1626065694
transform 1 0 10193 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_468
timestamp 1626065694
transform 1 0 13553 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_467
timestamp 1626065694
transform 1 0 8849 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_466
timestamp 1626065694
transform 1 0 9521 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_465
timestamp 1626065694
transform 1 0 20945 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_464
timestamp 1626065694
transform 1 0 18929 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_463
timestamp 1626065694
transform 1 0 21281 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_462
timestamp 1626065694
transform 1 0 21617 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_461
timestamp 1626065694
transform 1 0 21953 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_460
timestamp 1626065694
transform 1 0 17585 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_459
timestamp 1626065694
transform 1 0 22289 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_458
timestamp 1626065694
transform 1 0 19265 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_457
timestamp 1626065694
transform 1 0 22625 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_456
timestamp 1626065694
transform 1 0 19601 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_455
timestamp 1626065694
transform 1 0 22961 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_454
timestamp 1626065694
transform 1 0 23297 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_453
timestamp 1626065694
transform 1 0 23633 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_452
timestamp 1626065694
transform 1 0 23969 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_451
timestamp 1626065694
transform 1 0 24305 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_450
timestamp 1626065694
transform 1 0 24641 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_449
timestamp 1626065694
transform 1 0 24977 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_448
timestamp 1626065694
transform 1 0 25313 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_447
timestamp 1626065694
transform 1 0 25649 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_446
timestamp 1626065694
transform 1 0 19937 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_445
timestamp 1626065694
transform 1 0 20273 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_444
timestamp 1626065694
transform 1 0 20609 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_443
timestamp 1626065694
transform 1 0 17921 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_442
timestamp 1626065694
transform 1 0 18593 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_441
timestamp 1626065694
transform 1 0 18257 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_440
timestamp 1626065694
transform 1 0 33041 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_439
timestamp 1626065694
transform 1 0 29009 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_438
timestamp 1626065694
transform 1 0 33377 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_437
timestamp 1626065694
transform 1 0 33713 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_436
timestamp 1626065694
transform 1 0 34049 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_435
timestamp 1626065694
transform 1 0 29345 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_434
timestamp 1626065694
transform 1 0 29681 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_433
timestamp 1626065694
transform 1 0 30017 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_432
timestamp 1626065694
transform 1 0 25985 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_431
timestamp 1626065694
transform 1 0 30353 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_430
timestamp 1626065694
transform 1 0 30689 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_429
timestamp 1626065694
transform 1 0 26321 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_428
timestamp 1626065694
transform 1 0 31025 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_427
timestamp 1626065694
transform 1 0 26657 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_426
timestamp 1626065694
transform 1 0 31361 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_425
timestamp 1626065694
transform 1 0 31697 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_424
timestamp 1626065694
transform 1 0 26993 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_423
timestamp 1626065694
transform 1 0 27329 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_422
timestamp 1626065694
transform 1 0 32033 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_421
timestamp 1626065694
transform 1 0 28337 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_420
timestamp 1626065694
transform 1 0 32369 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_419
timestamp 1626065694
transform 1 0 32705 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_418
timestamp 1626065694
transform 1 0 28673 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_417
timestamp 1626065694
transform 1 0 27665 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_416
timestamp 1626065694
transform 1 0 28001 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_415
timestamp 1626065694
transform 1 0 42785 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_414
timestamp 1626065694
transform 1 0 39761 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_413
timestamp 1626065694
transform 1 0 40097 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_412
timestamp 1626065694
transform 1 0 40433 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_411
timestamp 1626065694
transform 1 0 40769 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_410
timestamp 1626065694
transform 1 0 41105 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_409
timestamp 1626065694
transform 1 0 41441 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_408
timestamp 1626065694
transform 1 0 41777 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_407
timestamp 1626065694
transform 1 0 42113 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_406
timestamp 1626065694
transform 1 0 42449 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_405
timestamp 1626065694
transform 1 0 39425 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_404
timestamp 1626065694
transform 1 0 34385 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_403
timestamp 1626065694
transform 1 0 34721 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_402
timestamp 1626065694
transform 1 0 35057 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_401
timestamp 1626065694
transform 1 0 35393 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_400
timestamp 1626065694
transform 1 0 35729 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_399
timestamp 1626065694
transform 1 0 36065 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_398
timestamp 1626065694
transform 1 0 36401 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_397
timestamp 1626065694
transform 1 0 36737 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_396
timestamp 1626065694
transform 1 0 37073 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_395
timestamp 1626065694
transform 1 0 37409 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_394
timestamp 1626065694
transform 1 0 37745 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_393
timestamp 1626065694
transform 1 0 38081 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_392
timestamp 1626065694
transform 1 0 38417 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_391
timestamp 1626065694
transform 1 0 38753 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_390
timestamp 1626065694
transform 1 0 39089 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_389
timestamp 1626065694
transform 1 0 48161 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_388
timestamp 1626065694
transform 1 0 48497 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_387
timestamp 1626065694
transform 1 0 48833 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_386
timestamp 1626065694
transform 1 0 49169 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_385
timestamp 1626065694
transform 1 0 49505 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_384
timestamp 1626065694
transform 1 0 44465 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_383
timestamp 1626065694
transform 1 0 44801 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_382
timestamp 1626065694
transform 1 0 49841 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_381
timestamp 1626065694
transform 1 0 50177 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_380
timestamp 1626065694
transform 1 0 50513 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_379
timestamp 1626065694
transform 1 0 50849 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_378
timestamp 1626065694
transform 1 0 45137 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_377
timestamp 1626065694
transform 1 0 45473 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_376
timestamp 1626065694
transform 1 0 45809 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_375
timestamp 1626065694
transform 1 0 51185 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_374
timestamp 1626065694
transform 1 0 46145 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_373
timestamp 1626065694
transform 1 0 43121 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_372
timestamp 1626065694
transform 1 0 43457 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_371
timestamp 1626065694
transform 1 0 46481 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_370
timestamp 1626065694
transform 1 0 46817 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_369
timestamp 1626065694
transform 1 0 47153 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_368
timestamp 1626065694
transform 1 0 47489 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_367
timestamp 1626065694
transform 1 0 43793 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_366
timestamp 1626065694
transform 1 0 44129 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_365
timestamp 1626065694
transform 1 0 47825 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_364
timestamp 1626065694
transform 1 0 58241 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_363
timestamp 1626065694
transform 1 0 58577 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_362
timestamp 1626065694
transform 1 0 57905 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_361
timestamp 1626065694
transform 1 0 51521 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_360
timestamp 1626065694
transform 1 0 51857 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_359
timestamp 1626065694
transform 1 0 52193 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_358
timestamp 1626065694
transform 1 0 52529 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_357
timestamp 1626065694
transform 1 0 52865 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_356
timestamp 1626065694
transform 1 0 53201 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_355
timestamp 1626065694
transform 1 0 53537 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_354
timestamp 1626065694
transform 1 0 53873 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_353
timestamp 1626065694
transform 1 0 54209 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_352
timestamp 1626065694
transform 1 0 54545 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_351
timestamp 1626065694
transform 1 0 54881 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_350
timestamp 1626065694
transform 1 0 59585 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_349
timestamp 1626065694
transform 1 0 57569 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_348
timestamp 1626065694
transform 1 0 55217 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_347
timestamp 1626065694
transform 1 0 59249 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_346
timestamp 1626065694
transform 1 0 55553 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_345
timestamp 1626065694
transform 1 0 55889 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_344
timestamp 1626065694
transform 1 0 56225 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_343
timestamp 1626065694
transform 1 0 56561 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_342
timestamp 1626065694
transform 1 0 56897 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_341
timestamp 1626065694
transform 1 0 58913 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_340
timestamp 1626065694
transform 1 0 57233 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_339
timestamp 1626065694
transform 1 0 63281 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_338
timestamp 1626065694
transform 1 0 60929 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_337
timestamp 1626065694
transform 1 0 62273 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_336
timestamp 1626065694
transform 1 0 66305 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_335
timestamp 1626065694
transform 1 0 65633 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_334
timestamp 1626065694
transform 1 0 66641 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_333
timestamp 1626065694
transform 1 0 66977 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_332
timestamp 1626065694
transform 1 0 65969 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_331
timestamp 1626065694
transform 1 0 64961 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_330
timestamp 1626065694
transform 1 0 67985 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_329
timestamp 1626065694
transform 1 0 67313 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_328
timestamp 1626065694
transform 1 0 64289 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_327
timestamp 1626065694
transform 1 0 60257 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_326
timestamp 1626065694
transform 1 0 61265 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_325
timestamp 1626065694
transform 1 0 67649 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_324
timestamp 1626065694
transform 1 0 59921 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_323
timestamp 1626065694
transform 1 0 63617 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_322
timestamp 1626065694
transform 1 0 62609 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_321
timestamp 1626065694
transform 1 0 61937 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_320
timestamp 1626065694
transform 1 0 61601 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_319
timestamp 1626065694
transform 1 0 60593 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_318
timestamp 1626065694
transform 1 0 62945 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_317
timestamp 1626065694
transform 1 0 65297 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_316
timestamp 1626065694
transform 1 0 64625 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_315
timestamp 1626065694
transform 1 0 63953 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_314
timestamp 1626065694
transform 1 0 134843 0 1 31259
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_313
timestamp 1626065694
transform 1 0 134843 0 1 36635
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_312
timestamp 1626065694
transform 1 0 134843 0 1 36971
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_311
timestamp 1626065694
transform 1 0 134843 0 1 37307
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_310
timestamp 1626065694
transform 1 0 134843 0 1 37643
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_309
timestamp 1626065694
transform 1 0 134843 0 1 37979
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_308
timestamp 1626065694
transform 1 0 134843 0 1 38315
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_307
timestamp 1626065694
transform 1 0 134843 0 1 38651
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_306
timestamp 1626065694
transform 1 0 134843 0 1 38987
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_305
timestamp 1626065694
transform 1 0 134843 0 1 39323
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_304
timestamp 1626065694
transform 1 0 134843 0 1 39659
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_303
timestamp 1626065694
transform 1 0 134843 0 1 39995
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_302
timestamp 1626065694
transform 1 0 134843 0 1 40331
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_301
timestamp 1626065694
transform 1 0 134843 0 1 40667
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_300
timestamp 1626065694
transform 1 0 134843 0 1 41003
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_299
timestamp 1626065694
transform 1 0 134843 0 1 41339
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_298
timestamp 1626065694
transform 1 0 134843 0 1 31931
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_297
timestamp 1626065694
transform 1 0 134843 0 1 32267
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_296
timestamp 1626065694
transform 1 0 134843 0 1 32603
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_295
timestamp 1626065694
transform 1 0 134843 0 1 32939
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_294
timestamp 1626065694
transform 1 0 134843 0 1 33275
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_293
timestamp 1626065694
transform 1 0 134843 0 1 33611
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_292
timestamp 1626065694
transform 1 0 134843 0 1 33947
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_291
timestamp 1626065694
transform 1 0 134843 0 1 34283
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_290
timestamp 1626065694
transform 1 0 134843 0 1 34619
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_289
timestamp 1626065694
transform 1 0 134843 0 1 34955
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_288
timestamp 1626065694
transform 1 0 134843 0 1 35291
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_287
timestamp 1626065694
transform 1 0 134843 0 1 35627
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_286
timestamp 1626065694
transform 1 0 134843 0 1 35963
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_285
timestamp 1626065694
transform 1 0 134843 0 1 36299
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_284
timestamp 1626065694
transform 1 0 134843 0 1 31595
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_283
timestamp 1626065694
transform 1 0 134843 0 1 27563
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_282
timestamp 1626065694
transform 1 0 134843 0 1 27899
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_281
timestamp 1626065694
transform 1 0 134843 0 1 28235
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_280
timestamp 1626065694
transform 1 0 134843 0 1 28571
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_279
timestamp 1626065694
transform 1 0 134843 0 1 28907
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_278
timestamp 1626065694
transform 1 0 134843 0 1 29243
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_277
timestamp 1626065694
transform 1 0 134843 0 1 29579
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_276
timestamp 1626065694
transform 1 0 134843 0 1 29915
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_275
timestamp 1626065694
transform 1 0 134843 0 1 30251
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_274
timestamp 1626065694
transform 1 0 134843 0 1 30587
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_273
timestamp 1626065694
transform 1 0 134843 0 1 30923
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_272
timestamp 1626065694
transform 1 0 134843 0 1 26219
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_271
timestamp 1626065694
transform 1 0 134843 0 1 26555
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_270
timestamp 1626065694
transform 1 0 134843 0 1 26891
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_269
timestamp 1626065694
transform 1 0 134843 0 1 27227
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_268
timestamp 1626065694
transform 1 0 134843 0 1 21515
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_267
timestamp 1626065694
transform 1 0 134843 0 1 22859
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_266
timestamp 1626065694
transform 1 0 134843 0 1 21851
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_265
timestamp 1626065694
transform 1 0 134843 0 1 22187
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_264
timestamp 1626065694
transform 1 0 134843 0 1 23195
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_263
timestamp 1626065694
transform 1 0 134843 0 1 25211
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_262
timestamp 1626065694
transform 1 0 134843 0 1 25547
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_261
timestamp 1626065694
transform 1 0 134843 0 1 25883
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_260
timestamp 1626065694
transform 1 0 134843 0 1 23531
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_259
timestamp 1626065694
transform 1 0 134843 0 1 23867
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_258
timestamp 1626065694
transform 1 0 134843 0 1 24203
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_257
timestamp 1626065694
transform 1 0 134843 0 1 24539
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_256
timestamp 1626065694
transform 1 0 134843 0 1 24875
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_255
timestamp 1626065694
transform 1 0 134843 0 1 22523
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_254
timestamp 1626065694
transform 1 0 134843 0 1 21179
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_253
timestamp 1626065694
transform 1 0 75377 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_252
timestamp 1626065694
transform 1 0 68321 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_251
timestamp 1626065694
transform 1 0 68657 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_250
timestamp 1626065694
transform 1 0 68993 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_249
timestamp 1626065694
transform 1 0 69329 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_248
timestamp 1626065694
transform 1 0 69665 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_247
timestamp 1626065694
transform 1 0 70001 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_246
timestamp 1626065694
transform 1 0 70337 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_245
timestamp 1626065694
transform 1 0 70673 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_244
timestamp 1626065694
transform 1 0 71009 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_243
timestamp 1626065694
transform 1 0 71345 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_242
timestamp 1626065694
transform 1 0 71681 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_241
timestamp 1626065694
transform 1 0 72017 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_240
timestamp 1626065694
transform 1 0 72353 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_239
timestamp 1626065694
transform 1 0 72689 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_238
timestamp 1626065694
transform 1 0 73025 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_237
timestamp 1626065694
transform 1 0 73361 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_236
timestamp 1626065694
transform 1 0 73697 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_235
timestamp 1626065694
transform 1 0 74033 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_234
timestamp 1626065694
transform 1 0 76385 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_233
timestamp 1626065694
transform 1 0 76721 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_232
timestamp 1626065694
transform 1 0 75713 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_231
timestamp 1626065694
transform 1 0 76049 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_230
timestamp 1626065694
transform 1 0 74369 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_229
timestamp 1626065694
transform 1 0 74705 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_228
timestamp 1626065694
transform 1 0 75041 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_227
timestamp 1626065694
transform 1 0 80417 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_226
timestamp 1626065694
transform 1 0 83105 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_225
timestamp 1626065694
transform 1 0 80753 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_224
timestamp 1626065694
transform 1 0 81089 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_223
timestamp 1626065694
transform 1 0 82433 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_222
timestamp 1626065694
transform 1 0 83777 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_221
timestamp 1626065694
transform 1 0 81425 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_220
timestamp 1626065694
transform 1 0 77393 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_219
timestamp 1626065694
transform 1 0 77057 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_218
timestamp 1626065694
transform 1 0 84113 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_217
timestamp 1626065694
transform 1 0 78065 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_216
timestamp 1626065694
transform 1 0 84449 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_215
timestamp 1626065694
transform 1 0 82769 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_214
timestamp 1626065694
transform 1 0 81761 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_213
timestamp 1626065694
transform 1 0 82097 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_212
timestamp 1626065694
transform 1 0 77729 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_211
timestamp 1626065694
transform 1 0 79745 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_210
timestamp 1626065694
transform 1 0 83441 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_209
timestamp 1626065694
transform 1 0 78737 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_208
timestamp 1626065694
transform 1 0 84785 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_207
timestamp 1626065694
transform 1 0 85121 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_206
timestamp 1626065694
transform 1 0 78401 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_205
timestamp 1626065694
transform 1 0 79073 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_204
timestamp 1626065694
transform 1 0 80081 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_203
timestamp 1626065694
transform 1 0 79409 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_202
timestamp 1626065694
transform 1 0 86801 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_201
timestamp 1626065694
transform 1 0 87137 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_200
timestamp 1626065694
transform 1 0 87473 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_199
timestamp 1626065694
transform 1 0 87809 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_198
timestamp 1626065694
transform 1 0 90161 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_197
timestamp 1626065694
transform 1 0 90497 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_196
timestamp 1626065694
transform 1 0 93185 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_195
timestamp 1626065694
transform 1 0 90833 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_194
timestamp 1626065694
transform 1 0 88145 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_193
timestamp 1626065694
transform 1 0 91169 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_192
timestamp 1626065694
transform 1 0 88481 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_191
timestamp 1626065694
transform 1 0 88817 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_190
timestamp 1626065694
transform 1 0 93521 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_189
timestamp 1626065694
transform 1 0 86465 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_188
timestamp 1626065694
transform 1 0 89153 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_187
timestamp 1626065694
transform 1 0 89489 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_186
timestamp 1626065694
transform 1 0 91505 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_185
timestamp 1626065694
transform 1 0 89825 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_184
timestamp 1626065694
transform 1 0 92513 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_183
timestamp 1626065694
transform 1 0 91841 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_182
timestamp 1626065694
transform 1 0 92849 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_181
timestamp 1626065694
transform 1 0 85457 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_180
timestamp 1626065694
transform 1 0 92177 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_179
timestamp 1626065694
transform 1 0 85793 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_178
timestamp 1626065694
transform 1 0 86129 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_177
timestamp 1626065694
transform 1 0 99569 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_176
timestamp 1626065694
transform 1 0 102257 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_175
timestamp 1626065694
transform 1 0 94865 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_174
timestamp 1626065694
transform 1 0 98225 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_173
timestamp 1626065694
transform 1 0 98561 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_172
timestamp 1626065694
transform 1 0 95201 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_171
timestamp 1626065694
transform 1 0 95537 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_170
timestamp 1626065694
transform 1 0 99905 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_169
timestamp 1626065694
transform 1 0 95873 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_168
timestamp 1626065694
transform 1 0 96209 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_167
timestamp 1626065694
transform 1 0 100241 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_166
timestamp 1626065694
transform 1 0 100577 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_165
timestamp 1626065694
transform 1 0 98897 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_164
timestamp 1626065694
transform 1 0 100913 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_163
timestamp 1626065694
transform 1 0 101249 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_162
timestamp 1626065694
transform 1 0 93857 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_161
timestamp 1626065694
transform 1 0 99233 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_160
timestamp 1626065694
transform 1 0 94193 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_159
timestamp 1626065694
transform 1 0 96545 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_158
timestamp 1626065694
transform 1 0 101585 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_157
timestamp 1626065694
transform 1 0 101921 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_156
timestamp 1626065694
transform 1 0 94529 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_155
timestamp 1626065694
transform 1 0 96881 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_154
timestamp 1626065694
transform 1 0 97217 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_153
timestamp 1626065694
transform 1 0 97553 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_152
timestamp 1626065694
transform 1 0 97889 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_151
timestamp 1626065694
transform 1 0 134843 0 1 15803
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_150
timestamp 1626065694
transform 1 0 134843 0 1 16139
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_149
timestamp 1626065694
transform 1 0 134843 0 1 16475
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_148
timestamp 1626065694
transform 1 0 134843 0 1 16811
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_147
timestamp 1626065694
transform 1 0 134843 0 1 17147
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_146
timestamp 1626065694
transform 1 0 134843 0 1 17483
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_145
timestamp 1626065694
transform 1 0 134843 0 1 17819
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_144
timestamp 1626065694
transform 1 0 134843 0 1 18155
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_143
timestamp 1626065694
transform 1 0 134843 0 1 18491
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_142
timestamp 1626065694
transform 1 0 134843 0 1 18827
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_141
timestamp 1626065694
transform 1 0 134843 0 1 19163
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_140
timestamp 1626065694
transform 1 0 134843 0 1 19499
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_139
timestamp 1626065694
transform 1 0 134843 0 1 19835
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_138
timestamp 1626065694
transform 1 0 134843 0 1 20171
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_137
timestamp 1626065694
transform 1 0 134843 0 1 20507
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_136
timestamp 1626065694
transform 1 0 134843 0 1 20843
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_135
timestamp 1626065694
transform 1 0 134843 0 1 15467
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_134
timestamp 1626065694
transform 1 0 134843 0 1 10763
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_133
timestamp 1626065694
transform 1 0 134843 0 1 11099
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_132
timestamp 1626065694
transform 1 0 134843 0 1 11435
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_131
timestamp 1626065694
transform 1 0 134843 0 1 11771
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_130
timestamp 1626065694
transform 1 0 134843 0 1 12107
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_129
timestamp 1626065694
transform 1 0 134843 0 1 12443
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_128
timestamp 1626065694
transform 1 0 134843 0 1 12779
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_127
timestamp 1626065694
transform 1 0 134843 0 1 13115
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_126
timestamp 1626065694
transform 1 0 134843 0 1 13451
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_125
timestamp 1626065694
transform 1 0 134843 0 1 13787
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_124
timestamp 1626065694
transform 1 0 134843 0 1 14123
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_123
timestamp 1626065694
transform 1 0 134843 0 1 14459
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_122
timestamp 1626065694
transform 1 0 134843 0 1 14795
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_121
timestamp 1626065694
transform 1 0 134843 0 1 15131
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_120
timestamp 1626065694
transform 1 0 109313 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_119
timestamp 1626065694
transform 1 0 109649 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_118
timestamp 1626065694
transform 1 0 106289 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_117
timestamp 1626065694
transform 1 0 109985 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_116
timestamp 1626065694
transform 1 0 107969 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_115
timestamp 1626065694
transform 1 0 110321 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_114
timestamp 1626065694
transform 1 0 110657 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_113
timestamp 1626065694
transform 1 0 106625 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_112
timestamp 1626065694
transform 1 0 106961 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_111
timestamp 1626065694
transform 1 0 104945 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_110
timestamp 1626065694
transform 1 0 105281 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_109
timestamp 1626065694
transform 1 0 102593 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_108
timestamp 1626065694
transform 1 0 102929 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_107
timestamp 1626065694
transform 1 0 103265 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_106
timestamp 1626065694
transform 1 0 104609 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_105
timestamp 1626065694
transform 1 0 103601 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_104
timestamp 1626065694
transform 1 0 103937 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_103
timestamp 1626065694
transform 1 0 107297 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_102
timestamp 1626065694
transform 1 0 105617 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_101
timestamp 1626065694
transform 1 0 108305 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_100
timestamp 1626065694
transform 1 0 107633 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_99
timestamp 1626065694
transform 1 0 108641 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_98
timestamp 1626065694
transform 1 0 105953 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_97
timestamp 1626065694
transform 1 0 108977 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_96
timestamp 1626065694
transform 1 0 104273 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_95
timestamp 1626065694
transform 1 0 117713 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_94
timestamp 1626065694
transform 1 0 115361 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_93
timestamp 1626065694
transform 1 0 112001 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_92
timestamp 1626065694
transform 1 0 118049 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_91
timestamp 1626065694
transform 1 0 112337 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_90
timestamp 1626065694
transform 1 0 112673 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_89
timestamp 1626065694
transform 1 0 113009 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_88
timestamp 1626065694
transform 1 0 116033 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_87
timestamp 1626065694
transform 1 0 113345 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_86
timestamp 1626065694
transform 1 0 118385 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_85
timestamp 1626065694
transform 1 0 116705 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_84
timestamp 1626065694
transform 1 0 116369 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_83
timestamp 1626065694
transform 1 0 117041 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_82
timestamp 1626065694
transform 1 0 113681 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_81
timestamp 1626065694
transform 1 0 118721 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_80
timestamp 1626065694
transform 1 0 119057 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_79
timestamp 1626065694
transform 1 0 110993 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_78
timestamp 1626065694
transform 1 0 114017 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_77
timestamp 1626065694
transform 1 0 115697 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_76
timestamp 1626065694
transform 1 0 111329 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_75
timestamp 1626065694
transform 1 0 117377 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_74
timestamp 1626065694
transform 1 0 114353 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_73
timestamp 1626065694
transform 1 0 114689 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_72
timestamp 1626065694
transform 1 0 111665 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_71
timestamp 1626065694
transform 1 0 115025 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_70
timestamp 1626065694
transform 1 0 127793 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_69
timestamp 1626065694
transform 1 0 134843 0 1 5387
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_68
timestamp 1626065694
transform 1 0 134843 0 1 5723
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_67
timestamp 1626065694
transform 1 0 134843 0 1 6059
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_66
timestamp 1626065694
transform 1 0 134843 0 1 6395
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_65
timestamp 1626065694
transform 1 0 134843 0 1 6731
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_64
timestamp 1626065694
transform 1 0 134843 0 1 7067
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_63
timestamp 1626065694
transform 1 0 134843 0 1 7403
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_62
timestamp 1626065694
transform 1 0 134843 0 1 7739
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_61
timestamp 1626065694
transform 1 0 134843 0 1 8075
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_60
timestamp 1626065694
transform 1 0 134843 0 1 8411
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_59
timestamp 1626065694
transform 1 0 134843 0 1 8747
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_58
timestamp 1626065694
transform 1 0 134843 0 1 9083
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_57
timestamp 1626065694
transform 1 0 134843 0 1 9419
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_56
timestamp 1626065694
transform 1 0 134843 0 1 9755
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_55
timestamp 1626065694
transform 1 0 134843 0 1 10091
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_54
timestamp 1626065694
transform 1 0 134843 0 1 10427
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_53
timestamp 1626065694
transform 1 0 126785 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_52
timestamp 1626065694
transform 1 0 127121 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_51
timestamp 1626065694
transform 1 0 127457 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_50
timestamp 1626065694
transform 1 0 119393 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_49
timestamp 1626065694
transform 1 0 119729 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_48
timestamp 1626065694
transform 1 0 120065 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_47
timestamp 1626065694
transform 1 0 120401 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_46
timestamp 1626065694
transform 1 0 120737 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_45
timestamp 1626065694
transform 1 0 121073 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_44
timestamp 1626065694
transform 1 0 121409 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_43
timestamp 1626065694
transform 1 0 121745 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_42
timestamp 1626065694
transform 1 0 122081 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_41
timestamp 1626065694
transform 1 0 122417 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_40
timestamp 1626065694
transform 1 0 122753 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_39
timestamp 1626065694
transform 1 0 123089 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_38
timestamp 1626065694
transform 1 0 123425 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_37
timestamp 1626065694
transform 1 0 123761 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_36
timestamp 1626065694
transform 1 0 124097 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_35
timestamp 1626065694
transform 1 0 124433 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_34
timestamp 1626065694
transform 1 0 124769 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_33
timestamp 1626065694
transform 1 0 125105 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_32
timestamp 1626065694
transform 1 0 125441 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_31
timestamp 1626065694
transform 1 0 125777 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_30
timestamp 1626065694
transform 1 0 126113 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_29
timestamp 1626065694
transform 1 0 126449 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_28
timestamp 1626065694
transform 1 0 134843 0 1 4379
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_27
timestamp 1626065694
transform 1 0 134843 0 1 4715
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_26
timestamp 1626065694
transform 1 0 134843 0 1 5051
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_25
timestamp 1626065694
transform 1 0 134843 0 1 3371
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_24
timestamp 1626065694
transform 1 0 134843 0 1 4043
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_23
timestamp 1626065694
transform 1 0 134843 0 1 3707
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_22
timestamp 1626065694
transform 1 0 134843 0 1 3035
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_21
timestamp 1626065694
transform 1 0 128465 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_20
timestamp 1626065694
transform 1 0 128801 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_19
timestamp 1626065694
transform 1 0 129137 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_18
timestamp 1626065694
transform 1 0 129473 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_17
timestamp 1626065694
transform 1 0 129809 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_16
timestamp 1626065694
transform 1 0 130145 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_15
timestamp 1626065694
transform 1 0 130481 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_14
timestamp 1626065694
transform 1 0 130817 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_13
timestamp 1626065694
transform 1 0 131153 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_12
timestamp 1626065694
transform 1 0 131489 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_11
timestamp 1626065694
transform 1 0 131825 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_10
timestamp 1626065694
transform 1 0 128129 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_9
timestamp 1626065694
transform 1 0 133169 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_8
timestamp 1626065694
transform 1 0 133505 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_7
timestamp 1626065694
transform 1 0 134843 0 1 2027
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_6
timestamp 1626065694
transform 1 0 133841 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_5
timestamp 1626065694
transform 1 0 134177 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_4
timestamp 1626065694
transform 1 0 132161 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_3
timestamp 1626065694
transform 1 0 132497 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_2
timestamp 1626065694
transform 1 0 132833 0 1 1691
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1
timestamp 1626065694
transform 1 0 134843 0 1 2363
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_0
timestamp 1626065694
transform 1 0 134843 0 1 2699
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3615
timestamp 1626065694
transform 1 0 68272 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3614
timestamp 1626065694
transform 1 0 21216 0 1 41621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3613
timestamp 1626065694
transform 1 0 21624 0 1 41621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3612
timestamp 1626065694
transform 1 0 22440 0 1 41621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3611
timestamp 1626065694
transform 1 0 114376 0 1 41621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3610
timestamp 1626065694
transform 1 0 115192 0 1 41621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3609
timestamp 1626065694
transform 1 0 115328 0 1 41621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3608
timestamp 1626065694
transform 1 0 20808 0 1 41621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3607
timestamp 1626065694
transform 1 0 22032 0 1 41621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3606
timestamp 1626065694
transform 1 0 114784 0 1 41621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3605
timestamp 1626065694
transform 1 0 115872 0 1 41621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3604
timestamp 1626065694
transform 1 0 109344 0 1 62293
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3603
timestamp 1626065694
transform 1 0 133144 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3602
timestamp 1626065694
transform 1 0 133144 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3601
timestamp 1626065694
transform 1 0 135320 0 1 80925
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3600
timestamp 1626065694
transform 1 0 128112 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3599
timestamp 1626065694
transform 1 0 128112 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3598
timestamp 1626065694
transform 1 0 129880 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3597
timestamp 1626065694
transform 1 0 129880 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3596
timestamp 1626065694
transform 1 0 131376 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3595
timestamp 1626065694
transform 1 0 131376 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3594
timestamp 1626065694
transform 1 0 130832 0 1 79157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3593
timestamp 1626065694
transform 1 0 134776 0 1 78341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3592
timestamp 1626065694
transform 1 0 135320 0 1 79429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3591
timestamp 1626065694
transform 1 0 136000 0 1 79837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3590
timestamp 1626065694
transform 1 0 119680 0 1 80245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3589
timestamp 1626065694
transform 1 0 119544 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3588
timestamp 1626065694
transform 1 0 119544 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3587
timestamp 1626065694
transform 1 0 121448 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3586
timestamp 1626065694
transform 1 0 121448 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3585
timestamp 1626065694
transform 1 0 122264 0 1 78341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3584
timestamp 1626065694
transform 1 0 122944 0 1 78477
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3583
timestamp 1626065694
transform 1 0 122944 0 1 81333
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3582
timestamp 1626065694
transform 1 0 123216 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3581
timestamp 1626065694
transform 1 0 123216 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3580
timestamp 1626065694
transform 1 0 124712 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3579
timestamp 1626065694
transform 1 0 124712 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3578
timestamp 1626065694
transform 1 0 126344 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3577
timestamp 1626065694
transform 1 0 126344 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3576
timestamp 1626065694
transform 1 0 122264 0 1 80653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3575
timestamp 1626065694
transform 1 0 122264 0 1 79837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3574
timestamp 1626065694
transform 1 0 122400 0 1 79701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3573
timestamp 1626065694
transform 1 0 122264 0 1 72765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3572
timestamp 1626065694
transform 1 0 122264 0 1 75485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3571
timestamp 1626065694
transform 1 0 122400 0 1 74261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3570
timestamp 1626065694
transform 1 0 122400 0 1 76845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3569
timestamp 1626065694
transform 1 0 122400 0 1 73989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3568
timestamp 1626065694
transform 1 0 122400 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3567
timestamp 1626065694
transform 1 0 122264 0 1 75621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3566
timestamp 1626065694
transform 1 0 134776 0 1 77661
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3565
timestamp 1626065694
transform 1 0 135320 0 1 76029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3564
timestamp 1626065694
transform 1 0 135320 0 1 77661
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3563
timestamp 1626065694
transform 1 0 135320 0 1 74125
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3562
timestamp 1626065694
transform 1 0 136000 0 1 72765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3561
timestamp 1626065694
transform 1 0 118456 0 1 80245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3560
timestamp 1626065694
transform 1 0 111384 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3559
timestamp 1626065694
transform 1 0 111384 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3558
timestamp 1626065694
transform 1 0 112880 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3557
timestamp 1626065694
transform 1 0 112880 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3556
timestamp 1626065694
transform 1 0 114648 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3555
timestamp 1626065694
transform 1 0 114648 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3554
timestamp 1626065694
transform 1 0 116416 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3553
timestamp 1626065694
transform 1 0 116416 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3552
timestamp 1626065694
transform 1 0 118048 0 1 79293
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3551
timestamp 1626065694
transform 1 0 118184 0 1 81333
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3550
timestamp 1626065694
transform 1 0 118184 0 1 79429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3549
timestamp 1626065694
transform 1 0 117912 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3548
timestamp 1626065694
transform 1 0 117912 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3547
timestamp 1626065694
transform 1 0 116552 0 1 78477
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3546
timestamp 1626065694
transform 1 0 117912 0 1 78613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3545
timestamp 1626065694
transform 1 0 117912 0 1 80653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3544
timestamp 1626065694
transform 1 0 118048 0 1 80789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3543
timestamp 1626065694
transform 1 0 118048 0 1 82693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3542
timestamp 1626065694
transform 1 0 102952 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3541
timestamp 1626065694
transform 1 0 102952 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3540
timestamp 1626065694
transform 1 0 104584 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3539
timestamp 1626065694
transform 1 0 104584 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3538
timestamp 1626065694
transform 1 0 106352 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3537
timestamp 1626065694
transform 1 0 106352 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3536
timestamp 1626065694
transform 1 0 107848 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3535
timestamp 1626065694
transform 1 0 107848 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3534
timestamp 1626065694
transform 1 0 109616 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3533
timestamp 1626065694
transform 1 0 109616 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3532
timestamp 1626065694
transform 1 0 106352 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3531
timestamp 1626065694
transform 1 0 106352 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3530
timestamp 1626065694
transform 1 0 106352 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3529
timestamp 1626065694
transform 1 0 109616 0 1 73037
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3528
timestamp 1626065694
transform 1 0 103360 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3527
timestamp 1626065694
transform 1 0 103768 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3526
timestamp 1626065694
transform 1 0 103768 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3525
timestamp 1626065694
transform 1 0 106080 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3524
timestamp 1626065694
transform 1 0 106216 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3523
timestamp 1626065694
transform 1 0 106216 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3522
timestamp 1626065694
transform 1 0 103904 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3521
timestamp 1626065694
transform 1 0 103904 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3520
timestamp 1626065694
transform 1 0 103904 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3519
timestamp 1626065694
transform 1 0 103904 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3518
timestamp 1626065694
transform 1 0 106352 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3517
timestamp 1626065694
transform 1 0 115328 0 1 74261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3516
timestamp 1626065694
transform 1 0 115328 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3515
timestamp 1626065694
transform 1 0 116552 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3514
timestamp 1626065694
transform 1 0 118048 0 1 77253
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3513
timestamp 1626065694
transform 1 0 115328 0 1 74397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3512
timestamp 1626065694
transform 1 0 115464 0 1 75621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3511
timestamp 1626065694
transform 1 0 115464 0 1 73037
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3510
timestamp 1626065694
transform 1 0 115872 0 1 72901
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3509
timestamp 1626065694
transform 1 0 115328 0 1 69637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3508
timestamp 1626065694
transform 1 0 115600 0 1 69229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3507
timestamp 1626065694
transform 1 0 115600 0 1 69501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3506
timestamp 1626065694
transform 1 0 115464 0 1 69637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3505
timestamp 1626065694
transform 1 0 115464 0 1 69909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3504
timestamp 1626065694
transform 1 0 115600 0 1 67597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3503
timestamp 1626065694
transform 1 0 114240 0 1 70453
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3502
timestamp 1626065694
transform 1 0 114240 0 1 70045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3501
timestamp 1626065694
transform 1 0 115328 0 1 70589
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3500
timestamp 1626065694
transform 1 0 114376 0 1 69909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3499
timestamp 1626065694
transform 1 0 114376 0 1 69637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3498
timestamp 1626065694
transform 1 0 114376 0 1 69093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3497
timestamp 1626065694
transform 1 0 114376 0 1 68821
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3496
timestamp 1626065694
transform 1 0 114240 0 1 69229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3495
timestamp 1626065694
transform 1 0 114240 0 1 69501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3494
timestamp 1626065694
transform 1 0 114376 0 1 68685
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3493
timestamp 1626065694
transform 1 0 114376 0 1 68413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3492
timestamp 1626065694
transform 1 0 114648 0 1 69501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3491
timestamp 1626065694
transform 1 0 114648 0 1 69229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3490
timestamp 1626065694
transform 1 0 114648 0 1 69637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3489
timestamp 1626065694
transform 1 0 114648 0 1 69909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3488
timestamp 1626065694
transform 1 0 114784 0 1 69093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3487
timestamp 1626065694
transform 1 0 114784 0 1 68821
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3486
timestamp 1626065694
transform 1 0 114648 0 1 68413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3485
timestamp 1626065694
transform 1 0 114648 0 1 68685
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3484
timestamp 1626065694
transform 1 0 115192 0 1 68821
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3483
timestamp 1626065694
transform 1 0 115872 0 1 70045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3482
timestamp 1626065694
transform 1 0 115872 0 1 68005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3481
timestamp 1626065694
transform 1 0 115872 0 1 67733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3480
timestamp 1626065694
transform 1 0 115192 0 1 69093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3479
timestamp 1626065694
transform 1 0 116008 0 1 69229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3478
timestamp 1626065694
transform 1 0 116008 0 1 69501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3477
timestamp 1626065694
transform 1 0 116008 0 1 68549
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3476
timestamp 1626065694
transform 1 0 116008 0 1 68821
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3475
timestamp 1626065694
transform 1 0 116008 0 1 67597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3474
timestamp 1626065694
transform 1 0 115056 0 1 69229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3473
timestamp 1626065694
transform 1 0 115056 0 1 69501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3472
timestamp 1626065694
transform 1 0 115328 0 1 68005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3471
timestamp 1626065694
transform 1 0 115328 0 1 68277
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3470
timestamp 1626065694
transform 1 0 115328 0 1 69909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3469
timestamp 1626065694
transform 1 0 109344 0 1 67733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3468
timestamp 1626065694
transform 1 0 104312 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3467
timestamp 1626065694
transform 1 0 102408 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3466
timestamp 1626065694
transform 1 0 103088 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3465
timestamp 1626065694
transform 1 0 104856 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3464
timestamp 1626065694
transform 1 0 104856 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3463
timestamp 1626065694
transform 1 0 105536 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3462
timestamp 1626065694
transform 1 0 103088 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3461
timestamp 1626065694
transform 1 0 103632 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3460
timestamp 1626065694
transform 1 0 102408 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3459
timestamp 1626065694
transform 1 0 105536 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3458
timestamp 1626065694
transform 1 0 107304 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3457
timestamp 1626065694
transform 1 0 107304 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3456
timestamp 1626065694
transform 1 0 103632 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3455
timestamp 1626065694
transform 1 0 104312 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3454
timestamp 1626065694
transform 1 0 108528 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3453
timestamp 1626065694
transform 1 0 108528 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3452
timestamp 1626065694
transform 1 0 110704 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3451
timestamp 1626065694
transform 1 0 110704 0 1 70589
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3450
timestamp 1626065694
transform 1 0 106080 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3449
timestamp 1626065694
transform 1 0 106080 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3448
timestamp 1626065694
transform 1 0 109616 0 1 70861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3447
timestamp 1626065694
transform 1 0 109480 0 1 68141
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3446
timestamp 1626065694
transform 1 0 109480 0 1 67869
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3445
timestamp 1626065694
transform 1 0 109344 0 1 64741
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3444
timestamp 1626065694
transform 1 0 109344 0 1 64333
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3443
timestamp 1626065694
transform 1 0 109480 0 1 67053
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3442
timestamp 1626065694
transform 1 0 109480 0 1 67325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3441
timestamp 1626065694
transform 1 0 109480 0 1 64197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3440
timestamp 1626065694
transform 1 0 109480 0 1 63925
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3439
timestamp 1626065694
transform 1 0 109344 0 1 62565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3438
timestamp 1626065694
transform 1 0 109344 0 1 63517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3437
timestamp 1626065694
transform 1 0 109344 0 1 63789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3436
timestamp 1626065694
transform 1 0 109208 0 1 63517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3435
timestamp 1626065694
transform 1 0 109208 0 1 63925
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3434
timestamp 1626065694
transform 1 0 109344 0 1 67325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3433
timestamp 1626065694
transform 1 0 114376 0 1 65285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3432
timestamp 1626065694
transform 1 0 115464 0 1 63381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3431
timestamp 1626065694
transform 1 0 115192 0 1 65557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3430
timestamp 1626065694
transform 1 0 115464 0 1 63653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3429
timestamp 1626065694
transform 1 0 114376 0 1 66917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3428
timestamp 1626065694
transform 1 0 114376 0 1 67189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3427
timestamp 1626065694
transform 1 0 114376 0 1 64469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3426
timestamp 1626065694
transform 1 0 114376 0 1 64741
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3425
timestamp 1626065694
transform 1 0 115464 0 1 64877
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3424
timestamp 1626065694
transform 1 0 115192 0 1 65285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3423
timestamp 1626065694
transform 1 0 114648 0 1 67189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3422
timestamp 1626065694
transform 1 0 114648 0 1 66917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3421
timestamp 1626065694
transform 1 0 114648 0 1 65285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3420
timestamp 1626065694
transform 1 0 114648 0 1 65557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3419
timestamp 1626065694
transform 1 0 114648 0 1 65149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3418
timestamp 1626065694
transform 1 0 114648 0 1 64877
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3417
timestamp 1626065694
transform 1 0 114648 0 1 66373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3416
timestamp 1626065694
transform 1 0 114648 0 1 66101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3415
timestamp 1626065694
transform 1 0 114784 0 1 66509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3414
timestamp 1626065694
transform 1 0 114784 0 1 66781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3413
timestamp 1626065694
transform 1 0 114648 0 1 65965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3412
timestamp 1626065694
transform 1 0 114648 0 1 65693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3411
timestamp 1626065694
transform 1 0 115600 0 1 67325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3410
timestamp 1626065694
transform 1 0 115464 0 1 65149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3409
timestamp 1626065694
transform 1 0 115464 0 1 62565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3408
timestamp 1626065694
transform 1 0 114376 0 1 62429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3407
timestamp 1626065694
transform 1 0 114784 0 1 63245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3406
timestamp 1626065694
transform 1 0 114784 0 1 62973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3405
timestamp 1626065694
transform 1 0 115464 0 1 62837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3404
timestamp 1626065694
transform 1 0 115600 0 1 65965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3403
timestamp 1626065694
transform 1 0 114240 0 1 62837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3402
timestamp 1626065694
transform 1 0 114240 0 1 62565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3401
timestamp 1626065694
transform 1 0 114648 0 1 62837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3400
timestamp 1626065694
transform 1 0 114648 0 1 62565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3399
timestamp 1626065694
transform 1 0 114784 0 1 62429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3398
timestamp 1626065694
transform 1 0 114648 0 1 64741
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3397
timestamp 1626065694
transform 1 0 114648 0 1 64469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3396
timestamp 1626065694
transform 1 0 115328 0 1 65557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3395
timestamp 1626065694
transform 1 0 115328 0 1 65285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3394
timestamp 1626065694
transform 1 0 114240 0 1 62973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3393
timestamp 1626065694
transform 1 0 114240 0 1 63245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3392
timestamp 1626065694
transform 1 0 115872 0 1 62565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3391
timestamp 1626065694
transform 1 0 115872 0 1 62837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3390
timestamp 1626065694
transform 1 0 115872 0 1 62429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3389
timestamp 1626065694
transform 1 0 114240 0 1 65149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3388
timestamp 1626065694
transform 1 0 114240 0 1 64877
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3387
timestamp 1626065694
transform 1 0 115600 0 1 65693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3386
timestamp 1626065694
transform 1 0 116008 0 1 62973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3385
timestamp 1626065694
transform 1 0 116008 0 1 63245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3384
timestamp 1626065694
transform 1 0 115872 0 1 66781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3383
timestamp 1626065694
transform 1 0 115872 0 1 66509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3382
timestamp 1626065694
transform 1 0 115872 0 1 66917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3381
timestamp 1626065694
transform 1 0 115872 0 1 67189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3380
timestamp 1626065694
transform 1 0 116008 0 1 66373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3379
timestamp 1626065694
transform 1 0 116008 0 1 66101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3378
timestamp 1626065694
transform 1 0 115872 0 1 63381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3377
timestamp 1626065694
transform 1 0 115872 0 1 63653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3376
timestamp 1626065694
transform 1 0 116008 0 1 64061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3375
timestamp 1626065694
transform 1 0 116008 0 1 63789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3374
timestamp 1626065694
transform 1 0 116008 0 1 65965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3373
timestamp 1626065694
transform 1 0 116008 0 1 65693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3372
timestamp 1626065694
transform 1 0 115600 0 1 66509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3371
timestamp 1626065694
transform 1 0 115192 0 1 62429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3370
timestamp 1626065694
transform 1 0 115600 0 1 66781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3369
timestamp 1626065694
transform 1 0 114376 0 1 66509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3368
timestamp 1626065694
transform 1 0 116008 0 1 67325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3367
timestamp 1626065694
transform 1 0 114376 0 1 66781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3366
timestamp 1626065694
transform 1 0 115872 0 1 65557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3365
timestamp 1626065694
transform 1 0 115872 0 1 65285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3364
timestamp 1626065694
transform 1 0 114240 0 1 66373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3363
timestamp 1626065694
transform 1 0 114240 0 1 66101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3362
timestamp 1626065694
transform 1 0 115328 0 1 64333
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3361
timestamp 1626065694
transform 1 0 115328 0 1 64061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3360
timestamp 1626065694
transform 1 0 115056 0 1 64877
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3359
timestamp 1626065694
transform 1 0 115056 0 1 65149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3358
timestamp 1626065694
transform 1 0 115056 0 1 62837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3357
timestamp 1626065694
transform 1 0 115056 0 1 62565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3356
timestamp 1626065694
transform 1 0 115056 0 1 66373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3355
timestamp 1626065694
transform 1 0 115056 0 1 66101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3354
timestamp 1626065694
transform 1 0 115328 0 1 66373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3353
timestamp 1626065694
transform 1 0 115328 0 1 66101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3352
timestamp 1626065694
transform 1 0 114376 0 1 65693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3351
timestamp 1626065694
transform 1 0 114376 0 1 65965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3350
timestamp 1626065694
transform 1 0 114376 0 1 65557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3349
timestamp 1626065694
transform 1 0 135320 0 1 67597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3348
timestamp 1626065694
transform 1 0 135320 0 1 72493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3347
timestamp 1626065694
transform 1 0 134087 0 1 72293
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3346
timestamp 1626065694
transform 1 0 135320 0 1 69365
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3345
timestamp 1626065694
transform 1 0 134776 0 1 68549
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3344
timestamp 1626065694
transform 1 0 134776 0 1 69093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3343
timestamp 1626065694
transform 1 0 134776 0 1 71269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3342
timestamp 1626065694
transform 1 0 134776 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3341
timestamp 1626065694
transform 1 0 133144 0 1 69773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3340
timestamp 1626065694
transform 1 0 135320 0 1 70861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3339
timestamp 1626065694
transform 1 0 122400 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3338
timestamp 1626065694
transform 1 0 135320 0 1 64061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3337
timestamp 1626065694
transform 1 0 135320 0 1 65829
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3336
timestamp 1626065694
transform 1 0 132600 0 1 64333
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3335
timestamp 1626065694
transform 1 0 132600 0 1 66917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3334
timestamp 1626065694
transform 1 0 133144 0 1 67053
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3333
timestamp 1626065694
transform 1 0 133416 0 1 64197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3332
timestamp 1626065694
transform 1 0 136000 0 1 64469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3331
timestamp 1626065694
transform 1 0 135320 0 1 62429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3330
timestamp 1626065694
transform 1 0 94384 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3329
timestamp 1626065694
transform 1 0 96288 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3328
timestamp 1626065694
transform 1 0 96288 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3327
timestamp 1626065694
transform 1 0 97920 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3326
timestamp 1626065694
transform 1 0 97920 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3325
timestamp 1626065694
transform 1 0 99688 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3324
timestamp 1626065694
transform 1 0 99688 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3323
timestamp 1626065694
transform 1 0 101320 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3322
timestamp 1626065694
transform 1 0 101320 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3321
timestamp 1626065694
transform 1 0 94384 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3320
timestamp 1626065694
transform 1 0 86224 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3319
timestamp 1626065694
transform 1 0 86224 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3318
timestamp 1626065694
transform 1 0 87720 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3317
timestamp 1626065694
transform 1 0 87720 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3316
timestamp 1626065694
transform 1 0 89352 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3315
timestamp 1626065694
transform 1 0 89352 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3314
timestamp 1626065694
transform 1 0 91120 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3313
timestamp 1626065694
transform 1 0 91120 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3312
timestamp 1626065694
transform 1 0 92888 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3311
timestamp 1626065694
transform 1 0 92888 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3310
timestamp 1626065694
transform 1 0 88536 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3309
timestamp 1626065694
transform 1 0 86360 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3308
timestamp 1626065694
transform 1 0 86224 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3307
timestamp 1626065694
transform 1 0 86496 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3306
timestamp 1626065694
transform 1 0 86496 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3305
timestamp 1626065694
transform 1 0 88944 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3304
timestamp 1626065694
transform 1 0 88944 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3303
timestamp 1626065694
transform 1 0 88944 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3302
timestamp 1626065694
transform 1 0 88944 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3301
timestamp 1626065694
transform 1 0 91256 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3300
timestamp 1626065694
transform 1 0 91256 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3299
timestamp 1626065694
transform 1 0 91392 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3298
timestamp 1626065694
transform 1 0 91392 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3297
timestamp 1626065694
transform 1 0 93704 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3296
timestamp 1626065694
transform 1 0 93704 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3295
timestamp 1626065694
transform 1 0 93704 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3294
timestamp 1626065694
transform 1 0 85952 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3293
timestamp 1626065694
transform 1 0 88400 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3292
timestamp 1626065694
transform 1 0 90984 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3291
timestamp 1626065694
transform 1 0 93568 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3290
timestamp 1626065694
transform 1 0 88536 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3289
timestamp 1626065694
transform 1 0 86360 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3288
timestamp 1626065694
transform 1 0 86360 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3287
timestamp 1626065694
transform 1 0 91392 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3286
timestamp 1626065694
transform 1 0 91392 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3285
timestamp 1626065694
transform 1 0 93568 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3284
timestamp 1626065694
transform 1 0 93568 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3283
timestamp 1626065694
transform 1 0 88808 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3282
timestamp 1626065694
transform 1 0 88808 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3281
timestamp 1626065694
transform 1 0 93840 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3280
timestamp 1626065694
transform 1 0 96288 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3279
timestamp 1626065694
transform 1 0 96288 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3278
timestamp 1626065694
transform 1 0 96424 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3277
timestamp 1626065694
transform 1 0 96424 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3276
timestamp 1626065694
transform 1 0 98872 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3275
timestamp 1626065694
transform 1 0 98872 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3274
timestamp 1626065694
transform 1 0 98872 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3273
timestamp 1626065694
transform 1 0 98872 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3272
timestamp 1626065694
transform 1 0 101320 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3271
timestamp 1626065694
transform 1 0 101320 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3270
timestamp 1626065694
transform 1 0 101456 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3269
timestamp 1626065694
transform 1 0 101456 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3268
timestamp 1626065694
transform 1 0 98600 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3267
timestamp 1626065694
transform 1 0 93840 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3266
timestamp 1626065694
transform 1 0 93840 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3265
timestamp 1626065694
transform 1 0 96016 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3264
timestamp 1626065694
transform 1 0 98464 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3263
timestamp 1626065694
transform 1 0 101048 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3262
timestamp 1626065694
transform 1 0 98736 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3261
timestamp 1626065694
transform 1 0 98736 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3260
timestamp 1626065694
transform 1 0 96152 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3259
timestamp 1626065694
transform 1 0 96152 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3258
timestamp 1626065694
transform 1 0 101184 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3257
timestamp 1626065694
transform 1 0 101184 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3256
timestamp 1626065694
transform 1 0 98600 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3255
timestamp 1626065694
transform 1 0 77656 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3254
timestamp 1626065694
transform 1 0 79424 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3253
timestamp 1626065694
transform 1 0 77656 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3252
timestamp 1626065694
transform 1 0 79424 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3251
timestamp 1626065694
transform 1 0 81328 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3250
timestamp 1626065694
transform 1 0 81328 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3249
timestamp 1626065694
transform 1 0 82688 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3248
timestamp 1626065694
transform 1 0 82688 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3247
timestamp 1626065694
transform 1 0 84456 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3246
timestamp 1626065694
transform 1 0 84456 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3245
timestamp 1626065694
transform 1 0 69224 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3244
timestamp 1626065694
transform 1 0 69224 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3243
timestamp 1626065694
transform 1 0 70856 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3242
timestamp 1626065694
transform 1 0 70856 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3241
timestamp 1626065694
transform 1 0 72624 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3240
timestamp 1626065694
transform 1 0 72624 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3239
timestamp 1626065694
transform 1 0 74392 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3238
timestamp 1626065694
transform 1 0 74392 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3237
timestamp 1626065694
transform 1 0 76160 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3236
timestamp 1626065694
transform 1 0 76160 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3235
timestamp 1626065694
transform 1 0 71400 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3234
timestamp 1626065694
transform 1 0 71264 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3233
timestamp 1626065694
transform 1 0 71400 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3232
timestamp 1626065694
transform 1 0 71400 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3231
timestamp 1626065694
transform 1 0 73848 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3230
timestamp 1626065694
transform 1 0 73848 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3229
timestamp 1626065694
transform 1 0 73984 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3228
timestamp 1626065694
transform 1 0 73984 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3227
timestamp 1626065694
transform 1 0 76432 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3226
timestamp 1626065694
transform 1 0 76432 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3225
timestamp 1626065694
transform 1 0 76432 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3224
timestamp 1626065694
transform 1 0 76432 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3223
timestamp 1626065694
transform 1 0 71128 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3222
timestamp 1626065694
transform 1 0 71400 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3221
timestamp 1626065694
transform 1 0 71400 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3220
timestamp 1626065694
transform 1 0 68544 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3219
timestamp 1626065694
transform 1 0 70992 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3218
timestamp 1626065694
transform 1 0 73576 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3217
timestamp 1626065694
transform 1 0 75888 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3216
timestamp 1626065694
transform 1 0 73712 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3215
timestamp 1626065694
transform 1 0 73712 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3214
timestamp 1626065694
transform 1 0 68952 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3213
timestamp 1626065694
transform 1 0 68952 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3212
timestamp 1626065694
transform 1 0 76160 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3211
timestamp 1626065694
transform 1 0 76160 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3210
timestamp 1626065694
transform 1 0 68952 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3209
timestamp 1626065694
transform 1 0 68952 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3208
timestamp 1626065694
transform 1 0 68816 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3207
timestamp 1626065694
transform 1 0 68816 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3206
timestamp 1626065694
transform 1 0 71128 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3205
timestamp 1626065694
transform 1 0 83912 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3204
timestamp 1626065694
transform 1 0 83912 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3203
timestamp 1626065694
transform 1 0 83912 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3202
timestamp 1626065694
transform 1 0 83912 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3201
timestamp 1626065694
transform 1 0 78880 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3200
timestamp 1626065694
transform 1 0 78608 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3199
timestamp 1626065694
transform 1 0 81056 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3198
timestamp 1626065694
transform 1 0 83504 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3197
timestamp 1626065694
transform 1 0 78880 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3196
timestamp 1626065694
transform 1 0 78880 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3195
timestamp 1626065694
transform 1 0 78880 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3194
timestamp 1626065694
transform 1 0 81328 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3193
timestamp 1626065694
transform 1 0 81328 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3192
timestamp 1626065694
transform 1 0 81464 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3191
timestamp 1626065694
transform 1 0 78608 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3190
timestamp 1626065694
transform 1 0 78608 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3189
timestamp 1626065694
transform 1 0 81464 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3188
timestamp 1626065694
transform 1 0 81464 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3187
timestamp 1626065694
transform 1 0 78744 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3186
timestamp 1626065694
transform 1 0 83776 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3185
timestamp 1626065694
transform 1 0 83776 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3184
timestamp 1626065694
transform 1 0 78744 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3183
timestamp 1626065694
transform 1 0 81464 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3182
timestamp 1626065694
transform 1 0 79424 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3181
timestamp 1626065694
transform 1 0 74392 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3180
timestamp 1626065694
transform 1 0 74392 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3179
timestamp 1626065694
transform 1 0 79968 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3178
timestamp 1626065694
transform 1 0 79968 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3177
timestamp 1626065694
transform 1 0 80648 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3176
timestamp 1626065694
transform 1 0 80648 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3175
timestamp 1626065694
transform 1 0 69904 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3174
timestamp 1626065694
transform 1 0 69904 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3173
timestamp 1626065694
transform 1 0 74936 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3172
timestamp 1626065694
transform 1 0 74936 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3171
timestamp 1626065694
transform 1 0 81872 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3170
timestamp 1626065694
transform 1 0 81872 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3169
timestamp 1626065694
transform 1 0 82416 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3168
timestamp 1626065694
transform 1 0 82416 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3167
timestamp 1626065694
transform 1 0 75616 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3166
timestamp 1626065694
transform 1 0 75616 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3165
timestamp 1626065694
transform 1 0 83096 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3164
timestamp 1626065694
transform 1 0 83096 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3163
timestamp 1626065694
transform 1 0 83640 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3162
timestamp 1626065694
transform 1 0 83640 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3161
timestamp 1626065694
transform 1 0 72216 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3160
timestamp 1626065694
transform 1 0 72216 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3159
timestamp 1626065694
transform 1 0 76160 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3158
timestamp 1626065694
transform 1 0 76160 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3157
timestamp 1626065694
transform 1 0 84592 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3156
timestamp 1626065694
transform 1 0 84592 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3155
timestamp 1626065694
transform 1 0 72080 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3154
timestamp 1626065694
transform 1 0 72080 0 1 70861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3153
timestamp 1626065694
transform 1 0 70584 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3152
timestamp 1626065694
transform 1 0 70584 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3151
timestamp 1626065694
transform 1 0 76840 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3150
timestamp 1626065694
transform 1 0 76840 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3149
timestamp 1626065694
transform 1 0 77384 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3148
timestamp 1626065694
transform 1 0 77384 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3147
timestamp 1626065694
transform 1 0 73712 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3146
timestamp 1626065694
transform 1 0 73712 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3145
timestamp 1626065694
transform 1 0 78200 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3144
timestamp 1626065694
transform 1 0 78200 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3143
timestamp 1626065694
transform 1 0 78472 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3142
timestamp 1626065694
transform 1 0 78472 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3141
timestamp 1626065694
transform 1 0 68680 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3140
timestamp 1626065694
transform 1 0 68680 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3139
timestamp 1626065694
transform 1 0 79424 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3138
timestamp 1626065694
transform 1 0 94928 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3137
timestamp 1626065694
transform 1 0 95608 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3136
timestamp 1626065694
transform 1 0 95608 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3135
timestamp 1626065694
transform 1 0 90712 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3134
timestamp 1626065694
transform 1 0 90712 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3133
timestamp 1626065694
transform 1 0 91120 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3132
timestamp 1626065694
transform 1 0 91120 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3131
timestamp 1626065694
transform 1 0 88128 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3130
timestamp 1626065694
transform 1 0 88128 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3129
timestamp 1626065694
transform 1 0 96832 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3128
timestamp 1626065694
transform 1 0 96832 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3127
timestamp 1626065694
transform 1 0 97376 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3126
timestamp 1626065694
transform 1 0 97376 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3125
timestamp 1626065694
transform 1 0 88672 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3124
timestamp 1626065694
transform 1 0 88672 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3123
timestamp 1626065694
transform 1 0 98600 0 1 71269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3122
timestamp 1626065694
transform 1 0 98600 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3121
timestamp 1626065694
transform 1 0 86904 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3120
timestamp 1626065694
transform 1 0 86904 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3119
timestamp 1626065694
transform 1 0 92344 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3118
timestamp 1626065694
transform 1 0 92344 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3117
timestamp 1626065694
transform 1 0 99824 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3116
timestamp 1626065694
transform 1 0 99824 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3115
timestamp 1626065694
transform 1 0 100912 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3114
timestamp 1626065694
transform 1 0 100912 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3113
timestamp 1626065694
transform 1 0 89352 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3112
timestamp 1626065694
transform 1 0 89352 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3111
timestamp 1626065694
transform 1 0 93296 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3110
timestamp 1626065694
transform 1 0 93296 0 1 70861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3109
timestamp 1626065694
transform 1 0 101864 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3108
timestamp 1626065694
transform 1 0 101864 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3107
timestamp 1626065694
transform 1 0 86088 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3106
timestamp 1626065694
transform 1 0 86088 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3105
timestamp 1626065694
transform 1 0 89896 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3104
timestamp 1626065694
transform 1 0 89896 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3103
timestamp 1626065694
transform 1 0 94928 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3102
timestamp 1626065694
transform 1 0 116008 0 1 51957
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3101
timestamp 1626065694
transform 1 0 134087 0 1 62058
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3100
timestamp 1626065694
transform 1 0 135320 0 1 60797
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3099
timestamp 1626065694
transform 1 0 135320 0 1 57533
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3098
timestamp 1626065694
transform 1 0 135320 0 1 59165
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3097
timestamp 1626065694
transform 1 0 133416 0 1 61477
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3096
timestamp 1626065694
transform 1 0 135320 0 1 52365
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3095
timestamp 1626065694
transform 1 0 135320 0 1 55901
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3094
timestamp 1626065694
transform 1 0 135320 0 1 53997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3093
timestamp 1626065694
transform 1 0 115056 0 1 58213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3092
timestamp 1626065694
transform 1 0 115328 0 1 58213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3091
timestamp 1626065694
transform 1 0 115328 0 1 58485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3090
timestamp 1626065694
transform 1 0 115464 0 1 62021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3089
timestamp 1626065694
transform 1 0 115464 0 1 61749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3088
timestamp 1626065694
transform 1 0 115600 0 1 61613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3087
timestamp 1626065694
transform 1 0 115600 0 1 61341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3086
timestamp 1626065694
transform 1 0 115464 0 1 59709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3085
timestamp 1626065694
transform 1 0 115464 0 1 59437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3084
timestamp 1626065694
transform 1 0 115600 0 1 57397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3083
timestamp 1626065694
transform 1 0 115600 0 1 57669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3082
timestamp 1626065694
transform 1 0 115600 0 1 57261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3081
timestamp 1626065694
transform 1 0 115464 0 1 58621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3080
timestamp 1626065694
transform 1 0 115464 0 1 58893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3079
timestamp 1626065694
transform 1 0 114240 0 1 57397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3078
timestamp 1626065694
transform 1 0 114240 0 1 57669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3077
timestamp 1626065694
transform 1 0 114240 0 1 57261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3076
timestamp 1626065694
transform 1 0 114240 0 1 60933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3075
timestamp 1626065694
transform 1 0 114240 0 1 61205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3074
timestamp 1626065694
transform 1 0 114376 0 1 57805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3073
timestamp 1626065694
transform 1 0 114376 0 1 58077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3072
timestamp 1626065694
transform 1 0 115192 0 1 57805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3071
timestamp 1626065694
transform 1 0 115192 0 1 58077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3070
timestamp 1626065694
transform 1 0 115328 0 1 57805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3069
timestamp 1626065694
transform 1 0 115328 0 1 58077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3068
timestamp 1626065694
transform 1 0 115192 0 1 62157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3067
timestamp 1626065694
transform 1 0 114240 0 1 58485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3066
timestamp 1626065694
transform 1 0 114240 0 1 58213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3065
timestamp 1626065694
transform 1 0 115056 0 1 61613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3064
timestamp 1626065694
transform 1 0 115056 0 1 61341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3063
timestamp 1626065694
transform 1 0 115192 0 1 60117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3062
timestamp 1626065694
transform 1 0 115192 0 1 60389
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3061
timestamp 1626065694
transform 1 0 115328 0 1 60117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3060
timestamp 1626065694
transform 1 0 115328 0 1 60389
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3059
timestamp 1626065694
transform 1 0 115328 0 1 61205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3058
timestamp 1626065694
transform 1 0 115328 0 1 60933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3057
timestamp 1626065694
transform 1 0 115192 0 1 57261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3056
timestamp 1626065694
transform 1 0 114376 0 1 59029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3055
timestamp 1626065694
transform 1 0 114376 0 1 59301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3054
timestamp 1626065694
transform 1 0 114376 0 1 58893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3053
timestamp 1626065694
transform 1 0 114376 0 1 58621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3052
timestamp 1626065694
transform 1 0 114784 0 1 59029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3051
timestamp 1626065694
transform 1 0 114784 0 1 59301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3050
timestamp 1626065694
transform 1 0 114784 0 1 58893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3049
timestamp 1626065694
transform 1 0 114784 0 1 58621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3048
timestamp 1626065694
transform 1 0 114648 0 1 61749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3047
timestamp 1626065694
transform 1 0 114648 0 1 62021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3046
timestamp 1626065694
transform 1 0 114648 0 1 61613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3045
timestamp 1626065694
transform 1 0 114648 0 1 61341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3044
timestamp 1626065694
transform 1 0 114648 0 1 57397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3043
timestamp 1626065694
transform 1 0 114648 0 1 57669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3042
timestamp 1626065694
transform 1 0 114648 0 1 57261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3041
timestamp 1626065694
transform 1 0 114784 0 1 58077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3040
timestamp 1626065694
transform 1 0 114784 0 1 57805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3039
timestamp 1626065694
transform 1 0 114784 0 1 58213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3038
timestamp 1626065694
transform 1 0 114784 0 1 58485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3037
timestamp 1626065694
transform 1 0 114648 0 1 60389
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3036
timestamp 1626065694
transform 1 0 114648 0 1 60117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3035
timestamp 1626065694
transform 1 0 114648 0 1 60525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3034
timestamp 1626065694
transform 1 0 114648 0 1 60797
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3033
timestamp 1626065694
transform 1 0 114784 0 1 62157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3032
timestamp 1626065694
transform 1 0 114648 0 1 60933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3031
timestamp 1626065694
transform 1 0 114648 0 1 61205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3030
timestamp 1626065694
transform 1 0 115872 0 1 58893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3029
timestamp 1626065694
transform 1 0 115872 0 1 58621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3028
timestamp 1626065694
transform 1 0 115872 0 1 59029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3027
timestamp 1626065694
transform 1 0 115872 0 1 59301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3026
timestamp 1626065694
transform 1 0 115872 0 1 62157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3025
timestamp 1626065694
transform 1 0 116008 0 1 58485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3024
timestamp 1626065694
transform 1 0 116008 0 1 58213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3023
timestamp 1626065694
transform 1 0 116008 0 1 59845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3022
timestamp 1626065694
transform 1 0 116008 0 1 60117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3021
timestamp 1626065694
transform 1 0 116008 0 1 59709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3020
timestamp 1626065694
transform 1 0 116008 0 1 59437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3019
timestamp 1626065694
transform 1 0 115872 0 1 61341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3018
timestamp 1626065694
transform 1 0 115872 0 1 61613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3017
timestamp 1626065694
transform 1 0 115872 0 1 57805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3016
timestamp 1626065694
transform 1 0 115872 0 1 58077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3015
timestamp 1626065694
transform 1 0 116008 0 1 57669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3014
timestamp 1626065694
transform 1 0 116008 0 1 57397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3013
timestamp 1626065694
transform 1 0 114240 0 1 62021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3012
timestamp 1626065694
transform 1 0 114240 0 1 61749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3011
timestamp 1626065694
transform 1 0 114376 0 1 62157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3010
timestamp 1626065694
transform 1 0 116008 0 1 62021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3009
timestamp 1626065694
transform 1 0 116008 0 1 61749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3008
timestamp 1626065694
transform 1 0 114240 0 1 61613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3007
timestamp 1626065694
transform 1 0 114240 0 1 61341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3006
timestamp 1626065694
transform 1 0 114376 0 1 60117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3005
timestamp 1626065694
transform 1 0 114376 0 1 60389
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3004
timestamp 1626065694
transform 1 0 115056 0 1 58485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3003
timestamp 1626065694
transform 1 0 114240 0 1 60525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3002
timestamp 1626065694
transform 1 0 114240 0 1 60797
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3001
timestamp 1626065694
transform 1 0 109480 0 1 59573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3000
timestamp 1626065694
transform 1 0 109480 0 1 60797
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2999
timestamp 1626065694
transform 1 0 109480 0 1 61069
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2998
timestamp 1626065694
transform 1 0 109480 0 1 58621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2997
timestamp 1626065694
transform 1 0 109480 0 1 58349
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2996
timestamp 1626065694
transform 1 0 109480 0 1 59845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2995
timestamp 1626065694
transform 1 0 109480 0 1 55221
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2994
timestamp 1626065694
transform 1 0 109344 0 1 56037
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2993
timestamp 1626065694
transform 1 0 109344 0 1 55629
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2992
timestamp 1626065694
transform 1 0 109480 0 1 55901
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2991
timestamp 1626065694
transform 1 0 109480 0 1 55629
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2990
timestamp 1626065694
transform 1 0 109480 0 1 55493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2989
timestamp 1626065694
transform 1 0 115464 0 1 54541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2988
timestamp 1626065694
transform 1 0 115464 0 1 53045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2987
timestamp 1626065694
transform 1 0 115600 0 1 52637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2986
timestamp 1626065694
transform 1 0 115600 0 1 52909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2985
timestamp 1626065694
transform 1 0 114376 0 1 53453
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2984
timestamp 1626065694
transform 1 0 114648 0 1 52093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2983
timestamp 1626065694
transform 1 0 114784 0 1 53861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2982
timestamp 1626065694
transform 1 0 114784 0 1 54133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2981
timestamp 1626065694
transform 1 0 114784 0 1 53725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2980
timestamp 1626065694
transform 1 0 114784 0 1 53453
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2979
timestamp 1626065694
transform 1 0 114784 0 1 54541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2978
timestamp 1626065694
transform 1 0 114784 0 1 54269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2977
timestamp 1626065694
transform 1 0 114784 0 1 54677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2976
timestamp 1626065694
transform 1 0 114784 0 1 54949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2975
timestamp 1626065694
transform 1 0 114240 0 1 54269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2974
timestamp 1626065694
transform 1 0 114240 0 1 54541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2973
timestamp 1626065694
transform 1 0 115192 0 1 53861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2972
timestamp 1626065694
transform 1 0 114784 0 1 52637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2971
timestamp 1626065694
transform 1 0 114784 0 1 52909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2970
timestamp 1626065694
transform 1 0 114784 0 1 52501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2969
timestamp 1626065694
transform 1 0 114784 0 1 52229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2968
timestamp 1626065694
transform 1 0 114648 0 1 53317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2967
timestamp 1626065694
transform 1 0 114648 0 1 53045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2966
timestamp 1626065694
transform 1 0 115192 0 1 54133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2965
timestamp 1626065694
transform 1 0 115328 0 1 53861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2964
timestamp 1626065694
transform 1 0 114648 0 1 56173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2963
timestamp 1626065694
transform 1 0 114648 0 1 56445
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2962
timestamp 1626065694
transform 1 0 114784 0 1 56853
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2961
timestamp 1626065694
transform 1 0 114784 0 1 56581
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2960
timestamp 1626065694
transform 1 0 115328 0 1 54133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2959
timestamp 1626065694
transform 1 0 115328 0 1 55765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2958
timestamp 1626065694
transform 1 0 115328 0 1 55493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2957
timestamp 1626065694
transform 1 0 115192 0 1 54949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2956
timestamp 1626065694
transform 1 0 116008 0 1 55357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2955
timestamp 1626065694
transform 1 0 116008 0 1 55085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2954
timestamp 1626065694
transform 1 0 116008 0 1 55493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2953
timestamp 1626065694
transform 1 0 116008 0 1 55765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2952
timestamp 1626065694
transform 1 0 115192 0 1 54677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2951
timestamp 1626065694
transform 1 0 115872 0 1 52637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2950
timestamp 1626065694
transform 1 0 115872 0 1 52909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2949
timestamp 1626065694
transform 1 0 114240 0 1 56989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2948
timestamp 1626065694
transform 1 0 115056 0 1 56173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2947
timestamp 1626065694
transform 1 0 116008 0 1 56173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2946
timestamp 1626065694
transform 1 0 116008 0 1 55901
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2945
timestamp 1626065694
transform 1 0 115056 0 1 56445
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2944
timestamp 1626065694
transform 1 0 115192 0 1 55901
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2943
timestamp 1626065694
transform 1 0 115328 0 1 56037
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2942
timestamp 1626065694
transform 1 0 114376 0 1 52501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2941
timestamp 1626065694
transform 1 0 116008 0 1 52229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2940
timestamp 1626065694
transform 1 0 115192 0 1 52229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2939
timestamp 1626065694
transform 1 0 115192 0 1 56989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2938
timestamp 1626065694
transform 1 0 114376 0 1 52229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2937
timestamp 1626065694
transform 1 0 115328 0 1 54677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2936
timestamp 1626065694
transform 1 0 114240 0 1 56445
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2935
timestamp 1626065694
transform 1 0 115328 0 1 54949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2934
timestamp 1626065694
transform 1 0 115192 0 1 52637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2933
timestamp 1626065694
transform 1 0 116008 0 1 54269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2932
timestamp 1626065694
transform 1 0 116008 0 1 54541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2931
timestamp 1626065694
transform 1 0 116008 0 1 54133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2930
timestamp 1626065694
transform 1 0 116008 0 1 53861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2929
timestamp 1626065694
transform 1 0 115872 0 1 54949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2928
timestamp 1626065694
transform 1 0 115872 0 1 54677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2927
timestamp 1626065694
transform 1 0 115872 0 1 53453
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2926
timestamp 1626065694
transform 1 0 115872 0 1 53725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2925
timestamp 1626065694
transform 1 0 114240 0 1 52093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2924
timestamp 1626065694
transform 1 0 115192 0 1 52909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2923
timestamp 1626065694
transform 1 0 114648 0 1 56989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2922
timestamp 1626065694
transform 1 0 114240 0 1 56173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2921
timestamp 1626065694
transform 1 0 114240 0 1 56581
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2920
timestamp 1626065694
transform 1 0 114240 0 1 56853
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2919
timestamp 1626065694
transform 1 0 114376 0 1 54677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2918
timestamp 1626065694
transform 1 0 114376 0 1 54949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2917
timestamp 1626065694
transform 1 0 114376 0 1 53861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2916
timestamp 1626065694
transform 1 0 114376 0 1 54133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2915
timestamp 1626065694
transform 1 0 114376 0 1 53725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2914
timestamp 1626065694
transform 1 0 115192 0 1 52501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2913
timestamp 1626065694
transform 1 0 114240 0 1 53045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2912
timestamp 1626065694
transform 1 0 114240 0 1 53317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2911
timestamp 1626065694
transform 1 0 114240 0 1 52909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2910
timestamp 1626065694
transform 1 0 114240 0 1 52637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2909
timestamp 1626065694
transform 1 0 115464 0 1 53317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2908
timestamp 1626065694
transform 1 0 115600 0 1 56989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2907
timestamp 1626065694
transform 1 0 115464 0 1 54269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2906
timestamp 1626065694
transform 1 0 109480 0 1 46789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2905
timestamp 1626065694
transform 1 0 115872 0 1 46789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2904
timestamp 1626065694
transform 1 0 115328 0 1 46789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2903
timestamp 1626065694
transform 1 0 114784 0 1 50597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2902
timestamp 1626065694
transform 1 0 114648 0 1 51821
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2901
timestamp 1626065694
transform 1 0 115464 0 1 51005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2900
timestamp 1626065694
transform 1 0 115464 0 1 50733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2899
timestamp 1626065694
transform 1 0 114648 0 1 49781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2898
timestamp 1626065694
transform 1 0 114648 0 1 49509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2897
timestamp 1626065694
transform 1 0 114648 0 1 48557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2896
timestamp 1626065694
transform 1 0 114648 0 1 48285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2895
timestamp 1626065694
transform 1 0 114648 0 1 48693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2894
timestamp 1626065694
transform 1 0 114648 0 1 48965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2893
timestamp 1626065694
transform 1 0 114240 0 1 49781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2892
timestamp 1626065694
transform 1 0 114784 0 1 48149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2891
timestamp 1626065694
transform 1 0 114784 0 1 47877
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2890
timestamp 1626065694
transform 1 0 114648 0 1 49101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2889
timestamp 1626065694
transform 1 0 114648 0 1 49373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2888
timestamp 1626065694
transform 1 0 114784 0 1 50189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2887
timestamp 1626065694
transform 1 0 114648 0 1 50733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2886
timestamp 1626065694
transform 1 0 114648 0 1 51005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2885
timestamp 1626065694
transform 1 0 114240 0 1 49509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2884
timestamp 1626065694
transform 1 0 115872 0 1 47197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2883
timestamp 1626065694
transform 1 0 115872 0 1 47469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2882
timestamp 1626065694
transform 1 0 115872 0 1 47061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2881
timestamp 1626065694
transform 1 0 114784 0 1 49917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2880
timestamp 1626065694
transform 1 0 114240 0 1 49917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2879
timestamp 1626065694
transform 1 0 115192 0 1 49509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2878
timestamp 1626065694
transform 1 0 115192 0 1 49781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2877
timestamp 1626065694
transform 1 0 115328 0 1 49509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2876
timestamp 1626065694
transform 1 0 115872 0 1 48285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2875
timestamp 1626065694
transform 1 0 115872 0 1 48013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2874
timestamp 1626065694
transform 1 0 114240 0 1 50733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2873
timestamp 1626065694
transform 1 0 114240 0 1 51005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2872
timestamp 1626065694
transform 1 0 114376 0 1 50597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2871
timestamp 1626065694
transform 1 0 115328 0 1 49781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2870
timestamp 1626065694
transform 1 0 115872 0 1 51413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2869
timestamp 1626065694
transform 1 0 115872 0 1 51141
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2868
timestamp 1626065694
transform 1 0 114376 0 1 50325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2867
timestamp 1626065694
transform 1 0 115056 0 1 48557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2866
timestamp 1626065694
transform 1 0 115056 0 1 48285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2865
timestamp 1626065694
transform 1 0 115328 0 1 47061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2864
timestamp 1626065694
transform 1 0 114784 0 1 50325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2863
timestamp 1626065694
transform 1 0 114240 0 1 50189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2862
timestamp 1626065694
transform 1 0 115872 0 1 49373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2861
timestamp 1626065694
transform 1 0 115872 0 1 49101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2860
timestamp 1626065694
transform 1 0 115872 0 1 49509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2859
timestamp 1626065694
transform 1 0 115872 0 1 49781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2858
timestamp 1626065694
transform 1 0 116008 0 1 51005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2857
timestamp 1626065694
transform 1 0 116008 0 1 50733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2856
timestamp 1626065694
transform 1 0 115872 0 1 50325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2855
timestamp 1626065694
transform 1 0 115872 0 1 50597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2854
timestamp 1626065694
transform 1 0 115872 0 1 50189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2853
timestamp 1626065694
transform 1 0 115872 0 1 49917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2852
timestamp 1626065694
transform 1 0 114376 0 1 49101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2851
timestamp 1626065694
transform 1 0 115192 0 1 51413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2850
timestamp 1626065694
transform 1 0 114376 0 1 49373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2849
timestamp 1626065694
transform 1 0 114240 0 1 48965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2848
timestamp 1626065694
transform 1 0 114240 0 1 48693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2847
timestamp 1626065694
transform 1 0 115192 0 1 51685
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2846
timestamp 1626065694
transform 1 0 115464 0 1 48285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2845
timestamp 1626065694
transform 1 0 115464 0 1 48557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2844
timestamp 1626065694
transform 1 0 115600 0 1 48693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2843
timestamp 1626065694
transform 1 0 115600 0 1 48965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2842
timestamp 1626065694
transform 1 0 115056 0 1 50733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2841
timestamp 1626065694
transform 1 0 115056 0 1 51005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2840
timestamp 1626065694
transform 1 0 114240 0 1 51821
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2839
timestamp 1626065694
transform 1 0 116008 0 1 48965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2838
timestamp 1626065694
transform 1 0 116008 0 1 48693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2837
timestamp 1626065694
transform 1 0 114240 0 1 47877
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2836
timestamp 1626065694
transform 1 0 114240 0 1 48149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2835
timestamp 1626065694
transform 1 0 115600 0 1 50189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2834
timestamp 1626065694
transform 1 0 115600 0 1 49917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2833
timestamp 1626065694
transform 1 0 115056 0 1 47469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2832
timestamp 1626065694
transform 1 0 115056 0 1 47741
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2831
timestamp 1626065694
transform 1 0 115328 0 1 48285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2830
timestamp 1626065694
transform 1 0 115328 0 1 48013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2829
timestamp 1626065694
transform 1 0 114376 0 1 48285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2828
timestamp 1626065694
transform 1 0 114376 0 1 48557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2827
timestamp 1626065694
transform 1 0 109344 0 1 47197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2826
timestamp 1626065694
transform 1 0 109344 0 1 46925
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2825
timestamp 1626065694
transform 1 0 109344 0 1 42573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2824
timestamp 1626065694
transform 1 0 109344 0 1 42981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2823
timestamp 1626065694
transform 1 0 109480 0 1 46517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2822
timestamp 1626065694
transform 1 0 109344 0 1 43253
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2821
timestamp 1626065694
transform 1 0 109344 0 1 42845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2820
timestamp 1626065694
transform 1 0 109344 0 1 43661
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2819
timestamp 1626065694
transform 1 0 109344 0 1 43389
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2818
timestamp 1626065694
transform 1 0 115464 0 1 44341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2817
timestamp 1626065694
transform 1 0 115328 0 1 45157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2816
timestamp 1626065694
transform 1 0 114784 0 1 42437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2815
timestamp 1626065694
transform 1 0 114240 0 1 44341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2814
timestamp 1626065694
transform 1 0 114240 0 1 46381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2813
timestamp 1626065694
transform 1 0 114240 0 1 46653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2812
timestamp 1626065694
transform 1 0 115192 0 1 43797
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2811
timestamp 1626065694
transform 1 0 112336 0 1 44613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2810
timestamp 1626065694
transform 1 0 112336 0 1 45021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2809
timestamp 1626065694
transform 1 0 114784 0 1 41893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2808
timestamp 1626065694
transform 1 0 116008 0 1 43253
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2807
timestamp 1626065694
transform 1 0 116008 0 1 43525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2806
timestamp 1626065694
transform 1 0 116008 0 1 43117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2805
timestamp 1626065694
transform 1 0 116008 0 1 42845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2804
timestamp 1626065694
transform 1 0 115192 0 1 43525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2803
timestamp 1626065694
transform 1 0 114376 0 1 44749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2802
timestamp 1626065694
transform 1 0 114784 0 1 43933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2801
timestamp 1626065694
transform 1 0 113696 0 1 45157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2800
timestamp 1626065694
transform 1 0 113696 0 1 45429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2799
timestamp 1626065694
transform 1 0 114784 0 1 44205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2798
timestamp 1626065694
transform 1 0 115464 0 1 46245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2797
timestamp 1626065694
transform 1 0 114376 0 1 45157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2796
timestamp 1626065694
transform 1 0 114376 0 1 45429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2795
timestamp 1626065694
transform 1 0 114784 0 1 45157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2794
timestamp 1626065694
transform 1 0 114240 0 1 44613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2793
timestamp 1626065694
transform 1 0 115872 0 1 41893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2792
timestamp 1626065694
transform 1 0 114784 0 1 45429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2791
timestamp 1626065694
transform 1 0 114648 0 1 45565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2790
timestamp 1626065694
transform 1 0 114648 0 1 45837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2789
timestamp 1626065694
transform 1 0 115328 0 1 41893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2788
timestamp 1626065694
transform 1 0 115464 0 1 45973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2787
timestamp 1626065694
transform 1 0 115192 0 1 41893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2786
timestamp 1626065694
transform 1 0 115192 0 1 46245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2785
timestamp 1626065694
transform 1 0 115192 0 1 45973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2784
timestamp 1626065694
transform 1 0 114240 0 1 42437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2783
timestamp 1626065694
transform 1 0 114240 0 1 42709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2782
timestamp 1626065694
transform 1 0 114376 0 1 45021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2781
timestamp 1626065694
transform 1 0 114784 0 1 42709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2780
timestamp 1626065694
transform 1 0 115872 0 1 44749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2779
timestamp 1626065694
transform 1 0 115872 0 1 45021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2778
timestamp 1626065694
transform 1 0 114376 0 1 43933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2777
timestamp 1626065694
transform 1 0 114376 0 1 44205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2776
timestamp 1626065694
transform 1 0 114376 0 1 43797
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2775
timestamp 1626065694
transform 1 0 115328 0 1 45973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2774
timestamp 1626065694
transform 1 0 114376 0 1 41893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2773
timestamp 1626065694
transform 1 0 115872 0 1 45157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2772
timestamp 1626065694
transform 1 0 115872 0 1 45429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2771
timestamp 1626065694
transform 1 0 115328 0 1 46245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2770
timestamp 1626065694
transform 1 0 114376 0 1 43525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2769
timestamp 1626065694
transform 1 0 114240 0 1 42029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2768
timestamp 1626065694
transform 1 0 114240 0 1 42301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2767
timestamp 1626065694
transform 1 0 115872 0 1 42709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2766
timestamp 1626065694
transform 1 0 115872 0 1 42437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2765
timestamp 1626065694
transform 1 0 114376 0 1 46245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2764
timestamp 1626065694
transform 1 0 115056 0 1 43117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2763
timestamp 1626065694
transform 1 0 114648 0 1 44749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2762
timestamp 1626065694
transform 1 0 115056 0 1 42845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2761
timestamp 1626065694
transform 1 0 116008 0 1 45565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2760
timestamp 1626065694
transform 1 0 116008 0 1 45837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2759
timestamp 1626065694
transform 1 0 114648 0 1 45021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2758
timestamp 1626065694
transform 1 0 114648 0 1 44613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2757
timestamp 1626065694
transform 1 0 114648 0 1 44341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2756
timestamp 1626065694
transform 1 0 115192 0 1 45157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2755
timestamp 1626065694
transform 1 0 116008 0 1 42301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2754
timestamp 1626065694
transform 1 0 116008 0 1 42029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2753
timestamp 1626065694
transform 1 0 114648 0 1 46381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2752
timestamp 1626065694
transform 1 0 114648 0 1 46653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2751
timestamp 1626065694
transform 1 0 114784 0 1 46245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2750
timestamp 1626065694
transform 1 0 114784 0 1 45973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2749
timestamp 1626065694
transform 1 0 114376 0 1 45973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2748
timestamp 1626065694
transform 1 0 115192 0 1 45429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2747
timestamp 1626065694
transform 1 0 114648 0 1 42029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2746
timestamp 1626065694
transform 1 0 114648 0 1 42301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2745
timestamp 1626065694
transform 1 0 115464 0 1 44613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2744
timestamp 1626065694
transform 1 0 115328 0 1 45429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2743
timestamp 1626065694
transform 1 0 116008 0 1 46381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2742
timestamp 1626065694
transform 1 0 114376 0 1 45837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2741
timestamp 1626065694
transform 1 0 114376 0 1 45565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2740
timestamp 1626065694
transform 1 0 116008 0 1 46653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2739
timestamp 1626065694
transform 1 0 115056 0 1 42029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2738
timestamp 1626065694
transform 1 0 115056 0 1 42301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2737
timestamp 1626065694
transform 1 0 115464 0 1 45565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2736
timestamp 1626065694
transform 1 0 115872 0 1 46245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2735
timestamp 1626065694
transform 1 0 115464 0 1 45837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2734
timestamp 1626065694
transform 1 0 115872 0 1 45973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2733
timestamp 1626065694
transform 1 0 114784 0 1 43797
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2732
timestamp 1626065694
transform 1 0 114784 0 1 43525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2731
timestamp 1626065694
transform 1 0 135320 0 1 48965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2730
timestamp 1626065694
transform 1 0 135320 0 1 47469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2729
timestamp 1626065694
transform 1 0 135320 0 1 50733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2728
timestamp 1626065694
transform 1 0 135320 0 1 42301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2727
timestamp 1626065694
transform 1 0 135320 0 1 45701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2726
timestamp 1626065694
transform 1 0 135320 0 1 43933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2725
timestamp 1626065694
transform 1 0 51272 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2724
timestamp 1626065694
transform 1 0 51272 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2723
timestamp 1626065694
transform 1 0 51272 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2722
timestamp 1626065694
transform 1 0 60792 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2721
timestamp 1626065694
transform 1 0 60792 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2720
timestamp 1626065694
transform 1 0 62696 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2719
timestamp 1626065694
transform 1 0 62696 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2718
timestamp 1626065694
transform 1 0 64192 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2717
timestamp 1626065694
transform 1 0 64192 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2716
timestamp 1626065694
transform 1 0 65824 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2715
timestamp 1626065694
transform 1 0 65824 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2714
timestamp 1626065694
transform 1 0 67592 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2713
timestamp 1626065694
transform 1 0 67592 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2712
timestamp 1626065694
transform 1 0 52632 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2711
timestamp 1626065694
transform 1 0 52632 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2710
timestamp 1626065694
transform 1 0 54128 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2709
timestamp 1626065694
transform 1 0 54128 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2708
timestamp 1626065694
transform 1 0 55896 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2707
timestamp 1626065694
transform 1 0 55896 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2706
timestamp 1626065694
transform 1 0 57664 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2705
timestamp 1626065694
transform 1 0 57664 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2704
timestamp 1626065694
transform 1 0 59160 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2703
timestamp 1626065694
transform 1 0 59160 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2702
timestamp 1626065694
transform 1 0 51408 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2701
timestamp 1626065694
transform 1 0 51408 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2700
timestamp 1626065694
transform 1 0 53720 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2699
timestamp 1626065694
transform 1 0 53720 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2698
timestamp 1626065694
transform 1 0 56304 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2697
timestamp 1626065694
transform 1 0 56304 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2696
timestamp 1626065694
transform 1 0 56168 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2695
timestamp 1626065694
transform 1 0 56168 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2694
timestamp 1626065694
transform 1 0 58752 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2693
timestamp 1626065694
transform 1 0 58752 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2692
timestamp 1626065694
transform 1 0 51408 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2691
timestamp 1626065694
transform 1 0 59432 0 1 75757
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2690
timestamp 1626065694
transform 1 0 51544 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2689
timestamp 1626065694
transform 1 0 51544 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2688
timestamp 1626065694
transform 1 0 53856 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2687
timestamp 1626065694
transform 1 0 53856 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2686
timestamp 1626065694
transform 1 0 53992 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2685
timestamp 1626065694
transform 1 0 53992 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2684
timestamp 1626065694
transform 1 0 56304 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2683
timestamp 1626065694
transform 1 0 56304 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2682
timestamp 1626065694
transform 1 0 56440 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2681
timestamp 1626065694
transform 1 0 56440 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2680
timestamp 1626065694
transform 1 0 58888 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2679
timestamp 1626065694
transform 1 0 58888 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2678
timestamp 1626065694
transform 1 0 59024 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2677
timestamp 1626065694
transform 1 0 59024 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2676
timestamp 1626065694
transform 1 0 53584 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2675
timestamp 1626065694
transform 1 0 56168 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2674
timestamp 1626065694
transform 1 0 58480 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2673
timestamp 1626065694
transform 1 0 61336 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2672
timestamp 1626065694
transform 1 0 61336 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2671
timestamp 1626065694
transform 1 0 63784 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2670
timestamp 1626065694
transform 1 0 61472 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2669
timestamp 1626065694
transform 1 0 61472 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2668
timestamp 1626065694
transform 1 0 61472 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2667
timestamp 1626065694
transform 1 0 61472 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2666
timestamp 1626065694
transform 1 0 63920 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2665
timestamp 1626065694
transform 1 0 63920 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2664
timestamp 1626065694
transform 1 0 63920 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2663
timestamp 1626065694
transform 1 0 63920 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2662
timestamp 1626065694
transform 1 0 66504 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2661
timestamp 1626065694
transform 1 0 66504 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2660
timestamp 1626065694
transform 1 0 66504 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2659
timestamp 1626065694
transform 1 0 66504 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2658
timestamp 1626065694
transform 1 0 63784 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2657
timestamp 1626065694
transform 1 0 66368 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2656
timestamp 1626065694
transform 1 0 66368 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2655
timestamp 1626065694
transform 1 0 60928 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2654
timestamp 1626065694
transform 1 0 63648 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2653
timestamp 1626065694
transform 1 0 66096 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2652
timestamp 1626065694
transform 1 0 50728 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2651
timestamp 1626065694
transform 1 0 50728 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2650
timestamp 1626065694
transform 1 0 44200 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2649
timestamp 1626065694
transform 1 0 44200 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2648
timestamp 1626065694
transform 1 0 49232 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2647
timestamp 1626065694
transform 1 0 49232 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2646
timestamp 1626065694
transform 1 0 45696 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2645
timestamp 1626065694
transform 1 0 45696 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2644
timestamp 1626065694
transform 1 0 47464 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2643
timestamp 1626065694
transform 1 0 47464 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2642
timestamp 1626065694
transform 1 0 37536 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2641
timestamp 1626065694
transform 1 0 37536 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2640
timestamp 1626065694
transform 1 0 39168 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2639
timestamp 1626065694
transform 1 0 39168 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2638
timestamp 1626065694
transform 1 0 40664 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2637
timestamp 1626065694
transform 1 0 40664 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2636
timestamp 1626065694
transform 1 0 42432 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2635
timestamp 1626065694
transform 1 0 42432 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2634
timestamp 1626065694
transform 1 0 35632 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2633
timestamp 1626065694
transform 1 0 35632 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2632
timestamp 1626065694
transform 1 0 38896 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2631
timestamp 1626065694
transform 1 0 38896 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2630
timestamp 1626065694
transform 1 0 39032 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2629
timestamp 1626065694
transform 1 0 41480 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2628
timestamp 1626065694
transform 1 0 41480 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2627
timestamp 1626065694
transform 1 0 41480 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2626
timestamp 1626065694
transform 1 0 41344 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2625
timestamp 1626065694
transform 1 0 41344 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2624
timestamp 1626065694
transform 1 0 41480 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2623
timestamp 1626065694
transform 1 0 36448 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2622
timestamp 1626065694
transform 1 0 36448 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2621
timestamp 1626065694
transform 1 0 36448 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2620
timestamp 1626065694
transform 1 0 36448 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2619
timestamp 1626065694
transform 1 0 36176 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2618
timestamp 1626065694
transform 1 0 38488 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2617
timestamp 1626065694
transform 1 0 41072 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2616
timestamp 1626065694
transform 1 0 39032 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2615
timestamp 1626065694
transform 1 0 36312 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2614
timestamp 1626065694
transform 1 0 36312 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2613
timestamp 1626065694
transform 1 0 38624 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2612
timestamp 1626065694
transform 1 0 38624 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2611
timestamp 1626065694
transform 1 0 39032 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2610
timestamp 1626065694
transform 1 0 39032 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2609
timestamp 1626065694
transform 1 0 48688 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2608
timestamp 1626065694
transform 1 0 43656 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2607
timestamp 1626065694
transform 1 0 43656 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2606
timestamp 1626065694
transform 1 0 43928 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2605
timestamp 1626065694
transform 1 0 43928 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2604
timestamp 1626065694
transform 1 0 43928 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2603
timestamp 1626065694
transform 1 0 43792 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2602
timestamp 1626065694
transform 1 0 44064 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2601
timestamp 1626065694
transform 1 0 44064 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2600
timestamp 1626065694
transform 1 0 46512 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2599
timestamp 1626065694
transform 1 0 46512 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2598
timestamp 1626065694
transform 1 0 46512 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2597
timestamp 1626065694
transform 1 0 43520 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2596
timestamp 1626065694
transform 1 0 46104 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2595
timestamp 1626065694
transform 1 0 48552 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2594
timestamp 1626065694
transform 1 0 51136 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2593
timestamp 1626065694
transform 1 0 46512 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2592
timestamp 1626065694
transform 1 0 48960 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2591
timestamp 1626065694
transform 1 0 46376 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2590
timestamp 1626065694
transform 1 0 46376 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2589
timestamp 1626065694
transform 1 0 48960 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2588
timestamp 1626065694
transform 1 0 48960 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2587
timestamp 1626065694
transform 1 0 48960 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2586
timestamp 1626065694
transform 1 0 48688 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2585
timestamp 1626065694
transform 1 0 45696 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2584
timestamp 1626065694
transform 1 0 34952 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2583
timestamp 1626065694
transform 1 0 34952 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2582
timestamp 1626065694
transform 1 0 46240 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2581
timestamp 1626065694
transform 1 0 46240 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2580
timestamp 1626065694
transform 1 0 39984 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2579
timestamp 1626065694
transform 1 0 39984 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2578
timestamp 1626065694
transform 1 0 46920 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2577
timestamp 1626065694
transform 1 0 46920 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2576
timestamp 1626065694
transform 1 0 40664 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2575
timestamp 1626065694
transform 1 0 40664 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2574
timestamp 1626065694
transform 1 0 48688 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2573
timestamp 1626065694
transform 1 0 48688 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2572
timestamp 1626065694
transform 1 0 35768 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2571
timestamp 1626065694
transform 1 0 35768 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2570
timestamp 1626065694
transform 1 0 41208 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2569
timestamp 1626065694
transform 1 0 41208 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2568
timestamp 1626065694
transform 1 0 49912 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2567
timestamp 1626065694
transform 1 0 49912 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2566
timestamp 1626065694
transform 1 0 50728 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2565
timestamp 1626065694
transform 1 0 50728 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2564
timestamp 1626065694
transform 1 0 36992 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2563
timestamp 1626065694
transform 1 0 36992 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2562
timestamp 1626065694
transform 1 0 34408 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2561
timestamp 1626065694
transform 1 0 34408 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2560
timestamp 1626065694
transform 1 0 41888 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2559
timestamp 1626065694
transform 1 0 41888 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2558
timestamp 1626065694
transform 1 0 42432 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2557
timestamp 1626065694
transform 1 0 42432 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2556
timestamp 1626065694
transform 1 0 37536 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2555
timestamp 1626065694
transform 1 0 37536 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2554
timestamp 1626065694
transform 1 0 43248 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2553
timestamp 1626065694
transform 1 0 43248 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2552
timestamp 1626065694
transform 1 0 38216 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2551
timestamp 1626065694
transform 1 0 38216 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2550
timestamp 1626065694
transform 1 0 36176 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2549
timestamp 1626065694
transform 1 0 36176 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2548
timestamp 1626065694
transform 1 0 44608 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2547
timestamp 1626065694
transform 1 0 44608 0 1 70861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2546
timestamp 1626065694
transform 1 0 45696 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2545
timestamp 1626065694
transform 1 0 61880 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2544
timestamp 1626065694
transform 1 0 61880 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2543
timestamp 1626065694
transform 1 0 62424 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2542
timestamp 1626065694
transform 1 0 62424 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2541
timestamp 1626065694
transform 1 0 53176 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2540
timestamp 1626065694
transform 1 0 57392 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2539
timestamp 1626065694
transform 1 0 63104 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2538
timestamp 1626065694
transform 1 0 63104 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2537
timestamp 1626065694
transform 1 0 63648 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2536
timestamp 1626065694
transform 1 0 63648 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2535
timestamp 1626065694
transform 1 0 57392 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2534
timestamp 1626065694
transform 1 0 53312 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2533
timestamp 1626065694
transform 1 0 53312 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2532
timestamp 1626065694
transform 1 0 58616 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2531
timestamp 1626065694
transform 1 0 65008 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2530
timestamp 1626065694
transform 1 0 65008 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2529
timestamp 1626065694
transform 1 0 58616 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2528
timestamp 1626065694
transform 1 0 54400 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2527
timestamp 1626065694
transform 1 0 66096 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2526
timestamp 1626065694
transform 1 0 66096 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2525
timestamp 1626065694
transform 1 0 54400 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2524
timestamp 1626065694
transform 1 0 54944 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2523
timestamp 1626065694
transform 1 0 66912 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2522
timestamp 1626065694
transform 1 0 66912 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2521
timestamp 1626065694
transform 1 0 67456 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2520
timestamp 1626065694
transform 1 0 67456 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2519
timestamp 1626065694
transform 1 0 59432 0 1 71541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2518
timestamp 1626065694
transform 1 0 54944 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2517
timestamp 1626065694
transform 1 0 68136 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2516
timestamp 1626065694
transform 1 0 68136 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2515
timestamp 1626065694
transform 1 0 56032 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2514
timestamp 1626065694
transform 1 0 59432 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2513
timestamp 1626065694
transform 1 0 59432 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2512
timestamp 1626065694
transform 1 0 59976 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2511
timestamp 1626065694
transform 1 0 59976 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2510
timestamp 1626065694
transform 1 0 56032 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2509
timestamp 1626065694
transform 1 0 52496 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2508
timestamp 1626065694
transform 1 0 61200 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2507
timestamp 1626065694
transform 1 0 61200 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2506
timestamp 1626065694
transform 1 0 52496 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2505
timestamp 1626065694
transform 1 0 53176 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2504
timestamp 1626065694
transform 1 0 1224 0 1 72629
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2503
timestamp 1626065694
transform 1 0 27200 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2502
timestamp 1626065694
transform 1 0 27200 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2501
timestamp 1626065694
transform 1 0 28968 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2500
timestamp 1626065694
transform 1 0 28968 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2499
timestamp 1626065694
transform 1 0 30600 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2498
timestamp 1626065694
transform 1 0 30600 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2497
timestamp 1626065694
transform 1 0 32368 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2496
timestamp 1626065694
transform 1 0 32368 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2495
timestamp 1626065694
transform 1 0 34136 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2494
timestamp 1626065694
transform 1 0 34136 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2493
timestamp 1626065694
transform 1 0 25704 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2492
timestamp 1626065694
transform 1 0 25704 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2491
timestamp 1626065694
transform 1 0 23936 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2490
timestamp 1626065694
transform 1 0 22168 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2489
timestamp 1626065694
transform 1 0 22168 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2488
timestamp 1626065694
transform 1 0 23936 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2487
timestamp 1626065694
transform 1 0 18904 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2486
timestamp 1626065694
transform 1 0 18904 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2485
timestamp 1626065694
transform 1 0 20672 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2484
timestamp 1626065694
transform 1 0 20672 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2483
timestamp 1626065694
transform 1 0 28832 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2482
timestamp 1626065694
transform 1 0 28968 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2481
timestamp 1626065694
transform 1 0 28968 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2480
timestamp 1626065694
transform 1 0 31416 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2479
timestamp 1626065694
transform 1 0 31416 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2478
timestamp 1626065694
transform 1 0 31552 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2477
timestamp 1626065694
transform 1 0 31552 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2476
timestamp 1626065694
transform 1 0 34000 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2475
timestamp 1626065694
transform 1 0 34000 0 1 75213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2474
timestamp 1626065694
transform 1 0 34000 0 1 75077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2473
timestamp 1626065694
transform 1 0 34000 0 1 73173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2472
timestamp 1626065694
transform 1 0 28968 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2471
timestamp 1626065694
transform 1 0 28968 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2470
timestamp 1626065694
transform 1 0 33728 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2469
timestamp 1626065694
transform 1 0 33728 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2468
timestamp 1626065694
transform 1 0 31280 0 1 75893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2467
timestamp 1626065694
transform 1 0 31280 0 1 76573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2466
timestamp 1626065694
transform 1 0 28968 0 1 73037
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2465
timestamp 1626065694
transform 1 0 28968 0 1 76981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2464
timestamp 1626065694
transform 1 0 28696 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2463
timestamp 1626065694
transform 1 0 31008 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2462
timestamp 1626065694
transform 1 0 33456 0 1 77117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2461
timestamp 1626065694
transform 1 0 8704 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2460
timestamp 1626065694
transform 1 0 8704 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2459
timestamp 1626065694
transform 1 0 10472 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2458
timestamp 1626065694
transform 1 0 10472 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2457
timestamp 1626065694
transform 1 0 12104 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2456
timestamp 1626065694
transform 1 0 12104 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2455
timestamp 1626065694
transform 1 0 14008 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2454
timestamp 1626065694
transform 1 0 14008 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2453
timestamp 1626065694
transform 1 0 15640 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2452
timestamp 1626065694
transform 1 0 15640 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2451
timestamp 1626065694
transform 1 0 17136 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2450
timestamp 1626065694
transform 1 0 17136 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2449
timestamp 1626065694
transform 1 0 5440 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2448
timestamp 1626065694
transform 1 0 5440 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2447
timestamp 1626065694
transform 1 0 7208 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2446
timestamp 1626065694
transform 1 0 7208 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2445
timestamp 1626065694
transform 1 0 2040 0 1 81061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2444
timestamp 1626065694
transform 1 0 2040 0 1 81333
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2443
timestamp 1626065694
transform 1 0 2176 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2442
timestamp 1626065694
transform 1 0 2176 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2441
timestamp 1626065694
transform 1 0 3944 0 1 81469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2440
timestamp 1626065694
transform 1 0 3944 0 1 82013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2439
timestamp 1626065694
transform 1 0 1224 0 1 79429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2438
timestamp 1626065694
transform 1 0 1224 0 1 77525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2437
timestamp 1626065694
transform 1 0 1224 0 1 76029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2436
timestamp 1626065694
transform 1 0 1224 0 1 74125
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2435
timestamp 1626065694
transform 1 0 1224 0 1 67461
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2434
timestamp 1626065694
transform 1 0 1224 0 1 69229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2433
timestamp 1626065694
transform 1 0 1224 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2432
timestamp 1626065694
transform 1 0 1224 0 1 65965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2431
timestamp 1626065694
transform 1 0 1224 0 1 62565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2430
timestamp 1626065694
transform 1 0 1224 0 1 64061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2429
timestamp 1626065694
transform 1 0 31280 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2428
timestamp 1626065694
transform 1 0 28968 0 1 70725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2427
timestamp 1626065694
transform 1 0 27472 0 1 67869
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2426
timestamp 1626065694
transform 1 0 27472 0 1 68141
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2425
timestamp 1626065694
transform 1 0 27336 0 1 67869
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2424
timestamp 1626065694
transform 1 0 27336 0 1 67597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2423
timestamp 1626065694
transform 1 0 31960 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2422
timestamp 1626065694
transform 1 0 31960 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2421
timestamp 1626065694
transform 1 0 32504 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2420
timestamp 1626065694
transform 1 0 32504 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2419
timestamp 1626065694
transform 1 0 33728 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2418
timestamp 1626065694
transform 1 0 33728 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2417
timestamp 1626065694
transform 1 0 28560 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2416
timestamp 1626065694
transform 1 0 28560 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2415
timestamp 1626065694
transform 1 0 28696 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2414
timestamp 1626065694
transform 1 0 28696 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2413
timestamp 1626065694
transform 1 0 29784 0 1 70997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2412
timestamp 1626065694
transform 1 0 29784 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2411
timestamp 1626065694
transform 1 0 31280 0 1 71405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2410
timestamp 1626065694
transform 1 0 21624 0 1 67597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2409
timestamp 1626065694
transform 1 0 21760 0 1 68821
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2408
timestamp 1626065694
transform 1 0 21760 0 1 69093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2407
timestamp 1626065694
transform 1 0 21624 0 1 69229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2406
timestamp 1626065694
transform 1 0 21624 0 1 69501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2405
timestamp 1626065694
transform 1 0 22168 0 1 69637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2404
timestamp 1626065694
transform 1 0 22168 0 1 69909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2403
timestamp 1626065694
transform 1 0 20808 0 1 69501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2402
timestamp 1626065694
transform 1 0 20808 0 1 69229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2401
timestamp 1626065694
transform 1 0 20808 0 1 68821
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2400
timestamp 1626065694
transform 1 0 20808 0 1 68549
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2399
timestamp 1626065694
transform 1 0 20808 0 1 67597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2398
timestamp 1626065694
transform 1 0 22440 0 1 68413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2397
timestamp 1626065694
transform 1 0 22440 0 1 68685
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2396
timestamp 1626065694
transform 1 0 20808 0 1 68005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2395
timestamp 1626065694
transform 1 0 20808 0 1 67733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2394
timestamp 1626065694
transform 1 0 22032 0 1 69093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2393
timestamp 1626065694
transform 1 0 22032 0 1 68821
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2392
timestamp 1626065694
transform 1 0 22168 0 1 69229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2391
timestamp 1626065694
transform 1 0 22168 0 1 69501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2390
timestamp 1626065694
transform 1 0 22440 0 1 69637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2389
timestamp 1626065694
transform 1 0 22440 0 1 69909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2388
timestamp 1626065694
transform 1 0 22440 0 1 69501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2387
timestamp 1626065694
transform 1 0 22440 0 1 69229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2386
timestamp 1626065694
transform 1 0 22032 0 1 68685
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2385
timestamp 1626065694
transform 1 0 22032 0 1 68413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2384
timestamp 1626065694
transform 1 0 21216 0 1 67597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2383
timestamp 1626065694
transform 1 0 21352 0 1 69501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2382
timestamp 1626065694
transform 1 0 21352 0 1 69229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2381
timestamp 1626065694
transform 1 0 21896 0 1 68005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2380
timestamp 1626065694
transform 1 0 22440 0 1 69093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2379
timestamp 1626065694
transform 1 0 22440 0 1 68821
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2378
timestamp 1626065694
transform 1 0 21896 0 1 68277
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2377
timestamp 1626065694
transform 1 0 20808 0 1 62565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2376
timestamp 1626065694
transform 1 0 21352 0 1 66373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2375
timestamp 1626065694
transform 1 0 21352 0 1 66101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2374
timestamp 1626065694
transform 1 0 21488 0 1 66373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2373
timestamp 1626065694
transform 1 0 21488 0 1 66101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2372
timestamp 1626065694
transform 1 0 21216 0 1 67325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2371
timestamp 1626065694
transform 1 0 20808 0 1 62973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2370
timestamp 1626065694
transform 1 0 21488 0 1 67189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2369
timestamp 1626065694
transform 1 0 21488 0 1 66917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2368
timestamp 1626065694
transform 1 0 21216 0 1 62429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2367
timestamp 1626065694
transform 1 0 20808 0 1 63245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2366
timestamp 1626065694
transform 1 0 20808 0 1 63653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2365
timestamp 1626065694
transform 1 0 20808 0 1 63381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2364
timestamp 1626065694
transform 1 0 20808 0 1 62429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2363
timestamp 1626065694
transform 1 0 22032 0 1 62429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2362
timestamp 1626065694
transform 1 0 21760 0 1 65965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2361
timestamp 1626065694
transform 1 0 21760 0 1 65693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2360
timestamp 1626065694
transform 1 0 21896 0 1 63653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2359
timestamp 1626065694
transform 1 0 21896 0 1 63381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2358
timestamp 1626065694
transform 1 0 21760 0 1 64061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2357
timestamp 1626065694
transform 1 0 21760 0 1 64333
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2356
timestamp 1626065694
transform 1 0 21624 0 1 67325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2355
timestamp 1626065694
transform 1 0 20808 0 1 66917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2354
timestamp 1626065694
transform 1 0 20808 0 1 67189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2353
timestamp 1626065694
transform 1 0 20808 0 1 66781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2352
timestamp 1626065694
transform 1 0 20808 0 1 66509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2351
timestamp 1626065694
transform 1 0 20944 0 1 66101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2350
timestamp 1626065694
transform 1 0 21624 0 1 66781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2349
timestamp 1626065694
transform 1 0 21624 0 1 66509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2348
timestamp 1626065694
transform 1 0 21896 0 1 65149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2347
timestamp 1626065694
transform 1 0 21896 0 1 64877
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2346
timestamp 1626065694
transform 1 0 21760 0 1 62837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2345
timestamp 1626065694
transform 1 0 22032 0 1 62565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2344
timestamp 1626065694
transform 1 0 22032 0 1 62837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2343
timestamp 1626065694
transform 1 0 22032 0 1 65557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2342
timestamp 1626065694
transform 1 0 22032 0 1 65285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2341
timestamp 1626065694
transform 1 0 22032 0 1 65693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2340
timestamp 1626065694
transform 1 0 22032 0 1 65965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2339
timestamp 1626065694
transform 1 0 21760 0 1 62565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2338
timestamp 1626065694
transform 1 0 20944 0 1 66373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2337
timestamp 1626065694
transform 1 0 22576 0 1 62429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2336
timestamp 1626065694
transform 1 0 20808 0 1 64061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2335
timestamp 1626065694
transform 1 0 22576 0 1 65965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2334
timestamp 1626065694
transform 1 0 20808 0 1 67325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2333
timestamp 1626065694
transform 1 0 20808 0 1 63789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2332
timestamp 1626065694
transform 1 0 22032 0 1 65013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2331
timestamp 1626065694
transform 1 0 22032 0 1 64469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2330
timestamp 1626065694
transform 1 0 22576 0 1 65693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2329
timestamp 1626065694
transform 1 0 22576 0 1 66101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2328
timestamp 1626065694
transform 1 0 22576 0 1 66373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2327
timestamp 1626065694
transform 1 0 22440 0 1 62565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2326
timestamp 1626065694
transform 1 0 22440 0 1 62837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2325
timestamp 1626065694
transform 1 0 22576 0 1 64469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2324
timestamp 1626065694
transform 1 0 22576 0 1 64741
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2323
timestamp 1626065694
transform 1 0 22032 0 1 63245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2322
timestamp 1626065694
transform 1 0 22032 0 1 62973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2321
timestamp 1626065694
transform 1 0 22576 0 1 63245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2320
timestamp 1626065694
transform 1 0 22576 0 1 62973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2319
timestamp 1626065694
transform 1 0 21624 0 1 62429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2318
timestamp 1626065694
transform 1 0 22032 0 1 66509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2317
timestamp 1626065694
transform 1 0 22032 0 1 66781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2316
timestamp 1626065694
transform 1 0 22440 0 1 66917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2315
timestamp 1626065694
transform 1 0 22440 0 1 67189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2314
timestamp 1626065694
transform 1 0 22168 0 1 66373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2313
timestamp 1626065694
transform 1 0 22168 0 1 66101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2312
timestamp 1626065694
transform 1 0 22168 0 1 64877
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2311
timestamp 1626065694
transform 1 0 22168 0 1 65149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2310
timestamp 1626065694
transform 1 0 22440 0 1 66781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2309
timestamp 1626065694
transform 1 0 22440 0 1 66509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2308
timestamp 1626065694
transform 1 0 22168 0 1 64741
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2307
timestamp 1626065694
transform 1 0 22168 0 1 64469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2306
timestamp 1626065694
transform 1 0 20944 0 1 65557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2305
timestamp 1626065694
transform 1 0 20944 0 1 65285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2304
timestamp 1626065694
transform 1 0 20808 0 1 65693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2303
timestamp 1626065694
transform 1 0 20808 0 1 65965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2302
timestamp 1626065694
transform 1 0 22032 0 1 66917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2301
timestamp 1626065694
transform 1 0 22032 0 1 67189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2300
timestamp 1626065694
transform 1 0 22440 0 1 65285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2299
timestamp 1626065694
transform 1 0 22440 0 1 65557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2298
timestamp 1626065694
transform 1 0 22440 0 1 65149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2297
timestamp 1626065694
transform 1 0 22440 0 1 64877
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2296
timestamp 1626065694
transform 1 0 20808 0 1 62837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2295
timestamp 1626065694
transform 1 0 21352 0 1 65285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2294
timestamp 1626065694
transform 1 0 21352 0 1 65557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2293
timestamp 1626065694
transform 1 0 21488 0 1 65285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2292
timestamp 1626065694
transform 1 0 21488 0 1 65557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2291
timestamp 1626065694
transform 1 0 27608 0 1 64741
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2290
timestamp 1626065694
transform 1 0 27472 0 1 63517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2289
timestamp 1626065694
transform 1 0 27472 0 1 63789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2288
timestamp 1626065694
transform 1 0 27336 0 1 64197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2287
timestamp 1626065694
transform 1 0 27336 0 1 64469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2286
timestamp 1626065694
transform 1 0 27608 0 1 64197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2285
timestamp 1626065694
transform 1 0 27608 0 1 63925
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2284
timestamp 1626065694
transform 1 0 27608 0 1 65013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2283
timestamp 1626065694
transform 1 0 20808 0 1 51957
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2282
timestamp 1626065694
transform 1 0 27336 0 1 59573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2281
timestamp 1626065694
transform 1 0 27336 0 1 59845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2280
timestamp 1626065694
transform 1 0 27608 0 1 58621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2279
timestamp 1626065694
transform 1 0 27608 0 1 58349
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2278
timestamp 1626065694
transform 1 0 22168 0 1 60797
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2277
timestamp 1626065694
transform 1 0 22168 0 1 60525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2276
timestamp 1626065694
transform 1 0 22168 0 1 60933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2275
timestamp 1626065694
transform 1 0 22168 0 1 61205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2274
timestamp 1626065694
transform 1 0 22168 0 1 58485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2273
timestamp 1626065694
transform 1 0 22168 0 1 58213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2272
timestamp 1626065694
transform 1 0 22168 0 1 58621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2271
timestamp 1626065694
transform 1 0 22168 0 1 58893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2270
timestamp 1626065694
transform 1 0 22032 0 1 60389
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2269
timestamp 1626065694
transform 1 0 22032 0 1 60117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2268
timestamp 1626065694
transform 1 0 22032 0 1 58077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2267
timestamp 1626065694
transform 1 0 22032 0 1 57805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2266
timestamp 1626065694
transform 1 0 22032 0 1 62157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2265
timestamp 1626065694
transform 1 0 22168 0 1 57669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2264
timestamp 1626065694
transform 1 0 22168 0 1 57397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2263
timestamp 1626065694
transform 1 0 22168 0 1 62021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2262
timestamp 1626065694
transform 1 0 22168 0 1 61749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2261
timestamp 1626065694
transform 1 0 22032 0 1 57261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2260
timestamp 1626065694
transform 1 0 22032 0 1 61341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2259
timestamp 1626065694
transform 1 0 22032 0 1 61613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2258
timestamp 1626065694
transform 1 0 20808 0 1 58213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2257
timestamp 1626065694
transform 1 0 20808 0 1 58485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2256
timestamp 1626065694
transform 1 0 22032 0 1 59301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2255
timestamp 1626065694
transform 1 0 22032 0 1 59029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2254
timestamp 1626065694
transform 1 0 21216 0 1 57261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2253
timestamp 1626065694
transform 1 0 22440 0 1 61341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2252
timestamp 1626065694
transform 1 0 22440 0 1 61613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2251
timestamp 1626065694
transform 1 0 22440 0 1 61205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2250
timestamp 1626065694
transform 1 0 22440 0 1 60933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2249
timestamp 1626065694
transform 1 0 22440 0 1 59301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2248
timestamp 1626065694
transform 1 0 22440 0 1 59029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2247
timestamp 1626065694
transform 1 0 22440 0 1 62021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2246
timestamp 1626065694
transform 1 0 22440 0 1 61749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2245
timestamp 1626065694
transform 1 0 22576 0 1 62157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2244
timestamp 1626065694
transform 1 0 22440 0 1 57261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2243
timestamp 1626065694
transform 1 0 22576 0 1 57397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2242
timestamp 1626065694
transform 1 0 22576 0 1 57669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2241
timestamp 1626065694
transform 1 0 22440 0 1 58485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2240
timestamp 1626065694
transform 1 0 22440 0 1 58213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2239
timestamp 1626065694
transform 1 0 22440 0 1 58621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2238
timestamp 1626065694
transform 1 0 22440 0 1 58893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2237
timestamp 1626065694
transform 1 0 21488 0 1 57805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2236
timestamp 1626065694
transform 1 0 21488 0 1 58077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2235
timestamp 1626065694
transform 1 0 22440 0 1 58077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2234
timestamp 1626065694
transform 1 0 22440 0 1 57805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2233
timestamp 1626065694
transform 1 0 22576 0 1 60525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2232
timestamp 1626065694
transform 1 0 22576 0 1 60797
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2231
timestamp 1626065694
transform 1 0 22440 0 1 60389
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2230
timestamp 1626065694
transform 1 0 22440 0 1 60117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2229
timestamp 1626065694
transform 1 0 21216 0 1 62157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2228
timestamp 1626065694
transform 1 0 21352 0 1 60933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2227
timestamp 1626065694
transform 1 0 21352 0 1 61205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2226
timestamp 1626065694
transform 1 0 21352 0 1 58485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2225
timestamp 1626065694
transform 1 0 21352 0 1 58213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2224
timestamp 1626065694
transform 1 0 21352 0 1 61749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2223
timestamp 1626065694
transform 1 0 21352 0 1 62021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2222
timestamp 1626065694
transform 1 0 21760 0 1 61613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2221
timestamp 1626065694
transform 1 0 21760 0 1 61341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2220
timestamp 1626065694
transform 1 0 21760 0 1 58485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2219
timestamp 1626065694
transform 1 0 21760 0 1 58213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2218
timestamp 1626065694
transform 1 0 21760 0 1 59709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2217
timestamp 1626065694
transform 1 0 21760 0 1 59437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2216
timestamp 1626065694
transform 1 0 21896 0 1 60389
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2215
timestamp 1626065694
transform 1 0 21896 0 1 60117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2214
timestamp 1626065694
transform 1 0 21760 0 1 57261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2213
timestamp 1626065694
transform 1 0 21216 0 1 58893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2212
timestamp 1626065694
transform 1 0 21624 0 1 62157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2211
timestamp 1626065694
transform 1 0 21216 0 1 58621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2210
timestamp 1626065694
transform 1 0 20808 0 1 59709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2209
timestamp 1626065694
transform 1 0 20808 0 1 59437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2208
timestamp 1626065694
transform 1 0 20808 0 1 59845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2207
timestamp 1626065694
transform 1 0 20808 0 1 60117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2206
timestamp 1626065694
transform 1 0 20808 0 1 57669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2205
timestamp 1626065694
transform 1 0 20808 0 1 57397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2204
timestamp 1626065694
transform 1 0 20944 0 1 57805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2203
timestamp 1626065694
transform 1 0 20944 0 1 58077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2202
timestamp 1626065694
transform 1 0 20808 0 1 59301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2201
timestamp 1626065694
transform 1 0 20808 0 1 59029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2200
timestamp 1626065694
transform 1 0 20808 0 1 62157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2199
timestamp 1626065694
transform 1 0 20944 0 1 61749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2198
timestamp 1626065694
transform 1 0 20944 0 1 62021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2197
timestamp 1626065694
transform 1 0 20944 0 1 61613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2196
timestamp 1626065694
transform 1 0 20944 0 1 61341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2195
timestamp 1626065694
transform 1 0 20808 0 1 58621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2194
timestamp 1626065694
transform 1 0 20808 0 1 58893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2193
timestamp 1626065694
transform 1 0 21216 0 1 52909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2192
timestamp 1626065694
transform 1 0 22168 0 1 56445
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2191
timestamp 1626065694
transform 1 0 22168 0 1 56173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2190
timestamp 1626065694
transform 1 0 22032 0 1 54677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2189
timestamp 1626065694
transform 1 0 22032 0 1 54949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2188
timestamp 1626065694
transform 1 0 22576 0 1 54541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2187
timestamp 1626065694
transform 1 0 22576 0 1 54269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2186
timestamp 1626065694
transform 1 0 22168 0 1 53861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2185
timestamp 1626065694
transform 1 0 22168 0 1 54269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2184
timestamp 1626065694
transform 1 0 22168 0 1 54541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2183
timestamp 1626065694
transform 1 0 20944 0 1 56173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2182
timestamp 1626065694
transform 1 0 22440 0 1 56445
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2181
timestamp 1626065694
transform 1 0 22440 0 1 56173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2180
timestamp 1626065694
transform 1 0 21352 0 1 56173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2179
timestamp 1626065694
transform 1 0 22440 0 1 53317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2178
timestamp 1626065694
transform 1 0 22440 0 1 53045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2177
timestamp 1626065694
transform 1 0 22576 0 1 52093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2176
timestamp 1626065694
transform 1 0 21352 0 1 56445
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2175
timestamp 1626065694
transform 1 0 21216 0 1 56989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2174
timestamp 1626065694
transform 1 0 20944 0 1 55901
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2173
timestamp 1626065694
transform 1 0 22440 0 1 54949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2172
timestamp 1626065694
transform 1 0 22440 0 1 54677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2171
timestamp 1626065694
transform 1 0 22576 0 1 52637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2170
timestamp 1626065694
transform 1 0 22576 0 1 52909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2169
timestamp 1626065694
transform 1 0 22440 0 1 52501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2168
timestamp 1626065694
transform 1 0 21488 0 1 55493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2167
timestamp 1626065694
transform 1 0 21488 0 1 55765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2166
timestamp 1626065694
transform 1 0 21624 0 1 56173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2165
timestamp 1626065694
transform 1 0 21624 0 1 56445
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2164
timestamp 1626065694
transform 1 0 22440 0 1 52229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2163
timestamp 1626065694
transform 1 0 20808 0 1 55765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2162
timestamp 1626065694
transform 1 0 22168 0 1 52093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2161
timestamp 1626065694
transform 1 0 22168 0 1 52229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2160
timestamp 1626065694
transform 1 0 22168 0 1 52501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2159
timestamp 1626065694
transform 1 0 20808 0 1 52229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2158
timestamp 1626065694
transform 1 0 21624 0 1 54677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2157
timestamp 1626065694
transform 1 0 21624 0 1 54949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2156
timestamp 1626065694
transform 1 0 21352 0 1 53317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2155
timestamp 1626065694
transform 1 0 22168 0 1 52909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2154
timestamp 1626065694
transform 1 0 22168 0 1 52637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2153
timestamp 1626065694
transform 1 0 21352 0 1 53045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2152
timestamp 1626065694
transform 1 0 21488 0 1 53317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2151
timestamp 1626065694
transform 1 0 22168 0 1 53045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2150
timestamp 1626065694
transform 1 0 21760 0 1 56989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2149
timestamp 1626065694
transform 1 0 21488 0 1 53045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2148
timestamp 1626065694
transform 1 0 21760 0 1 54133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2147
timestamp 1626065694
transform 1 0 21760 0 1 53861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2146
timestamp 1626065694
transform 1 0 21760 0 1 52909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2145
timestamp 1626065694
transform 1 0 21760 0 1 52637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2144
timestamp 1626065694
transform 1 0 22032 0 1 56989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2143
timestamp 1626065694
transform 1 0 21352 0 1 54269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2142
timestamp 1626065694
transform 1 0 22440 0 1 56989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2141
timestamp 1626065694
transform 1 0 21624 0 1 53453
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2140
timestamp 1626065694
transform 1 0 21624 0 1 53725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2139
timestamp 1626065694
transform 1 0 20944 0 1 55085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2138
timestamp 1626065694
transform 1 0 20944 0 1 55357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2137
timestamp 1626065694
transform 1 0 20808 0 1 54949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2136
timestamp 1626065694
transform 1 0 20808 0 1 54677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2135
timestamp 1626065694
transform 1 0 20808 0 1 54133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2134
timestamp 1626065694
transform 1 0 20808 0 1 53861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2133
timestamp 1626065694
transform 1 0 20944 0 1 54269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2132
timestamp 1626065694
transform 1 0 20944 0 1 54541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2131
timestamp 1626065694
transform 1 0 22168 0 1 53317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2130
timestamp 1626065694
transform 1 0 22440 0 1 56853
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2129
timestamp 1626065694
transform 1 0 22440 0 1 56581
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2128
timestamp 1626065694
transform 1 0 22032 0 1 56853
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2127
timestamp 1626065694
transform 1 0 22032 0 1 56581
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2126
timestamp 1626065694
transform 1 0 22440 0 1 53861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2125
timestamp 1626065694
transform 1 0 22440 0 1 54133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2124
timestamp 1626065694
transform 1 0 22440 0 1 53725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2123
timestamp 1626065694
transform 1 0 20944 0 1 52909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2122
timestamp 1626065694
transform 1 0 20944 0 1 52637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2121
timestamp 1626065694
transform 1 0 22440 0 1 53453
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2120
timestamp 1626065694
transform 1 0 22032 0 1 53725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2119
timestamp 1626065694
transform 1 0 22032 0 1 53453
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2118
timestamp 1626065694
transform 1 0 20808 0 1 53725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2117
timestamp 1626065694
transform 1 0 20808 0 1 53453
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2116
timestamp 1626065694
transform 1 0 20808 0 1 55493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2115
timestamp 1626065694
transform 1 0 22168 0 1 54133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2114
timestamp 1626065694
transform 1 0 21352 0 1 54541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2113
timestamp 1626065694
transform 1 0 21488 0 1 54269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2112
timestamp 1626065694
transform 1 0 21488 0 1 54541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2111
timestamp 1626065694
transform 1 0 21216 0 1 52637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2110
timestamp 1626065694
transform 1 0 27472 0 1 55493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2109
timestamp 1626065694
transform 1 0 27472 0 1 52365
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2108
timestamp 1626065694
transform 1 0 27472 0 1 52093
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2107
timestamp 1626065694
transform 1 0 27608 0 1 55493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2106
timestamp 1626065694
transform 1 0 27608 0 1 55221
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2105
timestamp 1626065694
transform 1 0 27472 0 1 55901
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2104
timestamp 1626065694
transform 1 0 1224 0 1 57533
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2103
timestamp 1626065694
transform 1 0 1224 0 1 60933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2102
timestamp 1626065694
transform 1 0 1224 0 1 59165
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2101
timestamp 1626065694
transform 1 0 1224 0 1 52501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2100
timestamp 1626065694
transform 1 0 1224 0 1 55901
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2099
timestamp 1626065694
transform 1 0 1224 0 1 54133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2098
timestamp 1626065694
transform 1 0 1224 0 1 48965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2097
timestamp 1626065694
transform 1 0 1224 0 1 47469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2096
timestamp 1626065694
transform 1 0 1224 0 1 50869
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2095
timestamp 1626065694
transform 1 0 1224 0 1 45565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2094
timestamp 1626065694
transform 1 0 1224 0 1 44069
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2093
timestamp 1626065694
transform 1 0 1224 0 1 42437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2092
timestamp 1626065694
transform 1 0 21760 0 1 46789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2091
timestamp 1626065694
transform 1 0 21352 0 1 46789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2090
timestamp 1626065694
transform 1 0 20944 0 1 46789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2089
timestamp 1626065694
transform 1 0 27336 0 1 46789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2088
timestamp 1626065694
transform 1 0 27336 0 1 51277
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2087
timestamp 1626065694
transform 1 0 27336 0 1 51005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2086
timestamp 1626065694
transform 1 0 27336 0 1 46925
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2085
timestamp 1626065694
transform 1 0 27336 0 1 47197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2084
timestamp 1626065694
transform 1 0 21760 0 1 51685
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2083
timestamp 1626065694
transform 1 0 22440 0 1 47877
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2082
timestamp 1626065694
transform 1 0 22440 0 1 48149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2081
timestamp 1626065694
transform 1 0 21760 0 1 47061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2080
timestamp 1626065694
transform 1 0 22168 0 1 50733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2079
timestamp 1626065694
transform 1 0 22440 0 1 50597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2078
timestamp 1626065694
transform 1 0 22440 0 1 50325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2077
timestamp 1626065694
transform 1 0 22576 0 1 50733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2076
timestamp 1626065694
transform 1 0 22576 0 1 51005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2075
timestamp 1626065694
transform 1 0 21760 0 1 48557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2074
timestamp 1626065694
transform 1 0 21760 0 1 48285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2073
timestamp 1626065694
transform 1 0 21624 0 1 49101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2072
timestamp 1626065694
transform 1 0 21216 0 1 49373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2071
timestamp 1626065694
transform 1 0 21352 0 1 47061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2070
timestamp 1626065694
transform 1 0 22440 0 1 48285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2069
timestamp 1626065694
transform 1 0 21216 0 1 49101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2068
timestamp 1626065694
transform 1 0 22440 0 1 48557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2067
timestamp 1626065694
transform 1 0 21624 0 1 49373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2066
timestamp 1626065694
transform 1 0 21760 0 1 49781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2065
timestamp 1626065694
transform 1 0 22032 0 1 49373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2064
timestamp 1626065694
transform 1 0 22032 0 1 49101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2063
timestamp 1626065694
transform 1 0 22168 0 1 47877
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2062
timestamp 1626065694
transform 1 0 22168 0 1 48149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2061
timestamp 1626065694
transform 1 0 22168 0 1 51821
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2060
timestamp 1626065694
transform 1 0 22032 0 1 50325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2059
timestamp 1626065694
transform 1 0 22032 0 1 50597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2058
timestamp 1626065694
transform 1 0 22168 0 1 49917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2057
timestamp 1626065694
transform 1 0 22168 0 1 48557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2056
timestamp 1626065694
transform 1 0 22440 0 1 49509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2055
timestamp 1626065694
transform 1 0 22440 0 1 49781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2054
timestamp 1626065694
transform 1 0 22440 0 1 49373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2053
timestamp 1626065694
transform 1 0 22440 0 1 49101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2052
timestamp 1626065694
transform 1 0 22168 0 1 48285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2051
timestamp 1626065694
transform 1 0 22168 0 1 48693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2050
timestamp 1626065694
transform 1 0 22168 0 1 48965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2049
timestamp 1626065694
transform 1 0 22168 0 1 50189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2048
timestamp 1626065694
transform 1 0 20944 0 1 50189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2047
timestamp 1626065694
transform 1 0 21760 0 1 49509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2046
timestamp 1626065694
transform 1 0 21216 0 1 50189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2045
timestamp 1626065694
transform 1 0 20944 0 1 49917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2044
timestamp 1626065694
transform 1 0 22168 0 1 49781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2043
timestamp 1626065694
transform 1 0 22576 0 1 50189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2042
timestamp 1626065694
transform 1 0 22576 0 1 49917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2041
timestamp 1626065694
transform 1 0 20944 0 1 47061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2040
timestamp 1626065694
transform 1 0 21216 0 1 49917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2039
timestamp 1626065694
transform 1 0 20808 0 1 47197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2038
timestamp 1626065694
transform 1 0 20808 0 1 47469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2037
timestamp 1626065694
transform 1 0 20808 0 1 48285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2036
timestamp 1626065694
transform 1 0 20808 0 1 48013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2035
timestamp 1626065694
transform 1 0 22576 0 1 48693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2034
timestamp 1626065694
transform 1 0 22576 0 1 48965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2033
timestamp 1626065694
transform 1 0 22576 0 1 51821
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2032
timestamp 1626065694
transform 1 0 22168 0 1 49509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2031
timestamp 1626065694
transform 1 0 21488 0 1 49917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2030
timestamp 1626065694
transform 1 0 21488 0 1 50189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2029
timestamp 1626065694
transform 1 0 21760 0 1 51413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2028
timestamp 1626065694
transform 1 0 21352 0 1 51005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2027
timestamp 1626065694
transform 1 0 21352 0 1 50733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2026
timestamp 1626065694
transform 1 0 20808 0 1 51413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2025
timestamp 1626065694
transform 1 0 20808 0 1 51141
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2024
timestamp 1626065694
transform 1 0 20944 0 1 49101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2023
timestamp 1626065694
transform 1 0 20944 0 1 49373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2022
timestamp 1626065694
transform 1 0 20808 0 1 48965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2021
timestamp 1626065694
transform 1 0 20808 0 1 48693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2020
timestamp 1626065694
transform 1 0 21352 0 1 48693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2019
timestamp 1626065694
transform 1 0 21352 0 1 48965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2018
timestamp 1626065694
transform 1 0 21488 0 1 47741
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2017
timestamp 1626065694
transform 1 0 21488 0 1 47469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2016
timestamp 1626065694
transform 1 0 21488 0 1 48693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2015
timestamp 1626065694
transform 1 0 21488 0 1 48965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2014
timestamp 1626065694
transform 1 0 20808 0 1 51005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2013
timestamp 1626065694
transform 1 0 20808 0 1 50733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2012
timestamp 1626065694
transform 1 0 20808 0 1 49509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2011
timestamp 1626065694
transform 1 0 20808 0 1 49781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2010
timestamp 1626065694
transform 1 0 20808 0 1 50597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2009
timestamp 1626065694
transform 1 0 20808 0 1 50325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2008
timestamp 1626065694
transform 1 0 21896 0 1 50597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2007
timestamp 1626065694
transform 1 0 21896 0 1 50325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2006
timestamp 1626065694
transform 1 0 21896 0 1 50733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2005
timestamp 1626065694
transform 1 0 21896 0 1 51005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2004
timestamp 1626065694
transform 1 0 22168 0 1 51005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2003
timestamp 1626065694
transform 1 0 20808 0 1 41893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2002
timestamp 1626065694
transform 1 0 22032 0 1 45837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2001
timestamp 1626065694
transform 1 0 20944 0 1 42029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2000
timestamp 1626065694
transform 1 0 20944 0 1 42301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1999
timestamp 1626065694
transform 1 0 20808 0 1 42709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1998
timestamp 1626065694
transform 1 0 20808 0 1 42437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1997
timestamp 1626065694
transform 1 0 20808 0 1 42845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1996
timestamp 1626065694
transform 1 0 20808 0 1 43117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1995
timestamp 1626065694
transform 1 0 20944 0 1 45837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1994
timestamp 1626065694
transform 1 0 20944 0 1 45565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1993
timestamp 1626065694
transform 1 0 20944 0 1 45973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1992
timestamp 1626065694
transform 1 0 20944 0 1 46245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1991
timestamp 1626065694
transform 1 0 22032 0 1 45565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1990
timestamp 1626065694
transform 1 0 22032 0 1 45973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1989
timestamp 1626065694
transform 1 0 22032 0 1 41893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1988
timestamp 1626065694
transform 1 0 22168 0 1 44205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1987
timestamp 1626065694
transform 1 0 22168 0 1 43933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1986
timestamp 1626065694
transform 1 0 21352 0 1 44341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1985
timestamp 1626065694
transform 1 0 22168 0 1 42709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1984
timestamp 1626065694
transform 1 0 22168 0 1 44341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1983
timestamp 1626065694
transform 1 0 22032 0 1 46245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1982
timestamp 1626065694
transform 1 0 21352 0 1 45565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1981
timestamp 1626065694
transform 1 0 21760 0 1 42301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1980
timestamp 1626065694
transform 1 0 22032 0 1 44749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1979
timestamp 1626065694
transform 1 0 20808 0 1 45429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1978
timestamp 1626065694
transform 1 0 20808 0 1 45157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1977
timestamp 1626065694
transform 1 0 21352 0 1 45837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1976
timestamp 1626065694
transform 1 0 22440 0 1 44613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1975
timestamp 1626065694
transform 1 0 22032 0 1 45021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1974
timestamp 1626065694
transform 1 0 22168 0 1 46653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1973
timestamp 1626065694
transform 1 0 21760 0 1 42029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1972
timestamp 1626065694
transform 1 0 22440 0 1 44341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1971
timestamp 1626065694
transform 1 0 22576 0 1 44749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1970
timestamp 1626065694
transform 1 0 22576 0 1 45021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1969
timestamp 1626065694
transform 1 0 22440 0 1 42437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1968
timestamp 1626065694
transform 1 0 22440 0 1 42709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1967
timestamp 1626065694
transform 1 0 23256 0 1 44749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1966
timestamp 1626065694
transform 1 0 23256 0 1 45021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1965
timestamp 1626065694
transform 1 0 21488 0 1 44749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1964
timestamp 1626065694
transform 1 0 22168 0 1 42301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1963
timestamp 1626065694
transform 1 0 21216 0 1 44749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1962
timestamp 1626065694
transform 1 0 21216 0 1 45021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1961
timestamp 1626065694
transform 1 0 21488 0 1 45021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1960
timestamp 1626065694
transform 1 0 22168 0 1 46381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1959
timestamp 1626065694
transform 1 0 20808 0 1 43525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1958
timestamp 1626065694
transform 1 0 20808 0 1 43253
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1957
timestamp 1626065694
transform 1 0 22576 0 1 45973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1956
timestamp 1626065694
transform 1 0 22440 0 1 41893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1955
timestamp 1626065694
transform 1 0 22576 0 1 46245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1954
timestamp 1626065694
transform 1 0 22576 0 1 42029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1953
timestamp 1626065694
transform 1 0 22576 0 1 42301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1952
timestamp 1626065694
transform 1 0 21488 0 1 43117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1951
timestamp 1626065694
transform 1 0 21624 0 1 43389
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1950
timestamp 1626065694
transform 1 0 22576 0 1 44205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1949
timestamp 1626065694
transform 1 0 22576 0 1 43933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1948
timestamp 1626065694
transform 1 0 21216 0 1 42845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1947
timestamp 1626065694
transform 1 0 22440 0 1 45565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1946
timestamp 1626065694
transform 1 0 22440 0 1 45837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1945
timestamp 1626065694
transform 1 0 22440 0 1 45429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1944
timestamp 1626065694
transform 1 0 22440 0 1 45157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1943
timestamp 1626065694
transform 1 0 21216 0 1 46245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1942
timestamp 1626065694
transform 1 0 20808 0 1 46653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1941
timestamp 1626065694
transform 1 0 20808 0 1 46381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1940
timestamp 1626065694
transform 1 0 21216 0 1 45973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1939
timestamp 1626065694
transform 1 0 22032 0 1 43797
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1938
timestamp 1626065694
transform 1 0 22032 0 1 43525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1937
timestamp 1626065694
transform 1 0 21216 0 1 43117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1936
timestamp 1626065694
transform 1 0 22440 0 1 43797
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1935
timestamp 1626065694
transform 1 0 22440 0 1 43525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1934
timestamp 1626065694
transform 1 0 22576 0 1 46381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1933
timestamp 1626065694
transform 1 0 22576 0 1 46653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1932
timestamp 1626065694
transform 1 0 21760 0 1 43525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1931
timestamp 1626065694
transform 1 0 21760 0 1 43797
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1930
timestamp 1626065694
transform 1 0 22168 0 1 42029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1929
timestamp 1626065694
transform 1 0 21624 0 1 41893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1928
timestamp 1626065694
transform 1 0 20944 0 1 44749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1927
timestamp 1626065694
transform 1 0 20944 0 1 45021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1926
timestamp 1626065694
transform 1 0 21760 0 1 45157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1925
timestamp 1626065694
transform 1 0 21760 0 1 45429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1924
timestamp 1626065694
transform 1 0 21216 0 1 41893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1923
timestamp 1626065694
transform 1 0 21352 0 1 44613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1922
timestamp 1626065694
transform 1 0 22168 0 1 44613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1921
timestamp 1626065694
transform 1 0 22032 0 1 45157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1920
timestamp 1626065694
transform 1 0 22168 0 1 42437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1919
timestamp 1626065694
transform 1 0 22032 0 1 45429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1918
timestamp 1626065694
transform 1 0 27608 0 1 42981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1917
timestamp 1626065694
transform 1 0 27472 0 1 43389
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1916
timestamp 1626065694
transform 1 0 27336 0 1 46517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1915
timestamp 1626065694
transform 1 0 25840 0 1 45157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1914
timestamp 1626065694
transform 1 0 25840 0 1 45429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1913
timestamp 1626065694
transform 1 0 27472 0 1 43661
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1912
timestamp 1626065694
transform 1 0 27608 0 1 43253
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1911
timestamp 1626065694
transform 1 0 17816 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1910
timestamp 1626065694
transform 1 0 18632 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1909
timestamp 1626065694
transform 1 0 20808 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1908
timestamp 1626065694
transform 1 0 18360 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1907
timestamp 1626065694
transform 1 0 19176 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1906
timestamp 1626065694
transform 1 0 21352 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1905
timestamp 1626065694
transform 1 0 22032 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1904
timestamp 1626065694
transform 1 0 21760 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1903
timestamp 1626065694
transform 1 0 22440 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1902
timestamp 1626065694
transform 1 0 22168 0 1 31285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1901
timestamp 1626065694
transform 1 0 22440 0 1 31285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1900
timestamp 1626065694
transform 1 0 22032 0 1 36453
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1899
timestamp 1626065694
transform 1 0 21760 0 1 36453
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1898
timestamp 1626065694
transform 1 0 22440 0 1 36453
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1897
timestamp 1626065694
transform 1 0 27472 0 1 40533
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1896
timestamp 1626065694
transform 1 0 27472 0 1 40261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1895
timestamp 1626065694
transform 1 0 27472 0 1 39037
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1894
timestamp 1626065694
transform 1 0 27472 0 1 39309
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1893
timestamp 1626065694
transform 1 0 27336 0 1 37813
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1892
timestamp 1626065694
transform 1 0 27336 0 1 38085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1891
timestamp 1626065694
transform 1 0 20808 0 1 39309
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1890
timestamp 1626065694
transform 1 0 20808 0 1 36861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1889
timestamp 1626065694
transform 1 0 20808 0 1 37133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1888
timestamp 1626065694
transform 1 0 20808 0 1 39173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1887
timestamp 1626065694
transform 1 0 20808 0 1 38901
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1886
timestamp 1626065694
transform 1 0 20808 0 1 37541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1885
timestamp 1626065694
transform 1 0 20808 0 1 37269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1884
timestamp 1626065694
transform 1 0 20944 0 1 37677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1883
timestamp 1626065694
transform 1 0 20944 0 1 37949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1882
timestamp 1626065694
transform 1 0 22032 0 1 40669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1881
timestamp 1626065694
transform 1 0 22032 0 1 40397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1880
timestamp 1626065694
transform 1 0 22032 0 1 40805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1879
timestamp 1626065694
transform 1 0 22032 0 1 41077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1878
timestamp 1626065694
transform 1 0 22032 0 1 37541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1877
timestamp 1626065694
transform 1 0 22032 0 1 37269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1876
timestamp 1626065694
transform 1 0 22168 0 1 37677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1875
timestamp 1626065694
transform 1 0 22168 0 1 37949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1874
timestamp 1626065694
transform 1 0 22032 0 1 38357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1873
timestamp 1626065694
transform 1 0 22032 0 1 38085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1872
timestamp 1626065694
transform 1 0 20808 0 1 41213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1871
timestamp 1626065694
transform 1 0 22032 0 1 36725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1870
timestamp 1626065694
transform 1 0 22032 0 1 39581
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1869
timestamp 1626065694
transform 1 0 22032 0 1 39853
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1868
timestamp 1626065694
transform 1 0 22168 0 1 40261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1867
timestamp 1626065694
transform 1 0 22168 0 1 39989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1866
timestamp 1626065694
transform 1 0 22168 0 1 36861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1865
timestamp 1626065694
transform 1 0 22168 0 1 37133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1864
timestamp 1626065694
transform 1 0 22032 0 1 41485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1863
timestamp 1626065694
transform 1 0 22032 0 1 41213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1862
timestamp 1626065694
transform 1 0 21352 0 1 36861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1861
timestamp 1626065694
transform 1 0 21352 0 1 37133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1860
timestamp 1626065694
transform 1 0 21488 0 1 36861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1859
timestamp 1626065694
transform 1 0 21488 0 1 37133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1858
timestamp 1626065694
transform 1 0 21488 0 1 38901
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1857
timestamp 1626065694
transform 1 0 21488 0 1 39173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1856
timestamp 1626065694
transform 1 0 21216 0 1 37541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1855
timestamp 1626065694
transform 1 0 21216 0 1 37269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1854
timestamp 1626065694
transform 1 0 20808 0 1 41485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1853
timestamp 1626065694
transform 1 0 20808 0 1 41077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1852
timestamp 1626065694
transform 1 0 20808 0 1 40805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1851
timestamp 1626065694
transform 1 0 20808 0 1 38493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1850
timestamp 1626065694
transform 1 0 20808 0 1 38765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1849
timestamp 1626065694
transform 1 0 20808 0 1 38357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1848
timestamp 1626065694
transform 1 0 21352 0 1 38085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1847
timestamp 1626065694
transform 1 0 21352 0 1 38357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1846
timestamp 1626065694
transform 1 0 21352 0 1 41213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1845
timestamp 1626065694
transform 1 0 21352 0 1 41485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1844
timestamp 1626065694
transform 1 0 21216 0 1 40669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1843
timestamp 1626065694
transform 1 0 21216 0 1 40397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1842
timestamp 1626065694
transform 1 0 21760 0 1 41077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1841
timestamp 1626065694
transform 1 0 21760 0 1 40805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1840
timestamp 1626065694
transform 1 0 21760 0 1 39853
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1839
timestamp 1626065694
transform 1 0 21760 0 1 39581
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1838
timestamp 1626065694
transform 1 0 21624 0 1 40397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1837
timestamp 1626065694
transform 1 0 21624 0 1 40669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1836
timestamp 1626065694
transform 1 0 21624 0 1 37269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1835
timestamp 1626065694
transform 1 0 21624 0 1 37541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1834
timestamp 1626065694
transform 1 0 21760 0 1 36725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1833
timestamp 1626065694
transform 1 0 20808 0 1 38085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1832
timestamp 1626065694
transform 1 0 21760 0 1 37949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1831
timestamp 1626065694
transform 1 0 21760 0 1 37677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1830
timestamp 1626065694
transform 1 0 22576 0 1 40397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1829
timestamp 1626065694
transform 1 0 22576 0 1 40669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1828
timestamp 1626065694
transform 1 0 22440 0 1 40261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1827
timestamp 1626065694
transform 1 0 22440 0 1 39989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1826
timestamp 1626065694
transform 1 0 20808 0 1 39581
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1825
timestamp 1626065694
transform 1 0 22440 0 1 36725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1824
timestamp 1626065694
transform 1 0 22440 0 1 37949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1823
timestamp 1626065694
transform 1 0 22440 0 1 37677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1822
timestamp 1626065694
transform 1 0 22440 0 1 38085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1821
timestamp 1626065694
transform 1 0 22440 0 1 38357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1820
timestamp 1626065694
transform 1 0 22576 0 1 41485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1819
timestamp 1626065694
transform 1 0 22576 0 1 41213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1818
timestamp 1626065694
transform 1 0 22576 0 1 37269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1817
timestamp 1626065694
transform 1 0 22576 0 1 37541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1816
timestamp 1626065694
transform 1 0 22576 0 1 37133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1815
timestamp 1626065694
transform 1 0 22576 0 1 36861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1814
timestamp 1626065694
transform 1 0 22440 0 1 41077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1813
timestamp 1626065694
transform 1 0 22440 0 1 40805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1812
timestamp 1626065694
transform 1 0 22576 0 1 39581
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1811
timestamp 1626065694
transform 1 0 22576 0 1 39853
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1810
timestamp 1626065694
transform 1 0 22032 0 1 36045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1809
timestamp 1626065694
transform 1 0 20944 0 1 36045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1808
timestamp 1626065694
transform 1 0 20944 0 1 32373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1807
timestamp 1626065694
transform 1 0 20808 0 1 34005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1806
timestamp 1626065694
transform 1 0 20808 0 1 33733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1805
timestamp 1626065694
transform 1 0 22032 0 1 31965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1804
timestamp 1626065694
transform 1 0 21352 0 1 33733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1803
timestamp 1626065694
transform 1 0 21352 0 1 34005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1802
timestamp 1626065694
transform 1 0 21352 0 1 33597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1801
timestamp 1626065694
transform 1 0 21352 0 1 33325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1800
timestamp 1626065694
transform 1 0 21216 0 1 34141
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1799
timestamp 1626065694
transform 1 0 21216 0 1 34413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1798
timestamp 1626065694
transform 1 0 21488 0 1 35909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1797
timestamp 1626065694
transform 1 0 21488 0 1 35637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1796
timestamp 1626065694
transform 1 0 22032 0 1 31693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1795
timestamp 1626065694
transform 1 0 22032 0 1 32101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1794
timestamp 1626065694
transform 1 0 21352 0 1 35501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1793
timestamp 1626065694
transform 1 0 21624 0 1 35501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1792
timestamp 1626065694
transform 1 0 21216 0 1 31965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1791
timestamp 1626065694
transform 1 0 21216 0 1 31693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1790
timestamp 1626065694
transform 1 0 22032 0 1 32373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1789
timestamp 1626065694
transform 1 0 22032 0 1 34141
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1788
timestamp 1626065694
transform 1 0 21488 0 1 36317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1787
timestamp 1626065694
transform 1 0 21488 0 1 36045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1786
timestamp 1626065694
transform 1 0 22032 0 1 34413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1785
timestamp 1626065694
transform 1 0 22032 0 1 34005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1784
timestamp 1626065694
transform 1 0 22032 0 1 33733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1783
timestamp 1626065694
transform 1 0 20944 0 1 32101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1782
timestamp 1626065694
transform 1 0 21760 0 1 32373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1781
timestamp 1626065694
transform 1 0 21760 0 1 32101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1780
timestamp 1626065694
transform 1 0 21624 0 1 36045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1779
timestamp 1626065694
transform 1 0 21624 0 1 36317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1778
timestamp 1626065694
transform 1 0 21760 0 1 33597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1777
timestamp 1626065694
transform 1 0 21760 0 1 33325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1776
timestamp 1626065694
transform 1 0 21624 0 1 31965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1775
timestamp 1626065694
transform 1 0 21624 0 1 31693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1774
timestamp 1626065694
transform 1 0 20944 0 1 32509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1773
timestamp 1626065694
transform 1 0 20808 0 1 34141
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1772
timestamp 1626065694
transform 1 0 20944 0 1 32781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1771
timestamp 1626065694
transform 1 0 20808 0 1 35365
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1770
timestamp 1626065694
transform 1 0 22168 0 1 31557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1769
timestamp 1626065694
transform 1 0 20808 0 1 34413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1768
timestamp 1626065694
transform 1 0 21896 0 1 35229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1767
timestamp 1626065694
transform 1 0 21896 0 1 34821
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1766
timestamp 1626065694
transform 1 0 20808 0 1 35637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1765
timestamp 1626065694
transform 1 0 20808 0 1 33325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1764
timestamp 1626065694
transform 1 0 21624 0 1 32917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1763
timestamp 1626065694
transform 1 0 21624 0 1 33189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1762
timestamp 1626065694
transform 1 0 22440 0 1 33733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1761
timestamp 1626065694
transform 1 0 22440 0 1 34005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1760
timestamp 1626065694
transform 1 0 22440 0 1 33597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1759
timestamp 1626065694
transform 1 0 22440 0 1 33325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1758
timestamp 1626065694
transform 1 0 22168 0 1 33597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1757
timestamp 1626065694
transform 1 0 22168 0 1 33325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1756
timestamp 1626065694
transform 1 0 22032 0 1 32781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1755
timestamp 1626065694
transform 1 0 22032 0 1 32509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1754
timestamp 1626065694
transform 1 0 22440 0 1 34141
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1753
timestamp 1626065694
transform 1 0 22440 0 1 34413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1752
timestamp 1626065694
transform 1 0 22032 0 1 32917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1751
timestamp 1626065694
transform 1 0 22032 0 1 33189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1750
timestamp 1626065694
transform 1 0 22440 0 1 36317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1749
timestamp 1626065694
transform 1 0 22440 0 1 36045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1748
timestamp 1626065694
transform 1 0 20944 0 1 31421
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1747
timestamp 1626065694
transform 1 0 20808 0 1 33597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1746
timestamp 1626065694
transform 1 0 21216 0 1 32781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1745
timestamp 1626065694
transform 1 0 21216 0 1 32509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1744
timestamp 1626065694
transform 1 0 22440 0 1 33189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1743
timestamp 1626065694
transform 1 0 22440 0 1 32917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1742
timestamp 1626065694
transform 1 0 22440 0 1 31557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1741
timestamp 1626065694
transform 1 0 20944 0 1 31693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1740
timestamp 1626065694
transform 1 0 22576 0 1 31693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1739
timestamp 1626065694
transform 1 0 22576 0 1 31965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1738
timestamp 1626065694
transform 1 0 20944 0 1 34957
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1737
timestamp 1626065694
transform 1 0 20944 0 1 35229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1736
timestamp 1626065694
transform 1 0 20808 0 1 34821
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1735
timestamp 1626065694
transform 1 0 20808 0 1 34549
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1734
timestamp 1626065694
transform 1 0 20808 0 1 33189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1733
timestamp 1626065694
transform 1 0 20808 0 1 32917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1732
timestamp 1626065694
transform 1 0 20944 0 1 36317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1731
timestamp 1626065694
transform 1 0 22168 0 1 35637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1730
timestamp 1626065694
transform 1 0 22576 0 1 32781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1729
timestamp 1626065694
transform 1 0 22576 0 1 32509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1728
timestamp 1626065694
transform 1 0 22440 0 1 35909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1727
timestamp 1626065694
transform 1 0 22440 0 1 35637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1726
timestamp 1626065694
transform 1 0 22440 0 1 32373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1725
timestamp 1626065694
transform 1 0 22440 0 1 32101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1724
timestamp 1626065694
transform 1 0 22168 0 1 35909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1723
timestamp 1626065694
transform 1 0 22032 0 1 36317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1722
timestamp 1626065694
transform 1 0 27472 0 1 34957
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1721
timestamp 1626065694
transform 1 0 27472 0 1 35229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1720
timestamp 1626065694
transform 1 0 14144 0 1 37541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1719
timestamp 1626065694
transform 1 0 1224 0 1 39037
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1718
timestamp 1626065694
transform 1 0 1224 0 1 40805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1717
timestamp 1626065694
transform 1 0 1224 0 1 37269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1716
timestamp 1626065694
transform 1 0 1224 0 1 34005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1715
timestamp 1626065694
transform 1 0 1224 0 1 32373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1714
timestamp 1626065694
transform 1 0 1224 0 1 35637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1713
timestamp 1626065694
transform 1 0 14008 0 1 34685
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1712
timestamp 1626065694
transform 1 0 14144 0 1 31829
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1711
timestamp 1626065694
transform 1 0 14008 0 1 32101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1710
timestamp 1626065694
transform 1 0 14144 0 1 34821
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1709
timestamp 1626065694
transform 1 0 14144 0 1 33325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1708
timestamp 1626065694
transform 1 0 14280 0 1 33461
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1707
timestamp 1626065694
transform 1 0 14280 0 1 36181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1706
timestamp 1626065694
transform 1 0 14144 0 1 29245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1705
timestamp 1626065694
transform 1 0 14008 0 1 27749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1704
timestamp 1626065694
transform 1 0 14008 0 1 30469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1703
timestamp 1626065694
transform 1 0 15912 0 1 27613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1702
timestamp 1626065694
transform 1 0 14008 0 1 30605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1701
timestamp 1626065694
transform 1 0 1224 0 1 30469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1700
timestamp 1626065694
transform 1 0 1224 0 1 28973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1699
timestamp 1626065694
transform 1 0 1224 0 1 27205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1698
timestamp 1626065694
transform 1 0 3128 0 1 22173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1697
timestamp 1626065694
transform 1 0 3128 0 1 21765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1696
timestamp 1626065694
transform 1 0 1224 0 1 22309
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1695
timestamp 1626065694
transform 1 0 1224 0 1 25573
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1694
timestamp 1626065694
transform 1 0 3808 0 1 23125
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1693
timestamp 1626065694
transform 1 0 3808 0 1 23261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1692
timestamp 1626065694
transform 1 0 3808 0 1 25845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1691
timestamp 1626065694
transform 1 0 544 0 1 23125
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1690
timestamp 1626065694
transform 1 0 2312 0 1 23941
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1689
timestamp 1626065694
transform 1 0 2312 0 1 24485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1688
timestamp 1626065694
transform 1 0 1224 0 1 23941
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1687
timestamp 1626065694
transform 1 0 2531 0 1 25300
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1686
timestamp 1626065694
transform 1 0 15912 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1685
timestamp 1626065694
transform 1 0 22168 0 1 26117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1684
timestamp 1626065694
transform 1 0 20808 0 1 26117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1683
timestamp 1626065694
transform 1 0 22576 0 1 26117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1682
timestamp 1626065694
transform 1 0 27336 0 1 26661
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1681
timestamp 1626065694
transform 1 0 27336 0 1 26389
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1680
timestamp 1626065694
transform 1 0 27336 0 1 31013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1679
timestamp 1626065694
transform 1 0 27336 0 1 30741
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1678
timestamp 1626065694
transform 1 0 27472 0 1 26253
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1677
timestamp 1626065694
transform 1 0 27472 0 1 30605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1676
timestamp 1626065694
transform 1 0 27472 0 1 30333
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1675
timestamp 1626065694
transform 1 0 22032 0 1 27749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1674
timestamp 1626065694
transform 1 0 22032 0 1 28021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1673
timestamp 1626065694
transform 1 0 22032 0 1 27613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1672
timestamp 1626065694
transform 1 0 22032 0 1 27341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1671
timestamp 1626065694
transform 1 0 21216 0 1 28837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1670
timestamp 1626065694
transform 1 0 21216 0 1 28565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1669
timestamp 1626065694
transform 1 0 22168 0 1 28157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1668
timestamp 1626065694
transform 1 0 21352 0 1 26933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1667
timestamp 1626065694
transform 1 0 21352 0 1 27205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1666
timestamp 1626065694
transform 1 0 21488 0 1 26933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1665
timestamp 1626065694
transform 1 0 21488 0 1 27205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1664
timestamp 1626065694
transform 1 0 22168 0 1 28429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1663
timestamp 1626065694
transform 1 0 19040 0 1 26661
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1662
timestamp 1626065694
transform 1 0 19040 0 1 27205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1661
timestamp 1626065694
transform 1 0 18632 0 1 26661
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1660
timestamp 1626065694
transform 1 0 18632 0 1 27205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1659
timestamp 1626065694
transform 1 0 20808 0 1 30469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1658
timestamp 1626065694
transform 1 0 20672 0 1 27205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1657
timestamp 1626065694
transform 1 0 20672 0 1 26797
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1656
timestamp 1626065694
transform 1 0 20808 0 1 30197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1655
timestamp 1626065694
transform 1 0 18632 0 1 26389
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1654
timestamp 1626065694
transform 1 0 22032 0 1 29653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1653
timestamp 1626065694
transform 1 0 22032 0 1 29381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1652
timestamp 1626065694
transform 1 0 21488 0 1 29381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1651
timestamp 1626065694
transform 1 0 21488 0 1 29653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1650
timestamp 1626065694
transform 1 0 20808 0 1 30877
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1649
timestamp 1626065694
transform 1 0 20808 0 1 30605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1648
timestamp 1626065694
transform 1 0 18904 0 1 27341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1647
timestamp 1626065694
transform 1 0 18904 0 1 28021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1646
timestamp 1626065694
transform 1 0 21352 0 1 28157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1645
timestamp 1626065694
transform 1 0 21760 0 1 29653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1644
timestamp 1626065694
transform 1 0 21760 0 1 29381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1643
timestamp 1626065694
transform 1 0 20808 0 1 26661
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1642
timestamp 1626065694
transform 1 0 21352 0 1 30197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1641
timestamp 1626065694
transform 1 0 21352 0 1 30469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1640
timestamp 1626065694
transform 1 0 20808 0 1 26933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1639
timestamp 1626065694
transform 1 0 20808 0 1 26525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1638
timestamp 1626065694
transform 1 0 20808 0 1 26253
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1637
timestamp 1626065694
transform 1 0 21896 0 1 26253
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1636
timestamp 1626065694
transform 1 0 21896 0 1 26525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1635
timestamp 1626065694
transform 1 0 17816 0 1 29109
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1634
timestamp 1626065694
transform 1 0 21760 0 1 27749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1633
timestamp 1626065694
transform 1 0 21760 0 1 28021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1632
timestamp 1626065694
transform 1 0 17816 0 1 27477
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1631
timestamp 1626065694
transform 1 0 20944 0 1 30061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1630
timestamp 1626065694
transform 1 0 20944 0 1 29789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1629
timestamp 1626065694
transform 1 0 21760 0 1 29245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1628
timestamp 1626065694
transform 1 0 21760 0 1 28973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1627
timestamp 1626065694
transform 1 0 21760 0 1 31149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1626
timestamp 1626065694
transform 1 0 21760 0 1 30877
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1625
timestamp 1626065694
transform 1 0 22032 0 1 28837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1624
timestamp 1626065694
transform 1 0 21624 0 1 28565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1623
timestamp 1626065694
transform 1 0 21624 0 1 28837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1622
timestamp 1626065694
transform 1 0 22032 0 1 28565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1621
timestamp 1626065694
transform 1 0 21488 0 1 28157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1620
timestamp 1626065694
transform 1 0 21488 0 1 28429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1619
timestamp 1626065694
transform 1 0 21216 0 1 26525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1618
timestamp 1626065694
transform 1 0 21216 0 1 26253
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1617
timestamp 1626065694
transform 1 0 22168 0 1 28973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1616
timestamp 1626065694
transform 1 0 22168 0 1 29245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1615
timestamp 1626065694
transform 1 0 17408 0 1 27205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1614
timestamp 1626065694
transform 1 0 20808 0 1 29381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1613
timestamp 1626065694
transform 1 0 22440 0 1 28157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1612
timestamp 1626065694
transform 1 0 22440 0 1 28429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1611
timestamp 1626065694
transform 1 0 22440 0 1 28021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1610
timestamp 1626065694
transform 1 0 22440 0 1 27749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1609
timestamp 1626065694
transform 1 0 20808 0 1 29653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1608
timestamp 1626065694
transform 1 0 20808 0 1 29245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1607
timestamp 1626065694
transform 1 0 20808 0 1 28973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1606
timestamp 1626065694
transform 1 0 17408 0 1 26661
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1605
timestamp 1626065694
transform 1 0 18224 0 1 26389
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1604
timestamp 1626065694
transform 1 0 17544 0 1 26525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1603
timestamp 1626065694
transform 1 0 20944 0 1 28429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1602
timestamp 1626065694
transform 1 0 20944 0 1 28157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1601
timestamp 1626065694
transform 1 0 22576 0 1 28565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1600
timestamp 1626065694
transform 1 0 22576 0 1 28837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1599
timestamp 1626065694
transform 1 0 20944 0 1 28565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1598
timestamp 1626065694
transform 1 0 20944 0 1 28837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1597
timestamp 1626065694
transform 1 0 22576 0 1 27341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1596
timestamp 1626065694
transform 1 0 22576 0 1 27613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1595
timestamp 1626065694
transform 1 0 22576 0 1 30061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1594
timestamp 1626065694
transform 1 0 22576 0 1 29789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1593
timestamp 1626065694
transform 1 0 22576 0 1 28973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1592
timestamp 1626065694
transform 1 0 22576 0 1 29245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1591
timestamp 1626065694
transform 1 0 21352 0 1 28429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1590
timestamp 1626065694
transform 1 0 18360 0 1 26661
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1589
timestamp 1626065694
transform 1 0 17680 0 1 26525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1588
timestamp 1626065694
transform 1 0 18360 0 1 27205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1587
timestamp 1626065694
transform 1 0 17680 0 1 26253
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1586
timestamp 1626065694
transform 1 0 22168 0 1 30061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1585
timestamp 1626065694
transform 1 0 22440 0 1 29381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1584
timestamp 1626065694
transform 1 0 22440 0 1 29653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1583
timestamp 1626065694
transform 1 0 22168 0 1 29789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1582
timestamp 1626065694
transform 1 0 21488 0 1 21493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1581
timestamp 1626065694
transform 1 0 21488 0 1 21765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1580
timestamp 1626065694
transform 1 0 21488 0 1 22989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1579
timestamp 1626065694
transform 1 0 21488 0 1 22717
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1578
timestamp 1626065694
transform 1 0 21488 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1577
timestamp 1626065694
transform 1 0 21488 0 1 23805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1576
timestamp 1626065694
transform 1 0 21488 0 1 24077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1575
timestamp 1626065694
transform 1 0 21488 0 1 25301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1574
timestamp 1626065694
transform 1 0 22168 0 1 25845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1573
timestamp 1626065694
transform 1 0 22168 0 1 25437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1572
timestamp 1626065694
transform 1 0 21624 0 1 24213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1571
timestamp 1626065694
transform 1 0 21624 0 1 24485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1570
timestamp 1626065694
transform 1 0 21760 0 1 25301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1569
timestamp 1626065694
transform 1 0 21760 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1568
timestamp 1626065694
transform 1 0 21896 0 1 24621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1567
timestamp 1626065694
transform 1 0 21896 0 1 24893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1566
timestamp 1626065694
transform 1 0 22032 0 1 24213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1565
timestamp 1626065694
transform 1 0 22576 0 1 25437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1564
timestamp 1626065694
transform 1 0 22576 0 1 25709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1563
timestamp 1626065694
transform 1 0 22440 0 1 25301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1562
timestamp 1626065694
transform 1 0 22440 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1561
timestamp 1626065694
transform 1 0 22032 0 1 24485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1560
timestamp 1626065694
transform 1 0 22576 0 1 24621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1559
timestamp 1626065694
transform 1 0 22576 0 1 24893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1558
timestamp 1626065694
transform 1 0 22440 0 1 24485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1557
timestamp 1626065694
transform 1 0 22440 0 1 24213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1556
timestamp 1626065694
transform 1 0 22168 0 1 24893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1555
timestamp 1626065694
transform 1 0 22168 0 1 23669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1554
timestamp 1626065694
transform 1 0 22168 0 1 24621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1553
timestamp 1626065694
transform 1 0 22168 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1552
timestamp 1626065694
transform 1 0 22440 0 1 23669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1551
timestamp 1626065694
transform 1 0 22576 0 1 25845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1550
timestamp 1626065694
transform 1 0 22168 0 1 25301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1549
timestamp 1626065694
transform 1 0 22032 0 1 24077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1548
timestamp 1626065694
transform 1 0 22032 0 1 23805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1547
timestamp 1626065694
transform 1 0 22440 0 1 23805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1546
timestamp 1626065694
transform 1 0 22440 0 1 24077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1545
timestamp 1626065694
transform 1 0 22168 0 1 25709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1544
timestamp 1626065694
transform 1 0 17680 0 1 24893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1543
timestamp 1626065694
transform 1 0 19176 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1542
timestamp 1626065694
transform 1 0 19176 0 1 25709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1541
timestamp 1626065694
transform 1 0 18224 0 1 25709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1540
timestamp 1626065694
transform 1 0 18224 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1539
timestamp 1626065694
transform 1 0 18224 0 1 24893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1538
timestamp 1626065694
transform 1 0 20808 0 1 25437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1537
timestamp 1626065694
transform 1 0 20944 0 1 24213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1536
timestamp 1626065694
transform 1 0 21352 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1535
timestamp 1626065694
transform 1 0 18632 0 1 25845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1534
timestamp 1626065694
transform 1 0 17408 0 1 25709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1533
timestamp 1626065694
transform 1 0 20944 0 1 24485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1532
timestamp 1626065694
transform 1 0 17544 0 1 25845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1531
timestamp 1626065694
transform 1 0 20808 0 1 25709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1530
timestamp 1626065694
transform 1 0 21216 0 1 24077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1529
timestamp 1626065694
transform 1 0 21216 0 1 23805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1528
timestamp 1626065694
transform 1 0 21352 0 1 25301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1527
timestamp 1626065694
transform 1 0 20808 0 1 25845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1526
timestamp 1626065694
transform 1 0 17408 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1525
timestamp 1626065694
transform 1 0 18768 0 1 25709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1524
timestamp 1626065694
transform 1 0 18768 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1523
timestamp 1626065694
transform 1 0 20808 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1522
timestamp 1626065694
transform 1 0 20808 0 1 25301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1521
timestamp 1626065694
transform 1 0 18224 0 1 25845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1520
timestamp 1626065694
transform 1 0 20808 0 1 24893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1519
timestamp 1626065694
transform 1 0 20808 0 1 24621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1518
timestamp 1626065694
transform 1 0 20944 0 1 21085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1517
timestamp 1626065694
transform 1 0 20944 0 1 21493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1516
timestamp 1626065694
transform 1 0 20944 0 1 21765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1515
timestamp 1626065694
transform 1 0 19040 0 1 22717
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1514
timestamp 1626065694
transform 1 0 20944 0 1 21901
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1513
timestamp 1626065694
transform 1 0 20944 0 1 22173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1512
timestamp 1626065694
transform 1 0 18224 0 1 22717
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1511
timestamp 1626065694
transform 1 0 20808 0 1 22581
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1510
timestamp 1626065694
transform 1 0 18632 0 1 21085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1509
timestamp 1626065694
transform 1 0 18632 0 1 22445
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1508
timestamp 1626065694
transform 1 0 18224 0 1 23261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1507
timestamp 1626065694
transform 1 0 20808 0 1 22309
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1506
timestamp 1626065694
transform 1 0 20944 0 1 22989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1505
timestamp 1626065694
transform 1 0 17680 0 1 23397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1504
timestamp 1626065694
transform 1 0 20944 0 1 22717
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1503
timestamp 1626065694
transform 1 0 18632 0 1 22717
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1502
timestamp 1626065694
transform 1 0 21352 0 1 21765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1501
timestamp 1626065694
transform 1 0 18632 0 1 23261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1500
timestamp 1626065694
transform 1 0 18360 0 1 22445
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1499
timestamp 1626065694
transform 1 0 21352 0 1 23261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1498
timestamp 1626065694
transform 1 0 18224 0 1 23397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1497
timestamp 1626065694
transform 1 0 18360 0 1 21085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1496
timestamp 1626065694
transform 1 0 21352 0 1 22989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1495
timestamp 1626065694
transform 1 0 19040 0 1 23261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1494
timestamp 1626065694
transform 1 0 21352 0 1 21493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1493
timestamp 1626065694
transform 1 0 20944 0 1 21357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1492
timestamp 1626065694
transform 1 0 21624 0 1 22309
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1491
timestamp 1626065694
transform 1 0 22032 0 1 22989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1490
timestamp 1626065694
transform 1 0 22032 0 1 23261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1489
timestamp 1626065694
transform 1 0 22576 0 1 22989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1488
timestamp 1626065694
transform 1 0 22576 0 1 23261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1487
timestamp 1626065694
transform 1 0 22168 0 1 23397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1486
timestamp 1626065694
transform 1 0 21624 0 1 22581
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1485
timestamp 1626065694
transform 1 0 21624 0 1 23261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1484
timestamp 1626065694
transform 1 0 22440 0 1 23397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1483
timestamp 1626065694
transform 1 0 21624 0 1 22989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1482
timestamp 1626065694
transform 1 0 22168 0 1 21765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1481
timestamp 1626065694
transform 1 0 22440 0 1 21765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1480
timestamp 1626065694
transform 1 0 22440 0 1 21085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1479
timestamp 1626065694
transform 1 0 22440 0 1 21357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1478
timestamp 1626065694
transform 1 0 22440 0 1 21493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1477
timestamp 1626065694
transform 1 0 22168 0 1 21357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1476
timestamp 1626065694
transform 1 0 22168 0 1 21085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1475
timestamp 1626065694
transform 1 0 22168 0 1 21493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1474
timestamp 1626065694
transform 1 0 21624 0 1 21357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1473
timestamp 1626065694
transform 1 0 21624 0 1 21085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1472
timestamp 1626065694
transform 1 0 21760 0 1 21493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1471
timestamp 1626065694
transform 1 0 21760 0 1 21765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1470
timestamp 1626065694
transform 1 0 27472 0 1 22717
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1469
timestamp 1626065694
transform 1 0 27472 0 1 25981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1468
timestamp 1626065694
transform 1 0 27336 0 1 23125
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1467
timestamp 1626065694
transform 1 0 27336 0 1 22309
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1466
timestamp 1626065694
transform 1 0 27336 0 1 22853
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1465
timestamp 1626065694
transform 1 0 27336 0 1 22037
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1464
timestamp 1626065694
transform 1 0 27472 0 1 23669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1463
timestamp 1626065694
transform 1 0 27472 0 1 23261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1462
timestamp 1626065694
transform 1 0 27608 0 1 23669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1461
timestamp 1626065694
transform 1 0 27608 0 1 23941
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1460
timestamp 1626065694
transform 1 0 27472 0 1 22445
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1459
timestamp 1626065694
transform 1 0 28560 0 1 10613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1458
timestamp 1626065694
transform 1 0 21216 0 1 15781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1457
timestamp 1626065694
transform 1 0 22440 0 1 15781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1456
timestamp 1626065694
transform 1 0 28968 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1455
timestamp 1626065694
transform 1 0 31688 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1454
timestamp 1626065694
transform 1 0 34000 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1453
timestamp 1626065694
transform 1 0 28968 0 1 19725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1452
timestamp 1626065694
transform 1 0 28968 0 1 17141
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1451
timestamp 1626065694
transform 1 0 28288 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1450
timestamp 1626065694
transform 1 0 28560 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1449
timestamp 1626065694
transform 1 0 28560 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1448
timestamp 1626065694
transform 1 0 29512 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1447
timestamp 1626065694
transform 1 0 29512 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1446
timestamp 1626065694
transform 1 0 30736 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1445
timestamp 1626065694
transform 1 0 30736 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1444
timestamp 1626065694
transform 1 0 32504 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1443
timestamp 1626065694
transform 1 0 32504 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1442
timestamp 1626065694
transform 1 0 33184 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1441
timestamp 1626065694
transform 1 0 33184 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1440
timestamp 1626065694
transform 1 0 33728 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1439
timestamp 1626065694
transform 1 0 33728 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1438
timestamp 1626065694
transform 1 0 26928 0 1 19589
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1437
timestamp 1626065694
transform 1 0 26928 0 1 19317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1436
timestamp 1626065694
transform 1 0 28288 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1435
timestamp 1626065694
transform 1 0 20808 0 1 20677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1434
timestamp 1626065694
transform 1 0 22032 0 1 20677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1433
timestamp 1626065694
transform 1 0 21080 0 1 20133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1432
timestamp 1626065694
transform 1 0 21760 0 1 20677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1431
timestamp 1626065694
transform 1 0 21760 0 1 20541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1430
timestamp 1626065694
transform 1 0 21760 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1429
timestamp 1626065694
transform 1 0 21216 0 1 17277
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1428
timestamp 1626065694
transform 1 0 21352 0 1 17141
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1427
timestamp 1626065694
transform 1 0 17816 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1426
timestamp 1626065694
transform 1 0 22440 0 1 20677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1425
timestamp 1626065694
transform 1 0 18360 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1424
timestamp 1626065694
transform 1 0 18632 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1423
timestamp 1626065694
transform 1 0 22168 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1422
timestamp 1626065694
transform 1 0 22168 0 1 20541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1421
timestamp 1626065694
transform 1 0 19176 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1420
timestamp 1626065694
transform 1 0 22440 0 1 19589
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1419
timestamp 1626065694
transform 1 0 21352 0 1 20541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1418
timestamp 1626065694
transform 1 0 20944 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1417
timestamp 1626065694
transform 1 0 22440 0 1 20541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1416
timestamp 1626065694
transform 1 0 22440 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1415
timestamp 1626065694
transform 1 0 22440 0 1 20133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1414
timestamp 1626065694
transform 1 0 22440 0 1 19725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1413
timestamp 1626065694
transform 1 0 21352 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1412
timestamp 1626065694
transform 1 0 21352 0 1 20677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1411
timestamp 1626065694
transform 1 0 20944 0 1 20541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1410
timestamp 1626065694
transform 1 0 21352 0 1 14557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1409
timestamp 1626065694
transform 1 0 21216 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1408
timestamp 1626065694
transform 1 0 20264 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1407
timestamp 1626065694
transform 1 0 20264 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1406
timestamp 1626065694
transform 1 0 28968 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1405
timestamp 1626065694
transform 1 0 28288 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1404
timestamp 1626065694
transform 1 0 30736 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1403
timestamp 1626065694
transform 1 0 33592 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1402
timestamp 1626065694
transform 1 0 28152 0 1 11293
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1401
timestamp 1626065694
transform 1 0 31416 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1400
timestamp 1626065694
transform 1 0 28696 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1399
timestamp 1626065694
transform 1 0 28696 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1398
timestamp 1626065694
transform 1 0 28968 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1397
timestamp 1626065694
transform 1 0 28968 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1396
timestamp 1626065694
transform 1 0 31416 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1395
timestamp 1626065694
transform 1 0 31416 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1394
timestamp 1626065694
transform 1 0 28832 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1393
timestamp 1626065694
transform 1 0 28832 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1392
timestamp 1626065694
transform 1 0 31416 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1391
timestamp 1626065694
transform 1 0 31552 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1390
timestamp 1626065694
transform 1 0 31552 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1389
timestamp 1626065694
transform 1 0 31688 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1388
timestamp 1626065694
transform 1 0 28832 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1387
timestamp 1626065694
transform 1 0 33456 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1386
timestamp 1626065694
transform 1 0 33456 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1385
timestamp 1626065694
transform 1 0 31144 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1384
timestamp 1626065694
transform 1 0 31144 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1383
timestamp 1626065694
transform 1 0 31280 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1382
timestamp 1626065694
transform 1 0 31280 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1381
timestamp 1626065694
transform 1 0 31416 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1380
timestamp 1626065694
transform 1 0 33864 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1379
timestamp 1626065694
transform 1 0 31416 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1378
timestamp 1626065694
transform 1 0 33592 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1377
timestamp 1626065694
transform 1 0 33864 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1376
timestamp 1626065694
transform 1 0 33592 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1375
timestamp 1626065694
transform 1 0 34136 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1374
timestamp 1626065694
transform 1 0 34136 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1373
timestamp 1626065694
transform 1 0 34000 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1372
timestamp 1626065694
transform 1 0 28832 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1371
timestamp 1626065694
transform 1 0 29104 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1370
timestamp 1626065694
transform 1 0 29104 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1369
timestamp 1626065694
transform 1 0 29104 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1368
timestamp 1626065694
transform 1 0 33864 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1367
timestamp 1626065694
transform 1 0 29104 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1366
timestamp 1626065694
transform 1 0 33864 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1365
timestamp 1626065694
transform 1 0 34000 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1364
timestamp 1626065694
transform 1 0 34000 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1363
timestamp 1626065694
transform 1 0 33864 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1362
timestamp 1626065694
transform 1 0 33864 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1361
timestamp 1626065694
transform 1 0 28560 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1360
timestamp 1626065694
transform 1 0 17000 0 1 17549
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1359
timestamp 1626065694
transform 1 0 17000 0 1 20133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1358
timestamp 1626065694
transform 1 0 14688 0 1 16053
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1357
timestamp 1626065694
transform 1 0 14688 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1356
timestamp 1626065694
transform 1 0 14688 0 1 16189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1355
timestamp 1626065694
transform 1 0 16592 0 1 19045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1354
timestamp 1626065694
transform 1 0 16592 0 1 20133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1353
timestamp 1626065694
transform 1 0 14552 0 1 17413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1352
timestamp 1626065694
transform 1 0 3808 0 1 20405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1351
timestamp 1626065694
transform 1 0 3672 0 1 20405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1350
timestamp 1626065694
transform 1 0 3672 0 1 17549
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1349
timestamp 1626065694
transform 1 0 2531 0 1 17893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1348
timestamp 1626065694
transform 1 0 1224 0 1 20541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1347
timestamp 1626065694
transform 1 0 3128 0 1 16053
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1346
timestamp 1626065694
transform 1 0 1224 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1345
timestamp 1626065694
transform 1 0 1224 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1344
timestamp 1626065694
transform 1 0 544 0 1 14693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1343
timestamp 1626065694
transform 1 0 1224 0 1 13877
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1342
timestamp 1626065694
transform 1 0 1224 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1341
timestamp 1626065694
transform 1 0 3128 0 1 15509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1340
timestamp 1626065694
transform 1 0 1224 0 1 15509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1339
timestamp 1626065694
transform 1 0 3128 0 1 13741
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1338
timestamp 1626065694
transform 1 0 3128 0 1 13333
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1337
timestamp 1626065694
transform 1 0 14552 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1336
timestamp 1626065694
transform 1 0 14688 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1335
timestamp 1626065694
transform 1 0 14688 0 1 13333
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1334
timestamp 1626065694
transform 1 0 14552 0 1 14693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1333
timestamp 1626065694
transform 1 0 14552 0 1 14557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1332
timestamp 1626065694
transform 1 0 14552 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1331
timestamp 1626065694
transform 1 0 1224 0 1 5445
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1330
timestamp 1626065694
transform 1 0 8704 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1329
timestamp 1626065694
transform 1 0 8704 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1328
timestamp 1626065694
transform 1 0 14552 0 1 9117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1327
timestamp 1626065694
transform 1 0 16320 0 1 8981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1326
timestamp 1626065694
transform 1 0 14688 0 1 7621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1325
timestamp 1626065694
transform 1 0 14688 0 1 10341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1324
timestamp 1626065694
transform 1 0 14688 0 1 10477
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1323
timestamp 1626065694
transform 1 0 544 0 1 7621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1322
timestamp 1626065694
transform 1 0 544 0 1 10205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1321
timestamp 1626065694
transform 1 0 1224 0 1 8709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1320
timestamp 1626065694
transform 1 0 1224 0 1 7213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1319
timestamp 1626065694
transform 1 0 1224 0 1 10477
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1318
timestamp 1626065694
transform 1 0 1224 0 1 3813
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1317
timestamp 1626065694
transform 1 0 2040 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1316
timestamp 1626065694
transform 1 0 2040 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1315
timestamp 1626065694
transform 1 0 3808 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1314
timestamp 1626065694
transform 1 0 3808 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1313
timestamp 1626065694
transform 1 0 5576 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1312
timestamp 1626065694
transform 1 0 5576 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1311
timestamp 1626065694
transform 1 0 7072 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1310
timestamp 1626065694
transform 1 0 7072 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1309
timestamp 1626065694
transform 1 0 10472 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1308
timestamp 1626065694
transform 1 0 10472 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1307
timestamp 1626065694
transform 1 0 12104 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1306
timestamp 1626065694
transform 1 0 12104 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1305
timestamp 1626065694
transform 1 0 14008 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1304
timestamp 1626065694
transform 1 0 14008 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1303
timestamp 1626065694
transform 1 0 16320 0 1 3813
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1302
timestamp 1626065694
transform 1 0 16048 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1301
timestamp 1626065694
transform 1 0 17136 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1300
timestamp 1626065694
transform 1 0 15504 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1299
timestamp 1626065694
transform 1 0 15504 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1298
timestamp 1626065694
transform 1 0 28152 0 1 9525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1297
timestamp 1626065694
transform 1 0 19040 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1296
timestamp 1626065694
transform 1 0 19040 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1295
timestamp 1626065694
transform 1 0 20264 0 1 3677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1294
timestamp 1626065694
transform 1 0 20264 0 1 1773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1293
timestamp 1626065694
transform 1 0 20808 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1292
timestamp 1626065694
transform 1 0 20808 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1291
timestamp 1626065694
transform 1 0 22168 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1290
timestamp 1626065694
transform 1 0 22168 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1289
timestamp 1626065694
transform 1 0 17408 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1288
timestamp 1626065694
transform 1 0 23120 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1287
timestamp 1626065694
transform 1 0 24208 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1286
timestamp 1626065694
transform 1 0 25432 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1285
timestamp 1626065694
transform 1 0 17408 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1284
timestamp 1626065694
transform 1 0 18224 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1283
timestamp 1626065694
transform 1 0 19584 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1282
timestamp 1626065694
transform 1 0 20536 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1281
timestamp 1626065694
transform 1 0 21760 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1280
timestamp 1626065694
transform 1 0 23936 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1279
timestamp 1626065694
transform 1 0 23936 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1278
timestamp 1626065694
transform 1 0 25704 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1277
timestamp 1626065694
transform 1 0 25704 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1276
timestamp 1626065694
transform 1 0 30464 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1275
timestamp 1626065694
transform 1 0 30464 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1274
timestamp 1626065694
transform 1 0 32096 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1273
timestamp 1626065694
transform 1 0 32096 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1272
timestamp 1626065694
transform 1 0 28968 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1271
timestamp 1626065694
transform 1 0 28968 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1270
timestamp 1626065694
transform 1 0 34000 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1269
timestamp 1626065694
transform 1 0 34000 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1268
timestamp 1626065694
transform 1 0 26520 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1267
timestamp 1626065694
transform 1 0 27608 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1266
timestamp 1626065694
transform 1 0 28696 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1265
timestamp 1626065694
transform 1 0 30056 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1264
timestamp 1626065694
transform 1 0 31280 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1263
timestamp 1626065694
transform 1 0 32368 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1262
timestamp 1626065694
transform 1 0 33456 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1261
timestamp 1626065694
transform 1 0 27336 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1260
timestamp 1626065694
transform 1 0 27336 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1259
timestamp 1626065694
transform 1 0 51272 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1258
timestamp 1626065694
transform 1 0 51272 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1257
timestamp 1626065694
transform 1 0 51272 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1256
timestamp 1626065694
transform 1 0 51272 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1255
timestamp 1626065694
transform 1 0 59976 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1254
timestamp 1626065694
transform 1 0 59976 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1253
timestamp 1626065694
transform 1 0 60656 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1252
timestamp 1626065694
transform 1 0 60656 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1251
timestamp 1626065694
transform 1 0 60792 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1250
timestamp 1626065694
transform 1 0 60792 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1249
timestamp 1626065694
transform 1 0 61880 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1248
timestamp 1626065694
transform 1 0 61880 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1247
timestamp 1626065694
transform 1 0 62424 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1246
timestamp 1626065694
transform 1 0 62424 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1245
timestamp 1626065694
transform 1 0 63104 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1244
timestamp 1626065694
transform 1 0 63104 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1243
timestamp 1626065694
transform 1 0 64464 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1242
timestamp 1626065694
transform 1 0 64464 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1241
timestamp 1626065694
transform 1 0 66232 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1240
timestamp 1626065694
transform 1 0 66232 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1239
timestamp 1626065694
transform 1 0 66912 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1238
timestamp 1626065694
transform 1 0 66912 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1237
timestamp 1626065694
transform 1 0 67456 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1236
timestamp 1626065694
transform 1 0 67456 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1235
timestamp 1626065694
transform 1 0 61608 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1234
timestamp 1626065694
transform 1 0 63920 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1233
timestamp 1626065694
transform 1 0 66640 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1232
timestamp 1626065694
transform 1 0 55624 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1231
timestamp 1626065694
transform 1 0 56168 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1230
timestamp 1626065694
transform 1 0 56168 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1229
timestamp 1626065694
transform 1 0 57392 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1228
timestamp 1626065694
transform 1 0 57392 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1227
timestamp 1626065694
transform 1 0 58208 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1226
timestamp 1626065694
transform 1 0 58208 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1225
timestamp 1626065694
transform 1 0 58344 0 1 18637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1224
timestamp 1626065694
transform 1 0 54400 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1223
timestamp 1626065694
transform 1 0 54400 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1222
timestamp 1626065694
transform 1 0 51544 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1221
timestamp 1626065694
transform 1 0 54128 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1220
timestamp 1626065694
transform 1 0 56440 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1219
timestamp 1626065694
transform 1 0 59160 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1218
timestamp 1626065694
transform 1 0 59432 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1217
timestamp 1626065694
transform 1 0 59432 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1216
timestamp 1626065694
transform 1 0 55624 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1215
timestamp 1626065694
transform 1 0 54944 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1214
timestamp 1626065694
transform 1 0 54944 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1213
timestamp 1626065694
transform 1 0 51952 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1212
timestamp 1626065694
transform 1 0 51952 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1211
timestamp 1626065694
transform 1 0 53176 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1210
timestamp 1626065694
transform 1 0 53176 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1209
timestamp 1626065694
transform 1 0 53720 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1208
timestamp 1626065694
transform 1 0 53720 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1207
timestamp 1626065694
transform 1 0 51544 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1206
timestamp 1626065694
transform 1 0 51544 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1205
timestamp 1626065694
transform 1 0 51544 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1204
timestamp 1626065694
transform 1 0 51544 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1203
timestamp 1626065694
transform 1 0 51408 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1202
timestamp 1626065694
transform 1 0 58752 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1201
timestamp 1626065694
transform 1 0 53992 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1200
timestamp 1626065694
transform 1 0 53992 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1199
timestamp 1626065694
transform 1 0 53992 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1198
timestamp 1626065694
transform 1 0 53992 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1197
timestamp 1626065694
transform 1 0 53992 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1196
timestamp 1626065694
transform 1 0 53992 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1195
timestamp 1626065694
transform 1 0 54128 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1194
timestamp 1626065694
transform 1 0 58752 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1193
timestamp 1626065694
transform 1 0 56440 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1192
timestamp 1626065694
transform 1 0 56440 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1191
timestamp 1626065694
transform 1 0 56440 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1190
timestamp 1626065694
transform 1 0 56440 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1189
timestamp 1626065694
transform 1 0 56576 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1188
timestamp 1626065694
transform 1 0 56576 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1187
timestamp 1626065694
transform 1 0 56440 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1186
timestamp 1626065694
transform 1 0 58888 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1185
timestamp 1626065694
transform 1 0 59024 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1184
timestamp 1626065694
transform 1 0 59024 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1183
timestamp 1626065694
transform 1 0 59024 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1182
timestamp 1626065694
transform 1 0 59024 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1181
timestamp 1626065694
transform 1 0 59024 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1180
timestamp 1626065694
transform 1 0 59024 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1179
timestamp 1626065694
transform 1 0 59160 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1178
timestamp 1626065694
transform 1 0 58888 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1177
timestamp 1626065694
transform 1 0 58888 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1176
timestamp 1626065694
transform 1 0 58888 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1175
timestamp 1626065694
transform 1 0 56440 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1174
timestamp 1626065694
transform 1 0 53584 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1173
timestamp 1626065694
transform 1 0 56032 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1172
timestamp 1626065694
transform 1 0 58480 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1171
timestamp 1626065694
transform 1 0 58616 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1170
timestamp 1626065694
transform 1 0 58616 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1169
timestamp 1626065694
transform 1 0 51408 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1168
timestamp 1626065694
transform 1 0 51408 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1167
timestamp 1626065694
transform 1 0 51408 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1166
timestamp 1626065694
transform 1 0 51408 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1165
timestamp 1626065694
transform 1 0 56304 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1164
timestamp 1626065694
transform 1 0 56304 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1163
timestamp 1626065694
transform 1 0 56304 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1162
timestamp 1626065694
transform 1 0 56304 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1161
timestamp 1626065694
transform 1 0 56440 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1160
timestamp 1626065694
transform 1 0 58344 0 1 14421
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1159
timestamp 1626065694
transform 1 0 53856 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1158
timestamp 1626065694
transform 1 0 53856 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1157
timestamp 1626065694
transform 1 0 53856 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1156
timestamp 1626065694
transform 1 0 53856 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1155
timestamp 1626065694
transform 1 0 53856 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1154
timestamp 1626065694
transform 1 0 53856 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1153
timestamp 1626065694
transform 1 0 63648 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1152
timestamp 1626065694
transform 1 0 63648 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1151
timestamp 1626065694
transform 1 0 64056 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1150
timestamp 1626065694
transform 1 0 64056 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1149
timestamp 1626065694
transform 1 0 64056 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1148
timestamp 1626065694
transform 1 0 64056 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1147
timestamp 1626065694
transform 1 0 63920 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1146
timestamp 1626065694
transform 1 0 63648 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1145
timestamp 1626065694
transform 1 0 66232 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1144
timestamp 1626065694
transform 1 0 66232 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1143
timestamp 1626065694
transform 1 0 66504 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1142
timestamp 1626065694
transform 1 0 66504 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1141
timestamp 1626065694
transform 1 0 66504 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1140
timestamp 1626065694
transform 1 0 66504 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1139
timestamp 1626065694
transform 1 0 66640 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1138
timestamp 1626065694
transform 1 0 66096 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1137
timestamp 1626065694
transform 1 0 66096 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1136
timestamp 1626065694
transform 1 0 66368 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1135
timestamp 1626065694
transform 1 0 66368 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1134
timestamp 1626065694
transform 1 0 60928 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1133
timestamp 1626065694
transform 1 0 63512 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1132
timestamp 1626065694
transform 1 0 65960 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1131
timestamp 1626065694
transform 1 0 66232 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1130
timestamp 1626065694
transform 1 0 66232 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1129
timestamp 1626065694
transform 1 0 61064 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1128
timestamp 1626065694
transform 1 0 61064 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1127
timestamp 1626065694
transform 1 0 61200 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1126
timestamp 1626065694
transform 1 0 61200 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1125
timestamp 1626065694
transform 1 0 61200 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1124
timestamp 1626065694
transform 1 0 61200 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1123
timestamp 1626065694
transform 1 0 63784 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1122
timestamp 1626065694
transform 1 0 63784 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1121
timestamp 1626065694
transform 1 0 63920 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1120
timestamp 1626065694
transform 1 0 63920 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1119
timestamp 1626065694
transform 1 0 63784 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1118
timestamp 1626065694
transform 1 0 63784 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1117
timestamp 1626065694
transform 1 0 61336 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1116
timestamp 1626065694
transform 1 0 61336 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1115
timestamp 1626065694
transform 1 0 61336 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1114
timestamp 1626065694
transform 1 0 61336 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1113
timestamp 1626065694
transform 1 0 61336 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1112
timestamp 1626065694
transform 1 0 61336 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1111
timestamp 1626065694
transform 1 0 61472 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1110
timestamp 1626065694
transform 1 0 61472 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1109
timestamp 1626065694
transform 1 0 61608 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1108
timestamp 1626065694
transform 1 0 63648 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1107
timestamp 1626065694
transform 1 0 44064 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1106
timestamp 1626065694
transform 1 0 43248 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1105
timestamp 1626065694
transform 1 0 43248 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1104
timestamp 1626065694
transform 1 0 43384 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1103
timestamp 1626065694
transform 1 0 43384 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1102
timestamp 1626065694
transform 1 0 44472 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1101
timestamp 1626065694
transform 1 0 44472 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1100
timestamp 1626065694
transform 1 0 45696 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1099
timestamp 1626065694
transform 1 0 45696 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1098
timestamp 1626065694
transform 1 0 46920 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1097
timestamp 1626065694
transform 1 0 46920 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1096
timestamp 1626065694
transform 1 0 47464 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1095
timestamp 1626065694
transform 1 0 47464 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1094
timestamp 1626065694
transform 1 0 48144 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1093
timestamp 1626065694
transform 1 0 48144 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1092
timestamp 1626065694
transform 1 0 46648 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1091
timestamp 1626065694
transform 1 0 49912 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1090
timestamp 1626065694
transform 1 0 49912 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1089
timestamp 1626065694
transform 1 0 48960 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1088
timestamp 1626065694
transform 1 0 42432 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1087
timestamp 1626065694
transform 1 0 38216 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1086
timestamp 1626065694
transform 1 0 41616 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1085
timestamp 1626065694
transform 1 0 38760 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1084
timestamp 1626065694
transform 1 0 34544 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1083
timestamp 1626065694
transform 1 0 39168 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1082
timestamp 1626065694
transform 1 0 37264 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1081
timestamp 1626065694
transform 1 0 38760 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1080
timestamp 1626065694
transform 1 0 39440 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1079
timestamp 1626065694
transform 1 0 39440 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1078
timestamp 1626065694
transform 1 0 39984 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1077
timestamp 1626065694
transform 1 0 39984 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1076
timestamp 1626065694
transform 1 0 40664 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1075
timestamp 1626065694
transform 1 0 40664 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1074
timestamp 1626065694
transform 1 0 41208 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1073
timestamp 1626065694
transform 1 0 41208 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1072
timestamp 1626065694
transform 1 0 42024 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1071
timestamp 1626065694
transform 1 0 42024 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1070
timestamp 1626065694
transform 1 0 42432 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1069
timestamp 1626065694
transform 1 0 35632 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1068
timestamp 1626065694
transform 1 0 34544 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1067
timestamp 1626065694
transform 1 0 35632 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1066
timestamp 1626065694
transform 1 0 36448 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1065
timestamp 1626065694
transform 1 0 38216 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1064
timestamp 1626065694
transform 1 0 37264 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1063
timestamp 1626065694
transform 1 0 41480 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1062
timestamp 1626065694
transform 1 0 38760 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1061
timestamp 1626065694
transform 1 0 38760 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1060
timestamp 1626065694
transform 1 0 41616 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1059
timestamp 1626065694
transform 1 0 41480 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1058
timestamp 1626065694
transform 1 0 38896 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1057
timestamp 1626065694
transform 1 0 41072 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1056
timestamp 1626065694
transform 1 0 41072 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1055
timestamp 1626065694
transform 1 0 41344 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1054
timestamp 1626065694
transform 1 0 41344 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1053
timestamp 1626065694
transform 1 0 41344 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1052
timestamp 1626065694
transform 1 0 36040 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1051
timestamp 1626065694
transform 1 0 38488 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1050
timestamp 1626065694
transform 1 0 41072 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1049
timestamp 1626065694
transform 1 0 41344 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1048
timestamp 1626065694
transform 1 0 41208 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1047
timestamp 1626065694
transform 1 0 41208 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1046
timestamp 1626065694
transform 1 0 41480 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1045
timestamp 1626065694
transform 1 0 36448 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1044
timestamp 1626065694
transform 1 0 36448 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1043
timestamp 1626065694
transform 1 0 41480 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1042
timestamp 1626065694
transform 1 0 36176 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1041
timestamp 1626065694
transform 1 0 36176 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1040
timestamp 1626065694
transform 1 0 36584 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1039
timestamp 1626065694
transform 1 0 36584 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1038
timestamp 1626065694
transform 1 0 36584 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1037
timestamp 1626065694
transform 1 0 36584 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1036
timestamp 1626065694
transform 1 0 36312 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1035
timestamp 1626065694
transform 1 0 36448 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1034
timestamp 1626065694
transform 1 0 38896 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1033
timestamp 1626065694
transform 1 0 38896 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1032
timestamp 1626065694
transform 1 0 36448 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1031
timestamp 1626065694
transform 1 0 36312 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1030
timestamp 1626065694
transform 1 0 38624 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1029
timestamp 1626065694
transform 1 0 38624 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1028
timestamp 1626065694
transform 1 0 39032 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1027
timestamp 1626065694
transform 1 0 39032 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1026
timestamp 1626065694
transform 1 0 39032 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1025
timestamp 1626065694
transform 1 0 39032 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1024
timestamp 1626065694
transform 1 0 36448 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1023
timestamp 1626065694
transform 1 0 38896 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1022
timestamp 1626065694
transform 1 0 41480 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1021
timestamp 1626065694
transform 1 0 41480 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1020
timestamp 1626065694
transform 1 0 39168 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1019
timestamp 1626065694
transform 1 0 43792 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1018
timestamp 1626065694
transform 1 0 43520 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1017
timestamp 1626065694
transform 1 0 45968 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1016
timestamp 1626065694
transform 1 0 48280 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1015
timestamp 1626065694
transform 1 0 51000 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1014
timestamp 1626065694
transform 1 0 46648 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1013
timestamp 1626065694
transform 1 0 46512 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1012
timestamp 1626065694
transform 1 0 48824 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1011
timestamp 1626065694
transform 1 0 48824 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1010
timestamp 1626065694
transform 1 0 48824 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1009
timestamp 1626065694
transform 1 0 48824 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1008
timestamp 1626065694
transform 1 0 46512 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1007
timestamp 1626065694
transform 1 0 46512 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1006
timestamp 1626065694
transform 1 0 49096 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1005
timestamp 1626065694
transform 1 0 49096 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1004
timestamp 1626065694
transform 1 0 48960 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1003
timestamp 1626065694
transform 1 0 51136 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1002
timestamp 1626065694
transform 1 0 51136 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1001
timestamp 1626065694
transform 1 0 44064 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1000
timestamp 1626065694
transform 1 0 46240 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_999
timestamp 1626065694
transform 1 0 46240 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_998
timestamp 1626065694
transform 1 0 46376 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_997
timestamp 1626065694
transform 1 0 46376 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_996
timestamp 1626065694
transform 1 0 46240 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_995
timestamp 1626065694
transform 1 0 46240 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_994
timestamp 1626065694
transform 1 0 44064 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_993
timestamp 1626065694
transform 1 0 43928 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_992
timestamp 1626065694
transform 1 0 44064 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_991
timestamp 1626065694
transform 1 0 43384 0 1 11429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_990
timestamp 1626065694
transform 1 0 43384 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_989
timestamp 1626065694
transform 1 0 44064 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_988
timestamp 1626065694
transform 1 0 46512 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_987
timestamp 1626065694
transform 1 0 46512 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_986
timestamp 1626065694
transform 1 0 46512 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_985
timestamp 1626065694
transform 1 0 48688 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_984
timestamp 1626065694
transform 1 0 48688 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_983
timestamp 1626065694
transform 1 0 48960 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_982
timestamp 1626065694
transform 1 0 48960 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_981
timestamp 1626065694
transform 1 0 43792 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_980
timestamp 1626065694
transform 1 0 43792 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_979
timestamp 1626065694
transform 1 0 48824 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_978
timestamp 1626065694
transform 1 0 48824 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_977
timestamp 1626065694
transform 1 0 43928 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_976
timestamp 1626065694
transform 1 0 43928 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_975
timestamp 1626065694
transform 1 0 43792 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_974
timestamp 1626065694
transform 1 0 40800 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_973
timestamp 1626065694
transform 1 0 40800 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_972
timestamp 1626065694
transform 1 0 39168 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_971
timestamp 1626065694
transform 1 0 39712 0 1 2317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_970
timestamp 1626065694
transform 1 0 39712 0 1 549
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_969
timestamp 1626065694
transform 1 0 39168 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_968
timestamp 1626065694
transform 1 0 35768 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_967
timestamp 1626065694
transform 1 0 35768 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_966
timestamp 1626065694
transform 1 0 42432 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_965
timestamp 1626065694
transform 1 0 42432 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_964
timestamp 1626065694
transform 1 0 37400 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_963
timestamp 1626065694
transform 1 0 37400 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_962
timestamp 1626065694
transform 1 0 34544 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_961
timestamp 1626065694
transform 1 0 35904 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_960
timestamp 1626065694
transform 1 0 36992 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_959
timestamp 1626065694
transform 1 0 38080 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_958
timestamp 1626065694
transform 1 0 39440 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_957
timestamp 1626065694
transform 1 0 40664 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_956
timestamp 1626065694
transform 1 0 41752 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_955
timestamp 1626065694
transform 1 0 49096 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_954
timestamp 1626065694
transform 1 0 49096 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_953
timestamp 1626065694
transform 1 0 44200 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_952
timestamp 1626065694
transform 1 0 44200 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_951
timestamp 1626065694
transform 1 0 45696 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_950
timestamp 1626065694
transform 1 0 45696 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_949
timestamp 1626065694
transform 1 0 47328 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_948
timestamp 1626065694
transform 1 0 47328 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_947
timestamp 1626065694
transform 1 0 50728 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_946
timestamp 1626065694
transform 1 0 50728 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_945
timestamp 1626065694
transform 1 0 42840 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_944
timestamp 1626065694
transform 1 0 43928 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_943
timestamp 1626065694
transform 1 0 45288 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_942
timestamp 1626065694
transform 1 0 46376 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_941
timestamp 1626065694
transform 1 0 47600 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_940
timestamp 1626065694
transform 1 0 48688 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_939
timestamp 1626065694
transform 1 0 49776 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_938
timestamp 1626065694
transform 1 0 51136 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_937
timestamp 1626065694
transform 1 0 59432 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_936
timestamp 1626065694
transform 1 0 59432 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_935
timestamp 1626065694
transform 1 0 52224 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_934
timestamp 1626065694
transform 1 0 53312 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_933
timestamp 1626065694
transform 1 0 54400 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_932
timestamp 1626065694
transform 1 0 55760 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_931
timestamp 1626065694
transform 1 0 56984 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_930
timestamp 1626065694
transform 1 0 58072 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_929
timestamp 1626065694
transform 1 0 59160 0 1 2861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_928
timestamp 1626065694
transform 1 0 57528 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_927
timestamp 1626065694
transform 1 0 57528 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_926
timestamp 1626065694
transform 1 0 55488 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_925
timestamp 1626065694
transform 1 0 55488 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_924
timestamp 1626065694
transform 1 0 52496 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_923
timestamp 1626065694
transform 1 0 52496 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_922
timestamp 1626065694
transform 1 0 54128 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_921
timestamp 1626065694
transform 1 0 54128 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_920
timestamp 1626065694
transform 1 0 64328 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_919
timestamp 1626065694
transform 1 0 64328 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_918
timestamp 1626065694
transform 1 0 65824 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_917
timestamp 1626065694
transform 1 0 65824 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_916
timestamp 1626065694
transform 1 0 60792 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_915
timestamp 1626065694
transform 1 0 67592 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_914
timestamp 1626065694
transform 1 0 67592 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_913
timestamp 1626065694
transform 1 0 60792 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_912
timestamp 1626065694
transform 1 0 62560 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_911
timestamp 1626065694
transform 1 0 62560 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_910
timestamp 1626065694
transform 1 0 115192 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_909
timestamp 1626065694
transform 1 0 115328 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_908
timestamp 1626065694
transform 1 0 117640 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_907
timestamp 1626065694
transform 1 0 118592 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_906
timestamp 1626065694
transform 1 0 114648 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_905
timestamp 1626065694
transform 1 0 116008 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_904
timestamp 1626065694
transform 1 0 114240 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_903
timestamp 1626065694
transform 1 0 118184 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_902
timestamp 1626065694
transform 1 0 119000 0 1 20949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_901
timestamp 1626065694
transform 1 0 114648 0 1 31285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_900
timestamp 1626065694
transform 1 0 114240 0 1 31285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_899
timestamp 1626065694
transform 1 0 119272 0 1 26525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_898
timestamp 1626065694
transform 1 0 119272 0 1 25845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_897
timestamp 1626065694
transform 1 0 119272 0 1 26661
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_896
timestamp 1626065694
transform 1 0 119272 0 1 27205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_895
timestamp 1626065694
transform 1 0 135320 0 1 37405
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_894
timestamp 1626065694
transform 1 0 135320 0 1 40805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_893
timestamp 1626065694
transform 1 0 135320 0 1 39037
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_892
timestamp 1626065694
transform 1 0 135320 0 1 32237
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_891
timestamp 1626065694
transform 1 0 135320 0 1 33869
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_890
timestamp 1626065694
transform 1 0 135320 0 1 35501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_889
timestamp 1626065694
transform 1 0 114648 0 1 36453
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_888
timestamp 1626065694
transform 1 0 115192 0 1 36453
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_887
timestamp 1626065694
transform 1 0 114240 0 1 36453
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_886
timestamp 1626065694
transform 1 0 115464 0 1 36453
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_885
timestamp 1626065694
transform 1 0 114648 0 1 39581
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_884
timestamp 1626065694
transform 1 0 115056 0 1 37949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_883
timestamp 1626065694
transform 1 0 114648 0 1 41077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_882
timestamp 1626065694
transform 1 0 114648 0 1 40805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_881
timestamp 1626065694
transform 1 0 114648 0 1 36725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_880
timestamp 1626065694
transform 1 0 115056 0 1 37677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_879
timestamp 1626065694
transform 1 0 114648 0 1 39989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_878
timestamp 1626065694
transform 1 0 115192 0 1 36725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_877
timestamp 1626065694
transform 1 0 115192 0 1 40805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_876
timestamp 1626065694
transform 1 0 115192 0 1 41077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_875
timestamp 1626065694
transform 1 0 115328 0 1 40805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_874
timestamp 1626065694
transform 1 0 114648 0 1 40397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_873
timestamp 1626065694
transform 1 0 114648 0 1 40669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_872
timestamp 1626065694
transform 1 0 115328 0 1 41077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_871
timestamp 1626065694
transform 1 0 115328 0 1 40397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_870
timestamp 1626065694
transform 1 0 115328 0 1 40669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_869
timestamp 1626065694
transform 1 0 114240 0 1 39853
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_868
timestamp 1626065694
transform 1 0 115192 0 1 40261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_867
timestamp 1626065694
transform 1 0 114240 0 1 39581
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_866
timestamp 1626065694
transform 1 0 114240 0 1 39989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_865
timestamp 1626065694
transform 1 0 114240 0 1 40261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_864
timestamp 1626065694
transform 1 0 115328 0 1 40125
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_863
timestamp 1626065694
transform 1 0 115464 0 1 37949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_862
timestamp 1626065694
transform 1 0 115464 0 1 37677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_861
timestamp 1626065694
transform 1 0 115464 0 1 39173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_860
timestamp 1626065694
transform 1 0 115464 0 1 38901
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_859
timestamp 1626065694
transform 1 0 115600 0 1 41485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_858
timestamp 1626065694
transform 1 0 114240 0 1 36861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_857
timestamp 1626065694
transform 1 0 114240 0 1 37133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_856
timestamp 1626065694
transform 1 0 114240 0 1 36725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_855
timestamp 1626065694
transform 1 0 114648 0 1 40261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_854
timestamp 1626065694
transform 1 0 115600 0 1 41213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_853
timestamp 1626065694
transform 1 0 115464 0 1 40805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_852
timestamp 1626065694
transform 1 0 115464 0 1 41077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_851
timestamp 1626065694
transform 1 0 114648 0 1 39853
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_850
timestamp 1626065694
transform 1 0 115464 0 1 36725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_849
timestamp 1626065694
transform 1 0 116008 0 1 41077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_848
timestamp 1626065694
transform 1 0 116008 0 1 40805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_847
timestamp 1626065694
transform 1 0 116008 0 1 41213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_846
timestamp 1626065694
transform 1 0 116008 0 1 41485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_845
timestamp 1626065694
transform 1 0 115600 0 1 37133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_844
timestamp 1626065694
transform 1 0 115600 0 1 36861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_843
timestamp 1626065694
transform 1 0 114376 0 1 38357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_842
timestamp 1626065694
transform 1 0 116008 0 1 38765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_841
timestamp 1626065694
transform 1 0 116008 0 1 38493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_840
timestamp 1626065694
transform 1 0 116008 0 1 38901
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_839
timestamp 1626065694
transform 1 0 116008 0 1 39173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_838
timestamp 1626065694
transform 1 0 114376 0 1 38085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_837
timestamp 1626065694
transform 1 0 115872 0 1 38357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_836
timestamp 1626065694
transform 1 0 115872 0 1 38085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_835
timestamp 1626065694
transform 1 0 114648 0 1 38085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_834
timestamp 1626065694
transform 1 0 114648 0 1 38357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_833
timestamp 1626065694
transform 1 0 114648 0 1 37949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_832
timestamp 1626065694
transform 1 0 114648 0 1 37677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_831
timestamp 1626065694
transform 1 0 114784 0 1 41485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_830
timestamp 1626065694
transform 1 0 114376 0 1 37269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_829
timestamp 1626065694
transform 1 0 114376 0 1 37541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_828
timestamp 1626065694
transform 1 0 114376 0 1 40805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_827
timestamp 1626065694
transform 1 0 114376 0 1 41077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_826
timestamp 1626065694
transform 1 0 114376 0 1 40669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_825
timestamp 1626065694
transform 1 0 115872 0 1 39309
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_824
timestamp 1626065694
transform 1 0 115872 0 1 39581
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_823
timestamp 1626065694
transform 1 0 114376 0 1 40397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_822
timestamp 1626065694
transform 1 0 114784 0 1 41213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_821
timestamp 1626065694
transform 1 0 115192 0 1 39581
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_820
timestamp 1626065694
transform 1 0 115192 0 1 39853
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_819
timestamp 1626065694
transform 1 0 115192 0 1 38357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_818
timestamp 1626065694
transform 1 0 115192 0 1 38085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_817
timestamp 1626065694
transform 1 0 115872 0 1 37133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_816
timestamp 1626065694
transform 1 0 115872 0 1 36861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_815
timestamp 1626065694
transform 1 0 115872 0 1 37269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_814
timestamp 1626065694
transform 1 0 115872 0 1 37541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_813
timestamp 1626065694
transform 1 0 115328 0 1 38357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_812
timestamp 1626065694
transform 1 0 116008 0 1 37949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_811
timestamp 1626065694
transform 1 0 116008 0 1 37677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_810
timestamp 1626065694
transform 1 0 115328 0 1 38085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_809
timestamp 1626065694
transform 1 0 114784 0 1 37133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_808
timestamp 1626065694
transform 1 0 114784 0 1 36861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_807
timestamp 1626065694
transform 1 0 114376 0 1 41485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_806
timestamp 1626065694
transform 1 0 114376 0 1 41213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_805
timestamp 1626065694
transform 1 0 114784 0 1 37269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_804
timestamp 1626065694
transform 1 0 114784 0 1 37541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_803
timestamp 1626065694
transform 1 0 114240 0 1 37677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_802
timestamp 1626065694
transform 1 0 114240 0 1 37949
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_801
timestamp 1626065694
transform 1 0 109344 0 1 40261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_800
timestamp 1626065694
transform 1 0 109344 0 1 39853
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_799
timestamp 1626065694
transform 1 0 109480 0 1 38085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_798
timestamp 1626065694
transform 1 0 109480 0 1 37813
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_797
timestamp 1626065694
transform 1 0 109480 0 1 40261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_796
timestamp 1626065694
transform 1 0 109480 0 1 40533
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_795
timestamp 1626065694
transform 1 0 109480 0 1 39037
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_794
timestamp 1626065694
transform 1 0 109480 0 1 39309
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_793
timestamp 1626065694
transform 1 0 109480 0 1 34685
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_792
timestamp 1626065694
transform 1 0 109480 0 1 34413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_791
timestamp 1626065694
transform 1 0 109344 0 1 31557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_790
timestamp 1626065694
transform 1 0 109480 0 1 31557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_789
timestamp 1626065694
transform 1 0 109480 0 1 31829
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_788
timestamp 1626065694
transform 1 0 109344 0 1 34685
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_787
timestamp 1626065694
transform 1 0 109344 0 1 34957
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_786
timestamp 1626065694
transform 1 0 109480 0 1 34141
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_785
timestamp 1626065694
transform 1 0 109480 0 1 33869
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_784
timestamp 1626065694
transform 1 0 114784 0 1 36045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_783
timestamp 1626065694
transform 1 0 114240 0 1 33597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_782
timestamp 1626065694
transform 1 0 114240 0 1 33325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_781
timestamp 1626065694
transform 1 0 114240 0 1 33733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_780
timestamp 1626065694
transform 1 0 114240 0 1 34005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_779
timestamp 1626065694
transform 1 0 114784 0 1 36317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_778
timestamp 1626065694
transform 1 0 116008 0 1 34413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_777
timestamp 1626065694
transform 1 0 116008 0 1 34141
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_776
timestamp 1626065694
transform 1 0 115328 0 1 33733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_775
timestamp 1626065694
transform 1 0 115192 0 1 33189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_774
timestamp 1626065694
transform 1 0 115192 0 1 34413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_773
timestamp 1626065694
transform 1 0 115192 0 1 34141
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_772
timestamp 1626065694
transform 1 0 116008 0 1 33733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_771
timestamp 1626065694
transform 1 0 116008 0 1 34005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_770
timestamp 1626065694
transform 1 0 116008 0 1 33597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_769
timestamp 1626065694
transform 1 0 116008 0 1 33325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_768
timestamp 1626065694
transform 1 0 115464 0 1 35909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_767
timestamp 1626065694
transform 1 0 115464 0 1 35637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_766
timestamp 1626065694
transform 1 0 115464 0 1 34821
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_765
timestamp 1626065694
transform 1 0 115464 0 1 35229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_764
timestamp 1626065694
transform 1 0 115872 0 1 35365
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_763
timestamp 1626065694
transform 1 0 115872 0 1 35637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_762
timestamp 1626065694
transform 1 0 114648 0 1 32373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_761
timestamp 1626065694
transform 1 0 115600 0 1 32781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_760
timestamp 1626065694
transform 1 0 115600 0 1 32509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_759
timestamp 1626065694
transform 1 0 115600 0 1 33325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_758
timestamp 1626065694
transform 1 0 115600 0 1 34005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_757
timestamp 1626065694
transform 1 0 115600 0 1 33733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_756
timestamp 1626065694
transform 1 0 115600 0 1 33597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_755
timestamp 1626065694
transform 1 0 114648 0 1 32101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_754
timestamp 1626065694
transform 1 0 114240 0 1 32373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_753
timestamp 1626065694
transform 1 0 116008 0 1 34821
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_752
timestamp 1626065694
transform 1 0 116008 0 1 34549
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_751
timestamp 1626065694
transform 1 0 115872 0 1 34957
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_750
timestamp 1626065694
transform 1 0 115872 0 1 35229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_749
timestamp 1626065694
transform 1 0 114240 0 1 32101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_748
timestamp 1626065694
transform 1 0 115328 0 1 32101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_747
timestamp 1626065694
transform 1 0 115328 0 1 32373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_746
timestamp 1626065694
transform 1 0 114648 0 1 31557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_745
timestamp 1626065694
transform 1 0 114240 0 1 34413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_744
timestamp 1626065694
transform 1 0 115600 0 1 34413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_743
timestamp 1626065694
transform 1 0 115600 0 1 34141
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_742
timestamp 1626065694
transform 1 0 115872 0 1 31421
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_741
timestamp 1626065694
transform 1 0 115872 0 1 31693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_740
timestamp 1626065694
transform 1 0 115192 0 1 32917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_739
timestamp 1626065694
transform 1 0 114784 0 1 31693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_738
timestamp 1626065694
transform 1 0 114240 0 1 34141
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_737
timestamp 1626065694
transform 1 0 114784 0 1 34005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_736
timestamp 1626065694
transform 1 0 115056 0 1 33597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_735
timestamp 1626065694
transform 1 0 115056 0 1 33325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_734
timestamp 1626065694
transform 1 0 114648 0 1 35637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_733
timestamp 1626065694
transform 1 0 114648 0 1 35909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_732
timestamp 1626065694
transform 1 0 114784 0 1 32781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_731
timestamp 1626065694
transform 1 0 114784 0 1 32509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_730
timestamp 1626065694
transform 1 0 114784 0 1 32917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_729
timestamp 1626065694
transform 1 0 114784 0 1 33189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_728
timestamp 1626065694
transform 1 0 114784 0 1 33733
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_727
timestamp 1626065694
transform 1 0 114376 0 1 36045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_726
timestamp 1626065694
transform 1 0 114376 0 1 36317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_725
timestamp 1626065694
transform 1 0 115872 0 1 32101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_724
timestamp 1626065694
transform 1 0 115872 0 1 32373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_723
timestamp 1626065694
transform 1 0 116008 0 1 36317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_722
timestamp 1626065694
transform 1 0 116008 0 1 36045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_721
timestamp 1626065694
transform 1 0 114240 0 1 35909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_720
timestamp 1626065694
transform 1 0 115192 0 1 36045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_719
timestamp 1626065694
transform 1 0 115192 0 1 36317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_718
timestamp 1626065694
transform 1 0 115328 0 1 36045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_717
timestamp 1626065694
transform 1 0 115872 0 1 32781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_716
timestamp 1626065694
transform 1 0 115872 0 1 32509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_715
timestamp 1626065694
transform 1 0 115872 0 1 32917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_714
timestamp 1626065694
transform 1 0 115872 0 1 33189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_713
timestamp 1626065694
transform 1 0 114376 0 1 32781
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_712
timestamp 1626065694
transform 1 0 114376 0 1 32509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_711
timestamp 1626065694
transform 1 0 114376 0 1 32917
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_710
timestamp 1626065694
transform 1 0 114376 0 1 33189
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_709
timestamp 1626065694
transform 1 0 114240 0 1 35637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_708
timestamp 1626065694
transform 1 0 115192 0 1 32101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_707
timestamp 1626065694
transform 1 0 114240 0 1 31557
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_706
timestamp 1626065694
transform 1 0 114784 0 1 31965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_705
timestamp 1626065694
transform 1 0 115192 0 1 32373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_704
timestamp 1626065694
transform 1 0 114376 0 1 31693
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_703
timestamp 1626065694
transform 1 0 114376 0 1 31965
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_702
timestamp 1626065694
transform 1 0 114648 0 1 33325
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_701
timestamp 1626065694
transform 1 0 114648 0 1 34413
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_700
timestamp 1626065694
transform 1 0 114648 0 1 34141
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_699
timestamp 1626065694
transform 1 0 115328 0 1 36317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_698
timestamp 1626065694
transform 1 0 114648 0 1 33597
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_697
timestamp 1626065694
transform 1 0 115328 0 1 34005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_696
timestamp 1626065694
transform 1 0 114240 0 1 26117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_695
timestamp 1626065694
transform 1 0 116008 0 1 26117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_694
timestamp 1626065694
transform 1 0 114648 0 1 26117
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_693
timestamp 1626065694
transform 1 0 114784 0 1 28837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_692
timestamp 1626065694
transform 1 0 115328 0 1 29653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_691
timestamp 1626065694
transform 1 0 115328 0 1 29381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_690
timestamp 1626065694
transform 1 0 115872 0 1 29789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_689
timestamp 1626065694
transform 1 0 115872 0 1 30061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_688
timestamp 1626065694
transform 1 0 115872 0 1 29653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_687
timestamp 1626065694
transform 1 0 115872 0 1 29381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_686
timestamp 1626065694
transform 1 0 114376 0 1 27341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_685
timestamp 1626065694
transform 1 0 114376 0 1 27613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_684
timestamp 1626065694
transform 1 0 114784 0 1 27341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_683
timestamp 1626065694
transform 1 0 114784 0 1 27613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_682
timestamp 1626065694
transform 1 0 115464 0 1 30469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_681
timestamp 1626065694
transform 1 0 115464 0 1 30197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_680
timestamp 1626065694
transform 1 0 115872 0 1 26661
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_679
timestamp 1626065694
transform 1 0 115872 0 1 26933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_678
timestamp 1626065694
transform 1 0 115872 0 1 26525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_677
timestamp 1626065694
transform 1 0 115872 0 1 26253
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_676
timestamp 1626065694
transform 1 0 115464 0 1 26525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_675
timestamp 1626065694
transform 1 0 115464 0 1 26253
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_674
timestamp 1626065694
transform 1 0 115464 0 1 30877
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_673
timestamp 1626065694
transform 1 0 115464 0 1 31149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_672
timestamp 1626065694
transform 1 0 115328 0 1 28973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_671
timestamp 1626065694
transform 1 0 115328 0 1 29245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_670
timestamp 1626065694
transform 1 0 115872 0 1 28837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_669
timestamp 1626065694
transform 1 0 115872 0 1 28565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_668
timestamp 1626065694
transform 1 0 116008 0 1 28973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_667
timestamp 1626065694
transform 1 0 116008 0 1 29245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_666
timestamp 1626065694
transform 1 0 117776 0 1 27205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_665
timestamp 1626065694
transform 1 0 117776 0 1 26661
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_664
timestamp 1626065694
transform 1 0 115600 0 1 27205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_663
timestamp 1626065694
transform 1 0 117640 0 1 26389
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_662
timestamp 1626065694
transform 1 0 116008 0 1 30197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_661
timestamp 1626065694
transform 1 0 116008 0 1 30469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_660
timestamp 1626065694
transform 1 0 115600 0 1 26933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_659
timestamp 1626065694
transform 1 0 114784 0 1 28429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_658
timestamp 1626065694
transform 1 0 114648 0 1 30061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_657
timestamp 1626065694
transform 1 0 114648 0 1 29789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_656
timestamp 1626065694
transform 1 0 114376 0 1 28429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_655
timestamp 1626065694
transform 1 0 114376 0 1 28157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_654
timestamp 1626065694
transform 1 0 114376 0 1 28565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_653
timestamp 1626065694
transform 1 0 114376 0 1 28837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_652
timestamp 1626065694
transform 1 0 118728 0 1 26661
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_651
timestamp 1626065694
transform 1 0 118864 0 1 27205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_650
timestamp 1626065694
transform 1 0 119000 0 1 26525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_649
timestamp 1626065694
transform 1 0 114648 0 1 29381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_648
timestamp 1626065694
transform 1 0 114648 0 1 29653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_647
timestamp 1626065694
transform 1 0 114648 0 1 29245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_646
timestamp 1626065694
transform 1 0 114648 0 1 28973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_645
timestamp 1626065694
transform 1 0 115872 0 1 28429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_644
timestamp 1626065694
transform 1 0 115872 0 1 28157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_643
timestamp 1626065694
transform 1 0 114784 0 1 28157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_642
timestamp 1626065694
transform 1 0 115736 0 1 27205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_641
timestamp 1626065694
transform 1 0 114784 0 1 27749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_640
timestamp 1626065694
transform 1 0 114784 0 1 28021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_639
timestamp 1626065694
transform 1 0 115736 0 1 26797
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_638
timestamp 1626065694
transform 1 0 117640 0 1 26797
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_637
timestamp 1626065694
transform 1 0 117640 0 1 27205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_636
timestamp 1626065694
transform 1 0 115192 0 1 28565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_635
timestamp 1626065694
transform 1 0 115192 0 1 28837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_634
timestamp 1626065694
transform 1 0 115464 0 1 29381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_633
timestamp 1626065694
transform 1 0 115464 0 1 29653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_632
timestamp 1626065694
transform 1 0 115056 0 1 29245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_631
timestamp 1626065694
transform 1 0 115056 0 1 28973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_630
timestamp 1626065694
transform 1 0 114376 0 1 27749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_629
timestamp 1626065694
transform 1 0 115192 0 1 27749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_628
timestamp 1626065694
transform 1 0 115192 0 1 28021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_627
timestamp 1626065694
transform 1 0 115600 0 1 28429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_626
timestamp 1626065694
transform 1 0 114376 0 1 28021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_625
timestamp 1626065694
transform 1 0 115872 0 1 30605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_624
timestamp 1626065694
transform 1 0 115872 0 1 30877
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_623
timestamp 1626065694
transform 1 0 114784 0 1 28565
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_622
timestamp 1626065694
transform 1 0 114240 0 1 29381
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_621
timestamp 1626065694
transform 1 0 114240 0 1 29653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_620
timestamp 1626065694
transform 1 0 114240 0 1 29245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_619
timestamp 1626065694
transform 1 0 115600 0 1 28157
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_618
timestamp 1626065694
transform 1 0 114240 0 1 28973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_617
timestamp 1626065694
transform 1 0 118184 0 1 26389
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_616
timestamp 1626065694
transform 1 0 118184 0 1 26661
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_615
timestamp 1626065694
transform 1 0 118184 0 1 27205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_614
timestamp 1626065694
transform 1 0 114240 0 1 30061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_613
timestamp 1626065694
transform 1 0 114240 0 1 29789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_612
timestamp 1626065694
transform 1 0 109344 0 1 31149
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_611
timestamp 1626065694
transform 1 0 109344 0 1 29925
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_610
timestamp 1626065694
transform 1 0 109344 0 1 30197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_609
timestamp 1626065694
transform 1 0 109344 0 1 26253
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_608
timestamp 1626065694
transform 1 0 109344 0 1 26389
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_607
timestamp 1626065694
transform 1 0 109344 0 1 30605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_606
timestamp 1626065694
transform 1 0 109344 0 1 30333
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_605
timestamp 1626065694
transform 1 0 109344 0 1 26661
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_604
timestamp 1626065694
transform 1 0 109344 0 1 25981
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_603
timestamp 1626065694
transform 1 0 109480 0 1 22445
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_602
timestamp 1626065694
transform 1 0 109344 0 1 21221
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_601
timestamp 1626065694
transform 1 0 109344 0 1 21493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_600
timestamp 1626065694
transform 1 0 109344 0 1 22037
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_599
timestamp 1626065694
transform 1 0 109344 0 1 23125
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_598
timestamp 1626065694
transform 1 0 109480 0 1 22717
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_597
timestamp 1626065694
transform 1 0 109344 0 1 22309
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_596
timestamp 1626065694
transform 1 0 109344 0 1 22853
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_595
timestamp 1626065694
transform 1 0 115056 0 1 25709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_594
timestamp 1626065694
transform 1 0 115056 0 1 25437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_593
timestamp 1626065694
transform 1 0 115056 0 1 24893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_592
timestamp 1626065694
transform 1 0 115056 0 1 22581
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_591
timestamp 1626065694
transform 1 0 115056 0 1 22309
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_590
timestamp 1626065694
transform 1 0 115056 0 1 21765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_589
timestamp 1626065694
transform 1 0 115056 0 1 21493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_588
timestamp 1626065694
transform 1 0 115056 0 1 24621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_587
timestamp 1626065694
transform 1 0 115600 0 1 24077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_586
timestamp 1626065694
transform 1 0 119000 0 1 25845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_585
timestamp 1626065694
transform 1 0 116008 0 1 24621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_584
timestamp 1626065694
transform 1 0 116008 0 1 24893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_583
timestamp 1626065694
transform 1 0 117640 0 1 24893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_582
timestamp 1626065694
transform 1 0 117640 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_581
timestamp 1626065694
transform 1 0 117640 0 1 25709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_580
timestamp 1626065694
transform 1 0 115600 0 1 25709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_579
timestamp 1626065694
transform 1 0 115600 0 1 25437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_578
timestamp 1626065694
transform 1 0 116008 0 1 25709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_577
timestamp 1626065694
transform 1 0 115600 0 1 23805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_576
timestamp 1626065694
transform 1 0 115872 0 1 25301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_575
timestamp 1626065694
transform 1 0 115872 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_574
timestamp 1626065694
transform 1 0 117640 0 1 25845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_573
timestamp 1626065694
transform 1 0 115192 0 1 25301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_572
timestamp 1626065694
transform 1 0 115192 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_571
timestamp 1626065694
transform 1 0 116008 0 1 25437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_570
timestamp 1626065694
transform 1 0 115464 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_569
timestamp 1626065694
transform 1 0 115464 0 1 25301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_568
timestamp 1626065694
transform 1 0 115464 0 1 24893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_567
timestamp 1626065694
transform 1 0 118184 0 1 25845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_566
timestamp 1626065694
transform 1 0 115872 0 1 24485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_565
timestamp 1626065694
transform 1 0 115872 0 1 24213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_564
timestamp 1626065694
transform 1 0 115464 0 1 24621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_563
timestamp 1626065694
transform 1 0 118184 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_562
timestamp 1626065694
transform 1 0 118184 0 1 25709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_561
timestamp 1626065694
transform 1 0 118184 0 1 24893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_560
timestamp 1626065694
transform 1 0 116008 0 1 25845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_559
timestamp 1626065694
transform 1 0 115192 0 1 24077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_558
timestamp 1626065694
transform 1 0 115192 0 1 23805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_557
timestamp 1626065694
transform 1 0 119000 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_556
timestamp 1626065694
transform 1 0 119000 0 1 25709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_555
timestamp 1626065694
transform 1 0 114240 0 1 23669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_554
timestamp 1626065694
transform 1 0 114648 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_553
timestamp 1626065694
transform 1 0 114240 0 1 23805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_552
timestamp 1626065694
transform 1 0 114240 0 1 24077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_551
timestamp 1626065694
transform 1 0 114784 0 1 25437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_550
timestamp 1626065694
transform 1 0 114648 0 1 25301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_549
timestamp 1626065694
transform 1 0 114648 0 1 24893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_548
timestamp 1626065694
transform 1 0 114784 0 1 25709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_547
timestamp 1626065694
transform 1 0 114648 0 1 24621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_546
timestamp 1626065694
transform 1 0 114240 0 1 24621
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_545
timestamp 1626065694
transform 1 0 114784 0 1 24213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_544
timestamp 1626065694
transform 1 0 114784 0 1 23669
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_543
timestamp 1626065694
transform 1 0 114784 0 1 23805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_542
timestamp 1626065694
transform 1 0 114784 0 1 24485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_541
timestamp 1626065694
transform 1 0 114648 0 1 25845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_540
timestamp 1626065694
transform 1 0 114240 0 1 25845
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_539
timestamp 1626065694
transform 1 0 114784 0 1 24077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_538
timestamp 1626065694
transform 1 0 114240 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_537
timestamp 1626065694
transform 1 0 114240 0 1 25709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_536
timestamp 1626065694
transform 1 0 114240 0 1 25437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_535
timestamp 1626065694
transform 1 0 114376 0 1 24485
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_534
timestamp 1626065694
transform 1 0 114376 0 1 24213
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_533
timestamp 1626065694
transform 1 0 114240 0 1 25301
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_532
timestamp 1626065694
transform 1 0 114240 0 1 24893
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_531
timestamp 1626065694
transform 1 0 114648 0 1 21357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_530
timestamp 1626065694
transform 1 0 114648 0 1 21085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_529
timestamp 1626065694
transform 1 0 114648 0 1 21493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_528
timestamp 1626065694
transform 1 0 114784 0 1 23397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_527
timestamp 1626065694
transform 1 0 114240 0 1 21765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_526
timestamp 1626065694
transform 1 0 114240 0 1 21493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_525
timestamp 1626065694
transform 1 0 114240 0 1 23397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_524
timestamp 1626065694
transform 1 0 114376 0 1 22989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_523
timestamp 1626065694
transform 1 0 114376 0 1 23261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_522
timestamp 1626065694
transform 1 0 114240 0 1 21357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_521
timestamp 1626065694
transform 1 0 114784 0 1 23261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_520
timestamp 1626065694
transform 1 0 114784 0 1 22989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_519
timestamp 1626065694
transform 1 0 114648 0 1 21765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_518
timestamp 1626065694
transform 1 0 114240 0 1 21085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_517
timestamp 1626065694
transform 1 0 118592 0 1 23261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_516
timestamp 1626065694
transform 1 0 118456 0 1 21221
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_515
timestamp 1626065694
transform 1 0 115872 0 1 21085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_514
timestamp 1626065694
transform 1 0 118592 0 1 22717
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_513
timestamp 1626065694
transform 1 0 115872 0 1 21357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_512
timestamp 1626065694
transform 1 0 118048 0 1 22717
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_511
timestamp 1626065694
transform 1 0 118048 0 1 23261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_510
timestamp 1626065694
transform 1 0 118320 0 1 22717
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_509
timestamp 1626065694
transform 1 0 118320 0 1 22989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_508
timestamp 1626065694
transform 1 0 118864 0 1 22989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_507
timestamp 1626065694
transform 1 0 118864 0 1 22717
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_506
timestamp 1626065694
transform 1 0 118456 0 1 22445
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_505
timestamp 1626065694
transform 1 0 117640 0 1 23261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_504
timestamp 1626065694
transform 1 0 116008 0 1 22717
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_503
timestamp 1626065694
transform 1 0 118184 0 1 23397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_502
timestamp 1626065694
transform 1 0 118320 0 1 21085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_501
timestamp 1626065694
transform 1 0 118320 0 1 22173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_500
timestamp 1626065694
transform 1 0 118864 0 1 22173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_499
timestamp 1626065694
transform 1 0 118864 0 1 22445
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_498
timestamp 1626065694
transform 1 0 116008 0 1 22989
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_497
timestamp 1626065694
transform 1 0 115600 0 1 21493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_496
timestamp 1626065694
transform 1 0 115600 0 1 21357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_495
timestamp 1626065694
transform 1 0 119000 0 1 23261
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_494
timestamp 1626065694
transform 1 0 119000 0 1 22717
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_493
timestamp 1626065694
transform 1 0 116008 0 1 21765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_492
timestamp 1626065694
transform 1 0 116008 0 1 21493
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_491
timestamp 1626065694
transform 1 0 115872 0 1 22309
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_490
timestamp 1626065694
transform 1 0 115872 0 1 22581
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_489
timestamp 1626065694
transform 1 0 115872 0 1 22173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_488
timestamp 1626065694
transform 1 0 115872 0 1 21901
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_487
timestamp 1626065694
transform 1 0 118048 0 1 21357
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_486
timestamp 1626065694
transform 1 0 118048 0 1 21085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_485
timestamp 1626065694
transform 1 0 115600 0 1 21085
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_484
timestamp 1626065694
transform 1 0 115600 0 1 21765
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_483
timestamp 1626065694
transform 1 0 117640 0 1 23397
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_482
timestamp 1626065694
transform 1 0 117640 0 1 22717
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_481
timestamp 1626065694
transform 1 0 135320 0 1 30469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_480
timestamp 1626065694
transform 1 0 135320 0 1 28973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_479
timestamp 1626065694
transform 1 0 135320 0 1 27205
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_478
timestamp 1626065694
transform 1 0 120768 0 1 25709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_477
timestamp 1626065694
transform 1 0 120768 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_476
timestamp 1626065694
transform 1 0 119408 0 1 25709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_475
timestamp 1626065694
transform 1 0 119408 0 1 25029
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_474
timestamp 1626065694
transform 1 0 135320 0 1 22173
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_473
timestamp 1626065694
transform 1 0 135320 0 1 23805
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_472
timestamp 1626065694
transform 1 0 135320 0 1 25437
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_471
timestamp 1626065694
transform 1 0 94520 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_470
timestamp 1626065694
transform 1 0 94520 0 1 19317
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_469
timestamp 1626065694
transform 1 0 95608 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_468
timestamp 1626065694
transform 1 0 95608 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_467
timestamp 1626065694
transform 1 0 96152 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_466
timestamp 1626065694
transform 1 0 96152 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_465
timestamp 1626065694
transform 1 0 93976 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_464
timestamp 1626065694
transform 1 0 96832 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_463
timestamp 1626065694
transform 1 0 96560 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_462
timestamp 1626065694
transform 1 0 96832 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_461
timestamp 1626065694
transform 1 0 98872 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_460
timestamp 1626065694
transform 1 0 101592 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_459
timestamp 1626065694
transform 1 0 98192 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_458
timestamp 1626065694
transform 1 0 98192 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_457
timestamp 1626065694
transform 1 0 98600 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_456
timestamp 1626065694
transform 1 0 98600 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_455
timestamp 1626065694
transform 1 0 99824 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_454
timestamp 1626065694
transform 1 0 99824 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_453
timestamp 1626065694
transform 1 0 101184 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_452
timestamp 1626065694
transform 1 0 101184 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_451
timestamp 1626065694
transform 1 0 101864 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_450
timestamp 1626065694
transform 1 0 101864 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_449
timestamp 1626065694
transform 1 0 89080 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_448
timestamp 1626065694
transform 1 0 91392 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_447
timestamp 1626065694
transform 1 0 86360 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_446
timestamp 1626065694
transform 1 0 86088 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_445
timestamp 1626065694
transform 1 0 86088 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_444
timestamp 1626065694
transform 1 0 86904 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_443
timestamp 1626065694
transform 1 0 86904 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_442
timestamp 1626065694
transform 1 0 87312 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_441
timestamp 1626065694
transform 1 0 87312 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_440
timestamp 1626065694
transform 1 0 88128 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_439
timestamp 1626065694
transform 1 0 88128 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_438
timestamp 1626065694
transform 1 0 88264 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_437
timestamp 1626065694
transform 1 0 88264 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_436
timestamp 1626065694
transform 1 0 89352 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_435
timestamp 1626065694
transform 1 0 89352 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_434
timestamp 1626065694
transform 1 0 89896 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_433
timestamp 1626065694
transform 1 0 89896 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_432
timestamp 1626065694
transform 1 0 90712 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_431
timestamp 1626065694
transform 1 0 90712 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_430
timestamp 1626065694
transform 1 0 91800 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_429
timestamp 1626065694
transform 1 0 91800 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_428
timestamp 1626065694
transform 1 0 92344 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_427
timestamp 1626065694
transform 1 0 92344 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_426
timestamp 1626065694
transform 1 0 93432 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_425
timestamp 1626065694
transform 1 0 93432 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_424
timestamp 1626065694
transform 1 0 89080 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_423
timestamp 1626065694
transform 1 0 86496 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_422
timestamp 1626065694
transform 1 0 91256 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_421
timestamp 1626065694
transform 1 0 85952 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_420
timestamp 1626065694
transform 1 0 88536 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_419
timestamp 1626065694
transform 1 0 90984 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_418
timestamp 1626065694
transform 1 0 93432 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_417
timestamp 1626065694
transform 1 0 86088 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_416
timestamp 1626065694
transform 1 0 86088 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_415
timestamp 1626065694
transform 1 0 91256 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_414
timestamp 1626065694
transform 1 0 91256 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_413
timestamp 1626065694
transform 1 0 86224 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_412
timestamp 1626065694
transform 1 0 86224 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_411
timestamp 1626065694
transform 1 0 86360 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_410
timestamp 1626065694
transform 1 0 86360 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_409
timestamp 1626065694
transform 1 0 86224 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_408
timestamp 1626065694
transform 1 0 86224 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_407
timestamp 1626065694
transform 1 0 91256 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_406
timestamp 1626065694
transform 1 0 91528 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_405
timestamp 1626065694
transform 1 0 91528 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_404
timestamp 1626065694
transform 1 0 91392 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_403
timestamp 1626065694
transform 1 0 86496 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_402
timestamp 1626065694
transform 1 0 93704 0 1 11429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_401
timestamp 1626065694
transform 1 0 93704 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_400
timestamp 1626065694
transform 1 0 86496 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_399
timestamp 1626065694
transform 1 0 88808 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_398
timestamp 1626065694
transform 1 0 88808 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_397
timestamp 1626065694
transform 1 0 88808 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_396
timestamp 1626065694
transform 1 0 88808 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_395
timestamp 1626065694
transform 1 0 88672 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_394
timestamp 1626065694
transform 1 0 88672 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_393
timestamp 1626065694
transform 1 0 86496 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_392
timestamp 1626065694
transform 1 0 86496 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_391
timestamp 1626065694
transform 1 0 93568 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_390
timestamp 1626065694
transform 1 0 86360 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_389
timestamp 1626065694
transform 1 0 93568 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_388
timestamp 1626065694
transform 1 0 86496 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_387
timestamp 1626065694
transform 1 0 91120 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_386
timestamp 1626065694
transform 1 0 91120 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_385
timestamp 1626065694
transform 1 0 91392 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_384
timestamp 1626065694
transform 1 0 91392 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_383
timestamp 1626065694
transform 1 0 91256 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_382
timestamp 1626065694
transform 1 0 91256 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_381
timestamp 1626065694
transform 1 0 88944 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_380
timestamp 1626065694
transform 1 0 88944 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_379
timestamp 1626065694
transform 1 0 88944 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_378
timestamp 1626065694
transform 1 0 88944 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_377
timestamp 1626065694
transform 1 0 88944 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_376
timestamp 1626065694
transform 1 0 88944 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_375
timestamp 1626065694
transform 1 0 96424 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_374
timestamp 1626065694
transform 1 0 96560 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_373
timestamp 1626065694
transform 1 0 93840 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_372
timestamp 1626065694
transform 1 0 96288 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_371
timestamp 1626065694
transform 1 0 99008 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_370
timestamp 1626065694
transform 1 0 99008 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_369
timestamp 1626065694
transform 1 0 95880 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_368
timestamp 1626065694
transform 1 0 98464 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_367
timestamp 1626065694
transform 1 0 100912 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_366
timestamp 1626065694
transform 1 0 99008 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_365
timestamp 1626065694
transform 1 0 99008 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_364
timestamp 1626065694
transform 1 0 99008 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_363
timestamp 1626065694
transform 1 0 99008 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_362
timestamp 1626065694
transform 1 0 98872 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_361
timestamp 1626065694
transform 1 0 93840 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_360
timestamp 1626065694
transform 1 0 101456 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_359
timestamp 1626065694
transform 1 0 101456 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_358
timestamp 1626065694
transform 1 0 101456 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_357
timestamp 1626065694
transform 1 0 101456 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_356
timestamp 1626065694
transform 1 0 101456 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_355
timestamp 1626065694
transform 1 0 101456 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_354
timestamp 1626065694
transform 1 0 101592 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_353
timestamp 1626065694
transform 1 0 93840 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_352
timestamp 1626065694
transform 1 0 96288 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_351
timestamp 1626065694
transform 1 0 93840 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_350
timestamp 1626065694
transform 1 0 96152 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_349
timestamp 1626065694
transform 1 0 93976 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_348
timestamp 1626065694
transform 1 0 98736 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_347
timestamp 1626065694
transform 1 0 98736 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_346
timestamp 1626065694
transform 1 0 98872 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_345
timestamp 1626065694
transform 1 0 98872 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_344
timestamp 1626065694
transform 1 0 98872 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_343
timestamp 1626065694
transform 1 0 98872 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_342
timestamp 1626065694
transform 1 0 93976 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_341
timestamp 1626065694
transform 1 0 96288 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_340
timestamp 1626065694
transform 1 0 93976 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_339
timestamp 1626065694
transform 1 0 93976 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_338
timestamp 1626065694
transform 1 0 101184 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_337
timestamp 1626065694
transform 1 0 101184 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_336
timestamp 1626065694
transform 1 0 101320 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_335
timestamp 1626065694
transform 1 0 101320 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_334
timestamp 1626065694
transform 1 0 101320 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_333
timestamp 1626065694
transform 1 0 101320 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_332
timestamp 1626065694
transform 1 0 93840 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_331
timestamp 1626065694
transform 1 0 96288 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_330
timestamp 1626065694
transform 1 0 96016 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_329
timestamp 1626065694
transform 1 0 96016 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_328
timestamp 1626065694
transform 1 0 96424 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_327
timestamp 1626065694
transform 1 0 96424 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_326
timestamp 1626065694
transform 1 0 96152 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_325
timestamp 1626065694
transform 1 0 96424 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_324
timestamp 1626065694
transform 1 0 81600 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_323
timestamp 1626065694
transform 1 0 77384 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_322
timestamp 1626065694
transform 1 0 77384 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_321
timestamp 1626065694
transform 1 0 78064 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_320
timestamp 1626065694
transform 1 0 78064 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_319
timestamp 1626065694
transform 1 0 79696 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_318
timestamp 1626065694
transform 1 0 79696 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_317
timestamp 1626065694
transform 1 0 80648 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_316
timestamp 1626065694
transform 1 0 80648 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_315
timestamp 1626065694
transform 1 0 81192 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_314
timestamp 1626065694
transform 1 0 81192 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_313
timestamp 1626065694
transform 1 0 81872 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_312
timestamp 1626065694
transform 1 0 81872 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_311
timestamp 1626065694
transform 1 0 83640 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_310
timestamp 1626065694
transform 1 0 83640 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_309
timestamp 1626065694
transform 1 0 83912 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_308
timestamp 1626065694
transform 1 0 84320 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_307
timestamp 1626065694
transform 1 0 84320 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_306
timestamp 1626065694
transform 1 0 84864 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_305
timestamp 1626065694
transform 1 0 84864 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_304
timestamp 1626065694
transform 1 0 78880 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_303
timestamp 1626065694
transform 1 0 69360 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_302
timestamp 1626065694
transform 1 0 69360 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_301
timestamp 1626065694
transform 1 0 70992 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_300
timestamp 1626065694
transform 1 0 70992 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_299
timestamp 1626065694
transform 1 0 71944 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_298
timestamp 1626065694
transform 1 0 71944 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_297
timestamp 1626065694
transform 1 0 72352 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_296
timestamp 1626065694
transform 1 0 72352 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_295
timestamp 1626065694
transform 1 0 73168 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_294
timestamp 1626065694
transform 1 0 73168 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_293
timestamp 1626065694
transform 1 0 74936 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_292
timestamp 1626065694
transform 1 0 74936 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_291
timestamp 1626065694
transform 1 0 75616 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_290
timestamp 1626065694
transform 1 0 75616 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_289
timestamp 1626065694
transform 1 0 76160 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_288
timestamp 1626065694
transform 1 0 76160 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_287
timestamp 1626065694
transform 1 0 68680 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_286
timestamp 1626065694
transform 1 0 74120 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_285
timestamp 1626065694
transform 1 0 76432 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_284
timestamp 1626065694
transform 1 0 68680 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_283
timestamp 1626065694
transform 1 0 69088 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_282
timestamp 1626065694
transform 1 0 71400 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_281
timestamp 1626065694
transform 1 0 76432 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_280
timestamp 1626065694
transform 1 0 76296 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_279
timestamp 1626065694
transform 1 0 76296 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_278
timestamp 1626065694
transform 1 0 71264 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_277
timestamp 1626065694
transform 1 0 68680 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_276
timestamp 1626065694
transform 1 0 68816 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_275
timestamp 1626065694
transform 1 0 68816 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_274
timestamp 1626065694
transform 1 0 76160 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_273
timestamp 1626065694
transform 1 0 68816 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_272
timestamp 1626065694
transform 1 0 68816 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_271
timestamp 1626065694
transform 1 0 73712 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_270
timestamp 1626065694
transform 1 0 73712 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_269
timestamp 1626065694
transform 1 0 73848 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_268
timestamp 1626065694
transform 1 0 73848 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_267
timestamp 1626065694
transform 1 0 73848 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_266
timestamp 1626065694
transform 1 0 73848 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_265
timestamp 1626065694
transform 1 0 76024 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_264
timestamp 1626065694
transform 1 0 76024 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_263
timestamp 1626065694
transform 1 0 76160 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_262
timestamp 1626065694
transform 1 0 68680 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_261
timestamp 1626065694
transform 1 0 71264 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_260
timestamp 1626065694
transform 1 0 71264 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_259
timestamp 1626065694
transform 1 0 71400 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_258
timestamp 1626065694
transform 1 0 76296 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_257
timestamp 1626065694
transform 1 0 76296 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_256
timestamp 1626065694
transform 1 0 76568 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_255
timestamp 1626065694
transform 1 0 76568 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_254
timestamp 1626065694
transform 1 0 73984 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_253
timestamp 1626065694
transform 1 0 74120 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_252
timestamp 1626065694
transform 1 0 71400 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_251
timestamp 1626065694
transform 1 0 76432 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_250
timestamp 1626065694
transform 1 0 71264 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_249
timestamp 1626065694
transform 1 0 73984 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_248
timestamp 1626065694
transform 1 0 76296 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_247
timestamp 1626065694
transform 1 0 73984 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_246
timestamp 1626065694
transform 1 0 70992 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_245
timestamp 1626065694
transform 1 0 68544 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_244
timestamp 1626065694
transform 1 0 68544 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_243
timestamp 1626065694
transform 1 0 68816 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_242
timestamp 1626065694
transform 1 0 68816 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_241
timestamp 1626065694
transform 1 0 68952 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_240
timestamp 1626065694
transform 1 0 68952 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_239
timestamp 1626065694
transform 1 0 69088 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_238
timestamp 1626065694
transform 1 0 76296 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_237
timestamp 1626065694
transform 1 0 71536 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_236
timestamp 1626065694
transform 1 0 71536 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_235
timestamp 1626065694
transform 1 0 71536 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_234
timestamp 1626065694
transform 1 0 71536 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_233
timestamp 1626065694
transform 1 0 73440 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_232
timestamp 1626065694
transform 1 0 71536 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_231
timestamp 1626065694
transform 1 0 71536 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_230
timestamp 1626065694
transform 1 0 71400 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_229
timestamp 1626065694
transform 1 0 76432 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_228
timestamp 1626065694
transform 1 0 75888 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_227
timestamp 1626065694
transform 1 0 73304 0 1 11429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_226
timestamp 1626065694
transform 1 0 73304 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_225
timestamp 1626065694
transform 1 0 73984 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_224
timestamp 1626065694
transform 1 0 79016 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_223
timestamp 1626065694
transform 1 0 79016 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_222
timestamp 1626065694
transform 1 0 81192 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_221
timestamp 1626065694
transform 1 0 81192 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_220
timestamp 1626065694
transform 1 0 81328 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_219
timestamp 1626065694
transform 1 0 81328 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_218
timestamp 1626065694
transform 1 0 81328 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_217
timestamp 1626065694
transform 1 0 81328 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_216
timestamp 1626065694
transform 1 0 81464 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_215
timestamp 1626065694
transform 1 0 81600 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_214
timestamp 1626065694
transform 1 0 78472 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_213
timestamp 1626065694
transform 1 0 79016 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_212
timestamp 1626065694
transform 1 0 79016 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_211
timestamp 1626065694
transform 1 0 78880 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_210
timestamp 1626065694
transform 1 0 84048 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_209
timestamp 1626065694
transform 1 0 83776 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_208
timestamp 1626065694
transform 1 0 81056 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_207
timestamp 1626065694
transform 1 0 81056 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_206
timestamp 1626065694
transform 1 0 81464 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_205
timestamp 1626065694
transform 1 0 81464 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_204
timestamp 1626065694
transform 1 0 83776 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_203
timestamp 1626065694
transform 1 0 83912 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_202
timestamp 1626065694
transform 1 0 83912 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_201
timestamp 1626065694
transform 1 0 83640 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_200
timestamp 1626065694
transform 1 0 83640 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_199
timestamp 1626065694
transform 1 0 84048 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_198
timestamp 1626065694
transform 1 0 83776 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_197
timestamp 1626065694
transform 1 0 83776 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_196
timestamp 1626065694
transform 1 0 78744 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_195
timestamp 1626065694
transform 1 0 78744 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_194
timestamp 1626065694
transform 1 0 78880 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_193
timestamp 1626065694
transform 1 0 78880 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_192
timestamp 1626065694
transform 1 0 78880 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_191
timestamp 1626065694
transform 1 0 78880 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_190
timestamp 1626065694
transform 1 0 84048 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_189
timestamp 1626065694
transform 1 0 84048 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_188
timestamp 1626065694
transform 1 0 80920 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_187
timestamp 1626065694
transform 1 0 83912 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_186
timestamp 1626065694
transform 1 0 83504 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_185
timestamp 1626065694
transform 1 0 81464 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_184
timestamp 1626065694
transform 1 0 78608 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_183
timestamp 1626065694
transform 1 0 78608 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_182
timestamp 1626065694
transform 1 0 69224 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_181
timestamp 1626065694
transform 1 0 69224 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_180
timestamp 1626065694
transform 1 0 70856 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_179
timestamp 1626065694
transform 1 0 70856 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_178
timestamp 1626065694
transform 1 0 72760 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_177
timestamp 1626065694
transform 1 0 72760 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_176
timestamp 1626065694
transform 1 0 74256 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_175
timestamp 1626065694
transform 1 0 74256 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_174
timestamp 1626065694
transform 1 0 76160 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_173
timestamp 1626065694
transform 1 0 76160 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_172
timestamp 1626065694
transform 1 0 77656 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_171
timestamp 1626065694
transform 1 0 77656 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_170
timestamp 1626065694
transform 1 0 84320 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_169
timestamp 1626065694
transform 1 0 84320 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_168
timestamp 1626065694
transform 1 0 79288 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_167
timestamp 1626065694
transform 1 0 79288 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_166
timestamp 1626065694
transform 1 0 82824 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_165
timestamp 1626065694
transform 1 0 82824 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_164
timestamp 1626065694
transform 1 0 81056 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_163
timestamp 1626065694
transform 1 0 81056 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_162
timestamp 1626065694
transform 1 0 86224 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_161
timestamp 1626065694
transform 1 0 86224 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_160
timestamp 1626065694
transform 1 0 87720 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_159
timestamp 1626065694
transform 1 0 87720 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_158
timestamp 1626065694
transform 1 0 89352 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_157
timestamp 1626065694
transform 1 0 89352 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_156
timestamp 1626065694
transform 1 0 91256 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_155
timestamp 1626065694
transform 1 0 91256 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_154
timestamp 1626065694
transform 1 0 92752 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_153
timestamp 1626065694
transform 1 0 92752 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_152
timestamp 1626065694
transform 1 0 94384 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_151
timestamp 1626065694
transform 1 0 96152 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_150
timestamp 1626065694
transform 1 0 94384 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_149
timestamp 1626065694
transform 1 0 96152 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_148
timestamp 1626065694
transform 1 0 99552 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_147
timestamp 1626065694
transform 1 0 99552 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_146
timestamp 1626065694
transform 1 0 101320 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_145
timestamp 1626065694
transform 1 0 101320 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_144
timestamp 1626065694
transform 1 0 97784 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_143
timestamp 1626065694
transform 1 0 97784 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_142
timestamp 1626065694
transform 1 0 108256 0 1 10613
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_141
timestamp 1626065694
transform 1 0 135320 0 1 17141
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_140
timestamp 1626065694
transform 1 0 135320 0 1 20541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_139
timestamp 1626065694
transform 1 0 135320 0 1 18909
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_138
timestamp 1626065694
transform 1 0 119952 0 1 20133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_137
timestamp 1626065694
transform 1 0 119952 0 1 18501
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_136
timestamp 1626065694
transform 1 0 122944 0 1 18365
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_135
timestamp 1626065694
transform 1 0 122808 0 1 20133
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_134
timestamp 1626065694
transform 1 0 122808 0 1 19861
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_133
timestamp 1626065694
transform 1 0 122808 0 1 16869
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_132
timestamp 1626065694
transform 1 0 122808 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_131
timestamp 1626065694
transform 1 0 122808 0 1 19725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_130
timestamp 1626065694
transform 1 0 122944 0 1 12653
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_129
timestamp 1626065694
transform 1 0 123352 0 1 10749
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_128
timestamp 1626065694
transform 1 0 123216 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_127
timestamp 1626065694
transform 1 0 122944 0 1 15645
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_126
timestamp 1626065694
transform 1 0 122944 0 1 12789
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_125
timestamp 1626065694
transform 1 0 122944 0 1 15509
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_124
timestamp 1626065694
transform 1 0 122808 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_123
timestamp 1626065694
transform 1 0 122808 0 1 11429
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_122
timestamp 1626065694
transform 1 0 122808 0 1 14013
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_121
timestamp 1626065694
transform 1 0 135320 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_120
timestamp 1626065694
transform 1 0 135320 0 1 15373
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_119
timestamp 1626065694
transform 1 0 135320 0 1 13877
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_118
timestamp 1626065694
transform 1 0 103768 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_117
timestamp 1626065694
transform 1 0 107168 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_116
timestamp 1626065694
transform 1 0 107304 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_115
timestamp 1626065694
transform 1 0 103904 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_114
timestamp 1626065694
transform 1 0 103904 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_113
timestamp 1626065694
transform 1 0 107304 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_112
timestamp 1626065694
transform 1 0 104040 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_111
timestamp 1626065694
transform 1 0 114240 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_110
timestamp 1626065694
transform 1 0 104040 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_109
timestamp 1626065694
transform 1 0 108392 0 1 11293
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_108
timestamp 1626065694
transform 1 0 114240 0 1 20541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_107
timestamp 1626065694
transform 1 0 103088 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_106
timestamp 1626065694
transform 1 0 108528 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_105
timestamp 1626065694
transform 1 0 108528 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_104
timestamp 1626065694
transform 1 0 106080 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_103
timestamp 1626065694
transform 1 0 106080 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_102
timestamp 1626065694
transform 1 0 106488 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_101
timestamp 1626065694
transform 1 0 106488 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_100
timestamp 1626065694
transform 1 0 106488 0 1 13197
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_99
timestamp 1626065694
transform 1 0 106488 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_98
timestamp 1626065694
transform 1 0 114240 0 1 20677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_97
timestamp 1626065694
transform 1 0 103088 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_96
timestamp 1626065694
transform 1 0 115056 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_95
timestamp 1626065694
transform 1 0 117640 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_94
timestamp 1626065694
transform 1 0 115056 0 1 20541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_93
timestamp 1626065694
transform 1 0 103632 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_92
timestamp 1626065694
transform 1 0 103632 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_91
timestamp 1626065694
transform 1 0 103632 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_90
timestamp 1626065694
transform 1 0 103632 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_89
timestamp 1626065694
transform 1 0 103768 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_88
timestamp 1626065694
transform 1 0 103768 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_87
timestamp 1626065694
transform 1 0 106352 0 1 15101
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_86
timestamp 1626065694
transform 1 0 115464 0 1 20541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_85
timestamp 1626065694
transform 1 0 104312 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_84
timestamp 1626065694
transform 1 0 104312 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_83
timestamp 1626065694
transform 1 0 114648 0 1 20677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_82
timestamp 1626065694
transform 1 0 106352 0 1 17005
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_81
timestamp 1626065694
transform 1 0 103496 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_80
timestamp 1626065694
transform 1 0 104856 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_79
timestamp 1626065694
transform 1 0 104856 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_78
timestamp 1626065694
transform 1 0 103496 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_77
timestamp 1626065694
transform 1 0 109616 0 1 19997
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_76
timestamp 1626065694
transform 1 0 105536 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_75
timestamp 1626065694
transform 1 0 105536 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_74
timestamp 1626065694
transform 1 0 105808 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_73
timestamp 1626065694
transform 1 0 105808 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_72
timestamp 1626065694
transform 1 0 109616 0 1 19725
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_71
timestamp 1626065694
transform 1 0 115464 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_70
timestamp 1626065694
transform 1 0 115328 0 1 20677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_69
timestamp 1626065694
transform 1 0 118184 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_68
timestamp 1626065694
transform 1 0 103360 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_67
timestamp 1626065694
transform 1 0 105944 0 1 13061
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_66
timestamp 1626065694
transform 1 0 119000 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_65
timestamp 1626065694
transform 1 0 102408 0 1 18773
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_64
timestamp 1626065694
transform 1 0 106216 0 1 11837
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_63
timestamp 1626065694
transform 1 0 106216 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_62
timestamp 1626065694
transform 1 0 106352 0 1 11973
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_61
timestamp 1626065694
transform 1 0 106352 0 1 13469
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_60
timestamp 1626065694
transform 1 0 108256 0 1 11021
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_59
timestamp 1626065694
transform 1 0 102408 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_58
timestamp 1626065694
transform 1 0 106352 0 1 14285
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_57
timestamp 1626065694
transform 1 0 106352 0 1 13605
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_56
timestamp 1626065694
transform 1 0 115192 0 1 20677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_55
timestamp 1626065694
transform 1 0 114648 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_54
timestamp 1626065694
transform 1 0 114648 0 1 20541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_53
timestamp 1626065694
transform 1 0 118592 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_52
timestamp 1626065694
transform 1 0 107168 0 1 19181
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_51
timestamp 1626065694
transform 1 0 116008 0 1 20677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_50
timestamp 1626065694
transform 1 0 116008 0 1 20541
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_49
timestamp 1626065694
transform 1 0 116008 0 1 20269
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_48
timestamp 1626065694
transform 1 0 103768 0 1 12245
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_47
timestamp 1626065694
transform 1 0 103768 0 1 11701
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_46
timestamp 1626065694
transform 1 0 103768 0 1 12517
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_45
timestamp 1626065694
transform 1 0 108392 0 1 9525
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_44
timestamp 1626065694
transform 1 0 104584 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_43
timestamp 1626065694
transform 1 0 104584 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_42
timestamp 1626065694
transform 1 0 102816 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_41
timestamp 1626065694
transform 1 0 107848 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_40
timestamp 1626065694
transform 1 0 107848 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_39
timestamp 1626065694
transform 1 0 109752 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_38
timestamp 1626065694
transform 1 0 109752 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_37
timestamp 1626065694
transform 1 0 106216 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_36
timestamp 1626065694
transform 1 0 106216 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_35
timestamp 1626065694
transform 1 0 102816 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_34
timestamp 1626065694
transform 1 0 113016 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_33
timestamp 1626065694
transform 1 0 113016 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_32
timestamp 1626065694
transform 1 0 114784 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_31
timestamp 1626065694
transform 1 0 114784 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_30
timestamp 1626065694
transform 1 0 118048 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_29
timestamp 1626065694
transform 1 0 118048 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_28
timestamp 1626065694
transform 1 0 116280 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_27
timestamp 1626065694
transform 1 0 116280 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_26
timestamp 1626065694
transform 1 0 111248 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_25
timestamp 1626065694
transform 1 0 111248 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_24
timestamp 1626065694
transform 1 0 135320 0 1 10341
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_23
timestamp 1626065694
transform 1 0 135320 0 1 8709
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_22
timestamp 1626065694
transform 1 0 135320 0 1 7077
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_21
timestamp 1626065694
transform 1 0 122944 0 1 9933
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_20
timestamp 1626065694
transform 1 0 119816 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_19
timestamp 1626065694
transform 1 0 121312 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_18
timestamp 1626065694
transform 1 0 121312 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_17
timestamp 1626065694
transform 1 0 123080 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_16
timestamp 1626065694
transform 1 0 123080 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_15
timestamp 1626065694
transform 1 0 124712 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_14
timestamp 1626065694
transform 1 0 124712 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_13
timestamp 1626065694
transform 1 0 126344 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_12
timestamp 1626065694
transform 1 0 126344 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_11
timestamp 1626065694
transform 1 0 119816 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_10
timestamp 1626065694
transform 1 0 135320 0 1 5309
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_9
timestamp 1626065694
transform 1 0 135320 0 1 3677
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_8
timestamp 1626065694
transform 1 0 127976 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_7
timestamp 1626065694
transform 1 0 127976 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_6
timestamp 1626065694
transform 1 0 129744 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_5
timestamp 1626065694
transform 1 0 129744 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_4
timestamp 1626065694
transform 1 0 131512 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_3
timestamp 1626065694
transform 1 0 131512 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_2
timestamp 1626065694
transform 1 0 135320 0 1 2045
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_1
timestamp 1626065694
transform 1 0 133144 0 1 1637
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_33  sky130_sram_2kbyte_1rw1r_32x512_8_contact_33_0
timestamp 1626065694
transform 1 0 133144 0 1 1229
box 0 0 76 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1259
timestamp 1626065694
transform 1 0 68325 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1258
timestamp 1626065694
transform 1 0 68325 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1257
timestamp 1626065694
transform 1 0 1797 0 1 41667
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1256
timestamp 1626065694
transform 1 0 134847 0 1 41667
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1255
timestamp 1626065694
transform 1 0 102261 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1254
timestamp 1626065694
transform 1 0 119397 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1253
timestamp 1626065694
transform 1 0 134847 0 1 72579
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1252
timestamp 1626065694
transform 1 0 127797 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1251
timestamp 1626065694
transform 1 0 132165 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1250
timestamp 1626065694
transform 1 0 132501 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1249
timestamp 1626065694
transform 1 0 132837 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1248
timestamp 1626065694
transform 1 0 133173 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1247
timestamp 1626065694
transform 1 0 133509 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1246
timestamp 1626065694
transform 1 0 133845 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1245
timestamp 1626065694
transform 1 0 134181 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1244
timestamp 1626065694
transform 1 0 134847 0 1 80643
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1243
timestamp 1626065694
transform 1 0 134847 0 1 80979
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1242
timestamp 1626065694
transform 1 0 130149 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1241
timestamp 1626065694
transform 1 0 130485 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1240
timestamp 1626065694
transform 1 0 130821 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1239
timestamp 1626065694
transform 1 0 131157 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1238
timestamp 1626065694
transform 1 0 131493 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1237
timestamp 1626065694
transform 1 0 131829 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1236
timestamp 1626065694
transform 1 0 128133 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1235
timestamp 1626065694
transform 1 0 128469 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1234
timestamp 1626065694
transform 1 0 128805 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1233
timestamp 1626065694
transform 1 0 129141 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1232
timestamp 1626065694
transform 1 0 129477 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1231
timestamp 1626065694
transform 1 0 129813 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1230
timestamp 1626065694
transform 1 0 134847 0 1 79299
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1229
timestamp 1626065694
transform 1 0 134847 0 1 79635
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1228
timestamp 1626065694
transform 1 0 134847 0 1 79971
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1227
timestamp 1626065694
transform 1 0 134847 0 1 80307
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1226
timestamp 1626065694
transform 1 0 134847 0 1 77955
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1225
timestamp 1626065694
transform 1 0 134847 0 1 78291
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1224
timestamp 1626065694
transform 1 0 134847 0 1 78627
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1223
timestamp 1626065694
transform 1 0 134847 0 1 78963
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1222
timestamp 1626065694
transform 1 0 126789 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1221
timestamp 1626065694
transform 1 0 127125 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1220
timestamp 1626065694
transform 1 0 127461 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1219
timestamp 1626065694
transform 1 0 119733 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1218
timestamp 1626065694
transform 1 0 120069 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1217
timestamp 1626065694
transform 1 0 120405 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1216
timestamp 1626065694
transform 1 0 120741 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1215
timestamp 1626065694
transform 1 0 121077 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1214
timestamp 1626065694
transform 1 0 121413 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1213
timestamp 1626065694
transform 1 0 121749 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1212
timestamp 1626065694
transform 1 0 122085 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1211
timestamp 1626065694
transform 1 0 122421 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1210
timestamp 1626065694
transform 1 0 122757 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1209
timestamp 1626065694
transform 1 0 123093 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1208
timestamp 1626065694
transform 1 0 123429 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1207
timestamp 1626065694
transform 1 0 123765 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1206
timestamp 1626065694
transform 1 0 124101 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1205
timestamp 1626065694
transform 1 0 124437 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1204
timestamp 1626065694
transform 1 0 124773 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1203
timestamp 1626065694
transform 1 0 125109 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1202
timestamp 1626065694
transform 1 0 125445 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1201
timestamp 1626065694
transform 1 0 125781 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1200
timestamp 1626065694
transform 1 0 126117 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1199
timestamp 1626065694
transform 1 0 126453 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1198
timestamp 1626065694
transform 1 0 134847 0 1 77619
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1197
timestamp 1626065694
transform 1 0 134847 0 1 72915
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1196
timestamp 1626065694
transform 1 0 134847 0 1 73251
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1195
timestamp 1626065694
transform 1 0 134847 0 1 73587
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1194
timestamp 1626065694
transform 1 0 134847 0 1 73923
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1193
timestamp 1626065694
transform 1 0 134847 0 1 74259
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1192
timestamp 1626065694
transform 1 0 134847 0 1 74595
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1191
timestamp 1626065694
transform 1 0 134847 0 1 74931
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1190
timestamp 1626065694
transform 1 0 134847 0 1 75267
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1189
timestamp 1626065694
transform 1 0 134847 0 1 75603
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1188
timestamp 1626065694
transform 1 0 134847 0 1 75939
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1187
timestamp 1626065694
transform 1 0 134847 0 1 76275
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1186
timestamp 1626065694
transform 1 0 134847 0 1 76611
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1185
timestamp 1626065694
transform 1 0 134847 0 1 76947
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1184
timestamp 1626065694
transform 1 0 134847 0 1 77283
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1183
timestamp 1626065694
transform 1 0 111333 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1182
timestamp 1626065694
transform 1 0 111669 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1181
timestamp 1626065694
transform 1 0 112005 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1180
timestamp 1626065694
transform 1 0 112341 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1179
timestamp 1626065694
transform 1 0 112677 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1178
timestamp 1626065694
transform 1 0 113013 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1177
timestamp 1626065694
transform 1 0 113349 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1176
timestamp 1626065694
transform 1 0 113685 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1175
timestamp 1626065694
transform 1 0 114021 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1174
timestamp 1626065694
transform 1 0 114357 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1173
timestamp 1626065694
transform 1 0 114693 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1172
timestamp 1626065694
transform 1 0 115029 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1171
timestamp 1626065694
transform 1 0 115365 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1170
timestamp 1626065694
transform 1 0 115701 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1169
timestamp 1626065694
transform 1 0 116037 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1168
timestamp 1626065694
transform 1 0 116373 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1167
timestamp 1626065694
transform 1 0 116709 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1166
timestamp 1626065694
transform 1 0 117045 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1165
timestamp 1626065694
transform 1 0 117381 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1164
timestamp 1626065694
transform 1 0 117717 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1163
timestamp 1626065694
transform 1 0 118053 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1162
timestamp 1626065694
transform 1 0 118389 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1161
timestamp 1626065694
transform 1 0 110997 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1160
timestamp 1626065694
transform 1 0 118725 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1159
timestamp 1626065694
transform 1 0 119061 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1158
timestamp 1626065694
transform 1 0 106629 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1157
timestamp 1626065694
transform 1 0 106965 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1156
timestamp 1626065694
transform 1 0 107301 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1155
timestamp 1626065694
transform 1 0 107637 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1154
timestamp 1626065694
transform 1 0 107973 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1153
timestamp 1626065694
transform 1 0 108309 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1152
timestamp 1626065694
transform 1 0 108645 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1151
timestamp 1626065694
transform 1 0 108981 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1150
timestamp 1626065694
transform 1 0 109317 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1149
timestamp 1626065694
transform 1 0 109653 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1148
timestamp 1626065694
transform 1 0 109989 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1147
timestamp 1626065694
transform 1 0 110325 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1146
timestamp 1626065694
transform 1 0 110661 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1145
timestamp 1626065694
transform 1 0 103269 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1144
timestamp 1626065694
transform 1 0 103605 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1143
timestamp 1626065694
transform 1 0 103941 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1142
timestamp 1626065694
transform 1 0 104277 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1141
timestamp 1626065694
transform 1 0 104613 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1140
timestamp 1626065694
transform 1 0 104949 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1139
timestamp 1626065694
transform 1 0 105285 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1138
timestamp 1626065694
transform 1 0 105621 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1137
timestamp 1626065694
transform 1 0 105957 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1136
timestamp 1626065694
transform 1 0 106293 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1135
timestamp 1626065694
transform 1 0 102597 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1134
timestamp 1626065694
transform 1 0 102933 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1133
timestamp 1626065694
transform 1 0 134847 0 1 67539
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1132
timestamp 1626065694
transform 1 0 134847 0 1 68211
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1131
timestamp 1626065694
transform 1 0 134847 0 1 68547
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1130
timestamp 1626065694
transform 1 0 134847 0 1 68883
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1129
timestamp 1626065694
transform 1 0 134847 0 1 69219
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1128
timestamp 1626065694
transform 1 0 134847 0 1 69555
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1127
timestamp 1626065694
transform 1 0 134847 0 1 69891
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1126
timestamp 1626065694
transform 1 0 134847 0 1 70227
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1125
timestamp 1626065694
transform 1 0 134847 0 1 70563
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1124
timestamp 1626065694
transform 1 0 134847 0 1 70899
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1123
timestamp 1626065694
transform 1 0 134847 0 1 71235
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1122
timestamp 1626065694
transform 1 0 134847 0 1 71571
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1121
timestamp 1626065694
transform 1 0 134847 0 1 71907
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1120
timestamp 1626065694
transform 1 0 134847 0 1 72243
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1119
timestamp 1626065694
transform 1 0 134847 0 1 67875
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1118
timestamp 1626065694
transform 1 0 134847 0 1 63843
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1117
timestamp 1626065694
transform 1 0 134847 0 1 64179
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1116
timestamp 1626065694
transform 1 0 134847 0 1 64515
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1115
timestamp 1626065694
transform 1 0 134847 0 1 64851
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1114
timestamp 1626065694
transform 1 0 134847 0 1 65187
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1113
timestamp 1626065694
transform 1 0 134847 0 1 65523
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1112
timestamp 1626065694
transform 1 0 134847 0 1 65859
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1111
timestamp 1626065694
transform 1 0 134847 0 1 66195
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1110
timestamp 1626065694
transform 1 0 134847 0 1 66531
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1109
timestamp 1626065694
transform 1 0 134847 0 1 66867
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1108
timestamp 1626065694
transform 1 0 134847 0 1 67203
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1107
timestamp 1626065694
transform 1 0 134847 0 1 62835
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1106
timestamp 1626065694
transform 1 0 134847 0 1 63171
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1105
timestamp 1626065694
transform 1 0 134847 0 1 62499
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1104
timestamp 1626065694
transform 1 0 134847 0 1 63507
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1103
timestamp 1626065694
transform 1 0 93861 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1102
timestamp 1626065694
transform 1 0 94197 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1101
timestamp 1626065694
transform 1 0 94533 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1100
timestamp 1626065694
transform 1 0 94869 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1099
timestamp 1626065694
transform 1 0 95205 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1098
timestamp 1626065694
transform 1 0 95541 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1097
timestamp 1626065694
transform 1 0 95877 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1096
timestamp 1626065694
transform 1 0 96213 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1095
timestamp 1626065694
transform 1 0 96549 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1094
timestamp 1626065694
transform 1 0 96885 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1093
timestamp 1626065694
transform 1 0 97221 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1092
timestamp 1626065694
transform 1 0 97557 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1091
timestamp 1626065694
transform 1 0 97893 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1090
timestamp 1626065694
transform 1 0 98229 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1089
timestamp 1626065694
transform 1 0 98565 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1088
timestamp 1626065694
transform 1 0 98901 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1087
timestamp 1626065694
transform 1 0 99237 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1086
timestamp 1626065694
transform 1 0 99573 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1085
timestamp 1626065694
transform 1 0 99909 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1084
timestamp 1626065694
transform 1 0 100245 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1083
timestamp 1626065694
transform 1 0 100581 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1082
timestamp 1626065694
transform 1 0 100917 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1081
timestamp 1626065694
transform 1 0 101253 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1080
timestamp 1626065694
transform 1 0 101589 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1079
timestamp 1626065694
transform 1 0 101925 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1078
timestamp 1626065694
transform 1 0 86805 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1077
timestamp 1626065694
transform 1 0 87141 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1076
timestamp 1626065694
transform 1 0 87477 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1075
timestamp 1626065694
transform 1 0 87813 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1074
timestamp 1626065694
transform 1 0 88149 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1073
timestamp 1626065694
transform 1 0 88485 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1072
timestamp 1626065694
transform 1 0 88821 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1071
timestamp 1626065694
transform 1 0 89157 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1070
timestamp 1626065694
transform 1 0 89493 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1069
timestamp 1626065694
transform 1 0 89829 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1068
timestamp 1626065694
transform 1 0 90165 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1067
timestamp 1626065694
transform 1 0 90501 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1066
timestamp 1626065694
transform 1 0 90837 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1065
timestamp 1626065694
transform 1 0 91173 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1064
timestamp 1626065694
transform 1 0 91509 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1063
timestamp 1626065694
transform 1 0 91845 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1062
timestamp 1626065694
transform 1 0 92181 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1061
timestamp 1626065694
transform 1 0 92517 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1060
timestamp 1626065694
transform 1 0 92853 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1059
timestamp 1626065694
transform 1 0 93189 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1058
timestamp 1626065694
transform 1 0 93525 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1057
timestamp 1626065694
transform 1 0 85461 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1056
timestamp 1626065694
transform 1 0 85797 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1055
timestamp 1626065694
transform 1 0 86133 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1054
timestamp 1626065694
transform 1 0 86469 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1053
timestamp 1626065694
transform 1 0 76725 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1052
timestamp 1626065694
transform 1 0 77061 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1051
timestamp 1626065694
transform 1 0 77397 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1050
timestamp 1626065694
transform 1 0 77733 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1049
timestamp 1626065694
transform 1 0 78069 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1048
timestamp 1626065694
transform 1 0 78405 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1047
timestamp 1626065694
transform 1 0 78741 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1046
timestamp 1626065694
transform 1 0 79077 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1045
timestamp 1626065694
transform 1 0 79413 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1044
timestamp 1626065694
transform 1 0 79749 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1043
timestamp 1626065694
transform 1 0 80085 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1042
timestamp 1626065694
transform 1 0 80421 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1041
timestamp 1626065694
transform 1 0 80757 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1040
timestamp 1626065694
transform 1 0 81093 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1039
timestamp 1626065694
transform 1 0 81429 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1038
timestamp 1626065694
transform 1 0 81765 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1037
timestamp 1626065694
transform 1 0 82101 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1036
timestamp 1626065694
transform 1 0 82437 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1035
timestamp 1626065694
transform 1 0 82773 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1034
timestamp 1626065694
transform 1 0 83109 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1033
timestamp 1626065694
transform 1 0 83445 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1032
timestamp 1626065694
transform 1 0 83781 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1031
timestamp 1626065694
transform 1 0 84117 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1030
timestamp 1626065694
transform 1 0 84453 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1029
timestamp 1626065694
transform 1 0 84789 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1028
timestamp 1626065694
transform 1 0 85125 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1027
timestamp 1626065694
transform 1 0 68997 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1026
timestamp 1626065694
transform 1 0 69333 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1025
timestamp 1626065694
transform 1 0 69669 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1024
timestamp 1626065694
transform 1 0 70005 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1023
timestamp 1626065694
transform 1 0 70341 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1022
timestamp 1626065694
transform 1 0 70677 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1021
timestamp 1626065694
transform 1 0 71013 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1020
timestamp 1626065694
transform 1 0 71349 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1019
timestamp 1626065694
transform 1 0 71685 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1018
timestamp 1626065694
transform 1 0 72021 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1017
timestamp 1626065694
transform 1 0 72357 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1016
timestamp 1626065694
transform 1 0 72693 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1015
timestamp 1626065694
transform 1 0 73029 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1014
timestamp 1626065694
transform 1 0 73365 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1013
timestamp 1626065694
transform 1 0 68661 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1012
timestamp 1626065694
transform 1 0 73701 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1011
timestamp 1626065694
transform 1 0 74037 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1010
timestamp 1626065694
transform 1 0 74373 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1009
timestamp 1626065694
transform 1 0 74709 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1008
timestamp 1626065694
transform 1 0 75045 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1007
timestamp 1626065694
transform 1 0 75381 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1006
timestamp 1626065694
transform 1 0 75717 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1005
timestamp 1626065694
transform 1 0 76053 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1004
timestamp 1626065694
transform 1 0 76389 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1003
timestamp 1626065694
transform 1 0 134847 0 1 57123
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1002
timestamp 1626065694
transform 1 0 134847 0 1 57459
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1001
timestamp 1626065694
transform 1 0 134847 0 1 57795
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1000
timestamp 1626065694
transform 1 0 134847 0 1 58131
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_999
timestamp 1626065694
transform 1 0 134847 0 1 58467
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_998
timestamp 1626065694
transform 1 0 134847 0 1 58803
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_997
timestamp 1626065694
transform 1 0 134847 0 1 59139
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_996
timestamp 1626065694
transform 1 0 134847 0 1 59475
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_995
timestamp 1626065694
transform 1 0 134847 0 1 59811
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_994
timestamp 1626065694
transform 1 0 134847 0 1 60147
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_993
timestamp 1626065694
transform 1 0 134847 0 1 60483
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_992
timestamp 1626065694
transform 1 0 134847 0 1 60819
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_991
timestamp 1626065694
transform 1 0 134847 0 1 61155
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_990
timestamp 1626065694
transform 1 0 134847 0 1 61491
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_989
timestamp 1626065694
transform 1 0 134847 0 1 61827
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_988
timestamp 1626065694
transform 1 0 134847 0 1 62163
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_987
timestamp 1626065694
transform 1 0 134847 0 1 52755
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_986
timestamp 1626065694
transform 1 0 134847 0 1 53091
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_985
timestamp 1626065694
transform 1 0 134847 0 1 53427
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_984
timestamp 1626065694
transform 1 0 134847 0 1 53763
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_983
timestamp 1626065694
transform 1 0 134847 0 1 54099
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_982
timestamp 1626065694
transform 1 0 134847 0 1 54435
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_981
timestamp 1626065694
transform 1 0 134847 0 1 54771
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_980
timestamp 1626065694
transform 1 0 134847 0 1 55107
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_979
timestamp 1626065694
transform 1 0 134847 0 1 55443
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_978
timestamp 1626065694
transform 1 0 134847 0 1 55779
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_977
timestamp 1626065694
transform 1 0 134847 0 1 56115
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_976
timestamp 1626065694
transform 1 0 134847 0 1 56451
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_975
timestamp 1626065694
transform 1 0 134847 0 1 52083
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_974
timestamp 1626065694
transform 1 0 134847 0 1 56787
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_973
timestamp 1626065694
transform 1 0 134847 0 1 52419
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_972
timestamp 1626065694
transform 1 0 134847 0 1 46707
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_971
timestamp 1626065694
transform 1 0 134847 0 1 50067
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_970
timestamp 1626065694
transform 1 0 134847 0 1 49059
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_969
timestamp 1626065694
transform 1 0 134847 0 1 50739
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_968
timestamp 1626065694
transform 1 0 134847 0 1 51075
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_967
timestamp 1626065694
transform 1 0 134847 0 1 51411
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_966
timestamp 1626065694
transform 1 0 134847 0 1 50403
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_965
timestamp 1626065694
transform 1 0 134847 0 1 51747
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_964
timestamp 1626065694
transform 1 0 134847 0 1 48387
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_963
timestamp 1626065694
transform 1 0 134847 0 1 49395
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_962
timestamp 1626065694
transform 1 0 134847 0 1 49731
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_961
timestamp 1626065694
transform 1 0 134847 0 1 48051
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_960
timestamp 1626065694
transform 1 0 134847 0 1 47043
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_959
timestamp 1626065694
transform 1 0 134847 0 1 47379
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_958
timestamp 1626065694
transform 1 0 134847 0 1 48723
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_957
timestamp 1626065694
transform 1 0 134847 0 1 47715
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_956
timestamp 1626065694
transform 1 0 134847 0 1 45699
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_955
timestamp 1626065694
transform 1 0 134847 0 1 46371
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_954
timestamp 1626065694
transform 1 0 134847 0 1 44355
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_953
timestamp 1626065694
transform 1 0 134847 0 1 44691
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_952
timestamp 1626065694
transform 1 0 134847 0 1 42003
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_951
timestamp 1626065694
transform 1 0 134847 0 1 45363
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_950
timestamp 1626065694
transform 1 0 134847 0 1 42339
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_949
timestamp 1626065694
transform 1 0 134847 0 1 42675
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_948
timestamp 1626065694
transform 1 0 134847 0 1 46035
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_947
timestamp 1626065694
transform 1 0 134847 0 1 45027
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_946
timestamp 1626065694
transform 1 0 134847 0 1 43011
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_945
timestamp 1626065694
transform 1 0 134847 0 1 43347
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_944
timestamp 1626065694
transform 1 0 134847 0 1 43683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_943
timestamp 1626065694
transform 1 0 134847 0 1 44019
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_942
timestamp 1626065694
transform 1 0 59925 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_941
timestamp 1626065694
transform 1 0 60261 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_940
timestamp 1626065694
transform 1 0 60597 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_939
timestamp 1626065694
transform 1 0 60933 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_938
timestamp 1626065694
transform 1 0 61269 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_937
timestamp 1626065694
transform 1 0 61605 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_936
timestamp 1626065694
transform 1 0 61941 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_935
timestamp 1626065694
transform 1 0 62277 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_934
timestamp 1626065694
transform 1 0 62613 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_933
timestamp 1626065694
transform 1 0 62949 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_932
timestamp 1626065694
transform 1 0 63285 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_931
timestamp 1626065694
transform 1 0 63621 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_930
timestamp 1626065694
transform 1 0 63957 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_929
timestamp 1626065694
transform 1 0 64293 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_928
timestamp 1626065694
transform 1 0 64629 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_927
timestamp 1626065694
transform 1 0 64965 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_926
timestamp 1626065694
transform 1 0 65301 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_925
timestamp 1626065694
transform 1 0 65637 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_924
timestamp 1626065694
transform 1 0 65973 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_923
timestamp 1626065694
transform 1 0 66309 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_922
timestamp 1626065694
transform 1 0 66645 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_921
timestamp 1626065694
transform 1 0 66981 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_920
timestamp 1626065694
transform 1 0 67317 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_919
timestamp 1626065694
transform 1 0 67653 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_918
timestamp 1626065694
transform 1 0 67989 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_917
timestamp 1626065694
transform 1 0 58917 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_916
timestamp 1626065694
transform 1 0 59253 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_915
timestamp 1626065694
transform 1 0 59589 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_914
timestamp 1626065694
transform 1 0 51861 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_913
timestamp 1626065694
transform 1 0 52197 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_912
timestamp 1626065694
transform 1 0 52533 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_911
timestamp 1626065694
transform 1 0 52869 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_910
timestamp 1626065694
transform 1 0 53205 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_909
timestamp 1626065694
transform 1 0 53541 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_908
timestamp 1626065694
transform 1 0 53877 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_907
timestamp 1626065694
transform 1 0 54213 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_906
timestamp 1626065694
transform 1 0 54549 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_905
timestamp 1626065694
transform 1 0 54885 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_904
timestamp 1626065694
transform 1 0 55221 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_903
timestamp 1626065694
transform 1 0 55557 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_902
timestamp 1626065694
transform 1 0 55893 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_901
timestamp 1626065694
transform 1 0 56229 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_900
timestamp 1626065694
transform 1 0 56565 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_899
timestamp 1626065694
transform 1 0 56901 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_898
timestamp 1626065694
transform 1 0 57237 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_897
timestamp 1626065694
transform 1 0 57573 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_896
timestamp 1626065694
transform 1 0 57909 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_895
timestamp 1626065694
transform 1 0 58245 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_894
timestamp 1626065694
transform 1 0 58581 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_893
timestamp 1626065694
transform 1 0 51525 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_892
timestamp 1626065694
transform 1 0 42789 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_891
timestamp 1626065694
transform 1 0 47157 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_890
timestamp 1626065694
transform 1 0 47493 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_889
timestamp 1626065694
transform 1 0 47829 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_888
timestamp 1626065694
transform 1 0 48165 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_887
timestamp 1626065694
transform 1 0 48501 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_886
timestamp 1626065694
transform 1 0 48837 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_885
timestamp 1626065694
transform 1 0 49173 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_884
timestamp 1626065694
transform 1 0 49509 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_883
timestamp 1626065694
transform 1 0 49845 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_882
timestamp 1626065694
transform 1 0 50181 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_881
timestamp 1626065694
transform 1 0 50517 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_880
timestamp 1626065694
transform 1 0 50853 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_879
timestamp 1626065694
transform 1 0 51189 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_878
timestamp 1626065694
transform 1 0 46821 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_877
timestamp 1626065694
transform 1 0 43125 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_876
timestamp 1626065694
transform 1 0 43461 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_875
timestamp 1626065694
transform 1 0 43797 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_874
timestamp 1626065694
transform 1 0 44133 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_873
timestamp 1626065694
transform 1 0 44469 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_872
timestamp 1626065694
transform 1 0 44805 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_871
timestamp 1626065694
transform 1 0 45141 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_870
timestamp 1626065694
transform 1 0 45477 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_869
timestamp 1626065694
transform 1 0 45813 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_868
timestamp 1626065694
transform 1 0 46149 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_867
timestamp 1626065694
transform 1 0 46485 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_866
timestamp 1626065694
transform 1 0 37749 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_865
timestamp 1626065694
transform 1 0 38085 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_864
timestamp 1626065694
transform 1 0 38421 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_863
timestamp 1626065694
transform 1 0 38757 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_862
timestamp 1626065694
transform 1 0 39093 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_861
timestamp 1626065694
transform 1 0 39429 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_860
timestamp 1626065694
transform 1 0 39765 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_859
timestamp 1626065694
transform 1 0 40101 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_858
timestamp 1626065694
transform 1 0 40437 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_857
timestamp 1626065694
transform 1 0 40773 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_856
timestamp 1626065694
transform 1 0 41109 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_855
timestamp 1626065694
transform 1 0 41445 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_854
timestamp 1626065694
transform 1 0 41781 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_853
timestamp 1626065694
transform 1 0 42117 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_852
timestamp 1626065694
transform 1 0 42453 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_851
timestamp 1626065694
transform 1 0 34389 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_850
timestamp 1626065694
transform 1 0 34725 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_849
timestamp 1626065694
transform 1 0 35061 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_848
timestamp 1626065694
transform 1 0 35397 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_847
timestamp 1626065694
transform 1 0 35733 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_846
timestamp 1626065694
transform 1 0 36069 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_845
timestamp 1626065694
transform 1 0 36405 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_844
timestamp 1626065694
transform 1 0 36741 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_843
timestamp 1626065694
transform 1 0 37077 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_842
timestamp 1626065694
transform 1 0 37413 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_841
timestamp 1626065694
transform 1 0 1797 0 1 72579
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_840
timestamp 1626065694
transform 1 0 17253 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_839
timestamp 1626065694
transform 1 0 25989 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_838
timestamp 1626065694
transform 1 0 26325 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_837
timestamp 1626065694
transform 1 0 26661 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_836
timestamp 1626065694
transform 1 0 26997 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_835
timestamp 1626065694
transform 1 0 27333 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_834
timestamp 1626065694
transform 1 0 27669 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_833
timestamp 1626065694
transform 1 0 28005 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_832
timestamp 1626065694
transform 1 0 28341 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_831
timestamp 1626065694
transform 1 0 28677 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_830
timestamp 1626065694
transform 1 0 29013 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_829
timestamp 1626065694
transform 1 0 29349 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_828
timestamp 1626065694
transform 1 0 29685 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_827
timestamp 1626065694
transform 1 0 30021 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_826
timestamp 1626065694
transform 1 0 30357 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_825
timestamp 1626065694
transform 1 0 30693 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_824
timestamp 1626065694
transform 1 0 31029 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_823
timestamp 1626065694
transform 1 0 31365 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_822
timestamp 1626065694
transform 1 0 31701 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_821
timestamp 1626065694
transform 1 0 32037 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_820
timestamp 1626065694
transform 1 0 32373 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_819
timestamp 1626065694
transform 1 0 32709 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_818
timestamp 1626065694
transform 1 0 33045 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_817
timestamp 1626065694
transform 1 0 33381 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_816
timestamp 1626065694
transform 1 0 33717 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_815
timestamp 1626065694
transform 1 0 34053 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_814
timestamp 1626065694
transform 1 0 25317 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_813
timestamp 1626065694
transform 1 0 25653 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_812
timestamp 1626065694
transform 1 0 17589 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_811
timestamp 1626065694
transform 1 0 17925 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_810
timestamp 1626065694
transform 1 0 18261 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_809
timestamp 1626065694
transform 1 0 18597 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_808
timestamp 1626065694
transform 1 0 18933 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_807
timestamp 1626065694
transform 1 0 19269 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_806
timestamp 1626065694
transform 1 0 19605 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_805
timestamp 1626065694
transform 1 0 19941 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_804
timestamp 1626065694
transform 1 0 20277 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_803
timestamp 1626065694
transform 1 0 20613 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_802
timestamp 1626065694
transform 1 0 20949 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_801
timestamp 1626065694
transform 1 0 21285 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_800
timestamp 1626065694
transform 1 0 21621 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_799
timestamp 1626065694
transform 1 0 21957 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_798
timestamp 1626065694
transform 1 0 22293 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_797
timestamp 1626065694
transform 1 0 22629 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_796
timestamp 1626065694
transform 1 0 22965 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_795
timestamp 1626065694
transform 1 0 23301 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_794
timestamp 1626065694
transform 1 0 23637 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_793
timestamp 1626065694
transform 1 0 23973 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_792
timestamp 1626065694
transform 1 0 24309 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_791
timestamp 1626065694
transform 1 0 24645 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_790
timestamp 1626065694
transform 1 0 24981 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_789
timestamp 1626065694
transform 1 0 9189 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_788
timestamp 1626065694
transform 1 0 9525 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_787
timestamp 1626065694
transform 1 0 9861 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_786
timestamp 1626065694
transform 1 0 10197 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_785
timestamp 1626065694
transform 1 0 10533 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_784
timestamp 1626065694
transform 1 0 10869 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_783
timestamp 1626065694
transform 1 0 11205 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_782
timestamp 1626065694
transform 1 0 11541 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_781
timestamp 1626065694
transform 1 0 11877 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_780
timestamp 1626065694
transform 1 0 12213 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_779
timestamp 1626065694
transform 1 0 12549 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_778
timestamp 1626065694
transform 1 0 12885 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_777
timestamp 1626065694
transform 1 0 13221 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_776
timestamp 1626065694
transform 1 0 13557 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_775
timestamp 1626065694
transform 1 0 13893 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_774
timestamp 1626065694
transform 1 0 14229 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_773
timestamp 1626065694
transform 1 0 14565 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_772
timestamp 1626065694
transform 1 0 14901 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_771
timestamp 1626065694
transform 1 0 15237 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_770
timestamp 1626065694
transform 1 0 15573 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_769
timestamp 1626065694
transform 1 0 15909 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_768
timestamp 1626065694
transform 1 0 16245 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_767
timestamp 1626065694
transform 1 0 16581 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_766
timestamp 1626065694
transform 1 0 16917 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_765
timestamp 1626065694
transform 1 0 8853 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_764
timestamp 1626065694
transform 1 0 4485 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_763
timestamp 1626065694
transform 1 0 4821 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_762
timestamp 1626065694
transform 1 0 5157 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_761
timestamp 1626065694
transform 1 0 5493 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_760
timestamp 1626065694
transform 1 0 5829 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_759
timestamp 1626065694
transform 1 0 6165 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_758
timestamp 1626065694
transform 1 0 6501 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_757
timestamp 1626065694
transform 1 0 6837 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_756
timestamp 1626065694
transform 1 0 7173 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_755
timestamp 1626065694
transform 1 0 7509 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_754
timestamp 1626065694
transform 1 0 7845 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_753
timestamp 1626065694
transform 1 0 8181 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_752
timestamp 1626065694
transform 1 0 8517 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_751
timestamp 1626065694
transform 1 0 3813 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_750
timestamp 1626065694
transform 1 0 4149 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_749
timestamp 1626065694
transform 1 0 1797 0 1 80643
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_748
timestamp 1626065694
transform 1 0 1797 0 1 80979
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_747
timestamp 1626065694
transform 1 0 2133 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_746
timestamp 1626065694
transform 1 0 2469 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_745
timestamp 1626065694
transform 1 0 2805 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_744
timestamp 1626065694
transform 1 0 3141 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_743
timestamp 1626065694
transform 1 0 3477 0 1 81432
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_742
timestamp 1626065694
transform 1 0 1797 0 1 78963
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_741
timestamp 1626065694
transform 1 0 1797 0 1 79299
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_740
timestamp 1626065694
transform 1 0 1797 0 1 79635
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_739
timestamp 1626065694
transform 1 0 1797 0 1 79971
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_738
timestamp 1626065694
transform 1 0 1797 0 1 80307
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_737
timestamp 1626065694
transform 1 0 1797 0 1 77955
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_736
timestamp 1626065694
transform 1 0 1797 0 1 78291
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_735
timestamp 1626065694
transform 1 0 1797 0 1 78627
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_734
timestamp 1626065694
transform 1 0 1797 0 1 73251
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_733
timestamp 1626065694
transform 1 0 1797 0 1 73587
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_732
timestamp 1626065694
transform 1 0 1797 0 1 76947
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_731
timestamp 1626065694
transform 1 0 1797 0 1 73923
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_730
timestamp 1626065694
transform 1 0 1797 0 1 74259
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_729
timestamp 1626065694
transform 1 0 1797 0 1 74595
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_728
timestamp 1626065694
transform 1 0 1797 0 1 74931
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_727
timestamp 1626065694
transform 1 0 1797 0 1 75267
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_726
timestamp 1626065694
transform 1 0 1797 0 1 75603
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_725
timestamp 1626065694
transform 1 0 1797 0 1 75939
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_724
timestamp 1626065694
transform 1 0 1797 0 1 77283
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_723
timestamp 1626065694
transform 1 0 1797 0 1 76275
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_722
timestamp 1626065694
transform 1 0 1797 0 1 76611
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_721
timestamp 1626065694
transform 1 0 1797 0 1 72915
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_720
timestamp 1626065694
transform 1 0 1797 0 1 77619
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_719
timestamp 1626065694
transform 1 0 1797 0 1 67539
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_718
timestamp 1626065694
transform 1 0 1797 0 1 69555
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_717
timestamp 1626065694
transform 1 0 1797 0 1 69891
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_716
timestamp 1626065694
transform 1 0 1797 0 1 70227
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_715
timestamp 1626065694
transform 1 0 1797 0 1 70563
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_714
timestamp 1626065694
transform 1 0 1797 0 1 70899
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_713
timestamp 1626065694
transform 1 0 1797 0 1 71235
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_712
timestamp 1626065694
transform 1 0 1797 0 1 71571
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_711
timestamp 1626065694
transform 1 0 1797 0 1 71907
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_710
timestamp 1626065694
transform 1 0 1797 0 1 72243
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_709
timestamp 1626065694
transform 1 0 1797 0 1 68547
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_708
timestamp 1626065694
transform 1 0 1797 0 1 68883
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_707
timestamp 1626065694
transform 1 0 1797 0 1 69219
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_706
timestamp 1626065694
transform 1 0 1797 0 1 67875
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_705
timestamp 1626065694
transform 1 0 1797 0 1 68211
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_704
timestamp 1626065694
transform 1 0 1797 0 1 63843
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_703
timestamp 1626065694
transform 1 0 1797 0 1 64179
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_702
timestamp 1626065694
transform 1 0 1797 0 1 64515
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_701
timestamp 1626065694
transform 1 0 1797 0 1 64851
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_700
timestamp 1626065694
transform 1 0 1797 0 1 65187
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_699
timestamp 1626065694
transform 1 0 1797 0 1 65523
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_698
timestamp 1626065694
transform 1 0 1797 0 1 65859
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_697
timestamp 1626065694
transform 1 0 1797 0 1 66195
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_696
timestamp 1626065694
transform 1 0 1797 0 1 66531
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_695
timestamp 1626065694
transform 1 0 1797 0 1 62499
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_694
timestamp 1626065694
transform 1 0 1797 0 1 66867
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_693
timestamp 1626065694
transform 1 0 1797 0 1 67203
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_692
timestamp 1626065694
transform 1 0 1797 0 1 62835
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_691
timestamp 1626065694
transform 1 0 1797 0 1 63171
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_690
timestamp 1626065694
transform 1 0 1797 0 1 63507
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_689
timestamp 1626065694
transform 1 0 1797 0 1 57123
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_688
timestamp 1626065694
transform 1 0 1797 0 1 57459
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_687
timestamp 1626065694
transform 1 0 1797 0 1 57795
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_686
timestamp 1626065694
transform 1 0 1797 0 1 58131
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_685
timestamp 1626065694
transform 1 0 1797 0 1 58467
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_684
timestamp 1626065694
transform 1 0 1797 0 1 58803
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_683
timestamp 1626065694
transform 1 0 1797 0 1 59139
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_682
timestamp 1626065694
transform 1 0 1797 0 1 59475
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_681
timestamp 1626065694
transform 1 0 1797 0 1 59811
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_680
timestamp 1626065694
transform 1 0 1797 0 1 60147
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_679
timestamp 1626065694
transform 1 0 1797 0 1 60483
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_678
timestamp 1626065694
transform 1 0 1797 0 1 60819
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_677
timestamp 1626065694
transform 1 0 1797 0 1 61155
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_676
timestamp 1626065694
transform 1 0 1797 0 1 61491
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_675
timestamp 1626065694
transform 1 0 1797 0 1 61827
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_674
timestamp 1626065694
transform 1 0 1797 0 1 62163
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_673
timestamp 1626065694
transform 1 0 1797 0 1 56787
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_672
timestamp 1626065694
transform 1 0 1797 0 1 54435
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_671
timestamp 1626065694
transform 1 0 1797 0 1 54771
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_670
timestamp 1626065694
transform 1 0 1797 0 1 55107
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_669
timestamp 1626065694
transform 1 0 1797 0 1 55443
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_668
timestamp 1626065694
transform 1 0 1797 0 1 55779
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_667
timestamp 1626065694
transform 1 0 1797 0 1 56115
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_666
timestamp 1626065694
transform 1 0 1797 0 1 56451
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_665
timestamp 1626065694
transform 1 0 1797 0 1 52419
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_664
timestamp 1626065694
transform 1 0 1797 0 1 52083
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_663
timestamp 1626065694
transform 1 0 1797 0 1 52755
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_662
timestamp 1626065694
transform 1 0 1797 0 1 53091
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_661
timestamp 1626065694
transform 1 0 1797 0 1 53427
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_660
timestamp 1626065694
transform 1 0 1797 0 1 53763
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_659
timestamp 1626065694
transform 1 0 1797 0 1 54099
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_658
timestamp 1626065694
transform 1 0 1797 0 1 46707
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_657
timestamp 1626065694
transform 1 0 1797 0 1 50067
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_656
timestamp 1626065694
transform 1 0 1797 0 1 50739
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_655
timestamp 1626065694
transform 1 0 1797 0 1 51075
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_654
timestamp 1626065694
transform 1 0 1797 0 1 47043
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_653
timestamp 1626065694
transform 1 0 1797 0 1 47379
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_652
timestamp 1626065694
transform 1 0 1797 0 1 51411
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_651
timestamp 1626065694
transform 1 0 1797 0 1 51747
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_650
timestamp 1626065694
transform 1 0 1797 0 1 49395
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_649
timestamp 1626065694
transform 1 0 1797 0 1 47715
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_648
timestamp 1626065694
transform 1 0 1797 0 1 49731
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_647
timestamp 1626065694
transform 1 0 1797 0 1 50403
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_646
timestamp 1626065694
transform 1 0 1797 0 1 49059
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_645
timestamp 1626065694
transform 1 0 1797 0 1 48051
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_644
timestamp 1626065694
transform 1 0 1797 0 1 48387
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_643
timestamp 1626065694
transform 1 0 1797 0 1 48723
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_642
timestamp 1626065694
transform 1 0 1797 0 1 42003
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_641
timestamp 1626065694
transform 1 0 1797 0 1 46035
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_640
timestamp 1626065694
transform 1 0 1797 0 1 46371
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_639
timestamp 1626065694
transform 1 0 1797 0 1 42339
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_638
timestamp 1626065694
transform 1 0 1797 0 1 42675
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_637
timestamp 1626065694
transform 1 0 1797 0 1 43011
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_636
timestamp 1626065694
transform 1 0 1797 0 1 43347
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_635
timestamp 1626065694
transform 1 0 1797 0 1 43683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_634
timestamp 1626065694
transform 1 0 1797 0 1 44019
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_633
timestamp 1626065694
transform 1 0 1797 0 1 44355
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_632
timestamp 1626065694
transform 1 0 1797 0 1 44691
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_631
timestamp 1626065694
transform 1 0 1797 0 1 45027
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_630
timestamp 1626065694
transform 1 0 1797 0 1 45363
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_629
timestamp 1626065694
transform 1 0 1797 0 1 45699
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_628
timestamp 1626065694
transform 1 0 1797 0 1 31251
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_627
timestamp 1626065694
transform 1 0 1797 0 1 37635
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_626
timestamp 1626065694
transform 1 0 1797 0 1 37971
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_625
timestamp 1626065694
transform 1 0 1797 0 1 38307
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_624
timestamp 1626065694
transform 1 0 1797 0 1 38643
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_623
timestamp 1626065694
transform 1 0 1797 0 1 38979
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_622
timestamp 1626065694
transform 1 0 1797 0 1 39315
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_621
timestamp 1626065694
transform 1 0 1797 0 1 39651
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_620
timestamp 1626065694
transform 1 0 1797 0 1 39987
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_619
timestamp 1626065694
transform 1 0 1797 0 1 40323
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_618
timestamp 1626065694
transform 1 0 1797 0 1 40659
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_617
timestamp 1626065694
transform 1 0 1797 0 1 40995
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_616
timestamp 1626065694
transform 1 0 1797 0 1 41331
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_615
timestamp 1626065694
transform 1 0 1797 0 1 37299
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_614
timestamp 1626065694
transform 1 0 1797 0 1 36627
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_613
timestamp 1626065694
transform 1 0 1797 0 1 36963
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_612
timestamp 1626065694
transform 1 0 1797 0 1 32259
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_611
timestamp 1626065694
transform 1 0 1797 0 1 32595
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_610
timestamp 1626065694
transform 1 0 1797 0 1 32931
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_609
timestamp 1626065694
transform 1 0 1797 0 1 33267
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_608
timestamp 1626065694
transform 1 0 1797 0 1 33603
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_607
timestamp 1626065694
transform 1 0 1797 0 1 33939
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_606
timestamp 1626065694
transform 1 0 1797 0 1 34275
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_605
timestamp 1626065694
transform 1 0 1797 0 1 34611
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_604
timestamp 1626065694
transform 1 0 1797 0 1 34947
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_603
timestamp 1626065694
transform 1 0 1797 0 1 31587
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_602
timestamp 1626065694
transform 1 0 1797 0 1 35283
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_601
timestamp 1626065694
transform 1 0 1797 0 1 35619
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_600
timestamp 1626065694
transform 1 0 1797 0 1 35955
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_599
timestamp 1626065694
transform 1 0 1797 0 1 36291
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_598
timestamp 1626065694
transform 1 0 1797 0 1 31923
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_597
timestamp 1626065694
transform 1 0 1797 0 1 26547
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_596
timestamp 1626065694
transform 1 0 1797 0 1 26883
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_595
timestamp 1626065694
transform 1 0 1797 0 1 27219
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_594
timestamp 1626065694
transform 1 0 1797 0 1 27555
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_593
timestamp 1626065694
transform 1 0 1797 0 1 30915
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_592
timestamp 1626065694
transform 1 0 1797 0 1 27891
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_591
timestamp 1626065694
transform 1 0 1797 0 1 28227
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_590
timestamp 1626065694
transform 1 0 1797 0 1 30243
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_589
timestamp 1626065694
transform 1 0 1797 0 1 28563
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_588
timestamp 1626065694
transform 1 0 1797 0 1 28899
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_587
timestamp 1626065694
transform 1 0 1797 0 1 29235
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_586
timestamp 1626065694
transform 1 0 1797 0 1 29571
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_585
timestamp 1626065694
transform 1 0 1797 0 1 30579
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_584
timestamp 1626065694
transform 1 0 1797 0 1 29907
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_583
timestamp 1626065694
transform 1 0 1797 0 1 26211
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_582
timestamp 1626065694
transform 1 0 1797 0 1 22851
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_581
timestamp 1626065694
transform 1 0 1797 0 1 23187
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_580
timestamp 1626065694
transform 1 0 1797 0 1 21843
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_579
timestamp 1626065694
transform 1 0 1797 0 1 23523
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_578
timestamp 1626065694
transform 1 0 1797 0 1 23859
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_577
timestamp 1626065694
transform 1 0 1797 0 1 22179
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_576
timestamp 1626065694
transform 1 0 1797 0 1 25539
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_575
timestamp 1626065694
transform 1 0 1797 0 1 25875
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_574
timestamp 1626065694
transform 1 0 1797 0 1 24531
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_573
timestamp 1626065694
transform 1 0 1797 0 1 22515
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_572
timestamp 1626065694
transform 1 0 1797 0 1 25203
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_571
timestamp 1626065694
transform 1 0 1797 0 1 24867
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_570
timestamp 1626065694
transform 1 0 1797 0 1 21171
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_569
timestamp 1626065694
transform 1 0 1797 0 1 21507
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_568
timestamp 1626065694
transform 1 0 1797 0 1 24195
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_567
timestamp 1626065694
transform 1 0 17253 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_566
timestamp 1626065694
transform 1 0 1797 0 1 15795
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_565
timestamp 1626065694
transform 1 0 1797 0 1 17475
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_564
timestamp 1626065694
transform 1 0 1797 0 1 17811
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_563
timestamp 1626065694
transform 1 0 1797 0 1 18147
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_562
timestamp 1626065694
transform 1 0 1797 0 1 18483
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_561
timestamp 1626065694
transform 1 0 1797 0 1 18819
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_560
timestamp 1626065694
transform 1 0 1797 0 1 19155
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_559
timestamp 1626065694
transform 1 0 1797 0 1 19491
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_558
timestamp 1626065694
transform 1 0 1797 0 1 19827
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_557
timestamp 1626065694
transform 1 0 1797 0 1 20163
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_556
timestamp 1626065694
transform 1 0 1797 0 1 20499
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_555
timestamp 1626065694
transform 1 0 1797 0 1 20835
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_554
timestamp 1626065694
transform 1 0 1797 0 1 16467
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_553
timestamp 1626065694
transform 1 0 1797 0 1 16803
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_552
timestamp 1626065694
transform 1 0 1797 0 1 17139
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_551
timestamp 1626065694
transform 1 0 1797 0 1 16131
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_550
timestamp 1626065694
transform 1 0 1797 0 1 13779
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_549
timestamp 1626065694
transform 1 0 1797 0 1 11763
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_548
timestamp 1626065694
transform 1 0 1797 0 1 12099
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_547
timestamp 1626065694
transform 1 0 1797 0 1 14115
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_546
timestamp 1626065694
transform 1 0 1797 0 1 12435
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_545
timestamp 1626065694
transform 1 0 1797 0 1 12771
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_544
timestamp 1626065694
transform 1 0 1797 0 1 14451
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_543
timestamp 1626065694
transform 1 0 1797 0 1 13107
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_542
timestamp 1626065694
transform 1 0 1797 0 1 10755
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_541
timestamp 1626065694
transform 1 0 1797 0 1 14787
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_540
timestamp 1626065694
transform 1 0 1797 0 1 11091
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_539
timestamp 1626065694
transform 1 0 1797 0 1 11427
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_538
timestamp 1626065694
transform 1 0 1797 0 1 15123
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_537
timestamp 1626065694
transform 1 0 1797 0 1 15459
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_536
timestamp 1626065694
transform 1 0 1797 0 1 13443
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_535
timestamp 1626065694
transform 1 0 1797 0 1 5379
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_534
timestamp 1626065694
transform 1 0 1797 0 1 5715
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_533
timestamp 1626065694
transform 1 0 1797 0 1 6051
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_532
timestamp 1626065694
transform 1 0 1797 0 1 6387
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_531
timestamp 1626065694
transform 1 0 1797 0 1 6723
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_530
timestamp 1626065694
transform 1 0 1797 0 1 7059
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_529
timestamp 1626065694
transform 1 0 1797 0 1 7395
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_528
timestamp 1626065694
transform 1 0 1797 0 1 7731
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_527
timestamp 1626065694
transform 1 0 1797 0 1 8067
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_526
timestamp 1626065694
transform 1 0 1797 0 1 8403
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_525
timestamp 1626065694
transform 1 0 1797 0 1 8739
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_524
timestamp 1626065694
transform 1 0 1797 0 1 9075
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_523
timestamp 1626065694
transform 1 0 1797 0 1 9411
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_522
timestamp 1626065694
transform 1 0 1797 0 1 9747
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_521
timestamp 1626065694
transform 1 0 1797 0 1 10083
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_520
timestamp 1626065694
transform 1 0 1797 0 1 10419
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_519
timestamp 1626065694
transform 1 0 4485 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_518
timestamp 1626065694
transform 1 0 1797 0 1 4707
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_517
timestamp 1626065694
transform 1 0 1797 0 1 5043
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_516
timestamp 1626065694
transform 1 0 1797 0 1 3027
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_515
timestamp 1626065694
transform 1 0 1797 0 1 3363
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_514
timestamp 1626065694
transform 1 0 1797 0 1 3699
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_513
timestamp 1626065694
transform 1 0 1797 0 1 4035
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_512
timestamp 1626065694
transform 1 0 1797 0 1 4371
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_511
timestamp 1626065694
transform 1 0 1797 0 1 2019
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_510
timestamp 1626065694
transform 1 0 1797 0 1 2355
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_509
timestamp 1626065694
transform 1 0 1797 0 1 2691
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_508
timestamp 1626065694
transform 1 0 2133 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_507
timestamp 1626065694
transform 1 0 2469 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_506
timestamp 1626065694
transform 1 0 2805 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_505
timestamp 1626065694
transform 1 0 3141 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_504
timestamp 1626065694
transform 1 0 3477 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_503
timestamp 1626065694
transform 1 0 3813 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_502
timestamp 1626065694
transform 1 0 4149 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_501
timestamp 1626065694
transform 1 0 8181 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_500
timestamp 1626065694
transform 1 0 7509 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_499
timestamp 1626065694
transform 1 0 5493 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_498
timestamp 1626065694
transform 1 0 8517 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_497
timestamp 1626065694
transform 1 0 7845 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_496
timestamp 1626065694
transform 1 0 6501 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_495
timestamp 1626065694
transform 1 0 6837 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_494
timestamp 1626065694
transform 1 0 7173 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_493
timestamp 1626065694
transform 1 0 6165 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_492
timestamp 1626065694
transform 1 0 5157 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_491
timestamp 1626065694
transform 1 0 5829 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_490
timestamp 1626065694
transform 1 0 4821 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_489
timestamp 1626065694
transform 1 0 13893 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_488
timestamp 1626065694
transform 1 0 14229 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_487
timestamp 1626065694
transform 1 0 14565 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_486
timestamp 1626065694
transform 1 0 14901 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_485
timestamp 1626065694
transform 1 0 15237 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_484
timestamp 1626065694
transform 1 0 15573 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_483
timestamp 1626065694
transform 1 0 15909 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_482
timestamp 1626065694
transform 1 0 10533 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_481
timestamp 1626065694
transform 1 0 16245 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_480
timestamp 1626065694
transform 1 0 16581 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_479
timestamp 1626065694
transform 1 0 16917 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_478
timestamp 1626065694
transform 1 0 10869 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_477
timestamp 1626065694
transform 1 0 11205 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_476
timestamp 1626065694
transform 1 0 11541 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_475
timestamp 1626065694
transform 1 0 11877 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_474
timestamp 1626065694
transform 1 0 9861 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_473
timestamp 1626065694
transform 1 0 12213 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_472
timestamp 1626065694
transform 1 0 12549 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_471
timestamp 1626065694
transform 1 0 12885 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_470
timestamp 1626065694
transform 1 0 13221 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_469
timestamp 1626065694
transform 1 0 9525 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_468
timestamp 1626065694
transform 1 0 10197 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_467
timestamp 1626065694
transform 1 0 13557 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_466
timestamp 1626065694
transform 1 0 8853 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_465
timestamp 1626065694
transform 1 0 9189 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_464
timestamp 1626065694
transform 1 0 18933 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_463
timestamp 1626065694
transform 1 0 20949 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_462
timestamp 1626065694
transform 1 0 17589 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_461
timestamp 1626065694
transform 1 0 21285 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_460
timestamp 1626065694
transform 1 0 21621 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_459
timestamp 1626065694
transform 1 0 21957 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_458
timestamp 1626065694
transform 1 0 17925 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_457
timestamp 1626065694
transform 1 0 22293 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_456
timestamp 1626065694
transform 1 0 19269 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_455
timestamp 1626065694
transform 1 0 22629 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_454
timestamp 1626065694
transform 1 0 19605 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_453
timestamp 1626065694
transform 1 0 22965 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_452
timestamp 1626065694
transform 1 0 23301 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_451
timestamp 1626065694
transform 1 0 23637 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_450
timestamp 1626065694
transform 1 0 23973 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_449
timestamp 1626065694
transform 1 0 24309 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_448
timestamp 1626065694
transform 1 0 24645 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_447
timestamp 1626065694
transform 1 0 24981 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_446
timestamp 1626065694
transform 1 0 25317 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_445
timestamp 1626065694
transform 1 0 25653 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_444
timestamp 1626065694
transform 1 0 19941 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_443
timestamp 1626065694
transform 1 0 20277 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_442
timestamp 1626065694
transform 1 0 20613 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_441
timestamp 1626065694
transform 1 0 18261 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_440
timestamp 1626065694
transform 1 0 18597 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_439
timestamp 1626065694
transform 1 0 33381 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_438
timestamp 1626065694
transform 1 0 33717 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_437
timestamp 1626065694
transform 1 0 29349 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_436
timestamp 1626065694
transform 1 0 34053 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_435
timestamp 1626065694
transform 1 0 29685 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_434
timestamp 1626065694
transform 1 0 30021 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_433
timestamp 1626065694
transform 1 0 30357 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_432
timestamp 1626065694
transform 1 0 25989 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_431
timestamp 1626065694
transform 1 0 30693 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_430
timestamp 1626065694
transform 1 0 31029 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_429
timestamp 1626065694
transform 1 0 26325 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_428
timestamp 1626065694
transform 1 0 31365 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_427
timestamp 1626065694
transform 1 0 26661 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_426
timestamp 1626065694
transform 1 0 31701 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_425
timestamp 1626065694
transform 1 0 28341 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_424
timestamp 1626065694
transform 1 0 26997 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_423
timestamp 1626065694
transform 1 0 27333 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_422
timestamp 1626065694
transform 1 0 32037 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_421
timestamp 1626065694
transform 1 0 32373 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_420
timestamp 1626065694
transform 1 0 28677 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_419
timestamp 1626065694
transform 1 0 32709 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_418
timestamp 1626065694
transform 1 0 33045 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_417
timestamp 1626065694
transform 1 0 29013 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_416
timestamp 1626065694
transform 1 0 27669 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_415
timestamp 1626065694
transform 1 0 28005 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_414
timestamp 1626065694
transform 1 0 42789 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_413
timestamp 1626065694
transform 1 0 40101 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_412
timestamp 1626065694
transform 1 0 40437 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_411
timestamp 1626065694
transform 1 0 40773 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_410
timestamp 1626065694
transform 1 0 41109 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_409
timestamp 1626065694
transform 1 0 41445 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_408
timestamp 1626065694
transform 1 0 41781 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_407
timestamp 1626065694
transform 1 0 42117 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_406
timestamp 1626065694
transform 1 0 42453 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_405
timestamp 1626065694
transform 1 0 39765 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_404
timestamp 1626065694
transform 1 0 34725 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_403
timestamp 1626065694
transform 1 0 35061 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_402
timestamp 1626065694
transform 1 0 35397 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_401
timestamp 1626065694
transform 1 0 34389 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_400
timestamp 1626065694
transform 1 0 35733 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_399
timestamp 1626065694
transform 1 0 36069 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_398
timestamp 1626065694
transform 1 0 36405 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_397
timestamp 1626065694
transform 1 0 36741 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_396
timestamp 1626065694
transform 1 0 37077 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_395
timestamp 1626065694
transform 1 0 37413 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_394
timestamp 1626065694
transform 1 0 37749 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_393
timestamp 1626065694
transform 1 0 38085 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_392
timestamp 1626065694
transform 1 0 38421 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_391
timestamp 1626065694
transform 1 0 38757 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_390
timestamp 1626065694
transform 1 0 39093 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_389
timestamp 1626065694
transform 1 0 39429 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_388
timestamp 1626065694
transform 1 0 48165 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_387
timestamp 1626065694
transform 1 0 48501 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_386
timestamp 1626065694
transform 1 0 48837 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_385
timestamp 1626065694
transform 1 0 49173 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_384
timestamp 1626065694
transform 1 0 49509 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_383
timestamp 1626065694
transform 1 0 44469 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_382
timestamp 1626065694
transform 1 0 44805 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_381
timestamp 1626065694
transform 1 0 49845 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_380
timestamp 1626065694
transform 1 0 50181 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_379
timestamp 1626065694
transform 1 0 50517 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_378
timestamp 1626065694
transform 1 0 50853 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_377
timestamp 1626065694
transform 1 0 45141 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_376
timestamp 1626065694
transform 1 0 43125 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_375
timestamp 1626065694
transform 1 0 45477 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_374
timestamp 1626065694
transform 1 0 45813 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_373
timestamp 1626065694
transform 1 0 51189 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_372
timestamp 1626065694
transform 1 0 46149 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_371
timestamp 1626065694
transform 1 0 43461 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_370
timestamp 1626065694
transform 1 0 43797 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_369
timestamp 1626065694
transform 1 0 46485 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_368
timestamp 1626065694
transform 1 0 46821 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_367
timestamp 1626065694
transform 1 0 47157 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_366
timestamp 1626065694
transform 1 0 47493 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_365
timestamp 1626065694
transform 1 0 44133 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_364
timestamp 1626065694
transform 1 0 47829 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_363
timestamp 1626065694
transform 1 0 59253 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_362
timestamp 1626065694
transform 1 0 58581 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_361
timestamp 1626065694
transform 1 0 57909 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_360
timestamp 1626065694
transform 1 0 59589 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_359
timestamp 1626065694
transform 1 0 57573 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_358
timestamp 1626065694
transform 1 0 51525 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_357
timestamp 1626065694
transform 1 0 51861 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_356
timestamp 1626065694
transform 1 0 52197 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_355
timestamp 1626065694
transform 1 0 52533 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_354
timestamp 1626065694
transform 1 0 52869 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_353
timestamp 1626065694
transform 1 0 53205 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_352
timestamp 1626065694
transform 1 0 53541 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_351
timestamp 1626065694
transform 1 0 53877 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_350
timestamp 1626065694
transform 1 0 54213 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_349
timestamp 1626065694
transform 1 0 54549 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_348
timestamp 1626065694
transform 1 0 54885 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_347
timestamp 1626065694
transform 1 0 58245 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_346
timestamp 1626065694
transform 1 0 55221 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_345
timestamp 1626065694
transform 1 0 55557 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_344
timestamp 1626065694
transform 1 0 58917 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_343
timestamp 1626065694
transform 1 0 55893 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_342
timestamp 1626065694
transform 1 0 56229 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_341
timestamp 1626065694
transform 1 0 56565 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_340
timestamp 1626065694
transform 1 0 56901 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_339
timestamp 1626065694
transform 1 0 57237 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_338
timestamp 1626065694
transform 1 0 61605 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_337
timestamp 1626065694
transform 1 0 64965 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_336
timestamp 1626065694
transform 1 0 66309 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_335
timestamp 1626065694
transform 1 0 65637 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_334
timestamp 1626065694
transform 1 0 66645 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_333
timestamp 1626065694
transform 1 0 66981 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_332
timestamp 1626065694
transform 1 0 67989 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_331
timestamp 1626065694
transform 1 0 65973 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_330
timestamp 1626065694
transform 1 0 64293 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_329
timestamp 1626065694
transform 1 0 61941 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_328
timestamp 1626065694
transform 1 0 67317 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_327
timestamp 1626065694
transform 1 0 59925 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_326
timestamp 1626065694
transform 1 0 67653 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_325
timestamp 1626065694
transform 1 0 62613 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_324
timestamp 1626065694
transform 1 0 63621 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_323
timestamp 1626065694
transform 1 0 63957 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_322
timestamp 1626065694
transform 1 0 60597 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_321
timestamp 1626065694
transform 1 0 62277 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_320
timestamp 1626065694
transform 1 0 64629 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_319
timestamp 1626065694
transform 1 0 65301 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_318
timestamp 1626065694
transform 1 0 61269 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_317
timestamp 1626065694
transform 1 0 62949 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_316
timestamp 1626065694
transform 1 0 60933 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_315
timestamp 1626065694
transform 1 0 63285 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_314
timestamp 1626065694
transform 1 0 60261 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_313
timestamp 1626065694
transform 1 0 102261 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_312
timestamp 1626065694
transform 1 0 134847 0 1 31251
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_311
timestamp 1626065694
transform 1 0 134847 0 1 36627
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_310
timestamp 1626065694
transform 1 0 134847 0 1 36963
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_309
timestamp 1626065694
transform 1 0 134847 0 1 37299
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_308
timestamp 1626065694
transform 1 0 134847 0 1 37635
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_307
timestamp 1626065694
transform 1 0 134847 0 1 37971
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_306
timestamp 1626065694
transform 1 0 134847 0 1 38307
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_305
timestamp 1626065694
transform 1 0 134847 0 1 38643
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_304
timestamp 1626065694
transform 1 0 134847 0 1 38979
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_303
timestamp 1626065694
transform 1 0 134847 0 1 39315
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_302
timestamp 1626065694
transform 1 0 134847 0 1 39651
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_301
timestamp 1626065694
transform 1 0 134847 0 1 39987
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_300
timestamp 1626065694
transform 1 0 134847 0 1 40323
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_299
timestamp 1626065694
transform 1 0 134847 0 1 40659
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_298
timestamp 1626065694
transform 1 0 134847 0 1 40995
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_297
timestamp 1626065694
transform 1 0 134847 0 1 41331
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_296
timestamp 1626065694
transform 1 0 134847 0 1 31923
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_295
timestamp 1626065694
transform 1 0 134847 0 1 32259
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_294
timestamp 1626065694
transform 1 0 134847 0 1 32595
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_293
timestamp 1626065694
transform 1 0 134847 0 1 32931
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_292
timestamp 1626065694
transform 1 0 134847 0 1 33267
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_291
timestamp 1626065694
transform 1 0 134847 0 1 33603
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_290
timestamp 1626065694
transform 1 0 134847 0 1 33939
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_289
timestamp 1626065694
transform 1 0 134847 0 1 31587
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_288
timestamp 1626065694
transform 1 0 134847 0 1 34275
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_287
timestamp 1626065694
transform 1 0 134847 0 1 34611
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_286
timestamp 1626065694
transform 1 0 134847 0 1 34947
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_285
timestamp 1626065694
transform 1 0 134847 0 1 35283
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_284
timestamp 1626065694
transform 1 0 134847 0 1 35619
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_283
timestamp 1626065694
transform 1 0 134847 0 1 35955
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_282
timestamp 1626065694
transform 1 0 134847 0 1 36291
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_281
timestamp 1626065694
transform 1 0 134847 0 1 27555
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_280
timestamp 1626065694
transform 1 0 134847 0 1 27891
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_279
timestamp 1626065694
transform 1 0 134847 0 1 28227
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_278
timestamp 1626065694
transform 1 0 134847 0 1 28563
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_277
timestamp 1626065694
transform 1 0 134847 0 1 28899
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_276
timestamp 1626065694
transform 1 0 134847 0 1 29235
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_275
timestamp 1626065694
transform 1 0 134847 0 1 29571
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_274
timestamp 1626065694
transform 1 0 134847 0 1 29907
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_273
timestamp 1626065694
transform 1 0 134847 0 1 30243
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_272
timestamp 1626065694
transform 1 0 134847 0 1 30579
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_271
timestamp 1626065694
transform 1 0 134847 0 1 30915
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_270
timestamp 1626065694
transform 1 0 134847 0 1 26211
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_269
timestamp 1626065694
transform 1 0 134847 0 1 26547
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_268
timestamp 1626065694
transform 1 0 134847 0 1 26883
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_267
timestamp 1626065694
transform 1 0 134847 0 1 27219
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_266
timestamp 1626065694
transform 1 0 134847 0 1 21507
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_265
timestamp 1626065694
transform 1 0 134847 0 1 22851
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_264
timestamp 1626065694
transform 1 0 134847 0 1 21843
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_263
timestamp 1626065694
transform 1 0 134847 0 1 23187
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_262
timestamp 1626065694
transform 1 0 134847 0 1 22179
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_261
timestamp 1626065694
transform 1 0 134847 0 1 25203
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_260
timestamp 1626065694
transform 1 0 134847 0 1 25539
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_259
timestamp 1626065694
transform 1 0 134847 0 1 25875
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_258
timestamp 1626065694
transform 1 0 134847 0 1 23523
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_257
timestamp 1626065694
transform 1 0 134847 0 1 23859
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_256
timestamp 1626065694
transform 1 0 134847 0 1 24195
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_255
timestamp 1626065694
transform 1 0 134847 0 1 24531
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_254
timestamp 1626065694
transform 1 0 134847 0 1 24867
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_253
timestamp 1626065694
transform 1 0 134847 0 1 22515
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_252
timestamp 1626065694
transform 1 0 134847 0 1 21171
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_251
timestamp 1626065694
transform 1 0 76725 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_250
timestamp 1626065694
transform 1 0 76389 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_249
timestamp 1626065694
transform 1 0 75717 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_248
timestamp 1626065694
transform 1 0 68661 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_247
timestamp 1626065694
transform 1 0 68997 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_246
timestamp 1626065694
transform 1 0 69333 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_245
timestamp 1626065694
transform 1 0 69669 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_244
timestamp 1626065694
transform 1 0 70005 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_243
timestamp 1626065694
transform 1 0 70341 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_242
timestamp 1626065694
transform 1 0 70677 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_241
timestamp 1626065694
transform 1 0 71013 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_240
timestamp 1626065694
transform 1 0 71349 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_239
timestamp 1626065694
transform 1 0 71685 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_238
timestamp 1626065694
transform 1 0 72021 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_237
timestamp 1626065694
transform 1 0 72357 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_236
timestamp 1626065694
transform 1 0 72693 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_235
timestamp 1626065694
transform 1 0 73029 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_234
timestamp 1626065694
transform 1 0 73365 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_233
timestamp 1626065694
transform 1 0 73701 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_232
timestamp 1626065694
transform 1 0 74037 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_231
timestamp 1626065694
transform 1 0 76053 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_230
timestamp 1626065694
transform 1 0 74373 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_229
timestamp 1626065694
transform 1 0 74709 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_228
timestamp 1626065694
transform 1 0 75045 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_227
timestamp 1626065694
transform 1 0 75381 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_226
timestamp 1626065694
transform 1 0 78741 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_225
timestamp 1626065694
transform 1 0 83781 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_224
timestamp 1626065694
transform 1 0 77061 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_223
timestamp 1626065694
transform 1 0 79749 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_222
timestamp 1626065694
transform 1 0 80757 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_221
timestamp 1626065694
transform 1 0 82773 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_220
timestamp 1626065694
transform 1 0 81093 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_219
timestamp 1626065694
transform 1 0 78069 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_218
timestamp 1626065694
transform 1 0 81429 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_217
timestamp 1626065694
transform 1 0 84117 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_216
timestamp 1626065694
transform 1 0 81765 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_215
timestamp 1626065694
transform 1 0 77397 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_214
timestamp 1626065694
transform 1 0 84453 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_213
timestamp 1626065694
transform 1 0 77733 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_212
timestamp 1626065694
transform 1 0 82101 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_211
timestamp 1626065694
transform 1 0 83445 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_210
timestamp 1626065694
transform 1 0 83109 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_209
timestamp 1626065694
transform 1 0 84789 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_208
timestamp 1626065694
transform 1 0 82437 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_207
timestamp 1626065694
transform 1 0 78405 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_206
timestamp 1626065694
transform 1 0 79077 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_205
timestamp 1626065694
transform 1 0 85125 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_204
timestamp 1626065694
transform 1 0 80085 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_203
timestamp 1626065694
transform 1 0 79413 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_202
timestamp 1626065694
transform 1 0 80421 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_201
timestamp 1626065694
transform 1 0 93861 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_200
timestamp 1626065694
transform 1 0 86805 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_199
timestamp 1626065694
transform 1 0 87141 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_198
timestamp 1626065694
transform 1 0 87477 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_197
timestamp 1626065694
transform 1 0 87813 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_196
timestamp 1626065694
transform 1 0 90165 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_195
timestamp 1626065694
transform 1 0 90501 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_194
timestamp 1626065694
transform 1 0 90837 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_193
timestamp 1626065694
transform 1 0 93525 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_192
timestamp 1626065694
transform 1 0 88149 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_191
timestamp 1626065694
transform 1 0 91173 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_190
timestamp 1626065694
transform 1 0 88485 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_189
timestamp 1626065694
transform 1 0 91509 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_188
timestamp 1626065694
transform 1 0 88821 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_187
timestamp 1626065694
transform 1 0 89157 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_186
timestamp 1626065694
transform 1 0 89493 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_185
timestamp 1626065694
transform 1 0 91845 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_184
timestamp 1626065694
transform 1 0 89829 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_183
timestamp 1626065694
transform 1 0 93189 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_182
timestamp 1626065694
transform 1 0 92853 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_181
timestamp 1626065694
transform 1 0 92181 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_180
timestamp 1626065694
transform 1 0 85461 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_179
timestamp 1626065694
transform 1 0 85797 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_178
timestamp 1626065694
transform 1 0 86133 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_177
timestamp 1626065694
transform 1 0 86469 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_176
timestamp 1626065694
transform 1 0 92517 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_175
timestamp 1626065694
transform 1 0 99909 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_174
timestamp 1626065694
transform 1 0 99573 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_173
timestamp 1626065694
transform 1 0 94869 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_172
timestamp 1626065694
transform 1 0 98229 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_171
timestamp 1626065694
transform 1 0 98565 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_170
timestamp 1626065694
transform 1 0 98901 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_169
timestamp 1626065694
transform 1 0 95541 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_168
timestamp 1626065694
transform 1 0 95205 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_167
timestamp 1626065694
transform 1 0 95877 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_166
timestamp 1626065694
transform 1 0 100245 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_165
timestamp 1626065694
transform 1 0 96213 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_164
timestamp 1626065694
transform 1 0 100581 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_163
timestamp 1626065694
transform 1 0 99237 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_162
timestamp 1626065694
transform 1 0 100917 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_161
timestamp 1626065694
transform 1 0 101253 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_160
timestamp 1626065694
transform 1 0 94197 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_159
timestamp 1626065694
transform 1 0 101589 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_158
timestamp 1626065694
transform 1 0 96549 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_157
timestamp 1626065694
transform 1 0 96885 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_156
timestamp 1626065694
transform 1 0 101925 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_155
timestamp 1626065694
transform 1 0 94533 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_154
timestamp 1626065694
transform 1 0 97221 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_153
timestamp 1626065694
transform 1 0 97557 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_152
timestamp 1626065694
transform 1 0 97893 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_151
timestamp 1626065694
transform 1 0 119397 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_150
timestamp 1626065694
transform 1 0 134847 0 1 15795
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_149
timestamp 1626065694
transform 1 0 134847 0 1 16131
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_148
timestamp 1626065694
transform 1 0 134847 0 1 16467
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_147
timestamp 1626065694
transform 1 0 134847 0 1 16803
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_146
timestamp 1626065694
transform 1 0 134847 0 1 17139
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_145
timestamp 1626065694
transform 1 0 134847 0 1 17475
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_144
timestamp 1626065694
transform 1 0 134847 0 1 17811
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_143
timestamp 1626065694
transform 1 0 134847 0 1 18147
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_142
timestamp 1626065694
transform 1 0 134847 0 1 18483
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_141
timestamp 1626065694
transform 1 0 134847 0 1 18819
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_140
timestamp 1626065694
transform 1 0 134847 0 1 19155
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_139
timestamp 1626065694
transform 1 0 134847 0 1 19491
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_138
timestamp 1626065694
transform 1 0 134847 0 1 19827
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_137
timestamp 1626065694
transform 1 0 134847 0 1 20163
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_136
timestamp 1626065694
transform 1 0 134847 0 1 20499
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_135
timestamp 1626065694
transform 1 0 134847 0 1 20835
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_134
timestamp 1626065694
transform 1 0 134847 0 1 15459
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_133
timestamp 1626065694
transform 1 0 134847 0 1 10755
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_132
timestamp 1626065694
transform 1 0 134847 0 1 11091
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_131
timestamp 1626065694
transform 1 0 134847 0 1 11427
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_130
timestamp 1626065694
transform 1 0 134847 0 1 11763
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_129
timestamp 1626065694
transform 1 0 134847 0 1 12099
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_128
timestamp 1626065694
transform 1 0 134847 0 1 12435
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_127
timestamp 1626065694
transform 1 0 134847 0 1 12771
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_126
timestamp 1626065694
transform 1 0 134847 0 1 13107
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_125
timestamp 1626065694
transform 1 0 134847 0 1 13443
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_124
timestamp 1626065694
transform 1 0 134847 0 1 13779
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_123
timestamp 1626065694
transform 1 0 134847 0 1 14115
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_122
timestamp 1626065694
transform 1 0 134847 0 1 14451
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_121
timestamp 1626065694
transform 1 0 134847 0 1 14787
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_120
timestamp 1626065694
transform 1 0 134847 0 1 15123
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_119
timestamp 1626065694
transform 1 0 109317 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_118
timestamp 1626065694
transform 1 0 109653 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_117
timestamp 1626065694
transform 1 0 106293 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_116
timestamp 1626065694
transform 1 0 104613 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_115
timestamp 1626065694
transform 1 0 109989 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_114
timestamp 1626065694
transform 1 0 107973 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_113
timestamp 1626065694
transform 1 0 110325 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_112
timestamp 1626065694
transform 1 0 110661 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_111
timestamp 1626065694
transform 1 0 106629 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_110
timestamp 1626065694
transform 1 0 106965 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_109
timestamp 1626065694
transform 1 0 104949 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_108
timestamp 1626065694
transform 1 0 107301 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_107
timestamp 1626065694
transform 1 0 105285 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_106
timestamp 1626065694
transform 1 0 102597 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_105
timestamp 1626065694
transform 1 0 102933 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_104
timestamp 1626065694
transform 1 0 103269 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_103
timestamp 1626065694
transform 1 0 103605 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_102
timestamp 1626065694
transform 1 0 103941 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_101
timestamp 1626065694
transform 1 0 104277 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_100
timestamp 1626065694
transform 1 0 105621 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_99
timestamp 1626065694
transform 1 0 105957 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_98
timestamp 1626065694
transform 1 0 108309 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_97
timestamp 1626065694
transform 1 0 107637 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_96
timestamp 1626065694
transform 1 0 108645 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_95
timestamp 1626065694
transform 1 0 108981 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_94
timestamp 1626065694
transform 1 0 112005 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_93
timestamp 1626065694
transform 1 0 118053 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_92
timestamp 1626065694
transform 1 0 112341 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_91
timestamp 1626065694
transform 1 0 112677 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_90
timestamp 1626065694
transform 1 0 116037 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_89
timestamp 1626065694
transform 1 0 113013 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_88
timestamp 1626065694
transform 1 0 113349 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_87
timestamp 1626065694
transform 1 0 116709 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_86
timestamp 1626065694
transform 1 0 118389 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_85
timestamp 1626065694
transform 1 0 116373 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_84
timestamp 1626065694
transform 1 0 117045 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_83
timestamp 1626065694
transform 1 0 113685 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_82
timestamp 1626065694
transform 1 0 115701 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_81
timestamp 1626065694
transform 1 0 118725 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_80
timestamp 1626065694
transform 1 0 110997 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_79
timestamp 1626065694
transform 1 0 119061 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_78
timestamp 1626065694
transform 1 0 114021 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_77
timestamp 1626065694
transform 1 0 117381 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_76
timestamp 1626065694
transform 1 0 111333 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_75
timestamp 1626065694
transform 1 0 115365 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_74
timestamp 1626065694
transform 1 0 114357 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_73
timestamp 1626065694
transform 1 0 114693 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_72
timestamp 1626065694
transform 1 0 111669 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_71
timestamp 1626065694
transform 1 0 115029 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_70
timestamp 1626065694
transform 1 0 117717 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_69
timestamp 1626065694
transform 1 0 127797 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_68
timestamp 1626065694
transform 1 0 134847 0 1 5379
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_67
timestamp 1626065694
transform 1 0 134847 0 1 5715
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_66
timestamp 1626065694
transform 1 0 134847 0 1 6051
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_65
timestamp 1626065694
transform 1 0 134847 0 1 6387
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_64
timestamp 1626065694
transform 1 0 134847 0 1 6723
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_63
timestamp 1626065694
transform 1 0 134847 0 1 7059
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_62
timestamp 1626065694
transform 1 0 134847 0 1 7395
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_61
timestamp 1626065694
transform 1 0 134847 0 1 7731
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_60
timestamp 1626065694
transform 1 0 134847 0 1 8067
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_59
timestamp 1626065694
transform 1 0 134847 0 1 8403
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_58
timestamp 1626065694
transform 1 0 134847 0 1 8739
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_57
timestamp 1626065694
transform 1 0 134847 0 1 9075
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_56
timestamp 1626065694
transform 1 0 134847 0 1 9411
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_55
timestamp 1626065694
transform 1 0 134847 0 1 9747
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_54
timestamp 1626065694
transform 1 0 134847 0 1 10083
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_53
timestamp 1626065694
transform 1 0 134847 0 1 10419
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_52
timestamp 1626065694
transform 1 0 126789 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_51
timestamp 1626065694
transform 1 0 127125 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_50
timestamp 1626065694
transform 1 0 127461 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_49
timestamp 1626065694
transform 1 0 119733 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_48
timestamp 1626065694
transform 1 0 120069 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_47
timestamp 1626065694
transform 1 0 120405 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_46
timestamp 1626065694
transform 1 0 120741 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_45
timestamp 1626065694
transform 1 0 121077 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_44
timestamp 1626065694
transform 1 0 121413 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_43
timestamp 1626065694
transform 1 0 121749 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_42
timestamp 1626065694
transform 1 0 122085 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_41
timestamp 1626065694
transform 1 0 122421 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_40
timestamp 1626065694
transform 1 0 122757 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_39
timestamp 1626065694
transform 1 0 123093 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_38
timestamp 1626065694
transform 1 0 123429 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_37
timestamp 1626065694
transform 1 0 123765 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_36
timestamp 1626065694
transform 1 0 124101 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_35
timestamp 1626065694
transform 1 0 124437 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_34
timestamp 1626065694
transform 1 0 124773 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_33
timestamp 1626065694
transform 1 0 125109 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_32
timestamp 1626065694
transform 1 0 125445 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_31
timestamp 1626065694
transform 1 0 125781 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_30
timestamp 1626065694
transform 1 0 126117 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_29
timestamp 1626065694
transform 1 0 126453 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_28
timestamp 1626065694
transform 1 0 134847 0 1 4707
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_27
timestamp 1626065694
transform 1 0 134847 0 1 5043
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_26
timestamp 1626065694
transform 1 0 134847 0 1 4035
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_25
timestamp 1626065694
transform 1 0 134847 0 1 3699
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_24
timestamp 1626065694
transform 1 0 134847 0 1 4371
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_23
timestamp 1626065694
transform 1 0 134847 0 1 3363
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_22
timestamp 1626065694
transform 1 0 134847 0 1 3027
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_21
timestamp 1626065694
transform 1 0 128469 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_20
timestamp 1626065694
transform 1 0 128805 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_19
timestamp 1626065694
transform 1 0 129141 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_18
timestamp 1626065694
transform 1 0 129477 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_17
timestamp 1626065694
transform 1 0 129813 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_16
timestamp 1626065694
transform 1 0 130149 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_15
timestamp 1626065694
transform 1 0 130485 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_14
timestamp 1626065694
transform 1 0 130821 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_13
timestamp 1626065694
transform 1 0 131157 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_12
timestamp 1626065694
transform 1 0 131493 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_11
timestamp 1626065694
transform 1 0 131829 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_10
timestamp 1626065694
transform 1 0 128133 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_9
timestamp 1626065694
transform 1 0 133173 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_8
timestamp 1626065694
transform 1 0 133509 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_7
timestamp 1626065694
transform 1 0 134847 0 1 2019
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_6
timestamp 1626065694
transform 1 0 133845 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_5
timestamp 1626065694
transform 1 0 134181 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_4
timestamp 1626065694
transform 1 0 132165 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_3
timestamp 1626065694
transform 1 0 132501 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_2
timestamp 1626065694
transform 1 0 134847 0 1 2355
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_1
timestamp 1626065694
transform 1 0 132837 0 1 1683
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_0
timestamp 1626065694
transform 1 0 134847 0 1 2691
box -59 -43 109 125
use sky130_sram_2kbyte_1rw1r_32x512_8_bank  sky130_sram_2kbyte_1rw1r_32x512_8_bank_0
timestamp 1626065694
transform 1 0 14862 0 1 9422
box 0 0 107270 69282
<< labels >>
rlabel metal3 s 0 8024 212 8100 4 csb0
rlabel metal3 s 0 9928 212 10004 4 web0
rlabel metal3 s 0 8296 212 8372 4 clk0
rlabel metal3 s 0 28152 212 28228 4 addr0[2]
rlabel metal3 s 0 29920 212 29996 4 addr0[3]
rlabel metal3 s 0 31008 212 31084 4 addr0[4]
rlabel metal3 s 0 32776 212 32852 4 addr0[5]
rlabel metal3 s 0 33728 212 33804 4 addr0[6]
rlabel metal3 s 0 35904 212 35980 4 addr0[7]
rlabel metal3 s 0 36856 212 36932 4 addr0[8]
rlabel metal3 s 136408 79152 136620 79228 4 csb1
rlabel metal3 s 136408 19312 136620 19388 4 addr1[2]
rlabel metal3 s 136408 17680 136620 17756 4 addr1[3]
rlabel metal3 s 136408 16320 136620 16396 4 addr1[4]
rlabel metal3 s 136408 14824 136620 14900 4 addr1[5]
rlabel metal3 s 136408 13600 136620 13676 4 addr1[6]
rlabel metal3 s 952 82008 135668 82356 4 vccd1
rlabel metal3 s 952 952 135668 1300 4 vccd1
rlabel metal3 s 272 272 136348 620 4 vssd1
rlabel metal3 s 272 82688 136348 83036 4 vssd1
rlabel metal4 s 130832 83096 130908 83308 4 clk1
rlabel metal4 s 68544 83096 68620 83308 4 dout1[16]
rlabel metal4 s 70992 83096 71068 83308 4 dout1[17]
rlabel metal4 s 73576 83096 73652 83308 4 dout1[18]
rlabel metal4 s 75888 83096 75964 83308 4 dout1[19]
rlabel metal4 s 78608 83096 78684 83308 4 dout1[20]
rlabel metal4 s 81056 83096 81132 83308 4 dout1[21]
rlabel metal4 s 83504 83096 83580 83308 4 dout1[22]
rlabel metal4 s 85952 83096 86028 83308 4 dout1[23]
rlabel metal4 s 88400 83096 88476 83308 4 dout1[24]
rlabel metal4 s 90984 83096 91060 83308 4 dout1[25]
rlabel metal4 s 93568 83096 93644 83308 4 dout1[26]
rlabel metal4 s 96016 83096 96092 83308 4 dout1[27]
rlabel metal4 s 98464 83096 98540 83308 4 dout1[28]
rlabel metal4 s 101048 83096 101124 83308 4 dout1[29]
rlabel metal4 s 103360 83096 103436 83308 4 dout1[30]
rlabel metal4 s 106080 83096 106156 83308 4 dout1[31]
rlabel metal4 s 119680 83096 119756 83308 4 addr1[0]
rlabel metal4 s 118456 83096 118532 83308 4 addr1[1]
rlabel metal4 s 33456 83096 33532 83308 4 dout1[2]
rlabel metal4 s 36176 83096 36252 83308 4 dout1[3]
rlabel metal4 s 38488 83096 38564 83308 4 dout1[4]
rlabel metal4 s 41072 83096 41148 83308 4 dout1[5]
rlabel metal4 s 43520 83096 43596 83308 4 dout1[6]
rlabel metal4 s 46104 83096 46180 83308 4 dout1[7]
rlabel metal4 s 48552 83096 48628 83308 4 dout1[8]
rlabel metal4 s 51136 83096 51212 83308 4 dout1[9]
rlabel metal4 s 53584 83096 53660 83308 4 dout1[10]
rlabel metal4 s 56168 83096 56244 83308 4 dout1[11]
rlabel metal4 s 58480 83096 58556 83308 4 dout1[12]
rlabel metal4 s 60928 83096 61004 83308 4 dout1[13]
rlabel metal4 s 63648 83096 63724 83308 4 dout1[14]
rlabel metal4 s 66096 83096 66172 83308 4 dout1[15]
rlabel metal4 s 28696 83096 28772 83308 4 dout1[0]
rlabel metal4 s 31008 83096 31084 83308 4 dout1[1]
rlabel metal4 s 36040 0 36116 212 4 dout0[3]
rlabel metal4 s 38488 0 38564 212 4 dout0[4]
rlabel metal4 s 41072 0 41148 212 4 dout0[5]
rlabel metal4 s 43520 0 43596 212 4 dout0[6]
rlabel metal4 s 45968 0 46044 212 4 dout0[7]
rlabel metal4 s 48280 0 48356 212 4 dout0[8]
rlabel metal4 s 51000 0 51076 212 4 dout0[9]
rlabel metal4 s 53584 0 53660 212 4 dout0[10]
rlabel metal4 s 56032 0 56108 212 4 dout0[11]
rlabel metal4 s 58480 0 58556 212 4 dout0[12]
rlabel metal4 s 60928 0 61004 212 4 dout0[13]
rlabel metal4 s 63512 0 63588 212 4 dout0[14]
rlabel metal4 s 65960 0 66036 212 4 dout0[15]
rlabel metal4 s 68272 0 68348 212 4 dout0[16]
rlabel metal4 s 16048 0 16124 212 4 addr0[0]
rlabel metal4 s 17136 0 17212 212 4 addr0[1]
rlabel metal4 s 18224 0 18300 212 4 wmask0[0]
rlabel metal4 s 19584 0 19660 212 4 wmask0[1]
rlabel metal4 s 20536 0 20612 212 4 wmask0[2]
rlabel metal4 s 21760 0 21836 212 4 wmask0[3]
rlabel metal4 s 23120 0 23196 212 4 din0[0]
rlabel metal4 s 24208 0 24284 212 4 din0[1]
rlabel metal4 s 25432 0 25508 212 4 din0[2]
rlabel metal4 s 26520 0 26596 212 4 din0[3]
rlabel metal4 s 27608 0 27684 212 4 din0[4]
rlabel metal4 s 28696 0 28772 212 4 din0[5]
rlabel metal4 s 30056 0 30132 212 4 din0[6]
rlabel metal4 s 31280 0 31356 212 4 din0[7]
rlabel metal4 s 32368 0 32444 212 4 din0[8]
rlabel metal4 s 33456 0 33532 212 4 din0[9]
rlabel metal4 s 34544 0 34620 212 4 din0[10]
rlabel metal4 s 35904 0 35980 212 4 din0[11]
rlabel metal4 s 36992 0 37068 212 4 din0[12]
rlabel metal4 s 38080 0 38156 212 4 din0[13]
rlabel metal4 s 39440 0 39516 212 4 din0[14]
rlabel metal4 s 40664 0 40740 212 4 din0[15]
rlabel metal4 s 41752 0 41828 212 4 din0[16]
rlabel metal4 s 42840 0 42916 212 4 din0[17]
rlabel metal4 s 43928 0 44004 212 4 din0[18]
rlabel metal4 s 45288 0 45364 212 4 din0[19]
rlabel metal4 s 46376 0 46452 212 4 din0[20]
rlabel metal4 s 47600 0 47676 212 4 din0[21]
rlabel metal4 s 48688 0 48764 212 4 din0[22]
rlabel metal4 s 49776 0 49852 212 4 din0[23]
rlabel metal4 s 51136 0 51212 212 4 din0[24]
rlabel metal4 s 52224 0 52300 212 4 din0[25]
rlabel metal4 s 53312 0 53388 212 4 din0[26]
rlabel metal4 s 54400 0 54476 212 4 din0[27]
rlabel metal4 s 55760 0 55836 212 4 din0[28]
rlabel metal4 s 56984 0 57060 212 4 din0[29]
rlabel metal4 s 58072 0 58148 212 4 din0[30]
rlabel metal4 s 59160 0 59236 212 4 din0[31]
rlabel metal4 s 28288 0 28364 212 4 dout0[0]
rlabel metal4 s 30736 0 30812 212 4 dout0[1]
rlabel metal4 s 33592 0 33668 212 4 dout0[2]
rlabel metal4 s 952 952 1300 82356 4 vccd1
rlabel metal4 s 272 272 620 83036 4 vssd1
rlabel metal4 s 103360 0 103436 212 4 dout0[30]
rlabel metal4 s 105944 0 106020 212 4 dout0[31]
rlabel metal4 s 70992 0 71068 212 4 dout0[17]
rlabel metal4 s 73440 0 73516 212 4 dout0[18]
rlabel metal4 s 75888 0 75964 212 4 dout0[19]
rlabel metal4 s 78472 0 78548 212 4 dout0[20]
rlabel metal4 s 80920 0 80996 212 4 dout0[21]
rlabel metal4 s 83504 0 83580 212 4 dout0[22]
rlabel metal4 s 85952 0 86028 212 4 dout0[23]
rlabel metal4 s 88536 0 88612 212 4 dout0[24]
rlabel metal4 s 90984 0 91060 212 4 dout0[25]
rlabel metal4 s 93432 0 93508 212 4 dout0[26]
rlabel metal4 s 95880 0 95956 212 4 dout0[27]
rlabel metal4 s 123216 0 123292 212 4 addr1[7]
rlabel metal4 s 123352 0 123428 212 4 addr1[8]
rlabel metal4 s 98464 0 98540 212 4 dout0[28]
rlabel metal4 s 135320 952 135668 82356 4 vccd1
rlabel metal4 s 136000 272 136348 83036 4 vssd1
rlabel metal4 s 100912 0 100988 212 4 dout0[29]
<< properties >>
string FIXED_BBOX 0 0 136620 83308
<< end >>
