magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< locali >>
rect 4094 100983 4122 101017
rect 70 100804 136 100838
rect 70 100612 136 100646
rect 4094 100433 4122 100467
rect 4094 100193 4122 100227
rect 70 100014 136 100048
rect 70 99822 136 99856
rect 4094 99643 4122 99677
rect 4094 99403 4122 99437
rect 70 99224 136 99258
rect 70 99032 136 99066
rect 4094 98853 4122 98887
rect 4094 98613 4122 98647
rect 70 98434 136 98468
rect 70 98242 136 98276
rect 4094 98063 4122 98097
rect 4094 97823 4122 97857
rect 70 97644 136 97678
rect 70 97452 136 97486
rect 4094 97273 4122 97307
rect 4094 97033 4122 97067
rect 70 96854 136 96888
rect 70 96662 136 96696
rect 4094 96483 4122 96517
rect 4094 96243 4122 96277
rect 70 96064 136 96098
rect 70 95872 136 95906
rect 4094 95693 4122 95727
rect 4094 95453 4122 95487
rect 70 95274 136 95308
rect 70 95082 136 95116
rect 4094 94903 4122 94937
rect 4094 94663 4122 94697
rect 70 94484 136 94518
rect 70 94292 136 94326
rect 4094 94113 4122 94147
rect 4094 93873 4122 93907
rect 70 93694 136 93728
rect 70 93502 136 93536
rect 4094 93323 4122 93357
rect 4094 93083 4122 93117
rect 70 92904 136 92938
rect 70 92712 136 92746
rect 4094 92533 4122 92567
rect 4094 92293 4122 92327
rect 70 92114 136 92148
rect 70 91922 136 91956
rect 4094 91743 4122 91777
rect 4094 91503 4122 91537
rect 70 91324 136 91358
rect 70 91132 136 91166
rect 4094 90953 4122 90987
rect 4094 90713 4122 90747
rect 70 90534 136 90568
rect 70 90342 136 90376
rect 4094 90163 4122 90197
rect 4094 89923 4122 89957
rect 70 89744 136 89778
rect 70 89552 136 89586
rect 4094 89373 4122 89407
rect 4094 89133 4122 89167
rect 70 88954 136 88988
rect 70 88762 136 88796
rect 4094 88583 4122 88617
rect 4094 88343 4122 88377
rect 70 88164 136 88198
rect 70 87972 136 88006
rect 4094 87793 4122 87827
rect 4094 87553 4122 87587
rect 70 87374 136 87408
rect 70 87182 136 87216
rect 4094 87003 4122 87037
rect 4094 86763 4122 86797
rect 70 86584 136 86618
rect 70 86392 136 86426
rect 4094 86213 4122 86247
rect 4094 85973 4122 86007
rect 70 85794 136 85828
rect 70 85602 136 85636
rect 4094 85423 4122 85457
rect 4094 85183 4122 85217
rect 70 85004 136 85038
rect 70 84812 136 84846
rect 4094 84633 4122 84667
rect 4094 84393 4122 84427
rect 70 84214 136 84248
rect 70 84022 136 84056
rect 4094 83843 4122 83877
rect 4094 83603 4122 83637
rect 70 83424 136 83458
rect 70 83232 136 83266
rect 4094 83053 4122 83087
rect 4094 82813 4122 82847
rect 70 82634 136 82668
rect 70 82442 136 82476
rect 4094 82263 4122 82297
rect 4094 82023 4122 82057
rect 70 81844 136 81878
rect 70 81652 136 81686
rect 4094 81473 4122 81507
rect 4094 81233 4122 81267
rect 70 81054 136 81088
rect 70 80862 136 80896
rect 4094 80683 4122 80717
rect 4094 80443 4122 80477
rect 70 80264 136 80298
rect 70 80072 136 80106
rect 4094 79893 4122 79927
rect 4094 79653 4122 79687
rect 70 79474 136 79508
rect 70 79282 136 79316
rect 4094 79103 4122 79137
rect 4094 78863 4122 78897
rect 70 78684 136 78718
rect 70 78492 136 78526
rect 4094 78313 4122 78347
rect 4094 78073 4122 78107
rect 70 77894 136 77928
rect 70 77702 136 77736
rect 4094 77523 4122 77557
rect 4094 77283 4122 77317
rect 70 77104 136 77138
rect 70 76912 136 76946
rect 4094 76733 4122 76767
rect 4094 76493 4122 76527
rect 70 76314 136 76348
rect 70 76122 136 76156
rect 4094 75943 4122 75977
rect 4094 75703 4122 75737
rect 70 75524 136 75558
rect 70 75332 136 75366
rect 4094 75153 4122 75187
rect 4094 74913 4122 74947
rect 70 74734 136 74768
rect 70 74542 136 74576
rect 4094 74363 4122 74397
rect 4094 74123 4122 74157
rect 70 73944 136 73978
rect 70 73752 136 73786
rect 4094 73573 4122 73607
rect 4094 73333 4122 73367
rect 70 73154 136 73188
rect 70 72962 136 72996
rect 4094 72783 4122 72817
rect 4094 72543 4122 72577
rect 70 72364 136 72398
rect 70 72172 136 72206
rect 4094 71993 4122 72027
rect 4094 71753 4122 71787
rect 70 71574 136 71608
rect 70 71382 136 71416
rect 4094 71203 4122 71237
rect 4094 70963 4122 70997
rect 70 70784 136 70818
rect 70 70592 136 70626
rect 4094 70413 4122 70447
rect 4094 70173 4122 70207
rect 70 69994 136 70028
rect 70 69802 136 69836
rect 4094 69623 4122 69657
rect 4094 69383 4122 69417
rect 70 69204 136 69238
rect 70 69012 136 69046
rect 4094 68833 4122 68867
rect 4094 68593 4122 68627
rect 70 68414 136 68448
rect 70 68222 136 68256
rect 4094 68043 4122 68077
rect 4094 67803 4122 67837
rect 70 67624 136 67658
rect 70 67432 136 67466
rect 4094 67253 4122 67287
rect 4094 67013 4122 67047
rect 70 66834 136 66868
rect 70 66642 136 66676
rect 4094 66463 4122 66497
rect 4094 66223 4122 66257
rect 70 66044 136 66078
rect 70 65852 136 65886
rect 4094 65673 4122 65707
rect 4094 65433 4122 65467
rect 70 65254 136 65288
rect 70 65062 136 65096
rect 4094 64883 4122 64917
rect 4094 64643 4122 64677
rect 70 64464 136 64498
rect 70 64272 136 64306
rect 4094 64093 4122 64127
rect 4094 63853 4122 63887
rect 70 63674 136 63708
rect 70 63482 136 63516
rect 4094 63303 4122 63337
rect 4094 63063 4122 63097
rect 70 62884 136 62918
rect 70 62692 136 62726
rect 4094 62513 4122 62547
rect 4094 62273 4122 62307
rect 70 62094 136 62128
rect 70 61902 136 61936
rect 4094 61723 4122 61757
rect 4094 61483 4122 61517
rect 70 61304 136 61338
rect 70 61112 136 61146
rect 4094 60933 4122 60967
rect 4094 60693 4122 60727
rect 70 60514 136 60548
rect 70 60322 136 60356
rect 4094 60143 4122 60177
rect 4094 59903 4122 59937
rect 70 59724 136 59758
rect 70 59532 136 59566
rect 4094 59353 4122 59387
rect 4094 59113 4122 59147
rect 70 58934 136 58968
rect 70 58742 136 58776
rect 4094 58563 4122 58597
rect 4094 58323 4122 58357
rect 70 58144 136 58178
rect 70 57952 136 57986
rect 4094 57773 4122 57807
rect 4094 57533 4122 57567
rect 70 57354 136 57388
rect 70 57162 136 57196
rect 4094 56983 4122 57017
rect 4094 56743 4122 56777
rect 70 56564 136 56598
rect 70 56372 136 56406
rect 4094 56193 4122 56227
rect 4094 55953 4122 55987
rect 70 55774 136 55808
rect 70 55582 136 55616
rect 4094 55403 4122 55437
rect 4094 55163 4122 55197
rect 70 54984 136 55018
rect 70 54792 136 54826
rect 4094 54613 4122 54647
rect 4094 54373 4122 54407
rect 70 54194 136 54228
rect 70 54002 136 54036
rect 4094 53823 4122 53857
rect 4094 53583 4122 53617
rect 70 53404 136 53438
rect 70 53212 136 53246
rect 4094 53033 4122 53067
rect 4094 52793 4122 52827
rect 70 52614 136 52648
rect 70 52422 136 52456
rect 4094 52243 4122 52277
rect 4094 52003 4122 52037
rect 70 51824 136 51858
rect 70 51632 136 51666
rect 4094 51453 4122 51487
rect 4094 51213 4122 51247
rect 70 51034 136 51068
rect 70 50842 136 50876
rect 4094 50663 4122 50697
rect 4094 50423 4122 50457
rect 70 50244 136 50278
rect 70 50052 136 50086
rect 4094 49873 4122 49907
rect 4094 49633 4122 49667
rect 70 49454 136 49488
rect 70 49262 136 49296
rect 4094 49083 4122 49117
rect 4094 48843 4122 48877
rect 70 48664 136 48698
rect 70 48472 136 48506
rect 4094 48293 4122 48327
rect 4094 48053 4122 48087
rect 70 47874 136 47908
rect 70 47682 136 47716
rect 4094 47503 4122 47537
rect 4094 47263 4122 47297
rect 70 47084 136 47118
rect 70 46892 136 46926
rect 4094 46713 4122 46747
rect 4094 46473 4122 46507
rect 70 46294 136 46328
rect 70 46102 136 46136
rect 4094 45923 4122 45957
rect 4094 45683 4122 45717
rect 70 45504 136 45538
rect 70 45312 136 45346
rect 4094 45133 4122 45167
rect 4094 44893 4122 44927
rect 70 44714 136 44748
rect 70 44522 136 44556
rect 4094 44343 4122 44377
rect 4094 44103 4122 44137
rect 70 43924 136 43958
rect 70 43732 136 43766
rect 4094 43553 4122 43587
rect 4094 43313 4122 43347
rect 70 43134 136 43168
rect 70 42942 136 42976
rect 4094 42763 4122 42797
rect 4094 42523 4122 42557
rect 70 42344 136 42378
rect 70 42152 136 42186
rect 4094 41973 4122 42007
rect 4094 41733 4122 41767
rect 70 41554 136 41588
rect 70 41362 136 41396
rect 4094 41183 4122 41217
rect 4094 40943 4122 40977
rect 70 40764 136 40798
rect 70 40572 136 40606
rect 4094 40393 4122 40427
rect 4094 40153 4122 40187
rect 70 39974 136 40008
rect 70 39782 136 39816
rect 4094 39603 4122 39637
rect 4094 39363 4122 39397
rect 70 39184 136 39218
rect 70 38992 136 39026
rect 4094 38813 4122 38847
rect 4094 38573 4122 38607
rect 70 38394 136 38428
rect 70 38202 136 38236
rect 4094 38023 4122 38057
rect 4094 37783 4122 37817
rect 70 37604 136 37638
rect 70 37412 136 37446
rect 4094 37233 4122 37267
rect 4094 36993 4122 37027
rect 70 36814 136 36848
rect 70 36622 136 36656
rect 4094 36443 4122 36477
rect 4094 36203 4122 36237
rect 70 36024 136 36058
rect 70 35832 136 35866
rect 4094 35653 4122 35687
rect 4094 35413 4122 35447
rect 70 35234 136 35268
rect 70 35042 136 35076
rect 4094 34863 4122 34897
rect 4094 34623 4122 34657
rect 70 34444 136 34478
rect 70 34252 136 34286
rect 4094 34073 4122 34107
rect 4094 33833 4122 33867
rect 70 33654 136 33688
rect 70 33462 136 33496
rect 4094 33283 4122 33317
rect 4094 33043 4122 33077
rect 70 32864 136 32898
rect 70 32672 136 32706
rect 4094 32493 4122 32527
rect 4094 32253 4122 32287
rect 70 32074 136 32108
rect 70 31882 136 31916
rect 4094 31703 4122 31737
rect 4094 31463 4122 31497
rect 70 31284 136 31318
rect 70 31092 136 31126
rect 4094 30913 4122 30947
rect 4094 30673 4122 30707
rect 70 30494 136 30528
rect 70 30302 136 30336
rect 4094 30123 4122 30157
rect 4094 29883 4122 29917
rect 70 29704 136 29738
rect 70 29512 136 29546
rect 4094 29333 4122 29367
rect 4094 29093 4122 29127
rect 70 28914 136 28948
rect 70 28722 136 28756
rect 4094 28543 4122 28577
rect 4094 28303 4122 28337
rect 70 28124 136 28158
rect 70 27932 136 27966
rect 4094 27753 4122 27787
rect 4094 27513 4122 27547
rect 70 27334 136 27368
rect 70 27142 136 27176
rect 4094 26963 4122 26997
rect 4094 26723 4122 26757
rect 70 26544 136 26578
rect 70 26352 136 26386
rect 4094 26173 4122 26207
rect 4094 25933 4122 25967
rect 70 25754 136 25788
rect 70 25562 136 25596
rect 4094 25383 4122 25417
rect 4094 25143 4122 25177
rect 70 24964 136 24998
rect 70 24772 136 24806
rect 4094 24593 4122 24627
rect 4094 24353 4122 24387
rect 70 24174 136 24208
rect 70 23982 136 24016
rect 4094 23803 4122 23837
rect 4094 23563 4122 23597
rect 70 23384 136 23418
rect 70 23192 136 23226
rect 4094 23013 4122 23047
rect 4094 22773 4122 22807
rect 70 22594 136 22628
rect 70 22402 136 22436
rect 4094 22223 4122 22257
rect 4094 21983 4122 22017
rect 70 21804 136 21838
rect 70 21612 136 21646
rect 4094 21433 4122 21467
rect 4094 21193 4122 21227
rect 70 21014 136 21048
rect 70 20822 136 20856
rect 4094 20643 4122 20677
rect 4094 20403 4122 20437
rect 70 20224 136 20258
rect 70 20032 136 20066
rect 4094 19853 4122 19887
rect 4094 19613 4122 19647
rect 70 19434 136 19468
rect 70 19242 136 19276
rect 4094 19063 4122 19097
rect 4094 18823 4122 18857
rect 70 18644 136 18678
rect 70 18452 136 18486
rect 4094 18273 4122 18307
rect 4094 18033 4122 18067
rect 70 17854 136 17888
rect 70 17662 136 17696
rect 4094 17483 4122 17517
rect 4094 17243 4122 17277
rect 70 17064 136 17098
rect 70 16872 136 16906
rect 4094 16693 4122 16727
rect 4094 16453 4122 16487
rect 70 16274 136 16308
rect 70 16082 136 16116
rect 4094 15903 4122 15937
rect 4094 15663 4122 15697
rect 70 15484 136 15518
rect 70 15292 136 15326
rect 4094 15113 4122 15147
rect 4094 14873 4122 14907
rect 70 14694 136 14728
rect 70 14502 136 14536
rect 4094 14323 4122 14357
rect 4094 14083 4122 14117
rect 70 13904 136 13938
rect 70 13712 136 13746
rect 4094 13533 4122 13567
rect 4094 13293 4122 13327
rect 70 13114 136 13148
rect 70 12922 136 12956
rect 4094 12743 4122 12777
rect 4094 12503 4122 12537
rect 70 12324 136 12358
rect 70 12132 136 12166
rect 4094 11953 4122 11987
rect 4094 11713 4122 11747
rect 70 11534 136 11568
rect 70 11342 136 11376
rect 4094 11163 4122 11197
rect 4094 10923 4122 10957
rect 70 10744 136 10778
rect 70 10552 136 10586
rect 4094 10373 4122 10407
rect 4094 10133 4122 10167
rect 70 9954 136 9988
rect 70 9762 136 9796
rect 4094 9583 4122 9617
rect 4094 9343 4122 9377
rect 70 9164 136 9198
rect 70 8972 136 9006
rect 4094 8793 4122 8827
rect 4094 8553 4122 8587
rect 70 8374 136 8408
rect 70 8182 136 8216
rect 4094 8003 4122 8037
rect 4094 7763 4122 7797
rect 70 7584 136 7618
rect 70 7392 136 7426
rect 4094 7213 4122 7247
rect 4094 6973 4122 7007
rect 70 6794 136 6828
rect 70 6602 136 6636
rect 4094 6423 4122 6457
rect 4094 6183 4122 6217
rect 70 6004 136 6038
rect 70 5812 136 5846
rect 4094 5633 4122 5667
rect 4094 5393 4122 5427
rect 70 5214 136 5248
rect 70 5022 136 5056
rect 4094 4843 4122 4877
rect 4094 4603 4122 4637
rect 70 4424 136 4458
rect 70 4232 136 4266
rect 4094 4053 4122 4087
rect 4094 3813 4122 3847
rect 70 3634 136 3668
rect 70 3442 136 3476
rect 4094 3263 4122 3297
rect 4094 3023 4122 3057
rect 70 2844 136 2878
rect 70 2652 136 2686
rect 4094 2473 4122 2507
rect 4094 2233 4122 2267
rect 70 2054 136 2088
rect 70 1862 136 1896
rect 4094 1683 4122 1717
rect 4094 1443 4122 1477
rect 70 1264 136 1298
rect 70 1072 136 1106
rect 4094 893 4122 927
rect 4094 653 4122 687
rect 70 474 136 508
rect 70 282 136 316
rect 4094 103 4122 137
<< metal1 >>
rect 71 100903 135 100955
rect 71 100495 135 100547
rect 71 100113 135 100165
rect 71 99705 135 99757
rect 71 99323 135 99375
rect 71 98915 135 98967
rect 71 98533 135 98585
rect 71 98125 135 98177
rect 71 97743 135 97795
rect 71 97335 135 97387
rect 71 96953 135 97005
rect 71 96545 135 96597
rect 71 96163 135 96215
rect 71 95755 135 95807
rect 71 95373 135 95425
rect 71 94965 135 95017
rect 71 94583 135 94635
rect 71 94175 135 94227
rect 71 93793 135 93845
rect 71 93385 135 93437
rect 71 93003 135 93055
rect 71 92595 135 92647
rect 71 92213 135 92265
rect 71 91805 135 91857
rect 71 91423 135 91475
rect 71 91015 135 91067
rect 71 90633 135 90685
rect 71 90225 135 90277
rect 71 89843 135 89895
rect 71 89435 135 89487
rect 71 89053 135 89105
rect 71 88645 135 88697
rect 71 88263 135 88315
rect 71 87855 135 87907
rect 71 87473 135 87525
rect 71 87065 135 87117
rect 71 86683 135 86735
rect 71 86275 135 86327
rect 71 85893 135 85945
rect 71 85485 135 85537
rect 71 85103 135 85155
rect 71 84695 135 84747
rect 71 84313 135 84365
rect 71 83905 135 83957
rect 71 83523 135 83575
rect 71 83115 135 83167
rect 71 82733 135 82785
rect 71 82325 135 82377
rect 71 81943 135 81995
rect 71 81535 135 81587
rect 71 81153 135 81205
rect 71 80745 135 80797
rect 71 80363 135 80415
rect 71 79955 135 80007
rect 71 79573 135 79625
rect 71 79165 135 79217
rect 71 78783 135 78835
rect 71 78375 135 78427
rect 71 77993 135 78045
rect 71 77585 135 77637
rect 71 77203 135 77255
rect 71 76795 135 76847
rect 71 76413 135 76465
rect 71 76005 135 76057
rect 71 75623 135 75675
rect 71 75215 135 75267
rect 71 74833 135 74885
rect 71 74425 135 74477
rect 71 74043 135 74095
rect 71 73635 135 73687
rect 71 73253 135 73305
rect 71 72845 135 72897
rect 71 72463 135 72515
rect 71 72055 135 72107
rect 71 71673 135 71725
rect 71 71265 135 71317
rect 71 70883 135 70935
rect 71 70475 135 70527
rect 71 70093 135 70145
rect 71 69685 135 69737
rect 71 69303 135 69355
rect 71 68895 135 68947
rect 71 68513 135 68565
rect 71 68105 135 68157
rect 71 67723 135 67775
rect 71 67315 135 67367
rect 71 66933 135 66985
rect 71 66525 135 66577
rect 71 66143 135 66195
rect 71 65735 135 65787
rect 71 65353 135 65405
rect 71 64945 135 64997
rect 71 64563 135 64615
rect 71 64155 135 64207
rect 71 63773 135 63825
rect 71 63365 135 63417
rect 71 62983 135 63035
rect 71 62575 135 62627
rect 71 62193 135 62245
rect 71 61785 135 61837
rect 71 61403 135 61455
rect 71 60995 135 61047
rect 71 60613 135 60665
rect 71 60205 135 60257
rect 71 59823 135 59875
rect 71 59415 135 59467
rect 71 59033 135 59085
rect 71 58625 135 58677
rect 71 58243 135 58295
rect 71 57835 135 57887
rect 71 57453 135 57505
rect 71 57045 135 57097
rect 71 56663 135 56715
rect 71 56255 135 56307
rect 71 55873 135 55925
rect 71 55465 135 55517
rect 71 55083 135 55135
rect 71 54675 135 54727
rect 71 54293 135 54345
rect 71 53885 135 53937
rect 71 53503 135 53555
rect 71 53095 135 53147
rect 71 52713 135 52765
rect 71 52305 135 52357
rect 71 51923 135 51975
rect 71 51515 135 51567
rect 71 51133 135 51185
rect 71 50725 135 50777
rect 71 50343 135 50395
rect 71 49935 135 49987
rect 71 49553 135 49605
rect 71 49145 135 49197
rect 71 48763 135 48815
rect 71 48355 135 48407
rect 71 47973 135 48025
rect 71 47565 135 47617
rect 71 47183 135 47235
rect 71 46775 135 46827
rect 71 46393 135 46445
rect 71 45985 135 46037
rect 71 45603 135 45655
rect 71 45195 135 45247
rect 71 44813 135 44865
rect 71 44405 135 44457
rect 71 44023 135 44075
rect 71 43615 135 43667
rect 71 43233 135 43285
rect 71 42825 135 42877
rect 71 42443 135 42495
rect 71 42035 135 42087
rect 71 41653 135 41705
rect 71 41245 135 41297
rect 71 40863 135 40915
rect 71 40455 135 40507
rect 71 40073 135 40125
rect 71 39665 135 39717
rect 71 39283 135 39335
rect 71 38875 135 38927
rect 71 38493 135 38545
rect 71 38085 135 38137
rect 71 37703 135 37755
rect 71 37295 135 37347
rect 71 36913 135 36965
rect 71 36505 135 36557
rect 71 36123 135 36175
rect 71 35715 135 35767
rect 71 35333 135 35385
rect 71 34925 135 34977
rect 71 34543 135 34595
rect 71 34135 135 34187
rect 71 33753 135 33805
rect 71 33345 135 33397
rect 71 32963 135 33015
rect 71 32555 135 32607
rect 71 32173 135 32225
rect 71 31765 135 31817
rect 71 31383 135 31435
rect 71 30975 135 31027
rect 71 30593 135 30645
rect 71 30185 135 30237
rect 71 29803 135 29855
rect 71 29395 135 29447
rect 71 29013 135 29065
rect 71 28605 135 28657
rect 71 28223 135 28275
rect 71 27815 135 27867
rect 71 27433 135 27485
rect 71 27025 135 27077
rect 71 26643 135 26695
rect 71 26235 135 26287
rect 71 25853 135 25905
rect 71 25445 135 25497
rect 71 25063 135 25115
rect 71 24655 135 24707
rect 71 24273 135 24325
rect 71 23865 135 23917
rect 71 23483 135 23535
rect 71 23075 135 23127
rect 71 22693 135 22745
rect 71 22285 135 22337
rect 71 21903 135 21955
rect 71 21495 135 21547
rect 71 21113 135 21165
rect 71 20705 135 20757
rect 71 20323 135 20375
rect 71 19915 135 19967
rect 71 19533 135 19585
rect 71 19125 135 19177
rect 71 18743 135 18795
rect 71 18335 135 18387
rect 71 17953 135 18005
rect 71 17545 135 17597
rect 71 17163 135 17215
rect 71 16755 135 16807
rect 71 16373 135 16425
rect 71 15965 135 16017
rect 71 15583 135 15635
rect 71 15175 135 15227
rect 71 14793 135 14845
rect 71 14385 135 14437
rect 71 14003 135 14055
rect 71 13595 135 13647
rect 71 13213 135 13265
rect 71 12805 135 12857
rect 71 12423 135 12475
rect 71 12015 135 12067
rect 71 11633 135 11685
rect 71 11225 135 11277
rect 71 10843 135 10895
rect 71 10435 135 10487
rect 71 10053 135 10105
rect 71 9645 135 9697
rect 71 9263 135 9315
rect 71 8855 135 8907
rect 71 8473 135 8525
rect 71 8065 135 8117
rect 71 7683 135 7735
rect 71 7275 135 7327
rect 71 6893 135 6945
rect 71 6485 135 6537
rect 71 6103 135 6155
rect 71 5695 135 5747
rect 71 5313 135 5365
rect 71 4905 135 4957
rect 71 4523 135 4575
rect 71 4115 135 4167
rect 71 3733 135 3785
rect 71 3325 135 3377
rect 71 2943 135 2995
rect 71 2535 135 2587
rect 71 2153 135 2205
rect 71 1745 135 1797
rect 71 1363 135 1415
rect 71 955 135 1007
rect 71 573 135 625
rect 71 165 135 217
rect 256 -30 284 101120
rect 681 -32 709 101120
rect 1724 0 1752 101120
rect 3372 0 3400 101120
<< metal2 >>
rect 70 0 98 101120
use contact_7  contact_7_255
timestamp 1624494425
transform 1 0 74 0 1 158
box 0 0 58 66
use contact_8  contact_8_255
timestamp 1624494425
transform 1 0 71 0 1 159
box 0 0 64 64
use wordline_driver  wordline_driver_254
timestamp 1624494425
transform 1 0 0 0 -1 790
box 70 -56 4140 490
use wordline_driver  wordline_driver_255
timestamp 1624494425
transform 1 0 0 0 1 0
box 70 -56 4140 490
use contact_7  contact_7_254
timestamp 1624494425
transform 1 0 74 0 1 566
box 0 0 58 66
use contact_8  contact_8_254
timestamp 1624494425
transform 1 0 71 0 1 567
box 0 0 64 64
use contact_7  contact_7_253
timestamp 1624494425
transform 1 0 74 0 1 948
box 0 0 58 66
use contact_8  contact_8_253
timestamp 1624494425
transform 1 0 71 0 1 949
box 0 0 64 64
use wordline_driver  wordline_driver_253
timestamp 1624494425
transform 1 0 0 0 1 790
box 70 -56 4140 490
use contact_7  contact_7_252
timestamp 1624494425
transform 1 0 74 0 1 1356
box 0 0 58 66
use contact_8  contact_8_252
timestamp 1624494425
transform 1 0 71 0 1 1357
box 0 0 64 64
use wordline_driver  wordline_driver_251
timestamp 1624494425
transform 1 0 0 0 1 1580
box 70 -56 4140 490
use wordline_driver  wordline_driver_252
timestamp 1624494425
transform 1 0 0 0 -1 1580
box 70 -56 4140 490
use contact_7  contact_7_251
timestamp 1624494425
transform 1 0 74 0 1 1738
box 0 0 58 66
use contact_8  contact_8_251
timestamp 1624494425
transform 1 0 71 0 1 1739
box 0 0 64 64
use wordline_driver  wordline_driver_250
timestamp 1624494425
transform 1 0 0 0 -1 2370
box 70 -56 4140 490
use contact_7  contact_7_250
timestamp 1624494425
transform 1 0 74 0 1 2146
box 0 0 58 66
use contact_8  contact_8_250
timestamp 1624494425
transform 1 0 71 0 1 2147
box 0 0 64 64
use contact_7  contact_7_249
timestamp 1624494425
transform 1 0 74 0 1 2528
box 0 0 58 66
use contact_8  contact_8_249
timestamp 1624494425
transform 1 0 71 0 1 2529
box 0 0 64 64
use wordline_driver  wordline_driver_248
timestamp 1624494425
transform 1 0 0 0 -1 3160
box 70 -56 4140 490
use wordline_driver  wordline_driver_249
timestamp 1624494425
transform 1 0 0 0 1 2370
box 70 -56 4140 490
use contact_7  contact_7_248
timestamp 1624494425
transform 1 0 74 0 1 2936
box 0 0 58 66
use contact_8  contact_8_248
timestamp 1624494425
transform 1 0 71 0 1 2937
box 0 0 64 64
use wordline_driver  wordline_driver_247
timestamp 1624494425
transform 1 0 0 0 1 3160
box 70 -56 4140 490
use contact_7  contact_7_247
timestamp 1624494425
transform 1 0 74 0 1 3318
box 0 0 58 66
use contact_8  contact_8_247
timestamp 1624494425
transform 1 0 71 0 1 3319
box 0 0 64 64
use contact_7  contact_7_246
timestamp 1624494425
transform 1 0 74 0 1 3726
box 0 0 58 66
use contact_8  contact_8_246
timestamp 1624494425
transform 1 0 71 0 1 3727
box 0 0 64 64
use wordline_driver  wordline_driver_246
timestamp 1624494425
transform 1 0 0 0 -1 3950
box 70 -56 4140 490
use contact_7  contact_7_245
timestamp 1624494425
transform 1 0 74 0 1 4108
box 0 0 58 66
use contact_8  contact_8_245
timestamp 1624494425
transform 1 0 71 0 1 4109
box 0 0 64 64
use wordline_driver  wordline_driver_244
timestamp 1624494425
transform 1 0 0 0 -1 4740
box 70 -56 4140 490
use wordline_driver  wordline_driver_245
timestamp 1624494425
transform 1 0 0 0 1 3950
box 70 -56 4140 490
use contact_7  contact_7_244
timestamp 1624494425
transform 1 0 74 0 1 4516
box 0 0 58 66
use contact_8  contact_8_244
timestamp 1624494425
transform 1 0 71 0 1 4517
box 0 0 64 64
use wordline_driver  wordline_driver_243
timestamp 1624494425
transform 1 0 0 0 1 4740
box 70 -56 4140 490
use contact_7  contact_7_243
timestamp 1624494425
transform 1 0 74 0 1 4898
box 0 0 58 66
use contact_8  contact_8_243
timestamp 1624494425
transform 1 0 71 0 1 4899
box 0 0 64 64
use contact_7  contact_7_242
timestamp 1624494425
transform 1 0 74 0 1 5306
box 0 0 58 66
use contact_8  contact_8_242
timestamp 1624494425
transform 1 0 71 0 1 5307
box 0 0 64 64
use wordline_driver  wordline_driver_242
timestamp 1624494425
transform 1 0 0 0 -1 5530
box 70 -56 4140 490
use contact_7  contact_7_241
timestamp 1624494425
transform 1 0 74 0 1 5688
box 0 0 58 66
use contact_8  contact_8_241
timestamp 1624494425
transform 1 0 71 0 1 5689
box 0 0 64 64
use wordline_driver  wordline_driver_240
timestamp 1624494425
transform 1 0 0 0 -1 6320
box 70 -56 4140 490
use wordline_driver  wordline_driver_241
timestamp 1624494425
transform 1 0 0 0 1 5530
box 70 -56 4140 490
use contact_7  contact_7_240
timestamp 1624494425
transform 1 0 74 0 1 6096
box 0 0 58 66
use contact_8  contact_8_240
timestamp 1624494425
transform 1 0 71 0 1 6097
box 0 0 64 64
use contact_7  contact_7_239
timestamp 1624494425
transform 1 0 74 0 1 6478
box 0 0 58 66
use contact_8  contact_8_239
timestamp 1624494425
transform 1 0 71 0 1 6479
box 0 0 64 64
use wordline_driver  wordline_driver_239
timestamp 1624494425
transform 1 0 0 0 1 6320
box 70 -56 4140 490
use contact_7  contact_7_238
timestamp 1624494425
transform 1 0 74 0 1 6886
box 0 0 58 66
use contact_8  contact_8_238
timestamp 1624494425
transform 1 0 71 0 1 6887
box 0 0 64 64
use wordline_driver  wordline_driver_237
timestamp 1624494425
transform 1 0 0 0 1 7110
box 70 -56 4140 490
use wordline_driver  wordline_driver_238
timestamp 1624494425
transform 1 0 0 0 -1 7110
box 70 -56 4140 490
use contact_7  contact_7_237
timestamp 1624494425
transform 1 0 74 0 1 7268
box 0 0 58 66
use contact_8  contact_8_237
timestamp 1624494425
transform 1 0 71 0 1 7269
box 0 0 64 64
use wordline_driver  wordline_driver_236
timestamp 1624494425
transform 1 0 0 0 -1 7900
box 70 -56 4140 490
use contact_7  contact_7_236
timestamp 1624494425
transform 1 0 74 0 1 7676
box 0 0 58 66
use contact_8  contact_8_236
timestamp 1624494425
transform 1 0 71 0 1 7677
box 0 0 64 64
use contact_7  contact_7_235
timestamp 1624494425
transform 1 0 74 0 1 8058
box 0 0 58 66
use contact_8  contact_8_235
timestamp 1624494425
transform 1 0 71 0 1 8059
box 0 0 64 64
use wordline_driver  wordline_driver_235
timestamp 1624494425
transform 1 0 0 0 1 7900
box 70 -56 4140 490
use contact_7  contact_7_234
timestamp 1624494425
transform 1 0 74 0 1 8466
box 0 0 58 66
use contact_8  contact_8_234
timestamp 1624494425
transform 1 0 71 0 1 8467
box 0 0 64 64
use wordline_driver  wordline_driver_233
timestamp 1624494425
transform 1 0 0 0 1 8690
box 70 -56 4140 490
use wordline_driver  wordline_driver_234
timestamp 1624494425
transform 1 0 0 0 -1 8690
box 70 -56 4140 490
use contact_7  contact_7_233
timestamp 1624494425
transform 1 0 74 0 1 8848
box 0 0 58 66
use contact_8  contact_8_233
timestamp 1624494425
transform 1 0 71 0 1 8849
box 0 0 64 64
use wordline_driver  wordline_driver_232
timestamp 1624494425
transform 1 0 0 0 -1 9480
box 70 -56 4140 490
use contact_7  contact_7_232
timestamp 1624494425
transform 1 0 74 0 1 9256
box 0 0 58 66
use contact_8  contact_8_232
timestamp 1624494425
transform 1 0 71 0 1 9257
box 0 0 64 64
use contact_7  contact_7_231
timestamp 1624494425
transform 1 0 74 0 1 9638
box 0 0 58 66
use contact_8  contact_8_231
timestamp 1624494425
transform 1 0 71 0 1 9639
box 0 0 64 64
use wordline_driver  wordline_driver_230
timestamp 1624494425
transform 1 0 0 0 -1 10270
box 70 -56 4140 490
use wordline_driver  wordline_driver_231
timestamp 1624494425
transform 1 0 0 0 1 9480
box 70 -56 4140 490
use contact_7  contact_7_230
timestamp 1624494425
transform 1 0 74 0 1 10046
box 0 0 58 66
use contact_8  contact_8_230
timestamp 1624494425
transform 1 0 71 0 1 10047
box 0 0 64 64
use wordline_driver  wordline_driver_229
timestamp 1624494425
transform 1 0 0 0 1 10270
box 70 -56 4140 490
use contact_7  contact_7_229
timestamp 1624494425
transform 1 0 74 0 1 10428
box 0 0 58 66
use contact_8  contact_8_229
timestamp 1624494425
transform 1 0 71 0 1 10429
box 0 0 64 64
use contact_7  contact_7_228
timestamp 1624494425
transform 1 0 74 0 1 10836
box 0 0 58 66
use contact_8  contact_8_228
timestamp 1624494425
transform 1 0 71 0 1 10837
box 0 0 64 64
use wordline_driver  wordline_driver_228
timestamp 1624494425
transform 1 0 0 0 -1 11060
box 70 -56 4140 490
use contact_7  contact_7_227
timestamp 1624494425
transform 1 0 74 0 1 11218
box 0 0 58 66
use contact_8  contact_8_227
timestamp 1624494425
transform 1 0 71 0 1 11219
box 0 0 64 64
use wordline_driver  wordline_driver_226
timestamp 1624494425
transform 1 0 0 0 -1 11850
box 70 -56 4140 490
use wordline_driver  wordline_driver_227
timestamp 1624494425
transform 1 0 0 0 1 11060
box 70 -56 4140 490
use contact_7  contact_7_226
timestamp 1624494425
transform 1 0 74 0 1 11626
box 0 0 58 66
use contact_8  contact_8_226
timestamp 1624494425
transform 1 0 71 0 1 11627
box 0 0 64 64
use wordline_driver  wordline_driver_225
timestamp 1624494425
transform 1 0 0 0 1 11850
box 70 -56 4140 490
use contact_7  contact_7_225
timestamp 1624494425
transform 1 0 74 0 1 12008
box 0 0 58 66
use contact_8  contact_8_225
timestamp 1624494425
transform 1 0 71 0 1 12009
box 0 0 64 64
use contact_7  contact_7_224
timestamp 1624494425
transform 1 0 74 0 1 12416
box 0 0 58 66
use contact_8  contact_8_224
timestamp 1624494425
transform 1 0 71 0 1 12417
box 0 0 64 64
use wordline_driver  wordline_driver_224
timestamp 1624494425
transform 1 0 0 0 -1 12640
box 70 -56 4140 490
use contact_7  contact_7_223
timestamp 1624494425
transform 1 0 74 0 1 12798
box 0 0 58 66
use contact_8  contact_8_223
timestamp 1624494425
transform 1 0 71 0 1 12799
box 0 0 64 64
use wordline_driver  wordline_driver_222
timestamp 1624494425
transform 1 0 0 0 -1 13430
box 70 -56 4140 490
use wordline_driver  wordline_driver_223
timestamp 1624494425
transform 1 0 0 0 1 12640
box 70 -56 4140 490
use contact_7  contact_7_222
timestamp 1624494425
transform 1 0 74 0 1 13206
box 0 0 58 66
use contact_8  contact_8_222
timestamp 1624494425
transform 1 0 71 0 1 13207
box 0 0 64 64
use contact_7  contact_7_221
timestamp 1624494425
transform 1 0 74 0 1 13588
box 0 0 58 66
use contact_8  contact_8_221
timestamp 1624494425
transform 1 0 71 0 1 13589
box 0 0 64 64
use wordline_driver  wordline_driver_221
timestamp 1624494425
transform 1 0 0 0 1 13430
box 70 -56 4140 490
use contact_7  contact_7_220
timestamp 1624494425
transform 1 0 74 0 1 13996
box 0 0 58 66
use contact_8  contact_8_220
timestamp 1624494425
transform 1 0 71 0 1 13997
box 0 0 64 64
use wordline_driver  wordline_driver_219
timestamp 1624494425
transform 1 0 0 0 1 14220
box 70 -56 4140 490
use wordline_driver  wordline_driver_220
timestamp 1624494425
transform 1 0 0 0 -1 14220
box 70 -56 4140 490
use contact_7  contact_7_219
timestamp 1624494425
transform 1 0 74 0 1 14378
box 0 0 58 66
use contact_8  contact_8_219
timestamp 1624494425
transform 1 0 71 0 1 14379
box 0 0 64 64
use wordline_driver  wordline_driver_218
timestamp 1624494425
transform 1 0 0 0 -1 15010
box 70 -56 4140 490
use contact_7  contact_7_218
timestamp 1624494425
transform 1 0 74 0 1 14786
box 0 0 58 66
use contact_8  contact_8_218
timestamp 1624494425
transform 1 0 71 0 1 14787
box 0 0 64 64
use contact_7  contact_7_217
timestamp 1624494425
transform 1 0 74 0 1 15168
box 0 0 58 66
use contact_8  contact_8_217
timestamp 1624494425
transform 1 0 71 0 1 15169
box 0 0 64 64
use wordline_driver  wordline_driver_217
timestamp 1624494425
transform 1 0 0 0 1 15010
box 70 -56 4140 490
use contact_7  contact_7_216
timestamp 1624494425
transform 1 0 74 0 1 15576
box 0 0 58 66
use contact_8  contact_8_216
timestamp 1624494425
transform 1 0 71 0 1 15577
box 0 0 64 64
use wordline_driver  wordline_driver_215
timestamp 1624494425
transform 1 0 0 0 1 15800
box 70 -56 4140 490
use wordline_driver  wordline_driver_216
timestamp 1624494425
transform 1 0 0 0 -1 15800
box 70 -56 4140 490
use contact_7  contact_7_215
timestamp 1624494425
transform 1 0 74 0 1 15958
box 0 0 58 66
use contact_8  contact_8_215
timestamp 1624494425
transform 1 0 71 0 1 15959
box 0 0 64 64
use wordline_driver  wordline_driver_214
timestamp 1624494425
transform 1 0 0 0 -1 16590
box 70 -56 4140 490
use contact_7  contact_7_214
timestamp 1624494425
transform 1 0 74 0 1 16366
box 0 0 58 66
use contact_8  contact_8_214
timestamp 1624494425
transform 1 0 71 0 1 16367
box 0 0 64 64
use contact_7  contact_7_213
timestamp 1624494425
transform 1 0 74 0 1 16748
box 0 0 58 66
use contact_8  contact_8_213
timestamp 1624494425
transform 1 0 71 0 1 16749
box 0 0 64 64
use wordline_driver  wordline_driver_212
timestamp 1624494425
transform 1 0 0 0 -1 17380
box 70 -56 4140 490
use wordline_driver  wordline_driver_213
timestamp 1624494425
transform 1 0 0 0 1 16590
box 70 -56 4140 490
use contact_7  contact_7_212
timestamp 1624494425
transform 1 0 74 0 1 17156
box 0 0 58 66
use contact_8  contact_8_212
timestamp 1624494425
transform 1 0 71 0 1 17157
box 0 0 64 64
use wordline_driver  wordline_driver_211
timestamp 1624494425
transform 1 0 0 0 1 17380
box 70 -56 4140 490
use contact_7  contact_7_211
timestamp 1624494425
transform 1 0 74 0 1 17538
box 0 0 58 66
use contact_8  contact_8_211
timestamp 1624494425
transform 1 0 71 0 1 17539
box 0 0 64 64
use contact_7  contact_7_210
timestamp 1624494425
transform 1 0 74 0 1 17946
box 0 0 58 66
use contact_8  contact_8_210
timestamp 1624494425
transform 1 0 71 0 1 17947
box 0 0 64 64
use wordline_driver  wordline_driver_210
timestamp 1624494425
transform 1 0 0 0 -1 18170
box 70 -56 4140 490
use contact_7  contact_7_209
timestamp 1624494425
transform 1 0 74 0 1 18328
box 0 0 58 66
use contact_8  contact_8_209
timestamp 1624494425
transform 1 0 71 0 1 18329
box 0 0 64 64
use wordline_driver  wordline_driver_208
timestamp 1624494425
transform 1 0 0 0 -1 18960
box 70 -56 4140 490
use wordline_driver  wordline_driver_209
timestamp 1624494425
transform 1 0 0 0 1 18170
box 70 -56 4140 490
use contact_7  contact_7_208
timestamp 1624494425
transform 1 0 74 0 1 18736
box 0 0 58 66
use contact_8  contact_8_208
timestamp 1624494425
transform 1 0 71 0 1 18737
box 0 0 64 64
use wordline_driver  wordline_driver_207
timestamp 1624494425
transform 1 0 0 0 1 18960
box 70 -56 4140 490
use contact_7  contact_7_207
timestamp 1624494425
transform 1 0 74 0 1 19118
box 0 0 58 66
use contact_8  contact_8_207
timestamp 1624494425
transform 1 0 71 0 1 19119
box 0 0 64 64
use contact_7  contact_7_206
timestamp 1624494425
transform 1 0 74 0 1 19526
box 0 0 58 66
use contact_8  contact_8_206
timestamp 1624494425
transform 1 0 71 0 1 19527
box 0 0 64 64
use wordline_driver  wordline_driver_206
timestamp 1624494425
transform 1 0 0 0 -1 19750
box 70 -56 4140 490
use contact_7  contact_7_205
timestamp 1624494425
transform 1 0 74 0 1 19908
box 0 0 58 66
use contact_8  contact_8_205
timestamp 1624494425
transform 1 0 71 0 1 19909
box 0 0 64 64
use wordline_driver  wordline_driver_204
timestamp 1624494425
transform 1 0 0 0 -1 20540
box 70 -56 4140 490
use wordline_driver  wordline_driver_205
timestamp 1624494425
transform 1 0 0 0 1 19750
box 70 -56 4140 490
use contact_7  contact_7_204
timestamp 1624494425
transform 1 0 74 0 1 20316
box 0 0 58 66
use contact_8  contact_8_204
timestamp 1624494425
transform 1 0 71 0 1 20317
box 0 0 64 64
use contact_7  contact_7_203
timestamp 1624494425
transform 1 0 74 0 1 20698
box 0 0 58 66
use contact_8  contact_8_203
timestamp 1624494425
transform 1 0 71 0 1 20699
box 0 0 64 64
use wordline_driver  wordline_driver_203
timestamp 1624494425
transform 1 0 0 0 1 20540
box 70 -56 4140 490
use contact_7  contact_7_202
timestamp 1624494425
transform 1 0 74 0 1 21106
box 0 0 58 66
use contact_8  contact_8_202
timestamp 1624494425
transform 1 0 71 0 1 21107
box 0 0 64 64
use wordline_driver  wordline_driver_201
timestamp 1624494425
transform 1 0 0 0 1 21330
box 70 -56 4140 490
use wordline_driver  wordline_driver_202
timestamp 1624494425
transform 1 0 0 0 -1 21330
box 70 -56 4140 490
use contact_7  contact_7_201
timestamp 1624494425
transform 1 0 74 0 1 21488
box 0 0 58 66
use contact_8  contact_8_201
timestamp 1624494425
transform 1 0 71 0 1 21489
box 0 0 64 64
use wordline_driver  wordline_driver_200
timestamp 1624494425
transform 1 0 0 0 -1 22120
box 70 -56 4140 490
use contact_7  contact_7_200
timestamp 1624494425
transform 1 0 74 0 1 21896
box 0 0 58 66
use contact_8  contact_8_200
timestamp 1624494425
transform 1 0 71 0 1 21897
box 0 0 64 64
use contact_7  contact_7_199
timestamp 1624494425
transform 1 0 74 0 1 22278
box 0 0 58 66
use contact_8  contact_8_199
timestamp 1624494425
transform 1 0 71 0 1 22279
box 0 0 64 64
use wordline_driver  wordline_driver_199
timestamp 1624494425
transform 1 0 0 0 1 22120
box 70 -56 4140 490
use contact_7  contact_7_198
timestamp 1624494425
transform 1 0 74 0 1 22686
box 0 0 58 66
use contact_8  contact_8_198
timestamp 1624494425
transform 1 0 71 0 1 22687
box 0 0 64 64
use wordline_driver  wordline_driver_197
timestamp 1624494425
transform 1 0 0 0 1 22910
box 70 -56 4140 490
use wordline_driver  wordline_driver_198
timestamp 1624494425
transform 1 0 0 0 -1 22910
box 70 -56 4140 490
use contact_7  contact_7_197
timestamp 1624494425
transform 1 0 74 0 1 23068
box 0 0 58 66
use contact_8  contact_8_197
timestamp 1624494425
transform 1 0 71 0 1 23069
box 0 0 64 64
use wordline_driver  wordline_driver_196
timestamp 1624494425
transform 1 0 0 0 -1 23700
box 70 -56 4140 490
use contact_7  contact_7_196
timestamp 1624494425
transform 1 0 74 0 1 23476
box 0 0 58 66
use contact_8  contact_8_196
timestamp 1624494425
transform 1 0 71 0 1 23477
box 0 0 64 64
use contact_7  contact_7_195
timestamp 1624494425
transform 1 0 74 0 1 23858
box 0 0 58 66
use contact_8  contact_8_195
timestamp 1624494425
transform 1 0 71 0 1 23859
box 0 0 64 64
use wordline_driver  wordline_driver_194
timestamp 1624494425
transform 1 0 0 0 -1 24490
box 70 -56 4140 490
use wordline_driver  wordline_driver_195
timestamp 1624494425
transform 1 0 0 0 1 23700
box 70 -56 4140 490
use contact_7  contact_7_194
timestamp 1624494425
transform 1 0 74 0 1 24266
box 0 0 58 66
use contact_8  contact_8_194
timestamp 1624494425
transform 1 0 71 0 1 24267
box 0 0 64 64
use wordline_driver  wordline_driver_193
timestamp 1624494425
transform 1 0 0 0 1 24490
box 70 -56 4140 490
use contact_7  contact_7_193
timestamp 1624494425
transform 1 0 74 0 1 24648
box 0 0 58 66
use contact_8  contact_8_193
timestamp 1624494425
transform 1 0 71 0 1 24649
box 0 0 64 64
use contact_7  contact_7_192
timestamp 1624494425
transform 1 0 74 0 1 25056
box 0 0 58 66
use contact_8  contact_8_192
timestamp 1624494425
transform 1 0 71 0 1 25057
box 0 0 64 64
use wordline_driver  wordline_driver_192
timestamp 1624494425
transform 1 0 0 0 -1 25280
box 70 -56 4140 490
use contact_7  contact_7_191
timestamp 1624494425
transform 1 0 74 0 1 25438
box 0 0 58 66
use contact_8  contact_8_191
timestamp 1624494425
transform 1 0 71 0 1 25439
box 0 0 64 64
use wordline_driver  wordline_driver_190
timestamp 1624494425
transform 1 0 0 0 -1 26070
box 70 -56 4140 490
use wordline_driver  wordline_driver_191
timestamp 1624494425
transform 1 0 0 0 1 25280
box 70 -56 4140 490
use contact_7  contact_7_190
timestamp 1624494425
transform 1 0 74 0 1 25846
box 0 0 58 66
use contact_8  contact_8_190
timestamp 1624494425
transform 1 0 71 0 1 25847
box 0 0 64 64
use wordline_driver  wordline_driver_189
timestamp 1624494425
transform 1 0 0 0 1 26070
box 70 -56 4140 490
use contact_7  contact_7_189
timestamp 1624494425
transform 1 0 74 0 1 26228
box 0 0 58 66
use contact_8  contact_8_189
timestamp 1624494425
transform 1 0 71 0 1 26229
box 0 0 64 64
use contact_7  contact_7_188
timestamp 1624494425
transform 1 0 74 0 1 26636
box 0 0 58 66
use contact_8  contact_8_188
timestamp 1624494425
transform 1 0 71 0 1 26637
box 0 0 64 64
use wordline_driver  wordline_driver_188
timestamp 1624494425
transform 1 0 0 0 -1 26860
box 70 -56 4140 490
use contact_7  contact_7_187
timestamp 1624494425
transform 1 0 74 0 1 27018
box 0 0 58 66
use contact_8  contact_8_187
timestamp 1624494425
transform 1 0 71 0 1 27019
box 0 0 64 64
use wordline_driver  wordline_driver_186
timestamp 1624494425
transform 1 0 0 0 -1 27650
box 70 -56 4140 490
use wordline_driver  wordline_driver_187
timestamp 1624494425
transform 1 0 0 0 1 26860
box 70 -56 4140 490
use contact_7  contact_7_186
timestamp 1624494425
transform 1 0 74 0 1 27426
box 0 0 58 66
use contact_8  contact_8_186
timestamp 1624494425
transform 1 0 71 0 1 27427
box 0 0 64 64
use contact_7  contact_7_185
timestamp 1624494425
transform 1 0 74 0 1 27808
box 0 0 58 66
use contact_8  contact_8_185
timestamp 1624494425
transform 1 0 71 0 1 27809
box 0 0 64 64
use wordline_driver  wordline_driver_185
timestamp 1624494425
transform 1 0 0 0 1 27650
box 70 -56 4140 490
use contact_7  contact_7_184
timestamp 1624494425
transform 1 0 74 0 1 28216
box 0 0 58 66
use contact_8  contact_8_184
timestamp 1624494425
transform 1 0 71 0 1 28217
box 0 0 64 64
use wordline_driver  wordline_driver_183
timestamp 1624494425
transform 1 0 0 0 1 28440
box 70 -56 4140 490
use wordline_driver  wordline_driver_184
timestamp 1624494425
transform 1 0 0 0 -1 28440
box 70 -56 4140 490
use contact_7  contact_7_183
timestamp 1624494425
transform 1 0 74 0 1 28598
box 0 0 58 66
use contact_8  contact_8_183
timestamp 1624494425
transform 1 0 71 0 1 28599
box 0 0 64 64
use wordline_driver  wordline_driver_182
timestamp 1624494425
transform 1 0 0 0 -1 29230
box 70 -56 4140 490
use contact_7  contact_7_182
timestamp 1624494425
transform 1 0 74 0 1 29006
box 0 0 58 66
use contact_8  contact_8_182
timestamp 1624494425
transform 1 0 71 0 1 29007
box 0 0 64 64
use contact_7  contact_7_181
timestamp 1624494425
transform 1 0 74 0 1 29388
box 0 0 58 66
use contact_8  contact_8_181
timestamp 1624494425
transform 1 0 71 0 1 29389
box 0 0 64 64
use wordline_driver  wordline_driver_181
timestamp 1624494425
transform 1 0 0 0 1 29230
box 70 -56 4140 490
use contact_7  contact_7_180
timestamp 1624494425
transform 1 0 74 0 1 29796
box 0 0 58 66
use contact_8  contact_8_180
timestamp 1624494425
transform 1 0 71 0 1 29797
box 0 0 64 64
use wordline_driver  wordline_driver_179
timestamp 1624494425
transform 1 0 0 0 1 30020
box 70 -56 4140 490
use wordline_driver  wordline_driver_180
timestamp 1624494425
transform 1 0 0 0 -1 30020
box 70 -56 4140 490
use contact_7  contact_7_179
timestamp 1624494425
transform 1 0 74 0 1 30178
box 0 0 58 66
use contact_8  contact_8_179
timestamp 1624494425
transform 1 0 71 0 1 30179
box 0 0 64 64
use wordline_driver  wordline_driver_178
timestamp 1624494425
transform 1 0 0 0 -1 30810
box 70 -56 4140 490
use contact_7  contact_7_178
timestamp 1624494425
transform 1 0 74 0 1 30586
box 0 0 58 66
use contact_8  contact_8_178
timestamp 1624494425
transform 1 0 71 0 1 30587
box 0 0 64 64
use contact_7  contact_7_177
timestamp 1624494425
transform 1 0 74 0 1 30968
box 0 0 58 66
use contact_8  contact_8_177
timestamp 1624494425
transform 1 0 71 0 1 30969
box 0 0 64 64
use wordline_driver  wordline_driver_176
timestamp 1624494425
transform 1 0 0 0 -1 31600
box 70 -56 4140 490
use wordline_driver  wordline_driver_177
timestamp 1624494425
transform 1 0 0 0 1 30810
box 70 -56 4140 490
use contact_7  contact_7_176
timestamp 1624494425
transform 1 0 74 0 1 31376
box 0 0 58 66
use contact_8  contact_8_176
timestamp 1624494425
transform 1 0 71 0 1 31377
box 0 0 64 64
use wordline_driver  wordline_driver_175
timestamp 1624494425
transform 1 0 0 0 1 31600
box 70 -56 4140 490
use contact_7  contact_7_175
timestamp 1624494425
transform 1 0 74 0 1 31758
box 0 0 58 66
use contact_8  contact_8_175
timestamp 1624494425
transform 1 0 71 0 1 31759
box 0 0 64 64
use contact_7  contact_7_174
timestamp 1624494425
transform 1 0 74 0 1 32166
box 0 0 58 66
use contact_8  contact_8_174
timestamp 1624494425
transform 1 0 71 0 1 32167
box 0 0 64 64
use wordline_driver  wordline_driver_174
timestamp 1624494425
transform 1 0 0 0 -1 32390
box 70 -56 4140 490
use contact_7  contact_7_173
timestamp 1624494425
transform 1 0 74 0 1 32548
box 0 0 58 66
use contact_8  contact_8_173
timestamp 1624494425
transform 1 0 71 0 1 32549
box 0 0 64 64
use wordline_driver  wordline_driver_172
timestamp 1624494425
transform 1 0 0 0 -1 33180
box 70 -56 4140 490
use wordline_driver  wordline_driver_173
timestamp 1624494425
transform 1 0 0 0 1 32390
box 70 -56 4140 490
use contact_7  contact_7_172
timestamp 1624494425
transform 1 0 74 0 1 32956
box 0 0 58 66
use contact_8  contact_8_172
timestamp 1624494425
transform 1 0 71 0 1 32957
box 0 0 64 64
use wordline_driver  wordline_driver_171
timestamp 1624494425
transform 1 0 0 0 1 33180
box 70 -56 4140 490
use contact_7  contact_7_171
timestamp 1624494425
transform 1 0 74 0 1 33338
box 0 0 58 66
use contact_8  contact_8_171
timestamp 1624494425
transform 1 0 71 0 1 33339
box 0 0 64 64
use contact_7  contact_7_170
timestamp 1624494425
transform 1 0 74 0 1 33746
box 0 0 58 66
use contact_8  contact_8_170
timestamp 1624494425
transform 1 0 71 0 1 33747
box 0 0 64 64
use wordline_driver  wordline_driver_170
timestamp 1624494425
transform 1 0 0 0 -1 33970
box 70 -56 4140 490
use contact_7  contact_7_169
timestamp 1624494425
transform 1 0 74 0 1 34128
box 0 0 58 66
use contact_8  contact_8_169
timestamp 1624494425
transform 1 0 71 0 1 34129
box 0 0 64 64
use wordline_driver  wordline_driver_168
timestamp 1624494425
transform 1 0 0 0 -1 34760
box 70 -56 4140 490
use wordline_driver  wordline_driver_169
timestamp 1624494425
transform 1 0 0 0 1 33970
box 70 -56 4140 490
use contact_7  contact_7_168
timestamp 1624494425
transform 1 0 74 0 1 34536
box 0 0 58 66
use contact_8  contact_8_168
timestamp 1624494425
transform 1 0 71 0 1 34537
box 0 0 64 64
use contact_7  contact_7_167
timestamp 1624494425
transform 1 0 74 0 1 34918
box 0 0 58 66
use contact_8  contact_8_167
timestamp 1624494425
transform 1 0 71 0 1 34919
box 0 0 64 64
use wordline_driver  wordline_driver_167
timestamp 1624494425
transform 1 0 0 0 1 34760
box 70 -56 4140 490
use contact_7  contact_7_166
timestamp 1624494425
transform 1 0 74 0 1 35326
box 0 0 58 66
use contact_8  contact_8_166
timestamp 1624494425
transform 1 0 71 0 1 35327
box 0 0 64 64
use wordline_driver  wordline_driver_165
timestamp 1624494425
transform 1 0 0 0 1 35550
box 70 -56 4140 490
use wordline_driver  wordline_driver_166
timestamp 1624494425
transform 1 0 0 0 -1 35550
box 70 -56 4140 490
use contact_7  contact_7_165
timestamp 1624494425
transform 1 0 74 0 1 35708
box 0 0 58 66
use contact_8  contact_8_165
timestamp 1624494425
transform 1 0 71 0 1 35709
box 0 0 64 64
use wordline_driver  wordline_driver_164
timestamp 1624494425
transform 1 0 0 0 -1 36340
box 70 -56 4140 490
use contact_7  contact_7_164
timestamp 1624494425
transform 1 0 74 0 1 36116
box 0 0 58 66
use contact_8  contact_8_164
timestamp 1624494425
transform 1 0 71 0 1 36117
box 0 0 64 64
use contact_7  contact_7_163
timestamp 1624494425
transform 1 0 74 0 1 36498
box 0 0 58 66
use contact_8  contact_8_163
timestamp 1624494425
transform 1 0 71 0 1 36499
box 0 0 64 64
use wordline_driver  wordline_driver_163
timestamp 1624494425
transform 1 0 0 0 1 36340
box 70 -56 4140 490
use contact_7  contact_7_162
timestamp 1624494425
transform 1 0 74 0 1 36906
box 0 0 58 66
use contact_8  contact_8_162
timestamp 1624494425
transform 1 0 71 0 1 36907
box 0 0 64 64
use wordline_driver  wordline_driver_161
timestamp 1624494425
transform 1 0 0 0 1 37130
box 70 -56 4140 490
use wordline_driver  wordline_driver_162
timestamp 1624494425
transform 1 0 0 0 -1 37130
box 70 -56 4140 490
use contact_7  contact_7_161
timestamp 1624494425
transform 1 0 74 0 1 37288
box 0 0 58 66
use contact_8  contact_8_161
timestamp 1624494425
transform 1 0 71 0 1 37289
box 0 0 64 64
use wordline_driver  wordline_driver_160
timestamp 1624494425
transform 1 0 0 0 -1 37920
box 70 -56 4140 490
use contact_7  contact_7_160
timestamp 1624494425
transform 1 0 74 0 1 37696
box 0 0 58 66
use contact_8  contact_8_160
timestamp 1624494425
transform 1 0 71 0 1 37697
box 0 0 64 64
use contact_7  contact_7_159
timestamp 1624494425
transform 1 0 74 0 1 38078
box 0 0 58 66
use contact_8  contact_8_159
timestamp 1624494425
transform 1 0 71 0 1 38079
box 0 0 64 64
use wordline_driver  wordline_driver_158
timestamp 1624494425
transform 1 0 0 0 -1 38710
box 70 -56 4140 490
use wordline_driver  wordline_driver_159
timestamp 1624494425
transform 1 0 0 0 1 37920
box 70 -56 4140 490
use contact_7  contact_7_158
timestamp 1624494425
transform 1 0 74 0 1 38486
box 0 0 58 66
use contact_8  contact_8_158
timestamp 1624494425
transform 1 0 71 0 1 38487
box 0 0 64 64
use wordline_driver  wordline_driver_157
timestamp 1624494425
transform 1 0 0 0 1 38710
box 70 -56 4140 490
use contact_7  contact_7_157
timestamp 1624494425
transform 1 0 74 0 1 38868
box 0 0 58 66
use contact_8  contact_8_157
timestamp 1624494425
transform 1 0 71 0 1 38869
box 0 0 64 64
use contact_7  contact_7_156
timestamp 1624494425
transform 1 0 74 0 1 39276
box 0 0 58 66
use contact_8  contact_8_156
timestamp 1624494425
transform 1 0 71 0 1 39277
box 0 0 64 64
use wordline_driver  wordline_driver_156
timestamp 1624494425
transform 1 0 0 0 -1 39500
box 70 -56 4140 490
use contact_7  contact_7_155
timestamp 1624494425
transform 1 0 74 0 1 39658
box 0 0 58 66
use contact_8  contact_8_155
timestamp 1624494425
transform 1 0 71 0 1 39659
box 0 0 64 64
use wordline_driver  wordline_driver_154
timestamp 1624494425
transform 1 0 0 0 -1 40290
box 70 -56 4140 490
use wordline_driver  wordline_driver_155
timestamp 1624494425
transform 1 0 0 0 1 39500
box 70 -56 4140 490
use contact_7  contact_7_154
timestamp 1624494425
transform 1 0 74 0 1 40066
box 0 0 58 66
use contact_8  contact_8_154
timestamp 1624494425
transform 1 0 71 0 1 40067
box 0 0 64 64
use wordline_driver  wordline_driver_153
timestamp 1624494425
transform 1 0 0 0 1 40290
box 70 -56 4140 490
use contact_7  contact_7_153
timestamp 1624494425
transform 1 0 74 0 1 40448
box 0 0 58 66
use contact_8  contact_8_153
timestamp 1624494425
transform 1 0 71 0 1 40449
box 0 0 64 64
use contact_7  contact_7_152
timestamp 1624494425
transform 1 0 74 0 1 40856
box 0 0 58 66
use contact_8  contact_8_152
timestamp 1624494425
transform 1 0 71 0 1 40857
box 0 0 64 64
use wordline_driver  wordline_driver_152
timestamp 1624494425
transform 1 0 0 0 -1 41080
box 70 -56 4140 490
use contact_7  contact_7_151
timestamp 1624494425
transform 1 0 74 0 1 41238
box 0 0 58 66
use contact_8  contact_8_151
timestamp 1624494425
transform 1 0 71 0 1 41239
box 0 0 64 64
use wordline_driver  wordline_driver_150
timestamp 1624494425
transform 1 0 0 0 -1 41870
box 70 -56 4140 490
use wordline_driver  wordline_driver_151
timestamp 1624494425
transform 1 0 0 0 1 41080
box 70 -56 4140 490
use contact_7  contact_7_150
timestamp 1624494425
transform 1 0 74 0 1 41646
box 0 0 58 66
use contact_8  contact_8_150
timestamp 1624494425
transform 1 0 71 0 1 41647
box 0 0 64 64
use contact_7  contact_7_149
timestamp 1624494425
transform 1 0 74 0 1 42028
box 0 0 58 66
use contact_8  contact_8_149
timestamp 1624494425
transform 1 0 71 0 1 42029
box 0 0 64 64
use wordline_driver  wordline_driver_149
timestamp 1624494425
transform 1 0 0 0 1 41870
box 70 -56 4140 490
use contact_7  contact_7_148
timestamp 1624494425
transform 1 0 74 0 1 42436
box 0 0 58 66
use contact_8  contact_8_148
timestamp 1624494425
transform 1 0 71 0 1 42437
box 0 0 64 64
use wordline_driver  wordline_driver_147
timestamp 1624494425
transform 1 0 0 0 1 42660
box 70 -56 4140 490
use wordline_driver  wordline_driver_148
timestamp 1624494425
transform 1 0 0 0 -1 42660
box 70 -56 4140 490
use contact_7  contact_7_147
timestamp 1624494425
transform 1 0 74 0 1 42818
box 0 0 58 66
use contact_8  contact_8_147
timestamp 1624494425
transform 1 0 71 0 1 42819
box 0 0 64 64
use wordline_driver  wordline_driver_146
timestamp 1624494425
transform 1 0 0 0 -1 43450
box 70 -56 4140 490
use contact_7  contact_7_146
timestamp 1624494425
transform 1 0 74 0 1 43226
box 0 0 58 66
use contact_8  contact_8_146
timestamp 1624494425
transform 1 0 71 0 1 43227
box 0 0 64 64
use contact_7  contact_7_145
timestamp 1624494425
transform 1 0 74 0 1 43608
box 0 0 58 66
use contact_8  contact_8_145
timestamp 1624494425
transform 1 0 71 0 1 43609
box 0 0 64 64
use wordline_driver  wordline_driver_145
timestamp 1624494425
transform 1 0 0 0 1 43450
box 70 -56 4140 490
use contact_7  contact_7_144
timestamp 1624494425
transform 1 0 74 0 1 44016
box 0 0 58 66
use contact_8  contact_8_144
timestamp 1624494425
transform 1 0 71 0 1 44017
box 0 0 64 64
use wordline_driver  wordline_driver_143
timestamp 1624494425
transform 1 0 0 0 1 44240
box 70 -56 4140 490
use wordline_driver  wordline_driver_144
timestamp 1624494425
transform 1 0 0 0 -1 44240
box 70 -56 4140 490
use contact_7  contact_7_143
timestamp 1624494425
transform 1 0 74 0 1 44398
box 0 0 58 66
use contact_8  contact_8_143
timestamp 1624494425
transform 1 0 71 0 1 44399
box 0 0 64 64
use wordline_driver  wordline_driver_142
timestamp 1624494425
transform 1 0 0 0 -1 45030
box 70 -56 4140 490
use contact_7  contact_7_142
timestamp 1624494425
transform 1 0 74 0 1 44806
box 0 0 58 66
use contact_8  contact_8_142
timestamp 1624494425
transform 1 0 71 0 1 44807
box 0 0 64 64
use contact_7  contact_7_141
timestamp 1624494425
transform 1 0 74 0 1 45188
box 0 0 58 66
use contact_8  contact_8_141
timestamp 1624494425
transform 1 0 71 0 1 45189
box 0 0 64 64
use wordline_driver  wordline_driver_140
timestamp 1624494425
transform 1 0 0 0 -1 45820
box 70 -56 4140 490
use wordline_driver  wordline_driver_141
timestamp 1624494425
transform 1 0 0 0 1 45030
box 70 -56 4140 490
use contact_7  contact_7_140
timestamp 1624494425
transform 1 0 74 0 1 45596
box 0 0 58 66
use contact_8  contact_8_140
timestamp 1624494425
transform 1 0 71 0 1 45597
box 0 0 64 64
use wordline_driver  wordline_driver_139
timestamp 1624494425
transform 1 0 0 0 1 45820
box 70 -56 4140 490
use contact_7  contact_7_139
timestamp 1624494425
transform 1 0 74 0 1 45978
box 0 0 58 66
use contact_8  contact_8_139
timestamp 1624494425
transform 1 0 71 0 1 45979
box 0 0 64 64
use contact_7  contact_7_138
timestamp 1624494425
transform 1 0 74 0 1 46386
box 0 0 58 66
use contact_8  contact_8_138
timestamp 1624494425
transform 1 0 71 0 1 46387
box 0 0 64 64
use wordline_driver  wordline_driver_138
timestamp 1624494425
transform 1 0 0 0 -1 46610
box 70 -56 4140 490
use contact_7  contact_7_137
timestamp 1624494425
transform 1 0 74 0 1 46768
box 0 0 58 66
use contact_8  contact_8_137
timestamp 1624494425
transform 1 0 71 0 1 46769
box 0 0 64 64
use wordline_driver  wordline_driver_136
timestamp 1624494425
transform 1 0 0 0 -1 47400
box 70 -56 4140 490
use wordline_driver  wordline_driver_137
timestamp 1624494425
transform 1 0 0 0 1 46610
box 70 -56 4140 490
use contact_7  contact_7_136
timestamp 1624494425
transform 1 0 74 0 1 47176
box 0 0 58 66
use contact_8  contact_8_136
timestamp 1624494425
transform 1 0 71 0 1 47177
box 0 0 64 64
use wordline_driver  wordline_driver_135
timestamp 1624494425
transform 1 0 0 0 1 47400
box 70 -56 4140 490
use contact_7  contact_7_135
timestamp 1624494425
transform 1 0 74 0 1 47558
box 0 0 58 66
use contact_8  contact_8_135
timestamp 1624494425
transform 1 0 71 0 1 47559
box 0 0 64 64
use contact_7  contact_7_134
timestamp 1624494425
transform 1 0 74 0 1 47966
box 0 0 58 66
use contact_8  contact_8_134
timestamp 1624494425
transform 1 0 71 0 1 47967
box 0 0 64 64
use wordline_driver  wordline_driver_134
timestamp 1624494425
transform 1 0 0 0 -1 48190
box 70 -56 4140 490
use contact_7  contact_7_133
timestamp 1624494425
transform 1 0 74 0 1 48348
box 0 0 58 66
use contact_8  contact_8_133
timestamp 1624494425
transform 1 0 71 0 1 48349
box 0 0 64 64
use wordline_driver  wordline_driver_132
timestamp 1624494425
transform 1 0 0 0 -1 48980
box 70 -56 4140 490
use wordline_driver  wordline_driver_133
timestamp 1624494425
transform 1 0 0 0 1 48190
box 70 -56 4140 490
use contact_7  contact_7_132
timestamp 1624494425
transform 1 0 74 0 1 48756
box 0 0 58 66
use contact_8  contact_8_132
timestamp 1624494425
transform 1 0 71 0 1 48757
box 0 0 64 64
use contact_7  contact_7_131
timestamp 1624494425
transform 1 0 74 0 1 49138
box 0 0 58 66
use contact_8  contact_8_131
timestamp 1624494425
transform 1 0 71 0 1 49139
box 0 0 64 64
use wordline_driver  wordline_driver_131
timestamp 1624494425
transform 1 0 0 0 1 48980
box 70 -56 4140 490
use contact_7  contact_7_130
timestamp 1624494425
transform 1 0 74 0 1 49546
box 0 0 58 66
use contact_8  contact_8_130
timestamp 1624494425
transform 1 0 71 0 1 49547
box 0 0 64 64
use wordline_driver  wordline_driver_129
timestamp 1624494425
transform 1 0 0 0 1 49770
box 70 -56 4140 490
use wordline_driver  wordline_driver_130
timestamp 1624494425
transform 1 0 0 0 -1 49770
box 70 -56 4140 490
use contact_7  contact_7_129
timestamp 1624494425
transform 1 0 74 0 1 49928
box 0 0 58 66
use contact_8  contact_8_129
timestamp 1624494425
transform 1 0 71 0 1 49929
box 0 0 64 64
use wordline_driver  wordline_driver_128
timestamp 1624494425
transform 1 0 0 0 -1 50560
box 70 -56 4140 490
use contact_7  contact_7_128
timestamp 1624494425
transform 1 0 74 0 1 50336
box 0 0 58 66
use contact_8  contact_8_128
timestamp 1624494425
transform 1 0 71 0 1 50337
box 0 0 64 64
use contact_7  contact_7_127
timestamp 1624494425
transform 1 0 74 0 1 50718
box 0 0 58 66
use contact_8  contact_8_127
timestamp 1624494425
transform 1 0 71 0 1 50719
box 0 0 64 64
use wordline_driver  wordline_driver_127
timestamp 1624494425
transform 1 0 0 0 1 50560
box 70 -56 4140 490
use contact_7  contact_7_126
timestamp 1624494425
transform 1 0 74 0 1 51126
box 0 0 58 66
use contact_8  contact_8_126
timestamp 1624494425
transform 1 0 71 0 1 51127
box 0 0 64 64
use wordline_driver  wordline_driver_125
timestamp 1624494425
transform 1 0 0 0 1 51350
box 70 -56 4140 490
use wordline_driver  wordline_driver_126
timestamp 1624494425
transform 1 0 0 0 -1 51350
box 70 -56 4140 490
use contact_7  contact_7_125
timestamp 1624494425
transform 1 0 74 0 1 51508
box 0 0 58 66
use contact_8  contact_8_125
timestamp 1624494425
transform 1 0 71 0 1 51509
box 0 0 64 64
use wordline_driver  wordline_driver_124
timestamp 1624494425
transform 1 0 0 0 -1 52140
box 70 -56 4140 490
use contact_7  contact_7_124
timestamp 1624494425
transform 1 0 74 0 1 51916
box 0 0 58 66
use contact_8  contact_8_124
timestamp 1624494425
transform 1 0 71 0 1 51917
box 0 0 64 64
use contact_7  contact_7_123
timestamp 1624494425
transform 1 0 74 0 1 52298
box 0 0 58 66
use contact_8  contact_8_123
timestamp 1624494425
transform 1 0 71 0 1 52299
box 0 0 64 64
use wordline_driver  wordline_driver_122
timestamp 1624494425
transform 1 0 0 0 -1 52930
box 70 -56 4140 490
use wordline_driver  wordline_driver_123
timestamp 1624494425
transform 1 0 0 0 1 52140
box 70 -56 4140 490
use contact_7  contact_7_122
timestamp 1624494425
transform 1 0 74 0 1 52706
box 0 0 58 66
use contact_8  contact_8_122
timestamp 1624494425
transform 1 0 71 0 1 52707
box 0 0 64 64
use wordline_driver  wordline_driver_121
timestamp 1624494425
transform 1 0 0 0 1 52930
box 70 -56 4140 490
use contact_7  contact_7_121
timestamp 1624494425
transform 1 0 74 0 1 53088
box 0 0 58 66
use contact_8  contact_8_121
timestamp 1624494425
transform 1 0 71 0 1 53089
box 0 0 64 64
use contact_7  contact_7_120
timestamp 1624494425
transform 1 0 74 0 1 53496
box 0 0 58 66
use contact_8  contact_8_120
timestamp 1624494425
transform 1 0 71 0 1 53497
box 0 0 64 64
use wordline_driver  wordline_driver_120
timestamp 1624494425
transform 1 0 0 0 -1 53720
box 70 -56 4140 490
use contact_7  contact_7_119
timestamp 1624494425
transform 1 0 74 0 1 53878
box 0 0 58 66
use contact_8  contact_8_119
timestamp 1624494425
transform 1 0 71 0 1 53879
box 0 0 64 64
use wordline_driver  wordline_driver_118
timestamp 1624494425
transform 1 0 0 0 -1 54510
box 70 -56 4140 490
use wordline_driver  wordline_driver_119
timestamp 1624494425
transform 1 0 0 0 1 53720
box 70 -56 4140 490
use contact_7  contact_7_118
timestamp 1624494425
transform 1 0 74 0 1 54286
box 0 0 58 66
use contact_8  contact_8_118
timestamp 1624494425
transform 1 0 71 0 1 54287
box 0 0 64 64
use wordline_driver  wordline_driver_117
timestamp 1624494425
transform 1 0 0 0 1 54510
box 70 -56 4140 490
use contact_7  contact_7_117
timestamp 1624494425
transform 1 0 74 0 1 54668
box 0 0 58 66
use contact_8  contact_8_117
timestamp 1624494425
transform 1 0 71 0 1 54669
box 0 0 64 64
use contact_7  contact_7_116
timestamp 1624494425
transform 1 0 74 0 1 55076
box 0 0 58 66
use contact_8  contact_8_116
timestamp 1624494425
transform 1 0 71 0 1 55077
box 0 0 64 64
use wordline_driver  wordline_driver_116
timestamp 1624494425
transform 1 0 0 0 -1 55300
box 70 -56 4140 490
use contact_7  contact_7_115
timestamp 1624494425
transform 1 0 74 0 1 55458
box 0 0 58 66
use contact_8  contact_8_115
timestamp 1624494425
transform 1 0 71 0 1 55459
box 0 0 64 64
use wordline_driver  wordline_driver_114
timestamp 1624494425
transform 1 0 0 0 -1 56090
box 70 -56 4140 490
use wordline_driver  wordline_driver_115
timestamp 1624494425
transform 1 0 0 0 1 55300
box 70 -56 4140 490
use contact_7  contact_7_114
timestamp 1624494425
transform 1 0 74 0 1 55866
box 0 0 58 66
use contact_8  contact_8_114
timestamp 1624494425
transform 1 0 71 0 1 55867
box 0 0 64 64
use contact_7  contact_7_113
timestamp 1624494425
transform 1 0 74 0 1 56248
box 0 0 58 66
use contact_8  contact_8_113
timestamp 1624494425
transform 1 0 71 0 1 56249
box 0 0 64 64
use wordline_driver  wordline_driver_113
timestamp 1624494425
transform 1 0 0 0 1 56090
box 70 -56 4140 490
use contact_7  contact_7_112
timestamp 1624494425
transform 1 0 74 0 1 56656
box 0 0 58 66
use contact_8  contact_8_112
timestamp 1624494425
transform 1 0 71 0 1 56657
box 0 0 64 64
use wordline_driver  wordline_driver_111
timestamp 1624494425
transform 1 0 0 0 1 56880
box 70 -56 4140 490
use wordline_driver  wordline_driver_112
timestamp 1624494425
transform 1 0 0 0 -1 56880
box 70 -56 4140 490
use contact_7  contact_7_111
timestamp 1624494425
transform 1 0 74 0 1 57038
box 0 0 58 66
use contact_8  contact_8_111
timestamp 1624494425
transform 1 0 71 0 1 57039
box 0 0 64 64
use wordline_driver  wordline_driver_110
timestamp 1624494425
transform 1 0 0 0 -1 57670
box 70 -56 4140 490
use contact_7  contact_7_110
timestamp 1624494425
transform 1 0 74 0 1 57446
box 0 0 58 66
use contact_8  contact_8_110
timestamp 1624494425
transform 1 0 71 0 1 57447
box 0 0 64 64
use contact_7  contact_7_109
timestamp 1624494425
transform 1 0 74 0 1 57828
box 0 0 58 66
use contact_8  contact_8_109
timestamp 1624494425
transform 1 0 71 0 1 57829
box 0 0 64 64
use wordline_driver  wordline_driver_109
timestamp 1624494425
transform 1 0 0 0 1 57670
box 70 -56 4140 490
use contact_7  contact_7_108
timestamp 1624494425
transform 1 0 74 0 1 58236
box 0 0 58 66
use contact_8  contact_8_108
timestamp 1624494425
transform 1 0 71 0 1 58237
box 0 0 64 64
use wordline_driver  wordline_driver_107
timestamp 1624494425
transform 1 0 0 0 1 58460
box 70 -56 4140 490
use wordline_driver  wordline_driver_108
timestamp 1624494425
transform 1 0 0 0 -1 58460
box 70 -56 4140 490
use contact_7  contact_7_107
timestamp 1624494425
transform 1 0 74 0 1 58618
box 0 0 58 66
use contact_8  contact_8_107
timestamp 1624494425
transform 1 0 71 0 1 58619
box 0 0 64 64
use wordline_driver  wordline_driver_106
timestamp 1624494425
transform 1 0 0 0 -1 59250
box 70 -56 4140 490
use contact_7  contact_7_106
timestamp 1624494425
transform 1 0 74 0 1 59026
box 0 0 58 66
use contact_8  contact_8_106
timestamp 1624494425
transform 1 0 71 0 1 59027
box 0 0 64 64
use contact_7  contact_7_105
timestamp 1624494425
transform 1 0 74 0 1 59408
box 0 0 58 66
use contact_8  contact_8_105
timestamp 1624494425
transform 1 0 71 0 1 59409
box 0 0 64 64
use wordline_driver  wordline_driver_104
timestamp 1624494425
transform 1 0 0 0 -1 60040
box 70 -56 4140 490
use wordline_driver  wordline_driver_105
timestamp 1624494425
transform 1 0 0 0 1 59250
box 70 -56 4140 490
use contact_7  contact_7_104
timestamp 1624494425
transform 1 0 74 0 1 59816
box 0 0 58 66
use contact_8  contact_8_104
timestamp 1624494425
transform 1 0 71 0 1 59817
box 0 0 64 64
use wordline_driver  wordline_driver_103
timestamp 1624494425
transform 1 0 0 0 1 60040
box 70 -56 4140 490
use contact_7  contact_7_103
timestamp 1624494425
transform 1 0 74 0 1 60198
box 0 0 58 66
use contact_8  contact_8_103
timestamp 1624494425
transform 1 0 71 0 1 60199
box 0 0 64 64
use contact_7  contact_7_102
timestamp 1624494425
transform 1 0 74 0 1 60606
box 0 0 58 66
use contact_8  contact_8_102
timestamp 1624494425
transform 1 0 71 0 1 60607
box 0 0 64 64
use wordline_driver  wordline_driver_102
timestamp 1624494425
transform 1 0 0 0 -1 60830
box 70 -56 4140 490
use contact_7  contact_7_101
timestamp 1624494425
transform 1 0 74 0 1 60988
box 0 0 58 66
use contact_8  contact_8_101
timestamp 1624494425
transform 1 0 71 0 1 60989
box 0 0 64 64
use wordline_driver  wordline_driver_100
timestamp 1624494425
transform 1 0 0 0 -1 61620
box 70 -56 4140 490
use wordline_driver  wordline_driver_101
timestamp 1624494425
transform 1 0 0 0 1 60830
box 70 -56 4140 490
use contact_7  contact_7_100
timestamp 1624494425
transform 1 0 74 0 1 61396
box 0 0 58 66
use contact_8  contact_8_100
timestamp 1624494425
transform 1 0 71 0 1 61397
box 0 0 64 64
use wordline_driver  wordline_driver_99
timestamp 1624494425
transform 1 0 0 0 1 61620
box 70 -56 4140 490
use contact_7  contact_7_99
timestamp 1624494425
transform 1 0 74 0 1 61778
box 0 0 58 66
use contact_8  contact_8_99
timestamp 1624494425
transform 1 0 71 0 1 61779
box 0 0 64 64
use contact_7  contact_7_98
timestamp 1624494425
transform 1 0 74 0 1 62186
box 0 0 58 66
use contact_8  contact_8_98
timestamp 1624494425
transform 1 0 71 0 1 62187
box 0 0 64 64
use wordline_driver  wordline_driver_98
timestamp 1624494425
transform 1 0 0 0 -1 62410
box 70 -56 4140 490
use contact_7  contact_7_97
timestamp 1624494425
transform 1 0 74 0 1 62568
box 0 0 58 66
use contact_8  contact_8_97
timestamp 1624494425
transform 1 0 71 0 1 62569
box 0 0 64 64
use wordline_driver  wordline_driver_96
timestamp 1624494425
transform 1 0 0 0 -1 63200
box 70 -56 4140 490
use wordline_driver  wordline_driver_97
timestamp 1624494425
transform 1 0 0 0 1 62410
box 70 -56 4140 490
use contact_7  contact_7_96
timestamp 1624494425
transform 1 0 74 0 1 62976
box 0 0 58 66
use contact_8  contact_8_96
timestamp 1624494425
transform 1 0 71 0 1 62977
box 0 0 64 64
use contact_7  contact_7_95
timestamp 1624494425
transform 1 0 74 0 1 63358
box 0 0 58 66
use contact_8  contact_8_95
timestamp 1624494425
transform 1 0 71 0 1 63359
box 0 0 64 64
use wordline_driver  wordline_driver_95
timestamp 1624494425
transform 1 0 0 0 1 63200
box 70 -56 4140 490
use contact_7  contact_7_94
timestamp 1624494425
transform 1 0 74 0 1 63766
box 0 0 58 66
use contact_8  contact_8_94
timestamp 1624494425
transform 1 0 71 0 1 63767
box 0 0 64 64
use wordline_driver  wordline_driver_93
timestamp 1624494425
transform 1 0 0 0 1 63990
box 70 -56 4140 490
use wordline_driver  wordline_driver_94
timestamp 1624494425
transform 1 0 0 0 -1 63990
box 70 -56 4140 490
use contact_7  contact_7_93
timestamp 1624494425
transform 1 0 74 0 1 64148
box 0 0 58 66
use contact_8  contact_8_93
timestamp 1624494425
transform 1 0 71 0 1 64149
box 0 0 64 64
use wordline_driver  wordline_driver_92
timestamp 1624494425
transform 1 0 0 0 -1 64780
box 70 -56 4140 490
use contact_7  contact_7_92
timestamp 1624494425
transform 1 0 74 0 1 64556
box 0 0 58 66
use contact_8  contact_8_92
timestamp 1624494425
transform 1 0 71 0 1 64557
box 0 0 64 64
use contact_7  contact_7_91
timestamp 1624494425
transform 1 0 74 0 1 64938
box 0 0 58 66
use contact_8  contact_8_91
timestamp 1624494425
transform 1 0 71 0 1 64939
box 0 0 64 64
use wordline_driver  wordline_driver_91
timestamp 1624494425
transform 1 0 0 0 1 64780
box 70 -56 4140 490
use contact_7  contact_7_90
timestamp 1624494425
transform 1 0 74 0 1 65346
box 0 0 58 66
use contact_8  contact_8_90
timestamp 1624494425
transform 1 0 71 0 1 65347
box 0 0 64 64
use wordline_driver  wordline_driver_89
timestamp 1624494425
transform 1 0 0 0 1 65570
box 70 -56 4140 490
use wordline_driver  wordline_driver_90
timestamp 1624494425
transform 1 0 0 0 -1 65570
box 70 -56 4140 490
use contact_7  contact_7_89
timestamp 1624494425
transform 1 0 74 0 1 65728
box 0 0 58 66
use contact_8  contact_8_89
timestamp 1624494425
transform 1 0 71 0 1 65729
box 0 0 64 64
use wordline_driver  wordline_driver_88
timestamp 1624494425
transform 1 0 0 0 -1 66360
box 70 -56 4140 490
use contact_7  contact_7_88
timestamp 1624494425
transform 1 0 74 0 1 66136
box 0 0 58 66
use contact_8  contact_8_88
timestamp 1624494425
transform 1 0 71 0 1 66137
box 0 0 64 64
use contact_7  contact_7_87
timestamp 1624494425
transform 1 0 74 0 1 66518
box 0 0 58 66
use contact_8  contact_8_87
timestamp 1624494425
transform 1 0 71 0 1 66519
box 0 0 64 64
use wordline_driver  wordline_driver_86
timestamp 1624494425
transform 1 0 0 0 -1 67150
box 70 -56 4140 490
use wordline_driver  wordline_driver_87
timestamp 1624494425
transform 1 0 0 0 1 66360
box 70 -56 4140 490
use contact_7  contact_7_86
timestamp 1624494425
transform 1 0 74 0 1 66926
box 0 0 58 66
use contact_8  contact_8_86
timestamp 1624494425
transform 1 0 71 0 1 66927
box 0 0 64 64
use wordline_driver  wordline_driver_85
timestamp 1624494425
transform 1 0 0 0 1 67150
box 70 -56 4140 490
use contact_7  contact_7_85
timestamp 1624494425
transform 1 0 74 0 1 67308
box 0 0 58 66
use contact_8  contact_8_85
timestamp 1624494425
transform 1 0 71 0 1 67309
box 0 0 64 64
use contact_7  contact_7_84
timestamp 1624494425
transform 1 0 74 0 1 67716
box 0 0 58 66
use contact_8  contact_8_84
timestamp 1624494425
transform 1 0 71 0 1 67717
box 0 0 64 64
use wordline_driver  wordline_driver_84
timestamp 1624494425
transform 1 0 0 0 -1 67940
box 70 -56 4140 490
use contact_7  contact_7_83
timestamp 1624494425
transform 1 0 74 0 1 68098
box 0 0 58 66
use contact_8  contact_8_83
timestamp 1624494425
transform 1 0 71 0 1 68099
box 0 0 64 64
use wordline_driver  wordline_driver_82
timestamp 1624494425
transform 1 0 0 0 -1 68730
box 70 -56 4140 490
use wordline_driver  wordline_driver_83
timestamp 1624494425
transform 1 0 0 0 1 67940
box 70 -56 4140 490
use contact_7  contact_7_82
timestamp 1624494425
transform 1 0 74 0 1 68506
box 0 0 58 66
use contact_8  contact_8_82
timestamp 1624494425
transform 1 0 71 0 1 68507
box 0 0 64 64
use wordline_driver  wordline_driver_81
timestamp 1624494425
transform 1 0 0 0 1 68730
box 70 -56 4140 490
use contact_7  contact_7_81
timestamp 1624494425
transform 1 0 74 0 1 68888
box 0 0 58 66
use contact_8  contact_8_81
timestamp 1624494425
transform 1 0 71 0 1 68889
box 0 0 64 64
use contact_7  contact_7_80
timestamp 1624494425
transform 1 0 74 0 1 69296
box 0 0 58 66
use contact_8  contact_8_80
timestamp 1624494425
transform 1 0 71 0 1 69297
box 0 0 64 64
use wordline_driver  wordline_driver_80
timestamp 1624494425
transform 1 0 0 0 -1 69520
box 70 -56 4140 490
use contact_7  contact_7_79
timestamp 1624494425
transform 1 0 74 0 1 69678
box 0 0 58 66
use contact_8  contact_8_79
timestamp 1624494425
transform 1 0 71 0 1 69679
box 0 0 64 64
use wordline_driver  wordline_driver_78
timestamp 1624494425
transform 1 0 0 0 -1 70310
box 70 -56 4140 490
use wordline_driver  wordline_driver_79
timestamp 1624494425
transform 1 0 0 0 1 69520
box 70 -56 4140 490
use contact_7  contact_7_78
timestamp 1624494425
transform 1 0 74 0 1 70086
box 0 0 58 66
use contact_8  contact_8_78
timestamp 1624494425
transform 1 0 71 0 1 70087
box 0 0 64 64
use contact_7  contact_7_77
timestamp 1624494425
transform 1 0 74 0 1 70468
box 0 0 58 66
use contact_8  contact_8_77
timestamp 1624494425
transform 1 0 71 0 1 70469
box 0 0 64 64
use wordline_driver  wordline_driver_77
timestamp 1624494425
transform 1 0 0 0 1 70310
box 70 -56 4140 490
use contact_7  contact_7_76
timestamp 1624494425
transform 1 0 74 0 1 70876
box 0 0 58 66
use contact_8  contact_8_76
timestamp 1624494425
transform 1 0 71 0 1 70877
box 0 0 64 64
use wordline_driver  wordline_driver_75
timestamp 1624494425
transform 1 0 0 0 1 71100
box 70 -56 4140 490
use wordline_driver  wordline_driver_76
timestamp 1624494425
transform 1 0 0 0 -1 71100
box 70 -56 4140 490
use contact_7  contact_7_75
timestamp 1624494425
transform 1 0 74 0 1 71258
box 0 0 58 66
use contact_8  contact_8_75
timestamp 1624494425
transform 1 0 71 0 1 71259
box 0 0 64 64
use wordline_driver  wordline_driver_74
timestamp 1624494425
transform 1 0 0 0 -1 71890
box 70 -56 4140 490
use contact_7  contact_7_74
timestamp 1624494425
transform 1 0 74 0 1 71666
box 0 0 58 66
use contact_8  contact_8_74
timestamp 1624494425
transform 1 0 71 0 1 71667
box 0 0 64 64
use contact_7  contact_7_73
timestamp 1624494425
transform 1 0 74 0 1 72048
box 0 0 58 66
use contact_8  contact_8_73
timestamp 1624494425
transform 1 0 71 0 1 72049
box 0 0 64 64
use wordline_driver  wordline_driver_73
timestamp 1624494425
transform 1 0 0 0 1 71890
box 70 -56 4140 490
use contact_7  contact_7_72
timestamp 1624494425
transform 1 0 74 0 1 72456
box 0 0 58 66
use contact_8  contact_8_72
timestamp 1624494425
transform 1 0 71 0 1 72457
box 0 0 64 64
use wordline_driver  wordline_driver_71
timestamp 1624494425
transform 1 0 0 0 1 72680
box 70 -56 4140 490
use wordline_driver  wordline_driver_72
timestamp 1624494425
transform 1 0 0 0 -1 72680
box 70 -56 4140 490
use contact_7  contact_7_71
timestamp 1624494425
transform 1 0 74 0 1 72838
box 0 0 58 66
use contact_8  contact_8_71
timestamp 1624494425
transform 1 0 71 0 1 72839
box 0 0 64 64
use wordline_driver  wordline_driver_70
timestamp 1624494425
transform 1 0 0 0 -1 73470
box 70 -56 4140 490
use contact_7  contact_7_70
timestamp 1624494425
transform 1 0 74 0 1 73246
box 0 0 58 66
use contact_8  contact_8_70
timestamp 1624494425
transform 1 0 71 0 1 73247
box 0 0 64 64
use contact_7  contact_7_69
timestamp 1624494425
transform 1 0 74 0 1 73628
box 0 0 58 66
use contact_8  contact_8_69
timestamp 1624494425
transform 1 0 71 0 1 73629
box 0 0 64 64
use wordline_driver  wordline_driver_68
timestamp 1624494425
transform 1 0 0 0 -1 74260
box 70 -56 4140 490
use wordline_driver  wordline_driver_69
timestamp 1624494425
transform 1 0 0 0 1 73470
box 70 -56 4140 490
use contact_7  contact_7_68
timestamp 1624494425
transform 1 0 74 0 1 74036
box 0 0 58 66
use contact_8  contact_8_68
timestamp 1624494425
transform 1 0 71 0 1 74037
box 0 0 64 64
use wordline_driver  wordline_driver_67
timestamp 1624494425
transform 1 0 0 0 1 74260
box 70 -56 4140 490
use contact_7  contact_7_67
timestamp 1624494425
transform 1 0 74 0 1 74418
box 0 0 58 66
use contact_8  contact_8_67
timestamp 1624494425
transform 1 0 71 0 1 74419
box 0 0 64 64
use contact_7  contact_7_66
timestamp 1624494425
transform 1 0 74 0 1 74826
box 0 0 58 66
use contact_8  contact_8_66
timestamp 1624494425
transform 1 0 71 0 1 74827
box 0 0 64 64
use wordline_driver  wordline_driver_66
timestamp 1624494425
transform 1 0 0 0 -1 75050
box 70 -56 4140 490
use contact_7  contact_7_65
timestamp 1624494425
transform 1 0 74 0 1 75208
box 0 0 58 66
use contact_8  contact_8_65
timestamp 1624494425
transform 1 0 71 0 1 75209
box 0 0 64 64
use wordline_driver  wordline_driver_64
timestamp 1624494425
transform 1 0 0 0 -1 75840
box 70 -56 4140 490
use wordline_driver  wordline_driver_65
timestamp 1624494425
transform 1 0 0 0 1 75050
box 70 -56 4140 490
use contact_7  contact_7_64
timestamp 1624494425
transform 1 0 74 0 1 75616
box 0 0 58 66
use contact_8  contact_8_64
timestamp 1624494425
transform 1 0 71 0 1 75617
box 0 0 64 64
use wordline_driver  wordline_driver_63
timestamp 1624494425
transform 1 0 0 0 1 75840
box 70 -56 4140 490
use contact_7  contact_7_63
timestamp 1624494425
transform 1 0 74 0 1 75998
box 0 0 58 66
use contact_8  contact_8_63
timestamp 1624494425
transform 1 0 71 0 1 75999
box 0 0 64 64
use contact_7  contact_7_62
timestamp 1624494425
transform 1 0 74 0 1 76406
box 0 0 58 66
use contact_8  contact_8_62
timestamp 1624494425
transform 1 0 71 0 1 76407
box 0 0 64 64
use wordline_driver  wordline_driver_62
timestamp 1624494425
transform 1 0 0 0 -1 76630
box 70 -56 4140 490
use contact_7  contact_7_61
timestamp 1624494425
transform 1 0 74 0 1 76788
box 0 0 58 66
use contact_8  contact_8_61
timestamp 1624494425
transform 1 0 71 0 1 76789
box 0 0 64 64
use wordline_driver  wordline_driver_60
timestamp 1624494425
transform 1 0 0 0 -1 77420
box 70 -56 4140 490
use wordline_driver  wordline_driver_61
timestamp 1624494425
transform 1 0 0 0 1 76630
box 70 -56 4140 490
use contact_7  contact_7_60
timestamp 1624494425
transform 1 0 74 0 1 77196
box 0 0 58 66
use contact_8  contact_8_60
timestamp 1624494425
transform 1 0 71 0 1 77197
box 0 0 64 64
use contact_7  contact_7_59
timestamp 1624494425
transform 1 0 74 0 1 77578
box 0 0 58 66
use contact_8  contact_8_59
timestamp 1624494425
transform 1 0 71 0 1 77579
box 0 0 64 64
use wordline_driver  wordline_driver_59
timestamp 1624494425
transform 1 0 0 0 1 77420
box 70 -56 4140 490
use contact_7  contact_7_58
timestamp 1624494425
transform 1 0 74 0 1 77986
box 0 0 58 66
use contact_8  contact_8_58
timestamp 1624494425
transform 1 0 71 0 1 77987
box 0 0 64 64
use wordline_driver  wordline_driver_57
timestamp 1624494425
transform 1 0 0 0 1 78210
box 70 -56 4140 490
use wordline_driver  wordline_driver_58
timestamp 1624494425
transform 1 0 0 0 -1 78210
box 70 -56 4140 490
use contact_7  contact_7_57
timestamp 1624494425
transform 1 0 74 0 1 78368
box 0 0 58 66
use contact_8  contact_8_57
timestamp 1624494425
transform 1 0 71 0 1 78369
box 0 0 64 64
use wordline_driver  wordline_driver_56
timestamp 1624494425
transform 1 0 0 0 -1 79000
box 70 -56 4140 490
use contact_7  contact_7_56
timestamp 1624494425
transform 1 0 74 0 1 78776
box 0 0 58 66
use contact_8  contact_8_56
timestamp 1624494425
transform 1 0 71 0 1 78777
box 0 0 64 64
use contact_7  contact_7_55
timestamp 1624494425
transform 1 0 74 0 1 79158
box 0 0 58 66
use contact_8  contact_8_55
timestamp 1624494425
transform 1 0 71 0 1 79159
box 0 0 64 64
use wordline_driver  wordline_driver_55
timestamp 1624494425
transform 1 0 0 0 1 79000
box 70 -56 4140 490
use contact_7  contact_7_54
timestamp 1624494425
transform 1 0 74 0 1 79566
box 0 0 58 66
use contact_8  contact_8_54
timestamp 1624494425
transform 1 0 71 0 1 79567
box 0 0 64 64
use wordline_driver  wordline_driver_53
timestamp 1624494425
transform 1 0 0 0 1 79790
box 70 -56 4140 490
use wordline_driver  wordline_driver_54
timestamp 1624494425
transform 1 0 0 0 -1 79790
box 70 -56 4140 490
use contact_7  contact_7_53
timestamp 1624494425
transform 1 0 74 0 1 79948
box 0 0 58 66
use contact_8  contact_8_53
timestamp 1624494425
transform 1 0 71 0 1 79949
box 0 0 64 64
use wordline_driver  wordline_driver_52
timestamp 1624494425
transform 1 0 0 0 -1 80580
box 70 -56 4140 490
use contact_7  contact_7_52
timestamp 1624494425
transform 1 0 74 0 1 80356
box 0 0 58 66
use contact_8  contact_8_52
timestamp 1624494425
transform 1 0 71 0 1 80357
box 0 0 64 64
use contact_7  contact_7_51
timestamp 1624494425
transform 1 0 74 0 1 80738
box 0 0 58 66
use contact_8  contact_8_51
timestamp 1624494425
transform 1 0 71 0 1 80739
box 0 0 64 64
use wordline_driver  wordline_driver_50
timestamp 1624494425
transform 1 0 0 0 -1 81370
box 70 -56 4140 490
use wordline_driver  wordline_driver_51
timestamp 1624494425
transform 1 0 0 0 1 80580
box 70 -56 4140 490
use contact_7  contact_7_50
timestamp 1624494425
transform 1 0 74 0 1 81146
box 0 0 58 66
use contact_8  contact_8_50
timestamp 1624494425
transform 1 0 71 0 1 81147
box 0 0 64 64
use wordline_driver  wordline_driver_49
timestamp 1624494425
transform 1 0 0 0 1 81370
box 70 -56 4140 490
use contact_7  contact_7_49
timestamp 1624494425
transform 1 0 74 0 1 81528
box 0 0 58 66
use contact_8  contact_8_49
timestamp 1624494425
transform 1 0 71 0 1 81529
box 0 0 64 64
use contact_7  contact_7_48
timestamp 1624494425
transform 1 0 74 0 1 81936
box 0 0 58 66
use contact_8  contact_8_48
timestamp 1624494425
transform 1 0 71 0 1 81937
box 0 0 64 64
use wordline_driver  wordline_driver_48
timestamp 1624494425
transform 1 0 0 0 -1 82160
box 70 -56 4140 490
use contact_7  contact_7_47
timestamp 1624494425
transform 1 0 74 0 1 82318
box 0 0 58 66
use contact_8  contact_8_47
timestamp 1624494425
transform 1 0 71 0 1 82319
box 0 0 64 64
use wordline_driver  wordline_driver_46
timestamp 1624494425
transform 1 0 0 0 -1 82950
box 70 -56 4140 490
use wordline_driver  wordline_driver_47
timestamp 1624494425
transform 1 0 0 0 1 82160
box 70 -56 4140 490
use contact_7  contact_7_46
timestamp 1624494425
transform 1 0 74 0 1 82726
box 0 0 58 66
use contact_8  contact_8_46
timestamp 1624494425
transform 1 0 71 0 1 82727
box 0 0 64 64
use wordline_driver  wordline_driver_45
timestamp 1624494425
transform 1 0 0 0 1 82950
box 70 -56 4140 490
use contact_7  contact_7_45
timestamp 1624494425
transform 1 0 74 0 1 83108
box 0 0 58 66
use contact_8  contact_8_45
timestamp 1624494425
transform 1 0 71 0 1 83109
box 0 0 64 64
use contact_7  contact_7_44
timestamp 1624494425
transform 1 0 74 0 1 83516
box 0 0 58 66
use contact_8  contact_8_44
timestamp 1624494425
transform 1 0 71 0 1 83517
box 0 0 64 64
use wordline_driver  wordline_driver_44
timestamp 1624494425
transform 1 0 0 0 -1 83740
box 70 -56 4140 490
use contact_7  contact_7_43
timestamp 1624494425
transform 1 0 74 0 1 83898
box 0 0 58 66
use contact_8  contact_8_43
timestamp 1624494425
transform 1 0 71 0 1 83899
box 0 0 64 64
use wordline_driver  wordline_driver_42
timestamp 1624494425
transform 1 0 0 0 -1 84530
box 70 -56 4140 490
use wordline_driver  wordline_driver_43
timestamp 1624494425
transform 1 0 0 0 1 83740
box 70 -56 4140 490
use contact_7  contact_7_42
timestamp 1624494425
transform 1 0 74 0 1 84306
box 0 0 58 66
use contact_8  contact_8_42
timestamp 1624494425
transform 1 0 71 0 1 84307
box 0 0 64 64
use contact_7  contact_7_41
timestamp 1624494425
transform 1 0 74 0 1 84688
box 0 0 58 66
use contact_8  contact_8_41
timestamp 1624494425
transform 1 0 71 0 1 84689
box 0 0 64 64
use wordline_driver  wordline_driver_41
timestamp 1624494425
transform 1 0 0 0 1 84530
box 70 -56 4140 490
use contact_7  contact_7_40
timestamp 1624494425
transform 1 0 74 0 1 85096
box 0 0 58 66
use contact_8  contact_8_40
timestamp 1624494425
transform 1 0 71 0 1 85097
box 0 0 64 64
use wordline_driver  wordline_driver_39
timestamp 1624494425
transform 1 0 0 0 1 85320
box 70 -56 4140 490
use wordline_driver  wordline_driver_40
timestamp 1624494425
transform 1 0 0 0 -1 85320
box 70 -56 4140 490
use contact_7  contact_7_39
timestamp 1624494425
transform 1 0 74 0 1 85478
box 0 0 58 66
use contact_8  contact_8_39
timestamp 1624494425
transform 1 0 71 0 1 85479
box 0 0 64 64
use wordline_driver  wordline_driver_38
timestamp 1624494425
transform 1 0 0 0 -1 86110
box 70 -56 4140 490
use contact_7  contact_7_38
timestamp 1624494425
transform 1 0 74 0 1 85886
box 0 0 58 66
use contact_8  contact_8_38
timestamp 1624494425
transform 1 0 71 0 1 85887
box 0 0 64 64
use contact_7  contact_7_37
timestamp 1624494425
transform 1 0 74 0 1 86268
box 0 0 58 66
use contact_8  contact_8_37
timestamp 1624494425
transform 1 0 71 0 1 86269
box 0 0 64 64
use wordline_driver  wordline_driver_37
timestamp 1624494425
transform 1 0 0 0 1 86110
box 70 -56 4140 490
use contact_7  contact_7_36
timestamp 1624494425
transform 1 0 74 0 1 86676
box 0 0 58 66
use contact_8  contact_8_36
timestamp 1624494425
transform 1 0 71 0 1 86677
box 0 0 64 64
use wordline_driver  wordline_driver_35
timestamp 1624494425
transform 1 0 0 0 1 86900
box 70 -56 4140 490
use wordline_driver  wordline_driver_36
timestamp 1624494425
transform 1 0 0 0 -1 86900
box 70 -56 4140 490
use contact_7  contact_7_35
timestamp 1624494425
transform 1 0 74 0 1 87058
box 0 0 58 66
use contact_8  contact_8_35
timestamp 1624494425
transform 1 0 71 0 1 87059
box 0 0 64 64
use wordline_driver  wordline_driver_34
timestamp 1624494425
transform 1 0 0 0 -1 87690
box 70 -56 4140 490
use contact_7  contact_7_34
timestamp 1624494425
transform 1 0 74 0 1 87466
box 0 0 58 66
use contact_8  contact_8_34
timestamp 1624494425
transform 1 0 71 0 1 87467
box 0 0 64 64
use contact_7  contact_7_33
timestamp 1624494425
transform 1 0 74 0 1 87848
box 0 0 58 66
use contact_8  contact_8_33
timestamp 1624494425
transform 1 0 71 0 1 87849
box 0 0 64 64
use wordline_driver  wordline_driver_32
timestamp 1624494425
transform 1 0 0 0 -1 88480
box 70 -56 4140 490
use wordline_driver  wordline_driver_33
timestamp 1624494425
transform 1 0 0 0 1 87690
box 70 -56 4140 490
use contact_7  contact_7_32
timestamp 1624494425
transform 1 0 74 0 1 88256
box 0 0 58 66
use contact_8  contact_8_32
timestamp 1624494425
transform 1 0 71 0 1 88257
box 0 0 64 64
use wordline_driver  wordline_driver_31
timestamp 1624494425
transform 1 0 0 0 1 88480
box 70 -56 4140 490
use contact_7  contact_7_31
timestamp 1624494425
transform 1 0 74 0 1 88638
box 0 0 58 66
use contact_8  contact_8_31
timestamp 1624494425
transform 1 0 71 0 1 88639
box 0 0 64 64
use contact_7  contact_7_30
timestamp 1624494425
transform 1 0 74 0 1 89046
box 0 0 58 66
use contact_8  contact_8_30
timestamp 1624494425
transform 1 0 71 0 1 89047
box 0 0 64 64
use wordline_driver  wordline_driver_30
timestamp 1624494425
transform 1 0 0 0 -1 89270
box 70 -56 4140 490
use contact_7  contact_7_29
timestamp 1624494425
transform 1 0 74 0 1 89428
box 0 0 58 66
use contact_8  contact_8_29
timestamp 1624494425
transform 1 0 71 0 1 89429
box 0 0 64 64
use wordline_driver  wordline_driver_28
timestamp 1624494425
transform 1 0 0 0 -1 90060
box 70 -56 4140 490
use wordline_driver  wordline_driver_29
timestamp 1624494425
transform 1 0 0 0 1 89270
box 70 -56 4140 490
use contact_7  contact_7_28
timestamp 1624494425
transform 1 0 74 0 1 89836
box 0 0 58 66
use contact_8  contact_8_28
timestamp 1624494425
transform 1 0 71 0 1 89837
box 0 0 64 64
use wordline_driver  wordline_driver_27
timestamp 1624494425
transform 1 0 0 0 1 90060
box 70 -56 4140 490
use contact_7  contact_7_27
timestamp 1624494425
transform 1 0 74 0 1 90218
box 0 0 58 66
use contact_8  contact_8_27
timestamp 1624494425
transform 1 0 71 0 1 90219
box 0 0 64 64
use contact_7  contact_7_26
timestamp 1624494425
transform 1 0 74 0 1 90626
box 0 0 58 66
use contact_8  contact_8_26
timestamp 1624494425
transform 1 0 71 0 1 90627
box 0 0 64 64
use wordline_driver  wordline_driver_26
timestamp 1624494425
transform 1 0 0 0 -1 90850
box 70 -56 4140 490
use contact_7  contact_7_25
timestamp 1624494425
transform 1 0 74 0 1 91008
box 0 0 58 66
use contact_8  contact_8_25
timestamp 1624494425
transform 1 0 71 0 1 91009
box 0 0 64 64
use wordline_driver  wordline_driver_24
timestamp 1624494425
transform 1 0 0 0 -1 91640
box 70 -56 4140 490
use wordline_driver  wordline_driver_25
timestamp 1624494425
transform 1 0 0 0 1 90850
box 70 -56 4140 490
use contact_7  contact_7_24
timestamp 1624494425
transform 1 0 74 0 1 91416
box 0 0 58 66
use contact_8  contact_8_24
timestamp 1624494425
transform 1 0 71 0 1 91417
box 0 0 64 64
use contact_7  contact_7_23
timestamp 1624494425
transform 1 0 74 0 1 91798
box 0 0 58 66
use contact_8  contact_8_23
timestamp 1624494425
transform 1 0 71 0 1 91799
box 0 0 64 64
use wordline_driver  wordline_driver_23
timestamp 1624494425
transform 1 0 0 0 1 91640
box 70 -56 4140 490
use contact_7  contact_7_22
timestamp 1624494425
transform 1 0 74 0 1 92206
box 0 0 58 66
use contact_8  contact_8_22
timestamp 1624494425
transform 1 0 71 0 1 92207
box 0 0 64 64
use wordline_driver  wordline_driver_21
timestamp 1624494425
transform 1 0 0 0 1 92430
box 70 -56 4140 490
use wordline_driver  wordline_driver_22
timestamp 1624494425
transform 1 0 0 0 -1 92430
box 70 -56 4140 490
use contact_7  contact_7_21
timestamp 1624494425
transform 1 0 74 0 1 92588
box 0 0 58 66
use contact_8  contact_8_21
timestamp 1624494425
transform 1 0 71 0 1 92589
box 0 0 64 64
use wordline_driver  wordline_driver_20
timestamp 1624494425
transform 1 0 0 0 -1 93220
box 70 -56 4140 490
use contact_7  contact_7_20
timestamp 1624494425
transform 1 0 74 0 1 92996
box 0 0 58 66
use contact_8  contact_8_20
timestamp 1624494425
transform 1 0 71 0 1 92997
box 0 0 64 64
use contact_7  contact_7_19
timestamp 1624494425
transform 1 0 74 0 1 93378
box 0 0 58 66
use contact_8  contact_8_19
timestamp 1624494425
transform 1 0 71 0 1 93379
box 0 0 64 64
use wordline_driver  wordline_driver_19
timestamp 1624494425
transform 1 0 0 0 1 93220
box 70 -56 4140 490
use contact_7  contact_7_18
timestamp 1624494425
transform 1 0 74 0 1 93786
box 0 0 58 66
use contact_8  contact_8_18
timestamp 1624494425
transform 1 0 71 0 1 93787
box 0 0 64 64
use wordline_driver  wordline_driver_17
timestamp 1624494425
transform 1 0 0 0 1 94010
box 70 -56 4140 490
use wordline_driver  wordline_driver_18
timestamp 1624494425
transform 1 0 0 0 -1 94010
box 70 -56 4140 490
use contact_7  contact_7_17
timestamp 1624494425
transform 1 0 74 0 1 94168
box 0 0 58 66
use contact_8  contact_8_17
timestamp 1624494425
transform 1 0 71 0 1 94169
box 0 0 64 64
use wordline_driver  wordline_driver_16
timestamp 1624494425
transform 1 0 0 0 -1 94800
box 70 -56 4140 490
use contact_7  contact_7_16
timestamp 1624494425
transform 1 0 74 0 1 94576
box 0 0 58 66
use contact_8  contact_8_16
timestamp 1624494425
transform 1 0 71 0 1 94577
box 0 0 64 64
use contact_7  contact_7_15
timestamp 1624494425
transform 1 0 74 0 1 94958
box 0 0 58 66
use contact_8  contact_8_15
timestamp 1624494425
transform 1 0 71 0 1 94959
box 0 0 64 64
use wordline_driver  wordline_driver_14
timestamp 1624494425
transform 1 0 0 0 -1 95590
box 70 -56 4140 490
use wordline_driver  wordline_driver_15
timestamp 1624494425
transform 1 0 0 0 1 94800
box 70 -56 4140 490
use contact_7  contact_7_14
timestamp 1624494425
transform 1 0 74 0 1 95366
box 0 0 58 66
use contact_8  contact_8_14
timestamp 1624494425
transform 1 0 71 0 1 95367
box 0 0 64 64
use wordline_driver  wordline_driver_13
timestamp 1624494425
transform 1 0 0 0 1 95590
box 70 -56 4140 490
use contact_7  contact_7_13
timestamp 1624494425
transform 1 0 74 0 1 95748
box 0 0 58 66
use contact_8  contact_8_13
timestamp 1624494425
transform 1 0 71 0 1 95749
box 0 0 64 64
use contact_7  contact_7_12
timestamp 1624494425
transform 1 0 74 0 1 96156
box 0 0 58 66
use contact_8  contact_8_12
timestamp 1624494425
transform 1 0 71 0 1 96157
box 0 0 64 64
use wordline_driver  wordline_driver_12
timestamp 1624494425
transform 1 0 0 0 -1 96380
box 70 -56 4140 490
use contact_7  contact_7_11
timestamp 1624494425
transform 1 0 74 0 1 96538
box 0 0 58 66
use contact_8  contact_8_11
timestamp 1624494425
transform 1 0 71 0 1 96539
box 0 0 64 64
use wordline_driver  wordline_driver_10
timestamp 1624494425
transform 1 0 0 0 -1 97170
box 70 -56 4140 490
use wordline_driver  wordline_driver_11
timestamp 1624494425
transform 1 0 0 0 1 96380
box 70 -56 4140 490
use contact_7  contact_7_10
timestamp 1624494425
transform 1 0 74 0 1 96946
box 0 0 58 66
use contact_8  contact_8_10
timestamp 1624494425
transform 1 0 71 0 1 96947
box 0 0 64 64
use wordline_driver  wordline_driver_9
timestamp 1624494425
transform 1 0 0 0 1 97170
box 70 -56 4140 490
use contact_7  contact_7_9
timestamp 1624494425
transform 1 0 74 0 1 97328
box 0 0 58 66
use contact_8  contact_8_9
timestamp 1624494425
transform 1 0 71 0 1 97329
box 0 0 64 64
use contact_7  contact_7_8
timestamp 1624494425
transform 1 0 74 0 1 97736
box 0 0 58 66
use contact_8  contact_8_8
timestamp 1624494425
transform 1 0 71 0 1 97737
box 0 0 64 64
use wordline_driver  wordline_driver_8
timestamp 1624494425
transform 1 0 0 0 -1 97960
box 70 -56 4140 490
use contact_7  contact_7_7
timestamp 1624494425
transform 1 0 74 0 1 98118
box 0 0 58 66
use contact_8  contact_8_7
timestamp 1624494425
transform 1 0 71 0 1 98119
box 0 0 64 64
use wordline_driver  wordline_driver_6
timestamp 1624494425
transform 1 0 0 0 -1 98750
box 70 -56 4140 490
use wordline_driver  wordline_driver_7
timestamp 1624494425
transform 1 0 0 0 1 97960
box 70 -56 4140 490
use contact_7  contact_7_6
timestamp 1624494425
transform 1 0 74 0 1 98526
box 0 0 58 66
use contact_8  contact_8_6
timestamp 1624494425
transform 1 0 71 0 1 98527
box 0 0 64 64
use contact_7  contact_7_5
timestamp 1624494425
transform 1 0 74 0 1 98908
box 0 0 58 66
use contact_8  contact_8_5
timestamp 1624494425
transform 1 0 71 0 1 98909
box 0 0 64 64
use wordline_driver  wordline_driver_5
timestamp 1624494425
transform 1 0 0 0 1 98750
box 70 -56 4140 490
use contact_7  contact_7_4
timestamp 1624494425
transform 1 0 74 0 1 99316
box 0 0 58 66
use contact_8  contact_8_4
timestamp 1624494425
transform 1 0 71 0 1 99317
box 0 0 64 64
use wordline_driver  wordline_driver_3
timestamp 1624494425
transform 1 0 0 0 1 99540
box 70 -56 4140 490
use wordline_driver  wordline_driver_4
timestamp 1624494425
transform 1 0 0 0 -1 99540
box 70 -56 4140 490
use contact_7  contact_7_3
timestamp 1624494425
transform 1 0 74 0 1 99698
box 0 0 58 66
use contact_8  contact_8_3
timestamp 1624494425
transform 1 0 71 0 1 99699
box 0 0 64 64
use wordline_driver  wordline_driver_2
timestamp 1624494425
transform 1 0 0 0 -1 100330
box 70 -56 4140 490
use contact_7  contact_7_2
timestamp 1624494425
transform 1 0 74 0 1 100106
box 0 0 58 66
use contact_8  contact_8_2
timestamp 1624494425
transform 1 0 71 0 1 100107
box 0 0 64 64
use contact_7  contact_7_1
timestamp 1624494425
transform 1 0 74 0 1 100488
box 0 0 58 66
use contact_8  contact_8_1
timestamp 1624494425
transform 1 0 71 0 1 100489
box 0 0 64 64
use wordline_driver  wordline_driver_1
timestamp 1624494425
transform 1 0 0 0 1 100330
box 70 -56 4140 490
use contact_7  contact_7_0
timestamp 1624494425
transform 1 0 74 0 1 100896
box 0 0 58 66
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 71 0 1 100897
box 0 0 64 64
use wordline_driver  wordline_driver_0
timestamp 1624494425
transform 1 0 0 0 -1 101120
box 70 -56 4140 490
<< labels >>
rlabel metal2 s 70 0 98 101120 4 en
rlabel locali s 103 299 103 299 4 in_0
rlabel locali s 4108 120 4108 120 4 wl_0
rlabel locali s 103 491 103 491 4 in_1
rlabel locali s 4108 670 4108 670 4 wl_1
rlabel locali s 103 1089 103 1089 4 in_2
rlabel locali s 4108 910 4108 910 4 wl_2
rlabel locali s 103 1281 103 1281 4 in_3
rlabel locali s 4108 1460 4108 1460 4 wl_3
rlabel locali s 103 1879 103 1879 4 in_4
rlabel locali s 4108 1700 4108 1700 4 wl_4
rlabel locali s 103 2071 103 2071 4 in_5
rlabel locali s 4108 2250 4108 2250 4 wl_5
rlabel locali s 103 2669 103 2669 4 in_6
rlabel locali s 4108 2490 4108 2490 4 wl_6
rlabel locali s 103 2861 103 2861 4 in_7
rlabel locali s 4108 3040 4108 3040 4 wl_7
rlabel locali s 103 3459 103 3459 4 in_8
rlabel locali s 4108 3280 4108 3280 4 wl_8
rlabel locali s 103 3651 103 3651 4 in_9
rlabel locali s 4108 3830 4108 3830 4 wl_9
rlabel locali s 103 4249 103 4249 4 in_10
rlabel locali s 4108 4070 4108 4070 4 wl_10
rlabel locali s 103 4441 103 4441 4 in_11
rlabel locali s 4108 4620 4108 4620 4 wl_11
rlabel locali s 103 5039 103 5039 4 in_12
rlabel locali s 4108 4860 4108 4860 4 wl_12
rlabel locali s 103 5231 103 5231 4 in_13
rlabel locali s 4108 5410 4108 5410 4 wl_13
rlabel locali s 103 5829 103 5829 4 in_14
rlabel locali s 4108 5650 4108 5650 4 wl_14
rlabel locali s 103 6021 103 6021 4 in_15
rlabel locali s 4108 6200 4108 6200 4 wl_15
rlabel locali s 103 6619 103 6619 4 in_16
rlabel locali s 4108 6440 4108 6440 4 wl_16
rlabel locali s 103 6811 103 6811 4 in_17
rlabel locali s 4108 6990 4108 6990 4 wl_17
rlabel locali s 103 7409 103 7409 4 in_18
rlabel locali s 4108 7230 4108 7230 4 wl_18
rlabel locali s 103 7601 103 7601 4 in_19
rlabel locali s 4108 7780 4108 7780 4 wl_19
rlabel locali s 103 8199 103 8199 4 in_20
rlabel locali s 4108 8020 4108 8020 4 wl_20
rlabel locali s 103 8391 103 8391 4 in_21
rlabel locali s 4108 8570 4108 8570 4 wl_21
rlabel locali s 103 8989 103 8989 4 in_22
rlabel locali s 4108 8810 4108 8810 4 wl_22
rlabel locali s 103 9181 103 9181 4 in_23
rlabel locali s 4108 9360 4108 9360 4 wl_23
rlabel locali s 103 9779 103 9779 4 in_24
rlabel locali s 4108 9600 4108 9600 4 wl_24
rlabel locali s 103 9971 103 9971 4 in_25
rlabel locali s 4108 10150 4108 10150 4 wl_25
rlabel locali s 103 10569 103 10569 4 in_26
rlabel locali s 4108 10390 4108 10390 4 wl_26
rlabel locali s 103 10761 103 10761 4 in_27
rlabel locali s 4108 10940 4108 10940 4 wl_27
rlabel locali s 103 11359 103 11359 4 in_28
rlabel locali s 4108 11180 4108 11180 4 wl_28
rlabel locali s 103 11551 103 11551 4 in_29
rlabel locali s 4108 11730 4108 11730 4 wl_29
rlabel locali s 103 12149 103 12149 4 in_30
rlabel locali s 4108 11970 4108 11970 4 wl_30
rlabel locali s 103 12341 103 12341 4 in_31
rlabel locali s 4108 12520 4108 12520 4 wl_31
rlabel locali s 103 12939 103 12939 4 in_32
rlabel locali s 4108 12760 4108 12760 4 wl_32
rlabel locali s 103 13131 103 13131 4 in_33
rlabel locali s 4108 13310 4108 13310 4 wl_33
rlabel locali s 103 13729 103 13729 4 in_34
rlabel locali s 4108 13550 4108 13550 4 wl_34
rlabel locali s 103 13921 103 13921 4 in_35
rlabel locali s 4108 14100 4108 14100 4 wl_35
rlabel locali s 103 14519 103 14519 4 in_36
rlabel locali s 4108 14340 4108 14340 4 wl_36
rlabel locali s 103 14711 103 14711 4 in_37
rlabel locali s 4108 14890 4108 14890 4 wl_37
rlabel locali s 103 15309 103 15309 4 in_38
rlabel locali s 4108 15130 4108 15130 4 wl_38
rlabel locali s 103 15501 103 15501 4 in_39
rlabel locali s 4108 15680 4108 15680 4 wl_39
rlabel locali s 103 16099 103 16099 4 in_40
rlabel locali s 4108 15920 4108 15920 4 wl_40
rlabel locali s 103 16291 103 16291 4 in_41
rlabel locali s 4108 16470 4108 16470 4 wl_41
rlabel locali s 103 16889 103 16889 4 in_42
rlabel locali s 4108 16710 4108 16710 4 wl_42
rlabel locali s 103 17081 103 17081 4 in_43
rlabel locali s 4108 17260 4108 17260 4 wl_43
rlabel locali s 103 17679 103 17679 4 in_44
rlabel locali s 4108 17500 4108 17500 4 wl_44
rlabel locali s 103 17871 103 17871 4 in_45
rlabel locali s 4108 18050 4108 18050 4 wl_45
rlabel locali s 103 18469 103 18469 4 in_46
rlabel locali s 4108 18290 4108 18290 4 wl_46
rlabel locali s 103 18661 103 18661 4 in_47
rlabel locali s 4108 18840 4108 18840 4 wl_47
rlabel locali s 103 19259 103 19259 4 in_48
rlabel locali s 4108 19080 4108 19080 4 wl_48
rlabel locali s 103 19451 103 19451 4 in_49
rlabel locali s 4108 19630 4108 19630 4 wl_49
rlabel locali s 103 20049 103 20049 4 in_50
rlabel locali s 4108 19870 4108 19870 4 wl_50
rlabel locali s 103 20241 103 20241 4 in_51
rlabel locali s 4108 20420 4108 20420 4 wl_51
rlabel locali s 103 20839 103 20839 4 in_52
rlabel locali s 4108 20660 4108 20660 4 wl_52
rlabel locali s 103 21031 103 21031 4 in_53
rlabel locali s 4108 21210 4108 21210 4 wl_53
rlabel locali s 103 21629 103 21629 4 in_54
rlabel locali s 4108 21450 4108 21450 4 wl_54
rlabel locali s 103 21821 103 21821 4 in_55
rlabel locali s 4108 22000 4108 22000 4 wl_55
rlabel locali s 103 22419 103 22419 4 in_56
rlabel locali s 4108 22240 4108 22240 4 wl_56
rlabel locali s 103 22611 103 22611 4 in_57
rlabel locali s 4108 22790 4108 22790 4 wl_57
rlabel locali s 103 23209 103 23209 4 in_58
rlabel locali s 4108 23030 4108 23030 4 wl_58
rlabel locali s 103 23401 103 23401 4 in_59
rlabel locali s 4108 23580 4108 23580 4 wl_59
rlabel locali s 103 23999 103 23999 4 in_60
rlabel locali s 4108 23820 4108 23820 4 wl_60
rlabel locali s 103 24191 103 24191 4 in_61
rlabel locali s 4108 24370 4108 24370 4 wl_61
rlabel locali s 103 24789 103 24789 4 in_62
rlabel locali s 4108 24610 4108 24610 4 wl_62
rlabel locali s 103 24981 103 24981 4 in_63
rlabel locali s 4108 25160 4108 25160 4 wl_63
rlabel locali s 103 25579 103 25579 4 in_64
rlabel locali s 4108 25400 4108 25400 4 wl_64
rlabel locali s 103 25771 103 25771 4 in_65
rlabel locali s 4108 25950 4108 25950 4 wl_65
rlabel locali s 103 26369 103 26369 4 in_66
rlabel locali s 4108 26190 4108 26190 4 wl_66
rlabel locali s 103 26561 103 26561 4 in_67
rlabel locali s 4108 26740 4108 26740 4 wl_67
rlabel locali s 103 27159 103 27159 4 in_68
rlabel locali s 4108 26980 4108 26980 4 wl_68
rlabel locali s 103 27351 103 27351 4 in_69
rlabel locali s 4108 27530 4108 27530 4 wl_69
rlabel locali s 103 27949 103 27949 4 in_70
rlabel locali s 4108 27770 4108 27770 4 wl_70
rlabel locali s 103 28141 103 28141 4 in_71
rlabel locali s 4108 28320 4108 28320 4 wl_71
rlabel locali s 103 28739 103 28739 4 in_72
rlabel locali s 4108 28560 4108 28560 4 wl_72
rlabel locali s 103 28931 103 28931 4 in_73
rlabel locali s 4108 29110 4108 29110 4 wl_73
rlabel locali s 103 29529 103 29529 4 in_74
rlabel locali s 4108 29350 4108 29350 4 wl_74
rlabel locali s 103 29721 103 29721 4 in_75
rlabel locali s 4108 29900 4108 29900 4 wl_75
rlabel locali s 103 30319 103 30319 4 in_76
rlabel locali s 4108 30140 4108 30140 4 wl_76
rlabel locali s 103 30511 103 30511 4 in_77
rlabel locali s 4108 30690 4108 30690 4 wl_77
rlabel locali s 103 31109 103 31109 4 in_78
rlabel locali s 4108 30930 4108 30930 4 wl_78
rlabel locali s 103 31301 103 31301 4 in_79
rlabel locali s 4108 31480 4108 31480 4 wl_79
rlabel locali s 103 31899 103 31899 4 in_80
rlabel locali s 4108 31720 4108 31720 4 wl_80
rlabel locali s 103 32091 103 32091 4 in_81
rlabel locali s 4108 32270 4108 32270 4 wl_81
rlabel locali s 103 32689 103 32689 4 in_82
rlabel locali s 4108 32510 4108 32510 4 wl_82
rlabel locali s 103 32881 103 32881 4 in_83
rlabel locali s 4108 33060 4108 33060 4 wl_83
rlabel locali s 103 33479 103 33479 4 in_84
rlabel locali s 4108 33300 4108 33300 4 wl_84
rlabel locali s 103 33671 103 33671 4 in_85
rlabel locali s 4108 33850 4108 33850 4 wl_85
rlabel locali s 103 34269 103 34269 4 in_86
rlabel locali s 4108 34090 4108 34090 4 wl_86
rlabel locali s 103 34461 103 34461 4 in_87
rlabel locali s 4108 34640 4108 34640 4 wl_87
rlabel locali s 103 35059 103 35059 4 in_88
rlabel locali s 4108 34880 4108 34880 4 wl_88
rlabel locali s 103 35251 103 35251 4 in_89
rlabel locali s 4108 35430 4108 35430 4 wl_89
rlabel locali s 103 35849 103 35849 4 in_90
rlabel locali s 4108 35670 4108 35670 4 wl_90
rlabel locali s 103 36041 103 36041 4 in_91
rlabel locali s 4108 36220 4108 36220 4 wl_91
rlabel locali s 103 36639 103 36639 4 in_92
rlabel locali s 4108 36460 4108 36460 4 wl_92
rlabel locali s 103 36831 103 36831 4 in_93
rlabel locali s 4108 37010 4108 37010 4 wl_93
rlabel locali s 103 37429 103 37429 4 in_94
rlabel locali s 4108 37250 4108 37250 4 wl_94
rlabel locali s 103 37621 103 37621 4 in_95
rlabel locali s 4108 37800 4108 37800 4 wl_95
rlabel locali s 103 38219 103 38219 4 in_96
rlabel locali s 4108 38040 4108 38040 4 wl_96
rlabel locali s 103 38411 103 38411 4 in_97
rlabel locali s 4108 38590 4108 38590 4 wl_97
rlabel locali s 103 39009 103 39009 4 in_98
rlabel locali s 4108 38830 4108 38830 4 wl_98
rlabel locali s 103 39201 103 39201 4 in_99
rlabel locali s 4108 39380 4108 39380 4 wl_99
rlabel locali s 103 39799 103 39799 4 in_100
rlabel locali s 4108 39620 4108 39620 4 wl_100
rlabel locali s 103 39991 103 39991 4 in_101
rlabel locali s 4108 40170 4108 40170 4 wl_101
rlabel locali s 103 40589 103 40589 4 in_102
rlabel locali s 4108 40410 4108 40410 4 wl_102
rlabel locali s 103 40781 103 40781 4 in_103
rlabel locali s 4108 40960 4108 40960 4 wl_103
rlabel locali s 103 41379 103 41379 4 in_104
rlabel locali s 4108 41200 4108 41200 4 wl_104
rlabel locali s 103 41571 103 41571 4 in_105
rlabel locali s 4108 41750 4108 41750 4 wl_105
rlabel locali s 103 42169 103 42169 4 in_106
rlabel locali s 4108 41990 4108 41990 4 wl_106
rlabel locali s 103 42361 103 42361 4 in_107
rlabel locali s 4108 42540 4108 42540 4 wl_107
rlabel locali s 103 42959 103 42959 4 in_108
rlabel locali s 4108 42780 4108 42780 4 wl_108
rlabel locali s 103 43151 103 43151 4 in_109
rlabel locali s 4108 43330 4108 43330 4 wl_109
rlabel locali s 103 43749 103 43749 4 in_110
rlabel locali s 4108 43570 4108 43570 4 wl_110
rlabel locali s 103 43941 103 43941 4 in_111
rlabel locali s 4108 44120 4108 44120 4 wl_111
rlabel locali s 103 44539 103 44539 4 in_112
rlabel locali s 4108 44360 4108 44360 4 wl_112
rlabel locali s 103 44731 103 44731 4 in_113
rlabel locali s 4108 44910 4108 44910 4 wl_113
rlabel locali s 103 45329 103 45329 4 in_114
rlabel locali s 4108 45150 4108 45150 4 wl_114
rlabel locali s 103 45521 103 45521 4 in_115
rlabel locali s 4108 45700 4108 45700 4 wl_115
rlabel locali s 103 46119 103 46119 4 in_116
rlabel locali s 4108 45940 4108 45940 4 wl_116
rlabel locali s 103 46311 103 46311 4 in_117
rlabel locali s 4108 46490 4108 46490 4 wl_117
rlabel locali s 103 46909 103 46909 4 in_118
rlabel locali s 4108 46730 4108 46730 4 wl_118
rlabel locali s 103 47101 103 47101 4 in_119
rlabel locali s 4108 47280 4108 47280 4 wl_119
rlabel locali s 103 47699 103 47699 4 in_120
rlabel locali s 4108 47520 4108 47520 4 wl_120
rlabel locali s 103 47891 103 47891 4 in_121
rlabel locali s 4108 48070 4108 48070 4 wl_121
rlabel locali s 103 48489 103 48489 4 in_122
rlabel locali s 4108 48310 4108 48310 4 wl_122
rlabel locali s 103 48681 103 48681 4 in_123
rlabel locali s 4108 48860 4108 48860 4 wl_123
rlabel locali s 103 49279 103 49279 4 in_124
rlabel locali s 4108 49100 4108 49100 4 wl_124
rlabel locali s 103 49471 103 49471 4 in_125
rlabel locali s 4108 49650 4108 49650 4 wl_125
rlabel locali s 103 50069 103 50069 4 in_126
rlabel locali s 4108 49890 4108 49890 4 wl_126
rlabel locali s 103 50261 103 50261 4 in_127
rlabel locali s 4108 50440 4108 50440 4 wl_127
rlabel locali s 103 50859 103 50859 4 in_128
rlabel locali s 4108 50680 4108 50680 4 wl_128
rlabel locali s 103 51051 103 51051 4 in_129
rlabel locali s 4108 51230 4108 51230 4 wl_129
rlabel locali s 103 51649 103 51649 4 in_130
rlabel locali s 4108 51470 4108 51470 4 wl_130
rlabel locali s 103 51841 103 51841 4 in_131
rlabel locali s 4108 52020 4108 52020 4 wl_131
rlabel locali s 103 52439 103 52439 4 in_132
rlabel locali s 4108 52260 4108 52260 4 wl_132
rlabel locali s 103 52631 103 52631 4 in_133
rlabel locali s 4108 52810 4108 52810 4 wl_133
rlabel locali s 103 53229 103 53229 4 in_134
rlabel locali s 4108 53050 4108 53050 4 wl_134
rlabel locali s 103 53421 103 53421 4 in_135
rlabel locali s 4108 53600 4108 53600 4 wl_135
rlabel locali s 103 54019 103 54019 4 in_136
rlabel locali s 4108 53840 4108 53840 4 wl_136
rlabel locali s 103 54211 103 54211 4 in_137
rlabel locali s 4108 54390 4108 54390 4 wl_137
rlabel locali s 103 54809 103 54809 4 in_138
rlabel locali s 4108 54630 4108 54630 4 wl_138
rlabel locali s 103 55001 103 55001 4 in_139
rlabel locali s 4108 55180 4108 55180 4 wl_139
rlabel locali s 103 55599 103 55599 4 in_140
rlabel locali s 4108 55420 4108 55420 4 wl_140
rlabel locali s 103 55791 103 55791 4 in_141
rlabel locali s 4108 55970 4108 55970 4 wl_141
rlabel locali s 103 56389 103 56389 4 in_142
rlabel locali s 4108 56210 4108 56210 4 wl_142
rlabel locali s 103 56581 103 56581 4 in_143
rlabel locali s 4108 56760 4108 56760 4 wl_143
rlabel locali s 103 57179 103 57179 4 in_144
rlabel locali s 4108 57000 4108 57000 4 wl_144
rlabel locali s 103 57371 103 57371 4 in_145
rlabel locali s 4108 57550 4108 57550 4 wl_145
rlabel locali s 103 57969 103 57969 4 in_146
rlabel locali s 4108 57790 4108 57790 4 wl_146
rlabel locali s 103 58161 103 58161 4 in_147
rlabel locali s 4108 58340 4108 58340 4 wl_147
rlabel locali s 103 58759 103 58759 4 in_148
rlabel locali s 4108 58580 4108 58580 4 wl_148
rlabel locali s 103 58951 103 58951 4 in_149
rlabel locali s 4108 59130 4108 59130 4 wl_149
rlabel locali s 103 59549 103 59549 4 in_150
rlabel locali s 4108 59370 4108 59370 4 wl_150
rlabel locali s 103 59741 103 59741 4 in_151
rlabel locali s 4108 59920 4108 59920 4 wl_151
rlabel locali s 103 60339 103 60339 4 in_152
rlabel locali s 4108 60160 4108 60160 4 wl_152
rlabel locali s 103 60531 103 60531 4 in_153
rlabel locali s 4108 60710 4108 60710 4 wl_153
rlabel locali s 103 61129 103 61129 4 in_154
rlabel locali s 4108 60950 4108 60950 4 wl_154
rlabel locali s 103 61321 103 61321 4 in_155
rlabel locali s 4108 61500 4108 61500 4 wl_155
rlabel locali s 103 61919 103 61919 4 in_156
rlabel locali s 4108 61740 4108 61740 4 wl_156
rlabel locali s 103 62111 103 62111 4 in_157
rlabel locali s 4108 62290 4108 62290 4 wl_157
rlabel locali s 103 62709 103 62709 4 in_158
rlabel locali s 4108 62530 4108 62530 4 wl_158
rlabel locali s 103 62901 103 62901 4 in_159
rlabel locali s 4108 63080 4108 63080 4 wl_159
rlabel locali s 103 63499 103 63499 4 in_160
rlabel locali s 4108 63320 4108 63320 4 wl_160
rlabel locali s 103 63691 103 63691 4 in_161
rlabel locali s 4108 63870 4108 63870 4 wl_161
rlabel locali s 103 64289 103 64289 4 in_162
rlabel locali s 4108 64110 4108 64110 4 wl_162
rlabel locali s 103 64481 103 64481 4 in_163
rlabel locali s 4108 64660 4108 64660 4 wl_163
rlabel locali s 103 65079 103 65079 4 in_164
rlabel locali s 4108 64900 4108 64900 4 wl_164
rlabel locali s 103 65271 103 65271 4 in_165
rlabel locali s 4108 65450 4108 65450 4 wl_165
rlabel locali s 103 65869 103 65869 4 in_166
rlabel locali s 4108 65690 4108 65690 4 wl_166
rlabel locali s 103 66061 103 66061 4 in_167
rlabel locali s 4108 66240 4108 66240 4 wl_167
rlabel locali s 103 66659 103 66659 4 in_168
rlabel locali s 4108 66480 4108 66480 4 wl_168
rlabel locali s 103 66851 103 66851 4 in_169
rlabel locali s 4108 67030 4108 67030 4 wl_169
rlabel locali s 103 67449 103 67449 4 in_170
rlabel locali s 4108 67270 4108 67270 4 wl_170
rlabel locali s 103 67641 103 67641 4 in_171
rlabel locali s 4108 67820 4108 67820 4 wl_171
rlabel locali s 103 68239 103 68239 4 in_172
rlabel locali s 4108 68060 4108 68060 4 wl_172
rlabel locali s 103 68431 103 68431 4 in_173
rlabel locali s 4108 68610 4108 68610 4 wl_173
rlabel locali s 103 69029 103 69029 4 in_174
rlabel locali s 4108 68850 4108 68850 4 wl_174
rlabel locali s 103 69221 103 69221 4 in_175
rlabel locali s 4108 69400 4108 69400 4 wl_175
rlabel locali s 103 69819 103 69819 4 in_176
rlabel locali s 4108 69640 4108 69640 4 wl_176
rlabel locali s 103 70011 103 70011 4 in_177
rlabel locali s 4108 70190 4108 70190 4 wl_177
rlabel locali s 103 70609 103 70609 4 in_178
rlabel locali s 4108 70430 4108 70430 4 wl_178
rlabel locali s 103 70801 103 70801 4 in_179
rlabel locali s 4108 70980 4108 70980 4 wl_179
rlabel locali s 103 71399 103 71399 4 in_180
rlabel locali s 4108 71220 4108 71220 4 wl_180
rlabel locali s 103 71591 103 71591 4 in_181
rlabel locali s 4108 71770 4108 71770 4 wl_181
rlabel locali s 103 72189 103 72189 4 in_182
rlabel locali s 4108 72010 4108 72010 4 wl_182
rlabel locali s 103 72381 103 72381 4 in_183
rlabel locali s 4108 72560 4108 72560 4 wl_183
rlabel locali s 103 72979 103 72979 4 in_184
rlabel locali s 4108 72800 4108 72800 4 wl_184
rlabel locali s 103 73171 103 73171 4 in_185
rlabel locali s 4108 73350 4108 73350 4 wl_185
rlabel locali s 103 73769 103 73769 4 in_186
rlabel locali s 4108 73590 4108 73590 4 wl_186
rlabel locali s 103 73961 103 73961 4 in_187
rlabel locali s 4108 74140 4108 74140 4 wl_187
rlabel locali s 103 74559 103 74559 4 in_188
rlabel locali s 4108 74380 4108 74380 4 wl_188
rlabel locali s 103 74751 103 74751 4 in_189
rlabel locali s 4108 74930 4108 74930 4 wl_189
rlabel locali s 103 75349 103 75349 4 in_190
rlabel locali s 4108 75170 4108 75170 4 wl_190
rlabel locali s 103 75541 103 75541 4 in_191
rlabel locali s 4108 75720 4108 75720 4 wl_191
rlabel locali s 103 76139 103 76139 4 in_192
rlabel locali s 4108 75960 4108 75960 4 wl_192
rlabel locali s 103 76331 103 76331 4 in_193
rlabel locali s 4108 76510 4108 76510 4 wl_193
rlabel locali s 103 76929 103 76929 4 in_194
rlabel locali s 4108 76750 4108 76750 4 wl_194
rlabel locali s 103 77121 103 77121 4 in_195
rlabel locali s 4108 77300 4108 77300 4 wl_195
rlabel locali s 103 77719 103 77719 4 in_196
rlabel locali s 4108 77540 4108 77540 4 wl_196
rlabel locali s 103 77911 103 77911 4 in_197
rlabel locali s 4108 78090 4108 78090 4 wl_197
rlabel locali s 103 78509 103 78509 4 in_198
rlabel locali s 4108 78330 4108 78330 4 wl_198
rlabel locali s 103 78701 103 78701 4 in_199
rlabel locali s 4108 78880 4108 78880 4 wl_199
rlabel locali s 103 79299 103 79299 4 in_200
rlabel locali s 4108 79120 4108 79120 4 wl_200
rlabel locali s 103 79491 103 79491 4 in_201
rlabel locali s 4108 79670 4108 79670 4 wl_201
rlabel locali s 103 80089 103 80089 4 in_202
rlabel locali s 4108 79910 4108 79910 4 wl_202
rlabel locali s 103 80281 103 80281 4 in_203
rlabel locali s 4108 80460 4108 80460 4 wl_203
rlabel locali s 103 80879 103 80879 4 in_204
rlabel locali s 4108 80700 4108 80700 4 wl_204
rlabel locali s 103 81071 103 81071 4 in_205
rlabel locali s 4108 81250 4108 81250 4 wl_205
rlabel locali s 103 81669 103 81669 4 in_206
rlabel locali s 4108 81490 4108 81490 4 wl_206
rlabel locali s 103 81861 103 81861 4 in_207
rlabel locali s 4108 82040 4108 82040 4 wl_207
rlabel locali s 103 82459 103 82459 4 in_208
rlabel locali s 4108 82280 4108 82280 4 wl_208
rlabel locali s 103 82651 103 82651 4 in_209
rlabel locali s 4108 82830 4108 82830 4 wl_209
rlabel locali s 103 83249 103 83249 4 in_210
rlabel locali s 4108 83070 4108 83070 4 wl_210
rlabel locali s 103 83441 103 83441 4 in_211
rlabel locali s 4108 83620 4108 83620 4 wl_211
rlabel locali s 103 84039 103 84039 4 in_212
rlabel locali s 4108 83860 4108 83860 4 wl_212
rlabel locali s 103 84231 103 84231 4 in_213
rlabel locali s 4108 84410 4108 84410 4 wl_213
rlabel locali s 103 84829 103 84829 4 in_214
rlabel locali s 4108 84650 4108 84650 4 wl_214
rlabel locali s 103 85021 103 85021 4 in_215
rlabel locali s 4108 85200 4108 85200 4 wl_215
rlabel locali s 103 85619 103 85619 4 in_216
rlabel locali s 4108 85440 4108 85440 4 wl_216
rlabel locali s 103 85811 103 85811 4 in_217
rlabel locali s 4108 85990 4108 85990 4 wl_217
rlabel locali s 103 86409 103 86409 4 in_218
rlabel locali s 4108 86230 4108 86230 4 wl_218
rlabel locali s 103 86601 103 86601 4 in_219
rlabel locali s 4108 86780 4108 86780 4 wl_219
rlabel locali s 103 87199 103 87199 4 in_220
rlabel locali s 4108 87020 4108 87020 4 wl_220
rlabel locali s 103 87391 103 87391 4 in_221
rlabel locali s 4108 87570 4108 87570 4 wl_221
rlabel locali s 103 87989 103 87989 4 in_222
rlabel locali s 4108 87810 4108 87810 4 wl_222
rlabel locali s 103 88181 103 88181 4 in_223
rlabel locali s 4108 88360 4108 88360 4 wl_223
rlabel locali s 103 88779 103 88779 4 in_224
rlabel locali s 4108 88600 4108 88600 4 wl_224
rlabel locali s 103 88971 103 88971 4 in_225
rlabel locali s 4108 89150 4108 89150 4 wl_225
rlabel locali s 103 89569 103 89569 4 in_226
rlabel locali s 4108 89390 4108 89390 4 wl_226
rlabel locali s 103 89761 103 89761 4 in_227
rlabel locali s 4108 89940 4108 89940 4 wl_227
rlabel locali s 103 90359 103 90359 4 in_228
rlabel locali s 4108 90180 4108 90180 4 wl_228
rlabel locali s 103 90551 103 90551 4 in_229
rlabel locali s 4108 90730 4108 90730 4 wl_229
rlabel locali s 103 91149 103 91149 4 in_230
rlabel locali s 4108 90970 4108 90970 4 wl_230
rlabel locali s 103 91341 103 91341 4 in_231
rlabel locali s 4108 91520 4108 91520 4 wl_231
rlabel locali s 103 91939 103 91939 4 in_232
rlabel locali s 4108 91760 4108 91760 4 wl_232
rlabel locali s 103 92131 103 92131 4 in_233
rlabel locali s 4108 92310 4108 92310 4 wl_233
rlabel locali s 103 92729 103 92729 4 in_234
rlabel locali s 4108 92550 4108 92550 4 wl_234
rlabel locali s 103 92921 103 92921 4 in_235
rlabel locali s 4108 93100 4108 93100 4 wl_235
rlabel locali s 103 93519 103 93519 4 in_236
rlabel locali s 4108 93340 4108 93340 4 wl_236
rlabel locali s 103 93711 103 93711 4 in_237
rlabel locali s 4108 93890 4108 93890 4 wl_237
rlabel locali s 103 94309 103 94309 4 in_238
rlabel locali s 4108 94130 4108 94130 4 wl_238
rlabel locali s 103 94501 103 94501 4 in_239
rlabel locali s 4108 94680 4108 94680 4 wl_239
rlabel locali s 103 95099 103 95099 4 in_240
rlabel locali s 4108 94920 4108 94920 4 wl_240
rlabel locali s 103 95291 103 95291 4 in_241
rlabel locali s 4108 95470 4108 95470 4 wl_241
rlabel locali s 103 95889 103 95889 4 in_242
rlabel locali s 4108 95710 4108 95710 4 wl_242
rlabel locali s 103 96081 103 96081 4 in_243
rlabel locali s 4108 96260 4108 96260 4 wl_243
rlabel locali s 103 96679 103 96679 4 in_244
rlabel locali s 4108 96500 4108 96500 4 wl_244
rlabel locali s 103 96871 103 96871 4 in_245
rlabel locali s 4108 97050 4108 97050 4 wl_245
rlabel locali s 103 97469 103 97469 4 in_246
rlabel locali s 4108 97290 4108 97290 4 wl_246
rlabel locali s 103 97661 103 97661 4 in_247
rlabel locali s 4108 97840 4108 97840 4 wl_247
rlabel locali s 103 98259 103 98259 4 in_248
rlabel locali s 4108 98080 4108 98080 4 wl_248
rlabel locali s 103 98451 103 98451 4 in_249
rlabel locali s 4108 98630 4108 98630 4 wl_249
rlabel locali s 103 99049 103 99049 4 in_250
rlabel locali s 4108 98870 4108 98870 4 wl_250
rlabel locali s 103 99241 103 99241 4 in_251
rlabel locali s 4108 99420 4108 99420 4 wl_251
rlabel locali s 103 99839 103 99839 4 in_252
rlabel locali s 4108 99660 4108 99660 4 wl_252
rlabel locali s 103 100031 103 100031 4 in_253
rlabel locali s 4108 100210 4108 100210 4 wl_253
rlabel locali s 103 100629 103 100629 4 in_254
rlabel locali s 4108 100450 4108 100450 4 wl_254
rlabel locali s 103 100821 103 100821 4 in_255
rlabel locali s 4108 101000 4108 101000 4 wl_255
rlabel metal1 s 681 -32 709 101120 4 vdd
rlabel metal1 s 3372 0 3400 101120 4 vdd
rlabel metal1 s 1724 0 1752 101120 4 gnd
rlabel metal1 s 256 -30 284 101120 4 gnd
<< properties >>
string FIXED_BBOX 0 0 4158 101120
<< end >>
