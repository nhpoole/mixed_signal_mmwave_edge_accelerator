magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1190 51852 5400 51876
rect -1260 -1292 5400 51852
rect -1190 -1316 5400 -1292
<< locali >>
rect 4094 50423 4122 50457
rect 70 50244 136 50278
rect 70 50052 136 50086
rect 4094 49873 4122 49907
rect 4094 49633 4122 49667
rect 70 49454 136 49488
rect 70 49262 136 49296
rect 4094 49083 4122 49117
rect 4094 48843 4122 48877
rect 70 48664 136 48698
rect 70 48472 136 48506
rect 4094 48293 4122 48327
rect 4094 48053 4122 48087
rect 70 47874 136 47908
rect 70 47682 136 47716
rect 4094 47503 4122 47537
rect 4094 47263 4122 47297
rect 70 47084 136 47118
rect 70 46892 136 46926
rect 4094 46713 4122 46747
rect 4094 46473 4122 46507
rect 70 46294 136 46328
rect 70 46102 136 46136
rect 4094 45923 4122 45957
rect 4094 45683 4122 45717
rect 70 45504 136 45538
rect 70 45312 136 45346
rect 4094 45133 4122 45167
rect 4094 44893 4122 44927
rect 70 44714 136 44748
rect 70 44522 136 44556
rect 4094 44343 4122 44377
rect 4094 44103 4122 44137
rect 70 43924 136 43958
rect 70 43732 136 43766
rect 4094 43553 4122 43587
rect 4094 43313 4122 43347
rect 70 43134 136 43168
rect 70 42942 136 42976
rect 4094 42763 4122 42797
rect 4094 42523 4122 42557
rect 70 42344 136 42378
rect 70 42152 136 42186
rect 4094 41973 4122 42007
rect 4094 41733 4122 41767
rect 70 41554 136 41588
rect 70 41362 136 41396
rect 4094 41183 4122 41217
rect 4094 40943 4122 40977
rect 70 40764 136 40798
rect 70 40572 136 40606
rect 4094 40393 4122 40427
rect 4094 40153 4122 40187
rect 70 39974 136 40008
rect 70 39782 136 39816
rect 4094 39603 4122 39637
rect 4094 39363 4122 39397
rect 70 39184 136 39218
rect 70 38992 136 39026
rect 4094 38813 4122 38847
rect 4094 38573 4122 38607
rect 70 38394 136 38428
rect 70 38202 136 38236
rect 4094 38023 4122 38057
rect 4094 37783 4122 37817
rect 70 37604 136 37638
rect 70 37412 136 37446
rect 4094 37233 4122 37267
rect 4094 36993 4122 37027
rect 70 36814 136 36848
rect 70 36622 136 36656
rect 4094 36443 4122 36477
rect 4094 36203 4122 36237
rect 70 36024 136 36058
rect 70 35832 136 35866
rect 4094 35653 4122 35687
rect 4094 35413 4122 35447
rect 70 35234 136 35268
rect 70 35042 136 35076
rect 4094 34863 4122 34897
rect 4094 34623 4122 34657
rect 70 34444 136 34478
rect 70 34252 136 34286
rect 4094 34073 4122 34107
rect 4094 33833 4122 33867
rect 70 33654 136 33688
rect 70 33462 136 33496
rect 4094 33283 4122 33317
rect 4094 33043 4122 33077
rect 70 32864 136 32898
rect 70 32672 136 32706
rect 4094 32493 4122 32527
rect 4094 32253 4122 32287
rect 70 32074 136 32108
rect 70 31882 136 31916
rect 4094 31703 4122 31737
rect 4094 31463 4122 31497
rect 70 31284 136 31318
rect 70 31092 136 31126
rect 4094 30913 4122 30947
rect 4094 30673 4122 30707
rect 70 30494 136 30528
rect 70 30302 136 30336
rect 4094 30123 4122 30157
rect 4094 29883 4122 29917
rect 70 29704 136 29738
rect 70 29512 136 29546
rect 4094 29333 4122 29367
rect 4094 29093 4122 29127
rect 70 28914 136 28948
rect 70 28722 136 28756
rect 4094 28543 4122 28577
rect 4094 28303 4122 28337
rect 70 28124 136 28158
rect 70 27932 136 27966
rect 4094 27753 4122 27787
rect 4094 27513 4122 27547
rect 70 27334 136 27368
rect 70 27142 136 27176
rect 4094 26963 4122 26997
rect 4094 26723 4122 26757
rect 70 26544 136 26578
rect 70 26352 136 26386
rect 4094 26173 4122 26207
rect 4094 25933 4122 25967
rect 70 25754 136 25788
rect 70 25562 136 25596
rect 4094 25383 4122 25417
rect 4094 25143 4122 25177
rect 70 24964 136 24998
rect 70 24772 136 24806
rect 4094 24593 4122 24627
rect 4094 24353 4122 24387
rect 70 24174 136 24208
rect 70 23982 136 24016
rect 4094 23803 4122 23837
rect 4094 23563 4122 23597
rect 70 23384 136 23418
rect 70 23192 136 23226
rect 4094 23013 4122 23047
rect 4094 22773 4122 22807
rect 70 22594 136 22628
rect 70 22402 136 22436
rect 4094 22223 4122 22257
rect 4094 21983 4122 22017
rect 70 21804 136 21838
rect 70 21612 136 21646
rect 4094 21433 4122 21467
rect 4094 21193 4122 21227
rect 70 21014 136 21048
rect 70 20822 136 20856
rect 4094 20643 4122 20677
rect 4094 20403 4122 20437
rect 70 20224 136 20258
rect 70 20032 136 20066
rect 4094 19853 4122 19887
rect 4094 19613 4122 19647
rect 70 19434 136 19468
rect 70 19242 136 19276
rect 4094 19063 4122 19097
rect 4094 18823 4122 18857
rect 70 18644 136 18678
rect 70 18452 136 18486
rect 4094 18273 4122 18307
rect 4094 18033 4122 18067
rect 70 17854 136 17888
rect 70 17662 136 17696
rect 4094 17483 4122 17517
rect 4094 17243 4122 17277
rect 70 17064 136 17098
rect 70 16872 136 16906
rect 4094 16693 4122 16727
rect 4094 16453 4122 16487
rect 70 16274 136 16308
rect 70 16082 136 16116
rect 4094 15903 4122 15937
rect 4094 15663 4122 15697
rect 70 15484 136 15518
rect 70 15292 136 15326
rect 4094 15113 4122 15147
rect 4094 14873 4122 14907
rect 70 14694 136 14728
rect 70 14502 136 14536
rect 4094 14323 4122 14357
rect 4094 14083 4122 14117
rect 70 13904 136 13938
rect 70 13712 136 13746
rect 4094 13533 4122 13567
rect 4094 13293 4122 13327
rect 70 13114 136 13148
rect 70 12922 136 12956
rect 4094 12743 4122 12777
rect 4094 12503 4122 12537
rect 70 12324 136 12358
rect 70 12132 136 12166
rect 4094 11953 4122 11987
rect 4094 11713 4122 11747
rect 70 11534 136 11568
rect 70 11342 136 11376
rect 4094 11163 4122 11197
rect 4094 10923 4122 10957
rect 70 10744 136 10778
rect 70 10552 136 10586
rect 4094 10373 4122 10407
rect 4094 10133 4122 10167
rect 70 9954 136 9988
rect 70 9762 136 9796
rect 4094 9583 4122 9617
rect 4094 9343 4122 9377
rect 70 9164 136 9198
rect 70 8972 136 9006
rect 4094 8793 4122 8827
rect 4094 8553 4122 8587
rect 70 8374 136 8408
rect 70 8182 136 8216
rect 4094 8003 4122 8037
rect 4094 7763 4122 7797
rect 70 7584 136 7618
rect 70 7392 136 7426
rect 4094 7213 4122 7247
rect 4094 6973 4122 7007
rect 70 6794 136 6828
rect 70 6602 136 6636
rect 4094 6423 4122 6457
rect 4094 6183 4122 6217
rect 70 6004 136 6038
rect 70 5812 136 5846
rect 4094 5633 4122 5667
rect 4094 5393 4122 5427
rect 70 5214 136 5248
rect 70 5022 136 5056
rect 4094 4843 4122 4877
rect 4094 4603 4122 4637
rect 70 4424 136 4458
rect 70 4232 136 4266
rect 4094 4053 4122 4087
rect 4094 3813 4122 3847
rect 70 3634 136 3668
rect 70 3442 136 3476
rect 4094 3263 4122 3297
rect 4094 3023 4122 3057
rect 70 2844 136 2878
rect 70 2652 136 2686
rect 4094 2473 4122 2507
rect 4094 2233 4122 2267
rect 70 2054 136 2088
rect 70 1862 136 1896
rect 4094 1683 4122 1717
rect 4094 1443 4122 1477
rect 70 1264 136 1298
rect 70 1072 136 1106
rect 4094 893 4122 927
rect 4094 653 4122 687
rect 70 474 136 508
rect 70 282 136 316
rect 4094 103 4122 137
<< metal1 >>
rect 71 50343 135 50395
rect 71 49935 135 49987
rect 71 49553 135 49605
rect 71 49145 135 49197
rect 71 48763 135 48815
rect 71 48355 135 48407
rect 71 47973 135 48025
rect 71 47565 135 47617
rect 71 47183 135 47235
rect 71 46775 135 46827
rect 71 46393 135 46445
rect 71 45985 135 46037
rect 71 45603 135 45655
rect 71 45195 135 45247
rect 71 44813 135 44865
rect 71 44405 135 44457
rect 71 44023 135 44075
rect 71 43615 135 43667
rect 71 43233 135 43285
rect 71 42825 135 42877
rect 71 42443 135 42495
rect 71 42035 135 42087
rect 71 41653 135 41705
rect 71 41245 135 41297
rect 71 40863 135 40915
rect 71 40455 135 40507
rect 71 40073 135 40125
rect 71 39665 135 39717
rect 71 39283 135 39335
rect 71 38875 135 38927
rect 71 38493 135 38545
rect 71 38085 135 38137
rect 71 37703 135 37755
rect 71 37295 135 37347
rect 71 36913 135 36965
rect 71 36505 135 36557
rect 71 36123 135 36175
rect 71 35715 135 35767
rect 71 35333 135 35385
rect 71 34925 135 34977
rect 71 34543 135 34595
rect 71 34135 135 34187
rect 71 33753 135 33805
rect 71 33345 135 33397
rect 71 32963 135 33015
rect 71 32555 135 32607
rect 71 32173 135 32225
rect 71 31765 135 31817
rect 71 31383 135 31435
rect 71 30975 135 31027
rect 71 30593 135 30645
rect 71 30185 135 30237
rect 71 29803 135 29855
rect 71 29395 135 29447
rect 71 29013 135 29065
rect 71 28605 135 28657
rect 71 28223 135 28275
rect 71 27815 135 27867
rect 71 27433 135 27485
rect 71 27025 135 27077
rect 71 26643 135 26695
rect 71 26235 135 26287
rect 71 25853 135 25905
rect 71 25445 135 25497
rect 71 25063 135 25115
rect 71 24655 135 24707
rect 71 24273 135 24325
rect 71 23865 135 23917
rect 71 23483 135 23535
rect 71 23075 135 23127
rect 71 22693 135 22745
rect 71 22285 135 22337
rect 71 21903 135 21955
rect 71 21495 135 21547
rect 71 21113 135 21165
rect 71 20705 135 20757
rect 71 20323 135 20375
rect 71 19915 135 19967
rect 71 19533 135 19585
rect 71 19125 135 19177
rect 71 18743 135 18795
rect 71 18335 135 18387
rect 71 17953 135 18005
rect 71 17545 135 17597
rect 71 17163 135 17215
rect 71 16755 135 16807
rect 71 16373 135 16425
rect 71 15965 135 16017
rect 71 15583 135 15635
rect 71 15175 135 15227
rect 71 14793 135 14845
rect 71 14385 135 14437
rect 71 14003 135 14055
rect 71 13595 135 13647
rect 71 13213 135 13265
rect 71 12805 135 12857
rect 71 12423 135 12475
rect 71 12015 135 12067
rect 71 11633 135 11685
rect 71 11225 135 11277
rect 71 10843 135 10895
rect 71 10435 135 10487
rect 71 10053 135 10105
rect 71 9645 135 9697
rect 71 9263 135 9315
rect 71 8855 135 8907
rect 71 8473 135 8525
rect 71 8065 135 8117
rect 71 7683 135 7735
rect 71 7275 135 7327
rect 71 6893 135 6945
rect 71 6485 135 6537
rect 71 6103 135 6155
rect 71 5695 135 5747
rect 71 5313 135 5365
rect 71 4905 135 4957
rect 71 4523 135 4575
rect 71 4115 135 4167
rect 71 3733 135 3785
rect 71 3325 135 3377
rect 71 2943 135 2995
rect 71 2535 135 2587
rect 71 2153 135 2205
rect 71 1745 135 1797
rect 71 1363 135 1415
rect 71 955 135 1007
rect 71 573 135 625
rect 71 165 135 217
rect 256 -30 284 50560
rect 681 -32 709 50560
rect 1724 0 1752 50560
rect 3372 0 3400 50560
<< metal2 >>
rect 70 0 98 50560
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_31
timestamp 1626486988
transform 1 0 74 0 1 158
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_31
timestamp 1626486988
transform 1 0 71 0 1 159
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_1
timestamp 1626486988
transform 1 0 0 0 -1 790
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_2
timestamp 1626486988
transform 1 0 0 0 1 0
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_30
timestamp 1626486988
transform 1 0 74 0 1 566
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_30
timestamp 1626486988
transform 1 0 71 0 1 567
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_29
timestamp 1626486988
transform 1 0 74 0 1 948
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_29
timestamp 1626486988
transform 1 0 71 0 1 949
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_5
timestamp 1626486988
transform 1 0 0 0 1 790
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_28
timestamp 1626486988
transform 1 0 74 0 1 1356
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_28
timestamp 1626486988
transform 1 0 71 0 1 1357
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_3
timestamp 1626486988
transform 1 0 0 0 1 1580
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_4
timestamp 1626486988
transform 1 0 0 0 -1 1580
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_27
timestamp 1626486988
transform 1 0 74 0 1 1738
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_27
timestamp 1626486988
transform 1 0 71 0 1 1739
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_0
timestamp 1626486988
transform 1 0 0 0 -1 2370
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_26
timestamp 1626486988
transform 1 0 74 0 1 2146
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_26
timestamp 1626486988
transform 1 0 71 0 1 2147
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_25
timestamp 1626486988
transform 1 0 74 0 1 2528
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_25
timestamp 1626486988
transform 1 0 71 0 1 2529
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_29
timestamp 1626486988
transform 1 0 0 0 -1 3160
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_30
timestamp 1626486988
transform 1 0 0 0 1 2370
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_24
timestamp 1626486988
transform 1 0 74 0 1 2936
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_24
timestamp 1626486988
transform 1 0 71 0 1 2937
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_28
timestamp 1626486988
transform 1 0 0 0 1 3160
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_23
timestamp 1626486988
transform 1 0 74 0 1 3318
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_23
timestamp 1626486988
transform 1 0 71 0 1 3319
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_22
timestamp 1626486988
transform 1 0 74 0 1 3726
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_22
timestamp 1626486988
transform 1 0 71 0 1 3727
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_27
timestamp 1626486988
transform 1 0 0 0 -1 3950
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_21
timestamp 1626486988
transform 1 0 74 0 1 4108
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_21
timestamp 1626486988
transform 1 0 71 0 1 4109
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_25
timestamp 1626486988
transform 1 0 0 0 -1 4740
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_26
timestamp 1626486988
transform 1 0 0 0 1 3950
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_20
timestamp 1626486988
transform 1 0 74 0 1 4516
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_20
timestamp 1626486988
transform 1 0 71 0 1 4517
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_24
timestamp 1626486988
transform 1 0 0 0 1 4740
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_19
timestamp 1626486988
transform 1 0 74 0 1 4898
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_19
timestamp 1626486988
transform 1 0 71 0 1 4899
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_18
timestamp 1626486988
transform 1 0 74 0 1 5306
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_18
timestamp 1626486988
transform 1 0 71 0 1 5307
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_23
timestamp 1626486988
transform 1 0 0 0 -1 5530
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_17
timestamp 1626486988
transform 1 0 74 0 1 5688
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_17
timestamp 1626486988
transform 1 0 71 0 1 5689
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_21
timestamp 1626486988
transform 1 0 0 0 -1 6320
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_22
timestamp 1626486988
transform 1 0 0 0 1 5530
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_16
timestamp 1626486988
transform 1 0 74 0 1 6096
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_16
timestamp 1626486988
transform 1 0 71 0 1 6097
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_15
timestamp 1626486988
transform 1 0 74 0 1 6478
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_15
timestamp 1626486988
transform 1 0 71 0 1 6479
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_20
timestamp 1626486988
transform 1 0 0 0 1 6320
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_14
timestamp 1626486988
transform 1 0 74 0 1 6886
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_14
timestamp 1626486988
transform 1 0 71 0 1 6887
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_18
timestamp 1626486988
transform 1 0 0 0 1 7110
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_19
timestamp 1626486988
transform 1 0 0 0 -1 7110
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_13
timestamp 1626486988
transform 1 0 74 0 1 7268
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_13
timestamp 1626486988
transform 1 0 71 0 1 7269
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_17
timestamp 1626486988
transform 1 0 0 0 -1 7900
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_12
timestamp 1626486988
transform 1 0 74 0 1 7676
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_12
timestamp 1626486988
transform 1 0 71 0 1 7677
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_11
timestamp 1626486988
transform 1 0 74 0 1 8058
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_11
timestamp 1626486988
transform 1 0 71 0 1 8059
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_16
timestamp 1626486988
transform 1 0 0 0 1 7900
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_10
timestamp 1626486988
transform 1 0 74 0 1 8466
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_10
timestamp 1626486988
transform 1 0 71 0 1 8467
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_14
timestamp 1626486988
transform 1 0 0 0 1 8690
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_15
timestamp 1626486988
transform 1 0 0 0 -1 8690
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_9
timestamp 1626486988
transform 1 0 74 0 1 8848
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_9
timestamp 1626486988
transform 1 0 71 0 1 8849
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_13
timestamp 1626486988
transform 1 0 0 0 -1 9480
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_8
timestamp 1626486988
transform 1 0 74 0 1 9256
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_8
timestamp 1626486988
transform 1 0 71 0 1 9257
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_7
timestamp 1626486988
transform 1 0 74 0 1 9638
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_7
timestamp 1626486988
transform 1 0 71 0 1 9639
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_11
timestamp 1626486988
transform 1 0 0 0 -1 10270
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_12
timestamp 1626486988
transform 1 0 0 0 1 9480
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_6
timestamp 1626486988
transform 1 0 74 0 1 10046
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_6
timestamp 1626486988
transform 1 0 71 0 1 10047
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_10
timestamp 1626486988
transform 1 0 0 0 1 10270
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_5
timestamp 1626486988
transform 1 0 74 0 1 10428
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_5
timestamp 1626486988
transform 1 0 71 0 1 10429
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_4
timestamp 1626486988
transform 1 0 74 0 1 10836
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_4
timestamp 1626486988
transform 1 0 71 0 1 10837
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_9
timestamp 1626486988
transform 1 0 0 0 -1 11060
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_3
timestamp 1626486988
transform 1 0 74 0 1 11218
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_3
timestamp 1626486988
transform 1 0 71 0 1 11219
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_7
timestamp 1626486988
transform 1 0 0 0 -1 11850
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_8
timestamp 1626486988
transform 1 0 0 0 1 11060
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_2
timestamp 1626486988
transform 1 0 74 0 1 11626
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1626486988
transform 1 0 71 0 1 11627
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_6
timestamp 1626486988
transform 1 0 0 0 1 11850
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1
timestamp 1626486988
transform 1 0 74 0 1 12008
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1626486988
transform 1 0 71 0 1 12009
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_0
timestamp 1626486988
transform 1 0 74 0 1 12416
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1626486988
transform 1 0 71 0 1 12417
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_62
timestamp 1626486988
transform 1 0 0 0 -1 12640
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_32
timestamp 1626486988
transform 1 0 71 0 1 12799
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_32
timestamp 1626486988
transform 1 0 74 0 1 12798
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_60
timestamp 1626486988
transform 1 0 0 0 -1 13430
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_61
timestamp 1626486988
transform 1 0 0 0 1 12640
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_63
timestamp 1626486988
transform 1 0 71 0 1 13207
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_63
timestamp 1626486988
transform 1 0 74 0 1 13588
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_62
timestamp 1626486988
transform 1 0 71 0 1 13589
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_33
timestamp 1626486988
transform 1 0 74 0 1 13206
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_59
timestamp 1626486988
transform 1 0 0 0 1 13430
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_62
timestamp 1626486988
transform 1 0 74 0 1 13996
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_61
timestamp 1626486988
transform 1 0 71 0 1 13997
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_57
timestamp 1626486988
transform 1 0 0 0 1 14220
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_58
timestamp 1626486988
transform 1 0 0 0 -1 14220
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_61
timestamp 1626486988
transform 1 0 74 0 1 14378
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_60
timestamp 1626486988
transform 1 0 71 0 1 14379
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_56
timestamp 1626486988
transform 1 0 0 0 -1 15010
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_60
timestamp 1626486988
transform 1 0 74 0 1 14786
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_59
timestamp 1626486988
transform 1 0 71 0 1 14787
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_59
timestamp 1626486988
transform 1 0 74 0 1 15168
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_58
timestamp 1626486988
transform 1 0 71 0 1 15169
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_55
timestamp 1626486988
transform 1 0 0 0 1 15010
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_58
timestamp 1626486988
transform 1 0 74 0 1 15576
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_57
timestamp 1626486988
transform 1 0 71 0 1 15577
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_53
timestamp 1626486988
transform 1 0 0 0 1 15800
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_54
timestamp 1626486988
transform 1 0 0 0 -1 15800
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_57
timestamp 1626486988
transform 1 0 74 0 1 15958
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_56
timestamp 1626486988
transform 1 0 71 0 1 15959
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_52
timestamp 1626486988
transform 1 0 0 0 -1 16590
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_56
timestamp 1626486988
transform 1 0 74 0 1 16366
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_55
timestamp 1626486988
transform 1 0 71 0 1 16367
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_55
timestamp 1626486988
transform 1 0 74 0 1 16748
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_54
timestamp 1626486988
transform 1 0 71 0 1 16749
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_50
timestamp 1626486988
transform 1 0 0 0 -1 17380
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_51
timestamp 1626486988
transform 1 0 0 0 1 16590
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_54
timestamp 1626486988
transform 1 0 74 0 1 17156
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_53
timestamp 1626486988
transform 1 0 71 0 1 17157
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_49
timestamp 1626486988
transform 1 0 0 0 1 17380
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_53
timestamp 1626486988
transform 1 0 74 0 1 17538
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_52
timestamp 1626486988
transform 1 0 71 0 1 17539
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_52
timestamp 1626486988
transform 1 0 74 0 1 17946
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_51
timestamp 1626486988
transform 1 0 71 0 1 17947
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_48
timestamp 1626486988
transform 1 0 0 0 -1 18170
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_51
timestamp 1626486988
transform 1 0 74 0 1 18328
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_50
timestamp 1626486988
transform 1 0 71 0 1 18329
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_46
timestamp 1626486988
transform 1 0 0 0 -1 18960
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_47
timestamp 1626486988
transform 1 0 0 0 1 18170
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_50
timestamp 1626486988
transform 1 0 74 0 1 18736
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_49
timestamp 1626486988
transform 1 0 71 0 1 18737
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_45
timestamp 1626486988
transform 1 0 0 0 1 18960
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_49
timestamp 1626486988
transform 1 0 74 0 1 19118
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_48
timestamp 1626486988
transform 1 0 71 0 1 19119
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_48
timestamp 1626486988
transform 1 0 74 0 1 19526
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_47
timestamp 1626486988
transform 1 0 71 0 1 19527
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_44
timestamp 1626486988
transform 1 0 0 0 -1 19750
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_47
timestamp 1626486988
transform 1 0 74 0 1 19908
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_46
timestamp 1626486988
transform 1 0 71 0 1 19909
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_42
timestamp 1626486988
transform 1 0 0 0 -1 20540
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_43
timestamp 1626486988
transform 1 0 0 0 1 19750
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_46
timestamp 1626486988
transform 1 0 74 0 1 20316
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_45
timestamp 1626486988
transform 1 0 71 0 1 20317
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_45
timestamp 1626486988
transform 1 0 74 0 1 20698
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_44
timestamp 1626486988
transform 1 0 71 0 1 20699
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_41
timestamp 1626486988
transform 1 0 0 0 1 20540
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_44
timestamp 1626486988
transform 1 0 74 0 1 21106
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_43
timestamp 1626486988
transform 1 0 71 0 1 21107
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_39
timestamp 1626486988
transform 1 0 0 0 1 21330
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_40
timestamp 1626486988
transform 1 0 0 0 -1 21330
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_43
timestamp 1626486988
transform 1 0 74 0 1 21488
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_42
timestamp 1626486988
transform 1 0 71 0 1 21489
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_38
timestamp 1626486988
transform 1 0 0 0 -1 22120
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_42
timestamp 1626486988
transform 1 0 74 0 1 21896
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_41
timestamp 1626486988
transform 1 0 71 0 1 21897
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_41
timestamp 1626486988
transform 1 0 74 0 1 22278
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_40
timestamp 1626486988
transform 1 0 71 0 1 22279
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_37
timestamp 1626486988
transform 1 0 0 0 1 22120
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_40
timestamp 1626486988
transform 1 0 74 0 1 22686
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_39
timestamp 1626486988
transform 1 0 71 0 1 22687
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_35
timestamp 1626486988
transform 1 0 0 0 1 22910
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_36
timestamp 1626486988
transform 1 0 0 0 -1 22910
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_39
timestamp 1626486988
transform 1 0 74 0 1 23068
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_38
timestamp 1626486988
transform 1 0 71 0 1 23069
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_34
timestamp 1626486988
transform 1 0 0 0 -1 23700
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_38
timestamp 1626486988
transform 1 0 74 0 1 23476
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_37
timestamp 1626486988
transform 1 0 71 0 1 23477
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_37
timestamp 1626486988
transform 1 0 74 0 1 23858
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_36
timestamp 1626486988
transform 1 0 71 0 1 23859
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_32
timestamp 1626486988
transform 1 0 0 0 -1 24490
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_33
timestamp 1626486988
transform 1 0 0 0 1 23700
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_36
timestamp 1626486988
transform 1 0 74 0 1 24266
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_35
timestamp 1626486988
transform 1 0 71 0 1 24267
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_31
timestamp 1626486988
transform 1 0 0 0 1 24490
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_35
timestamp 1626486988
transform 1 0 74 0 1 24648
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_34
timestamp 1626486988
transform 1 0 71 0 1 24649
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_34
timestamp 1626486988
transform 1 0 74 0 1 25056
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_33
timestamp 1626486988
transform 1 0 71 0 1 25057
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_127
timestamp 1626486988
transform 1 0 0 0 -1 25280
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_80
timestamp 1626486988
transform 1 0 74 0 1 25438
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_80
timestamp 1626486988
transform 1 0 71 0 1 25439
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_65
timestamp 1626486988
transform 1 0 0 0 -1 26070
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_126
timestamp 1626486988
transform 1 0 0 0 1 25280
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_79
timestamp 1626486988
transform 1 0 74 0 1 25846
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_79
timestamp 1626486988
transform 1 0 71 0 1 25847
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_64
timestamp 1626486988
transform 1 0 0 0 1 26070
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_78
timestamp 1626486988
transform 1 0 74 0 1 26228
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_78
timestamp 1626486988
transform 1 0 71 0 1 26229
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_77
timestamp 1626486988
transform 1 0 74 0 1 26636
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_77
timestamp 1626486988
transform 1 0 71 0 1 26637
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_63
timestamp 1626486988
transform 1 0 0 0 -1 26860
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_76
timestamp 1626486988
transform 1 0 74 0 1 27018
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_76
timestamp 1626486988
transform 1 0 71 0 1 27019
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_91
timestamp 1626486988
transform 1 0 0 0 -1 27650
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_92
timestamp 1626486988
transform 1 0 0 0 1 26860
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_75
timestamp 1626486988
transform 1 0 74 0 1 27426
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_75
timestamp 1626486988
transform 1 0 71 0 1 27427
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_74
timestamp 1626486988
transform 1 0 74 0 1 27808
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_74
timestamp 1626486988
transform 1 0 71 0 1 27809
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_90
timestamp 1626486988
transform 1 0 0 0 1 27650
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_73
timestamp 1626486988
transform 1 0 74 0 1 28216
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_73
timestamp 1626486988
transform 1 0 71 0 1 28217
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_88
timestamp 1626486988
transform 1 0 0 0 1 28440
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_89
timestamp 1626486988
transform 1 0 0 0 -1 28440
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_72
timestamp 1626486988
transform 1 0 74 0 1 28598
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_72
timestamp 1626486988
transform 1 0 71 0 1 28599
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_87
timestamp 1626486988
transform 1 0 0 0 -1 29230
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_71
timestamp 1626486988
transform 1 0 74 0 1 29006
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_71
timestamp 1626486988
transform 1 0 71 0 1 29007
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_70
timestamp 1626486988
transform 1 0 74 0 1 29388
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_70
timestamp 1626486988
transform 1 0 71 0 1 29389
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_86
timestamp 1626486988
transform 1 0 0 0 1 29230
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_69
timestamp 1626486988
transform 1 0 74 0 1 29796
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_69
timestamp 1626486988
transform 1 0 71 0 1 29797
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_84
timestamp 1626486988
transform 1 0 0 0 1 30020
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_85
timestamp 1626486988
transform 1 0 0 0 -1 30020
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_68
timestamp 1626486988
transform 1 0 74 0 1 30178
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_68
timestamp 1626486988
transform 1 0 71 0 1 30179
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_83
timestamp 1626486988
transform 1 0 0 0 -1 30810
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_67
timestamp 1626486988
transform 1 0 74 0 1 30586
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_67
timestamp 1626486988
transform 1 0 71 0 1 30587
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_66
timestamp 1626486988
transform 1 0 74 0 1 30968
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_66
timestamp 1626486988
transform 1 0 71 0 1 30969
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_81
timestamp 1626486988
transform 1 0 0 0 -1 31600
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_82
timestamp 1626486988
transform 1 0 0 0 1 30810
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_65
timestamp 1626486988
transform 1 0 74 0 1 31376
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_65
timestamp 1626486988
transform 1 0 71 0 1 31377
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_80
timestamp 1626486988
transform 1 0 0 0 1 31600
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_95
timestamp 1626486988
transform 1 0 74 0 1 32166
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_95
timestamp 1626486988
transform 1 0 71 0 1 32167
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_64
timestamp 1626486988
transform 1 0 74 0 1 31758
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_64
timestamp 1626486988
transform 1 0 71 0 1 31759
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_79
timestamp 1626486988
transform 1 0 0 0 -1 32390
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_94
timestamp 1626486988
transform 1 0 74 0 1 32548
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_94
timestamp 1626486988
transform 1 0 71 0 1 32549
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_77
timestamp 1626486988
transform 1 0 0 0 -1 33180
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_78
timestamp 1626486988
transform 1 0 0 0 1 32390
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_93
timestamp 1626486988
transform 1 0 74 0 1 32956
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_93
timestamp 1626486988
transform 1 0 71 0 1 32957
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_76
timestamp 1626486988
transform 1 0 0 0 1 33180
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_92
timestamp 1626486988
transform 1 0 74 0 1 33338
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_92
timestamp 1626486988
transform 1 0 71 0 1 33339
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_91
timestamp 1626486988
transform 1 0 74 0 1 33746
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_91
timestamp 1626486988
transform 1 0 71 0 1 33747
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_75
timestamp 1626486988
transform 1 0 0 0 -1 33970
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_90
timestamp 1626486988
transform 1 0 74 0 1 34128
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_90
timestamp 1626486988
transform 1 0 71 0 1 34129
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_73
timestamp 1626486988
transform 1 0 0 0 -1 34760
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_74
timestamp 1626486988
transform 1 0 0 0 1 33970
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_89
timestamp 1626486988
transform 1 0 74 0 1 34536
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_89
timestamp 1626486988
transform 1 0 71 0 1 34537
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_88
timestamp 1626486988
transform 1 0 74 0 1 34918
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_88
timestamp 1626486988
transform 1 0 71 0 1 34919
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_72
timestamp 1626486988
transform 1 0 0 0 1 34760
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_87
timestamp 1626486988
transform 1 0 74 0 1 35326
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_87
timestamp 1626486988
transform 1 0 71 0 1 35327
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_70
timestamp 1626486988
transform 1 0 0 0 1 35550
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_71
timestamp 1626486988
transform 1 0 0 0 -1 35550
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_86
timestamp 1626486988
transform 1 0 74 0 1 35708
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_86
timestamp 1626486988
transform 1 0 71 0 1 35709
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_69
timestamp 1626486988
transform 1 0 0 0 -1 36340
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_85
timestamp 1626486988
transform 1 0 74 0 1 36116
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_85
timestamp 1626486988
transform 1 0 71 0 1 36117
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_84
timestamp 1626486988
transform 1 0 74 0 1 36498
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_84
timestamp 1626486988
transform 1 0 71 0 1 36499
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_68
timestamp 1626486988
transform 1 0 0 0 1 36340
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_83
timestamp 1626486988
transform 1 0 74 0 1 36906
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_83
timestamp 1626486988
transform 1 0 71 0 1 36907
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_66
timestamp 1626486988
transform 1 0 0 0 1 37130
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_67
timestamp 1626486988
transform 1 0 0 0 -1 37130
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_82
timestamp 1626486988
transform 1 0 74 0 1 37288
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_82
timestamp 1626486988
transform 1 0 71 0 1 37289
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_125
timestamp 1626486988
transform 1 0 0 0 -1 37920
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_127
timestamp 1626486988
transform 1 0 74 0 1 38078
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_127
timestamp 1626486988
transform 1 0 71 0 1 38079
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_81
timestamp 1626486988
transform 1 0 74 0 1 37696
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_81
timestamp 1626486988
transform 1 0 71 0 1 37697
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_123
timestamp 1626486988
transform 1 0 0 0 -1 38710
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_124
timestamp 1626486988
transform 1 0 0 0 1 37920
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_126
timestamp 1626486988
transform 1 0 74 0 1 38486
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_126
timestamp 1626486988
transform 1 0 71 0 1 38487
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_122
timestamp 1626486988
transform 1 0 0 0 1 38710
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_125
timestamp 1626486988
transform 1 0 74 0 1 38868
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_125
timestamp 1626486988
transform 1 0 71 0 1 38869
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_124
timestamp 1626486988
transform 1 0 74 0 1 39276
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_124
timestamp 1626486988
transform 1 0 71 0 1 39277
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_121
timestamp 1626486988
transform 1 0 0 0 -1 39500
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_123
timestamp 1626486988
transform 1 0 74 0 1 39658
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_123
timestamp 1626486988
transform 1 0 71 0 1 39659
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_119
timestamp 1626486988
transform 1 0 0 0 -1 40290
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_120
timestamp 1626486988
transform 1 0 0 0 1 39500
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_122
timestamp 1626486988
transform 1 0 74 0 1 40066
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_122
timestamp 1626486988
transform 1 0 71 0 1 40067
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_118
timestamp 1626486988
transform 1 0 0 0 1 40290
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_121
timestamp 1626486988
transform 1 0 74 0 1 40448
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_121
timestamp 1626486988
transform 1 0 71 0 1 40449
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_120
timestamp 1626486988
transform 1 0 74 0 1 40856
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_120
timestamp 1626486988
transform 1 0 71 0 1 40857
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_117
timestamp 1626486988
transform 1 0 0 0 -1 41080
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_119
timestamp 1626486988
transform 1 0 74 0 1 41238
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_119
timestamp 1626486988
transform 1 0 71 0 1 41239
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_115
timestamp 1626486988
transform 1 0 0 0 -1 41870
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_116
timestamp 1626486988
transform 1 0 0 0 1 41080
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_118
timestamp 1626486988
transform 1 0 74 0 1 41646
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_118
timestamp 1626486988
transform 1 0 71 0 1 41647
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_117
timestamp 1626486988
transform 1 0 74 0 1 42028
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_117
timestamp 1626486988
transform 1 0 71 0 1 42029
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_114
timestamp 1626486988
transform 1 0 0 0 1 41870
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_116
timestamp 1626486988
transform 1 0 74 0 1 42436
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_116
timestamp 1626486988
transform 1 0 71 0 1 42437
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_112
timestamp 1626486988
transform 1 0 0 0 1 42660
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_113
timestamp 1626486988
transform 1 0 0 0 -1 42660
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_115
timestamp 1626486988
transform 1 0 74 0 1 42818
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_115
timestamp 1626486988
transform 1 0 71 0 1 42819
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_111
timestamp 1626486988
transform 1 0 0 0 -1 43450
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_114
timestamp 1626486988
transform 1 0 74 0 1 43226
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_114
timestamp 1626486988
transform 1 0 71 0 1 43227
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_113
timestamp 1626486988
transform 1 0 74 0 1 43608
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_113
timestamp 1626486988
transform 1 0 71 0 1 43609
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_110
timestamp 1626486988
transform 1 0 0 0 1 43450
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_112
timestamp 1626486988
transform 1 0 74 0 1 44016
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_112
timestamp 1626486988
transform 1 0 71 0 1 44017
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_108
timestamp 1626486988
transform 1 0 0 0 1 44240
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_109
timestamp 1626486988
transform 1 0 0 0 -1 44240
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_111
timestamp 1626486988
transform 1 0 74 0 1 44398
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_111
timestamp 1626486988
transform 1 0 71 0 1 44399
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_107
timestamp 1626486988
transform 1 0 0 0 -1 45030
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_110
timestamp 1626486988
transform 1 0 74 0 1 44806
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_110
timestamp 1626486988
transform 1 0 71 0 1 44807
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_109
timestamp 1626486988
transform 1 0 74 0 1 45188
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_109
timestamp 1626486988
transform 1 0 71 0 1 45189
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_105
timestamp 1626486988
transform 1 0 0 0 -1 45820
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_106
timestamp 1626486988
transform 1 0 0 0 1 45030
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_108
timestamp 1626486988
transform 1 0 74 0 1 45596
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_108
timestamp 1626486988
transform 1 0 71 0 1 45597
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_104
timestamp 1626486988
transform 1 0 0 0 1 45820
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_107
timestamp 1626486988
transform 1 0 74 0 1 45978
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_107
timestamp 1626486988
transform 1 0 71 0 1 45979
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_106
timestamp 1626486988
transform 1 0 74 0 1 46386
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_106
timestamp 1626486988
transform 1 0 71 0 1 46387
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_103
timestamp 1626486988
transform 1 0 0 0 -1 46610
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_105
timestamp 1626486988
transform 1 0 74 0 1 46768
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_105
timestamp 1626486988
transform 1 0 71 0 1 46769
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_101
timestamp 1626486988
transform 1 0 0 0 -1 47400
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_102
timestamp 1626486988
transform 1 0 0 0 1 46610
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_104
timestamp 1626486988
transform 1 0 74 0 1 47176
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_104
timestamp 1626486988
transform 1 0 71 0 1 47177
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_100
timestamp 1626486988
transform 1 0 0 0 1 47400
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_103
timestamp 1626486988
transform 1 0 74 0 1 47558
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_103
timestamp 1626486988
transform 1 0 71 0 1 47559
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_102
timestamp 1626486988
transform 1 0 74 0 1 47966
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_102
timestamp 1626486988
transform 1 0 71 0 1 47967
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_99
timestamp 1626486988
transform 1 0 0 0 -1 48190
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_101
timestamp 1626486988
transform 1 0 74 0 1 48348
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_101
timestamp 1626486988
transform 1 0 71 0 1 48349
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_97
timestamp 1626486988
transform 1 0 0 0 -1 48980
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_98
timestamp 1626486988
transform 1 0 0 0 1 48190
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_100
timestamp 1626486988
transform 1 0 74 0 1 48756
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_100
timestamp 1626486988
transform 1 0 71 0 1 48757
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_99
timestamp 1626486988
transform 1 0 74 0 1 49138
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_99
timestamp 1626486988
transform 1 0 71 0 1 49139
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_96
timestamp 1626486988
transform 1 0 0 0 1 48980
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_98
timestamp 1626486988
transform 1 0 74 0 1 49546
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_98
timestamp 1626486988
transform 1 0 71 0 1 49547
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_94
timestamp 1626486988
transform 1 0 0 0 1 49770
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_95
timestamp 1626486988
transform 1 0 0 0 -1 49770
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_97
timestamp 1626486988
transform 1 0 74 0 1 49928
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_97
timestamp 1626486988
transform 1 0 71 0 1 49929
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver  sky130_sram_2kbyte_1rw1r_32x512_8_wordline_driver_93
timestamp 1626486988
transform 1 0 0 0 -1 50560
box 70 -56 4140 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_96
timestamp 1626486988
transform 1 0 74 0 1 50336
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_96
timestamp 1626486988
transform 1 0 71 0 1 50337
box 0 0 64 64
<< labels >>
rlabel metal2 s 70 0 98 50560 4 en
rlabel metal1 s 681 -32 709 50560 4 vdd
rlabel metal1 s 3372 0 3400 50560 4 vdd
rlabel metal1 s 256 -30 284 50560 4 gnd
rlabel metal1 s 1724 0 1752 50560 4 gnd
rlabel locali s 4108 25400 4108 25400 4 wl_64
rlabel locali s 4108 25950 4108 25950 4 wl_65
rlabel locali s 4108 26190 4108 26190 4 wl_66
rlabel locali s 4108 26740 4108 26740 4 wl_67
rlabel locali s 4108 26980 4108 26980 4 wl_68
rlabel locali s 4108 27530 4108 27530 4 wl_69
rlabel locali s 4108 27770 4108 27770 4 wl_70
rlabel locali s 4108 28320 4108 28320 4 wl_71
rlabel locali s 4108 28560 4108 28560 4 wl_72
rlabel locali s 4108 29110 4108 29110 4 wl_73
rlabel locali s 4108 29350 4108 29350 4 wl_74
rlabel locali s 4108 29900 4108 29900 4 wl_75
rlabel locali s 4108 30140 4108 30140 4 wl_76
rlabel locali s 4108 30690 4108 30690 4 wl_77
rlabel locali s 4108 30930 4108 30930 4 wl_78
rlabel locali s 4108 31480 4108 31480 4 wl_79
rlabel locali s 4108 31720 4108 31720 4 wl_80
rlabel locali s 4108 32270 4108 32270 4 wl_81
rlabel locali s 4108 32510 4108 32510 4 wl_82
rlabel locali s 4108 33060 4108 33060 4 wl_83
rlabel locali s 4108 33300 4108 33300 4 wl_84
rlabel locali s 4108 33850 4108 33850 4 wl_85
rlabel locali s 4108 34090 4108 34090 4 wl_86
rlabel locali s 4108 34640 4108 34640 4 wl_87
rlabel locali s 4108 34880 4108 34880 4 wl_88
rlabel locali s 4108 35430 4108 35430 4 wl_89
rlabel locali s 4108 35670 4108 35670 4 wl_90
rlabel locali s 4108 36220 4108 36220 4 wl_91
rlabel locali s 4108 36460 4108 36460 4 wl_92
rlabel locali s 4108 37010 4108 37010 4 wl_93
rlabel locali s 4108 37250 4108 37250 4 wl_94
rlabel locali s 4108 37800 4108 37800 4 wl_95
rlabel locali s 4108 38040 4108 38040 4 wl_96
rlabel locali s 4108 38590 4108 38590 4 wl_97
rlabel locali s 4108 38830 4108 38830 4 wl_98
rlabel locali s 4108 39380 4108 39380 4 wl_99
rlabel locali s 4108 39620 4108 39620 4 wl_100
rlabel locali s 4108 40170 4108 40170 4 wl_101
rlabel locali s 4108 40410 4108 40410 4 wl_102
rlabel locali s 4108 40960 4108 40960 4 wl_103
rlabel locali s 4108 41200 4108 41200 4 wl_104
rlabel locali s 4108 41750 4108 41750 4 wl_105
rlabel locali s 4108 41990 4108 41990 4 wl_106
rlabel locali s 4108 42540 4108 42540 4 wl_107
rlabel locali s 4108 42780 4108 42780 4 wl_108
rlabel locali s 4108 43330 4108 43330 4 wl_109
rlabel locali s 4108 43570 4108 43570 4 wl_110
rlabel locali s 4108 44120 4108 44120 4 wl_111
rlabel locali s 4108 44360 4108 44360 4 wl_112
rlabel locali s 4108 44910 4108 44910 4 wl_113
rlabel locali s 4108 45150 4108 45150 4 wl_114
rlabel locali s 4108 45700 4108 45700 4 wl_115
rlabel locali s 4108 45940 4108 45940 4 wl_116
rlabel locali s 4108 46490 4108 46490 4 wl_117
rlabel locali s 4108 46730 4108 46730 4 wl_118
rlabel locali s 4108 47280 4108 47280 4 wl_119
rlabel locali s 4108 47520 4108 47520 4 wl_120
rlabel locali s 4108 48070 4108 48070 4 wl_121
rlabel locali s 4108 48310 4108 48310 4 wl_122
rlabel locali s 4108 48860 4108 48860 4 wl_123
rlabel locali s 4108 49100 4108 49100 4 wl_124
rlabel locali s 4108 49650 4108 49650 4 wl_125
rlabel locali s 4108 49890 4108 49890 4 wl_126
rlabel locali s 4108 50440 4108 50440 4 wl_127
rlabel locali s 103 38219 103 38219 4 in_96
rlabel locali s 103 31899 103 31899 4 in_80
rlabel locali s 103 38411 103 38411 4 in_97
rlabel locali s 103 28739 103 28739 4 in_72
rlabel locali s 103 39009 103 39009 4 in_98
rlabel locali s 103 32091 103 32091 4 in_81
rlabel locali s 103 39201 103 39201 4 in_99
rlabel locali s 103 27159 103 27159 4 in_68
rlabel locali s 103 39799 103 39799 4 in_100
rlabel locali s 103 32689 103 32689 4 in_82
rlabel locali s 103 39991 103 39991 4 in_101
rlabel locali s 103 28931 103 28931 4 in_73
rlabel locali s 103 40589 103 40589 4 in_102
rlabel locali s 103 32881 103 32881 4 in_83
rlabel locali s 103 40781 103 40781 4 in_103
rlabel locali s 103 26369 103 26369 4 in_66
rlabel locali s 103 41379 103 41379 4 in_104
rlabel locali s 103 33479 103 33479 4 in_84
rlabel locali s 103 41571 103 41571 4 in_105
rlabel locali s 103 29529 103 29529 4 in_74
rlabel locali s 103 42169 103 42169 4 in_106
rlabel locali s 103 33671 103 33671 4 in_85
rlabel locali s 103 42361 103 42361 4 in_107
rlabel locali s 103 27351 103 27351 4 in_69
rlabel locali s 103 42959 103 42959 4 in_108
rlabel locali s 103 34269 103 34269 4 in_86
rlabel locali s 103 43151 103 43151 4 in_109
rlabel locali s 103 29721 103 29721 4 in_75
rlabel locali s 103 43749 103 43749 4 in_110
rlabel locali s 103 34461 103 34461 4 in_87
rlabel locali s 103 43941 103 43941 4 in_111
rlabel locali s 103 25771 103 25771 4 in_65
rlabel locali s 103 44539 103 44539 4 in_112
rlabel locali s 103 35059 103 35059 4 in_88
rlabel locali s 103 44731 103 44731 4 in_113
rlabel locali s 103 30319 103 30319 4 in_76
rlabel locali s 103 45329 103 45329 4 in_114
rlabel locali s 103 35251 103 35251 4 in_89
rlabel locali s 103 45521 103 45521 4 in_115
rlabel locali s 103 27949 103 27949 4 in_70
rlabel locali s 103 46119 103 46119 4 in_116
rlabel locali s 103 35849 103 35849 4 in_90
rlabel locali s 103 46311 103 46311 4 in_117
rlabel locali s 103 30511 103 30511 4 in_77
rlabel locali s 103 46909 103 46909 4 in_118
rlabel locali s 103 36041 103 36041 4 in_91
rlabel locali s 103 47101 103 47101 4 in_119
rlabel locali s 103 26561 103 26561 4 in_67
rlabel locali s 103 47699 103 47699 4 in_120
rlabel locali s 103 36639 103 36639 4 in_92
rlabel locali s 103 47891 103 47891 4 in_121
rlabel locali s 103 31109 103 31109 4 in_78
rlabel locali s 103 48489 103 48489 4 in_122
rlabel locali s 103 36831 103 36831 4 in_93
rlabel locali s 103 48681 103 48681 4 in_123
rlabel locali s 103 28141 103 28141 4 in_71
rlabel locali s 103 49279 103 49279 4 in_124
rlabel locali s 103 37429 103 37429 4 in_94
rlabel locali s 103 49471 103 49471 4 in_125
rlabel locali s 103 31301 103 31301 4 in_79
rlabel locali s 103 50069 103 50069 4 in_126
rlabel locali s 103 37621 103 37621 4 in_95
rlabel locali s 103 50261 103 50261 4 in_127
rlabel locali s 103 25579 103 25579 4 in_64
rlabel locali s 103 299 103 299 4 in_0
rlabel locali s 103 491 103 491 4 in_1
rlabel locali s 103 1089 103 1089 4 in_2
rlabel locali s 103 1281 103 1281 4 in_3
rlabel locali s 103 1879 103 1879 4 in_4
rlabel locali s 103 2071 103 2071 4 in_5
rlabel locali s 103 2669 103 2669 4 in_6
rlabel locali s 103 2861 103 2861 4 in_7
rlabel locali s 103 3459 103 3459 4 in_8
rlabel locali s 103 3651 103 3651 4 in_9
rlabel locali s 103 4249 103 4249 4 in_10
rlabel locali s 103 4441 103 4441 4 in_11
rlabel locali s 103 5039 103 5039 4 in_12
rlabel locali s 103 5231 103 5231 4 in_13
rlabel locali s 103 5829 103 5829 4 in_14
rlabel locali s 103 6021 103 6021 4 in_15
rlabel locali s 103 6619 103 6619 4 in_16
rlabel locali s 103 6811 103 6811 4 in_17
rlabel locali s 103 7409 103 7409 4 in_18
rlabel locali s 103 7601 103 7601 4 in_19
rlabel locali s 103 8199 103 8199 4 in_20
rlabel locali s 103 8391 103 8391 4 in_21
rlabel locali s 103 8989 103 8989 4 in_22
rlabel locali s 103 9181 103 9181 4 in_23
rlabel locali s 103 9779 103 9779 4 in_24
rlabel locali s 103 9971 103 9971 4 in_25
rlabel locali s 103 10569 103 10569 4 in_26
rlabel locali s 103 10761 103 10761 4 in_27
rlabel locali s 103 11359 103 11359 4 in_28
rlabel locali s 103 11551 103 11551 4 in_29
rlabel locali s 103 12149 103 12149 4 in_30
rlabel locali s 103 12341 103 12341 4 in_31
rlabel locali s 103 12939 103 12939 4 in_32
rlabel locali s 103 13131 103 13131 4 in_33
rlabel locali s 103 13729 103 13729 4 in_34
rlabel locali s 103 13921 103 13921 4 in_35
rlabel locali s 103 14519 103 14519 4 in_36
rlabel locali s 103 14711 103 14711 4 in_37
rlabel locali s 103 15309 103 15309 4 in_38
rlabel locali s 103 15501 103 15501 4 in_39
rlabel locali s 103 16099 103 16099 4 in_40
rlabel locali s 103 16291 103 16291 4 in_41
rlabel locali s 103 16889 103 16889 4 in_42
rlabel locali s 103 17081 103 17081 4 in_43
rlabel locali s 103 17679 103 17679 4 in_44
rlabel locali s 103 17871 103 17871 4 in_45
rlabel locali s 103 18469 103 18469 4 in_46
rlabel locali s 103 18661 103 18661 4 in_47
rlabel locali s 103 19259 103 19259 4 in_48
rlabel locali s 103 19451 103 19451 4 in_49
rlabel locali s 103 20049 103 20049 4 in_50
rlabel locali s 103 20241 103 20241 4 in_51
rlabel locali s 103 20839 103 20839 4 in_52
rlabel locali s 103 21031 103 21031 4 in_53
rlabel locali s 103 21629 103 21629 4 in_54
rlabel locali s 103 21821 103 21821 4 in_55
rlabel locali s 103 22419 103 22419 4 in_56
rlabel locali s 103 22611 103 22611 4 in_57
rlabel locali s 103 23209 103 23209 4 in_58
rlabel locali s 103 23401 103 23401 4 in_59
rlabel locali s 103 23999 103 23999 4 in_60
rlabel locali s 103 24191 103 24191 4 in_61
rlabel locali s 103 24789 103 24789 4 in_62
rlabel locali s 103 24981 103 24981 4 in_63
rlabel locali s 4108 120 4108 120 4 wl_0
rlabel locali s 4108 12760 4108 12760 4 wl_32
rlabel locali s 4108 6440 4108 6440 4 wl_16
rlabel locali s 4108 13310 4108 13310 4 wl_33
rlabel locali s 4108 3280 4108 3280 4 wl_8
rlabel locali s 4108 13550 4108 13550 4 wl_34
rlabel locali s 4108 6990 4108 6990 4 wl_17
rlabel locali s 4108 14100 4108 14100 4 wl_35
rlabel locali s 4108 1700 4108 1700 4 wl_4
rlabel locali s 4108 14340 4108 14340 4 wl_36
rlabel locali s 4108 7230 4108 7230 4 wl_18
rlabel locali s 4108 14890 4108 14890 4 wl_37
rlabel locali s 4108 3830 4108 3830 4 wl_9
rlabel locali s 4108 15130 4108 15130 4 wl_38
rlabel locali s 4108 7780 4108 7780 4 wl_19
rlabel locali s 4108 15680 4108 15680 4 wl_39
rlabel locali s 4108 910 4108 910 4 wl_2
rlabel locali s 4108 15920 4108 15920 4 wl_40
rlabel locali s 4108 8020 4108 8020 4 wl_20
rlabel locali s 4108 16470 4108 16470 4 wl_41
rlabel locali s 4108 4070 4108 4070 4 wl_10
rlabel locali s 4108 16710 4108 16710 4 wl_42
rlabel locali s 4108 8570 4108 8570 4 wl_21
rlabel locali s 4108 17260 4108 17260 4 wl_43
rlabel locali s 4108 2250 4108 2250 4 wl_5
rlabel locali s 4108 17500 4108 17500 4 wl_44
rlabel locali s 4108 8810 4108 8810 4 wl_22
rlabel locali s 4108 18050 4108 18050 4 wl_45
rlabel locali s 4108 4620 4108 4620 4 wl_11
rlabel locali s 4108 18290 4108 18290 4 wl_46
rlabel locali s 4108 9360 4108 9360 4 wl_23
rlabel locali s 4108 18840 4108 18840 4 wl_47
rlabel locali s 4108 670 4108 670 4 wl_1
rlabel locali s 4108 19080 4108 19080 4 wl_48
rlabel locali s 4108 9600 4108 9600 4 wl_24
rlabel locali s 4108 19630 4108 19630 4 wl_49
rlabel locali s 4108 4860 4108 4860 4 wl_12
rlabel locali s 4108 19870 4108 19870 4 wl_50
rlabel locali s 4108 10150 4108 10150 4 wl_25
rlabel locali s 4108 20420 4108 20420 4 wl_51
rlabel locali s 4108 2490 4108 2490 4 wl_6
rlabel locali s 4108 20660 4108 20660 4 wl_52
rlabel locali s 4108 10390 4108 10390 4 wl_26
rlabel locali s 4108 21210 4108 21210 4 wl_53
rlabel locali s 4108 5410 4108 5410 4 wl_13
rlabel locali s 4108 21450 4108 21450 4 wl_54
rlabel locali s 4108 10940 4108 10940 4 wl_27
rlabel locali s 4108 22000 4108 22000 4 wl_55
rlabel locali s 4108 1460 4108 1460 4 wl_3
rlabel locali s 4108 22240 4108 22240 4 wl_56
rlabel locali s 4108 11180 4108 11180 4 wl_28
rlabel locali s 4108 22790 4108 22790 4 wl_57
rlabel locali s 4108 5650 4108 5650 4 wl_14
rlabel locali s 4108 23030 4108 23030 4 wl_58
rlabel locali s 4108 11730 4108 11730 4 wl_29
rlabel locali s 4108 23580 4108 23580 4 wl_59
rlabel locali s 4108 3040 4108 3040 4 wl_7
rlabel locali s 4108 23820 4108 23820 4 wl_60
rlabel locali s 4108 11970 4108 11970 4 wl_30
rlabel locali s 4108 24370 4108 24370 4 wl_61
rlabel locali s 4108 6200 4108 6200 4 wl_15
rlabel locali s 4108 24610 4108 24610 4 wl_62
rlabel locali s 4108 12520 4108 12520 4 wl_31
rlabel locali s 4108 25160 4108 25160 4 wl_63
<< properties >>
string FIXED_BBOX 0 0 4158 50560
<< end >>
