magic
tech sky130A
timestamp 1626486988
<< checkpaint >>
rect -854 -798 854 798
<< metal4 >>
rect -224 139 224 168
rect -224 -139 -139 139
rect 139 -139 224 139
rect -224 -168 224 -139
<< via4 >>
rect -139 -139 139 139
<< metal5 >>
rect -224 139 224 168
rect -224 -139 -139 139
rect 139 -139 224 139
rect -224 -168 224 -139
<< end >>
