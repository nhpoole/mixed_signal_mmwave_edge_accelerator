magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -14774 32200 37172 32258
rect -87761 -1968 37172 32200
rect -87761 -43940 12313 -1968
<< nwell >>
rect -11247 15506 -9306 16346
rect -7803 15507 -7200 15828
<< locali >>
rect -7288 15499 -7240 15506
rect -7288 15465 -7281 15499
rect -7247 15465 -7240 15499
rect -7288 15458 -7240 15465
rect -7184 15503 -7136 15510
rect -7184 15469 -7177 15503
rect -7143 15469 -7136 15503
rect -7184 15462 -7136 15469
<< viali >>
rect -7281 15465 -7247 15499
rect -7177 15469 -7143 15503
<< metal1 >>
rect -4458 30284 -4398 30294
rect -4458 30232 -4454 30284
rect -4402 30232 -4398 30284
rect -4458 16436 -4398 30232
rect -11018 16376 -9518 16436
rect -8284 16432 -7850 16436
rect -8284 16380 -7912 16432
rect -7860 16380 -7850 16432
rect -8284 16376 -7850 16380
rect -4464 16432 -4392 16436
rect -4464 16380 -4454 16432
rect -4402 16380 -4392 16432
rect -4464 16376 -4392 16380
rect -7540 15742 -7332 15838
rect -7490 15499 -7228 15512
rect -7490 15465 -7281 15499
rect -7247 15465 -7228 15499
rect -7490 15452 -7228 15465
rect -7196 15503 -7030 15516
rect -7196 15469 -7177 15503
rect -7143 15469 -7030 15503
rect -7196 15456 -7030 15469
rect -7528 15198 -7326 15294
rect -9694 14740 -9688 14760
rect -11068 14680 -9566 14740
rect -8452 14680 -1320 14740
rect 664 1564 1066 1624
<< via1 >>
rect -4454 30232 -4402 30284
rect -7912 16380 -7860 16432
rect -4454 16380 -4402 16432
<< metal2 >>
rect -4458 30288 -4398 30297
rect -4464 30286 -4392 30288
rect -4464 30230 -4456 30286
rect -4400 30230 -4392 30286
rect -4464 30228 -4392 30230
rect -4458 30219 -4398 30228
rect -7916 16436 -7856 16442
rect -4458 16436 -4398 16442
rect -7916 16432 -4398 16436
rect -7916 16380 -7912 16432
rect -7860 16380 -4454 16432
rect -4402 16380 -4398 16432
rect -7916 16376 -4398 16380
rect -7916 16370 -7856 16376
rect -4458 16370 -4398 16376
rect -13297 15560 -11530 15562
rect -13297 15504 -13286 15560
rect -13230 15504 -11530 15560
rect -13297 15502 -11530 15504
rect -9675 15560 -8926 15562
rect -9675 15504 -9664 15560
rect -9608 15504 -8926 15560
rect -9675 15502 -8926 15504
rect -12495 15411 -11732 15413
rect -12495 15355 -12484 15411
rect -12428 15355 -11732 15411
rect -12495 15353 -11732 15355
rect -9859 15411 -9164 15413
rect -9859 15355 -9848 15411
rect -9792 15355 -9164 15411
rect -9859 15353 -9164 15355
rect -10082 14806 -7716 14866
rect -13105 14576 -13015 14580
rect -9874 14576 -9774 14585
rect -13110 14554 -9766 14576
rect -13110 14498 -13088 14554
rect -13032 14498 -9852 14554
rect -9796 14498 -9766 14554
rect -13110 14476 -9766 14498
rect -13105 14472 -13015 14476
rect -9874 14467 -9774 14476
rect -13499 14354 -13409 14358
rect -9686 14354 -9586 14363
rect -13504 14332 -9586 14354
rect -13504 14276 -13482 14332
rect -13426 14276 -9664 14332
rect -9608 14276 -9586 14332
rect -13504 14254 -9586 14276
rect -13499 14250 -13409 14254
rect -9686 14245 -9586 14254
rect -11022 11009 -10932 11014
rect -11026 10997 -10928 11009
rect -6664 11001 -6578 11006
rect -11026 10941 -11005 10997
rect -10949 10941 -10928 10997
rect -11026 10929 -10928 10941
rect -6668 10991 -6574 11001
rect -6668 10935 -6649 10991
rect -6593 10935 -6574 10991
rect -11022 10869 -10932 10929
rect -6668 10925 -6574 10935
rect -6664 10871 -6578 10925
rect -11022 10779 -8595 10869
rect -6664 10785 -4371 10871
rect -8685 10686 -8595 10779
rect -8685 10630 -8668 10686
rect -8612 10630 -8595 10686
rect -8685 10604 -8595 10630
rect -4457 10674 -4371 10785
rect -4457 10618 -4442 10674
rect -4386 10618 -4371 10674
rect -4457 10594 -4371 10618
rect -1851 6516 480 6518
rect -1851 6460 -1840 6516
rect -1784 6460 480 6516
rect -1851 6458 480 6460
rect -1566 5556 -1506 5565
rect -1566 5554 2058 5556
rect -1566 5498 -1564 5554
rect -1508 5498 2058 5554
rect -1566 5496 2058 5498
rect -1566 5487 -1506 5496
rect -10744 3789 -10642 3794
rect -6568 3791 -6474 3796
rect -10748 3771 -10638 3789
rect -10748 3715 -10721 3771
rect -10665 3715 -10638 3771
rect -10748 3697 -10638 3715
rect -6572 3777 -6470 3791
rect -6572 3721 -6549 3777
rect -6493 3721 -6470 3777
rect -6572 3707 -6470 3721
rect -10744 3649 -10642 3697
rect -10744 3547 -8631 3649
rect -8733 3462 -8631 3547
rect -6568 3639 -6474 3707
rect -6568 3545 -4455 3639
rect -8733 3406 -8710 3462
rect -8654 3406 -8631 3462
rect -8733 3374 -8631 3406
rect -4549 3454 -4455 3545
rect -4549 3398 -4530 3454
rect -4474 3398 -4455 3454
rect -4549 3370 -4455 3398
<< via2 >>
rect -4456 30284 -4400 30286
rect -4456 30232 -4454 30284
rect -4454 30232 -4402 30284
rect -4402 30232 -4400 30284
rect -4456 30230 -4400 30232
rect -13286 15504 -13230 15560
rect -9664 15504 -9608 15560
rect -12484 15355 -12428 15411
rect -9848 15355 -9792 15411
rect -13088 14498 -13032 14554
rect -9852 14498 -9796 14554
rect -13482 14276 -13426 14332
rect -9664 14276 -9608 14332
rect -11005 10941 -10949 10997
rect -6649 10935 -6593 10991
rect -8668 10630 -8612 10686
rect -4442 10618 -4386 10674
rect -1840 6460 -1784 6516
rect -1564 5498 -1508 5554
rect -10721 3715 -10665 3771
rect -6549 3721 -6493 3777
rect -8710 3406 -8654 3462
rect -4530 3398 -4474 3454
<< metal3 >>
rect -4486 30293 -4350 30322
rect -4486 30229 -4460 30293
rect -4396 30229 -4350 30293
rect -4486 30192 -4350 30229
rect -13310 15560 -13210 15584
rect -13310 15504 -13286 15560
rect -13230 15504 -13210 15560
rect -13504 14332 -13404 14354
rect -13504 14276 -13482 14332
rect -13426 14276 -13404 14332
rect -13504 3497 -13404 14276
rect -13310 5903 -13210 15504
rect -9686 15560 -9586 15580
rect -9686 15504 -9664 15560
rect -9608 15504 -9586 15560
rect -12510 15411 -12410 15434
rect -12510 15355 -12484 15411
rect -12428 15355 -12410 15411
rect -12510 14670 -12410 15355
rect -12510 14606 -12492 14670
rect -12428 14606 -12410 14670
rect -12510 14582 -12410 14606
rect -9874 15411 -9774 15436
rect -9874 15355 -9848 15411
rect -9792 15355 -9774 15411
rect -9874 14581 -9774 15355
rect -13110 14554 -13010 14576
rect -13110 14498 -13088 14554
rect -13032 14498 -13010 14554
rect -13110 10725 -13010 14498
rect -9879 14554 -9769 14581
rect -9879 14498 -9852 14554
rect -9796 14498 -9769 14554
rect -9879 14471 -9769 14498
rect -9686 14359 -9586 15504
rect 10952 14470 11052 14476
rect -1600 14452 11052 14470
rect -1600 14388 10970 14452
rect 11034 14388 11052 14452
rect -1600 14370 11052 14388
rect -9691 14332 -9581 14359
rect -9691 14276 -9664 14332
rect -9608 14276 -9581 14332
rect -9691 14249 -9581 14276
rect -11124 14101 -10954 14120
rect -11124 14012 -11111 14101
rect -12012 14010 -11111 14012
rect -12572 13957 -11111 14010
rect -10967 14012 -10954 14101
rect -8772 14110 -8612 14124
rect -8772 14012 -8764 14110
rect -10967 13966 -8764 14012
rect -8620 14012 -8612 14110
rect -6398 14083 -6256 14128
rect -6398 14019 -6359 14083
rect -6295 14019 -6256 14083
rect -6398 14012 -6256 14019
rect -4024 14097 -3862 14112
rect -4024 14012 -4015 14097
rect -8620 13966 -4015 14012
rect -10967 13957 -4015 13966
rect -12572 13953 -4015 13957
rect -3871 14012 -3862 14097
rect -3871 14010 -2864 14012
rect -3871 13953 -2610 14010
rect -12572 13408 -2610 13953
rect -12572 11918 -11971 13408
rect -10026 13056 -7214 13156
rect -10026 12694 -9896 13056
rect -7314 12716 -7214 13056
rect -10026 12562 -9926 12694
rect -12700 11901 -11971 11918
rect -12700 11837 -12677 11901
rect -12613 11837 -11971 11901
rect -12700 11820 -11971 11837
rect -13115 10708 -13005 10725
rect -13115 10644 -13092 10708
rect -13028 10644 -13005 10708
rect -13115 10627 -13005 10644
rect -13110 10626 -13010 10627
rect -12572 9826 -11971 11820
rect -3213 11908 -2610 13408
rect -1858 12903 -1758 12904
rect -1863 12886 -1753 12903
rect -1863 12822 -1840 12886
rect -1776 12822 -1753 12886
rect -1863 12805 -1753 12822
rect -3213 11879 -2434 11908
rect -3213 11815 -2533 11879
rect -2469 11815 -2434 11879
rect -3213 11786 -2434 11815
rect -11022 10997 -10932 11046
rect -9332 11021 -9232 11294
rect -5192 11029 -5092 11278
rect -11022 10941 -11005 10997
rect -10949 10941 -10932 10997
rect -11022 10924 -10932 10941
rect -9337 11004 -9227 11021
rect -9337 10940 -9314 11004
rect -9250 10940 -9227 11004
rect -9337 10923 -9227 10940
rect -6664 10991 -6578 11028
rect -6664 10935 -6649 10991
rect -6593 10935 -6578 10991
rect -9332 10922 -9232 10923
rect -6664 10920 -6578 10935
rect -5197 11012 -5087 11029
rect -5197 10948 -5174 11012
rect -5110 10948 -5087 11012
rect -5197 10931 -5087 10948
rect -5192 10930 -5092 10931
rect -8101 10882 -8003 10887
rect -7570 10882 -7470 10888
rect -8102 10864 -7470 10882
rect -3901 10880 -3803 10885
rect -3400 10880 -3300 10886
rect -8102 10800 -8084 10864
rect -8020 10800 -7552 10864
rect -7488 10800 -7470 10864
rect -8102 10782 -7470 10800
rect -8101 10777 -8003 10782
rect -7570 10776 -7470 10782
rect -3902 10862 -3300 10880
rect -3902 10798 -3884 10862
rect -3820 10798 -3382 10862
rect -3318 10798 -3300 10862
rect -3902 10780 -3300 10798
rect -3901 10775 -3803 10780
rect -3400 10774 -3300 10780
rect -10156 10725 -10056 10726
rect -5956 10725 -5856 10726
rect -10161 10708 -10051 10725
rect -5961 10708 -5851 10725
rect -10161 10644 -10138 10708
rect -10074 10644 -10051 10708
rect -10161 10627 -10051 10644
rect -8690 10686 -8590 10708
rect -8690 10630 -8668 10686
rect -8612 10630 -8590 10686
rect -10156 10588 -10056 10627
rect -8690 10608 -8590 10630
rect -5961 10644 -5938 10708
rect -5874 10644 -5851 10708
rect -5961 10627 -5851 10644
rect -4462 10674 -4366 10694
rect -10156 10476 -10002 10588
rect -12678 9799 -11971 9826
rect -12678 9735 -12645 9799
rect -12581 9735 -11971 9799
rect -12678 9708 -11971 9735
rect -13100 8615 -13000 8616
rect -13105 8598 -12995 8615
rect -13105 8534 -13082 8598
rect -13018 8534 -12995 8598
rect -13105 8517 -12995 8534
rect -13315 5886 -13205 5903
rect -13315 5822 -13292 5886
rect -13228 5822 -13205 5886
rect -13315 5805 -13205 5822
rect -13310 5804 -13210 5805
rect -13509 3480 -13399 3497
rect -13509 3416 -13486 3480
rect -13422 3416 -13399 3480
rect -13509 3399 -13399 3416
rect -13504 3398 -13404 3399
rect -13100 1627 -13000 8517
rect -12572 8256 -11971 9708
rect -10102 8616 -10002 10476
rect -8685 10421 -8595 10608
rect -5956 10476 -5856 10627
rect -4462 10618 -4442 10674
rect -4386 10618 -4366 10674
rect -4462 10598 -4366 10618
rect -4457 10357 -4371 10598
rect -3213 9850 -2610 11786
rect -3213 9828 -2420 9850
rect -3213 9764 -2512 9828
rect -2448 9764 -2420 9828
rect -3213 9742 -2420 9764
rect -7192 8616 -7092 9154
rect -10510 8598 -7092 8616
rect -10510 8534 -10486 8598
rect -10422 8534 -7092 8598
rect -10510 8516 -7092 8534
rect -3213 8256 -2610 9742
rect -12572 7654 -2610 8256
rect -12572 7652 -2956 7654
rect -11068 7558 -10886 7652
rect -11068 7414 -11049 7558
rect -10905 7414 -10886 7558
rect -11068 7402 -10886 7414
rect -8768 7558 -8586 7652
rect -8768 7414 -8749 7558
rect -8605 7414 -8586 7558
rect -8768 7402 -8586 7414
rect -6468 7558 -6286 7652
rect -6468 7414 -6449 7558
rect -6305 7414 -6286 7558
rect -6468 7402 -6286 7414
rect -4048 7558 -3866 7652
rect -4048 7414 -4029 7558
rect -3885 7414 -3866 7558
rect -4048 7402 -3866 7414
rect -11062 7401 -10892 7402
rect -8762 7401 -8592 7402
rect -6462 7401 -6292 7402
rect -4042 7401 -3872 7402
rect -11062 6871 -10892 6890
rect -11062 6782 -11049 6871
rect -11950 6778 -11049 6782
rect -12509 6727 -11049 6778
rect -10905 6782 -10892 6871
rect -8762 6871 -8592 6890
rect -8762 6782 -8749 6871
rect -10905 6727 -8749 6782
rect -8605 6782 -8592 6871
rect -6462 6871 -6292 6890
rect -6462 6782 -6449 6871
rect -8605 6727 -6449 6782
rect -6305 6782 -6292 6871
rect -4042 6871 -3872 6890
rect -4042 6782 -4029 6871
rect -6305 6727 -4029 6782
rect -3885 6782 -3872 6871
rect -3885 6778 -2802 6782
rect -3885 6727 -2548 6778
rect -12509 6178 -2548 6727
rect -12509 4688 -11909 6178
rect -11530 5886 -7198 5904
rect -11530 5822 -11506 5886
rect -11442 5822 -7198 5886
rect -11530 5804 -7198 5822
rect -10006 5428 -9906 5804
rect -7298 5478 -7198 5804
rect -12638 4671 -11909 4688
rect -12638 4607 -12615 4671
rect -12551 4607 -11909 4671
rect -12638 4590 -11909 4607
rect -12509 2596 -11909 4590
rect -3151 4678 -2548 6178
rect -1858 6516 -1758 12805
rect -1600 8863 -1500 14370
rect 10952 14364 11052 14370
rect -1605 8846 -1495 8863
rect -1605 8782 -1582 8846
rect -1518 8782 -1495 8846
rect -1605 8765 -1495 8782
rect -1600 8764 -1500 8765
rect -1858 6460 -1840 6516
rect -1784 6460 -1758 6516
rect -1858 5665 -1758 6460
rect -1863 5648 -1753 5665
rect -1863 5584 -1840 5648
rect -1776 5584 -1753 5648
rect -1863 5567 -1753 5584
rect -1858 5566 -1758 5567
rect -1586 5554 -1486 5594
rect -1586 5498 -1564 5554
rect -1508 5498 -1486 5554
rect -3151 4649 -2372 4678
rect -3151 4585 -2471 4649
rect -2407 4585 -2372 4649
rect -3151 4556 -2372 4585
rect -10744 3771 -10642 3844
rect -9304 3797 -9204 4022
rect -10744 3715 -10721 3771
rect -10665 3715 -10642 3771
rect -10744 3692 -10642 3715
rect -9309 3780 -9199 3797
rect -9309 3716 -9286 3780
rect -9222 3716 -9199 3780
rect -9309 3699 -9199 3716
rect -6568 3777 -6474 3830
rect -5084 3801 -4984 4060
rect -6568 3721 -6549 3777
rect -6493 3721 -6474 3777
rect -6568 3702 -6474 3721
rect -5089 3784 -4979 3801
rect -5089 3720 -5066 3784
rect -5002 3720 -4979 3784
rect -5089 3703 -4979 3720
rect -5084 3702 -4984 3703
rect -9304 3698 -9204 3699
rect -8085 3644 -7987 3649
rect -7554 3644 -7454 3650
rect -3845 3644 -3747 3649
rect -3344 3644 -3244 3650
rect -8086 3626 -7454 3644
rect -8086 3562 -8068 3626
rect -8004 3562 -7536 3626
rect -7472 3562 -7454 3626
rect -8086 3544 -7454 3562
rect -3846 3626 -3244 3644
rect -3846 3562 -3828 3626
rect -3764 3562 -3326 3626
rect -3262 3562 -3244 3626
rect -3846 3544 -3244 3562
rect -8085 3539 -7987 3544
rect -7554 3538 -7454 3544
rect -3845 3539 -3747 3544
rect -3344 3538 -3244 3544
rect -5940 3501 -5840 3502
rect -10180 3497 -10080 3498
rect -10185 3480 -10075 3497
rect -10185 3416 -10162 3480
rect -10098 3416 -10075 3480
rect -10185 3399 -10075 3416
rect -8738 3462 -8626 3490
rect -8738 3406 -8710 3462
rect -8654 3406 -8626 3462
rect -5945 3484 -5835 3501
rect -10180 3350 -10080 3399
rect -8738 3378 -8626 3406
rect -10180 3238 -10026 3350
rect -12616 2569 -11909 2596
rect -12616 2505 -12583 2569
rect -12519 2505 -11909 2569
rect -12616 2478 -11909 2505
rect -13103 1610 -12993 1627
rect -13103 1546 -13080 1610
rect -13016 1546 -12993 1610
rect -13103 1529 -12993 1546
rect -13100 1528 -13000 1529
rect -12509 1028 -11909 2478
rect -10126 1378 -10026 3238
rect -8733 3109 -8631 3378
rect -7176 3254 -7174 3446
rect -5945 3420 -5922 3484
rect -5858 3420 -5835 3484
rect -5945 3403 -5835 3420
rect -4554 3454 -4450 3478
rect -5940 3238 -5840 3403
rect -4554 3398 -4530 3454
rect -4474 3398 -4450 3454
rect -4554 3374 -4450 3398
rect -4549 3065 -4455 3374
rect -3151 2620 -2548 4556
rect -3151 2598 -2358 2620
rect -3151 2534 -2450 2598
rect -2386 2534 -2358 2598
rect -3151 2512 -2358 2534
rect -7176 1378 -7076 1916
rect -10126 1278 -7076 1378
rect -3151 1028 -2548 2512
rect -1586 1625 -1486 5498
rect -1591 1608 -1481 1625
rect -1591 1544 -1568 1608
rect -1504 1544 -1481 1608
rect -1591 1527 -1481 1544
rect -1586 1526 -1486 1527
rect -12509 468 -2548 1028
rect -12509 422 -11078 468
rect -11094 324 -11078 422
rect -10934 422 -8666 468
rect -10934 324 -10918 422
rect -11094 302 -10918 324
rect -8682 324 -8666 422
rect -8522 422 -6346 468
rect -8522 324 -8506 422
rect -8682 302 -8506 324
rect -6362 324 -6346 422
rect -6202 422 -3946 468
rect -6202 324 -6186 422
rect -6362 302 -6186 324
rect -3962 324 -3946 422
rect -3802 424 -2548 468
rect -3802 422 -3061 424
rect -3802 324 -3786 422
rect -3962 302 -3786 324
<< via3 >>
rect -4460 30286 -4396 30293
rect -4460 30230 -4456 30286
rect -4456 30230 -4400 30286
rect -4400 30230 -4396 30286
rect -4460 30229 -4396 30230
rect -12492 14606 -12428 14670
rect 10970 14388 11034 14452
rect -11111 13957 -10967 14101
rect -8764 13966 -8620 14110
rect -6359 14019 -6295 14083
rect -4015 13953 -3871 14097
rect -12677 11837 -12613 11901
rect -13092 10644 -13028 10708
rect -1840 12822 -1776 12886
rect -2533 11815 -2469 11879
rect -9314 10940 -9250 11004
rect -5174 10948 -5110 11012
rect -8084 10800 -8020 10864
rect -7552 10800 -7488 10864
rect -3884 10798 -3820 10862
rect -3382 10798 -3318 10862
rect -10138 10644 -10074 10708
rect -5938 10644 -5874 10708
rect -12645 9735 -12581 9799
rect -13082 8534 -13018 8598
rect -13292 5822 -13228 5886
rect -13486 3416 -13422 3480
rect -2512 9764 -2448 9828
rect -10486 8534 -10422 8598
rect -11049 7414 -10905 7558
rect -8749 7414 -8605 7558
rect -6449 7414 -6305 7558
rect -4029 7414 -3885 7558
rect -11049 6727 -10905 6871
rect -8749 6727 -8605 6871
rect -6449 6727 -6305 6871
rect -4029 6727 -3885 6871
rect -11506 5822 -11442 5886
rect -12615 4607 -12551 4671
rect -1582 8782 -1518 8846
rect -1840 5584 -1776 5648
rect -2471 4585 -2407 4649
rect -9286 3716 -9222 3780
rect -5066 3720 -5002 3784
rect -8068 3562 -8004 3626
rect -7536 3562 -7472 3626
rect -3828 3562 -3764 3626
rect -3326 3562 -3262 3626
rect -10162 3416 -10098 3480
rect -12583 2505 -12519 2569
rect -13080 1546 -13016 1610
rect -5922 3420 -5858 3484
rect -2450 2534 -2386 2598
rect -1568 1544 -1504 1608
rect -11078 324 -10934 468
rect -8666 324 -8522 468
rect -6346 324 -6202 468
rect -3946 324 -3802 468
<< metal4 >>
rect -4928 30293 -3252 30940
rect -4928 30229 -4460 30293
rect -4396 30229 -3252 30293
rect -4928 30140 -3252 30229
rect -12511 14670 -12409 14689
rect -12511 14606 -12492 14670
rect -12428 14606 -12409 14670
rect -12511 14587 -12409 14606
rect -12510 13220 -12410 14587
rect 10952 14471 11052 15140
rect 10951 14452 11053 14471
rect 10951 14388 10970 14452
rect 11034 14388 11053 14452
rect 10951 14369 11053 14388
rect -11125 14101 -10953 14115
rect -11125 13957 -11111 14101
rect -10967 13957 -10953 14101
rect -8773 14110 -8611 14119
rect -8773 13966 -8764 14110
rect -8620 13966 -8611 14110
rect -6399 14083 -6255 14123
rect -6399 14019 -6359 14083
rect -6295 14019 -6255 14083
rect -6399 13979 -6255 14019
rect -4025 14097 -3861 14107
rect -8773 13957 -8611 13966
rect -11125 13943 -10953 13957
rect -11124 13605 -10954 13943
rect -8772 13654 -8612 13957
rect -6398 13705 -6256 13979
rect -4025 13953 -4015 14097
rect -3871 13953 -3861 14097
rect -4025 13943 -3861 13953
rect -4024 13667 -3862 13943
rect -12510 13120 -10034 13220
rect -10134 12904 -10034 13120
rect -10134 12886 -1758 12904
rect -10134 12822 -1840 12886
rect -1776 12822 -1758 12886
rect -10134 12804 -1758 12822
rect -10134 12450 -10034 12804
rect -12695 11918 -12595 11919
rect -12695 11901 -12243 11918
rect -12695 11837 -12677 11901
rect -12613 11837 -12243 11901
rect -12695 11820 -12243 11837
rect -12695 11819 -12595 11820
rect -8246 11784 -7706 11884
rect -9332 11004 -9232 11022
rect -9332 10940 -9314 11004
rect -9250 10940 -9232 11004
rect -9332 10726 -9232 10940
rect -13110 10708 -9232 10726
rect -13110 10644 -13092 10708
rect -13028 10644 -10138 10708
rect -10074 10644 -9232 10708
rect -13110 10626 -9232 10644
rect -8102 10864 -8002 10882
rect -8102 10800 -8084 10864
rect -8020 10800 -8002 10864
rect -8102 10382 -8002 10800
rect -12673 9826 -12553 9827
rect -12673 9799 -12205 9826
rect -12673 9735 -12645 9799
rect -12581 9735 -12205 9799
rect -12673 9708 -12205 9735
rect -12673 9707 -12553 9708
rect -10152 8864 -10052 9244
rect -7806 8864 -7706 11784
rect -7570 10883 -7470 12804
rect -5934 12450 -5834 12804
rect -4046 11784 -3506 11884
rect -5192 11012 -5092 11030
rect -5192 10948 -5174 11012
rect -5110 10948 -5092 11012
rect -7571 10864 -7469 10883
rect -7571 10800 -7552 10864
rect -7488 10800 -7469 10864
rect -7571 10781 -7469 10800
rect -5192 10726 -5092 10948
rect -5956 10708 -5092 10726
rect -5956 10644 -5938 10708
rect -5874 10644 -5092 10708
rect -5956 10626 -5092 10644
rect -3902 10862 -3802 10880
rect -3902 10798 -3884 10862
rect -3820 10798 -3802 10862
rect -3902 10382 -3802 10798
rect -5952 8864 -5852 9244
rect -3606 8864 -3506 11784
rect -3400 10881 -3300 12804
rect -2563 11908 -2439 11909
rect -2879 11879 -2439 11908
rect -2879 11815 -2533 11879
rect -2469 11815 -2439 11879
rect -2879 11786 -2439 11815
rect -2563 11785 -2439 11786
rect -3401 10862 -3299 10881
rect -3401 10798 -3382 10862
rect -3318 10798 -3299 10862
rect -3401 10779 -3299 10798
rect -2535 9850 -2425 9851
rect -2922 9828 -2425 9850
rect -2922 9764 -2512 9828
rect -2448 9764 -2425 9828
rect -2922 9742 -2425 9764
rect -2535 9741 -2425 9742
rect -10152 8846 -1500 8864
rect -10152 8782 -1582 8846
rect -1518 8782 -1500 8846
rect -10152 8764 -1500 8782
rect -10505 8616 -10403 8617
rect -13100 8598 -10403 8616
rect -13100 8534 -13082 8598
rect -13018 8534 -10486 8598
rect -10422 8534 -10403 8598
rect -13100 8516 -10403 8534
rect -10505 8515 -10403 8516
rect -11062 7558 -10892 7927
rect -11062 7414 -11049 7558
rect -10905 7414 -10892 7558
rect -11062 6885 -10892 7414
rect -8762 7558 -8592 7927
rect -8762 7414 -8749 7558
rect -8605 7414 -8592 7558
rect -8762 6885 -8592 7414
rect -6462 7558 -6292 7927
rect -6462 7414 -6449 7558
rect -6305 7414 -6292 7558
rect -6462 6885 -6292 7414
rect -4042 7558 -3872 7927
rect -4042 7414 -4029 7558
rect -3885 7414 -3872 7558
rect -4042 6885 -3872 7414
rect -11063 6871 -10891 6885
rect -11063 6727 -11049 6871
rect -10905 6727 -10891 6871
rect -11063 6713 -10891 6727
rect -8763 6871 -8591 6885
rect -8763 6727 -8749 6871
rect -8605 6727 -8591 6871
rect -8763 6713 -8591 6727
rect -6463 6871 -6291 6885
rect -6463 6727 -6449 6871
rect -6305 6727 -6291 6871
rect -6463 6713 -6291 6727
rect -4043 6871 -3871 6885
rect -4043 6727 -4029 6871
rect -3885 6727 -3871 6871
rect -4043 6713 -3871 6727
rect -11062 6375 -10892 6713
rect -8762 6375 -8592 6713
rect -6462 6375 -6292 6713
rect -4042 6375 -3872 6713
rect -11525 5904 -11423 5905
rect -13310 5886 -11423 5904
rect -13310 5822 -13292 5886
rect -13228 5822 -11506 5886
rect -11442 5822 -11423 5886
rect -13310 5804 -11423 5822
rect -11525 5803 -11423 5804
rect -10158 5648 -1758 5666
rect -10158 5584 -1840 5648
rect -1776 5584 -1758 5648
rect -10158 5566 -1758 5584
rect -10158 5212 -10058 5566
rect -12633 4688 -12533 4689
rect -12633 4671 -12181 4688
rect -12633 4607 -12615 4671
rect -12551 4607 -12181 4671
rect -12633 4590 -12181 4607
rect -12633 4589 -12533 4590
rect -8230 4546 -7690 4646
rect -9304 3780 -9204 3798
rect -9304 3716 -9286 3780
rect -9222 3716 -9204 3780
rect -9304 3498 -9204 3716
rect -13504 3480 -9204 3498
rect -13504 3416 -13486 3480
rect -13422 3416 -10162 3480
rect -10098 3416 -9204 3480
rect -13504 3398 -9204 3416
rect -8086 3626 -7986 3644
rect -8086 3562 -8068 3626
rect -8004 3562 -7986 3626
rect -8086 3144 -7986 3562
rect -12611 2596 -12491 2597
rect -12611 2569 -12143 2596
rect -12611 2505 -12583 2569
rect -12519 2505 -12143 2569
rect -12611 2478 -12143 2505
rect -12611 2477 -12491 2478
rect -10176 1628 -10076 2006
rect -13098 1626 -9512 1628
rect -7790 1626 -7690 4546
rect -7554 3645 -7454 5566
rect -5918 5212 -5818 5566
rect -3990 4546 -3450 4646
rect -5084 3784 -4984 3802
rect -5084 3720 -5066 3784
rect -5002 3720 -4984 3784
rect -7555 3626 -7453 3645
rect -7555 3562 -7536 3626
rect -7472 3562 -7453 3626
rect -7555 3543 -7453 3562
rect -5084 3502 -4984 3720
rect -5940 3484 -4984 3502
rect -5940 3420 -5922 3484
rect -5858 3420 -4984 3484
rect -5940 3402 -4984 3420
rect -3846 3626 -3746 3644
rect -3846 3562 -3828 3626
rect -3764 3562 -3746 3626
rect -3846 3144 -3746 3562
rect -5936 1626 -5836 2006
rect -3550 1626 -3450 4546
rect -3344 3645 -3244 5566
rect -2501 4678 -2377 4679
rect -2817 4649 -2377 4678
rect -2817 4585 -2471 4649
rect -2407 4585 -2377 4649
rect -2817 4556 -2377 4585
rect -2501 4555 -2377 4556
rect -3345 3626 -3243 3645
rect -3345 3562 -3326 3626
rect -3262 3562 -3243 3626
rect -3345 3543 -3243 3562
rect -2473 2620 -2363 2621
rect -2860 2598 -2363 2620
rect -2860 2534 -2450 2598
rect -2386 2534 -2363 2598
rect -2860 2512 -2363 2534
rect -2473 2511 -2363 2512
rect -13098 1610 -1486 1626
rect -13098 1546 -13080 1610
rect -13016 1608 -1486 1610
rect -13016 1546 -1568 1608
rect -13098 1544 -1568 1546
rect -1504 1544 -1486 1608
rect -13098 1528 -1486 1544
rect -10176 1526 -1486 1528
rect -11094 485 -10918 750
rect -8682 485 -8506 750
rect -6362 485 -6186 750
rect -3962 485 -3786 750
rect -11095 468 -10917 485
rect -11095 324 -11078 468
rect -10934 324 -10917 468
rect -11095 307 -10917 324
rect -8683 468 -8505 485
rect -8683 324 -8666 468
rect -8522 324 -8505 468
rect -8683 307 -8505 324
rect -6363 468 -6185 485
rect -6363 324 -6346 468
rect -6202 324 -6185 468
rect -6363 307 -6185 324
rect -3963 468 -3785 485
rect -3963 324 -3946 468
rect -3802 324 -3785 468
rect -3963 307 -3785 324
rect -11094 140 -10918 307
rect -8682 140 -8506 307
rect -6362 140 -6186 307
rect -3962 140 -3786 307
rect -13514 -660 -1808 140
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_7
timestamp 1626486988
transform -1 0 -11077 0 1 724
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_7
timestamp 1626486988
transform 1 0 -12158 0 1 2542
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_15
timestamp 1626486988
transform 1 0 -10672 0 1 2546
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_14
timestamp 1626486988
transform 1 0 -8632 0 1 2546
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_7
timestamp 1626486988
transform 1 0 -8594 0 1 724
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_6
timestamp 1626486988
transform 1 0 -3823 0 1 726
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_13
timestamp 1626486988
transform 1 0 -4392 0 1 2546
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_12
timestamp 1626486988
transform 1 0 -6432 0 1 2546
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_6
timestamp 1626486988
transform -1 0 -6306 0 1 726
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_6
timestamp 1626486988
transform -1 0 -2902 0 1 2544
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_5
timestamp 1626486988
transform -1 0 -11077 0 1 6480
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_4
timestamp 1626486988
transform -1 0 -11139 0 1 7954
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_5
timestamp 1626486988
transform 1 0 -12158 0 1 4646
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_11
timestamp 1626486988
transform 1 0 -10672 0 1 4646
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_10
timestamp 1626486988
transform 1 0 -8632 0 1 4646
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_5
timestamp 1626486988
transform 1 0 -8656 0 1 7954
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_4
timestamp 1626486988
transform 1 0 -8594 0 1 6480
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_3
timestamp 1626486988
transform 1 0 -3885 0 1 7956
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_2
timestamp 1626486988
transform 1 0 -3823 0 1 6482
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_9
timestamp 1626486988
transform 1 0 -4392 0 1 4646
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_8
timestamp 1626486988
transform 1 0 -6432 0 1 4646
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_3
timestamp 1626486988
transform -1 0 -6368 0 1 7956
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_2
timestamp 1626486988
transform -1 0 -6306 0 1 6482
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_4
timestamp 1626486988
transform -1 0 -2902 0 1 4648
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_3
timestamp 1626486988
transform 1 0 -12220 0 1 11876
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_2
timestamp 1626486988
transform 1 0 -12220 0 1 9772
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_7
timestamp 1626486988
transform 1 0 -8694 0 1 11876
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_6
timestamp 1626486988
transform 1 0 -10734 0 1 11876
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_5
timestamp 1626486988
transform 1 0 -8694 0 1 9776
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_4
timestamp 1626486988
transform 1 0 -10734 0 1 9776
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_3
timestamp 1626486988
transform 1 0 -4454 0 1 11876
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_2
timestamp 1626486988
transform 1 0 -6494 0 1 11876
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_1
timestamp 1626486988
transform 1 0 -4454 0 1 9776
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_0
timestamp 1626486988
transform 1 0 -6494 0 1 9776
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_1
timestamp 1626486988
transform -1 0 -2964 0 1 11878
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_0
timestamp 1626486988
transform -1 0 -2964 0 1 9774
box -350 -900 244 900
use txgate  txgate_1
timestamp 1626486988
transform 1 0 -83901 0 1 -42680
box 74185 57360 76542 59116
use txgate  txgate_0
timestamp 1626486988
transform 1 0 -86501 0 1 -42680
box 74185 57360 76542 59116
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_1
timestamp 1626486988
transform -1 0 -11139 0 1 13710
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_1
timestamp 1626486988
transform 1 0 -8656 0 1 13710
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_0
timestamp 1626486988
transform 1 0 -3885 0 1 13712
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_0
timestamp 1626486988
transform -1 0 -6368 0 1 13712
box -950 -300 818 300
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1626486988
transform -1 0 -7070 0 1 15246
box -38 -48 314 592
use se_fold_casc_wide_swing_ota  se_fold_casc_wide_swing_ota_0
timestamp 1626486988
transform 1 0 10912 0 1 26540
box -15168 -27248 25000 4400
<< labels >>
flabel metal4 s -5616 -342 -5562 -296 1 FreeSans 600 0 0 0 VSS
flabel metal4 s -9816 8794 -9798 8822 1 FreeSans 600 0 0 0 vse
flabel metal4 s -9746 12834 -9732 12846 1 FreeSans 600 0 0 0 vip
flabel metal1 s 704 1582 716 1600 1 FreeSans 600 0 0 0 ibiasn
flabel metal4 s -4738 30526 -4712 30558 1 FreeSans 600 0 0 0 VDD
flabel metal1 s -7056 15480 -7054 15484 1 FreeSans 600 0 0 0 rst_n
flabel metal1 s -7332 15474 -7328 15480 1 FreeSans 600 0 0 0 rst
flabel metal3 s -9542 5852 -9520 5872 1 FreeSans 600 0 0 0 vdiffp
flabel metal4 s -9702 5600 -9680 5618 1 FreeSans 600 0 0 0 vip
flabel metal4 s -9786 1568 -9770 1582 1 FreeSans 600 0 0 0 vim
flabel metal3 s -9812 1318 -9800 1332 1 FreeSans 600 0 0 0 vdiffm
flabel metal3 s -9752 13102 -9732 13118 1 FreeSans 600 0 0 0 vocm
flabel metal3 s -9862 8562 -9854 8578 1 FreeSans 600 0 0 0 vim
<< end >>
