magic
tech sky130A
magscale 1 2
timestamp 1621146761
<< nwell >>
rect -676 -519 676 519
<< pmoslvt >>
rect -480 -300 480 300
<< pdiff >>
rect -538 288 -480 300
rect -538 -288 -526 288
rect -492 -288 -480 288
rect -538 -300 -480 -288
rect 480 288 538 300
rect 480 -288 492 288
rect 526 -288 538 288
rect 480 -300 538 -288
<< pdiffc >>
rect -526 -288 -492 288
rect 492 -288 526 288
<< nsubdiff >>
rect -640 449 -544 483
rect 544 449 640 483
rect -640 387 -606 449
rect 606 387 640 449
rect -640 -449 -606 -387
rect 606 -449 640 -387
rect -640 -483 -544 -449
rect 544 -483 640 -449
<< nsubdiffcont >>
rect -544 449 544 483
rect -640 -387 -606 387
rect 606 -387 640 387
rect -544 -483 544 -449
<< poly >>
rect -294 381 294 397
rect -294 364 -278 381
rect -480 347 -278 364
rect 278 364 294 381
rect 278 347 480 364
rect -480 300 480 347
rect -480 -347 480 -300
rect -480 -364 -278 -347
rect -294 -381 -278 -364
rect 278 -364 480 -347
rect 278 -381 294 -364
rect -294 -397 294 -381
<< polycont >>
rect -278 347 278 381
rect -278 -381 278 -347
<< locali >>
rect -640 449 -544 483
rect 544 449 640 483
rect -640 387 -606 449
rect 606 387 640 449
rect -294 347 -278 381
rect 278 347 294 381
rect -526 288 -492 304
rect -526 -304 -492 -288
rect 492 288 526 304
rect 492 -304 526 -288
rect -294 -381 -278 -347
rect 278 -381 294 -347
rect -640 -449 -606 -387
rect 606 -449 640 -387
rect -640 -483 -544 -449
rect 544 -483 640 -449
<< viali >>
rect -232 347 232 381
rect -526 -288 -492 288
rect 492 -288 526 288
rect -232 -381 232 -347
<< metal1 >>
rect -244 381 244 387
rect -244 347 -232 381
rect 232 347 244 381
rect -244 341 244 347
rect -532 288 -486 300
rect -532 -288 -526 288
rect -492 -288 -486 288
rect -532 -300 -486 -288
rect 486 288 532 300
rect 486 -288 492 288
rect 526 -288 532 288
rect 486 -300 532 -288
rect -244 -347 244 -341
rect -244 -381 -232 -347
rect 232 -381 244 -347
rect -244 -387 244 -381
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -623 -466 623 466
string parameters w 3 l 4.8 m 1 nf 1 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
