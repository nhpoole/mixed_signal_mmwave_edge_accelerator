* Stimulus file.

.include ../layouts/gm_c_stage/gm_c_stage_pex.spice
.include gm_c_stage_lvs.spice

.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_01v8/sky130_fd_pr__esd_nfet_01v8__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_pfet_g5v0d10v5/sky130_fd_pr__esd_pfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d16v0/sky130_fd_pr__pfet_g5v0d16v0__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d16v0/sky130_fd_pr__nfet_g5v0d16v0__tt_discrete.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_g5v0d10v5/sky130_fd_pr__esd_nfet_g5v0d10v5__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/nonfet.spice
* Mismatch parameters
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__mismatch.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice
* Resistor~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/Capacitor
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical__lin.spice
* Special cells
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/specialized_cells.spice
* All models
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/all.spice
* Corner
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/rf.spice

.param vdd=1.8 ibias=10u vincm=1.1 vsig=0 vcmdes=1.1

vdd VDD VSS 'vdd'
vss VSS GND 0
vip vip VSS dc 'vincm+vsig' ac 1 0
vim vim VSS dc 'vincm-vsig'
vocm vocm VSS 'vcmdes'
i1 vdd ibiasn 'ibias'
x1 vip vim vocm vop vom ibiasn VDD VSS gm_c_stage_flat
*x1 vip vim vocm vop vom ibiasn VDD VSS gm_c_stage_lvs

*.op
*.print all
*write gm_c_stage_lvs_op.raw

* Control Block 1
*.control
*    op
*    print all
*    *ac dec 100 0.1 1g
*    noise v(vop, vom) vip dec 100 1 100k
*    run
*    *write gm_c_stage_lvs_ac.raw
*    *setplot noise1
*    *write gm_c_stage_lvs_noise1.raw v(onoise_spectrum) v(inoise_spectrum)
*    setplot noise2
*    write gm_c_stage_lvs_noise2.raw v(onoise_total) v(inoise_total)
*    quit
*.endc

* Control Block 2
.ac dec 100 0.1 1g
*.noise v(vop, vom) vip dec 100 1 100k
.control
    let incm = 0.4
    while incm < 1.6
        set incm = $&incm
        alter @vip[dc]=$incm
        alter @vim[dc]=$incm
        run
        write gm_c_stage_lvs_ac_{$incm}.raw
        *setplot noise1
        *write gm_c_stage_lvs_noise1_{$incm}.raw v(onoise_spectrum) v(inoise_spectrum)
        *setplot noise2
        *write gm_c_stage_lvs_noise2_{$incm}.raw v(onoise_total) v(inoise_total)
        let incm = incm + 0.1
    end
    alter @vip[dc]=0.7
    alter @vim[dc]=0.7
    op
    print all
    quit
.endc

* Control Block 3
*.ac dec 100 0.1 1g
*.control
*    let temperature = -40
*    while temperature < 130
*        set temp = $&temperature
*        run
*        write gm_c_stage_lvs_temp_{$temp}.raw
*        let temperature = temperature + 10
*    end
*    quit
*.endc

* Control Block 4
*.ac dec 100 0.1 1g
*.control
*    let supply = 1.62
*    while supply < 2
*        alterparam vdd = {$&supply}
*        reset
*        run
*        write gm_c_stage_lvs_vdd_{$&supply}.raw
*        let supply = supply + 0.04
*    end
*    quit
*.endc

