magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -6914 -1648 6914 1648
<< pwell >>
rect -5654 -326 5654 326
<< nmoslvt >>
rect -5570 -300 -4610 300
rect -4552 -300 -3592 300
rect -3534 -300 -2574 300
rect -2516 -300 -1556 300
rect -1498 -300 -538 300
rect -480 -300 480 300
rect 538 -300 1498 300
rect 1556 -300 2516 300
rect 2574 -300 3534 300
rect 3592 -300 4552 300
rect 4610 -300 5570 300
<< ndiff >>
rect -5628 255 -5570 300
rect -5628 221 -5616 255
rect -5582 221 -5570 255
rect -5628 187 -5570 221
rect -5628 153 -5616 187
rect -5582 153 -5570 187
rect -5628 119 -5570 153
rect -5628 85 -5616 119
rect -5582 85 -5570 119
rect -5628 51 -5570 85
rect -5628 17 -5616 51
rect -5582 17 -5570 51
rect -5628 -17 -5570 17
rect -5628 -51 -5616 -17
rect -5582 -51 -5570 -17
rect -5628 -85 -5570 -51
rect -5628 -119 -5616 -85
rect -5582 -119 -5570 -85
rect -5628 -153 -5570 -119
rect -5628 -187 -5616 -153
rect -5582 -187 -5570 -153
rect -5628 -221 -5570 -187
rect -5628 -255 -5616 -221
rect -5582 -255 -5570 -221
rect -5628 -300 -5570 -255
rect -4610 255 -4552 300
rect -4610 221 -4598 255
rect -4564 221 -4552 255
rect -4610 187 -4552 221
rect -4610 153 -4598 187
rect -4564 153 -4552 187
rect -4610 119 -4552 153
rect -4610 85 -4598 119
rect -4564 85 -4552 119
rect -4610 51 -4552 85
rect -4610 17 -4598 51
rect -4564 17 -4552 51
rect -4610 -17 -4552 17
rect -4610 -51 -4598 -17
rect -4564 -51 -4552 -17
rect -4610 -85 -4552 -51
rect -4610 -119 -4598 -85
rect -4564 -119 -4552 -85
rect -4610 -153 -4552 -119
rect -4610 -187 -4598 -153
rect -4564 -187 -4552 -153
rect -4610 -221 -4552 -187
rect -4610 -255 -4598 -221
rect -4564 -255 -4552 -221
rect -4610 -300 -4552 -255
rect -3592 255 -3534 300
rect -3592 221 -3580 255
rect -3546 221 -3534 255
rect -3592 187 -3534 221
rect -3592 153 -3580 187
rect -3546 153 -3534 187
rect -3592 119 -3534 153
rect -3592 85 -3580 119
rect -3546 85 -3534 119
rect -3592 51 -3534 85
rect -3592 17 -3580 51
rect -3546 17 -3534 51
rect -3592 -17 -3534 17
rect -3592 -51 -3580 -17
rect -3546 -51 -3534 -17
rect -3592 -85 -3534 -51
rect -3592 -119 -3580 -85
rect -3546 -119 -3534 -85
rect -3592 -153 -3534 -119
rect -3592 -187 -3580 -153
rect -3546 -187 -3534 -153
rect -3592 -221 -3534 -187
rect -3592 -255 -3580 -221
rect -3546 -255 -3534 -221
rect -3592 -300 -3534 -255
rect -2574 255 -2516 300
rect -2574 221 -2562 255
rect -2528 221 -2516 255
rect -2574 187 -2516 221
rect -2574 153 -2562 187
rect -2528 153 -2516 187
rect -2574 119 -2516 153
rect -2574 85 -2562 119
rect -2528 85 -2516 119
rect -2574 51 -2516 85
rect -2574 17 -2562 51
rect -2528 17 -2516 51
rect -2574 -17 -2516 17
rect -2574 -51 -2562 -17
rect -2528 -51 -2516 -17
rect -2574 -85 -2516 -51
rect -2574 -119 -2562 -85
rect -2528 -119 -2516 -85
rect -2574 -153 -2516 -119
rect -2574 -187 -2562 -153
rect -2528 -187 -2516 -153
rect -2574 -221 -2516 -187
rect -2574 -255 -2562 -221
rect -2528 -255 -2516 -221
rect -2574 -300 -2516 -255
rect -1556 255 -1498 300
rect -1556 221 -1544 255
rect -1510 221 -1498 255
rect -1556 187 -1498 221
rect -1556 153 -1544 187
rect -1510 153 -1498 187
rect -1556 119 -1498 153
rect -1556 85 -1544 119
rect -1510 85 -1498 119
rect -1556 51 -1498 85
rect -1556 17 -1544 51
rect -1510 17 -1498 51
rect -1556 -17 -1498 17
rect -1556 -51 -1544 -17
rect -1510 -51 -1498 -17
rect -1556 -85 -1498 -51
rect -1556 -119 -1544 -85
rect -1510 -119 -1498 -85
rect -1556 -153 -1498 -119
rect -1556 -187 -1544 -153
rect -1510 -187 -1498 -153
rect -1556 -221 -1498 -187
rect -1556 -255 -1544 -221
rect -1510 -255 -1498 -221
rect -1556 -300 -1498 -255
rect -538 255 -480 300
rect -538 221 -526 255
rect -492 221 -480 255
rect -538 187 -480 221
rect -538 153 -526 187
rect -492 153 -480 187
rect -538 119 -480 153
rect -538 85 -526 119
rect -492 85 -480 119
rect -538 51 -480 85
rect -538 17 -526 51
rect -492 17 -480 51
rect -538 -17 -480 17
rect -538 -51 -526 -17
rect -492 -51 -480 -17
rect -538 -85 -480 -51
rect -538 -119 -526 -85
rect -492 -119 -480 -85
rect -538 -153 -480 -119
rect -538 -187 -526 -153
rect -492 -187 -480 -153
rect -538 -221 -480 -187
rect -538 -255 -526 -221
rect -492 -255 -480 -221
rect -538 -300 -480 -255
rect 480 255 538 300
rect 480 221 492 255
rect 526 221 538 255
rect 480 187 538 221
rect 480 153 492 187
rect 526 153 538 187
rect 480 119 538 153
rect 480 85 492 119
rect 526 85 538 119
rect 480 51 538 85
rect 480 17 492 51
rect 526 17 538 51
rect 480 -17 538 17
rect 480 -51 492 -17
rect 526 -51 538 -17
rect 480 -85 538 -51
rect 480 -119 492 -85
rect 526 -119 538 -85
rect 480 -153 538 -119
rect 480 -187 492 -153
rect 526 -187 538 -153
rect 480 -221 538 -187
rect 480 -255 492 -221
rect 526 -255 538 -221
rect 480 -300 538 -255
rect 1498 255 1556 300
rect 1498 221 1510 255
rect 1544 221 1556 255
rect 1498 187 1556 221
rect 1498 153 1510 187
rect 1544 153 1556 187
rect 1498 119 1556 153
rect 1498 85 1510 119
rect 1544 85 1556 119
rect 1498 51 1556 85
rect 1498 17 1510 51
rect 1544 17 1556 51
rect 1498 -17 1556 17
rect 1498 -51 1510 -17
rect 1544 -51 1556 -17
rect 1498 -85 1556 -51
rect 1498 -119 1510 -85
rect 1544 -119 1556 -85
rect 1498 -153 1556 -119
rect 1498 -187 1510 -153
rect 1544 -187 1556 -153
rect 1498 -221 1556 -187
rect 1498 -255 1510 -221
rect 1544 -255 1556 -221
rect 1498 -300 1556 -255
rect 2516 255 2574 300
rect 2516 221 2528 255
rect 2562 221 2574 255
rect 2516 187 2574 221
rect 2516 153 2528 187
rect 2562 153 2574 187
rect 2516 119 2574 153
rect 2516 85 2528 119
rect 2562 85 2574 119
rect 2516 51 2574 85
rect 2516 17 2528 51
rect 2562 17 2574 51
rect 2516 -17 2574 17
rect 2516 -51 2528 -17
rect 2562 -51 2574 -17
rect 2516 -85 2574 -51
rect 2516 -119 2528 -85
rect 2562 -119 2574 -85
rect 2516 -153 2574 -119
rect 2516 -187 2528 -153
rect 2562 -187 2574 -153
rect 2516 -221 2574 -187
rect 2516 -255 2528 -221
rect 2562 -255 2574 -221
rect 2516 -300 2574 -255
rect 3534 255 3592 300
rect 3534 221 3546 255
rect 3580 221 3592 255
rect 3534 187 3592 221
rect 3534 153 3546 187
rect 3580 153 3592 187
rect 3534 119 3592 153
rect 3534 85 3546 119
rect 3580 85 3592 119
rect 3534 51 3592 85
rect 3534 17 3546 51
rect 3580 17 3592 51
rect 3534 -17 3592 17
rect 3534 -51 3546 -17
rect 3580 -51 3592 -17
rect 3534 -85 3592 -51
rect 3534 -119 3546 -85
rect 3580 -119 3592 -85
rect 3534 -153 3592 -119
rect 3534 -187 3546 -153
rect 3580 -187 3592 -153
rect 3534 -221 3592 -187
rect 3534 -255 3546 -221
rect 3580 -255 3592 -221
rect 3534 -300 3592 -255
rect 4552 255 4610 300
rect 4552 221 4564 255
rect 4598 221 4610 255
rect 4552 187 4610 221
rect 4552 153 4564 187
rect 4598 153 4610 187
rect 4552 119 4610 153
rect 4552 85 4564 119
rect 4598 85 4610 119
rect 4552 51 4610 85
rect 4552 17 4564 51
rect 4598 17 4610 51
rect 4552 -17 4610 17
rect 4552 -51 4564 -17
rect 4598 -51 4610 -17
rect 4552 -85 4610 -51
rect 4552 -119 4564 -85
rect 4598 -119 4610 -85
rect 4552 -153 4610 -119
rect 4552 -187 4564 -153
rect 4598 -187 4610 -153
rect 4552 -221 4610 -187
rect 4552 -255 4564 -221
rect 4598 -255 4610 -221
rect 4552 -300 4610 -255
rect 5570 255 5628 300
rect 5570 221 5582 255
rect 5616 221 5628 255
rect 5570 187 5628 221
rect 5570 153 5582 187
rect 5616 153 5628 187
rect 5570 119 5628 153
rect 5570 85 5582 119
rect 5616 85 5628 119
rect 5570 51 5628 85
rect 5570 17 5582 51
rect 5616 17 5628 51
rect 5570 -17 5628 17
rect 5570 -51 5582 -17
rect 5616 -51 5628 -17
rect 5570 -85 5628 -51
rect 5570 -119 5582 -85
rect 5616 -119 5628 -85
rect 5570 -153 5628 -119
rect 5570 -187 5582 -153
rect 5616 -187 5628 -153
rect 5570 -221 5628 -187
rect 5570 -255 5582 -221
rect 5616 -255 5628 -221
rect 5570 -300 5628 -255
<< ndiffc >>
rect -5616 221 -5582 255
rect -5616 153 -5582 187
rect -5616 85 -5582 119
rect -5616 17 -5582 51
rect -5616 -51 -5582 -17
rect -5616 -119 -5582 -85
rect -5616 -187 -5582 -153
rect -5616 -255 -5582 -221
rect -4598 221 -4564 255
rect -4598 153 -4564 187
rect -4598 85 -4564 119
rect -4598 17 -4564 51
rect -4598 -51 -4564 -17
rect -4598 -119 -4564 -85
rect -4598 -187 -4564 -153
rect -4598 -255 -4564 -221
rect -3580 221 -3546 255
rect -3580 153 -3546 187
rect -3580 85 -3546 119
rect -3580 17 -3546 51
rect -3580 -51 -3546 -17
rect -3580 -119 -3546 -85
rect -3580 -187 -3546 -153
rect -3580 -255 -3546 -221
rect -2562 221 -2528 255
rect -2562 153 -2528 187
rect -2562 85 -2528 119
rect -2562 17 -2528 51
rect -2562 -51 -2528 -17
rect -2562 -119 -2528 -85
rect -2562 -187 -2528 -153
rect -2562 -255 -2528 -221
rect -1544 221 -1510 255
rect -1544 153 -1510 187
rect -1544 85 -1510 119
rect -1544 17 -1510 51
rect -1544 -51 -1510 -17
rect -1544 -119 -1510 -85
rect -1544 -187 -1510 -153
rect -1544 -255 -1510 -221
rect -526 221 -492 255
rect -526 153 -492 187
rect -526 85 -492 119
rect -526 17 -492 51
rect -526 -51 -492 -17
rect -526 -119 -492 -85
rect -526 -187 -492 -153
rect -526 -255 -492 -221
rect 492 221 526 255
rect 492 153 526 187
rect 492 85 526 119
rect 492 17 526 51
rect 492 -51 526 -17
rect 492 -119 526 -85
rect 492 -187 526 -153
rect 492 -255 526 -221
rect 1510 221 1544 255
rect 1510 153 1544 187
rect 1510 85 1544 119
rect 1510 17 1544 51
rect 1510 -51 1544 -17
rect 1510 -119 1544 -85
rect 1510 -187 1544 -153
rect 1510 -255 1544 -221
rect 2528 221 2562 255
rect 2528 153 2562 187
rect 2528 85 2562 119
rect 2528 17 2562 51
rect 2528 -51 2562 -17
rect 2528 -119 2562 -85
rect 2528 -187 2562 -153
rect 2528 -255 2562 -221
rect 3546 221 3580 255
rect 3546 153 3580 187
rect 3546 85 3580 119
rect 3546 17 3580 51
rect 3546 -51 3580 -17
rect 3546 -119 3580 -85
rect 3546 -187 3580 -153
rect 3546 -255 3580 -221
rect 4564 221 4598 255
rect 4564 153 4598 187
rect 4564 85 4598 119
rect 4564 17 4598 51
rect 4564 -51 4598 -17
rect 4564 -119 4598 -85
rect 4564 -187 4598 -153
rect 4564 -255 4598 -221
rect 5582 221 5616 255
rect 5582 153 5616 187
rect 5582 85 5616 119
rect 5582 17 5616 51
rect 5582 -51 5616 -17
rect 5582 -119 5616 -85
rect 5582 -187 5616 -153
rect 5582 -255 5616 -221
<< poly >>
rect -5384 372 -4796 388
rect -5384 355 -5345 372
rect -5570 338 -5345 355
rect -5311 338 -5277 372
rect -5243 338 -5209 372
rect -5175 338 -5141 372
rect -5107 338 -5073 372
rect -5039 338 -5005 372
rect -4971 338 -4937 372
rect -4903 338 -4869 372
rect -4835 355 -4796 372
rect -4366 372 -3778 388
rect -4366 355 -4327 372
rect -4835 338 -4610 355
rect -5570 300 -4610 338
rect -4552 338 -4327 355
rect -4293 338 -4259 372
rect -4225 338 -4191 372
rect -4157 338 -4123 372
rect -4089 338 -4055 372
rect -4021 338 -3987 372
rect -3953 338 -3919 372
rect -3885 338 -3851 372
rect -3817 355 -3778 372
rect -3348 372 -2760 388
rect -3348 355 -3309 372
rect -3817 338 -3592 355
rect -4552 300 -3592 338
rect -3534 338 -3309 355
rect -3275 338 -3241 372
rect -3207 338 -3173 372
rect -3139 338 -3105 372
rect -3071 338 -3037 372
rect -3003 338 -2969 372
rect -2935 338 -2901 372
rect -2867 338 -2833 372
rect -2799 355 -2760 372
rect -2330 372 -1742 388
rect -2330 355 -2291 372
rect -2799 338 -2574 355
rect -3534 300 -2574 338
rect -2516 338 -2291 355
rect -2257 338 -2223 372
rect -2189 338 -2155 372
rect -2121 338 -2087 372
rect -2053 338 -2019 372
rect -1985 338 -1951 372
rect -1917 338 -1883 372
rect -1849 338 -1815 372
rect -1781 355 -1742 372
rect -1312 372 -724 388
rect -1312 355 -1273 372
rect -1781 338 -1556 355
rect -2516 300 -1556 338
rect -1498 338 -1273 355
rect -1239 338 -1205 372
rect -1171 338 -1137 372
rect -1103 338 -1069 372
rect -1035 338 -1001 372
rect -967 338 -933 372
rect -899 338 -865 372
rect -831 338 -797 372
rect -763 355 -724 372
rect -294 372 294 388
rect -294 355 -255 372
rect -763 338 -538 355
rect -1498 300 -538 338
rect -480 338 -255 355
rect -221 338 -187 372
rect -153 338 -119 372
rect -85 338 -51 372
rect -17 338 17 372
rect 51 338 85 372
rect 119 338 153 372
rect 187 338 221 372
rect 255 355 294 372
rect 724 372 1312 388
rect 724 355 763 372
rect 255 338 480 355
rect -480 300 480 338
rect 538 338 763 355
rect 797 338 831 372
rect 865 338 899 372
rect 933 338 967 372
rect 1001 338 1035 372
rect 1069 338 1103 372
rect 1137 338 1171 372
rect 1205 338 1239 372
rect 1273 355 1312 372
rect 1742 372 2330 388
rect 1742 355 1781 372
rect 1273 338 1498 355
rect 538 300 1498 338
rect 1556 338 1781 355
rect 1815 338 1849 372
rect 1883 338 1917 372
rect 1951 338 1985 372
rect 2019 338 2053 372
rect 2087 338 2121 372
rect 2155 338 2189 372
rect 2223 338 2257 372
rect 2291 355 2330 372
rect 2760 372 3348 388
rect 2760 355 2799 372
rect 2291 338 2516 355
rect 1556 300 2516 338
rect 2574 338 2799 355
rect 2833 338 2867 372
rect 2901 338 2935 372
rect 2969 338 3003 372
rect 3037 338 3071 372
rect 3105 338 3139 372
rect 3173 338 3207 372
rect 3241 338 3275 372
rect 3309 355 3348 372
rect 3778 372 4366 388
rect 3778 355 3817 372
rect 3309 338 3534 355
rect 2574 300 3534 338
rect 3592 338 3817 355
rect 3851 338 3885 372
rect 3919 338 3953 372
rect 3987 338 4021 372
rect 4055 338 4089 372
rect 4123 338 4157 372
rect 4191 338 4225 372
rect 4259 338 4293 372
rect 4327 355 4366 372
rect 4796 372 5384 388
rect 4796 355 4835 372
rect 4327 338 4552 355
rect 3592 300 4552 338
rect 4610 338 4835 355
rect 4869 338 4903 372
rect 4937 338 4971 372
rect 5005 338 5039 372
rect 5073 338 5107 372
rect 5141 338 5175 372
rect 5209 338 5243 372
rect 5277 338 5311 372
rect 5345 355 5384 372
rect 5345 338 5570 355
rect 4610 300 5570 338
rect -5570 -338 -4610 -300
rect -5570 -355 -5345 -338
rect -5384 -372 -5345 -355
rect -5311 -372 -5277 -338
rect -5243 -372 -5209 -338
rect -5175 -372 -5141 -338
rect -5107 -372 -5073 -338
rect -5039 -372 -5005 -338
rect -4971 -372 -4937 -338
rect -4903 -372 -4869 -338
rect -4835 -355 -4610 -338
rect -4552 -338 -3592 -300
rect -4552 -355 -4327 -338
rect -4835 -372 -4796 -355
rect -5384 -388 -4796 -372
rect -4366 -372 -4327 -355
rect -4293 -372 -4259 -338
rect -4225 -372 -4191 -338
rect -4157 -372 -4123 -338
rect -4089 -372 -4055 -338
rect -4021 -372 -3987 -338
rect -3953 -372 -3919 -338
rect -3885 -372 -3851 -338
rect -3817 -355 -3592 -338
rect -3534 -338 -2574 -300
rect -3534 -355 -3309 -338
rect -3817 -372 -3778 -355
rect -4366 -388 -3778 -372
rect -3348 -372 -3309 -355
rect -3275 -372 -3241 -338
rect -3207 -372 -3173 -338
rect -3139 -372 -3105 -338
rect -3071 -372 -3037 -338
rect -3003 -372 -2969 -338
rect -2935 -372 -2901 -338
rect -2867 -372 -2833 -338
rect -2799 -355 -2574 -338
rect -2516 -338 -1556 -300
rect -2516 -355 -2291 -338
rect -2799 -372 -2760 -355
rect -3348 -388 -2760 -372
rect -2330 -372 -2291 -355
rect -2257 -372 -2223 -338
rect -2189 -372 -2155 -338
rect -2121 -372 -2087 -338
rect -2053 -372 -2019 -338
rect -1985 -372 -1951 -338
rect -1917 -372 -1883 -338
rect -1849 -372 -1815 -338
rect -1781 -355 -1556 -338
rect -1498 -338 -538 -300
rect -1498 -355 -1273 -338
rect -1781 -372 -1742 -355
rect -2330 -388 -1742 -372
rect -1312 -372 -1273 -355
rect -1239 -372 -1205 -338
rect -1171 -372 -1137 -338
rect -1103 -372 -1069 -338
rect -1035 -372 -1001 -338
rect -967 -372 -933 -338
rect -899 -372 -865 -338
rect -831 -372 -797 -338
rect -763 -355 -538 -338
rect -480 -338 480 -300
rect -480 -355 -255 -338
rect -763 -372 -724 -355
rect -1312 -388 -724 -372
rect -294 -372 -255 -355
rect -221 -372 -187 -338
rect -153 -372 -119 -338
rect -85 -372 -51 -338
rect -17 -372 17 -338
rect 51 -372 85 -338
rect 119 -372 153 -338
rect 187 -372 221 -338
rect 255 -355 480 -338
rect 538 -338 1498 -300
rect 538 -355 763 -338
rect 255 -372 294 -355
rect -294 -388 294 -372
rect 724 -372 763 -355
rect 797 -372 831 -338
rect 865 -372 899 -338
rect 933 -372 967 -338
rect 1001 -372 1035 -338
rect 1069 -372 1103 -338
rect 1137 -372 1171 -338
rect 1205 -372 1239 -338
rect 1273 -355 1498 -338
rect 1556 -338 2516 -300
rect 1556 -355 1781 -338
rect 1273 -372 1312 -355
rect 724 -388 1312 -372
rect 1742 -372 1781 -355
rect 1815 -372 1849 -338
rect 1883 -372 1917 -338
rect 1951 -372 1985 -338
rect 2019 -372 2053 -338
rect 2087 -372 2121 -338
rect 2155 -372 2189 -338
rect 2223 -372 2257 -338
rect 2291 -355 2516 -338
rect 2574 -338 3534 -300
rect 2574 -355 2799 -338
rect 2291 -372 2330 -355
rect 1742 -388 2330 -372
rect 2760 -372 2799 -355
rect 2833 -372 2867 -338
rect 2901 -372 2935 -338
rect 2969 -372 3003 -338
rect 3037 -372 3071 -338
rect 3105 -372 3139 -338
rect 3173 -372 3207 -338
rect 3241 -372 3275 -338
rect 3309 -355 3534 -338
rect 3592 -338 4552 -300
rect 3592 -355 3817 -338
rect 3309 -372 3348 -355
rect 2760 -388 3348 -372
rect 3778 -372 3817 -355
rect 3851 -372 3885 -338
rect 3919 -372 3953 -338
rect 3987 -372 4021 -338
rect 4055 -372 4089 -338
rect 4123 -372 4157 -338
rect 4191 -372 4225 -338
rect 4259 -372 4293 -338
rect 4327 -355 4552 -338
rect 4610 -338 5570 -300
rect 4610 -355 4835 -338
rect 4327 -372 4366 -355
rect 3778 -388 4366 -372
rect 4796 -372 4835 -355
rect 4869 -372 4903 -338
rect 4937 -372 4971 -338
rect 5005 -372 5039 -338
rect 5073 -372 5107 -338
rect 5141 -372 5175 -338
rect 5209 -372 5243 -338
rect 5277 -372 5311 -338
rect 5345 -355 5570 -338
rect 5345 -372 5384 -355
rect 4796 -388 5384 -372
<< polycont >>
rect -5345 338 -5311 372
rect -5277 338 -5243 372
rect -5209 338 -5175 372
rect -5141 338 -5107 372
rect -5073 338 -5039 372
rect -5005 338 -4971 372
rect -4937 338 -4903 372
rect -4869 338 -4835 372
rect -4327 338 -4293 372
rect -4259 338 -4225 372
rect -4191 338 -4157 372
rect -4123 338 -4089 372
rect -4055 338 -4021 372
rect -3987 338 -3953 372
rect -3919 338 -3885 372
rect -3851 338 -3817 372
rect -3309 338 -3275 372
rect -3241 338 -3207 372
rect -3173 338 -3139 372
rect -3105 338 -3071 372
rect -3037 338 -3003 372
rect -2969 338 -2935 372
rect -2901 338 -2867 372
rect -2833 338 -2799 372
rect -2291 338 -2257 372
rect -2223 338 -2189 372
rect -2155 338 -2121 372
rect -2087 338 -2053 372
rect -2019 338 -1985 372
rect -1951 338 -1917 372
rect -1883 338 -1849 372
rect -1815 338 -1781 372
rect -1273 338 -1239 372
rect -1205 338 -1171 372
rect -1137 338 -1103 372
rect -1069 338 -1035 372
rect -1001 338 -967 372
rect -933 338 -899 372
rect -865 338 -831 372
rect -797 338 -763 372
rect -255 338 -221 372
rect -187 338 -153 372
rect -119 338 -85 372
rect -51 338 -17 372
rect 17 338 51 372
rect 85 338 119 372
rect 153 338 187 372
rect 221 338 255 372
rect 763 338 797 372
rect 831 338 865 372
rect 899 338 933 372
rect 967 338 1001 372
rect 1035 338 1069 372
rect 1103 338 1137 372
rect 1171 338 1205 372
rect 1239 338 1273 372
rect 1781 338 1815 372
rect 1849 338 1883 372
rect 1917 338 1951 372
rect 1985 338 2019 372
rect 2053 338 2087 372
rect 2121 338 2155 372
rect 2189 338 2223 372
rect 2257 338 2291 372
rect 2799 338 2833 372
rect 2867 338 2901 372
rect 2935 338 2969 372
rect 3003 338 3037 372
rect 3071 338 3105 372
rect 3139 338 3173 372
rect 3207 338 3241 372
rect 3275 338 3309 372
rect 3817 338 3851 372
rect 3885 338 3919 372
rect 3953 338 3987 372
rect 4021 338 4055 372
rect 4089 338 4123 372
rect 4157 338 4191 372
rect 4225 338 4259 372
rect 4293 338 4327 372
rect 4835 338 4869 372
rect 4903 338 4937 372
rect 4971 338 5005 372
rect 5039 338 5073 372
rect 5107 338 5141 372
rect 5175 338 5209 372
rect 5243 338 5277 372
rect 5311 338 5345 372
rect -5345 -372 -5311 -338
rect -5277 -372 -5243 -338
rect -5209 -372 -5175 -338
rect -5141 -372 -5107 -338
rect -5073 -372 -5039 -338
rect -5005 -372 -4971 -338
rect -4937 -372 -4903 -338
rect -4869 -372 -4835 -338
rect -4327 -372 -4293 -338
rect -4259 -372 -4225 -338
rect -4191 -372 -4157 -338
rect -4123 -372 -4089 -338
rect -4055 -372 -4021 -338
rect -3987 -372 -3953 -338
rect -3919 -372 -3885 -338
rect -3851 -372 -3817 -338
rect -3309 -372 -3275 -338
rect -3241 -372 -3207 -338
rect -3173 -372 -3139 -338
rect -3105 -372 -3071 -338
rect -3037 -372 -3003 -338
rect -2969 -372 -2935 -338
rect -2901 -372 -2867 -338
rect -2833 -372 -2799 -338
rect -2291 -372 -2257 -338
rect -2223 -372 -2189 -338
rect -2155 -372 -2121 -338
rect -2087 -372 -2053 -338
rect -2019 -372 -1985 -338
rect -1951 -372 -1917 -338
rect -1883 -372 -1849 -338
rect -1815 -372 -1781 -338
rect -1273 -372 -1239 -338
rect -1205 -372 -1171 -338
rect -1137 -372 -1103 -338
rect -1069 -372 -1035 -338
rect -1001 -372 -967 -338
rect -933 -372 -899 -338
rect -865 -372 -831 -338
rect -797 -372 -763 -338
rect -255 -372 -221 -338
rect -187 -372 -153 -338
rect -119 -372 -85 -338
rect -51 -372 -17 -338
rect 17 -372 51 -338
rect 85 -372 119 -338
rect 153 -372 187 -338
rect 221 -372 255 -338
rect 763 -372 797 -338
rect 831 -372 865 -338
rect 899 -372 933 -338
rect 967 -372 1001 -338
rect 1035 -372 1069 -338
rect 1103 -372 1137 -338
rect 1171 -372 1205 -338
rect 1239 -372 1273 -338
rect 1781 -372 1815 -338
rect 1849 -372 1883 -338
rect 1917 -372 1951 -338
rect 1985 -372 2019 -338
rect 2053 -372 2087 -338
rect 2121 -372 2155 -338
rect 2189 -372 2223 -338
rect 2257 -372 2291 -338
rect 2799 -372 2833 -338
rect 2867 -372 2901 -338
rect 2935 -372 2969 -338
rect 3003 -372 3037 -338
rect 3071 -372 3105 -338
rect 3139 -372 3173 -338
rect 3207 -372 3241 -338
rect 3275 -372 3309 -338
rect 3817 -372 3851 -338
rect 3885 -372 3919 -338
rect 3953 -372 3987 -338
rect 4021 -372 4055 -338
rect 4089 -372 4123 -338
rect 4157 -372 4191 -338
rect 4225 -372 4259 -338
rect 4293 -372 4327 -338
rect 4835 -372 4869 -338
rect 4903 -372 4937 -338
rect 4971 -372 5005 -338
rect 5039 -372 5073 -338
rect 5107 -372 5141 -338
rect 5175 -372 5209 -338
rect 5243 -372 5277 -338
rect 5311 -372 5345 -338
<< locali >>
rect -5384 338 -5345 372
rect -5311 338 -5287 372
rect -5243 338 -5215 372
rect -5175 338 -5143 372
rect -5107 338 -5073 372
rect -5037 338 -5005 372
rect -4965 338 -4937 372
rect -4893 338 -4869 372
rect -4835 338 -4796 372
rect -4366 338 -4327 372
rect -4293 338 -4269 372
rect -4225 338 -4197 372
rect -4157 338 -4125 372
rect -4089 338 -4055 372
rect -4019 338 -3987 372
rect -3947 338 -3919 372
rect -3875 338 -3851 372
rect -3817 338 -3778 372
rect -3348 338 -3309 372
rect -3275 338 -3251 372
rect -3207 338 -3179 372
rect -3139 338 -3107 372
rect -3071 338 -3037 372
rect -3001 338 -2969 372
rect -2929 338 -2901 372
rect -2857 338 -2833 372
rect -2799 338 -2760 372
rect -2330 338 -2291 372
rect -2257 338 -2233 372
rect -2189 338 -2161 372
rect -2121 338 -2089 372
rect -2053 338 -2019 372
rect -1983 338 -1951 372
rect -1911 338 -1883 372
rect -1839 338 -1815 372
rect -1781 338 -1742 372
rect -1312 338 -1273 372
rect -1239 338 -1215 372
rect -1171 338 -1143 372
rect -1103 338 -1071 372
rect -1035 338 -1001 372
rect -965 338 -933 372
rect -893 338 -865 372
rect -821 338 -797 372
rect -763 338 -724 372
rect -294 338 -255 372
rect -221 338 -197 372
rect -153 338 -125 372
rect -85 338 -53 372
rect -17 338 17 372
rect 53 338 85 372
rect 125 338 153 372
rect 197 338 221 372
rect 255 338 294 372
rect 724 338 763 372
rect 797 338 821 372
rect 865 338 893 372
rect 933 338 965 372
rect 1001 338 1035 372
rect 1071 338 1103 372
rect 1143 338 1171 372
rect 1215 338 1239 372
rect 1273 338 1312 372
rect 1742 338 1781 372
rect 1815 338 1839 372
rect 1883 338 1911 372
rect 1951 338 1983 372
rect 2019 338 2053 372
rect 2089 338 2121 372
rect 2161 338 2189 372
rect 2233 338 2257 372
rect 2291 338 2330 372
rect 2760 338 2799 372
rect 2833 338 2857 372
rect 2901 338 2929 372
rect 2969 338 3001 372
rect 3037 338 3071 372
rect 3107 338 3139 372
rect 3179 338 3207 372
rect 3251 338 3275 372
rect 3309 338 3348 372
rect 3778 338 3817 372
rect 3851 338 3875 372
rect 3919 338 3947 372
rect 3987 338 4019 372
rect 4055 338 4089 372
rect 4125 338 4157 372
rect 4197 338 4225 372
rect 4269 338 4293 372
rect 4327 338 4366 372
rect 4796 338 4835 372
rect 4869 338 4893 372
rect 4937 338 4965 372
rect 5005 338 5037 372
rect 5073 338 5107 372
rect 5143 338 5175 372
rect 5215 338 5243 372
rect 5287 338 5311 372
rect 5345 338 5384 372
rect -5616 269 -5582 304
rect -5616 197 -5582 221
rect -5616 125 -5582 153
rect -5616 53 -5582 85
rect -5616 -17 -5582 17
rect -5616 -85 -5582 -53
rect -5616 -153 -5582 -125
rect -5616 -221 -5582 -197
rect -5616 -304 -5582 -269
rect -4598 269 -4564 304
rect -4598 197 -4564 221
rect -4598 125 -4564 153
rect -4598 53 -4564 85
rect -4598 -17 -4564 17
rect -4598 -85 -4564 -53
rect -4598 -153 -4564 -125
rect -4598 -221 -4564 -197
rect -4598 -304 -4564 -269
rect -3580 269 -3546 304
rect -3580 197 -3546 221
rect -3580 125 -3546 153
rect -3580 53 -3546 85
rect -3580 -17 -3546 17
rect -3580 -85 -3546 -53
rect -3580 -153 -3546 -125
rect -3580 -221 -3546 -197
rect -3580 -304 -3546 -269
rect -2562 269 -2528 304
rect -2562 197 -2528 221
rect -2562 125 -2528 153
rect -2562 53 -2528 85
rect -2562 -17 -2528 17
rect -2562 -85 -2528 -53
rect -2562 -153 -2528 -125
rect -2562 -221 -2528 -197
rect -2562 -304 -2528 -269
rect -1544 269 -1510 304
rect -1544 197 -1510 221
rect -1544 125 -1510 153
rect -1544 53 -1510 85
rect -1544 -17 -1510 17
rect -1544 -85 -1510 -53
rect -1544 -153 -1510 -125
rect -1544 -221 -1510 -197
rect -1544 -304 -1510 -269
rect -526 269 -492 304
rect -526 197 -492 221
rect -526 125 -492 153
rect -526 53 -492 85
rect -526 -17 -492 17
rect -526 -85 -492 -53
rect -526 -153 -492 -125
rect -526 -221 -492 -197
rect -526 -304 -492 -269
rect 492 269 526 304
rect 492 197 526 221
rect 492 125 526 153
rect 492 53 526 85
rect 492 -17 526 17
rect 492 -85 526 -53
rect 492 -153 526 -125
rect 492 -221 526 -197
rect 492 -304 526 -269
rect 1510 269 1544 304
rect 1510 197 1544 221
rect 1510 125 1544 153
rect 1510 53 1544 85
rect 1510 -17 1544 17
rect 1510 -85 1544 -53
rect 1510 -153 1544 -125
rect 1510 -221 1544 -197
rect 1510 -304 1544 -269
rect 2528 269 2562 304
rect 2528 197 2562 221
rect 2528 125 2562 153
rect 2528 53 2562 85
rect 2528 -17 2562 17
rect 2528 -85 2562 -53
rect 2528 -153 2562 -125
rect 2528 -221 2562 -197
rect 2528 -304 2562 -269
rect 3546 269 3580 304
rect 3546 197 3580 221
rect 3546 125 3580 153
rect 3546 53 3580 85
rect 3546 -17 3580 17
rect 3546 -85 3580 -53
rect 3546 -153 3580 -125
rect 3546 -221 3580 -197
rect 3546 -304 3580 -269
rect 4564 269 4598 304
rect 4564 197 4598 221
rect 4564 125 4598 153
rect 4564 53 4598 85
rect 4564 -17 4598 17
rect 4564 -85 4598 -53
rect 4564 -153 4598 -125
rect 4564 -221 4598 -197
rect 4564 -304 4598 -269
rect 5582 269 5616 304
rect 5582 197 5616 221
rect 5582 125 5616 153
rect 5582 53 5616 85
rect 5582 -17 5616 17
rect 5582 -85 5616 -53
rect 5582 -153 5616 -125
rect 5582 -221 5616 -197
rect 5582 -304 5616 -269
rect -5384 -372 -5345 -338
rect -5311 -372 -5287 -338
rect -5243 -372 -5215 -338
rect -5175 -372 -5143 -338
rect -5107 -372 -5073 -338
rect -5037 -372 -5005 -338
rect -4965 -372 -4937 -338
rect -4893 -372 -4869 -338
rect -4835 -372 -4796 -338
rect -4366 -372 -4327 -338
rect -4293 -372 -4269 -338
rect -4225 -372 -4197 -338
rect -4157 -372 -4125 -338
rect -4089 -372 -4055 -338
rect -4019 -372 -3987 -338
rect -3947 -372 -3919 -338
rect -3875 -372 -3851 -338
rect -3817 -372 -3778 -338
rect -3348 -372 -3309 -338
rect -3275 -372 -3251 -338
rect -3207 -372 -3179 -338
rect -3139 -372 -3107 -338
rect -3071 -372 -3037 -338
rect -3001 -372 -2969 -338
rect -2929 -372 -2901 -338
rect -2857 -372 -2833 -338
rect -2799 -372 -2760 -338
rect -2330 -372 -2291 -338
rect -2257 -372 -2233 -338
rect -2189 -372 -2161 -338
rect -2121 -372 -2089 -338
rect -2053 -372 -2019 -338
rect -1983 -372 -1951 -338
rect -1911 -372 -1883 -338
rect -1839 -372 -1815 -338
rect -1781 -372 -1742 -338
rect -1312 -372 -1273 -338
rect -1239 -372 -1215 -338
rect -1171 -372 -1143 -338
rect -1103 -372 -1071 -338
rect -1035 -372 -1001 -338
rect -965 -372 -933 -338
rect -893 -372 -865 -338
rect -821 -372 -797 -338
rect -763 -372 -724 -338
rect -294 -372 -255 -338
rect -221 -372 -197 -338
rect -153 -372 -125 -338
rect -85 -372 -53 -338
rect -17 -372 17 -338
rect 53 -372 85 -338
rect 125 -372 153 -338
rect 197 -372 221 -338
rect 255 -372 294 -338
rect 724 -372 763 -338
rect 797 -372 821 -338
rect 865 -372 893 -338
rect 933 -372 965 -338
rect 1001 -372 1035 -338
rect 1071 -372 1103 -338
rect 1143 -372 1171 -338
rect 1215 -372 1239 -338
rect 1273 -372 1312 -338
rect 1742 -372 1781 -338
rect 1815 -372 1839 -338
rect 1883 -372 1911 -338
rect 1951 -372 1983 -338
rect 2019 -372 2053 -338
rect 2089 -372 2121 -338
rect 2161 -372 2189 -338
rect 2233 -372 2257 -338
rect 2291 -372 2330 -338
rect 2760 -372 2799 -338
rect 2833 -372 2857 -338
rect 2901 -372 2929 -338
rect 2969 -372 3001 -338
rect 3037 -372 3071 -338
rect 3107 -372 3139 -338
rect 3179 -372 3207 -338
rect 3251 -372 3275 -338
rect 3309 -372 3348 -338
rect 3778 -372 3817 -338
rect 3851 -372 3875 -338
rect 3919 -372 3947 -338
rect 3987 -372 4019 -338
rect 4055 -372 4089 -338
rect 4125 -372 4157 -338
rect 4197 -372 4225 -338
rect 4269 -372 4293 -338
rect 4327 -372 4366 -338
rect 4796 -372 4835 -338
rect 4869 -372 4893 -338
rect 4937 -372 4965 -338
rect 5005 -372 5037 -338
rect 5073 -372 5107 -338
rect 5143 -372 5175 -338
rect 5215 -372 5243 -338
rect 5287 -372 5311 -338
rect 5345 -372 5384 -338
<< viali >>
rect -5287 338 -5277 372
rect -5277 338 -5253 372
rect -5215 338 -5209 372
rect -5209 338 -5181 372
rect -5143 338 -5141 372
rect -5141 338 -5109 372
rect -5071 338 -5039 372
rect -5039 338 -5037 372
rect -4999 338 -4971 372
rect -4971 338 -4965 372
rect -4927 338 -4903 372
rect -4903 338 -4893 372
rect -4269 338 -4259 372
rect -4259 338 -4235 372
rect -4197 338 -4191 372
rect -4191 338 -4163 372
rect -4125 338 -4123 372
rect -4123 338 -4091 372
rect -4053 338 -4021 372
rect -4021 338 -4019 372
rect -3981 338 -3953 372
rect -3953 338 -3947 372
rect -3909 338 -3885 372
rect -3885 338 -3875 372
rect -3251 338 -3241 372
rect -3241 338 -3217 372
rect -3179 338 -3173 372
rect -3173 338 -3145 372
rect -3107 338 -3105 372
rect -3105 338 -3073 372
rect -3035 338 -3003 372
rect -3003 338 -3001 372
rect -2963 338 -2935 372
rect -2935 338 -2929 372
rect -2891 338 -2867 372
rect -2867 338 -2857 372
rect -2233 338 -2223 372
rect -2223 338 -2199 372
rect -2161 338 -2155 372
rect -2155 338 -2127 372
rect -2089 338 -2087 372
rect -2087 338 -2055 372
rect -2017 338 -1985 372
rect -1985 338 -1983 372
rect -1945 338 -1917 372
rect -1917 338 -1911 372
rect -1873 338 -1849 372
rect -1849 338 -1839 372
rect -1215 338 -1205 372
rect -1205 338 -1181 372
rect -1143 338 -1137 372
rect -1137 338 -1109 372
rect -1071 338 -1069 372
rect -1069 338 -1037 372
rect -999 338 -967 372
rect -967 338 -965 372
rect -927 338 -899 372
rect -899 338 -893 372
rect -855 338 -831 372
rect -831 338 -821 372
rect -197 338 -187 372
rect -187 338 -163 372
rect -125 338 -119 372
rect -119 338 -91 372
rect -53 338 -51 372
rect -51 338 -19 372
rect 19 338 51 372
rect 51 338 53 372
rect 91 338 119 372
rect 119 338 125 372
rect 163 338 187 372
rect 187 338 197 372
rect 821 338 831 372
rect 831 338 855 372
rect 893 338 899 372
rect 899 338 927 372
rect 965 338 967 372
rect 967 338 999 372
rect 1037 338 1069 372
rect 1069 338 1071 372
rect 1109 338 1137 372
rect 1137 338 1143 372
rect 1181 338 1205 372
rect 1205 338 1215 372
rect 1839 338 1849 372
rect 1849 338 1873 372
rect 1911 338 1917 372
rect 1917 338 1945 372
rect 1983 338 1985 372
rect 1985 338 2017 372
rect 2055 338 2087 372
rect 2087 338 2089 372
rect 2127 338 2155 372
rect 2155 338 2161 372
rect 2199 338 2223 372
rect 2223 338 2233 372
rect 2857 338 2867 372
rect 2867 338 2891 372
rect 2929 338 2935 372
rect 2935 338 2963 372
rect 3001 338 3003 372
rect 3003 338 3035 372
rect 3073 338 3105 372
rect 3105 338 3107 372
rect 3145 338 3173 372
rect 3173 338 3179 372
rect 3217 338 3241 372
rect 3241 338 3251 372
rect 3875 338 3885 372
rect 3885 338 3909 372
rect 3947 338 3953 372
rect 3953 338 3981 372
rect 4019 338 4021 372
rect 4021 338 4053 372
rect 4091 338 4123 372
rect 4123 338 4125 372
rect 4163 338 4191 372
rect 4191 338 4197 372
rect 4235 338 4259 372
rect 4259 338 4269 372
rect 4893 338 4903 372
rect 4903 338 4927 372
rect 4965 338 4971 372
rect 4971 338 4999 372
rect 5037 338 5039 372
rect 5039 338 5071 372
rect 5109 338 5141 372
rect 5141 338 5143 372
rect 5181 338 5209 372
rect 5209 338 5215 372
rect 5253 338 5277 372
rect 5277 338 5287 372
rect -5616 255 -5582 269
rect -5616 235 -5582 255
rect -5616 187 -5582 197
rect -5616 163 -5582 187
rect -5616 119 -5582 125
rect -5616 91 -5582 119
rect -5616 51 -5582 53
rect -5616 19 -5582 51
rect -5616 -51 -5582 -19
rect -5616 -53 -5582 -51
rect -5616 -119 -5582 -91
rect -5616 -125 -5582 -119
rect -5616 -187 -5582 -163
rect -5616 -197 -5582 -187
rect -5616 -255 -5582 -235
rect -5616 -269 -5582 -255
rect -4598 255 -4564 269
rect -4598 235 -4564 255
rect -4598 187 -4564 197
rect -4598 163 -4564 187
rect -4598 119 -4564 125
rect -4598 91 -4564 119
rect -4598 51 -4564 53
rect -4598 19 -4564 51
rect -4598 -51 -4564 -19
rect -4598 -53 -4564 -51
rect -4598 -119 -4564 -91
rect -4598 -125 -4564 -119
rect -4598 -187 -4564 -163
rect -4598 -197 -4564 -187
rect -4598 -255 -4564 -235
rect -4598 -269 -4564 -255
rect -3580 255 -3546 269
rect -3580 235 -3546 255
rect -3580 187 -3546 197
rect -3580 163 -3546 187
rect -3580 119 -3546 125
rect -3580 91 -3546 119
rect -3580 51 -3546 53
rect -3580 19 -3546 51
rect -3580 -51 -3546 -19
rect -3580 -53 -3546 -51
rect -3580 -119 -3546 -91
rect -3580 -125 -3546 -119
rect -3580 -187 -3546 -163
rect -3580 -197 -3546 -187
rect -3580 -255 -3546 -235
rect -3580 -269 -3546 -255
rect -2562 255 -2528 269
rect -2562 235 -2528 255
rect -2562 187 -2528 197
rect -2562 163 -2528 187
rect -2562 119 -2528 125
rect -2562 91 -2528 119
rect -2562 51 -2528 53
rect -2562 19 -2528 51
rect -2562 -51 -2528 -19
rect -2562 -53 -2528 -51
rect -2562 -119 -2528 -91
rect -2562 -125 -2528 -119
rect -2562 -187 -2528 -163
rect -2562 -197 -2528 -187
rect -2562 -255 -2528 -235
rect -2562 -269 -2528 -255
rect -1544 255 -1510 269
rect -1544 235 -1510 255
rect -1544 187 -1510 197
rect -1544 163 -1510 187
rect -1544 119 -1510 125
rect -1544 91 -1510 119
rect -1544 51 -1510 53
rect -1544 19 -1510 51
rect -1544 -51 -1510 -19
rect -1544 -53 -1510 -51
rect -1544 -119 -1510 -91
rect -1544 -125 -1510 -119
rect -1544 -187 -1510 -163
rect -1544 -197 -1510 -187
rect -1544 -255 -1510 -235
rect -1544 -269 -1510 -255
rect -526 255 -492 269
rect -526 235 -492 255
rect -526 187 -492 197
rect -526 163 -492 187
rect -526 119 -492 125
rect -526 91 -492 119
rect -526 51 -492 53
rect -526 19 -492 51
rect -526 -51 -492 -19
rect -526 -53 -492 -51
rect -526 -119 -492 -91
rect -526 -125 -492 -119
rect -526 -187 -492 -163
rect -526 -197 -492 -187
rect -526 -255 -492 -235
rect -526 -269 -492 -255
rect 492 255 526 269
rect 492 235 526 255
rect 492 187 526 197
rect 492 163 526 187
rect 492 119 526 125
rect 492 91 526 119
rect 492 51 526 53
rect 492 19 526 51
rect 492 -51 526 -19
rect 492 -53 526 -51
rect 492 -119 526 -91
rect 492 -125 526 -119
rect 492 -187 526 -163
rect 492 -197 526 -187
rect 492 -255 526 -235
rect 492 -269 526 -255
rect 1510 255 1544 269
rect 1510 235 1544 255
rect 1510 187 1544 197
rect 1510 163 1544 187
rect 1510 119 1544 125
rect 1510 91 1544 119
rect 1510 51 1544 53
rect 1510 19 1544 51
rect 1510 -51 1544 -19
rect 1510 -53 1544 -51
rect 1510 -119 1544 -91
rect 1510 -125 1544 -119
rect 1510 -187 1544 -163
rect 1510 -197 1544 -187
rect 1510 -255 1544 -235
rect 1510 -269 1544 -255
rect 2528 255 2562 269
rect 2528 235 2562 255
rect 2528 187 2562 197
rect 2528 163 2562 187
rect 2528 119 2562 125
rect 2528 91 2562 119
rect 2528 51 2562 53
rect 2528 19 2562 51
rect 2528 -51 2562 -19
rect 2528 -53 2562 -51
rect 2528 -119 2562 -91
rect 2528 -125 2562 -119
rect 2528 -187 2562 -163
rect 2528 -197 2562 -187
rect 2528 -255 2562 -235
rect 2528 -269 2562 -255
rect 3546 255 3580 269
rect 3546 235 3580 255
rect 3546 187 3580 197
rect 3546 163 3580 187
rect 3546 119 3580 125
rect 3546 91 3580 119
rect 3546 51 3580 53
rect 3546 19 3580 51
rect 3546 -51 3580 -19
rect 3546 -53 3580 -51
rect 3546 -119 3580 -91
rect 3546 -125 3580 -119
rect 3546 -187 3580 -163
rect 3546 -197 3580 -187
rect 3546 -255 3580 -235
rect 3546 -269 3580 -255
rect 4564 255 4598 269
rect 4564 235 4598 255
rect 4564 187 4598 197
rect 4564 163 4598 187
rect 4564 119 4598 125
rect 4564 91 4598 119
rect 4564 51 4598 53
rect 4564 19 4598 51
rect 4564 -51 4598 -19
rect 4564 -53 4598 -51
rect 4564 -119 4598 -91
rect 4564 -125 4598 -119
rect 4564 -187 4598 -163
rect 4564 -197 4598 -187
rect 4564 -255 4598 -235
rect 4564 -269 4598 -255
rect 5582 255 5616 269
rect 5582 235 5616 255
rect 5582 187 5616 197
rect 5582 163 5616 187
rect 5582 119 5616 125
rect 5582 91 5616 119
rect 5582 51 5616 53
rect 5582 19 5616 51
rect 5582 -51 5616 -19
rect 5582 -53 5616 -51
rect 5582 -119 5616 -91
rect 5582 -125 5616 -119
rect 5582 -187 5616 -163
rect 5582 -197 5616 -187
rect 5582 -255 5616 -235
rect 5582 -269 5616 -255
rect -5287 -372 -5277 -338
rect -5277 -372 -5253 -338
rect -5215 -372 -5209 -338
rect -5209 -372 -5181 -338
rect -5143 -372 -5141 -338
rect -5141 -372 -5109 -338
rect -5071 -372 -5039 -338
rect -5039 -372 -5037 -338
rect -4999 -372 -4971 -338
rect -4971 -372 -4965 -338
rect -4927 -372 -4903 -338
rect -4903 -372 -4893 -338
rect -4269 -372 -4259 -338
rect -4259 -372 -4235 -338
rect -4197 -372 -4191 -338
rect -4191 -372 -4163 -338
rect -4125 -372 -4123 -338
rect -4123 -372 -4091 -338
rect -4053 -372 -4021 -338
rect -4021 -372 -4019 -338
rect -3981 -372 -3953 -338
rect -3953 -372 -3947 -338
rect -3909 -372 -3885 -338
rect -3885 -372 -3875 -338
rect -3251 -372 -3241 -338
rect -3241 -372 -3217 -338
rect -3179 -372 -3173 -338
rect -3173 -372 -3145 -338
rect -3107 -372 -3105 -338
rect -3105 -372 -3073 -338
rect -3035 -372 -3003 -338
rect -3003 -372 -3001 -338
rect -2963 -372 -2935 -338
rect -2935 -372 -2929 -338
rect -2891 -372 -2867 -338
rect -2867 -372 -2857 -338
rect -2233 -372 -2223 -338
rect -2223 -372 -2199 -338
rect -2161 -372 -2155 -338
rect -2155 -372 -2127 -338
rect -2089 -372 -2087 -338
rect -2087 -372 -2055 -338
rect -2017 -372 -1985 -338
rect -1985 -372 -1983 -338
rect -1945 -372 -1917 -338
rect -1917 -372 -1911 -338
rect -1873 -372 -1849 -338
rect -1849 -372 -1839 -338
rect -1215 -372 -1205 -338
rect -1205 -372 -1181 -338
rect -1143 -372 -1137 -338
rect -1137 -372 -1109 -338
rect -1071 -372 -1069 -338
rect -1069 -372 -1037 -338
rect -999 -372 -967 -338
rect -967 -372 -965 -338
rect -927 -372 -899 -338
rect -899 -372 -893 -338
rect -855 -372 -831 -338
rect -831 -372 -821 -338
rect -197 -372 -187 -338
rect -187 -372 -163 -338
rect -125 -372 -119 -338
rect -119 -372 -91 -338
rect -53 -372 -51 -338
rect -51 -372 -19 -338
rect 19 -372 51 -338
rect 51 -372 53 -338
rect 91 -372 119 -338
rect 119 -372 125 -338
rect 163 -372 187 -338
rect 187 -372 197 -338
rect 821 -372 831 -338
rect 831 -372 855 -338
rect 893 -372 899 -338
rect 899 -372 927 -338
rect 965 -372 967 -338
rect 967 -372 999 -338
rect 1037 -372 1069 -338
rect 1069 -372 1071 -338
rect 1109 -372 1137 -338
rect 1137 -372 1143 -338
rect 1181 -372 1205 -338
rect 1205 -372 1215 -338
rect 1839 -372 1849 -338
rect 1849 -372 1873 -338
rect 1911 -372 1917 -338
rect 1917 -372 1945 -338
rect 1983 -372 1985 -338
rect 1985 -372 2017 -338
rect 2055 -372 2087 -338
rect 2087 -372 2089 -338
rect 2127 -372 2155 -338
rect 2155 -372 2161 -338
rect 2199 -372 2223 -338
rect 2223 -372 2233 -338
rect 2857 -372 2867 -338
rect 2867 -372 2891 -338
rect 2929 -372 2935 -338
rect 2935 -372 2963 -338
rect 3001 -372 3003 -338
rect 3003 -372 3035 -338
rect 3073 -372 3105 -338
rect 3105 -372 3107 -338
rect 3145 -372 3173 -338
rect 3173 -372 3179 -338
rect 3217 -372 3241 -338
rect 3241 -372 3251 -338
rect 3875 -372 3885 -338
rect 3885 -372 3909 -338
rect 3947 -372 3953 -338
rect 3953 -372 3981 -338
rect 4019 -372 4021 -338
rect 4021 -372 4053 -338
rect 4091 -372 4123 -338
rect 4123 -372 4125 -338
rect 4163 -372 4191 -338
rect 4191 -372 4197 -338
rect 4235 -372 4259 -338
rect 4259 -372 4269 -338
rect 4893 -372 4903 -338
rect 4903 -372 4927 -338
rect 4965 -372 4971 -338
rect 4971 -372 4999 -338
rect 5037 -372 5039 -338
rect 5039 -372 5071 -338
rect 5109 -372 5141 -338
rect 5141 -372 5143 -338
rect 5181 -372 5209 -338
rect 5209 -372 5215 -338
rect 5253 -372 5277 -338
rect 5277 -372 5287 -338
<< metal1 >>
rect -5334 372 -4846 378
rect -5334 338 -5287 372
rect -5253 338 -5215 372
rect -5181 338 -5143 372
rect -5109 338 -5071 372
rect -5037 338 -4999 372
rect -4965 338 -4927 372
rect -4893 338 -4846 372
rect -5334 332 -4846 338
rect -4316 372 -3828 378
rect -4316 338 -4269 372
rect -4235 338 -4197 372
rect -4163 338 -4125 372
rect -4091 338 -4053 372
rect -4019 338 -3981 372
rect -3947 338 -3909 372
rect -3875 338 -3828 372
rect -4316 332 -3828 338
rect -3298 372 -2810 378
rect -3298 338 -3251 372
rect -3217 338 -3179 372
rect -3145 338 -3107 372
rect -3073 338 -3035 372
rect -3001 338 -2963 372
rect -2929 338 -2891 372
rect -2857 338 -2810 372
rect -3298 332 -2810 338
rect -2280 372 -1792 378
rect -2280 338 -2233 372
rect -2199 338 -2161 372
rect -2127 338 -2089 372
rect -2055 338 -2017 372
rect -1983 338 -1945 372
rect -1911 338 -1873 372
rect -1839 338 -1792 372
rect -2280 332 -1792 338
rect -1262 372 -774 378
rect -1262 338 -1215 372
rect -1181 338 -1143 372
rect -1109 338 -1071 372
rect -1037 338 -999 372
rect -965 338 -927 372
rect -893 338 -855 372
rect -821 338 -774 372
rect -1262 332 -774 338
rect -244 372 244 378
rect -244 338 -197 372
rect -163 338 -125 372
rect -91 338 -53 372
rect -19 338 19 372
rect 53 338 91 372
rect 125 338 163 372
rect 197 338 244 372
rect -244 332 244 338
rect 774 372 1262 378
rect 774 338 821 372
rect 855 338 893 372
rect 927 338 965 372
rect 999 338 1037 372
rect 1071 338 1109 372
rect 1143 338 1181 372
rect 1215 338 1262 372
rect 774 332 1262 338
rect 1792 372 2280 378
rect 1792 338 1839 372
rect 1873 338 1911 372
rect 1945 338 1983 372
rect 2017 338 2055 372
rect 2089 338 2127 372
rect 2161 338 2199 372
rect 2233 338 2280 372
rect 1792 332 2280 338
rect 2810 372 3298 378
rect 2810 338 2857 372
rect 2891 338 2929 372
rect 2963 338 3001 372
rect 3035 338 3073 372
rect 3107 338 3145 372
rect 3179 338 3217 372
rect 3251 338 3298 372
rect 2810 332 3298 338
rect 3828 372 4316 378
rect 3828 338 3875 372
rect 3909 338 3947 372
rect 3981 338 4019 372
rect 4053 338 4091 372
rect 4125 338 4163 372
rect 4197 338 4235 372
rect 4269 338 4316 372
rect 3828 332 4316 338
rect 4846 372 5334 378
rect 4846 338 4893 372
rect 4927 338 4965 372
rect 4999 338 5037 372
rect 5071 338 5109 372
rect 5143 338 5181 372
rect 5215 338 5253 372
rect 5287 338 5334 372
rect 4846 332 5334 338
rect -5622 269 -5576 300
rect -5622 235 -5616 269
rect -5582 235 -5576 269
rect -5622 197 -5576 235
rect -5622 163 -5616 197
rect -5582 163 -5576 197
rect -5622 125 -5576 163
rect -5622 91 -5616 125
rect -5582 91 -5576 125
rect -5622 53 -5576 91
rect -5622 19 -5616 53
rect -5582 19 -5576 53
rect -5622 -19 -5576 19
rect -5622 -53 -5616 -19
rect -5582 -53 -5576 -19
rect -5622 -91 -5576 -53
rect -5622 -125 -5616 -91
rect -5582 -125 -5576 -91
rect -5622 -163 -5576 -125
rect -5622 -197 -5616 -163
rect -5582 -197 -5576 -163
rect -5622 -235 -5576 -197
rect -5622 -269 -5616 -235
rect -5582 -269 -5576 -235
rect -5622 -300 -5576 -269
rect -4604 269 -4558 300
rect -4604 235 -4598 269
rect -4564 235 -4558 269
rect -4604 197 -4558 235
rect -4604 163 -4598 197
rect -4564 163 -4558 197
rect -4604 125 -4558 163
rect -4604 91 -4598 125
rect -4564 91 -4558 125
rect -4604 53 -4558 91
rect -4604 19 -4598 53
rect -4564 19 -4558 53
rect -4604 -19 -4558 19
rect -4604 -53 -4598 -19
rect -4564 -53 -4558 -19
rect -4604 -91 -4558 -53
rect -4604 -125 -4598 -91
rect -4564 -125 -4558 -91
rect -4604 -163 -4558 -125
rect -4604 -197 -4598 -163
rect -4564 -197 -4558 -163
rect -4604 -235 -4558 -197
rect -4604 -269 -4598 -235
rect -4564 -269 -4558 -235
rect -4604 -300 -4558 -269
rect -3586 269 -3540 300
rect -3586 235 -3580 269
rect -3546 235 -3540 269
rect -3586 197 -3540 235
rect -3586 163 -3580 197
rect -3546 163 -3540 197
rect -3586 125 -3540 163
rect -3586 91 -3580 125
rect -3546 91 -3540 125
rect -3586 53 -3540 91
rect -3586 19 -3580 53
rect -3546 19 -3540 53
rect -3586 -19 -3540 19
rect -3586 -53 -3580 -19
rect -3546 -53 -3540 -19
rect -3586 -91 -3540 -53
rect -3586 -125 -3580 -91
rect -3546 -125 -3540 -91
rect -3586 -163 -3540 -125
rect -3586 -197 -3580 -163
rect -3546 -197 -3540 -163
rect -3586 -235 -3540 -197
rect -3586 -269 -3580 -235
rect -3546 -269 -3540 -235
rect -3586 -300 -3540 -269
rect -2568 269 -2522 300
rect -2568 235 -2562 269
rect -2528 235 -2522 269
rect -2568 197 -2522 235
rect -2568 163 -2562 197
rect -2528 163 -2522 197
rect -2568 125 -2522 163
rect -2568 91 -2562 125
rect -2528 91 -2522 125
rect -2568 53 -2522 91
rect -2568 19 -2562 53
rect -2528 19 -2522 53
rect -2568 -19 -2522 19
rect -2568 -53 -2562 -19
rect -2528 -53 -2522 -19
rect -2568 -91 -2522 -53
rect -2568 -125 -2562 -91
rect -2528 -125 -2522 -91
rect -2568 -163 -2522 -125
rect -2568 -197 -2562 -163
rect -2528 -197 -2522 -163
rect -2568 -235 -2522 -197
rect -2568 -269 -2562 -235
rect -2528 -269 -2522 -235
rect -2568 -300 -2522 -269
rect -1550 269 -1504 300
rect -1550 235 -1544 269
rect -1510 235 -1504 269
rect -1550 197 -1504 235
rect -1550 163 -1544 197
rect -1510 163 -1504 197
rect -1550 125 -1504 163
rect -1550 91 -1544 125
rect -1510 91 -1504 125
rect -1550 53 -1504 91
rect -1550 19 -1544 53
rect -1510 19 -1504 53
rect -1550 -19 -1504 19
rect -1550 -53 -1544 -19
rect -1510 -53 -1504 -19
rect -1550 -91 -1504 -53
rect -1550 -125 -1544 -91
rect -1510 -125 -1504 -91
rect -1550 -163 -1504 -125
rect -1550 -197 -1544 -163
rect -1510 -197 -1504 -163
rect -1550 -235 -1504 -197
rect -1550 -269 -1544 -235
rect -1510 -269 -1504 -235
rect -1550 -300 -1504 -269
rect -532 269 -486 300
rect -532 235 -526 269
rect -492 235 -486 269
rect -532 197 -486 235
rect -532 163 -526 197
rect -492 163 -486 197
rect -532 125 -486 163
rect -532 91 -526 125
rect -492 91 -486 125
rect -532 53 -486 91
rect -532 19 -526 53
rect -492 19 -486 53
rect -532 -19 -486 19
rect -532 -53 -526 -19
rect -492 -53 -486 -19
rect -532 -91 -486 -53
rect -532 -125 -526 -91
rect -492 -125 -486 -91
rect -532 -163 -486 -125
rect -532 -197 -526 -163
rect -492 -197 -486 -163
rect -532 -235 -486 -197
rect -532 -269 -526 -235
rect -492 -269 -486 -235
rect -532 -300 -486 -269
rect 486 269 532 300
rect 486 235 492 269
rect 526 235 532 269
rect 486 197 532 235
rect 486 163 492 197
rect 526 163 532 197
rect 486 125 532 163
rect 486 91 492 125
rect 526 91 532 125
rect 486 53 532 91
rect 486 19 492 53
rect 526 19 532 53
rect 486 -19 532 19
rect 486 -53 492 -19
rect 526 -53 532 -19
rect 486 -91 532 -53
rect 486 -125 492 -91
rect 526 -125 532 -91
rect 486 -163 532 -125
rect 486 -197 492 -163
rect 526 -197 532 -163
rect 486 -235 532 -197
rect 486 -269 492 -235
rect 526 -269 532 -235
rect 486 -300 532 -269
rect 1504 269 1550 300
rect 1504 235 1510 269
rect 1544 235 1550 269
rect 1504 197 1550 235
rect 1504 163 1510 197
rect 1544 163 1550 197
rect 1504 125 1550 163
rect 1504 91 1510 125
rect 1544 91 1550 125
rect 1504 53 1550 91
rect 1504 19 1510 53
rect 1544 19 1550 53
rect 1504 -19 1550 19
rect 1504 -53 1510 -19
rect 1544 -53 1550 -19
rect 1504 -91 1550 -53
rect 1504 -125 1510 -91
rect 1544 -125 1550 -91
rect 1504 -163 1550 -125
rect 1504 -197 1510 -163
rect 1544 -197 1550 -163
rect 1504 -235 1550 -197
rect 1504 -269 1510 -235
rect 1544 -269 1550 -235
rect 1504 -300 1550 -269
rect 2522 269 2568 300
rect 2522 235 2528 269
rect 2562 235 2568 269
rect 2522 197 2568 235
rect 2522 163 2528 197
rect 2562 163 2568 197
rect 2522 125 2568 163
rect 2522 91 2528 125
rect 2562 91 2568 125
rect 2522 53 2568 91
rect 2522 19 2528 53
rect 2562 19 2568 53
rect 2522 -19 2568 19
rect 2522 -53 2528 -19
rect 2562 -53 2568 -19
rect 2522 -91 2568 -53
rect 2522 -125 2528 -91
rect 2562 -125 2568 -91
rect 2522 -163 2568 -125
rect 2522 -197 2528 -163
rect 2562 -197 2568 -163
rect 2522 -235 2568 -197
rect 2522 -269 2528 -235
rect 2562 -269 2568 -235
rect 2522 -300 2568 -269
rect 3540 269 3586 300
rect 3540 235 3546 269
rect 3580 235 3586 269
rect 3540 197 3586 235
rect 3540 163 3546 197
rect 3580 163 3586 197
rect 3540 125 3586 163
rect 3540 91 3546 125
rect 3580 91 3586 125
rect 3540 53 3586 91
rect 3540 19 3546 53
rect 3580 19 3586 53
rect 3540 -19 3586 19
rect 3540 -53 3546 -19
rect 3580 -53 3586 -19
rect 3540 -91 3586 -53
rect 3540 -125 3546 -91
rect 3580 -125 3586 -91
rect 3540 -163 3586 -125
rect 3540 -197 3546 -163
rect 3580 -197 3586 -163
rect 3540 -235 3586 -197
rect 3540 -269 3546 -235
rect 3580 -269 3586 -235
rect 3540 -300 3586 -269
rect 4558 269 4604 300
rect 4558 235 4564 269
rect 4598 235 4604 269
rect 4558 197 4604 235
rect 4558 163 4564 197
rect 4598 163 4604 197
rect 4558 125 4604 163
rect 4558 91 4564 125
rect 4598 91 4604 125
rect 4558 53 4604 91
rect 4558 19 4564 53
rect 4598 19 4604 53
rect 4558 -19 4604 19
rect 4558 -53 4564 -19
rect 4598 -53 4604 -19
rect 4558 -91 4604 -53
rect 4558 -125 4564 -91
rect 4598 -125 4604 -91
rect 4558 -163 4604 -125
rect 4558 -197 4564 -163
rect 4598 -197 4604 -163
rect 4558 -235 4604 -197
rect 4558 -269 4564 -235
rect 4598 -269 4604 -235
rect 4558 -300 4604 -269
rect 5576 269 5622 300
rect 5576 235 5582 269
rect 5616 235 5622 269
rect 5576 197 5622 235
rect 5576 163 5582 197
rect 5616 163 5622 197
rect 5576 125 5622 163
rect 5576 91 5582 125
rect 5616 91 5622 125
rect 5576 53 5622 91
rect 5576 19 5582 53
rect 5616 19 5622 53
rect 5576 -19 5622 19
rect 5576 -53 5582 -19
rect 5616 -53 5622 -19
rect 5576 -91 5622 -53
rect 5576 -125 5582 -91
rect 5616 -125 5622 -91
rect 5576 -163 5622 -125
rect 5576 -197 5582 -163
rect 5616 -197 5622 -163
rect 5576 -235 5622 -197
rect 5576 -269 5582 -235
rect 5616 -269 5622 -235
rect 5576 -300 5622 -269
rect -5334 -338 -4846 -332
rect -5334 -372 -5287 -338
rect -5253 -372 -5215 -338
rect -5181 -372 -5143 -338
rect -5109 -372 -5071 -338
rect -5037 -372 -4999 -338
rect -4965 -372 -4927 -338
rect -4893 -372 -4846 -338
rect -5334 -378 -4846 -372
rect -4316 -338 -3828 -332
rect -4316 -372 -4269 -338
rect -4235 -372 -4197 -338
rect -4163 -372 -4125 -338
rect -4091 -372 -4053 -338
rect -4019 -372 -3981 -338
rect -3947 -372 -3909 -338
rect -3875 -372 -3828 -338
rect -4316 -378 -3828 -372
rect -3298 -338 -2810 -332
rect -3298 -372 -3251 -338
rect -3217 -372 -3179 -338
rect -3145 -372 -3107 -338
rect -3073 -372 -3035 -338
rect -3001 -372 -2963 -338
rect -2929 -372 -2891 -338
rect -2857 -372 -2810 -338
rect -3298 -378 -2810 -372
rect -2280 -338 -1792 -332
rect -2280 -372 -2233 -338
rect -2199 -372 -2161 -338
rect -2127 -372 -2089 -338
rect -2055 -372 -2017 -338
rect -1983 -372 -1945 -338
rect -1911 -372 -1873 -338
rect -1839 -372 -1792 -338
rect -2280 -378 -1792 -372
rect -1262 -338 -774 -332
rect -1262 -372 -1215 -338
rect -1181 -372 -1143 -338
rect -1109 -372 -1071 -338
rect -1037 -372 -999 -338
rect -965 -372 -927 -338
rect -893 -372 -855 -338
rect -821 -372 -774 -338
rect -1262 -378 -774 -372
rect -244 -338 244 -332
rect -244 -372 -197 -338
rect -163 -372 -125 -338
rect -91 -372 -53 -338
rect -19 -372 19 -338
rect 53 -372 91 -338
rect 125 -372 163 -338
rect 197 -372 244 -338
rect -244 -378 244 -372
rect 774 -338 1262 -332
rect 774 -372 821 -338
rect 855 -372 893 -338
rect 927 -372 965 -338
rect 999 -372 1037 -338
rect 1071 -372 1109 -338
rect 1143 -372 1181 -338
rect 1215 -372 1262 -338
rect 774 -378 1262 -372
rect 1792 -338 2280 -332
rect 1792 -372 1839 -338
rect 1873 -372 1911 -338
rect 1945 -372 1983 -338
rect 2017 -372 2055 -338
rect 2089 -372 2127 -338
rect 2161 -372 2199 -338
rect 2233 -372 2280 -338
rect 1792 -378 2280 -372
rect 2810 -338 3298 -332
rect 2810 -372 2857 -338
rect 2891 -372 2929 -338
rect 2963 -372 3001 -338
rect 3035 -372 3073 -338
rect 3107 -372 3145 -338
rect 3179 -372 3217 -338
rect 3251 -372 3298 -338
rect 2810 -378 3298 -372
rect 3828 -338 4316 -332
rect 3828 -372 3875 -338
rect 3909 -372 3947 -338
rect 3981 -372 4019 -338
rect 4053 -372 4091 -338
rect 4125 -372 4163 -338
rect 4197 -372 4235 -338
rect 4269 -372 4316 -338
rect 3828 -378 4316 -372
rect 4846 -338 5334 -332
rect 4846 -372 4893 -338
rect 4927 -372 4965 -338
rect 4999 -372 5037 -338
rect 5071 -372 5109 -338
rect 5143 -372 5181 -338
rect 5215 -372 5253 -338
rect 5287 -372 5334 -338
rect 4846 -378 5334 -372
<< end >>
