magic
tech sky130A
magscale 1 2
timestamp 1622263318
<< nwell >>
rect 402 846 2798 3698
rect 10 522 2798 846
<< pwell >>
rect 92 358 278 465
rect 90 279 2798 358
rect 79 245 2798 279
rect 90 214 2798 245
rect 402 -1758 2798 214
<< nmos >>
rect 826 -630 1026 -230
rect 1084 -630 1284 -230
rect 1342 -630 1542 -230
rect 1600 -630 1800 -230
rect 1858 -630 2058 -230
rect 2116 -630 2316 -230
<< scnmos >>
rect 170 309 200 439
<< scpmoshvt >>
rect 170 559 200 759
<< pmoshvt >>
rect 831 2063 1031 2463
rect 1089 2063 1289 2463
rect 1347 2063 1547 2463
rect 1605 2063 1805 2463
rect 1863 2063 2063 2463
rect 2121 2063 2321 2463
rect 831 1203 1031 1603
rect 1089 1203 1289 1603
rect 1347 1203 1547 1603
rect 1605 1203 1805 1603
rect 1863 1203 2063 1603
rect 2121 1203 2321 1603
<< ndiff >>
rect 118 427 170 439
rect 118 393 126 427
rect 160 393 170 427
rect 118 359 170 393
rect 118 325 126 359
rect 160 325 170 359
rect 118 309 170 325
rect 200 427 252 439
rect 200 393 210 427
rect 244 393 252 427
rect 200 359 252 393
rect 200 325 210 359
rect 244 325 252 359
rect 200 309 252 325
rect 768 -242 826 -230
rect 768 -618 780 -242
rect 814 -618 826 -242
rect 768 -630 826 -618
rect 1026 -242 1084 -230
rect 1026 -618 1038 -242
rect 1072 -618 1084 -242
rect 1026 -630 1084 -618
rect 1284 -242 1342 -230
rect 1284 -618 1296 -242
rect 1330 -618 1342 -242
rect 1284 -630 1342 -618
rect 1542 -242 1600 -230
rect 1542 -618 1554 -242
rect 1588 -618 1600 -242
rect 1542 -630 1600 -618
rect 1800 -242 1858 -230
rect 1800 -618 1812 -242
rect 1846 -618 1858 -242
rect 1800 -630 1858 -618
rect 2058 -242 2116 -230
rect 2058 -618 2070 -242
rect 2104 -618 2116 -242
rect 2058 -630 2116 -618
rect 2316 -242 2374 -230
rect 2316 -618 2328 -242
rect 2362 -618 2374 -242
rect 2316 -630 2374 -618
<< pdiff >>
rect 118 747 170 759
rect 118 713 126 747
rect 160 713 170 747
rect 118 679 170 713
rect 118 645 126 679
rect 160 645 170 679
rect 118 611 170 645
rect 118 577 126 611
rect 160 577 170 611
rect 118 559 170 577
rect 200 747 252 759
rect 200 713 210 747
rect 244 713 252 747
rect 200 679 252 713
rect 200 645 210 679
rect 244 645 252 679
rect 200 611 252 645
rect 200 577 210 611
rect 244 577 252 611
rect 200 559 252 577
rect 773 2451 831 2463
rect 773 2075 785 2451
rect 819 2075 831 2451
rect 773 2063 831 2075
rect 1031 2451 1089 2463
rect 1031 2075 1043 2451
rect 1077 2075 1089 2451
rect 1031 2063 1089 2075
rect 1289 2451 1347 2463
rect 1289 2075 1301 2451
rect 1335 2075 1347 2451
rect 1289 2063 1347 2075
rect 1547 2451 1605 2463
rect 1547 2075 1559 2451
rect 1593 2075 1605 2451
rect 1547 2063 1605 2075
rect 1805 2451 1863 2463
rect 1805 2075 1817 2451
rect 1851 2075 1863 2451
rect 1805 2063 1863 2075
rect 2063 2451 2121 2463
rect 2063 2075 2075 2451
rect 2109 2075 2121 2451
rect 2063 2063 2121 2075
rect 2321 2451 2379 2463
rect 2321 2075 2333 2451
rect 2367 2075 2379 2451
rect 2321 2063 2379 2075
rect 773 1591 831 1603
rect 773 1215 785 1591
rect 819 1215 831 1591
rect 773 1203 831 1215
rect 1031 1591 1089 1603
rect 1031 1215 1043 1591
rect 1077 1215 1089 1591
rect 1031 1203 1089 1215
rect 1289 1591 1347 1603
rect 1289 1215 1301 1591
rect 1335 1215 1347 1591
rect 1289 1203 1347 1215
rect 1547 1591 1605 1603
rect 1547 1215 1559 1591
rect 1593 1215 1605 1591
rect 1547 1203 1605 1215
rect 1805 1591 1863 1603
rect 1805 1215 1817 1591
rect 1851 1215 1863 1591
rect 1805 1203 1863 1215
rect 2063 1591 2121 1603
rect 2063 1215 2075 1591
rect 2109 1215 2121 1591
rect 2063 1203 2121 1215
rect 2321 1591 2379 1603
rect 2321 1215 2333 1591
rect 2367 1215 2379 1591
rect 2321 1203 2379 1215
<< ndiffc >>
rect 126 393 160 427
rect 126 325 160 359
rect 210 393 244 427
rect 210 325 244 359
rect 780 -618 814 -242
rect 1038 -618 1072 -242
rect 1296 -618 1330 -242
rect 1554 -618 1588 -242
rect 1812 -618 1846 -242
rect 2070 -618 2104 -242
rect 2328 -618 2362 -242
<< pdiffc >>
rect 126 713 160 747
rect 126 645 160 679
rect 126 577 160 611
rect 210 713 244 747
rect 210 645 244 679
rect 210 577 244 611
rect 785 2075 819 2451
rect 1043 2075 1077 2451
rect 1301 2075 1335 2451
rect 1559 2075 1593 2451
rect 1817 2075 1851 2451
rect 2075 2075 2109 2451
rect 2333 2075 2367 2451
rect 785 1215 819 1591
rect 1043 1215 1077 1591
rect 1301 1215 1335 1591
rect 1559 1215 1593 1591
rect 1817 1215 1851 1591
rect 2075 1215 2109 1591
rect 2333 1215 2367 1591
<< psubdiff >>
rect 438 222 600 322
rect 2600 222 2762 322
rect 438 160 538 222
rect 2662 160 2762 222
rect 438 -1622 538 -1560
rect 2662 -1622 2762 -1560
rect 438 -1722 600 -1622
rect 2600 -1722 2762 -1622
<< nsubdiff >>
rect 438 3562 600 3662
rect 2600 3562 2762 3662
rect 438 3500 538 3562
rect 2662 3500 2762 3562
rect 438 658 538 720
rect 2662 658 2762 720
rect 438 558 600 658
rect 2600 558 2762 658
<< psubdiffcont >>
rect 600 222 2600 322
rect 438 -1560 538 160
rect 2662 -1560 2762 160
rect 600 -1722 2600 -1622
<< nsubdiffcont >>
rect 600 3562 2600 3662
rect 438 720 538 3500
rect 2662 720 2762 3500
rect 600 558 2600 658
<< poly >>
rect 170 759 200 785
rect 865 2544 997 2560
rect 865 2527 881 2544
rect 831 2510 881 2527
rect 981 2527 997 2544
rect 1123 2544 1255 2560
rect 1123 2527 1139 2544
rect 981 2510 1031 2527
rect 831 2463 1031 2510
rect 1089 2510 1139 2527
rect 1239 2527 1255 2544
rect 1381 2544 1513 2560
rect 1381 2527 1397 2544
rect 1239 2510 1289 2527
rect 1089 2463 1289 2510
rect 1347 2510 1397 2527
rect 1497 2527 1513 2544
rect 1639 2544 1771 2560
rect 1639 2527 1655 2544
rect 1497 2510 1547 2527
rect 1347 2463 1547 2510
rect 1605 2510 1655 2527
rect 1755 2527 1771 2544
rect 1897 2544 2029 2560
rect 1897 2527 1913 2544
rect 1755 2510 1805 2527
rect 1605 2463 1805 2510
rect 1863 2510 1913 2527
rect 2013 2527 2029 2544
rect 2155 2544 2287 2560
rect 2155 2527 2171 2544
rect 2013 2510 2063 2527
rect 1863 2463 2063 2510
rect 2121 2510 2171 2527
rect 2271 2527 2287 2544
rect 2271 2510 2321 2527
rect 2121 2463 2321 2510
rect 831 2016 1031 2063
rect 831 1999 881 2016
rect 865 1982 881 1999
rect 981 1999 1031 2016
rect 1089 2016 1289 2063
rect 1089 1999 1139 2016
rect 981 1982 997 1999
rect 865 1966 997 1982
rect 1123 1982 1139 1999
rect 1239 1999 1289 2016
rect 1347 2016 1547 2063
rect 1347 1999 1397 2016
rect 1239 1982 1255 1999
rect 1123 1966 1255 1982
rect 1381 1982 1397 1999
rect 1497 1999 1547 2016
rect 1605 2016 1805 2063
rect 1605 1999 1655 2016
rect 1497 1982 1513 1999
rect 1381 1966 1513 1982
rect 1639 1982 1655 1999
rect 1755 1999 1805 2016
rect 1863 2016 2063 2063
rect 1863 1999 1913 2016
rect 1755 1982 1771 1999
rect 1639 1966 1771 1982
rect 1897 1982 1913 1999
rect 2013 1999 2063 2016
rect 2121 2016 2321 2063
rect 2121 1999 2171 2016
rect 2013 1982 2029 1999
rect 1897 1966 2029 1982
rect 2155 1982 2171 1999
rect 2271 1999 2321 2016
rect 2271 1982 2287 1999
rect 2155 1966 2287 1982
rect 865 1684 997 1700
rect 865 1667 881 1684
rect 831 1650 881 1667
rect 981 1667 997 1684
rect 1123 1684 1255 1700
rect 1123 1667 1139 1684
rect 981 1650 1031 1667
rect 831 1603 1031 1650
rect 1089 1650 1139 1667
rect 1239 1667 1255 1684
rect 1381 1684 1513 1700
rect 1381 1667 1397 1684
rect 1239 1650 1289 1667
rect 1089 1603 1289 1650
rect 1347 1650 1397 1667
rect 1497 1667 1513 1684
rect 1639 1684 1771 1700
rect 1639 1667 1655 1684
rect 1497 1650 1547 1667
rect 1347 1603 1547 1650
rect 1605 1650 1655 1667
rect 1755 1667 1771 1684
rect 1897 1684 2029 1700
rect 1897 1667 1913 1684
rect 1755 1650 1805 1667
rect 1605 1603 1805 1650
rect 1863 1650 1913 1667
rect 2013 1667 2029 1684
rect 2155 1684 2287 1700
rect 2155 1667 2171 1684
rect 2013 1650 2063 1667
rect 1863 1603 2063 1650
rect 2121 1650 2171 1667
rect 2271 1667 2287 1684
rect 2271 1650 2321 1667
rect 2121 1603 2321 1650
rect 831 1156 1031 1203
rect 831 1139 881 1156
rect 865 1122 881 1139
rect 981 1139 1031 1156
rect 1089 1156 1289 1203
rect 1089 1139 1139 1156
rect 981 1122 997 1139
rect 865 1106 997 1122
rect 1123 1122 1139 1139
rect 1239 1139 1289 1156
rect 1347 1156 1547 1203
rect 1347 1139 1397 1156
rect 1239 1122 1255 1139
rect 1123 1106 1255 1122
rect 1381 1122 1397 1139
rect 1497 1139 1547 1156
rect 1605 1156 1805 1203
rect 1605 1139 1655 1156
rect 1497 1122 1513 1139
rect 1381 1106 1513 1122
rect 1639 1122 1655 1139
rect 1755 1139 1805 1156
rect 1863 1156 2063 1203
rect 1863 1139 1913 1156
rect 1755 1122 1771 1139
rect 1639 1106 1771 1122
rect 1897 1122 1913 1139
rect 2013 1139 2063 1156
rect 2121 1156 2321 1203
rect 2121 1139 2171 1156
rect 2013 1122 2029 1139
rect 1897 1106 2029 1122
rect 2155 1122 2171 1139
rect 2271 1139 2321 1156
rect 2271 1122 2287 1139
rect 2155 1106 2287 1122
rect 170 527 200 559
rect 114 511 200 527
rect 114 477 130 511
rect 164 477 200 511
rect 114 461 200 477
rect 170 439 200 461
rect 170 283 200 309
rect 860 -158 992 -142
rect 860 -175 876 -158
rect 826 -192 876 -175
rect 976 -175 992 -158
rect 1118 -158 1250 -142
rect 1118 -175 1134 -158
rect 976 -192 1026 -175
rect 826 -230 1026 -192
rect 1084 -192 1134 -175
rect 1234 -175 1250 -158
rect 1376 -158 1508 -142
rect 1376 -175 1392 -158
rect 1234 -192 1284 -175
rect 1084 -230 1284 -192
rect 1342 -192 1392 -175
rect 1492 -175 1508 -158
rect 1634 -158 1766 -142
rect 1634 -175 1650 -158
rect 1492 -192 1542 -175
rect 1342 -230 1542 -192
rect 1600 -192 1650 -175
rect 1750 -175 1766 -158
rect 1892 -158 2024 -142
rect 1892 -175 1908 -158
rect 1750 -192 1800 -175
rect 1600 -230 1800 -192
rect 1858 -192 1908 -175
rect 2008 -175 2024 -158
rect 2150 -158 2282 -142
rect 2150 -175 2166 -158
rect 2008 -192 2058 -175
rect 1858 -230 2058 -192
rect 2116 -192 2166 -175
rect 2266 -175 2282 -158
rect 2266 -192 2316 -175
rect 2116 -230 2316 -192
rect 826 -668 1026 -630
rect 826 -685 876 -668
rect 860 -702 876 -685
rect 976 -685 1026 -668
rect 1084 -668 1284 -630
rect 1084 -685 1134 -668
rect 976 -702 992 -685
rect 860 -718 992 -702
rect 1118 -702 1134 -685
rect 1234 -685 1284 -668
rect 1342 -668 1542 -630
rect 1342 -685 1392 -668
rect 1234 -702 1250 -685
rect 1118 -718 1250 -702
rect 1376 -702 1392 -685
rect 1492 -685 1542 -668
rect 1600 -668 1800 -630
rect 1600 -685 1650 -668
rect 1492 -702 1508 -685
rect 1376 -718 1508 -702
rect 1634 -702 1650 -685
rect 1750 -685 1800 -668
rect 1858 -668 2058 -630
rect 1858 -685 1908 -668
rect 1750 -702 1766 -685
rect 1634 -718 1766 -702
rect 1892 -702 1908 -685
rect 2008 -685 2058 -668
rect 2116 -668 2316 -630
rect 2116 -685 2166 -668
rect 2008 -702 2024 -685
rect 1892 -718 2024 -702
rect 2150 -702 2166 -685
rect 2266 -685 2316 -668
rect 2266 -702 2282 -685
rect 2150 -718 2282 -702
<< polycont >>
rect 881 2510 981 2544
rect 1139 2510 1239 2544
rect 1397 2510 1497 2544
rect 1655 2510 1755 2544
rect 1913 2510 2013 2544
rect 2171 2510 2271 2544
rect 881 1982 981 2016
rect 1139 1982 1239 2016
rect 1397 1982 1497 2016
rect 1655 1982 1755 2016
rect 1913 1982 2013 2016
rect 2171 1982 2271 2016
rect 881 1650 981 1684
rect 1139 1650 1239 1684
rect 1397 1650 1497 1684
rect 1655 1650 1755 1684
rect 1913 1650 2013 1684
rect 2171 1650 2271 1684
rect 881 1122 981 1156
rect 1139 1122 1239 1156
rect 1397 1122 1497 1156
rect 1655 1122 1755 1156
rect 1913 1122 2013 1156
rect 2171 1122 2271 1156
rect 130 477 164 511
rect 876 -192 976 -158
rect 1134 -192 1234 -158
rect 1392 -192 1492 -158
rect 1650 -192 1750 -158
rect 1908 -192 2008 -158
rect 2166 -192 2266 -158
rect 876 -702 976 -668
rect 1134 -702 1234 -668
rect 1392 -702 1492 -668
rect 1650 -702 1750 -668
rect 1908 -702 2008 -668
rect 2166 -702 2266 -668
<< locali >>
rect 438 3500 538 3662
rect 50 789 79 823
rect 113 789 171 823
rect 205 789 263 823
rect 297 789 326 823
rect 2662 3500 2762 3662
rect 865 2510 881 2544
rect 981 2510 997 2544
rect 1123 2510 1139 2544
rect 1239 2510 1255 2544
rect 1381 2510 1397 2544
rect 1497 2510 1513 2544
rect 1639 2510 1655 2544
rect 1755 2510 1771 2544
rect 1897 2510 1913 2544
rect 2013 2510 2029 2544
rect 2155 2510 2171 2544
rect 2271 2510 2287 2544
rect 785 2451 819 2467
rect 785 2059 819 2075
rect 1043 2451 1077 2467
rect 1043 2059 1077 2075
rect 1301 2451 1335 2467
rect 1301 2059 1335 2075
rect 1559 2451 1593 2467
rect 1559 2059 1593 2075
rect 1817 2451 1851 2467
rect 1817 2059 1851 2075
rect 2075 2451 2109 2467
rect 2075 2059 2109 2075
rect 2333 2451 2367 2467
rect 2333 2059 2367 2075
rect 865 1982 881 2016
rect 981 1982 997 2016
rect 1123 1982 1139 2016
rect 1239 1982 1255 2016
rect 1381 1982 1397 2016
rect 1497 1982 1513 2016
rect 1639 1982 1655 2016
rect 1755 1982 1771 2016
rect 1897 1982 1913 2016
rect 2013 1982 2029 2016
rect 2155 1982 2171 2016
rect 2271 1982 2287 2016
rect 865 1650 881 1684
rect 981 1650 997 1684
rect 1123 1650 1139 1684
rect 1239 1650 1255 1684
rect 1381 1650 1397 1684
rect 1497 1650 1513 1684
rect 1639 1650 1655 1684
rect 1755 1650 1771 1684
rect 1897 1650 1913 1684
rect 2013 1650 2029 1684
rect 2155 1650 2171 1684
rect 2271 1650 2287 1684
rect 785 1591 819 1607
rect 785 1199 819 1215
rect 1043 1591 1077 1607
rect 1043 1199 1077 1215
rect 1301 1591 1335 1607
rect 1301 1199 1335 1215
rect 1559 1591 1593 1607
rect 1559 1199 1593 1215
rect 1817 1591 1851 1607
rect 1817 1199 1851 1215
rect 2075 1591 2109 1607
rect 2075 1199 2109 1215
rect 2333 1591 2367 1607
rect 2333 1199 2367 1215
rect 865 1122 881 1156
rect 981 1122 997 1156
rect 1123 1122 1139 1156
rect 1239 1122 1255 1156
rect 1381 1122 1397 1156
rect 1497 1122 1513 1156
rect 1639 1122 1655 1156
rect 1755 1122 1771 1156
rect 1897 1122 1913 1156
rect 2013 1122 2029 1156
rect 2155 1122 2171 1156
rect 2271 1122 2287 1156
rect 118 747 160 789
rect 118 713 126 747
rect 118 679 160 713
rect 118 645 126 679
rect 118 611 160 645
rect 118 577 126 611
rect 118 561 160 577
rect 194 747 260 755
rect 194 713 210 747
rect 244 713 260 747
rect 194 679 260 713
rect 194 645 210 679
rect 244 645 260 679
rect 194 611 260 645
rect 194 577 210 611
rect 244 577 260 611
rect 194 559 260 577
rect 114 478 118 525
rect 166 478 180 525
rect 114 477 130 478
rect 164 477 180 478
rect 214 468 260 559
rect 438 558 538 720
rect 2662 558 2762 720
rect 114 427 160 443
rect 214 439 220 468
rect 114 393 126 427
rect 114 359 160 393
rect 114 325 126 359
rect 114 279 160 325
rect 194 427 220 439
rect 194 393 210 427
rect 244 393 260 420
rect 194 359 260 393
rect 194 325 210 359
rect 244 325 260 359
rect 194 313 260 325
rect 50 245 79 279
rect 113 245 171 279
rect 205 245 263 279
rect 297 245 326 279
rect 438 160 538 322
rect 2662 160 2762 322
rect 860 -192 876 -158
rect 976 -192 992 -158
rect 1118 -192 1134 -158
rect 1234 -192 1250 -158
rect 1376 -192 1392 -158
rect 1492 -192 1508 -158
rect 1634 -192 1650 -158
rect 1750 -192 1766 -158
rect 1892 -192 1908 -158
rect 2008 -192 2024 -158
rect 2150 -192 2166 -158
rect 2266 -192 2282 -158
rect 780 -242 814 -226
rect 780 -634 814 -618
rect 1038 -242 1072 -226
rect 1038 -634 1072 -618
rect 1296 -242 1330 -226
rect 1296 -634 1330 -618
rect 1554 -242 1588 -226
rect 1554 -634 1588 -618
rect 1812 -242 1846 -226
rect 1812 -634 1846 -618
rect 2070 -242 2104 -226
rect 2070 -634 2104 -618
rect 2328 -242 2362 -226
rect 2328 -634 2362 -618
rect 860 -702 876 -668
rect 976 -702 992 -668
rect 1118 -702 1134 -668
rect 1234 -702 1250 -668
rect 1376 -702 1392 -668
rect 1492 -702 1508 -668
rect 1634 -702 1650 -668
rect 1750 -702 1766 -668
rect 1892 -702 1908 -668
rect 2008 -702 2024 -668
rect 2150 -702 2166 -668
rect 2266 -702 2282 -668
rect 438 -1722 538 -1560
rect 2662 -1722 2762 -1560
<< viali >>
rect 538 3562 600 3662
rect 600 3562 2600 3662
rect 2600 3562 2662 3662
rect 79 789 113 823
rect 171 789 205 823
rect 263 789 297 823
rect 438 798 538 3422
rect 889 2510 973 2544
rect 1147 2510 1231 2544
rect 1405 2510 1489 2544
rect 1663 2510 1747 2544
rect 1921 2510 2005 2544
rect 2179 2510 2263 2544
rect 785 2075 819 2451
rect 1043 2075 1077 2451
rect 1301 2075 1335 2451
rect 1559 2075 1593 2451
rect 1817 2075 1851 2451
rect 2075 2075 2109 2451
rect 2333 2075 2367 2451
rect 889 1982 973 2016
rect 1147 1982 1231 2016
rect 1405 1982 1489 2016
rect 1663 1982 1747 2016
rect 1921 1982 2005 2016
rect 2179 1982 2263 2016
rect 889 1650 973 1684
rect 1147 1650 1231 1684
rect 1405 1650 1489 1684
rect 1663 1650 1747 1684
rect 1921 1650 2005 1684
rect 2179 1650 2263 1684
rect 785 1215 819 1591
rect 1043 1215 1077 1591
rect 1301 1215 1335 1591
rect 1559 1215 1593 1591
rect 1817 1215 1851 1591
rect 2075 1215 2109 1591
rect 2333 1215 2367 1591
rect 889 1122 973 1156
rect 1147 1122 1231 1156
rect 1405 1122 1489 1156
rect 1663 1122 1747 1156
rect 1921 1122 2005 1156
rect 2179 1122 2263 1156
rect 118 511 166 526
rect 118 478 130 511
rect 130 478 164 511
rect 164 478 166 511
rect 2662 798 2762 3422
rect 538 558 600 658
rect 600 558 2600 658
rect 2600 558 2662 658
rect 220 427 268 468
rect 220 420 244 427
rect 244 420 268 427
rect 79 245 113 279
rect 171 245 205 279
rect 263 245 297 279
rect 538 222 600 322
rect 600 222 2600 322
rect 2600 222 2662 322
rect 438 -1530 538 130
rect 884 -192 968 -158
rect 1142 -192 1226 -158
rect 1400 -192 1484 -158
rect 1658 -192 1742 -158
rect 1916 -192 2000 -158
rect 2174 -192 2258 -158
rect 780 -618 814 -242
rect 1038 -618 1072 -242
rect 1296 -618 1330 -242
rect 1554 -618 1588 -242
rect 1812 -618 1846 -242
rect 2070 -618 2104 -242
rect 2328 -618 2362 -242
rect 884 -702 968 -668
rect 1142 -702 1226 -668
rect 1400 -702 1484 -668
rect 1658 -702 1742 -668
rect 1916 -702 2000 -668
rect 2174 -702 2258 -668
rect 2662 -1530 2762 130
rect 538 -1722 600 -1622
rect 600 -1722 2600 -1622
rect 2600 -1722 2662 -1622
<< metal1 >>
rect 432 3662 2768 3668
rect 432 3562 538 3662
rect 2662 3562 2768 3662
rect 432 3556 2768 3562
rect 432 3422 544 3556
rect 432 854 438 3422
rect 50 823 438 854
rect 50 789 79 823
rect 113 789 171 823
rect 205 789 263 823
rect 297 798 438 823
rect 538 798 544 3422
rect 1144 3256 1154 3556
rect 2046 3256 2056 3556
rect 2656 3422 2768 3556
rect 700 3052 2602 3082
rect 700 2988 734 3052
rect 2558 2988 2602 3052
rect 700 2958 2602 2988
rect 774 2694 834 2958
rect 904 2694 964 2958
rect 1282 2814 1288 2874
rect 1348 2814 1354 2874
rect 1800 2814 1806 2874
rect 1866 2814 1872 2874
rect 620 2582 626 2642
rect 686 2582 692 2642
rect 774 2634 964 2694
rect 626 2048 686 2582
rect 774 2451 834 2634
rect 904 2550 964 2634
rect 877 2544 985 2550
rect 877 2510 889 2544
rect 973 2510 985 2544
rect 877 2504 985 2510
rect 1135 2544 1243 2550
rect 1135 2510 1147 2544
rect 1231 2510 1243 2544
rect 1135 2504 1243 2510
rect 774 2418 785 2451
rect 779 2118 785 2418
rect 626 1068 686 1988
rect 774 2075 785 2118
rect 819 2418 834 2451
rect 1037 2451 1083 2463
rect 819 2118 825 2418
rect 819 2075 834 2118
rect 1037 2100 1043 2451
rect 774 1852 834 2075
rect 1030 2075 1043 2100
rect 1077 2100 1083 2451
rect 1288 2451 1348 2814
rect 1538 2702 1544 2762
rect 1604 2702 1610 2762
rect 1410 2582 1416 2642
rect 1476 2582 1482 2642
rect 1416 2550 1476 2582
rect 1393 2544 1501 2550
rect 1393 2510 1405 2544
rect 1489 2510 1501 2544
rect 1393 2504 1501 2510
rect 1077 2075 1090 2100
rect 877 2016 985 2022
rect 877 1982 889 2016
rect 973 1982 985 2016
rect 877 1976 985 1982
rect 904 1852 964 1976
rect 774 1792 964 1852
rect 1030 1804 1090 2075
rect 1288 2075 1301 2451
rect 1335 2075 1348 2451
rect 1544 2451 1604 2702
rect 1666 2582 1672 2642
rect 1732 2582 1738 2642
rect 1672 2550 1732 2582
rect 1651 2544 1759 2550
rect 1651 2510 1663 2544
rect 1747 2510 1759 2544
rect 1651 2504 1759 2510
rect 1544 2418 1559 2451
rect 1135 2016 1243 2022
rect 1135 1982 1147 2016
rect 1231 1982 1243 2016
rect 1135 1976 1243 1982
rect 1160 1918 1220 1976
rect 1154 1858 1160 1918
rect 1220 1858 1226 1918
rect 774 1591 834 1792
rect 904 1690 964 1792
rect 1024 1744 1030 1804
rect 1090 1744 1096 1804
rect 877 1684 985 1690
rect 877 1650 889 1684
rect 973 1650 985 1684
rect 877 1644 985 1650
rect 1135 1684 1243 1690
rect 1135 1650 1147 1684
rect 1231 1650 1243 1684
rect 1135 1644 1243 1650
rect 774 1538 785 1591
rect 779 1215 785 1538
rect 819 1538 834 1591
rect 1037 1591 1083 1603
rect 819 1215 825 1538
rect 1037 1260 1043 1591
rect 779 1203 825 1215
rect 1028 1215 1043 1260
rect 1077 1260 1083 1591
rect 1288 1591 1348 2075
rect 1553 2075 1559 2418
rect 1593 2418 1604 2451
rect 1806 2451 1866 2814
rect 2194 2682 2254 2958
rect 2322 2682 2382 2958
rect 2468 2702 2474 2762
rect 2534 2702 2540 2762
rect 2194 2622 2382 2682
rect 2194 2550 2254 2622
rect 1909 2544 2017 2550
rect 1909 2510 1921 2544
rect 2005 2510 2017 2544
rect 1909 2504 2017 2510
rect 2167 2544 2275 2550
rect 2167 2510 2179 2544
rect 2263 2510 2275 2544
rect 2167 2504 2275 2510
rect 1593 2075 1599 2418
rect 1806 2390 1817 2451
rect 1811 2132 1817 2390
rect 1553 2063 1599 2075
rect 1800 2075 1817 2132
rect 1851 2390 1866 2451
rect 2069 2451 2115 2463
rect 1851 2132 1857 2390
rect 1851 2075 1860 2132
rect 2069 2124 2075 2451
rect 1393 2016 1501 2022
rect 1393 1982 1405 2016
rect 1489 1982 1501 2016
rect 1393 1976 1501 1982
rect 1651 2016 1759 2022
rect 1651 1982 1663 2016
rect 1747 1982 1759 2016
rect 1651 1976 1759 1982
rect 1412 1858 1418 1918
rect 1478 1858 1484 1918
rect 1670 1858 1676 1918
rect 1736 1858 1742 1918
rect 1418 1690 1478 1858
rect 1542 1744 1548 1804
rect 1608 1744 1614 1804
rect 1393 1684 1501 1690
rect 1393 1650 1405 1684
rect 1489 1650 1501 1684
rect 1393 1644 1501 1650
rect 1077 1215 1088 1260
rect 1288 1252 1301 1591
rect 877 1156 985 1162
rect 877 1122 889 1156
rect 973 1122 985 1156
rect 877 1116 985 1122
rect 626 1008 876 1068
rect 936 1008 942 1068
rect 1028 956 1088 1215
rect 1295 1215 1301 1252
rect 1335 1252 1348 1591
rect 1548 1591 1608 1744
rect 1676 1690 1736 1858
rect 1651 1684 1759 1690
rect 1651 1650 1663 1684
rect 1747 1650 1759 1684
rect 1651 1644 1759 1650
rect 1548 1558 1559 1591
rect 1553 1254 1559 1558
rect 1335 1215 1341 1252
rect 1295 1203 1341 1215
rect 1544 1215 1559 1254
rect 1593 1558 1608 1591
rect 1800 1591 1860 2075
rect 2064 2075 2075 2124
rect 2109 2124 2115 2451
rect 2322 2451 2382 2622
rect 2109 2075 2124 2124
rect 1909 2016 2017 2022
rect 1909 1982 1921 2016
rect 2005 1982 2017 2016
rect 1909 1976 2017 1982
rect 1934 1918 1994 1976
rect 1928 1858 1934 1918
rect 1994 1858 2000 1918
rect 2064 1804 2124 2075
rect 2322 2075 2333 2451
rect 2367 2075 2382 2451
rect 2167 2016 2275 2022
rect 2167 1982 2179 2016
rect 2263 1982 2275 2016
rect 2167 1976 2275 1982
rect 2322 1860 2382 2075
rect 2058 1744 2064 1804
rect 2124 1744 2130 1804
rect 2190 1800 2382 1860
rect 2190 1690 2250 1800
rect 1909 1684 2017 1690
rect 1909 1650 1921 1684
rect 2005 1650 2017 1684
rect 1909 1644 2017 1650
rect 2167 1684 2275 1690
rect 2167 1650 2179 1684
rect 2263 1650 2275 1684
rect 2167 1644 2275 1650
rect 1593 1254 1599 1558
rect 1800 1546 1817 1591
rect 1811 1268 1817 1546
rect 1593 1215 1604 1254
rect 1135 1156 1243 1162
rect 1135 1122 1147 1156
rect 1231 1122 1243 1156
rect 1135 1116 1243 1122
rect 1393 1156 1501 1162
rect 1393 1122 1405 1156
rect 1489 1122 1501 1156
rect 1393 1116 1501 1122
rect 1160 1068 1220 1116
rect 1154 1008 1160 1068
rect 1220 1008 1226 1068
rect 1022 896 1028 956
rect 1088 896 1094 956
rect 1544 808 1604 1215
rect 1802 1215 1817 1268
rect 1851 1546 1860 1591
rect 2069 1591 2115 1603
rect 1851 1268 1857 1546
rect 2069 1292 2075 1591
rect 1851 1215 1862 1268
rect 1651 1156 1759 1162
rect 1651 1122 1663 1156
rect 1747 1122 1759 1156
rect 1651 1116 1759 1122
rect 1672 1062 1732 1116
rect 1802 848 1862 1215
rect 2064 1215 2075 1292
rect 2109 1292 2115 1591
rect 2322 1591 2382 1800
rect 2109 1215 2124 1292
rect 1909 1156 2017 1162
rect 1909 1122 1921 1156
rect 2005 1122 2017 1156
rect 1909 1116 2017 1122
rect 1936 1068 1996 1116
rect 1930 1008 1936 1068
rect 1996 1008 2002 1068
rect 2064 956 2124 1215
rect 2322 1215 2333 1591
rect 2367 1215 2382 1591
rect 2167 1156 2275 1162
rect 2167 1122 2179 1156
rect 2263 1122 2275 1156
rect 2167 1116 2275 1122
rect 2188 1070 2248 1116
rect 2322 1070 2382 1215
rect 2188 1010 2382 1070
rect 2058 896 2064 956
rect 2124 896 2130 956
rect 297 789 544 798
rect 50 758 544 789
rect 432 664 544 758
rect 1538 748 1544 808
rect 1604 748 1610 808
rect 1796 788 1802 848
rect 1862 788 1868 848
rect 2188 664 2248 1010
rect 2322 664 2382 1010
rect 2474 956 2534 2702
rect 2468 896 2474 956
rect 2534 896 2540 956
rect 2656 798 2662 3422
rect 2762 798 2768 3422
rect 2656 664 2768 798
rect 432 658 2768 664
rect 432 558 538 658
rect 2662 558 2768 658
rect 432 552 2768 558
rect -108 532 -48 538
rect -48 526 178 532
rect -48 478 118 526
rect 166 478 178 526
rect -48 472 178 478
rect 214 474 274 480
rect -108 466 -48 472
rect 208 414 214 474
rect 274 414 280 474
rect 214 408 274 414
rect 432 322 2768 328
rect 432 310 538 322
rect 50 279 538 310
rect 50 245 79 279
rect 113 245 171 279
rect 205 245 263 279
rect 297 245 538 279
rect 50 222 538 245
rect 2662 222 2768 322
rect 50 216 2768 222
rect 50 214 544 216
rect 432 130 544 214
rect 432 -1530 438 130
rect 538 -1530 544 130
rect 1544 168 1604 174
rect 1022 42 1028 102
rect 1088 42 1094 102
rect 872 -158 980 -152
rect 872 -192 884 -158
rect 968 -192 980 -158
rect 872 -198 980 -192
rect 774 -242 820 -230
rect 774 -564 780 -242
rect 766 -618 780 -564
rect 814 -564 820 -242
rect 1028 -242 1088 42
rect 1276 -2 1282 58
rect 1342 -2 1348 58
rect 1130 -158 1238 -152
rect 1130 -192 1142 -158
rect 1226 -192 1238 -158
rect 1130 -198 1238 -192
rect 1028 -312 1038 -242
rect 814 -618 826 -564
rect 1032 -582 1038 -312
rect 766 -738 826 -618
rect 1022 -618 1038 -582
rect 1072 -312 1088 -242
rect 1282 -242 1342 -2
rect 1408 -114 1414 -54
rect 1474 -114 1480 -54
rect 1414 -152 1474 -114
rect 1388 -158 1496 -152
rect 1388 -192 1400 -158
rect 1484 -192 1496 -158
rect 1388 -198 1496 -192
rect 1282 -278 1296 -242
rect 1072 -582 1078 -312
rect 1072 -618 1082 -582
rect 872 -668 980 -662
rect 872 -702 884 -668
rect 968 -702 980 -668
rect 872 -708 980 -702
rect 896 -738 956 -708
rect 766 -798 956 -738
rect 766 -1034 826 -798
rect 896 -1034 956 -798
rect 1022 -864 1082 -618
rect 1290 -618 1296 -278
rect 1330 -278 1342 -242
rect 1544 -242 1604 108
rect 2656 130 2768 216
rect 1796 -2 1802 58
rect 1862 -2 1868 58
rect 1664 -114 1670 -54
rect 1730 -114 1736 -54
rect 1670 -152 1730 -114
rect 1646 -158 1754 -152
rect 1646 -192 1658 -158
rect 1742 -192 1754 -158
rect 1646 -198 1754 -192
rect 1544 -274 1554 -242
rect 1330 -618 1336 -278
rect 1290 -630 1336 -618
rect 1548 -618 1554 -274
rect 1588 -274 1604 -242
rect 1802 -242 1862 -2
rect 1904 -158 2012 -152
rect 1904 -192 1916 -158
rect 2000 -192 2012 -158
rect 1904 -198 2012 -192
rect 2162 -158 2270 -152
rect 2162 -192 2174 -158
rect 2258 -192 2270 -158
rect 2162 -198 2270 -192
rect 1588 -618 1594 -274
rect 1802 -284 1812 -242
rect 1548 -630 1594 -618
rect 1806 -618 1812 -284
rect 1846 -284 1862 -242
rect 2064 -242 2110 -230
rect 1846 -618 1852 -284
rect 2064 -564 2070 -242
rect 1806 -630 1852 -618
rect 2058 -618 2070 -564
rect 2104 -564 2110 -242
rect 2322 -242 2368 -230
rect 2104 -618 2118 -564
rect 2322 -572 2328 -242
rect 1130 -668 1238 -662
rect 1130 -702 1142 -668
rect 1226 -702 1238 -668
rect 1130 -708 1238 -702
rect 1388 -668 1496 -662
rect 1388 -702 1400 -668
rect 1484 -702 1496 -668
rect 1388 -708 1496 -702
rect 1646 -668 1754 -662
rect 1646 -702 1658 -668
rect 1742 -702 1754 -668
rect 1646 -708 1754 -702
rect 1904 -668 2012 -662
rect 1904 -702 1916 -668
rect 2000 -702 2012 -668
rect 1904 -708 2012 -702
rect 1156 -750 1216 -708
rect 1930 -750 1990 -708
rect 1150 -810 1156 -750
rect 1216 -810 1222 -750
rect 1924 -810 1930 -750
rect 1990 -810 1996 -750
rect 2058 -864 2118 -618
rect 2314 -618 2328 -572
rect 2362 -572 2368 -242
rect 2362 -618 2374 -572
rect 2162 -668 2270 -662
rect 2162 -702 2174 -668
rect 2258 -702 2270 -668
rect 2162 -708 2270 -702
rect 2186 -744 2246 -708
rect 2314 -744 2374 -618
rect 2186 -804 2374 -744
rect 1016 -924 1022 -864
rect 1082 -924 1088 -864
rect 2052 -924 2058 -864
rect 2118 -924 2124 -864
rect 2186 -1034 2246 -804
rect 2314 -1034 2374 -804
rect 656 -1066 2434 -1034
rect 656 -1134 692 -1066
rect 2400 -1134 2434 -1066
rect 656 -1164 2434 -1134
rect 432 -1616 544 -1530
rect 1144 -1616 1154 -1316
rect 2046 -1616 2056 -1316
rect 2656 -1530 2662 130
rect 2762 -1530 2768 130
rect 2656 -1616 2768 -1530
rect 432 -1622 2768 -1616
rect 432 -1722 538 -1622
rect 2662 -1722 2768 -1622
rect 432 -1728 2768 -1722
<< via1 >>
rect 544 3256 1144 3556
rect 2056 3256 2656 3556
rect 734 2988 2558 3052
rect 1288 2814 1348 2874
rect 1806 2814 1866 2874
rect 626 2582 686 2642
rect 626 1988 686 2048
rect 1544 2702 1604 2762
rect 1416 2582 1476 2642
rect 1672 2582 1732 2642
rect 1160 1858 1220 1918
rect 1030 1744 1090 1804
rect 2474 2702 2534 2762
rect 1418 1858 1478 1918
rect 1676 1858 1736 1918
rect 1548 1744 1608 1804
rect 876 1008 936 1068
rect 1934 1858 1994 1918
rect 2064 1744 2124 1804
rect 1160 1008 1220 1068
rect 1028 896 1088 956
rect 1936 1008 1996 1068
rect 2064 896 2124 956
rect 1544 748 1604 808
rect 1802 788 1862 848
rect 2474 896 2534 956
rect -108 472 -48 532
rect 214 468 274 474
rect 214 420 220 468
rect 220 420 268 468
rect 268 420 274 468
rect 214 414 274 420
rect 1544 108 1604 168
rect 1028 42 1088 102
rect 1282 -2 1342 58
rect 1414 -114 1474 -54
rect 1802 -2 1862 58
rect 1670 -114 1730 -54
rect 1156 -810 1216 -750
rect 1930 -810 1990 -750
rect 1022 -924 1082 -864
rect 2058 -924 2118 -864
rect 692 -1134 2400 -1066
rect 544 -1616 1144 -1316
rect 2056 -1616 2656 -1316
<< metal2 >>
rect 544 3556 1144 3566
rect 544 3246 1144 3256
rect 2056 3556 2656 3566
rect 2056 3246 2656 3256
rect 700 3052 2602 3082
rect 700 2988 734 3052
rect 2558 2988 2602 3052
rect 700 2958 2602 2988
rect 1288 2874 1348 2880
rect 1806 2874 1866 2880
rect 1348 2814 1806 2874
rect 1288 2808 1348 2814
rect 1806 2808 1866 2814
rect 1544 2762 1604 2768
rect 2474 2762 2534 2768
rect 1604 2702 2474 2762
rect 1544 2696 1604 2702
rect 2474 2696 2534 2702
rect 626 2642 686 2648
rect 1416 2642 1476 2648
rect 1672 2642 1732 2648
rect 686 2582 1416 2642
rect 1476 2582 1672 2642
rect 626 2576 686 2582
rect 1416 2576 1476 2582
rect 1672 2576 1732 2582
rect -108 1988 626 2048
rect 686 1988 692 2048
rect -108 532 -48 1988
rect 1160 1918 1220 1924
rect 1418 1918 1478 1924
rect 1676 1918 1736 1924
rect 1934 1918 1994 1924
rect 628 1858 1160 1918
rect 1220 1858 1418 1918
rect 1478 1858 1676 1918
rect 1736 1858 1934 1918
rect -114 472 -108 532
rect -48 472 -42 532
rect 628 474 688 1858
rect 1160 1852 1220 1858
rect 1418 1852 1478 1858
rect 1676 1852 1736 1858
rect 1934 1852 1994 1858
rect 1030 1804 1090 1810
rect 1548 1804 1608 1810
rect 2064 1804 2124 1810
rect 1090 1744 1548 1804
rect 1608 1744 2064 1804
rect 1030 1738 1090 1744
rect 1548 1738 1608 1744
rect 2064 1738 2124 1744
rect 208 414 214 474
rect 274 414 688 474
rect 628 -750 688 414
rect 876 1068 936 1074
rect 1160 1068 1220 1074
rect 1936 1068 1996 1074
rect 936 1008 1160 1068
rect 1220 1008 1936 1068
rect 876 -54 936 1008
rect 1160 1002 1220 1008
rect 1936 1002 1996 1008
rect 1028 956 1088 962
rect 2064 956 2124 962
rect 2474 956 2534 962
rect 1088 896 2064 956
rect 2124 896 2474 956
rect 1028 102 1088 896
rect 2064 890 2124 896
rect 2474 890 2534 896
rect 1802 848 1862 854
rect 1544 808 1604 814
rect 1544 168 1604 748
rect 1538 108 1544 168
rect 1604 108 1610 168
rect 1028 36 1088 42
rect 1282 58 1342 64
rect 1802 58 1862 788
rect 1342 -2 1802 58
rect 1282 -8 1342 -2
rect 1802 -8 1862 -2
rect 1414 -54 1474 -48
rect 1670 -54 1730 -48
rect 876 -114 1414 -54
rect 1474 -114 1670 -54
rect 1414 -120 1474 -114
rect 1670 -120 1730 -114
rect 1156 -750 1216 -744
rect 1930 -750 1990 -744
rect 628 -810 1156 -750
rect 1216 -810 1930 -750
rect 1156 -816 1216 -810
rect 1930 -816 1990 -810
rect 1022 -864 1082 -858
rect 2058 -864 2118 -858
rect 1082 -924 2058 -864
rect 1022 -930 1082 -924
rect 2058 -930 2118 -924
rect 656 -1066 2434 -1034
rect 656 -1134 692 -1066
rect 2400 -1134 2434 -1066
rect 656 -1164 2434 -1134
rect 544 -1316 1144 -1306
rect 544 -1626 1144 -1616
rect 2056 -1316 2656 -1306
rect 2056 -1626 2656 -1616
<< via2 >>
rect 544 3256 1144 3556
rect 2056 3256 2656 3556
rect 734 2988 2558 3052
rect 692 -1134 2400 -1066
rect 544 -1616 1144 -1316
rect 2056 -1616 2656 -1316
<< metal3 >>
rect 534 3556 1154 3561
rect 534 3256 544 3556
rect 1144 3256 1154 3556
rect 534 3251 1154 3256
rect 2046 3556 2666 3561
rect 2046 3256 2056 3556
rect 2656 3256 2666 3556
rect 2046 3251 2666 3256
rect 700 3052 2602 3082
rect 700 2988 734 3052
rect 2558 2988 2602 3052
rect 700 2958 2602 2988
rect 656 -1066 2434 -1034
rect 656 -1134 692 -1066
rect 2400 -1134 2434 -1066
rect 656 -1164 2434 -1134
rect 534 -1316 1154 -1311
rect 534 -1616 544 -1316
rect 1144 -1616 1154 -1316
rect 534 -1621 1154 -1616
rect 2046 -1316 2666 -1311
rect 2046 -1616 2056 -1316
rect 2656 -1616 2666 -1316
rect 2046 -1621 2666 -1616
<< via3 >>
rect 544 3256 1144 3556
rect 2056 3256 2656 3556
rect 734 2988 2558 3052
rect 692 -1134 2400 -1066
rect 544 -1616 1144 -1316
rect 2056 -1616 2656 -1316
<< metal4 >>
rect 360 3556 2840 3740
rect 360 3256 544 3556
rect 1144 3256 2056 3556
rect 2656 3256 2840 3556
rect 360 3052 2840 3256
rect 360 2988 734 3052
rect 2558 2988 2840 3052
rect 360 2940 2840 2988
rect 360 -1066 2840 -1000
rect 360 -1134 692 -1066
rect 2400 -1134 2840 -1066
rect 360 -1316 2840 -1134
rect 360 -1616 544 -1316
rect 1144 -1616 2056 -1316
rect 2656 -1616 2840 -1316
rect 360 -1800 2840 -1616
<< labels >>
flabel metal1 -26 494 -20 498 1 FreeSans 480 0 0 0 SEL
port 3 n
flabel metal2 1570 420 1578 428 1 FreeSans 480 0 0 0 A
port 1 n
flabel metal2 1824 440 1832 446 1 FreeSans 480 0 0 0 Y
port 4 n
flabel metal2 1048 442 1058 448 1 FreeSans 480 0 0 0 B
port 2 n
flabel metal2 434 442 444 452 1 FreeSans 480 0 0 0 SELB
flabel metal4 1310 3714 1322 3724 1 FreeSans 480 0 0 0 VDD
port 5 n power bidirectional
flabel metal4 1382 -1784 1396 -1776 1 FreeSans 480 0 0 0 VSS
port 6 n ground bidirectional
flabel locali 214 551 248 585 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 214 483 248 517 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 122 483 156 517 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/A
flabel nwell 79 789 113 823 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 79 245 113 279 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 79 245 113 279 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 79 789 113 823 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 50 262 50 262 4 sky130_fd_sc_hd__inv_1_0/inv_1
<< end >>
