magic
tech sky130A
magscale 1 2
timestamp 1620700822
<< error_p >>
rect -3550 -5000 -3254 5000
rect -3230 4950 -2910 4951
rect -3230 2550 -2852 4950
rect -2796 2666 -2590 4834
rect -3230 2549 -2910 2550
rect -3230 2450 -2910 2451
rect -3230 50 -2852 2450
rect -2796 166 -2590 2334
rect -3230 49 -2910 50
rect -3230 -50 -2910 -49
rect -3230 -2450 -2852 -50
rect -2796 -2334 -2590 -166
rect -3230 -2451 -2910 -2450
rect -3230 -2550 -2910 -2549
rect -3230 -4950 -2852 -2550
rect -2796 -4834 -2590 -2666
rect -3230 -4951 -2910 -4950
rect -628 -5000 -332 5000
rect -308 4950 12 4951
rect -308 2550 70 4950
rect 126 2666 332 4834
rect -308 2549 12 2550
rect -308 2450 12 2451
rect -308 50 70 2450
rect 126 166 332 2334
rect -308 49 12 50
rect -308 -50 12 -49
rect -308 -2450 70 -50
rect 126 -2334 332 -166
rect -308 -2451 12 -2450
rect -308 -2550 12 -2549
rect -308 -4950 70 -2550
rect 126 -4834 332 -2666
rect -308 -4951 12 -4950
rect 2294 -5000 2590 5000
rect 2614 4950 2934 4951
rect 2614 2550 2992 4950
rect 3048 2666 3254 4834
rect 2614 2549 2934 2550
rect 2614 2450 2934 2451
rect 2614 50 2992 2450
rect 3048 166 3254 2334
rect 2614 49 2934 50
rect 2614 -50 2934 -49
rect 2614 -2450 2992 -50
rect 3048 -2334 3254 -166
rect 2614 -2451 2934 -2450
rect 2614 -2550 2934 -2549
rect 2614 -4950 2992 -2550
rect 3048 -4834 3254 -2666
rect 2614 -4951 2934 -4950
rect 5216 -5000 5512 5000
rect 5536 2771 5832 4951
rect 5536 2549 5856 2771
rect 5536 2229 5856 2451
rect 5536 271 5832 2229
rect 5536 49 5856 271
rect 5536 -271 5856 -49
rect 5536 -2229 5832 -271
rect 5536 -2451 5856 -2229
rect 5536 -2771 5856 -2549
rect 5536 -4951 5832 -2771
<< metal4 >>
rect -5834 4909 -2932 4950
rect -5834 2591 -3188 4909
rect -2952 2591 -2932 4909
rect -5834 2550 -2932 2591
rect -2912 4909 -10 4950
rect -2912 2591 -266 4909
rect -30 2591 -10 4909
rect -2912 2550 -10 2591
rect 10 4909 2912 4950
rect 10 2591 2656 4909
rect 2892 2591 2912 4909
rect 10 2550 2912 2591
rect 2932 4909 5834 4950
rect 2932 2591 5578 4909
rect 5814 2591 5834 4909
rect 2932 2550 5834 2591
rect -5834 2409 -2932 2450
rect -5834 91 -3188 2409
rect -2952 91 -2932 2409
rect -5834 50 -2932 91
rect -2912 2409 -10 2450
rect -2912 91 -266 2409
rect -30 91 -10 2409
rect -2912 50 -10 91
rect 10 2409 2912 2450
rect 10 91 2656 2409
rect 2892 91 2912 2409
rect 10 50 2912 91
rect 2932 2409 5834 2450
rect 2932 91 5578 2409
rect 5814 91 5834 2409
rect 2932 50 5834 91
rect -5834 -91 -2932 -50
rect -5834 -2409 -3188 -91
rect -2952 -2409 -2932 -91
rect -5834 -2450 -2932 -2409
rect -2912 -91 -10 -50
rect -2912 -2409 -266 -91
rect -30 -2409 -10 -91
rect -2912 -2450 -10 -2409
rect 10 -91 2912 -50
rect 10 -2409 2656 -91
rect 2892 -2409 2912 -91
rect 10 -2450 2912 -2409
rect 2932 -91 5834 -50
rect 2932 -2409 5578 -91
rect 5814 -2409 5834 -91
rect 2932 -2450 5834 -2409
rect -5834 -2591 -2932 -2550
rect -5834 -4909 -3188 -2591
rect -2952 -4909 -2932 -2591
rect -5834 -4950 -2932 -4909
rect -2912 -2591 -10 -2550
rect -2912 -4909 -266 -2591
rect -30 -4909 -10 -2591
rect -2912 -4950 -10 -4909
rect 10 -2591 2912 -2550
rect 10 -4909 2656 -2591
rect 2892 -4909 2912 -2591
rect 10 -4950 2912 -4909
rect 2932 -2591 5834 -2550
rect 2932 -4909 5578 -2591
rect 5814 -4909 5834 -2591
rect 2932 -4950 5834 -4909
<< via4 >>
rect -3188 2591 -2952 4909
rect -266 2591 -30 4909
rect 2656 2591 2892 4909
rect 5578 2591 5814 4909
rect -3188 91 -2952 2409
rect -266 91 -30 2409
rect 2656 91 2892 2409
rect 5578 91 5814 2409
rect -3188 -2409 -2952 -91
rect -266 -2409 -30 -91
rect 2656 -2409 2892 -91
rect 5578 -2409 5814 -91
rect -3188 -4909 -2952 -2591
rect -266 -4909 -30 -2591
rect 2656 -4909 2892 -2591
rect 5578 -4909 5814 -2591
<< mimcap2 >>
rect -5734 4810 -3534 4850
rect -5734 2690 -5694 4810
rect -3574 2690 -3534 4810
rect -5734 2650 -3534 2690
rect -2812 4810 -612 4850
rect -2812 2690 -2772 4810
rect -652 2690 -612 4810
rect -2812 2650 -612 2690
rect 110 4810 2310 4850
rect 110 2690 150 4810
rect 2270 2690 2310 4810
rect 110 2650 2310 2690
rect 3032 4810 5232 4850
rect 3032 2690 3072 4810
rect 5192 2690 5232 4810
rect 3032 2650 5232 2690
rect -5734 2310 -3534 2350
rect -5734 190 -5694 2310
rect -3574 190 -3534 2310
rect -5734 150 -3534 190
rect -2812 2310 -612 2350
rect -2812 190 -2772 2310
rect -652 190 -612 2310
rect -2812 150 -612 190
rect 110 2310 2310 2350
rect 110 190 150 2310
rect 2270 190 2310 2310
rect 110 150 2310 190
rect 3032 2310 5232 2350
rect 3032 190 3072 2310
rect 5192 190 5232 2310
rect 3032 150 5232 190
rect -5734 -190 -3534 -150
rect -5734 -2310 -5694 -190
rect -3574 -2310 -3534 -190
rect -5734 -2350 -3534 -2310
rect -2812 -190 -612 -150
rect -2812 -2310 -2772 -190
rect -652 -2310 -612 -190
rect -2812 -2350 -612 -2310
rect 110 -190 2310 -150
rect 110 -2310 150 -190
rect 2270 -2310 2310 -190
rect 110 -2350 2310 -2310
rect 3032 -190 5232 -150
rect 3032 -2310 3072 -190
rect 5192 -2310 5232 -190
rect 3032 -2350 5232 -2310
rect -5734 -2690 -3534 -2650
rect -5734 -4810 -5694 -2690
rect -3574 -4810 -3534 -2690
rect -5734 -4850 -3534 -4810
rect -2812 -2690 -612 -2650
rect -2812 -4810 -2772 -2690
rect -652 -4810 -612 -2690
rect -2812 -4850 -612 -4810
rect 110 -2690 2310 -2650
rect 110 -4810 150 -2690
rect 2270 -4810 2310 -2690
rect 110 -4850 2310 -4810
rect 3032 -2690 5232 -2650
rect 3032 -4810 3072 -2690
rect 5192 -4810 5232 -2690
rect 3032 -4850 5232 -4810
<< mimcap2contact >>
rect -5694 2690 -3574 4810
rect -2772 2690 -652 4810
rect 150 2690 2270 4810
rect 3072 2690 5192 4810
rect -5694 190 -3574 2310
rect -2772 190 -652 2310
rect 150 190 2270 2310
rect 3072 190 5192 2310
rect -5694 -2310 -3574 -190
rect -2772 -2310 -652 -190
rect 150 -2310 2270 -190
rect 3072 -2310 5192 -190
rect -5694 -4810 -3574 -2690
rect -2772 -4810 -652 -2690
rect 150 -4810 2270 -2690
rect 3072 -4810 5192 -2690
<< metal5 >>
rect -4794 4834 -4474 5000
rect -3574 4834 -3254 5000
rect -5718 4810 -3254 4834
rect -5718 2690 -5694 4810
rect -3574 2690 -3254 4810
rect -5718 2666 -3254 2690
rect -4794 2334 -4474 2666
rect -3574 2334 -3254 2666
rect -3230 4909 -2910 4951
rect -3230 2591 -3188 4909
rect -2952 2591 -2910 4909
rect -1872 4834 -1552 5000
rect -652 4834 -332 5000
rect -2796 4810 -332 4834
rect -2796 2690 -2772 4810
rect -652 2690 -332 4810
rect -2796 2666 -332 2690
rect -3230 2549 -2910 2591
rect -5718 2310 -3254 2334
rect -5718 190 -5694 2310
rect -3574 190 -3254 2310
rect -5718 166 -3254 190
rect -4794 -166 -4474 166
rect -3574 -166 -3254 166
rect -3230 2409 -2910 2451
rect -3230 91 -3188 2409
rect -2952 91 -2910 2409
rect -1872 2334 -1552 2666
rect -652 2334 -332 2666
rect -308 4909 12 4951
rect -308 2591 -266 4909
rect -30 2591 12 4909
rect 1050 4834 1370 5000
rect 2270 4834 2590 5000
rect 126 4810 2590 4834
rect 126 2690 150 4810
rect 2270 2690 2590 4810
rect 126 2666 2590 2690
rect -308 2549 12 2591
rect -2796 2310 -332 2334
rect -2796 190 -2772 2310
rect -652 190 -332 2310
rect -2796 166 -332 190
rect -3230 49 -2910 91
rect -5718 -190 -3254 -166
rect -5718 -2310 -5694 -190
rect -3574 -2310 -3254 -190
rect -5718 -2334 -3254 -2310
rect -4794 -2666 -4474 -2334
rect -3574 -2666 -3254 -2334
rect -3230 -91 -2910 -49
rect -3230 -2409 -3188 -91
rect -2952 -2409 -2910 -91
rect -1872 -166 -1552 166
rect -652 -166 -332 166
rect -308 2409 12 2451
rect -308 91 -266 2409
rect -30 91 12 2409
rect 1050 2334 1370 2666
rect 2270 2334 2590 2666
rect 2614 4909 2934 4951
rect 2614 2591 2656 4909
rect 2892 2591 2934 4909
rect 3972 4834 4292 5000
rect 5192 4834 5512 5000
rect 3048 4810 5512 4834
rect 3048 2690 3072 4810
rect 5192 2690 5512 4810
rect 3048 2666 5512 2690
rect 2614 2549 2934 2591
rect 126 2310 2590 2334
rect 126 190 150 2310
rect 2270 190 2590 2310
rect 126 166 2590 190
rect -308 49 12 91
rect -2796 -190 -332 -166
rect -2796 -2310 -2772 -190
rect -652 -2310 -332 -190
rect -2796 -2334 -332 -2310
rect -3230 -2451 -2910 -2409
rect -5718 -2690 -3254 -2666
rect -5718 -4810 -5694 -2690
rect -3574 -4810 -3254 -2690
rect -5718 -4834 -3254 -4810
rect -4794 -5000 -4474 -4834
rect -3574 -5000 -3254 -4834
rect -3230 -2591 -2910 -2549
rect -3230 -4909 -3188 -2591
rect -2952 -4909 -2910 -2591
rect -1872 -2666 -1552 -2334
rect -652 -2666 -332 -2334
rect -308 -91 12 -49
rect -308 -2409 -266 -91
rect -30 -2409 12 -91
rect 1050 -166 1370 166
rect 2270 -166 2590 166
rect 2614 2409 2934 2451
rect 2614 91 2656 2409
rect 2892 91 2934 2409
rect 3972 2334 4292 2666
rect 5192 2334 5512 2666
rect 5536 4909 5856 4951
rect 5536 2591 5578 4909
rect 5814 2591 5856 4909
rect 5536 2549 5856 2591
rect 3048 2310 5512 2334
rect 3048 190 3072 2310
rect 5192 190 5512 2310
rect 3048 166 5512 190
rect 2614 49 2934 91
rect 126 -190 2590 -166
rect 126 -2310 150 -190
rect 2270 -2310 2590 -190
rect 126 -2334 2590 -2310
rect -308 -2451 12 -2409
rect -2796 -2690 -332 -2666
rect -2796 -4810 -2772 -2690
rect -652 -4810 -332 -2690
rect -2796 -4834 -332 -4810
rect -3230 -4951 -2910 -4909
rect -1872 -5000 -1552 -4834
rect -652 -5000 -332 -4834
rect -308 -2591 12 -2549
rect -308 -4909 -266 -2591
rect -30 -4909 12 -2591
rect 1050 -2666 1370 -2334
rect 2270 -2666 2590 -2334
rect 2614 -91 2934 -49
rect 2614 -2409 2656 -91
rect 2892 -2409 2934 -91
rect 3972 -166 4292 166
rect 5192 -166 5512 166
rect 5536 2409 5856 2451
rect 5536 91 5578 2409
rect 5814 91 5856 2409
rect 5536 49 5856 91
rect 3048 -190 5512 -166
rect 3048 -2310 3072 -190
rect 5192 -2310 5512 -190
rect 3048 -2334 5512 -2310
rect 2614 -2451 2934 -2409
rect 126 -2690 2590 -2666
rect 126 -4810 150 -2690
rect 2270 -4810 2590 -2690
rect 126 -4834 2590 -4810
rect -308 -4951 12 -4909
rect 1050 -5000 1370 -4834
rect 2270 -5000 2590 -4834
rect 2614 -2591 2934 -2549
rect 2614 -4909 2656 -2591
rect 2892 -4909 2934 -2591
rect 3972 -2666 4292 -2334
rect 5192 -2666 5512 -2334
rect 5536 -91 5856 -49
rect 5536 -2409 5578 -91
rect 5814 -2409 5856 -91
rect 5536 -2451 5856 -2409
rect 3048 -2690 5512 -2666
rect 3048 -4810 3072 -2690
rect 5192 -4810 5512 -2690
rect 3048 -4834 5512 -4810
rect 2614 -4951 2934 -4909
rect 3972 -5000 4292 -4834
rect 5192 -5000 5512 -4834
rect 5536 -2591 5856 -2549
rect 5536 -4909 5578 -2591
rect 5814 -4909 5856 -2591
rect 5536 -4951 5856 -4909
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX 2932 2550 5332 4950
string parameters w 11.00 l 11.00 val 128.479 carea 1.00 cperi 0.17 nx 4 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
