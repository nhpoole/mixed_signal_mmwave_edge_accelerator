magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< error_p >>
rect -1119 -100 -1061 100
rect -901 -100 -843 100
rect -683 -100 -625 100
rect -465 -100 -407 100
rect -247 -100 -189 100
rect -29 -100 29 100
rect 189 -100 247 100
rect 407 -100 465 100
rect 625 -100 683 100
rect 843 -100 901 100
rect 1061 -100 1119 100
<< nmoslvt >>
rect -1061 -100 -901 100
rect -843 -100 -683 100
rect -625 -100 -465 100
rect -407 -100 -247 100
rect -189 -100 -29 100
rect 29 -100 189 100
rect 247 -100 407 100
rect 465 -100 625 100
rect 683 -100 843 100
rect 901 -100 1061 100
<< ndiff >>
rect -1119 88 -1061 100
rect -1119 -88 -1107 88
rect -1073 -88 -1061 88
rect -1119 -100 -1061 -88
rect -901 88 -843 100
rect -901 -88 -889 88
rect -855 -88 -843 88
rect -901 -100 -843 -88
rect -683 88 -625 100
rect -683 -88 -671 88
rect -637 -88 -625 88
rect -683 -100 -625 -88
rect -465 88 -407 100
rect -465 -88 -453 88
rect -419 -88 -407 88
rect -465 -100 -407 -88
rect -247 88 -189 100
rect -247 -88 -235 88
rect -201 -88 -189 88
rect -247 -100 -189 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 189 88 247 100
rect 189 -88 201 88
rect 235 -88 247 88
rect 189 -100 247 -88
rect 407 88 465 100
rect 407 -88 419 88
rect 453 -88 465 88
rect 407 -100 465 -88
rect 625 88 683 100
rect 625 -88 637 88
rect 671 -88 683 88
rect 625 -100 683 -88
rect 843 88 901 100
rect 843 -88 855 88
rect 889 -88 901 88
rect 843 -100 901 -88
rect 1061 88 1119 100
rect 1061 -88 1073 88
rect 1107 -88 1119 88
rect 1061 -100 1119 -88
<< ndiffc >>
rect -1107 -88 -1073 88
rect -889 -88 -855 88
rect -671 -88 -637 88
rect -453 -88 -419 88
rect -235 -88 -201 88
rect -17 -88 17 88
rect 201 -88 235 88
rect 419 -88 453 88
rect 637 -88 671 88
rect 855 -88 889 88
rect 1073 -88 1107 88
<< poly >>
rect -1035 172 -927 188
rect -1035 155 -1019 172
rect -1061 138 -1019 155
rect -943 155 -927 172
rect -817 172 -709 188
rect -817 155 -801 172
rect -943 138 -901 155
rect -1061 100 -901 138
rect -843 138 -801 155
rect -725 155 -709 172
rect -599 172 -491 188
rect -599 155 -583 172
rect -725 138 -683 155
rect -843 100 -683 138
rect -625 138 -583 155
rect -507 155 -491 172
rect -381 172 -273 188
rect -381 155 -365 172
rect -507 138 -465 155
rect -625 100 -465 138
rect -407 138 -365 155
rect -289 155 -273 172
rect -163 172 -55 188
rect -163 155 -147 172
rect -289 138 -247 155
rect -407 100 -247 138
rect -189 138 -147 155
rect -71 155 -55 172
rect 55 172 163 188
rect 55 155 71 172
rect -71 138 -29 155
rect -189 100 -29 138
rect 29 138 71 155
rect 147 155 163 172
rect 273 172 381 188
rect 273 155 289 172
rect 147 138 189 155
rect 29 100 189 138
rect 247 138 289 155
rect 365 155 381 172
rect 491 172 599 188
rect 491 155 507 172
rect 365 138 407 155
rect 247 100 407 138
rect 465 138 507 155
rect 583 155 599 172
rect 709 172 817 188
rect 709 155 725 172
rect 583 138 625 155
rect 465 100 625 138
rect 683 138 725 155
rect 801 155 817 172
rect 927 172 1035 188
rect 927 155 943 172
rect 801 138 843 155
rect 683 100 843 138
rect 901 138 943 155
rect 1019 155 1035 172
rect 1019 138 1061 155
rect 901 100 1061 138
rect -1061 -138 -901 -100
rect -1061 -155 -1019 -138
rect -1035 -172 -1019 -155
rect -943 -155 -901 -138
rect -843 -138 -683 -100
rect -843 -155 -801 -138
rect -943 -172 -927 -155
rect -1035 -188 -927 -172
rect -817 -172 -801 -155
rect -725 -155 -683 -138
rect -625 -138 -465 -100
rect -625 -155 -583 -138
rect -725 -172 -709 -155
rect -817 -188 -709 -172
rect -599 -172 -583 -155
rect -507 -155 -465 -138
rect -407 -138 -247 -100
rect -407 -155 -365 -138
rect -507 -172 -491 -155
rect -599 -188 -491 -172
rect -381 -172 -365 -155
rect -289 -155 -247 -138
rect -189 -138 -29 -100
rect -189 -155 -147 -138
rect -289 -172 -273 -155
rect -381 -188 -273 -172
rect -163 -172 -147 -155
rect -71 -155 -29 -138
rect 29 -138 189 -100
rect 29 -155 71 -138
rect -71 -172 -55 -155
rect -163 -188 -55 -172
rect 55 -172 71 -155
rect 147 -155 189 -138
rect 247 -138 407 -100
rect 247 -155 289 -138
rect 147 -172 163 -155
rect 55 -188 163 -172
rect 273 -172 289 -155
rect 365 -155 407 -138
rect 465 -138 625 -100
rect 465 -155 507 -138
rect 365 -172 381 -155
rect 273 -188 381 -172
rect 491 -172 507 -155
rect 583 -155 625 -138
rect 683 -138 843 -100
rect 683 -155 725 -138
rect 583 -172 599 -155
rect 491 -188 599 -172
rect 709 -172 725 -155
rect 801 -155 843 -138
rect 901 -138 1061 -100
rect 901 -155 943 -138
rect 801 -172 817 -155
rect 709 -188 817 -172
rect 927 -172 943 -155
rect 1019 -155 1061 -138
rect 1019 -172 1035 -155
rect 927 -188 1035 -172
<< polycont >>
rect -1019 138 -943 172
rect -801 138 -725 172
rect -583 138 -507 172
rect -365 138 -289 172
rect -147 138 -71 172
rect 71 138 147 172
rect 289 138 365 172
rect 507 138 583 172
rect 725 138 801 172
rect 943 138 1019 172
rect -1019 -172 -943 -138
rect -801 -172 -725 -138
rect -583 -172 -507 -138
rect -365 -172 -289 -138
rect -147 -172 -71 -138
rect 71 -172 147 -138
rect 289 -172 365 -138
rect 507 -172 583 -138
rect 725 -172 801 -138
rect 943 -172 1019 -138
<< locali >>
rect -1035 138 -1019 172
rect -943 138 -927 172
rect -817 138 -801 172
rect -725 138 -709 172
rect -599 138 -583 172
rect -507 138 -491 172
rect -381 138 -365 172
rect -289 138 -273 172
rect -163 138 -147 172
rect -71 138 -55 172
rect 55 138 71 172
rect 147 138 163 172
rect 273 138 289 172
rect 365 138 381 172
rect 491 138 507 172
rect 583 138 599 172
rect 709 138 725 172
rect 801 138 817 172
rect 927 138 943 172
rect 1019 138 1035 172
rect -1107 88 -1073 104
rect -1107 -104 -1073 -88
rect -889 88 -855 104
rect -889 -104 -855 -88
rect -671 88 -637 104
rect -671 -104 -637 -88
rect -453 88 -419 104
rect -453 -104 -419 -88
rect -235 88 -201 104
rect -235 -104 -201 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 201 88 235 104
rect 201 -104 235 -88
rect 419 88 453 104
rect 419 -104 453 -88
rect 637 88 671 104
rect 637 -104 671 -88
rect 855 88 889 104
rect 855 -104 889 -88
rect 1073 88 1107 104
rect 1073 -104 1107 -88
rect -1035 -172 -1019 -138
rect -943 -172 -927 -138
rect -817 -172 -801 -138
rect -725 -172 -709 -138
rect -599 -172 -583 -138
rect -507 -172 -491 -138
rect -381 -172 -365 -138
rect -289 -172 -273 -138
rect -163 -172 -147 -138
rect -71 -172 -55 -138
rect 55 -172 71 -138
rect 147 -172 163 -138
rect 273 -172 289 -138
rect 365 -172 381 -138
rect 491 -172 507 -138
rect 583 -172 599 -138
rect 709 -172 725 -138
rect 801 -172 817 -138
rect 927 -172 943 -138
rect 1019 -172 1035 -138
<< viali >>
rect -1013 138 -949 172
rect -795 138 -731 172
rect -577 138 -513 172
rect -359 138 -295 172
rect -141 138 -77 172
rect 77 138 141 172
rect 295 138 359 172
rect 513 138 577 172
rect 731 138 795 172
rect 949 138 1013 172
rect -1107 -88 -1073 88
rect -889 -88 -855 88
rect -671 -88 -637 88
rect -453 -88 -419 88
rect -235 -88 -201 88
rect -17 -88 17 88
rect 201 -88 235 88
rect 419 -88 453 88
rect 637 -88 671 88
rect 855 -88 889 88
rect 1073 -88 1107 88
rect -1013 -172 -949 -138
rect -795 -172 -731 -138
rect -577 -172 -513 -138
rect -359 -172 -295 -138
rect -141 -172 -77 -138
rect 77 -172 141 -138
rect 295 -172 359 -138
rect 513 -172 577 -138
rect 731 -172 795 -138
rect 949 -172 1013 -138
<< metal1 >>
rect -1025 172 -937 178
rect -1025 138 -1013 172
rect -949 138 -937 172
rect -1025 132 -937 138
rect -807 172 -719 178
rect -807 138 -795 172
rect -731 138 -719 172
rect -807 132 -719 138
rect -589 172 -501 178
rect -589 138 -577 172
rect -513 138 -501 172
rect -589 132 -501 138
rect -371 172 -283 178
rect -371 138 -359 172
rect -295 138 -283 172
rect -371 132 -283 138
rect -153 172 -65 178
rect -153 138 -141 172
rect -77 138 -65 172
rect -153 132 -65 138
rect 65 172 153 178
rect 65 138 77 172
rect 141 138 153 172
rect 65 132 153 138
rect 283 172 371 178
rect 283 138 295 172
rect 359 138 371 172
rect 283 132 371 138
rect 501 172 589 178
rect 501 138 513 172
rect 577 138 589 172
rect 501 132 589 138
rect 719 172 807 178
rect 719 138 731 172
rect 795 138 807 172
rect 719 132 807 138
rect 937 172 1025 178
rect 937 138 949 172
rect 1013 138 1025 172
rect 937 132 1025 138
rect -1113 88 -1067 100
rect -1113 -88 -1107 88
rect -1073 -88 -1067 88
rect -1113 -100 -1067 -88
rect -895 88 -849 100
rect -895 -88 -889 88
rect -855 -88 -849 88
rect -895 -100 -849 -88
rect -677 88 -631 100
rect -677 -88 -671 88
rect -637 -88 -631 88
rect -677 -100 -631 -88
rect -459 88 -413 100
rect -459 -88 -453 88
rect -419 -88 -413 88
rect -459 -100 -413 -88
rect -241 88 -195 100
rect -241 -88 -235 88
rect -201 -88 -195 88
rect -241 -100 -195 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 195 88 241 100
rect 195 -88 201 88
rect 235 -88 241 88
rect 195 -100 241 -88
rect 413 88 459 100
rect 413 -88 419 88
rect 453 -88 459 88
rect 413 -100 459 -88
rect 631 88 677 100
rect 631 -88 637 88
rect 671 -88 677 88
rect 631 -100 677 -88
rect 849 88 895 100
rect 849 -88 855 88
rect 889 -88 895 88
rect 849 -100 895 -88
rect 1067 88 1113 100
rect 1067 -88 1073 88
rect 1107 -88 1113 88
rect 1067 -100 1113 -88
rect -1025 -138 -937 -132
rect -1025 -172 -1013 -138
rect -949 -172 -937 -138
rect -1025 -178 -937 -172
rect -807 -138 -719 -132
rect -807 -172 -795 -138
rect -731 -172 -719 -138
rect -807 -178 -719 -172
rect -589 -138 -501 -132
rect -589 -172 -577 -138
rect -513 -172 -501 -138
rect -589 -178 -501 -172
rect -371 -138 -283 -132
rect -371 -172 -359 -138
rect -295 -172 -283 -138
rect -371 -178 -283 -172
rect -153 -138 -65 -132
rect -153 -172 -141 -138
rect -77 -172 -65 -138
rect -153 -178 -65 -172
rect 65 -138 153 -132
rect 65 -172 77 -138
rect 141 -172 153 -138
rect 65 -178 153 -172
rect 283 -138 371 -132
rect 283 -172 295 -138
rect 359 -172 371 -138
rect 283 -178 371 -172
rect 501 -138 589 -132
rect 501 -172 513 -138
rect 577 -172 589 -138
rect 501 -178 589 -172
rect 719 -138 807 -132
rect 719 -172 731 -138
rect 795 -172 807 -138
rect 719 -178 807 -172
rect 937 -138 1025 -132
rect 937 -172 949 -138
rect 1013 -172 1025 -138
rect 937 -178 1025 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string parameters w 1 l 0.8 m 1 nf 10 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
