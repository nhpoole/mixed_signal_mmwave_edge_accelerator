magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1289 -1283 1289 1283
<< viali >>
rect -17 -17 17 17
<< metal1 >>
rect -29 17 29 23
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -23 29 -17
<< end >>
