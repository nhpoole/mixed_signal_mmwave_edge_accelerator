magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -2210 -1560 2078 1560
<< metal3 >>
rect -950 -300 818 300
<< mimcap >>
rect -850 152 750 200
rect -850 -152 -802 152
rect 702 -152 750 152
rect -850 -200 750 -152
<< mimcapcontact >>
rect -802 -152 702 152
<< metal4 >>
rect -811 152 711 161
rect -811 -152 -802 152
rect 702 -152 711 152
rect -811 -161 711 -152
<< properties >>
string FIXED_BBOX -950 -300 850 300
<< end >>
