magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1476 -1529 1476 1529
<< pwell >>
rect -216 -269 216 269
<< nmos >>
rect -30 -131 30 69
<< ndiff >>
rect -88 54 -30 69
rect -88 20 -76 54
rect -42 20 -30 54
rect -88 -14 -30 20
rect -88 -48 -76 -14
rect -42 -48 -30 -14
rect -88 -82 -30 -48
rect -88 -116 -76 -82
rect -42 -116 -30 -82
rect -88 -131 -30 -116
rect 30 54 88 69
rect 30 20 42 54
rect 76 20 88 54
rect 30 -14 88 20
rect 30 -48 42 -14
rect 76 -48 88 -14
rect 30 -82 88 -48
rect 30 -116 42 -82
rect 76 -116 88 -82
rect 30 -131 88 -116
<< ndiffc >>
rect -76 20 -42 54
rect -76 -48 -42 -14
rect -76 -116 -42 -82
rect 42 20 76 54
rect 42 -48 76 -14
rect 42 -116 76 -82
<< psubdiff >>
rect -190 209 -85 243
rect -51 209 -17 243
rect 17 209 51 243
rect 85 209 190 243
rect -190 119 -156 209
rect 156 119 190 209
rect -190 51 -156 85
rect -190 -17 -156 17
rect -190 -85 -156 -51
rect -190 -209 -156 -119
rect 156 51 190 85
rect 156 -17 190 17
rect 156 -85 190 -51
rect 156 -209 190 -119
rect -190 -243 -85 -209
rect -51 -243 -17 -209
rect 17 -243 51 -209
rect 85 -243 190 -209
<< psubdiffcont >>
rect -85 209 -51 243
rect -17 209 17 243
rect 51 209 85 243
rect -190 85 -156 119
rect 156 85 190 119
rect -190 17 -156 51
rect -190 -51 -156 -17
rect -190 -119 -156 -85
rect 156 17 190 51
rect 156 -51 190 -17
rect 156 -119 190 -85
rect -85 -243 -51 -209
rect -17 -243 17 -209
rect 51 -243 85 -209
<< poly >>
rect -33 141 33 157
rect -33 107 -17 141
rect 17 107 33 141
rect -33 91 33 107
rect -30 69 30 91
rect -30 -157 30 -131
<< polycont >>
rect -17 107 17 141
<< locali >>
rect -190 209 -85 243
rect -51 209 -17 243
rect 17 209 51 243
rect 85 209 190 243
rect -190 119 -156 209
rect -33 107 -17 141
rect 17 107 33 141
rect 156 119 190 209
rect -190 51 -156 85
rect -190 -17 -156 17
rect -190 -85 -156 -51
rect -190 -209 -156 -119
rect -76 54 -42 73
rect -76 -14 -42 -12
rect -76 -50 -42 -48
rect -76 -135 -42 -116
rect 42 54 76 73
rect 42 -14 76 -12
rect 42 -50 76 -48
rect 42 -135 76 -116
rect 156 51 190 85
rect 156 -17 190 17
rect 156 -85 190 -51
rect 156 -209 190 -119
rect -190 -243 -85 -209
rect -51 -243 -17 -209
rect 17 -243 51 -209
rect 85 -243 190 -209
<< viali >>
rect -17 107 17 141
rect -76 20 -42 22
rect -76 -12 -42 20
rect -76 -82 -42 -50
rect -76 -84 -42 -82
rect 42 20 76 22
rect 42 -12 76 20
rect 42 -82 76 -50
rect 42 -84 76 -82
<< metal1 >>
rect -29 141 29 147
rect -29 107 -17 141
rect 17 107 29 141
rect -29 101 29 107
rect -82 22 -36 69
rect -82 -12 -76 22
rect -42 -12 -36 22
rect -82 -50 -36 -12
rect -82 -84 -76 -50
rect -42 -84 -36 -50
rect -82 -131 -36 -84
rect 36 22 82 69
rect 36 -12 42 22
rect 76 -12 82 22
rect 36 -50 82 -12
rect 36 -84 42 -50
rect 76 -84 82 -50
rect 36 -131 82 -84
<< properties >>
string FIXED_BBOX -173 -226 173 226
<< end >>
