magic
tech sky130A
magscale 1 2
timestamp 1622323610
<< error_p >>
rect -160 -217 160 217
<< metal5 >>
rect -160 160 160 217
rect -160 -217 160 -160
<< rm5 >>
rect -160 -160 160 160
<< properties >>
string gencell sky130_fd_pr__res_generic_m5
string parameters w 1.600 l 1.600 m 1 nx 1 wmin 1.60 lmin 1.60 rho 0.029 val 29.0m dummy 0 dw 0.0 term 0.0 roverlap 0
string library sky130
<< end >>
