magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -3605 -1448 3605 1448
<< pwell >>
rect -2345 -126 2345 126
<< nmos >>
rect -2261 -100 -1861 100
rect -1803 -100 -1403 100
rect -1345 -100 -945 100
rect -887 -100 -487 100
rect -429 -100 -29 100
rect 29 -100 429 100
rect 487 -100 887 100
rect 945 -100 1345 100
rect 1403 -100 1803 100
rect 1861 -100 2261 100
<< ndiff >>
rect -2319 85 -2261 100
rect -2319 51 -2307 85
rect -2273 51 -2261 85
rect -2319 17 -2261 51
rect -2319 -17 -2307 17
rect -2273 -17 -2261 17
rect -2319 -51 -2261 -17
rect -2319 -85 -2307 -51
rect -2273 -85 -2261 -51
rect -2319 -100 -2261 -85
rect -1861 85 -1803 100
rect -1861 51 -1849 85
rect -1815 51 -1803 85
rect -1861 17 -1803 51
rect -1861 -17 -1849 17
rect -1815 -17 -1803 17
rect -1861 -51 -1803 -17
rect -1861 -85 -1849 -51
rect -1815 -85 -1803 -51
rect -1861 -100 -1803 -85
rect -1403 85 -1345 100
rect -1403 51 -1391 85
rect -1357 51 -1345 85
rect -1403 17 -1345 51
rect -1403 -17 -1391 17
rect -1357 -17 -1345 17
rect -1403 -51 -1345 -17
rect -1403 -85 -1391 -51
rect -1357 -85 -1345 -51
rect -1403 -100 -1345 -85
rect -945 85 -887 100
rect -945 51 -933 85
rect -899 51 -887 85
rect -945 17 -887 51
rect -945 -17 -933 17
rect -899 -17 -887 17
rect -945 -51 -887 -17
rect -945 -85 -933 -51
rect -899 -85 -887 -51
rect -945 -100 -887 -85
rect -487 85 -429 100
rect -487 51 -475 85
rect -441 51 -429 85
rect -487 17 -429 51
rect -487 -17 -475 17
rect -441 -17 -429 17
rect -487 -51 -429 -17
rect -487 -85 -475 -51
rect -441 -85 -429 -51
rect -487 -100 -429 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 429 85 487 100
rect 429 51 441 85
rect 475 51 487 85
rect 429 17 487 51
rect 429 -17 441 17
rect 475 -17 487 17
rect 429 -51 487 -17
rect 429 -85 441 -51
rect 475 -85 487 -51
rect 429 -100 487 -85
rect 887 85 945 100
rect 887 51 899 85
rect 933 51 945 85
rect 887 17 945 51
rect 887 -17 899 17
rect 933 -17 945 17
rect 887 -51 945 -17
rect 887 -85 899 -51
rect 933 -85 945 -51
rect 887 -100 945 -85
rect 1345 85 1403 100
rect 1345 51 1357 85
rect 1391 51 1403 85
rect 1345 17 1403 51
rect 1345 -17 1357 17
rect 1391 -17 1403 17
rect 1345 -51 1403 -17
rect 1345 -85 1357 -51
rect 1391 -85 1403 -51
rect 1345 -100 1403 -85
rect 1803 85 1861 100
rect 1803 51 1815 85
rect 1849 51 1861 85
rect 1803 17 1861 51
rect 1803 -17 1815 17
rect 1849 -17 1861 17
rect 1803 -51 1861 -17
rect 1803 -85 1815 -51
rect 1849 -85 1861 -51
rect 1803 -100 1861 -85
rect 2261 85 2319 100
rect 2261 51 2273 85
rect 2307 51 2319 85
rect 2261 17 2319 51
rect 2261 -17 2273 17
rect 2307 -17 2319 17
rect 2261 -51 2319 -17
rect 2261 -85 2273 -51
rect 2307 -85 2319 -51
rect 2261 -100 2319 -85
<< ndiffc >>
rect -2307 51 -2273 85
rect -2307 -17 -2273 17
rect -2307 -85 -2273 -51
rect -1849 51 -1815 85
rect -1849 -17 -1815 17
rect -1849 -85 -1815 -51
rect -1391 51 -1357 85
rect -1391 -17 -1357 17
rect -1391 -85 -1357 -51
rect -933 51 -899 85
rect -933 -17 -899 17
rect -933 -85 -899 -51
rect -475 51 -441 85
rect -475 -17 -441 17
rect -475 -85 -441 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 441 51 475 85
rect 441 -17 475 17
rect 441 -85 475 -51
rect 899 51 933 85
rect 899 -17 933 17
rect 899 -85 933 -51
rect 1357 51 1391 85
rect 1357 -17 1391 17
rect 1357 -85 1391 -51
rect 1815 51 1849 85
rect 1815 -17 1849 17
rect 1815 -85 1849 -51
rect 2273 51 2307 85
rect 2273 -17 2307 17
rect 2273 -85 2307 -51
<< poly >>
rect -2187 172 -1935 188
rect -2187 155 -2146 172
rect -2261 138 -2146 155
rect -2112 138 -2078 172
rect -2044 138 -2010 172
rect -1976 155 -1935 172
rect -1729 172 -1477 188
rect -1729 155 -1688 172
rect -1976 138 -1861 155
rect -2261 100 -1861 138
rect -1803 138 -1688 155
rect -1654 138 -1620 172
rect -1586 138 -1552 172
rect -1518 155 -1477 172
rect -1271 172 -1019 188
rect -1271 155 -1230 172
rect -1518 138 -1403 155
rect -1803 100 -1403 138
rect -1345 138 -1230 155
rect -1196 138 -1162 172
rect -1128 138 -1094 172
rect -1060 155 -1019 172
rect -813 172 -561 188
rect -813 155 -772 172
rect -1060 138 -945 155
rect -1345 100 -945 138
rect -887 138 -772 155
rect -738 138 -704 172
rect -670 138 -636 172
rect -602 155 -561 172
rect -355 172 -103 188
rect -355 155 -314 172
rect -602 138 -487 155
rect -887 100 -487 138
rect -429 138 -314 155
rect -280 138 -246 172
rect -212 138 -178 172
rect -144 155 -103 172
rect 103 172 355 188
rect 103 155 144 172
rect -144 138 -29 155
rect -429 100 -29 138
rect 29 138 144 155
rect 178 138 212 172
rect 246 138 280 172
rect 314 155 355 172
rect 561 172 813 188
rect 561 155 602 172
rect 314 138 429 155
rect 29 100 429 138
rect 487 138 602 155
rect 636 138 670 172
rect 704 138 738 172
rect 772 155 813 172
rect 1019 172 1271 188
rect 1019 155 1060 172
rect 772 138 887 155
rect 487 100 887 138
rect 945 138 1060 155
rect 1094 138 1128 172
rect 1162 138 1196 172
rect 1230 155 1271 172
rect 1477 172 1729 188
rect 1477 155 1518 172
rect 1230 138 1345 155
rect 945 100 1345 138
rect 1403 138 1518 155
rect 1552 138 1586 172
rect 1620 138 1654 172
rect 1688 155 1729 172
rect 1935 172 2187 188
rect 1935 155 1976 172
rect 1688 138 1803 155
rect 1403 100 1803 138
rect 1861 138 1976 155
rect 2010 138 2044 172
rect 2078 138 2112 172
rect 2146 155 2187 172
rect 2146 138 2261 155
rect 1861 100 2261 138
rect -2261 -138 -1861 -100
rect -2261 -155 -2146 -138
rect -2187 -172 -2146 -155
rect -2112 -172 -2078 -138
rect -2044 -172 -2010 -138
rect -1976 -155 -1861 -138
rect -1803 -138 -1403 -100
rect -1803 -155 -1688 -138
rect -1976 -172 -1935 -155
rect -2187 -188 -1935 -172
rect -1729 -172 -1688 -155
rect -1654 -172 -1620 -138
rect -1586 -172 -1552 -138
rect -1518 -155 -1403 -138
rect -1345 -138 -945 -100
rect -1345 -155 -1230 -138
rect -1518 -172 -1477 -155
rect -1729 -188 -1477 -172
rect -1271 -172 -1230 -155
rect -1196 -172 -1162 -138
rect -1128 -172 -1094 -138
rect -1060 -155 -945 -138
rect -887 -138 -487 -100
rect -887 -155 -772 -138
rect -1060 -172 -1019 -155
rect -1271 -188 -1019 -172
rect -813 -172 -772 -155
rect -738 -172 -704 -138
rect -670 -172 -636 -138
rect -602 -155 -487 -138
rect -429 -138 -29 -100
rect -429 -155 -314 -138
rect -602 -172 -561 -155
rect -813 -188 -561 -172
rect -355 -172 -314 -155
rect -280 -172 -246 -138
rect -212 -172 -178 -138
rect -144 -155 -29 -138
rect 29 -138 429 -100
rect 29 -155 144 -138
rect -144 -172 -103 -155
rect -355 -188 -103 -172
rect 103 -172 144 -155
rect 178 -172 212 -138
rect 246 -172 280 -138
rect 314 -155 429 -138
rect 487 -138 887 -100
rect 487 -155 602 -138
rect 314 -172 355 -155
rect 103 -188 355 -172
rect 561 -172 602 -155
rect 636 -172 670 -138
rect 704 -172 738 -138
rect 772 -155 887 -138
rect 945 -138 1345 -100
rect 945 -155 1060 -138
rect 772 -172 813 -155
rect 561 -188 813 -172
rect 1019 -172 1060 -155
rect 1094 -172 1128 -138
rect 1162 -172 1196 -138
rect 1230 -155 1345 -138
rect 1403 -138 1803 -100
rect 1403 -155 1518 -138
rect 1230 -172 1271 -155
rect 1019 -188 1271 -172
rect 1477 -172 1518 -155
rect 1552 -172 1586 -138
rect 1620 -172 1654 -138
rect 1688 -155 1803 -138
rect 1861 -138 2261 -100
rect 1861 -155 1976 -138
rect 1688 -172 1729 -155
rect 1477 -188 1729 -172
rect 1935 -172 1976 -155
rect 2010 -172 2044 -138
rect 2078 -172 2112 -138
rect 2146 -155 2261 -138
rect 2146 -172 2187 -155
rect 1935 -188 2187 -172
<< polycont >>
rect -2146 138 -2112 172
rect -2078 138 -2044 172
rect -2010 138 -1976 172
rect -1688 138 -1654 172
rect -1620 138 -1586 172
rect -1552 138 -1518 172
rect -1230 138 -1196 172
rect -1162 138 -1128 172
rect -1094 138 -1060 172
rect -772 138 -738 172
rect -704 138 -670 172
rect -636 138 -602 172
rect -314 138 -280 172
rect -246 138 -212 172
rect -178 138 -144 172
rect 144 138 178 172
rect 212 138 246 172
rect 280 138 314 172
rect 602 138 636 172
rect 670 138 704 172
rect 738 138 772 172
rect 1060 138 1094 172
rect 1128 138 1162 172
rect 1196 138 1230 172
rect 1518 138 1552 172
rect 1586 138 1620 172
rect 1654 138 1688 172
rect 1976 138 2010 172
rect 2044 138 2078 172
rect 2112 138 2146 172
rect -2146 -172 -2112 -138
rect -2078 -172 -2044 -138
rect -2010 -172 -1976 -138
rect -1688 -172 -1654 -138
rect -1620 -172 -1586 -138
rect -1552 -172 -1518 -138
rect -1230 -172 -1196 -138
rect -1162 -172 -1128 -138
rect -1094 -172 -1060 -138
rect -772 -172 -738 -138
rect -704 -172 -670 -138
rect -636 -172 -602 -138
rect -314 -172 -280 -138
rect -246 -172 -212 -138
rect -178 -172 -144 -138
rect 144 -172 178 -138
rect 212 -172 246 -138
rect 280 -172 314 -138
rect 602 -172 636 -138
rect 670 -172 704 -138
rect 738 -172 772 -138
rect 1060 -172 1094 -138
rect 1128 -172 1162 -138
rect 1196 -172 1230 -138
rect 1518 -172 1552 -138
rect 1586 -172 1620 -138
rect 1654 -172 1688 -138
rect 1976 -172 2010 -138
rect 2044 -172 2078 -138
rect 2112 -172 2146 -138
<< locali >>
rect -2187 138 -2150 172
rect -2112 138 -2078 172
rect -2044 138 -2010 172
rect -1972 138 -1935 172
rect -1729 138 -1692 172
rect -1654 138 -1620 172
rect -1586 138 -1552 172
rect -1514 138 -1477 172
rect -1271 138 -1234 172
rect -1196 138 -1162 172
rect -1128 138 -1094 172
rect -1056 138 -1019 172
rect -813 138 -776 172
rect -738 138 -704 172
rect -670 138 -636 172
rect -598 138 -561 172
rect -355 138 -318 172
rect -280 138 -246 172
rect -212 138 -178 172
rect -140 138 -103 172
rect 103 138 140 172
rect 178 138 212 172
rect 246 138 280 172
rect 318 138 355 172
rect 561 138 598 172
rect 636 138 670 172
rect 704 138 738 172
rect 776 138 813 172
rect 1019 138 1056 172
rect 1094 138 1128 172
rect 1162 138 1196 172
rect 1234 138 1271 172
rect 1477 138 1514 172
rect 1552 138 1586 172
rect 1620 138 1654 172
rect 1692 138 1729 172
rect 1935 138 1972 172
rect 2010 138 2044 172
rect 2078 138 2112 172
rect 2150 138 2187 172
rect -2307 85 -2273 104
rect -2307 17 -2273 19
rect -2307 -19 -2273 -17
rect -2307 -104 -2273 -85
rect -1849 85 -1815 104
rect -1849 17 -1815 19
rect -1849 -19 -1815 -17
rect -1849 -104 -1815 -85
rect -1391 85 -1357 104
rect -1391 17 -1357 19
rect -1391 -19 -1357 -17
rect -1391 -104 -1357 -85
rect -933 85 -899 104
rect -933 17 -899 19
rect -933 -19 -899 -17
rect -933 -104 -899 -85
rect -475 85 -441 104
rect -475 17 -441 19
rect -475 -19 -441 -17
rect -475 -104 -441 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 441 85 475 104
rect 441 17 475 19
rect 441 -19 475 -17
rect 441 -104 475 -85
rect 899 85 933 104
rect 899 17 933 19
rect 899 -19 933 -17
rect 899 -104 933 -85
rect 1357 85 1391 104
rect 1357 17 1391 19
rect 1357 -19 1391 -17
rect 1357 -104 1391 -85
rect 1815 85 1849 104
rect 1815 17 1849 19
rect 1815 -19 1849 -17
rect 1815 -104 1849 -85
rect 2273 85 2307 104
rect 2273 17 2307 19
rect 2273 -19 2307 -17
rect 2273 -104 2307 -85
rect -2187 -172 -2150 -138
rect -2112 -172 -2078 -138
rect -2044 -172 -2010 -138
rect -1972 -172 -1935 -138
rect -1729 -172 -1692 -138
rect -1654 -172 -1620 -138
rect -1586 -172 -1552 -138
rect -1514 -172 -1477 -138
rect -1271 -172 -1234 -138
rect -1196 -172 -1162 -138
rect -1128 -172 -1094 -138
rect -1056 -172 -1019 -138
rect -813 -172 -776 -138
rect -738 -172 -704 -138
rect -670 -172 -636 -138
rect -598 -172 -561 -138
rect -355 -172 -318 -138
rect -280 -172 -246 -138
rect -212 -172 -178 -138
rect -140 -172 -103 -138
rect 103 -172 140 -138
rect 178 -172 212 -138
rect 246 -172 280 -138
rect 318 -172 355 -138
rect 561 -172 598 -138
rect 636 -172 670 -138
rect 704 -172 738 -138
rect 776 -172 813 -138
rect 1019 -172 1056 -138
rect 1094 -172 1128 -138
rect 1162 -172 1196 -138
rect 1234 -172 1271 -138
rect 1477 -172 1514 -138
rect 1552 -172 1586 -138
rect 1620 -172 1654 -138
rect 1692 -172 1729 -138
rect 1935 -172 1972 -138
rect 2010 -172 2044 -138
rect 2078 -172 2112 -138
rect 2150 -172 2187 -138
<< viali >>
rect -2150 138 -2146 172
rect -2146 138 -2116 172
rect -2078 138 -2044 172
rect -2006 138 -1976 172
rect -1976 138 -1972 172
rect -1692 138 -1688 172
rect -1688 138 -1658 172
rect -1620 138 -1586 172
rect -1548 138 -1518 172
rect -1518 138 -1514 172
rect -1234 138 -1230 172
rect -1230 138 -1200 172
rect -1162 138 -1128 172
rect -1090 138 -1060 172
rect -1060 138 -1056 172
rect -776 138 -772 172
rect -772 138 -742 172
rect -704 138 -670 172
rect -632 138 -602 172
rect -602 138 -598 172
rect -318 138 -314 172
rect -314 138 -284 172
rect -246 138 -212 172
rect -174 138 -144 172
rect -144 138 -140 172
rect 140 138 144 172
rect 144 138 174 172
rect 212 138 246 172
rect 284 138 314 172
rect 314 138 318 172
rect 598 138 602 172
rect 602 138 632 172
rect 670 138 704 172
rect 742 138 772 172
rect 772 138 776 172
rect 1056 138 1060 172
rect 1060 138 1090 172
rect 1128 138 1162 172
rect 1200 138 1230 172
rect 1230 138 1234 172
rect 1514 138 1518 172
rect 1518 138 1548 172
rect 1586 138 1620 172
rect 1658 138 1688 172
rect 1688 138 1692 172
rect 1972 138 1976 172
rect 1976 138 2006 172
rect 2044 138 2078 172
rect 2116 138 2146 172
rect 2146 138 2150 172
rect -2307 51 -2273 53
rect -2307 19 -2273 51
rect -2307 -51 -2273 -19
rect -2307 -53 -2273 -51
rect -1849 51 -1815 53
rect -1849 19 -1815 51
rect -1849 -51 -1815 -19
rect -1849 -53 -1815 -51
rect -1391 51 -1357 53
rect -1391 19 -1357 51
rect -1391 -51 -1357 -19
rect -1391 -53 -1357 -51
rect -933 51 -899 53
rect -933 19 -899 51
rect -933 -51 -899 -19
rect -933 -53 -899 -51
rect -475 51 -441 53
rect -475 19 -441 51
rect -475 -51 -441 -19
rect -475 -53 -441 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 441 51 475 53
rect 441 19 475 51
rect 441 -51 475 -19
rect 441 -53 475 -51
rect 899 51 933 53
rect 899 19 933 51
rect 899 -51 933 -19
rect 899 -53 933 -51
rect 1357 51 1391 53
rect 1357 19 1391 51
rect 1357 -51 1391 -19
rect 1357 -53 1391 -51
rect 1815 51 1849 53
rect 1815 19 1849 51
rect 1815 -51 1849 -19
rect 1815 -53 1849 -51
rect 2273 51 2307 53
rect 2273 19 2307 51
rect 2273 -51 2307 -19
rect 2273 -53 2307 -51
rect -2150 -172 -2146 -138
rect -2146 -172 -2116 -138
rect -2078 -172 -2044 -138
rect -2006 -172 -1976 -138
rect -1976 -172 -1972 -138
rect -1692 -172 -1688 -138
rect -1688 -172 -1658 -138
rect -1620 -172 -1586 -138
rect -1548 -172 -1518 -138
rect -1518 -172 -1514 -138
rect -1234 -172 -1230 -138
rect -1230 -172 -1200 -138
rect -1162 -172 -1128 -138
rect -1090 -172 -1060 -138
rect -1060 -172 -1056 -138
rect -776 -172 -772 -138
rect -772 -172 -742 -138
rect -704 -172 -670 -138
rect -632 -172 -602 -138
rect -602 -172 -598 -138
rect -318 -172 -314 -138
rect -314 -172 -284 -138
rect -246 -172 -212 -138
rect -174 -172 -144 -138
rect -144 -172 -140 -138
rect 140 -172 144 -138
rect 144 -172 174 -138
rect 212 -172 246 -138
rect 284 -172 314 -138
rect 314 -172 318 -138
rect 598 -172 602 -138
rect 602 -172 632 -138
rect 670 -172 704 -138
rect 742 -172 772 -138
rect 772 -172 776 -138
rect 1056 -172 1060 -138
rect 1060 -172 1090 -138
rect 1128 -172 1162 -138
rect 1200 -172 1230 -138
rect 1230 -172 1234 -138
rect 1514 -172 1518 -138
rect 1518 -172 1548 -138
rect 1586 -172 1620 -138
rect 1658 -172 1688 -138
rect 1688 -172 1692 -138
rect 1972 -172 1976 -138
rect 1976 -172 2006 -138
rect 2044 -172 2078 -138
rect 2116 -172 2146 -138
rect 2146 -172 2150 -138
<< metal1 >>
rect -2165 172 -1957 178
rect -2165 138 -2150 172
rect -2116 138 -2078 172
rect -2044 138 -2006 172
rect -1972 138 -1957 172
rect -2165 132 -1957 138
rect -1707 172 -1499 178
rect -1707 138 -1692 172
rect -1658 138 -1620 172
rect -1586 138 -1548 172
rect -1514 138 -1499 172
rect -1707 132 -1499 138
rect -1249 172 -1041 178
rect -1249 138 -1234 172
rect -1200 138 -1162 172
rect -1128 138 -1090 172
rect -1056 138 -1041 172
rect -1249 132 -1041 138
rect -791 172 -583 178
rect -791 138 -776 172
rect -742 138 -704 172
rect -670 138 -632 172
rect -598 138 -583 172
rect -791 132 -583 138
rect -333 172 -125 178
rect -333 138 -318 172
rect -284 138 -246 172
rect -212 138 -174 172
rect -140 138 -125 172
rect -333 132 -125 138
rect 125 172 333 178
rect 125 138 140 172
rect 174 138 212 172
rect 246 138 284 172
rect 318 138 333 172
rect 125 132 333 138
rect 583 172 791 178
rect 583 138 598 172
rect 632 138 670 172
rect 704 138 742 172
rect 776 138 791 172
rect 583 132 791 138
rect 1041 172 1249 178
rect 1041 138 1056 172
rect 1090 138 1128 172
rect 1162 138 1200 172
rect 1234 138 1249 172
rect 1041 132 1249 138
rect 1499 172 1707 178
rect 1499 138 1514 172
rect 1548 138 1586 172
rect 1620 138 1658 172
rect 1692 138 1707 172
rect 1499 132 1707 138
rect 1957 172 2165 178
rect 1957 138 1972 172
rect 2006 138 2044 172
rect 2078 138 2116 172
rect 2150 138 2165 172
rect 1957 132 2165 138
rect -2313 53 -2267 100
rect -2313 19 -2307 53
rect -2273 19 -2267 53
rect -2313 -19 -2267 19
rect -2313 -53 -2307 -19
rect -2273 -53 -2267 -19
rect -2313 -100 -2267 -53
rect -1855 53 -1809 100
rect -1855 19 -1849 53
rect -1815 19 -1809 53
rect -1855 -19 -1809 19
rect -1855 -53 -1849 -19
rect -1815 -53 -1809 -19
rect -1855 -100 -1809 -53
rect -1397 53 -1351 100
rect -1397 19 -1391 53
rect -1357 19 -1351 53
rect -1397 -19 -1351 19
rect -1397 -53 -1391 -19
rect -1357 -53 -1351 -19
rect -1397 -100 -1351 -53
rect -939 53 -893 100
rect -939 19 -933 53
rect -899 19 -893 53
rect -939 -19 -893 19
rect -939 -53 -933 -19
rect -899 -53 -893 -19
rect -939 -100 -893 -53
rect -481 53 -435 100
rect -481 19 -475 53
rect -441 19 -435 53
rect -481 -19 -435 19
rect -481 -53 -475 -19
rect -441 -53 -435 -19
rect -481 -100 -435 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 435 53 481 100
rect 435 19 441 53
rect 475 19 481 53
rect 435 -19 481 19
rect 435 -53 441 -19
rect 475 -53 481 -19
rect 435 -100 481 -53
rect 893 53 939 100
rect 893 19 899 53
rect 933 19 939 53
rect 893 -19 939 19
rect 893 -53 899 -19
rect 933 -53 939 -19
rect 893 -100 939 -53
rect 1351 53 1397 100
rect 1351 19 1357 53
rect 1391 19 1397 53
rect 1351 -19 1397 19
rect 1351 -53 1357 -19
rect 1391 -53 1397 -19
rect 1351 -100 1397 -53
rect 1809 53 1855 100
rect 1809 19 1815 53
rect 1849 19 1855 53
rect 1809 -19 1855 19
rect 1809 -53 1815 -19
rect 1849 -53 1855 -19
rect 1809 -100 1855 -53
rect 2267 53 2313 100
rect 2267 19 2273 53
rect 2307 19 2313 53
rect 2267 -19 2313 19
rect 2267 -53 2273 -19
rect 2307 -53 2313 -19
rect 2267 -100 2313 -53
rect -2165 -138 -1957 -132
rect -2165 -172 -2150 -138
rect -2116 -172 -2078 -138
rect -2044 -172 -2006 -138
rect -1972 -172 -1957 -138
rect -2165 -178 -1957 -172
rect -1707 -138 -1499 -132
rect -1707 -172 -1692 -138
rect -1658 -172 -1620 -138
rect -1586 -172 -1548 -138
rect -1514 -172 -1499 -138
rect -1707 -178 -1499 -172
rect -1249 -138 -1041 -132
rect -1249 -172 -1234 -138
rect -1200 -172 -1162 -138
rect -1128 -172 -1090 -138
rect -1056 -172 -1041 -138
rect -1249 -178 -1041 -172
rect -791 -138 -583 -132
rect -791 -172 -776 -138
rect -742 -172 -704 -138
rect -670 -172 -632 -138
rect -598 -172 -583 -138
rect -791 -178 -583 -172
rect -333 -138 -125 -132
rect -333 -172 -318 -138
rect -284 -172 -246 -138
rect -212 -172 -174 -138
rect -140 -172 -125 -138
rect -333 -178 -125 -172
rect 125 -138 333 -132
rect 125 -172 140 -138
rect 174 -172 212 -138
rect 246 -172 284 -138
rect 318 -172 333 -138
rect 125 -178 333 -172
rect 583 -138 791 -132
rect 583 -172 598 -138
rect 632 -172 670 -138
rect 704 -172 742 -138
rect 776 -172 791 -138
rect 583 -178 791 -172
rect 1041 -138 1249 -132
rect 1041 -172 1056 -138
rect 1090 -172 1128 -138
rect 1162 -172 1200 -138
rect 1234 -172 1249 -138
rect 1041 -178 1249 -172
rect 1499 -138 1707 -132
rect 1499 -172 1514 -138
rect 1548 -172 1586 -138
rect 1620 -172 1658 -138
rect 1692 -172 1707 -138
rect 1499 -178 1707 -172
rect 1957 -138 2165 -132
rect 1957 -172 1972 -138
rect 2006 -172 2044 -138
rect 2078 -172 2116 -138
rect 2150 -172 2165 -138
rect 1957 -178 2165 -172
<< end >>
