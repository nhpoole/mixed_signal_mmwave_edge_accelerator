magic
tech sky130A
magscale 1 2
timestamp 1623661481
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 30 -17 64 17
<< locali >>
rect 18 197 66 325
rect 288 191 354 265
rect 1131 375 1185 493
rect 1151 300 1185 375
rect 1151 285 1271 300
rect 1152 283 1271 285
rect 1153 282 1271 283
rect 1155 277 1271 282
rect 896 207 1048 265
rect 896 199 963 207
rect 1157 178 1271 277
rect 1154 173 1271 178
rect 1151 153 1271 173
rect 1151 97 1185 153
rect 1119 51 1185 97
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 35 393 69 493
rect 103 427 169 527
rect 35 359 156 393
rect 122 280 156 359
rect 203 337 248 493
rect 122 214 168 280
rect 122 161 156 214
rect 17 127 156 161
rect 17 69 69 127
rect 103 17 169 93
rect 203 69 237 337
rect 287 333 357 483
rect 391 367 450 527
rect 554 451 716 485
rect 682 417 716 451
rect 750 435 818 527
rect 856 427 912 527
rect 682 400 721 417
rect 683 399 721 400
rect 581 382 635 399
rect 684 397 721 399
rect 581 356 653 382
rect 287 299 424 333
rect 390 219 424 299
rect 490 271 551 337
rect 586 314 653 356
rect 390 157 467 219
rect 586 208 620 314
rect 687 265 721 397
rect 960 373 994 493
rect 1028 375 1097 527
rect 755 341 994 373
rect 755 307 1117 341
rect 1083 265 1117 307
rect 1219 334 1271 527
rect 303 153 467 157
rect 303 123 424 153
rect 517 147 620 208
rect 654 199 844 265
rect 1083 199 1123 265
rect 303 69 341 123
rect 654 107 689 199
rect 1083 173 1117 199
rect 991 165 1117 173
rect 375 17 441 89
rect 554 73 689 107
rect 848 139 1117 165
rect 848 131 1019 139
rect 744 17 812 106
rect 848 51 916 131
rect 1051 17 1085 105
rect 1219 17 1271 119
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< obsm1 >>
rect 202 388 260 397
rect 573 388 631 397
rect 202 360 631 388
rect 202 351 260 360
rect 573 351 631 360
rect 110 320 168 329
rect 478 320 536 329
rect 110 292 536 320
rect 110 283 168 292
rect 478 283 536 292
<< labels >>
rlabel locali s 288 191 354 265 6 D
port 1 nsew signal input
rlabel locali s 1157 178 1271 277 6 Q
port 2 nsew signal output
rlabel locali s 1155 277 1271 282 6 Q
port 2 nsew signal output
rlabel locali s 1154 173 1271 178 6 Q
port 2 nsew signal output
rlabel locali s 1153 282 1271 283 6 Q
port 2 nsew signal output
rlabel locali s 1152 283 1271 285 6 Q
port 2 nsew signal output
rlabel locali s 1151 300 1185 375 6 Q
port 2 nsew signal output
rlabel locali s 1151 285 1271 300 6 Q
port 2 nsew signal output
rlabel locali s 1151 153 1271 173 6 Q
port 2 nsew signal output
rlabel locali s 1151 97 1185 153 6 Q
port 2 nsew signal output
rlabel locali s 1131 375 1185 493 6 Q
port 2 nsew signal output
rlabel locali s 1119 51 1185 97 6 Q
port 2 nsew signal output
rlabel locali s 896 207 1048 265 6 RESET_B
port 3 nsew signal input
rlabel locali s 896 199 963 207 6 RESET_B
port 3 nsew signal input
rlabel locali s 18 197 66 325 6 GATE
port 4 nsew clock input
rlabel metal1 s 0 -48 1288 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1326 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1288 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
