magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -3615 -1960 3615 1960
<< nwell >>
rect -2355 -700 2355 700
<< pmoshvt >>
rect -2261 -600 -1861 600
rect -1803 -600 -1403 600
rect -1345 -600 -945 600
rect -887 -600 -487 600
rect -429 -600 -29 600
rect 29 -600 429 600
rect 487 -600 887 600
rect 945 -600 1345 600
rect 1403 -600 1803 600
rect 1861 -600 2261 600
<< pdiff >>
rect -2319 561 -2261 600
rect -2319 527 -2307 561
rect -2273 527 -2261 561
rect -2319 493 -2261 527
rect -2319 459 -2307 493
rect -2273 459 -2261 493
rect -2319 425 -2261 459
rect -2319 391 -2307 425
rect -2273 391 -2261 425
rect -2319 357 -2261 391
rect -2319 323 -2307 357
rect -2273 323 -2261 357
rect -2319 289 -2261 323
rect -2319 255 -2307 289
rect -2273 255 -2261 289
rect -2319 221 -2261 255
rect -2319 187 -2307 221
rect -2273 187 -2261 221
rect -2319 153 -2261 187
rect -2319 119 -2307 153
rect -2273 119 -2261 153
rect -2319 85 -2261 119
rect -2319 51 -2307 85
rect -2273 51 -2261 85
rect -2319 17 -2261 51
rect -2319 -17 -2307 17
rect -2273 -17 -2261 17
rect -2319 -51 -2261 -17
rect -2319 -85 -2307 -51
rect -2273 -85 -2261 -51
rect -2319 -119 -2261 -85
rect -2319 -153 -2307 -119
rect -2273 -153 -2261 -119
rect -2319 -187 -2261 -153
rect -2319 -221 -2307 -187
rect -2273 -221 -2261 -187
rect -2319 -255 -2261 -221
rect -2319 -289 -2307 -255
rect -2273 -289 -2261 -255
rect -2319 -323 -2261 -289
rect -2319 -357 -2307 -323
rect -2273 -357 -2261 -323
rect -2319 -391 -2261 -357
rect -2319 -425 -2307 -391
rect -2273 -425 -2261 -391
rect -2319 -459 -2261 -425
rect -2319 -493 -2307 -459
rect -2273 -493 -2261 -459
rect -2319 -527 -2261 -493
rect -2319 -561 -2307 -527
rect -2273 -561 -2261 -527
rect -2319 -600 -2261 -561
rect -1861 561 -1803 600
rect -1861 527 -1849 561
rect -1815 527 -1803 561
rect -1861 493 -1803 527
rect -1861 459 -1849 493
rect -1815 459 -1803 493
rect -1861 425 -1803 459
rect -1861 391 -1849 425
rect -1815 391 -1803 425
rect -1861 357 -1803 391
rect -1861 323 -1849 357
rect -1815 323 -1803 357
rect -1861 289 -1803 323
rect -1861 255 -1849 289
rect -1815 255 -1803 289
rect -1861 221 -1803 255
rect -1861 187 -1849 221
rect -1815 187 -1803 221
rect -1861 153 -1803 187
rect -1861 119 -1849 153
rect -1815 119 -1803 153
rect -1861 85 -1803 119
rect -1861 51 -1849 85
rect -1815 51 -1803 85
rect -1861 17 -1803 51
rect -1861 -17 -1849 17
rect -1815 -17 -1803 17
rect -1861 -51 -1803 -17
rect -1861 -85 -1849 -51
rect -1815 -85 -1803 -51
rect -1861 -119 -1803 -85
rect -1861 -153 -1849 -119
rect -1815 -153 -1803 -119
rect -1861 -187 -1803 -153
rect -1861 -221 -1849 -187
rect -1815 -221 -1803 -187
rect -1861 -255 -1803 -221
rect -1861 -289 -1849 -255
rect -1815 -289 -1803 -255
rect -1861 -323 -1803 -289
rect -1861 -357 -1849 -323
rect -1815 -357 -1803 -323
rect -1861 -391 -1803 -357
rect -1861 -425 -1849 -391
rect -1815 -425 -1803 -391
rect -1861 -459 -1803 -425
rect -1861 -493 -1849 -459
rect -1815 -493 -1803 -459
rect -1861 -527 -1803 -493
rect -1861 -561 -1849 -527
rect -1815 -561 -1803 -527
rect -1861 -600 -1803 -561
rect -1403 561 -1345 600
rect -1403 527 -1391 561
rect -1357 527 -1345 561
rect -1403 493 -1345 527
rect -1403 459 -1391 493
rect -1357 459 -1345 493
rect -1403 425 -1345 459
rect -1403 391 -1391 425
rect -1357 391 -1345 425
rect -1403 357 -1345 391
rect -1403 323 -1391 357
rect -1357 323 -1345 357
rect -1403 289 -1345 323
rect -1403 255 -1391 289
rect -1357 255 -1345 289
rect -1403 221 -1345 255
rect -1403 187 -1391 221
rect -1357 187 -1345 221
rect -1403 153 -1345 187
rect -1403 119 -1391 153
rect -1357 119 -1345 153
rect -1403 85 -1345 119
rect -1403 51 -1391 85
rect -1357 51 -1345 85
rect -1403 17 -1345 51
rect -1403 -17 -1391 17
rect -1357 -17 -1345 17
rect -1403 -51 -1345 -17
rect -1403 -85 -1391 -51
rect -1357 -85 -1345 -51
rect -1403 -119 -1345 -85
rect -1403 -153 -1391 -119
rect -1357 -153 -1345 -119
rect -1403 -187 -1345 -153
rect -1403 -221 -1391 -187
rect -1357 -221 -1345 -187
rect -1403 -255 -1345 -221
rect -1403 -289 -1391 -255
rect -1357 -289 -1345 -255
rect -1403 -323 -1345 -289
rect -1403 -357 -1391 -323
rect -1357 -357 -1345 -323
rect -1403 -391 -1345 -357
rect -1403 -425 -1391 -391
rect -1357 -425 -1345 -391
rect -1403 -459 -1345 -425
rect -1403 -493 -1391 -459
rect -1357 -493 -1345 -459
rect -1403 -527 -1345 -493
rect -1403 -561 -1391 -527
rect -1357 -561 -1345 -527
rect -1403 -600 -1345 -561
rect -945 561 -887 600
rect -945 527 -933 561
rect -899 527 -887 561
rect -945 493 -887 527
rect -945 459 -933 493
rect -899 459 -887 493
rect -945 425 -887 459
rect -945 391 -933 425
rect -899 391 -887 425
rect -945 357 -887 391
rect -945 323 -933 357
rect -899 323 -887 357
rect -945 289 -887 323
rect -945 255 -933 289
rect -899 255 -887 289
rect -945 221 -887 255
rect -945 187 -933 221
rect -899 187 -887 221
rect -945 153 -887 187
rect -945 119 -933 153
rect -899 119 -887 153
rect -945 85 -887 119
rect -945 51 -933 85
rect -899 51 -887 85
rect -945 17 -887 51
rect -945 -17 -933 17
rect -899 -17 -887 17
rect -945 -51 -887 -17
rect -945 -85 -933 -51
rect -899 -85 -887 -51
rect -945 -119 -887 -85
rect -945 -153 -933 -119
rect -899 -153 -887 -119
rect -945 -187 -887 -153
rect -945 -221 -933 -187
rect -899 -221 -887 -187
rect -945 -255 -887 -221
rect -945 -289 -933 -255
rect -899 -289 -887 -255
rect -945 -323 -887 -289
rect -945 -357 -933 -323
rect -899 -357 -887 -323
rect -945 -391 -887 -357
rect -945 -425 -933 -391
rect -899 -425 -887 -391
rect -945 -459 -887 -425
rect -945 -493 -933 -459
rect -899 -493 -887 -459
rect -945 -527 -887 -493
rect -945 -561 -933 -527
rect -899 -561 -887 -527
rect -945 -600 -887 -561
rect -487 561 -429 600
rect -487 527 -475 561
rect -441 527 -429 561
rect -487 493 -429 527
rect -487 459 -475 493
rect -441 459 -429 493
rect -487 425 -429 459
rect -487 391 -475 425
rect -441 391 -429 425
rect -487 357 -429 391
rect -487 323 -475 357
rect -441 323 -429 357
rect -487 289 -429 323
rect -487 255 -475 289
rect -441 255 -429 289
rect -487 221 -429 255
rect -487 187 -475 221
rect -441 187 -429 221
rect -487 153 -429 187
rect -487 119 -475 153
rect -441 119 -429 153
rect -487 85 -429 119
rect -487 51 -475 85
rect -441 51 -429 85
rect -487 17 -429 51
rect -487 -17 -475 17
rect -441 -17 -429 17
rect -487 -51 -429 -17
rect -487 -85 -475 -51
rect -441 -85 -429 -51
rect -487 -119 -429 -85
rect -487 -153 -475 -119
rect -441 -153 -429 -119
rect -487 -187 -429 -153
rect -487 -221 -475 -187
rect -441 -221 -429 -187
rect -487 -255 -429 -221
rect -487 -289 -475 -255
rect -441 -289 -429 -255
rect -487 -323 -429 -289
rect -487 -357 -475 -323
rect -441 -357 -429 -323
rect -487 -391 -429 -357
rect -487 -425 -475 -391
rect -441 -425 -429 -391
rect -487 -459 -429 -425
rect -487 -493 -475 -459
rect -441 -493 -429 -459
rect -487 -527 -429 -493
rect -487 -561 -475 -527
rect -441 -561 -429 -527
rect -487 -600 -429 -561
rect -29 561 29 600
rect -29 527 -17 561
rect 17 527 29 561
rect -29 493 29 527
rect -29 459 -17 493
rect 17 459 29 493
rect -29 425 29 459
rect -29 391 -17 425
rect 17 391 29 425
rect -29 357 29 391
rect -29 323 -17 357
rect 17 323 29 357
rect -29 289 29 323
rect -29 255 -17 289
rect 17 255 29 289
rect -29 221 29 255
rect -29 187 -17 221
rect 17 187 29 221
rect -29 153 29 187
rect -29 119 -17 153
rect 17 119 29 153
rect -29 85 29 119
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -119 29 -85
rect -29 -153 -17 -119
rect 17 -153 29 -119
rect -29 -187 29 -153
rect -29 -221 -17 -187
rect 17 -221 29 -187
rect -29 -255 29 -221
rect -29 -289 -17 -255
rect 17 -289 29 -255
rect -29 -323 29 -289
rect -29 -357 -17 -323
rect 17 -357 29 -323
rect -29 -391 29 -357
rect -29 -425 -17 -391
rect 17 -425 29 -391
rect -29 -459 29 -425
rect -29 -493 -17 -459
rect 17 -493 29 -459
rect -29 -527 29 -493
rect -29 -561 -17 -527
rect 17 -561 29 -527
rect -29 -600 29 -561
rect 429 561 487 600
rect 429 527 441 561
rect 475 527 487 561
rect 429 493 487 527
rect 429 459 441 493
rect 475 459 487 493
rect 429 425 487 459
rect 429 391 441 425
rect 475 391 487 425
rect 429 357 487 391
rect 429 323 441 357
rect 475 323 487 357
rect 429 289 487 323
rect 429 255 441 289
rect 475 255 487 289
rect 429 221 487 255
rect 429 187 441 221
rect 475 187 487 221
rect 429 153 487 187
rect 429 119 441 153
rect 475 119 487 153
rect 429 85 487 119
rect 429 51 441 85
rect 475 51 487 85
rect 429 17 487 51
rect 429 -17 441 17
rect 475 -17 487 17
rect 429 -51 487 -17
rect 429 -85 441 -51
rect 475 -85 487 -51
rect 429 -119 487 -85
rect 429 -153 441 -119
rect 475 -153 487 -119
rect 429 -187 487 -153
rect 429 -221 441 -187
rect 475 -221 487 -187
rect 429 -255 487 -221
rect 429 -289 441 -255
rect 475 -289 487 -255
rect 429 -323 487 -289
rect 429 -357 441 -323
rect 475 -357 487 -323
rect 429 -391 487 -357
rect 429 -425 441 -391
rect 475 -425 487 -391
rect 429 -459 487 -425
rect 429 -493 441 -459
rect 475 -493 487 -459
rect 429 -527 487 -493
rect 429 -561 441 -527
rect 475 -561 487 -527
rect 429 -600 487 -561
rect 887 561 945 600
rect 887 527 899 561
rect 933 527 945 561
rect 887 493 945 527
rect 887 459 899 493
rect 933 459 945 493
rect 887 425 945 459
rect 887 391 899 425
rect 933 391 945 425
rect 887 357 945 391
rect 887 323 899 357
rect 933 323 945 357
rect 887 289 945 323
rect 887 255 899 289
rect 933 255 945 289
rect 887 221 945 255
rect 887 187 899 221
rect 933 187 945 221
rect 887 153 945 187
rect 887 119 899 153
rect 933 119 945 153
rect 887 85 945 119
rect 887 51 899 85
rect 933 51 945 85
rect 887 17 945 51
rect 887 -17 899 17
rect 933 -17 945 17
rect 887 -51 945 -17
rect 887 -85 899 -51
rect 933 -85 945 -51
rect 887 -119 945 -85
rect 887 -153 899 -119
rect 933 -153 945 -119
rect 887 -187 945 -153
rect 887 -221 899 -187
rect 933 -221 945 -187
rect 887 -255 945 -221
rect 887 -289 899 -255
rect 933 -289 945 -255
rect 887 -323 945 -289
rect 887 -357 899 -323
rect 933 -357 945 -323
rect 887 -391 945 -357
rect 887 -425 899 -391
rect 933 -425 945 -391
rect 887 -459 945 -425
rect 887 -493 899 -459
rect 933 -493 945 -459
rect 887 -527 945 -493
rect 887 -561 899 -527
rect 933 -561 945 -527
rect 887 -600 945 -561
rect 1345 561 1403 600
rect 1345 527 1357 561
rect 1391 527 1403 561
rect 1345 493 1403 527
rect 1345 459 1357 493
rect 1391 459 1403 493
rect 1345 425 1403 459
rect 1345 391 1357 425
rect 1391 391 1403 425
rect 1345 357 1403 391
rect 1345 323 1357 357
rect 1391 323 1403 357
rect 1345 289 1403 323
rect 1345 255 1357 289
rect 1391 255 1403 289
rect 1345 221 1403 255
rect 1345 187 1357 221
rect 1391 187 1403 221
rect 1345 153 1403 187
rect 1345 119 1357 153
rect 1391 119 1403 153
rect 1345 85 1403 119
rect 1345 51 1357 85
rect 1391 51 1403 85
rect 1345 17 1403 51
rect 1345 -17 1357 17
rect 1391 -17 1403 17
rect 1345 -51 1403 -17
rect 1345 -85 1357 -51
rect 1391 -85 1403 -51
rect 1345 -119 1403 -85
rect 1345 -153 1357 -119
rect 1391 -153 1403 -119
rect 1345 -187 1403 -153
rect 1345 -221 1357 -187
rect 1391 -221 1403 -187
rect 1345 -255 1403 -221
rect 1345 -289 1357 -255
rect 1391 -289 1403 -255
rect 1345 -323 1403 -289
rect 1345 -357 1357 -323
rect 1391 -357 1403 -323
rect 1345 -391 1403 -357
rect 1345 -425 1357 -391
rect 1391 -425 1403 -391
rect 1345 -459 1403 -425
rect 1345 -493 1357 -459
rect 1391 -493 1403 -459
rect 1345 -527 1403 -493
rect 1345 -561 1357 -527
rect 1391 -561 1403 -527
rect 1345 -600 1403 -561
rect 1803 561 1861 600
rect 1803 527 1815 561
rect 1849 527 1861 561
rect 1803 493 1861 527
rect 1803 459 1815 493
rect 1849 459 1861 493
rect 1803 425 1861 459
rect 1803 391 1815 425
rect 1849 391 1861 425
rect 1803 357 1861 391
rect 1803 323 1815 357
rect 1849 323 1861 357
rect 1803 289 1861 323
rect 1803 255 1815 289
rect 1849 255 1861 289
rect 1803 221 1861 255
rect 1803 187 1815 221
rect 1849 187 1861 221
rect 1803 153 1861 187
rect 1803 119 1815 153
rect 1849 119 1861 153
rect 1803 85 1861 119
rect 1803 51 1815 85
rect 1849 51 1861 85
rect 1803 17 1861 51
rect 1803 -17 1815 17
rect 1849 -17 1861 17
rect 1803 -51 1861 -17
rect 1803 -85 1815 -51
rect 1849 -85 1861 -51
rect 1803 -119 1861 -85
rect 1803 -153 1815 -119
rect 1849 -153 1861 -119
rect 1803 -187 1861 -153
rect 1803 -221 1815 -187
rect 1849 -221 1861 -187
rect 1803 -255 1861 -221
rect 1803 -289 1815 -255
rect 1849 -289 1861 -255
rect 1803 -323 1861 -289
rect 1803 -357 1815 -323
rect 1849 -357 1861 -323
rect 1803 -391 1861 -357
rect 1803 -425 1815 -391
rect 1849 -425 1861 -391
rect 1803 -459 1861 -425
rect 1803 -493 1815 -459
rect 1849 -493 1861 -459
rect 1803 -527 1861 -493
rect 1803 -561 1815 -527
rect 1849 -561 1861 -527
rect 1803 -600 1861 -561
rect 2261 561 2319 600
rect 2261 527 2273 561
rect 2307 527 2319 561
rect 2261 493 2319 527
rect 2261 459 2273 493
rect 2307 459 2319 493
rect 2261 425 2319 459
rect 2261 391 2273 425
rect 2307 391 2319 425
rect 2261 357 2319 391
rect 2261 323 2273 357
rect 2307 323 2319 357
rect 2261 289 2319 323
rect 2261 255 2273 289
rect 2307 255 2319 289
rect 2261 221 2319 255
rect 2261 187 2273 221
rect 2307 187 2319 221
rect 2261 153 2319 187
rect 2261 119 2273 153
rect 2307 119 2319 153
rect 2261 85 2319 119
rect 2261 51 2273 85
rect 2307 51 2319 85
rect 2261 17 2319 51
rect 2261 -17 2273 17
rect 2307 -17 2319 17
rect 2261 -51 2319 -17
rect 2261 -85 2273 -51
rect 2307 -85 2319 -51
rect 2261 -119 2319 -85
rect 2261 -153 2273 -119
rect 2307 -153 2319 -119
rect 2261 -187 2319 -153
rect 2261 -221 2273 -187
rect 2307 -221 2319 -187
rect 2261 -255 2319 -221
rect 2261 -289 2273 -255
rect 2307 -289 2319 -255
rect 2261 -323 2319 -289
rect 2261 -357 2273 -323
rect 2307 -357 2319 -323
rect 2261 -391 2319 -357
rect 2261 -425 2273 -391
rect 2307 -425 2319 -391
rect 2261 -459 2319 -425
rect 2261 -493 2273 -459
rect 2307 -493 2319 -459
rect 2261 -527 2319 -493
rect 2261 -561 2273 -527
rect 2307 -561 2319 -527
rect 2261 -600 2319 -561
<< pdiffc >>
rect -2307 527 -2273 561
rect -2307 459 -2273 493
rect -2307 391 -2273 425
rect -2307 323 -2273 357
rect -2307 255 -2273 289
rect -2307 187 -2273 221
rect -2307 119 -2273 153
rect -2307 51 -2273 85
rect -2307 -17 -2273 17
rect -2307 -85 -2273 -51
rect -2307 -153 -2273 -119
rect -2307 -221 -2273 -187
rect -2307 -289 -2273 -255
rect -2307 -357 -2273 -323
rect -2307 -425 -2273 -391
rect -2307 -493 -2273 -459
rect -2307 -561 -2273 -527
rect -1849 527 -1815 561
rect -1849 459 -1815 493
rect -1849 391 -1815 425
rect -1849 323 -1815 357
rect -1849 255 -1815 289
rect -1849 187 -1815 221
rect -1849 119 -1815 153
rect -1849 51 -1815 85
rect -1849 -17 -1815 17
rect -1849 -85 -1815 -51
rect -1849 -153 -1815 -119
rect -1849 -221 -1815 -187
rect -1849 -289 -1815 -255
rect -1849 -357 -1815 -323
rect -1849 -425 -1815 -391
rect -1849 -493 -1815 -459
rect -1849 -561 -1815 -527
rect -1391 527 -1357 561
rect -1391 459 -1357 493
rect -1391 391 -1357 425
rect -1391 323 -1357 357
rect -1391 255 -1357 289
rect -1391 187 -1357 221
rect -1391 119 -1357 153
rect -1391 51 -1357 85
rect -1391 -17 -1357 17
rect -1391 -85 -1357 -51
rect -1391 -153 -1357 -119
rect -1391 -221 -1357 -187
rect -1391 -289 -1357 -255
rect -1391 -357 -1357 -323
rect -1391 -425 -1357 -391
rect -1391 -493 -1357 -459
rect -1391 -561 -1357 -527
rect -933 527 -899 561
rect -933 459 -899 493
rect -933 391 -899 425
rect -933 323 -899 357
rect -933 255 -899 289
rect -933 187 -899 221
rect -933 119 -899 153
rect -933 51 -899 85
rect -933 -17 -899 17
rect -933 -85 -899 -51
rect -933 -153 -899 -119
rect -933 -221 -899 -187
rect -933 -289 -899 -255
rect -933 -357 -899 -323
rect -933 -425 -899 -391
rect -933 -493 -899 -459
rect -933 -561 -899 -527
rect -475 527 -441 561
rect -475 459 -441 493
rect -475 391 -441 425
rect -475 323 -441 357
rect -475 255 -441 289
rect -475 187 -441 221
rect -475 119 -441 153
rect -475 51 -441 85
rect -475 -17 -441 17
rect -475 -85 -441 -51
rect -475 -153 -441 -119
rect -475 -221 -441 -187
rect -475 -289 -441 -255
rect -475 -357 -441 -323
rect -475 -425 -441 -391
rect -475 -493 -441 -459
rect -475 -561 -441 -527
rect -17 527 17 561
rect -17 459 17 493
rect -17 391 17 425
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect -17 -425 17 -391
rect -17 -493 17 -459
rect -17 -561 17 -527
rect 441 527 475 561
rect 441 459 475 493
rect 441 391 475 425
rect 441 323 475 357
rect 441 255 475 289
rect 441 187 475 221
rect 441 119 475 153
rect 441 51 475 85
rect 441 -17 475 17
rect 441 -85 475 -51
rect 441 -153 475 -119
rect 441 -221 475 -187
rect 441 -289 475 -255
rect 441 -357 475 -323
rect 441 -425 475 -391
rect 441 -493 475 -459
rect 441 -561 475 -527
rect 899 527 933 561
rect 899 459 933 493
rect 899 391 933 425
rect 899 323 933 357
rect 899 255 933 289
rect 899 187 933 221
rect 899 119 933 153
rect 899 51 933 85
rect 899 -17 933 17
rect 899 -85 933 -51
rect 899 -153 933 -119
rect 899 -221 933 -187
rect 899 -289 933 -255
rect 899 -357 933 -323
rect 899 -425 933 -391
rect 899 -493 933 -459
rect 899 -561 933 -527
rect 1357 527 1391 561
rect 1357 459 1391 493
rect 1357 391 1391 425
rect 1357 323 1391 357
rect 1357 255 1391 289
rect 1357 187 1391 221
rect 1357 119 1391 153
rect 1357 51 1391 85
rect 1357 -17 1391 17
rect 1357 -85 1391 -51
rect 1357 -153 1391 -119
rect 1357 -221 1391 -187
rect 1357 -289 1391 -255
rect 1357 -357 1391 -323
rect 1357 -425 1391 -391
rect 1357 -493 1391 -459
rect 1357 -561 1391 -527
rect 1815 527 1849 561
rect 1815 459 1849 493
rect 1815 391 1849 425
rect 1815 323 1849 357
rect 1815 255 1849 289
rect 1815 187 1849 221
rect 1815 119 1849 153
rect 1815 51 1849 85
rect 1815 -17 1849 17
rect 1815 -85 1849 -51
rect 1815 -153 1849 -119
rect 1815 -221 1849 -187
rect 1815 -289 1849 -255
rect 1815 -357 1849 -323
rect 1815 -425 1849 -391
rect 1815 -493 1849 -459
rect 1815 -561 1849 -527
rect 2273 527 2307 561
rect 2273 459 2307 493
rect 2273 391 2307 425
rect 2273 323 2307 357
rect 2273 255 2307 289
rect 2273 187 2307 221
rect 2273 119 2307 153
rect 2273 51 2307 85
rect 2273 -17 2307 17
rect 2273 -85 2307 -51
rect 2273 -153 2307 -119
rect 2273 -221 2307 -187
rect 2273 -289 2307 -255
rect 2273 -357 2307 -323
rect 2273 -425 2307 -391
rect 2273 -493 2307 -459
rect 2273 -561 2307 -527
<< poly >>
rect -2187 681 -1935 697
rect -2187 664 -2146 681
rect -2261 647 -2146 664
rect -2112 647 -2078 681
rect -2044 647 -2010 681
rect -1976 664 -1935 681
rect -1729 681 -1477 697
rect -1729 664 -1688 681
rect -1976 647 -1861 664
rect -2261 600 -1861 647
rect -1803 647 -1688 664
rect -1654 647 -1620 681
rect -1586 647 -1552 681
rect -1518 664 -1477 681
rect -1271 681 -1019 697
rect -1271 664 -1230 681
rect -1518 647 -1403 664
rect -1803 600 -1403 647
rect -1345 647 -1230 664
rect -1196 647 -1162 681
rect -1128 647 -1094 681
rect -1060 664 -1019 681
rect -813 681 -561 697
rect -813 664 -772 681
rect -1060 647 -945 664
rect -1345 600 -945 647
rect -887 647 -772 664
rect -738 647 -704 681
rect -670 647 -636 681
rect -602 664 -561 681
rect -355 681 -103 697
rect -355 664 -314 681
rect -602 647 -487 664
rect -887 600 -487 647
rect -429 647 -314 664
rect -280 647 -246 681
rect -212 647 -178 681
rect -144 664 -103 681
rect 103 681 355 697
rect 103 664 144 681
rect -144 647 -29 664
rect -429 600 -29 647
rect 29 647 144 664
rect 178 647 212 681
rect 246 647 280 681
rect 314 664 355 681
rect 561 681 813 697
rect 561 664 602 681
rect 314 647 429 664
rect 29 600 429 647
rect 487 647 602 664
rect 636 647 670 681
rect 704 647 738 681
rect 772 664 813 681
rect 1019 681 1271 697
rect 1019 664 1060 681
rect 772 647 887 664
rect 487 600 887 647
rect 945 647 1060 664
rect 1094 647 1128 681
rect 1162 647 1196 681
rect 1230 664 1271 681
rect 1477 681 1729 697
rect 1477 664 1518 681
rect 1230 647 1345 664
rect 945 600 1345 647
rect 1403 647 1518 664
rect 1552 647 1586 681
rect 1620 647 1654 681
rect 1688 664 1729 681
rect 1935 681 2187 697
rect 1935 664 1976 681
rect 1688 647 1803 664
rect 1403 600 1803 647
rect 1861 647 1976 664
rect 2010 647 2044 681
rect 2078 647 2112 681
rect 2146 664 2187 681
rect 2146 647 2261 664
rect 1861 600 2261 647
rect -2261 -647 -1861 -600
rect -2261 -664 -2146 -647
rect -2187 -681 -2146 -664
rect -2112 -681 -2078 -647
rect -2044 -681 -2010 -647
rect -1976 -664 -1861 -647
rect -1803 -647 -1403 -600
rect -1803 -664 -1688 -647
rect -1976 -681 -1935 -664
rect -2187 -697 -1935 -681
rect -1729 -681 -1688 -664
rect -1654 -681 -1620 -647
rect -1586 -681 -1552 -647
rect -1518 -664 -1403 -647
rect -1345 -647 -945 -600
rect -1345 -664 -1230 -647
rect -1518 -681 -1477 -664
rect -1729 -697 -1477 -681
rect -1271 -681 -1230 -664
rect -1196 -681 -1162 -647
rect -1128 -681 -1094 -647
rect -1060 -664 -945 -647
rect -887 -647 -487 -600
rect -887 -664 -772 -647
rect -1060 -681 -1019 -664
rect -1271 -697 -1019 -681
rect -813 -681 -772 -664
rect -738 -681 -704 -647
rect -670 -681 -636 -647
rect -602 -664 -487 -647
rect -429 -647 -29 -600
rect -429 -664 -314 -647
rect -602 -681 -561 -664
rect -813 -697 -561 -681
rect -355 -681 -314 -664
rect -280 -681 -246 -647
rect -212 -681 -178 -647
rect -144 -664 -29 -647
rect 29 -647 429 -600
rect 29 -664 144 -647
rect -144 -681 -103 -664
rect -355 -697 -103 -681
rect 103 -681 144 -664
rect 178 -681 212 -647
rect 246 -681 280 -647
rect 314 -664 429 -647
rect 487 -647 887 -600
rect 487 -664 602 -647
rect 314 -681 355 -664
rect 103 -697 355 -681
rect 561 -681 602 -664
rect 636 -681 670 -647
rect 704 -681 738 -647
rect 772 -664 887 -647
rect 945 -647 1345 -600
rect 945 -664 1060 -647
rect 772 -681 813 -664
rect 561 -697 813 -681
rect 1019 -681 1060 -664
rect 1094 -681 1128 -647
rect 1162 -681 1196 -647
rect 1230 -664 1345 -647
rect 1403 -647 1803 -600
rect 1403 -664 1518 -647
rect 1230 -681 1271 -664
rect 1019 -697 1271 -681
rect 1477 -681 1518 -664
rect 1552 -681 1586 -647
rect 1620 -681 1654 -647
rect 1688 -664 1803 -647
rect 1861 -647 2261 -600
rect 1861 -664 1976 -647
rect 1688 -681 1729 -664
rect 1477 -697 1729 -681
rect 1935 -681 1976 -664
rect 2010 -681 2044 -647
rect 2078 -681 2112 -647
rect 2146 -664 2261 -647
rect 2146 -681 2187 -664
rect 1935 -697 2187 -681
<< polycont >>
rect -2146 647 -2112 681
rect -2078 647 -2044 681
rect -2010 647 -1976 681
rect -1688 647 -1654 681
rect -1620 647 -1586 681
rect -1552 647 -1518 681
rect -1230 647 -1196 681
rect -1162 647 -1128 681
rect -1094 647 -1060 681
rect -772 647 -738 681
rect -704 647 -670 681
rect -636 647 -602 681
rect -314 647 -280 681
rect -246 647 -212 681
rect -178 647 -144 681
rect 144 647 178 681
rect 212 647 246 681
rect 280 647 314 681
rect 602 647 636 681
rect 670 647 704 681
rect 738 647 772 681
rect 1060 647 1094 681
rect 1128 647 1162 681
rect 1196 647 1230 681
rect 1518 647 1552 681
rect 1586 647 1620 681
rect 1654 647 1688 681
rect 1976 647 2010 681
rect 2044 647 2078 681
rect 2112 647 2146 681
rect -2146 -681 -2112 -647
rect -2078 -681 -2044 -647
rect -2010 -681 -1976 -647
rect -1688 -681 -1654 -647
rect -1620 -681 -1586 -647
rect -1552 -681 -1518 -647
rect -1230 -681 -1196 -647
rect -1162 -681 -1128 -647
rect -1094 -681 -1060 -647
rect -772 -681 -738 -647
rect -704 -681 -670 -647
rect -636 -681 -602 -647
rect -314 -681 -280 -647
rect -246 -681 -212 -647
rect -178 -681 -144 -647
rect 144 -681 178 -647
rect 212 -681 246 -647
rect 280 -681 314 -647
rect 602 -681 636 -647
rect 670 -681 704 -647
rect 738 -681 772 -647
rect 1060 -681 1094 -647
rect 1128 -681 1162 -647
rect 1196 -681 1230 -647
rect 1518 -681 1552 -647
rect 1586 -681 1620 -647
rect 1654 -681 1688 -647
rect 1976 -681 2010 -647
rect 2044 -681 2078 -647
rect 2112 -681 2146 -647
<< locali >>
rect -2187 647 -2150 681
rect -2112 647 -2078 681
rect -2044 647 -2010 681
rect -1972 647 -1935 681
rect -1729 647 -1692 681
rect -1654 647 -1620 681
rect -1586 647 -1552 681
rect -1514 647 -1477 681
rect -1271 647 -1234 681
rect -1196 647 -1162 681
rect -1128 647 -1094 681
rect -1056 647 -1019 681
rect -813 647 -776 681
rect -738 647 -704 681
rect -670 647 -636 681
rect -598 647 -561 681
rect -355 647 -318 681
rect -280 647 -246 681
rect -212 647 -178 681
rect -140 647 -103 681
rect 103 647 140 681
rect 178 647 212 681
rect 246 647 280 681
rect 318 647 355 681
rect 561 647 598 681
rect 636 647 670 681
rect 704 647 738 681
rect 776 647 813 681
rect 1019 647 1056 681
rect 1094 647 1128 681
rect 1162 647 1196 681
rect 1234 647 1271 681
rect 1477 647 1514 681
rect 1552 647 1586 681
rect 1620 647 1654 681
rect 1692 647 1729 681
rect 1935 647 1972 681
rect 2010 647 2044 681
rect 2078 647 2112 681
rect 2150 647 2187 681
rect -2307 561 -2273 604
rect -2307 493 -2273 523
rect -2307 425 -2273 451
rect -2307 357 -2273 379
rect -2307 289 -2273 307
rect -2307 221 -2273 235
rect -2307 153 -2273 163
rect -2307 85 -2273 91
rect -2307 17 -2273 19
rect -2307 -19 -2273 -17
rect -2307 -91 -2273 -85
rect -2307 -163 -2273 -153
rect -2307 -235 -2273 -221
rect -2307 -307 -2273 -289
rect -2307 -379 -2273 -357
rect -2307 -451 -2273 -425
rect -2307 -523 -2273 -493
rect -2307 -604 -2273 -561
rect -1849 561 -1815 604
rect -1849 493 -1815 523
rect -1849 425 -1815 451
rect -1849 357 -1815 379
rect -1849 289 -1815 307
rect -1849 221 -1815 235
rect -1849 153 -1815 163
rect -1849 85 -1815 91
rect -1849 17 -1815 19
rect -1849 -19 -1815 -17
rect -1849 -91 -1815 -85
rect -1849 -163 -1815 -153
rect -1849 -235 -1815 -221
rect -1849 -307 -1815 -289
rect -1849 -379 -1815 -357
rect -1849 -451 -1815 -425
rect -1849 -523 -1815 -493
rect -1849 -604 -1815 -561
rect -1391 561 -1357 604
rect -1391 493 -1357 523
rect -1391 425 -1357 451
rect -1391 357 -1357 379
rect -1391 289 -1357 307
rect -1391 221 -1357 235
rect -1391 153 -1357 163
rect -1391 85 -1357 91
rect -1391 17 -1357 19
rect -1391 -19 -1357 -17
rect -1391 -91 -1357 -85
rect -1391 -163 -1357 -153
rect -1391 -235 -1357 -221
rect -1391 -307 -1357 -289
rect -1391 -379 -1357 -357
rect -1391 -451 -1357 -425
rect -1391 -523 -1357 -493
rect -1391 -604 -1357 -561
rect -933 561 -899 604
rect -933 493 -899 523
rect -933 425 -899 451
rect -933 357 -899 379
rect -933 289 -899 307
rect -933 221 -899 235
rect -933 153 -899 163
rect -933 85 -899 91
rect -933 17 -899 19
rect -933 -19 -899 -17
rect -933 -91 -899 -85
rect -933 -163 -899 -153
rect -933 -235 -899 -221
rect -933 -307 -899 -289
rect -933 -379 -899 -357
rect -933 -451 -899 -425
rect -933 -523 -899 -493
rect -933 -604 -899 -561
rect -475 561 -441 604
rect -475 493 -441 523
rect -475 425 -441 451
rect -475 357 -441 379
rect -475 289 -441 307
rect -475 221 -441 235
rect -475 153 -441 163
rect -475 85 -441 91
rect -475 17 -441 19
rect -475 -19 -441 -17
rect -475 -91 -441 -85
rect -475 -163 -441 -153
rect -475 -235 -441 -221
rect -475 -307 -441 -289
rect -475 -379 -441 -357
rect -475 -451 -441 -425
rect -475 -523 -441 -493
rect -475 -604 -441 -561
rect -17 561 17 604
rect -17 493 17 523
rect -17 425 17 451
rect -17 357 17 379
rect -17 289 17 307
rect -17 221 17 235
rect -17 153 17 163
rect -17 85 17 91
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -91 17 -85
rect -17 -163 17 -153
rect -17 -235 17 -221
rect -17 -307 17 -289
rect -17 -379 17 -357
rect -17 -451 17 -425
rect -17 -523 17 -493
rect -17 -604 17 -561
rect 441 561 475 604
rect 441 493 475 523
rect 441 425 475 451
rect 441 357 475 379
rect 441 289 475 307
rect 441 221 475 235
rect 441 153 475 163
rect 441 85 475 91
rect 441 17 475 19
rect 441 -19 475 -17
rect 441 -91 475 -85
rect 441 -163 475 -153
rect 441 -235 475 -221
rect 441 -307 475 -289
rect 441 -379 475 -357
rect 441 -451 475 -425
rect 441 -523 475 -493
rect 441 -604 475 -561
rect 899 561 933 604
rect 899 493 933 523
rect 899 425 933 451
rect 899 357 933 379
rect 899 289 933 307
rect 899 221 933 235
rect 899 153 933 163
rect 899 85 933 91
rect 899 17 933 19
rect 899 -19 933 -17
rect 899 -91 933 -85
rect 899 -163 933 -153
rect 899 -235 933 -221
rect 899 -307 933 -289
rect 899 -379 933 -357
rect 899 -451 933 -425
rect 899 -523 933 -493
rect 899 -604 933 -561
rect 1357 561 1391 604
rect 1357 493 1391 523
rect 1357 425 1391 451
rect 1357 357 1391 379
rect 1357 289 1391 307
rect 1357 221 1391 235
rect 1357 153 1391 163
rect 1357 85 1391 91
rect 1357 17 1391 19
rect 1357 -19 1391 -17
rect 1357 -91 1391 -85
rect 1357 -163 1391 -153
rect 1357 -235 1391 -221
rect 1357 -307 1391 -289
rect 1357 -379 1391 -357
rect 1357 -451 1391 -425
rect 1357 -523 1391 -493
rect 1357 -604 1391 -561
rect 1815 561 1849 604
rect 1815 493 1849 523
rect 1815 425 1849 451
rect 1815 357 1849 379
rect 1815 289 1849 307
rect 1815 221 1849 235
rect 1815 153 1849 163
rect 1815 85 1849 91
rect 1815 17 1849 19
rect 1815 -19 1849 -17
rect 1815 -91 1849 -85
rect 1815 -163 1849 -153
rect 1815 -235 1849 -221
rect 1815 -307 1849 -289
rect 1815 -379 1849 -357
rect 1815 -451 1849 -425
rect 1815 -523 1849 -493
rect 1815 -604 1849 -561
rect 2273 561 2307 604
rect 2273 493 2307 523
rect 2273 425 2307 451
rect 2273 357 2307 379
rect 2273 289 2307 307
rect 2273 221 2307 235
rect 2273 153 2307 163
rect 2273 85 2307 91
rect 2273 17 2307 19
rect 2273 -19 2307 -17
rect 2273 -91 2307 -85
rect 2273 -163 2307 -153
rect 2273 -235 2307 -221
rect 2273 -307 2307 -289
rect 2273 -379 2307 -357
rect 2273 -451 2307 -425
rect 2273 -523 2307 -493
rect 2273 -604 2307 -561
rect -2187 -681 -2150 -647
rect -2112 -681 -2078 -647
rect -2044 -681 -2010 -647
rect -1972 -681 -1935 -647
rect -1729 -681 -1692 -647
rect -1654 -681 -1620 -647
rect -1586 -681 -1552 -647
rect -1514 -681 -1477 -647
rect -1271 -681 -1234 -647
rect -1196 -681 -1162 -647
rect -1128 -681 -1094 -647
rect -1056 -681 -1019 -647
rect -813 -681 -776 -647
rect -738 -681 -704 -647
rect -670 -681 -636 -647
rect -598 -681 -561 -647
rect -355 -681 -318 -647
rect -280 -681 -246 -647
rect -212 -681 -178 -647
rect -140 -681 -103 -647
rect 103 -681 140 -647
rect 178 -681 212 -647
rect 246 -681 280 -647
rect 318 -681 355 -647
rect 561 -681 598 -647
rect 636 -681 670 -647
rect 704 -681 738 -647
rect 776 -681 813 -647
rect 1019 -681 1056 -647
rect 1094 -681 1128 -647
rect 1162 -681 1196 -647
rect 1234 -681 1271 -647
rect 1477 -681 1514 -647
rect 1552 -681 1586 -647
rect 1620 -681 1654 -647
rect 1692 -681 1729 -647
rect 1935 -681 1972 -647
rect 2010 -681 2044 -647
rect 2078 -681 2112 -647
rect 2150 -681 2187 -647
<< viali >>
rect -2150 647 -2146 681
rect -2146 647 -2116 681
rect -2078 647 -2044 681
rect -2006 647 -1976 681
rect -1976 647 -1972 681
rect -1692 647 -1688 681
rect -1688 647 -1658 681
rect -1620 647 -1586 681
rect -1548 647 -1518 681
rect -1518 647 -1514 681
rect -1234 647 -1230 681
rect -1230 647 -1200 681
rect -1162 647 -1128 681
rect -1090 647 -1060 681
rect -1060 647 -1056 681
rect -776 647 -772 681
rect -772 647 -742 681
rect -704 647 -670 681
rect -632 647 -602 681
rect -602 647 -598 681
rect -318 647 -314 681
rect -314 647 -284 681
rect -246 647 -212 681
rect -174 647 -144 681
rect -144 647 -140 681
rect 140 647 144 681
rect 144 647 174 681
rect 212 647 246 681
rect 284 647 314 681
rect 314 647 318 681
rect 598 647 602 681
rect 602 647 632 681
rect 670 647 704 681
rect 742 647 772 681
rect 772 647 776 681
rect 1056 647 1060 681
rect 1060 647 1090 681
rect 1128 647 1162 681
rect 1200 647 1230 681
rect 1230 647 1234 681
rect 1514 647 1518 681
rect 1518 647 1548 681
rect 1586 647 1620 681
rect 1658 647 1688 681
rect 1688 647 1692 681
rect 1972 647 1976 681
rect 1976 647 2006 681
rect 2044 647 2078 681
rect 2116 647 2146 681
rect 2146 647 2150 681
rect -2307 527 -2273 557
rect -2307 523 -2273 527
rect -2307 459 -2273 485
rect -2307 451 -2273 459
rect -2307 391 -2273 413
rect -2307 379 -2273 391
rect -2307 323 -2273 341
rect -2307 307 -2273 323
rect -2307 255 -2273 269
rect -2307 235 -2273 255
rect -2307 187 -2273 197
rect -2307 163 -2273 187
rect -2307 119 -2273 125
rect -2307 91 -2273 119
rect -2307 51 -2273 53
rect -2307 19 -2273 51
rect -2307 -51 -2273 -19
rect -2307 -53 -2273 -51
rect -2307 -119 -2273 -91
rect -2307 -125 -2273 -119
rect -2307 -187 -2273 -163
rect -2307 -197 -2273 -187
rect -2307 -255 -2273 -235
rect -2307 -269 -2273 -255
rect -2307 -323 -2273 -307
rect -2307 -341 -2273 -323
rect -2307 -391 -2273 -379
rect -2307 -413 -2273 -391
rect -2307 -459 -2273 -451
rect -2307 -485 -2273 -459
rect -2307 -527 -2273 -523
rect -2307 -557 -2273 -527
rect -1849 527 -1815 557
rect -1849 523 -1815 527
rect -1849 459 -1815 485
rect -1849 451 -1815 459
rect -1849 391 -1815 413
rect -1849 379 -1815 391
rect -1849 323 -1815 341
rect -1849 307 -1815 323
rect -1849 255 -1815 269
rect -1849 235 -1815 255
rect -1849 187 -1815 197
rect -1849 163 -1815 187
rect -1849 119 -1815 125
rect -1849 91 -1815 119
rect -1849 51 -1815 53
rect -1849 19 -1815 51
rect -1849 -51 -1815 -19
rect -1849 -53 -1815 -51
rect -1849 -119 -1815 -91
rect -1849 -125 -1815 -119
rect -1849 -187 -1815 -163
rect -1849 -197 -1815 -187
rect -1849 -255 -1815 -235
rect -1849 -269 -1815 -255
rect -1849 -323 -1815 -307
rect -1849 -341 -1815 -323
rect -1849 -391 -1815 -379
rect -1849 -413 -1815 -391
rect -1849 -459 -1815 -451
rect -1849 -485 -1815 -459
rect -1849 -527 -1815 -523
rect -1849 -557 -1815 -527
rect -1391 527 -1357 557
rect -1391 523 -1357 527
rect -1391 459 -1357 485
rect -1391 451 -1357 459
rect -1391 391 -1357 413
rect -1391 379 -1357 391
rect -1391 323 -1357 341
rect -1391 307 -1357 323
rect -1391 255 -1357 269
rect -1391 235 -1357 255
rect -1391 187 -1357 197
rect -1391 163 -1357 187
rect -1391 119 -1357 125
rect -1391 91 -1357 119
rect -1391 51 -1357 53
rect -1391 19 -1357 51
rect -1391 -51 -1357 -19
rect -1391 -53 -1357 -51
rect -1391 -119 -1357 -91
rect -1391 -125 -1357 -119
rect -1391 -187 -1357 -163
rect -1391 -197 -1357 -187
rect -1391 -255 -1357 -235
rect -1391 -269 -1357 -255
rect -1391 -323 -1357 -307
rect -1391 -341 -1357 -323
rect -1391 -391 -1357 -379
rect -1391 -413 -1357 -391
rect -1391 -459 -1357 -451
rect -1391 -485 -1357 -459
rect -1391 -527 -1357 -523
rect -1391 -557 -1357 -527
rect -933 527 -899 557
rect -933 523 -899 527
rect -933 459 -899 485
rect -933 451 -899 459
rect -933 391 -899 413
rect -933 379 -899 391
rect -933 323 -899 341
rect -933 307 -899 323
rect -933 255 -899 269
rect -933 235 -899 255
rect -933 187 -899 197
rect -933 163 -899 187
rect -933 119 -899 125
rect -933 91 -899 119
rect -933 51 -899 53
rect -933 19 -899 51
rect -933 -51 -899 -19
rect -933 -53 -899 -51
rect -933 -119 -899 -91
rect -933 -125 -899 -119
rect -933 -187 -899 -163
rect -933 -197 -899 -187
rect -933 -255 -899 -235
rect -933 -269 -899 -255
rect -933 -323 -899 -307
rect -933 -341 -899 -323
rect -933 -391 -899 -379
rect -933 -413 -899 -391
rect -933 -459 -899 -451
rect -933 -485 -899 -459
rect -933 -527 -899 -523
rect -933 -557 -899 -527
rect -475 527 -441 557
rect -475 523 -441 527
rect -475 459 -441 485
rect -475 451 -441 459
rect -475 391 -441 413
rect -475 379 -441 391
rect -475 323 -441 341
rect -475 307 -441 323
rect -475 255 -441 269
rect -475 235 -441 255
rect -475 187 -441 197
rect -475 163 -441 187
rect -475 119 -441 125
rect -475 91 -441 119
rect -475 51 -441 53
rect -475 19 -441 51
rect -475 -51 -441 -19
rect -475 -53 -441 -51
rect -475 -119 -441 -91
rect -475 -125 -441 -119
rect -475 -187 -441 -163
rect -475 -197 -441 -187
rect -475 -255 -441 -235
rect -475 -269 -441 -255
rect -475 -323 -441 -307
rect -475 -341 -441 -323
rect -475 -391 -441 -379
rect -475 -413 -441 -391
rect -475 -459 -441 -451
rect -475 -485 -441 -459
rect -475 -527 -441 -523
rect -475 -557 -441 -527
rect -17 527 17 557
rect -17 523 17 527
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect -17 -527 17 -523
rect -17 -557 17 -527
rect 441 527 475 557
rect 441 523 475 527
rect 441 459 475 485
rect 441 451 475 459
rect 441 391 475 413
rect 441 379 475 391
rect 441 323 475 341
rect 441 307 475 323
rect 441 255 475 269
rect 441 235 475 255
rect 441 187 475 197
rect 441 163 475 187
rect 441 119 475 125
rect 441 91 475 119
rect 441 51 475 53
rect 441 19 475 51
rect 441 -51 475 -19
rect 441 -53 475 -51
rect 441 -119 475 -91
rect 441 -125 475 -119
rect 441 -187 475 -163
rect 441 -197 475 -187
rect 441 -255 475 -235
rect 441 -269 475 -255
rect 441 -323 475 -307
rect 441 -341 475 -323
rect 441 -391 475 -379
rect 441 -413 475 -391
rect 441 -459 475 -451
rect 441 -485 475 -459
rect 441 -527 475 -523
rect 441 -557 475 -527
rect 899 527 933 557
rect 899 523 933 527
rect 899 459 933 485
rect 899 451 933 459
rect 899 391 933 413
rect 899 379 933 391
rect 899 323 933 341
rect 899 307 933 323
rect 899 255 933 269
rect 899 235 933 255
rect 899 187 933 197
rect 899 163 933 187
rect 899 119 933 125
rect 899 91 933 119
rect 899 51 933 53
rect 899 19 933 51
rect 899 -51 933 -19
rect 899 -53 933 -51
rect 899 -119 933 -91
rect 899 -125 933 -119
rect 899 -187 933 -163
rect 899 -197 933 -187
rect 899 -255 933 -235
rect 899 -269 933 -255
rect 899 -323 933 -307
rect 899 -341 933 -323
rect 899 -391 933 -379
rect 899 -413 933 -391
rect 899 -459 933 -451
rect 899 -485 933 -459
rect 899 -527 933 -523
rect 899 -557 933 -527
rect 1357 527 1391 557
rect 1357 523 1391 527
rect 1357 459 1391 485
rect 1357 451 1391 459
rect 1357 391 1391 413
rect 1357 379 1391 391
rect 1357 323 1391 341
rect 1357 307 1391 323
rect 1357 255 1391 269
rect 1357 235 1391 255
rect 1357 187 1391 197
rect 1357 163 1391 187
rect 1357 119 1391 125
rect 1357 91 1391 119
rect 1357 51 1391 53
rect 1357 19 1391 51
rect 1357 -51 1391 -19
rect 1357 -53 1391 -51
rect 1357 -119 1391 -91
rect 1357 -125 1391 -119
rect 1357 -187 1391 -163
rect 1357 -197 1391 -187
rect 1357 -255 1391 -235
rect 1357 -269 1391 -255
rect 1357 -323 1391 -307
rect 1357 -341 1391 -323
rect 1357 -391 1391 -379
rect 1357 -413 1391 -391
rect 1357 -459 1391 -451
rect 1357 -485 1391 -459
rect 1357 -527 1391 -523
rect 1357 -557 1391 -527
rect 1815 527 1849 557
rect 1815 523 1849 527
rect 1815 459 1849 485
rect 1815 451 1849 459
rect 1815 391 1849 413
rect 1815 379 1849 391
rect 1815 323 1849 341
rect 1815 307 1849 323
rect 1815 255 1849 269
rect 1815 235 1849 255
rect 1815 187 1849 197
rect 1815 163 1849 187
rect 1815 119 1849 125
rect 1815 91 1849 119
rect 1815 51 1849 53
rect 1815 19 1849 51
rect 1815 -51 1849 -19
rect 1815 -53 1849 -51
rect 1815 -119 1849 -91
rect 1815 -125 1849 -119
rect 1815 -187 1849 -163
rect 1815 -197 1849 -187
rect 1815 -255 1849 -235
rect 1815 -269 1849 -255
rect 1815 -323 1849 -307
rect 1815 -341 1849 -323
rect 1815 -391 1849 -379
rect 1815 -413 1849 -391
rect 1815 -459 1849 -451
rect 1815 -485 1849 -459
rect 1815 -527 1849 -523
rect 1815 -557 1849 -527
rect 2273 527 2307 557
rect 2273 523 2307 527
rect 2273 459 2307 485
rect 2273 451 2307 459
rect 2273 391 2307 413
rect 2273 379 2307 391
rect 2273 323 2307 341
rect 2273 307 2307 323
rect 2273 255 2307 269
rect 2273 235 2307 255
rect 2273 187 2307 197
rect 2273 163 2307 187
rect 2273 119 2307 125
rect 2273 91 2307 119
rect 2273 51 2307 53
rect 2273 19 2307 51
rect 2273 -51 2307 -19
rect 2273 -53 2307 -51
rect 2273 -119 2307 -91
rect 2273 -125 2307 -119
rect 2273 -187 2307 -163
rect 2273 -197 2307 -187
rect 2273 -255 2307 -235
rect 2273 -269 2307 -255
rect 2273 -323 2307 -307
rect 2273 -341 2307 -323
rect 2273 -391 2307 -379
rect 2273 -413 2307 -391
rect 2273 -459 2307 -451
rect 2273 -485 2307 -459
rect 2273 -527 2307 -523
rect 2273 -557 2307 -527
rect -2150 -681 -2146 -647
rect -2146 -681 -2116 -647
rect -2078 -681 -2044 -647
rect -2006 -681 -1976 -647
rect -1976 -681 -1972 -647
rect -1692 -681 -1688 -647
rect -1688 -681 -1658 -647
rect -1620 -681 -1586 -647
rect -1548 -681 -1518 -647
rect -1518 -681 -1514 -647
rect -1234 -681 -1230 -647
rect -1230 -681 -1200 -647
rect -1162 -681 -1128 -647
rect -1090 -681 -1060 -647
rect -1060 -681 -1056 -647
rect -776 -681 -772 -647
rect -772 -681 -742 -647
rect -704 -681 -670 -647
rect -632 -681 -602 -647
rect -602 -681 -598 -647
rect -318 -681 -314 -647
rect -314 -681 -284 -647
rect -246 -681 -212 -647
rect -174 -681 -144 -647
rect -144 -681 -140 -647
rect 140 -681 144 -647
rect 144 -681 174 -647
rect 212 -681 246 -647
rect 284 -681 314 -647
rect 314 -681 318 -647
rect 598 -681 602 -647
rect 602 -681 632 -647
rect 670 -681 704 -647
rect 742 -681 772 -647
rect 772 -681 776 -647
rect 1056 -681 1060 -647
rect 1060 -681 1090 -647
rect 1128 -681 1162 -647
rect 1200 -681 1230 -647
rect 1230 -681 1234 -647
rect 1514 -681 1518 -647
rect 1518 -681 1548 -647
rect 1586 -681 1620 -647
rect 1658 -681 1688 -647
rect 1688 -681 1692 -647
rect 1972 -681 1976 -647
rect 1976 -681 2006 -647
rect 2044 -681 2078 -647
rect 2116 -681 2146 -647
rect 2146 -681 2150 -647
<< metal1 >>
rect -2165 681 -1957 687
rect -2165 647 -2150 681
rect -2116 647 -2078 681
rect -2044 647 -2006 681
rect -1972 647 -1957 681
rect -2165 641 -1957 647
rect -1707 681 -1499 687
rect -1707 647 -1692 681
rect -1658 647 -1620 681
rect -1586 647 -1548 681
rect -1514 647 -1499 681
rect -1707 641 -1499 647
rect -1249 681 -1041 687
rect -1249 647 -1234 681
rect -1200 647 -1162 681
rect -1128 647 -1090 681
rect -1056 647 -1041 681
rect -1249 641 -1041 647
rect -791 681 -583 687
rect -791 647 -776 681
rect -742 647 -704 681
rect -670 647 -632 681
rect -598 647 -583 681
rect -791 641 -583 647
rect -333 681 -125 687
rect -333 647 -318 681
rect -284 647 -246 681
rect -212 647 -174 681
rect -140 647 -125 681
rect -333 641 -125 647
rect 125 681 333 687
rect 125 647 140 681
rect 174 647 212 681
rect 246 647 284 681
rect 318 647 333 681
rect 125 641 333 647
rect 583 681 791 687
rect 583 647 598 681
rect 632 647 670 681
rect 704 647 742 681
rect 776 647 791 681
rect 583 641 791 647
rect 1041 681 1249 687
rect 1041 647 1056 681
rect 1090 647 1128 681
rect 1162 647 1200 681
rect 1234 647 1249 681
rect 1041 641 1249 647
rect 1499 681 1707 687
rect 1499 647 1514 681
rect 1548 647 1586 681
rect 1620 647 1658 681
rect 1692 647 1707 681
rect 1499 641 1707 647
rect 1957 681 2165 687
rect 1957 647 1972 681
rect 2006 647 2044 681
rect 2078 647 2116 681
rect 2150 647 2165 681
rect 1957 641 2165 647
rect -2313 557 -2267 600
rect -2313 523 -2307 557
rect -2273 523 -2267 557
rect -2313 485 -2267 523
rect -2313 451 -2307 485
rect -2273 451 -2267 485
rect -2313 413 -2267 451
rect -2313 379 -2307 413
rect -2273 379 -2267 413
rect -2313 341 -2267 379
rect -2313 307 -2307 341
rect -2273 307 -2267 341
rect -2313 269 -2267 307
rect -2313 235 -2307 269
rect -2273 235 -2267 269
rect -2313 197 -2267 235
rect -2313 163 -2307 197
rect -2273 163 -2267 197
rect -2313 125 -2267 163
rect -2313 91 -2307 125
rect -2273 91 -2267 125
rect -2313 53 -2267 91
rect -2313 19 -2307 53
rect -2273 19 -2267 53
rect -2313 -19 -2267 19
rect -2313 -53 -2307 -19
rect -2273 -53 -2267 -19
rect -2313 -91 -2267 -53
rect -2313 -125 -2307 -91
rect -2273 -125 -2267 -91
rect -2313 -163 -2267 -125
rect -2313 -197 -2307 -163
rect -2273 -197 -2267 -163
rect -2313 -235 -2267 -197
rect -2313 -269 -2307 -235
rect -2273 -269 -2267 -235
rect -2313 -307 -2267 -269
rect -2313 -341 -2307 -307
rect -2273 -341 -2267 -307
rect -2313 -379 -2267 -341
rect -2313 -413 -2307 -379
rect -2273 -413 -2267 -379
rect -2313 -451 -2267 -413
rect -2313 -485 -2307 -451
rect -2273 -485 -2267 -451
rect -2313 -523 -2267 -485
rect -2313 -557 -2307 -523
rect -2273 -557 -2267 -523
rect -2313 -600 -2267 -557
rect -1855 557 -1809 600
rect -1855 523 -1849 557
rect -1815 523 -1809 557
rect -1855 485 -1809 523
rect -1855 451 -1849 485
rect -1815 451 -1809 485
rect -1855 413 -1809 451
rect -1855 379 -1849 413
rect -1815 379 -1809 413
rect -1855 341 -1809 379
rect -1855 307 -1849 341
rect -1815 307 -1809 341
rect -1855 269 -1809 307
rect -1855 235 -1849 269
rect -1815 235 -1809 269
rect -1855 197 -1809 235
rect -1855 163 -1849 197
rect -1815 163 -1809 197
rect -1855 125 -1809 163
rect -1855 91 -1849 125
rect -1815 91 -1809 125
rect -1855 53 -1809 91
rect -1855 19 -1849 53
rect -1815 19 -1809 53
rect -1855 -19 -1809 19
rect -1855 -53 -1849 -19
rect -1815 -53 -1809 -19
rect -1855 -91 -1809 -53
rect -1855 -125 -1849 -91
rect -1815 -125 -1809 -91
rect -1855 -163 -1809 -125
rect -1855 -197 -1849 -163
rect -1815 -197 -1809 -163
rect -1855 -235 -1809 -197
rect -1855 -269 -1849 -235
rect -1815 -269 -1809 -235
rect -1855 -307 -1809 -269
rect -1855 -341 -1849 -307
rect -1815 -341 -1809 -307
rect -1855 -379 -1809 -341
rect -1855 -413 -1849 -379
rect -1815 -413 -1809 -379
rect -1855 -451 -1809 -413
rect -1855 -485 -1849 -451
rect -1815 -485 -1809 -451
rect -1855 -523 -1809 -485
rect -1855 -557 -1849 -523
rect -1815 -557 -1809 -523
rect -1855 -600 -1809 -557
rect -1397 557 -1351 600
rect -1397 523 -1391 557
rect -1357 523 -1351 557
rect -1397 485 -1351 523
rect -1397 451 -1391 485
rect -1357 451 -1351 485
rect -1397 413 -1351 451
rect -1397 379 -1391 413
rect -1357 379 -1351 413
rect -1397 341 -1351 379
rect -1397 307 -1391 341
rect -1357 307 -1351 341
rect -1397 269 -1351 307
rect -1397 235 -1391 269
rect -1357 235 -1351 269
rect -1397 197 -1351 235
rect -1397 163 -1391 197
rect -1357 163 -1351 197
rect -1397 125 -1351 163
rect -1397 91 -1391 125
rect -1357 91 -1351 125
rect -1397 53 -1351 91
rect -1397 19 -1391 53
rect -1357 19 -1351 53
rect -1397 -19 -1351 19
rect -1397 -53 -1391 -19
rect -1357 -53 -1351 -19
rect -1397 -91 -1351 -53
rect -1397 -125 -1391 -91
rect -1357 -125 -1351 -91
rect -1397 -163 -1351 -125
rect -1397 -197 -1391 -163
rect -1357 -197 -1351 -163
rect -1397 -235 -1351 -197
rect -1397 -269 -1391 -235
rect -1357 -269 -1351 -235
rect -1397 -307 -1351 -269
rect -1397 -341 -1391 -307
rect -1357 -341 -1351 -307
rect -1397 -379 -1351 -341
rect -1397 -413 -1391 -379
rect -1357 -413 -1351 -379
rect -1397 -451 -1351 -413
rect -1397 -485 -1391 -451
rect -1357 -485 -1351 -451
rect -1397 -523 -1351 -485
rect -1397 -557 -1391 -523
rect -1357 -557 -1351 -523
rect -1397 -600 -1351 -557
rect -939 557 -893 600
rect -939 523 -933 557
rect -899 523 -893 557
rect -939 485 -893 523
rect -939 451 -933 485
rect -899 451 -893 485
rect -939 413 -893 451
rect -939 379 -933 413
rect -899 379 -893 413
rect -939 341 -893 379
rect -939 307 -933 341
rect -899 307 -893 341
rect -939 269 -893 307
rect -939 235 -933 269
rect -899 235 -893 269
rect -939 197 -893 235
rect -939 163 -933 197
rect -899 163 -893 197
rect -939 125 -893 163
rect -939 91 -933 125
rect -899 91 -893 125
rect -939 53 -893 91
rect -939 19 -933 53
rect -899 19 -893 53
rect -939 -19 -893 19
rect -939 -53 -933 -19
rect -899 -53 -893 -19
rect -939 -91 -893 -53
rect -939 -125 -933 -91
rect -899 -125 -893 -91
rect -939 -163 -893 -125
rect -939 -197 -933 -163
rect -899 -197 -893 -163
rect -939 -235 -893 -197
rect -939 -269 -933 -235
rect -899 -269 -893 -235
rect -939 -307 -893 -269
rect -939 -341 -933 -307
rect -899 -341 -893 -307
rect -939 -379 -893 -341
rect -939 -413 -933 -379
rect -899 -413 -893 -379
rect -939 -451 -893 -413
rect -939 -485 -933 -451
rect -899 -485 -893 -451
rect -939 -523 -893 -485
rect -939 -557 -933 -523
rect -899 -557 -893 -523
rect -939 -600 -893 -557
rect -481 557 -435 600
rect -481 523 -475 557
rect -441 523 -435 557
rect -481 485 -435 523
rect -481 451 -475 485
rect -441 451 -435 485
rect -481 413 -435 451
rect -481 379 -475 413
rect -441 379 -435 413
rect -481 341 -435 379
rect -481 307 -475 341
rect -441 307 -435 341
rect -481 269 -435 307
rect -481 235 -475 269
rect -441 235 -435 269
rect -481 197 -435 235
rect -481 163 -475 197
rect -441 163 -435 197
rect -481 125 -435 163
rect -481 91 -475 125
rect -441 91 -435 125
rect -481 53 -435 91
rect -481 19 -475 53
rect -441 19 -435 53
rect -481 -19 -435 19
rect -481 -53 -475 -19
rect -441 -53 -435 -19
rect -481 -91 -435 -53
rect -481 -125 -475 -91
rect -441 -125 -435 -91
rect -481 -163 -435 -125
rect -481 -197 -475 -163
rect -441 -197 -435 -163
rect -481 -235 -435 -197
rect -481 -269 -475 -235
rect -441 -269 -435 -235
rect -481 -307 -435 -269
rect -481 -341 -475 -307
rect -441 -341 -435 -307
rect -481 -379 -435 -341
rect -481 -413 -475 -379
rect -441 -413 -435 -379
rect -481 -451 -435 -413
rect -481 -485 -475 -451
rect -441 -485 -435 -451
rect -481 -523 -435 -485
rect -481 -557 -475 -523
rect -441 -557 -435 -523
rect -481 -600 -435 -557
rect -23 557 23 600
rect -23 523 -17 557
rect 17 523 23 557
rect -23 485 23 523
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -523 23 -485
rect -23 -557 -17 -523
rect 17 -557 23 -523
rect -23 -600 23 -557
rect 435 557 481 600
rect 435 523 441 557
rect 475 523 481 557
rect 435 485 481 523
rect 435 451 441 485
rect 475 451 481 485
rect 435 413 481 451
rect 435 379 441 413
rect 475 379 481 413
rect 435 341 481 379
rect 435 307 441 341
rect 475 307 481 341
rect 435 269 481 307
rect 435 235 441 269
rect 475 235 481 269
rect 435 197 481 235
rect 435 163 441 197
rect 475 163 481 197
rect 435 125 481 163
rect 435 91 441 125
rect 475 91 481 125
rect 435 53 481 91
rect 435 19 441 53
rect 475 19 481 53
rect 435 -19 481 19
rect 435 -53 441 -19
rect 475 -53 481 -19
rect 435 -91 481 -53
rect 435 -125 441 -91
rect 475 -125 481 -91
rect 435 -163 481 -125
rect 435 -197 441 -163
rect 475 -197 481 -163
rect 435 -235 481 -197
rect 435 -269 441 -235
rect 475 -269 481 -235
rect 435 -307 481 -269
rect 435 -341 441 -307
rect 475 -341 481 -307
rect 435 -379 481 -341
rect 435 -413 441 -379
rect 475 -413 481 -379
rect 435 -451 481 -413
rect 435 -485 441 -451
rect 475 -485 481 -451
rect 435 -523 481 -485
rect 435 -557 441 -523
rect 475 -557 481 -523
rect 435 -600 481 -557
rect 893 557 939 600
rect 893 523 899 557
rect 933 523 939 557
rect 893 485 939 523
rect 893 451 899 485
rect 933 451 939 485
rect 893 413 939 451
rect 893 379 899 413
rect 933 379 939 413
rect 893 341 939 379
rect 893 307 899 341
rect 933 307 939 341
rect 893 269 939 307
rect 893 235 899 269
rect 933 235 939 269
rect 893 197 939 235
rect 893 163 899 197
rect 933 163 939 197
rect 893 125 939 163
rect 893 91 899 125
rect 933 91 939 125
rect 893 53 939 91
rect 893 19 899 53
rect 933 19 939 53
rect 893 -19 939 19
rect 893 -53 899 -19
rect 933 -53 939 -19
rect 893 -91 939 -53
rect 893 -125 899 -91
rect 933 -125 939 -91
rect 893 -163 939 -125
rect 893 -197 899 -163
rect 933 -197 939 -163
rect 893 -235 939 -197
rect 893 -269 899 -235
rect 933 -269 939 -235
rect 893 -307 939 -269
rect 893 -341 899 -307
rect 933 -341 939 -307
rect 893 -379 939 -341
rect 893 -413 899 -379
rect 933 -413 939 -379
rect 893 -451 939 -413
rect 893 -485 899 -451
rect 933 -485 939 -451
rect 893 -523 939 -485
rect 893 -557 899 -523
rect 933 -557 939 -523
rect 893 -600 939 -557
rect 1351 557 1397 600
rect 1351 523 1357 557
rect 1391 523 1397 557
rect 1351 485 1397 523
rect 1351 451 1357 485
rect 1391 451 1397 485
rect 1351 413 1397 451
rect 1351 379 1357 413
rect 1391 379 1397 413
rect 1351 341 1397 379
rect 1351 307 1357 341
rect 1391 307 1397 341
rect 1351 269 1397 307
rect 1351 235 1357 269
rect 1391 235 1397 269
rect 1351 197 1397 235
rect 1351 163 1357 197
rect 1391 163 1397 197
rect 1351 125 1397 163
rect 1351 91 1357 125
rect 1391 91 1397 125
rect 1351 53 1397 91
rect 1351 19 1357 53
rect 1391 19 1397 53
rect 1351 -19 1397 19
rect 1351 -53 1357 -19
rect 1391 -53 1397 -19
rect 1351 -91 1397 -53
rect 1351 -125 1357 -91
rect 1391 -125 1397 -91
rect 1351 -163 1397 -125
rect 1351 -197 1357 -163
rect 1391 -197 1397 -163
rect 1351 -235 1397 -197
rect 1351 -269 1357 -235
rect 1391 -269 1397 -235
rect 1351 -307 1397 -269
rect 1351 -341 1357 -307
rect 1391 -341 1397 -307
rect 1351 -379 1397 -341
rect 1351 -413 1357 -379
rect 1391 -413 1397 -379
rect 1351 -451 1397 -413
rect 1351 -485 1357 -451
rect 1391 -485 1397 -451
rect 1351 -523 1397 -485
rect 1351 -557 1357 -523
rect 1391 -557 1397 -523
rect 1351 -600 1397 -557
rect 1809 557 1855 600
rect 1809 523 1815 557
rect 1849 523 1855 557
rect 1809 485 1855 523
rect 1809 451 1815 485
rect 1849 451 1855 485
rect 1809 413 1855 451
rect 1809 379 1815 413
rect 1849 379 1855 413
rect 1809 341 1855 379
rect 1809 307 1815 341
rect 1849 307 1855 341
rect 1809 269 1855 307
rect 1809 235 1815 269
rect 1849 235 1855 269
rect 1809 197 1855 235
rect 1809 163 1815 197
rect 1849 163 1855 197
rect 1809 125 1855 163
rect 1809 91 1815 125
rect 1849 91 1855 125
rect 1809 53 1855 91
rect 1809 19 1815 53
rect 1849 19 1855 53
rect 1809 -19 1855 19
rect 1809 -53 1815 -19
rect 1849 -53 1855 -19
rect 1809 -91 1855 -53
rect 1809 -125 1815 -91
rect 1849 -125 1855 -91
rect 1809 -163 1855 -125
rect 1809 -197 1815 -163
rect 1849 -197 1855 -163
rect 1809 -235 1855 -197
rect 1809 -269 1815 -235
rect 1849 -269 1855 -235
rect 1809 -307 1855 -269
rect 1809 -341 1815 -307
rect 1849 -341 1855 -307
rect 1809 -379 1855 -341
rect 1809 -413 1815 -379
rect 1849 -413 1855 -379
rect 1809 -451 1855 -413
rect 1809 -485 1815 -451
rect 1849 -485 1855 -451
rect 1809 -523 1855 -485
rect 1809 -557 1815 -523
rect 1849 -557 1855 -523
rect 1809 -600 1855 -557
rect 2267 557 2313 600
rect 2267 523 2273 557
rect 2307 523 2313 557
rect 2267 485 2313 523
rect 2267 451 2273 485
rect 2307 451 2313 485
rect 2267 413 2313 451
rect 2267 379 2273 413
rect 2307 379 2313 413
rect 2267 341 2313 379
rect 2267 307 2273 341
rect 2307 307 2313 341
rect 2267 269 2313 307
rect 2267 235 2273 269
rect 2307 235 2313 269
rect 2267 197 2313 235
rect 2267 163 2273 197
rect 2307 163 2313 197
rect 2267 125 2313 163
rect 2267 91 2273 125
rect 2307 91 2313 125
rect 2267 53 2313 91
rect 2267 19 2273 53
rect 2307 19 2313 53
rect 2267 -19 2313 19
rect 2267 -53 2273 -19
rect 2307 -53 2313 -19
rect 2267 -91 2313 -53
rect 2267 -125 2273 -91
rect 2307 -125 2313 -91
rect 2267 -163 2313 -125
rect 2267 -197 2273 -163
rect 2307 -197 2313 -163
rect 2267 -235 2313 -197
rect 2267 -269 2273 -235
rect 2307 -269 2313 -235
rect 2267 -307 2313 -269
rect 2267 -341 2273 -307
rect 2307 -341 2313 -307
rect 2267 -379 2313 -341
rect 2267 -413 2273 -379
rect 2307 -413 2313 -379
rect 2267 -451 2313 -413
rect 2267 -485 2273 -451
rect 2307 -485 2313 -451
rect 2267 -523 2313 -485
rect 2267 -557 2273 -523
rect 2307 -557 2313 -523
rect 2267 -600 2313 -557
rect -2165 -647 -1957 -641
rect -2165 -681 -2150 -647
rect -2116 -681 -2078 -647
rect -2044 -681 -2006 -647
rect -1972 -681 -1957 -647
rect -2165 -687 -1957 -681
rect -1707 -647 -1499 -641
rect -1707 -681 -1692 -647
rect -1658 -681 -1620 -647
rect -1586 -681 -1548 -647
rect -1514 -681 -1499 -647
rect -1707 -687 -1499 -681
rect -1249 -647 -1041 -641
rect -1249 -681 -1234 -647
rect -1200 -681 -1162 -647
rect -1128 -681 -1090 -647
rect -1056 -681 -1041 -647
rect -1249 -687 -1041 -681
rect -791 -647 -583 -641
rect -791 -681 -776 -647
rect -742 -681 -704 -647
rect -670 -681 -632 -647
rect -598 -681 -583 -647
rect -791 -687 -583 -681
rect -333 -647 -125 -641
rect -333 -681 -318 -647
rect -284 -681 -246 -647
rect -212 -681 -174 -647
rect -140 -681 -125 -647
rect -333 -687 -125 -681
rect 125 -647 333 -641
rect 125 -681 140 -647
rect 174 -681 212 -647
rect 246 -681 284 -647
rect 318 -681 333 -647
rect 125 -687 333 -681
rect 583 -647 791 -641
rect 583 -681 598 -647
rect 632 -681 670 -647
rect 704 -681 742 -647
rect 776 -681 791 -647
rect 583 -687 791 -681
rect 1041 -647 1249 -641
rect 1041 -681 1056 -647
rect 1090 -681 1128 -647
rect 1162 -681 1200 -647
rect 1234 -681 1249 -647
rect 1041 -687 1249 -681
rect 1499 -647 1707 -641
rect 1499 -681 1514 -647
rect 1548 -681 1586 -647
rect 1620 -681 1658 -647
rect 1692 -681 1707 -647
rect 1499 -687 1707 -681
rect 1957 -647 2165 -641
rect 1957 -681 1972 -647
rect 2006 -681 2044 -647
rect 2078 -681 2116 -647
rect 2150 -681 2165 -647
rect 1957 -687 2165 -681
<< end >>
