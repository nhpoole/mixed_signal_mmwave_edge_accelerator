magic
tech sky130A
timestamp 1625948044
<< metal3 >>
rect -61 16 61 24
rect -61 -16 -56 16
rect -24 -16 -16 16
rect 16 -16 24 16
rect 56 -16 61 16
rect -61 -24 61 -16
<< via3 >>
rect -56 -16 -24 16
rect -16 -16 16 16
rect 24 -16 56 16
<< metal4 >>
rect -61 16 61 24
rect -61 -16 -56 16
rect -24 -16 -16 16
rect 16 -16 24 16
rect 56 -16 61 16
rect -61 -24 61 -16
<< end >>
