magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -2410 -1560 2409 1560
<< metal3 >>
rect -1150 272 1149 300
rect -1150 208 1065 272
rect 1129 208 1149 272
rect -1150 192 1149 208
rect -1150 128 1065 192
rect 1129 128 1149 192
rect -1150 112 1149 128
rect -1150 48 1065 112
rect 1129 48 1149 112
rect -1150 32 1149 48
rect -1150 -32 1065 32
rect 1129 -32 1149 32
rect -1150 -48 1149 -32
rect -1150 -112 1065 -48
rect 1129 -112 1149 -48
rect -1150 -128 1149 -112
rect -1150 -192 1065 -128
rect 1129 -192 1149 -128
rect -1150 -208 1149 -192
rect -1150 -272 1065 -208
rect 1129 -272 1149 -208
rect -1150 -300 1149 -272
<< via3 >>
rect 1065 208 1129 272
rect 1065 128 1129 192
rect 1065 48 1129 112
rect 1065 -32 1129 32
rect 1065 -112 1129 -48
rect 1065 -192 1129 -128
rect 1065 -272 1129 -208
<< mimcap >>
rect -1050 152 950 200
rect -1050 -152 -1002 152
rect 902 -152 950 152
rect -1050 -200 950 -152
<< mimcapcontact >>
rect -1002 -152 902 152
<< metal4 >>
rect 1049 272 1145 288
rect 1049 208 1065 272
rect 1129 208 1145 272
rect 1049 192 1145 208
rect -1011 152 911 161
rect -1011 -152 -1002 152
rect 902 -152 911 152
rect -1011 -161 911 -152
rect 1049 128 1065 192
rect 1129 128 1145 192
rect 1049 112 1145 128
rect 1049 48 1065 112
rect 1129 48 1145 112
rect 1049 32 1145 48
rect 1049 -32 1065 32
rect 1129 -32 1145 32
rect 1049 -48 1145 -32
rect 1049 -112 1065 -48
rect 1129 -112 1145 -48
rect 1049 -128 1145 -112
rect 1049 -192 1065 -128
rect 1129 -192 1145 -128
rect 1049 -208 1145 -192
rect 1049 -272 1065 -208
rect 1129 -272 1145 -208
rect 1049 -288 1145 -272
<< properties >>
string FIXED_BBOX -1150 -300 1050 300
<< end >>
