magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1332 -1786 5948 1930
<< locali >>
rect 4104 453 4152 460
rect 4104 419 4111 453
rect 4145 419 4152 453
rect 4104 412 4152 419
rect 2274 377 2322 384
rect 520 369 568 376
rect 288 329 336 336
rect 288 295 295 329
rect 329 295 336 329
rect 520 335 527 369
rect 561 335 568 369
rect 2274 343 2281 377
rect 2315 343 2322 377
rect 2274 336 2322 343
rect 520 328 568 335
rect 288 288 336 295
rect 4026 325 4074 332
rect 780 285 828 292
rect 780 251 787 285
rect 821 251 828 285
rect 4026 291 4033 325
rect 4067 291 4074 325
rect 4026 284 4074 291
rect 4198 325 4246 332
rect 4198 291 4205 325
rect 4239 291 4246 325
rect 4198 284 4246 291
rect 4340 329 4388 336
rect 4340 295 4347 329
rect 4381 295 4388 329
rect 4340 288 4388 295
rect 4442 325 4490 332
rect 4442 291 4449 325
rect 4483 291 4490 325
rect 4442 284 4490 291
rect 780 244 828 251
rect 2526 273 2574 280
rect 384 235 432 242
rect 384 201 391 235
rect 425 201 432 235
rect 2526 239 2533 273
rect 2567 239 2574 273
rect 2526 232 2574 239
rect 384 194 432 201
rect 1886 223 1934 230
rect 1886 189 1893 223
rect 1927 189 1934 223
rect 1886 182 1934 189
rect 3634 223 3682 230
rect 3634 189 3641 223
rect 3675 189 3682 223
rect 3634 182 3682 189
rect 2186 -37 2234 -30
rect 2186 -71 2193 -37
rect 2227 -71 2234 -37
rect 2186 -78 2234 -71
rect 3636 -41 3684 -34
rect 3636 -75 3643 -41
rect 3677 -75 3684 -41
rect 780 -85 828 -78
rect 3636 -82 3684 -75
rect 780 -119 787 -85
rect 821 -119 828 -85
rect 780 -126 828 -119
rect 2526 -91 2574 -84
rect 2526 -125 2533 -91
rect 2567 -125 2574 -91
rect 2526 -132 2574 -125
rect 520 -145 568 -138
rect 520 -179 527 -145
rect 561 -179 568 -145
rect 520 -186 568 -179
rect 2280 -149 2328 -142
rect 2280 -183 2287 -149
rect 2321 -183 2328 -149
rect 2280 -190 2328 -183
<< viali >>
rect 4111 419 4145 453
rect 295 295 329 329
rect 527 335 561 369
rect 2281 343 2315 377
rect 787 251 821 285
rect 4033 291 4067 325
rect 4205 291 4239 325
rect 4347 295 4381 329
rect 4449 291 4483 325
rect 391 201 425 235
rect 2533 239 2567 273
rect 1893 189 1927 223
rect 3641 189 3675 223
rect 2193 -71 2227 -37
rect 3643 -75 3677 -41
rect 787 -119 821 -85
rect 2533 -125 2567 -91
rect 527 -179 561 -145
rect 2287 -183 2321 -149
<< metal1 >>
rect -10 664 86 670
rect -10 642 132 664
rect -10 590 12 642
rect 64 590 132 642
rect -10 568 132 590
rect -10 562 86 568
rect -72 462 580 466
rect -72 410 518 462
rect 570 410 580 462
rect -72 406 580 410
rect 4092 453 4394 466
rect 4092 419 4111 453
rect 4145 419 4394 453
rect 4092 406 4394 419
rect 514 369 574 406
rect 2268 390 2328 396
rect -72 329 348 342
rect -72 295 295 329
rect 329 295 348 329
rect 514 335 527 369
rect 561 335 574 369
rect 514 316 574 335
rect 2262 386 2334 390
rect 2262 334 2272 386
rect 2324 334 2334 386
rect 4192 338 4252 344
rect 2262 330 2334 334
rect 2268 324 2328 330
rect 3934 325 4086 338
rect -72 282 348 295
rect 774 285 834 304
rect 774 251 787 285
rect 821 251 834 285
rect 774 248 834 251
rect 372 235 834 248
rect 2520 273 2580 292
rect 2520 239 2533 273
rect 2567 239 2580 273
rect 3934 291 4033 325
rect 4067 291 4086 325
rect 3934 278 4086 291
rect 4186 334 4258 338
rect 4186 282 4196 334
rect 4248 282 4258 334
rect 4186 278 4258 282
rect 4334 329 4394 406
rect 4334 295 4347 329
rect 4381 295 4394 329
rect 2520 236 2580 239
rect 3624 236 3684 242
rect 3934 236 3994 278
rect 4192 272 4252 278
rect 4334 276 4394 295
rect 4430 325 4688 338
rect 4430 291 4449 325
rect 4483 291 4688 325
rect 4430 278 4688 291
rect 372 201 391 235
rect 425 201 834 235
rect 372 188 834 201
rect 1874 223 2580 236
rect 1874 189 1893 223
rect 1927 189 2580 223
rect 1874 176 2580 189
rect 3622 232 3994 236
rect 3622 180 3628 232
rect 3680 180 3994 232
rect 3622 176 3994 180
rect 3624 170 3684 176
rect -10 24 232 120
rect 2174 -37 2580 -24
rect 3934 -28 3994 -22
rect 774 -72 834 -66
rect 2174 -71 2193 -37
rect 2227 -71 2580 -37
rect 768 -76 840 -72
rect 514 -132 574 -126
rect 768 -128 778 -76
rect 830 -128 840 -76
rect 2174 -84 2580 -71
rect 768 -132 840 -128
rect 2520 -91 2580 -84
rect 3624 -32 3994 -28
rect 3624 -41 3938 -32
rect 3624 -75 3643 -41
rect 3677 -75 3938 -41
rect 3624 -84 3938 -75
rect 3990 -84 3994 -32
rect 3624 -88 3994 -84
rect 2520 -125 2533 -91
rect 2567 -125 2580 -91
rect 3934 -94 3994 -88
rect 508 -136 580 -132
rect 508 -188 518 -136
rect 570 -188 580 -136
rect 774 -138 834 -132
rect 2274 -136 2334 -130
rect 508 -192 580 -188
rect 2268 -140 2340 -136
rect 2268 -192 2278 -140
rect 2330 -192 2340 -140
rect 2520 -144 2580 -125
rect 514 -198 574 -192
rect 2268 -196 2340 -192
rect 2274 -202 2334 -196
rect -10 -424 86 -418
rect -10 -446 480 -424
rect -10 -498 12 -446
rect 64 -498 480 -446
rect -10 -520 480 -498
rect -10 -526 86 -520
<< via1 >>
rect 12 590 64 642
rect 518 410 570 462
rect 2272 377 2324 386
rect 2272 343 2281 377
rect 2281 343 2315 377
rect 2315 343 2324 377
rect 2272 334 2324 343
rect 4196 325 4248 334
rect 4196 291 4205 325
rect 4205 291 4239 325
rect 4239 291 4248 325
rect 4196 282 4248 291
rect 3628 223 3680 232
rect 3628 189 3641 223
rect 3641 189 3675 223
rect 3675 189 3680 223
rect 3628 180 3680 189
rect 778 -85 830 -76
rect 778 -119 787 -85
rect 787 -119 821 -85
rect 821 -119 830 -85
rect 778 -128 830 -119
rect 3938 -84 3990 -32
rect 518 -145 570 -136
rect 518 -179 527 -145
rect 527 -179 561 -145
rect 561 -179 570 -145
rect 518 -188 570 -179
rect 2278 -149 2330 -140
rect 2278 -183 2287 -149
rect 2287 -183 2321 -149
rect 2321 -183 2330 -149
rect 2278 -192 2330 -183
rect 12 -498 64 -446
<< metal2 >>
rect -16 642 92 664
rect -16 590 12 642
rect 64 590 92 642
rect -16 568 92 590
rect -10 -424 86 568
rect 514 466 574 472
rect 510 462 2332 466
rect 510 410 518 462
rect 570 410 2332 462
rect 510 406 2332 410
rect 514 -136 574 406
rect 2268 386 2328 406
rect 2268 334 2272 386
rect 2324 334 2328 386
rect 2268 324 2328 334
rect 3934 334 4258 338
rect 3934 282 4196 334
rect 4248 282 4258 334
rect 3934 278 4258 282
rect 3618 232 3690 236
rect 3618 180 3628 232
rect 3680 180 3690 232
rect 3618 176 3690 180
rect 3624 102 3684 176
rect 514 -188 518 -136
rect 570 -188 574 -136
rect 774 42 3684 102
rect 774 -76 834 42
rect 3934 -28 3994 278
rect 774 -128 778 -76
rect 830 -128 834 -76
rect 3928 -32 4000 -28
rect 3928 -84 3938 -32
rect 3990 -84 4000 -32
rect 3928 -88 4000 -84
rect 774 -138 834 -128
rect 514 -214 574 -188
rect 2274 -140 2334 -130
rect 2274 -192 2278 -140
rect 2330 -192 2334 -140
rect 2274 -214 2334 -192
rect 514 -274 2334 -214
rect -16 -446 92 -424
rect -16 -498 12 -446
rect 64 -498 92 -446
rect -16 -520 92 -498
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_3
timestamp 1626486988
transform 1 0 500 0 -1 72
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_2
timestamp 1626486988
transform 1 0 500 0 1 72
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_1
timestamp 1626486988
transform 1 0 2248 0 -1 72
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_0
timestamp 1626486988
transform 1 0 2248 0 1 72
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1626486988
transform 1 0 224 0 1 72
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1626486988
transform 1 0 4272 0 1 72
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0
timestamp 1626486988
transform -1 0 4272 0 1 72
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1626486988
transform 1 0 408 0 -1 72
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1626486988
transform 1 0 132 0 1 72
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1626486988
transform 1 0 3996 0 -1 72
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1626486988
transform 1 0 4548 0 1 72
box -38 -48 130 592
<< labels >>
flabel metal2 s 20 502 26 506 1 FreeSans 600 0 0 0 VDD
flabel metal1 s 94 100 96 104 1 FreeSans 600 0 0 0 VSS
flabel metal1 s -52 310 -44 318 1 FreeSans 600 0 0 0 trigb
flabel metal1 s -52 434 -42 442 1 FreeSans 600 0 0 0 clk
flabel metal1 s 4644 304 4650 308 1 FreeSans 600 0 0 0 pulse
<< end >>
