magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< metal1 >>
rect 552 1388 616 1440
rect 1720 1388 1784 1440
rect 2888 1388 2952 1440
rect 4056 1388 4120 1440
rect 5224 1388 5288 1440
rect 6392 1388 6456 1440
rect 7560 1388 7624 1440
rect 8728 1388 8792 1440
rect 9896 1388 9960 1440
rect 11064 1388 11128 1440
rect 12232 1388 12296 1440
rect 13400 1388 13464 1440
rect 14568 1388 14632 1440
rect 15736 1388 15800 1440
rect 16904 1388 16968 1440
rect 18072 1388 18136 1440
rect 19240 1388 19304 1440
rect 20408 1388 20472 1440
rect 21576 1388 21640 1440
rect 22744 1388 22808 1440
rect 23912 1388 23976 1440
rect 25080 1388 25144 1440
rect 26248 1388 26312 1440
rect 27416 1388 27480 1440
rect 28584 1388 28648 1440
rect 29752 1388 29816 1440
rect 30920 1388 30984 1440
rect 32088 1388 32152 1440
rect 33256 1388 33320 1440
rect 34424 1388 34488 1440
rect 35592 1388 35656 1440
rect 36760 1388 36824 1440
rect 552 -26 616 26
rect 1720 -26 1784 26
rect 2888 -26 2952 26
rect 4056 -26 4120 26
rect 5224 -26 5288 26
rect 6392 -26 6456 26
rect 7560 -26 7624 26
rect 8728 -26 8792 26
rect 9896 -26 9960 26
rect 11064 -26 11128 26
rect 12232 -26 12296 26
rect 13400 -26 13464 26
rect 14568 -26 14632 26
rect 15736 -26 15800 26
rect 16904 -26 16968 26
rect 18072 -26 18136 26
rect 19240 -26 19304 26
rect 20408 -26 20472 26
rect 21576 -26 21640 26
rect 22744 -26 22808 26
rect 23912 -26 23976 26
rect 25080 -26 25144 26
rect 26248 -26 26312 26
rect 27416 -26 27480 26
rect 28584 -26 28648 26
rect 29752 -26 29816 26
rect 30920 -26 30984 26
rect 32088 -26 32152 26
rect 33256 -26 33320 26
rect 34424 -26 34488 26
rect 35592 -26 35656 26
rect 36760 -26 36824 26
<< metal2 >>
rect 137 538 203 590
rect 369 0 397 1414
rect 556 1390 612 1438
rect 1082 609 1148 661
rect 1305 538 1371 590
rect 556 -24 612 24
rect 1537 0 1565 1414
rect 1724 1390 1780 1438
rect 2250 609 2316 661
rect 2473 538 2539 590
rect 1724 -24 1780 24
rect 2705 0 2733 1414
rect 2892 1390 2948 1438
rect 3418 609 3484 661
rect 3641 538 3707 590
rect 2892 -24 2948 24
rect 3873 0 3901 1414
rect 4060 1390 4116 1438
rect 4586 609 4652 661
rect 4809 538 4875 590
rect 4060 -24 4116 24
rect 5041 0 5069 1414
rect 5228 1390 5284 1438
rect 5754 609 5820 661
rect 5977 538 6043 590
rect 5228 -24 5284 24
rect 6209 0 6237 1414
rect 6396 1390 6452 1438
rect 6922 609 6988 661
rect 7145 538 7211 590
rect 6396 -24 6452 24
rect 7377 0 7405 1414
rect 7564 1390 7620 1438
rect 8090 609 8156 661
rect 8313 538 8379 590
rect 7564 -24 7620 24
rect 8545 0 8573 1414
rect 8732 1390 8788 1438
rect 9258 609 9324 661
rect 9481 538 9547 590
rect 8732 -24 8788 24
rect 9713 0 9741 1414
rect 9900 1390 9956 1438
rect 10426 609 10492 661
rect 10649 538 10715 590
rect 9900 -24 9956 24
rect 10881 0 10909 1414
rect 11068 1390 11124 1438
rect 11594 609 11660 661
rect 11817 538 11883 590
rect 11068 -24 11124 24
rect 12049 0 12077 1414
rect 12236 1390 12292 1438
rect 12762 609 12828 661
rect 12985 538 13051 590
rect 12236 -24 12292 24
rect 13217 0 13245 1414
rect 13404 1390 13460 1438
rect 13930 609 13996 661
rect 14153 538 14219 590
rect 13404 -24 13460 24
rect 14385 0 14413 1414
rect 14572 1390 14628 1438
rect 15098 609 15164 661
rect 15321 538 15387 590
rect 14572 -24 14628 24
rect 15553 0 15581 1414
rect 15740 1390 15796 1438
rect 16266 609 16332 661
rect 16489 538 16555 590
rect 15740 -24 15796 24
rect 16721 0 16749 1414
rect 16908 1390 16964 1438
rect 17434 609 17500 661
rect 17657 538 17723 590
rect 16908 -24 16964 24
rect 17889 0 17917 1414
rect 18076 1390 18132 1438
rect 18602 609 18668 661
rect 18825 538 18891 590
rect 18076 -24 18132 24
rect 19057 0 19085 1414
rect 19244 1390 19300 1438
rect 19770 609 19836 661
rect 19993 538 20059 590
rect 19244 -24 19300 24
rect 20225 0 20253 1414
rect 20412 1390 20468 1438
rect 20938 609 21004 661
rect 21161 538 21227 590
rect 20412 -24 20468 24
rect 21393 0 21421 1414
rect 21580 1390 21636 1438
rect 22106 609 22172 661
rect 22329 538 22395 590
rect 21580 -24 21636 24
rect 22561 0 22589 1414
rect 22748 1390 22804 1438
rect 23274 609 23340 661
rect 23497 538 23563 590
rect 22748 -24 22804 24
rect 23729 0 23757 1414
rect 23916 1390 23972 1438
rect 24442 609 24508 661
rect 24665 538 24731 590
rect 23916 -24 23972 24
rect 24897 0 24925 1414
rect 25084 1390 25140 1438
rect 25610 609 25676 661
rect 25833 538 25899 590
rect 25084 -24 25140 24
rect 26065 0 26093 1414
rect 26252 1390 26308 1438
rect 26778 609 26844 661
rect 27001 538 27067 590
rect 26252 -24 26308 24
rect 27233 0 27261 1414
rect 27420 1390 27476 1438
rect 27946 609 28012 661
rect 28169 538 28235 590
rect 27420 -24 27476 24
rect 28401 0 28429 1414
rect 28588 1390 28644 1438
rect 29114 609 29180 661
rect 29337 538 29403 590
rect 28588 -24 28644 24
rect 29569 0 29597 1414
rect 29756 1390 29812 1438
rect 30282 609 30348 661
rect 30505 538 30571 590
rect 29756 -24 29812 24
rect 30737 0 30765 1414
rect 30924 1390 30980 1438
rect 31450 609 31516 661
rect 31673 538 31739 590
rect 30924 -24 30980 24
rect 31905 0 31933 1414
rect 32092 1390 32148 1438
rect 32618 609 32684 661
rect 32841 538 32907 590
rect 32092 -24 32148 24
rect 33073 0 33101 1414
rect 33260 1390 33316 1438
rect 33786 609 33852 661
rect 34009 538 34075 590
rect 33260 -24 33316 24
rect 34241 0 34269 1414
rect 34428 1390 34484 1438
rect 34954 609 35020 661
rect 35177 538 35243 590
rect 34428 -24 34484 24
rect 35409 0 35437 1414
rect 35596 1390 35652 1438
rect 36122 609 36188 661
rect 36345 538 36411 590
rect 35596 -24 35652 24
rect 36577 0 36605 1414
rect 36764 1390 36820 1438
rect 37290 609 37356 661
rect 36764 -24 36820 24
<< metal3 >>
rect 535 1365 633 1463
rect 1703 1365 1801 1463
rect 2871 1365 2969 1463
rect 4039 1365 4137 1463
rect 5207 1365 5305 1463
rect 6375 1365 6473 1463
rect 7543 1365 7641 1463
rect 8711 1365 8809 1463
rect 9879 1365 9977 1463
rect 11047 1365 11145 1463
rect 12215 1365 12313 1463
rect 13383 1365 13481 1463
rect 14551 1365 14649 1463
rect 15719 1365 15817 1463
rect 16887 1365 16985 1463
rect 18055 1365 18153 1463
rect 19223 1365 19321 1463
rect 20391 1365 20489 1463
rect 21559 1365 21657 1463
rect 22727 1365 22825 1463
rect 23895 1365 23993 1463
rect 25063 1365 25161 1463
rect 26231 1365 26329 1463
rect 27399 1365 27497 1463
rect 28567 1365 28665 1463
rect 29735 1365 29833 1463
rect 30903 1365 31001 1463
rect 32071 1365 32169 1463
rect 33239 1365 33337 1463
rect 34407 1365 34505 1463
rect 35575 1365 35673 1463
rect 36743 1365 36841 1463
rect 0 278 37376 338
rect 535 -49 633 49
rect 1703 -49 1801 49
rect 2871 -49 2969 49
rect 4039 -49 4137 49
rect 5207 -49 5305 49
rect 6375 -49 6473 49
rect 7543 -49 7641 49
rect 8711 -49 8809 49
rect 9879 -49 9977 49
rect 11047 -49 11145 49
rect 12215 -49 12313 49
rect 13383 -49 13481 49
rect 14551 -49 14649 49
rect 15719 -49 15817 49
rect 16887 -49 16985 49
rect 18055 -49 18153 49
rect 19223 -49 19321 49
rect 20391 -49 20489 49
rect 21559 -49 21657 49
rect 22727 -49 22825 49
rect 23895 -49 23993 49
rect 25063 -49 25161 49
rect 26231 -49 26329 49
rect 27399 -49 27497 49
rect 28567 -49 28665 49
rect 29735 -49 29833 49
rect 30903 -49 31001 49
rect 32071 -49 32169 49
rect 33239 -49 33337 49
rect 34407 -49 34505 49
rect 35575 -49 35673 49
rect 36743 -49 36841 49
use contact_9  contact_9_31
timestamp 1624494425
transform 1 0 363 0 1 271
box 0 0 66 74
use contact_9  contact_9_94
timestamp 1624494425
transform 1 0 551 0 1 -37
box 0 0 66 74
use contact_9  contact_9_95
timestamp 1624494425
transform 1 0 551 0 1 1377
box 0 0 66 74
use contact_8  contact_8_62
timestamp 1624494425
transform 1 0 552 0 1 -32
box 0 0 64 64
use contact_8  contact_8_63
timestamp 1624494425
transform 1 0 552 0 1 1382
box 0 0 64 64
use contact_7  contact_7_62
timestamp 1624494425
transform 1 0 555 0 1 -33
box 0 0 58 66
use contact_7  contact_7_63
timestamp 1624494425
transform 1 0 555 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_30
timestamp 1624494425
transform 1 0 1168 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_31
timestamp 1624494425
transform 1 0 0 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_30
timestamp 1624494425
transform 1 0 1531 0 1 271
box 0 0 66 74
use contact_9  contact_9_92
timestamp 1624494425
transform 1 0 1719 0 1 -37
box 0 0 66 74
use contact_9  contact_9_93
timestamp 1624494425
transform 1 0 1719 0 1 1377
box 0 0 66 74
use contact_8  contact_8_60
timestamp 1624494425
transform 1 0 1720 0 1 -32
box 0 0 64 64
use contact_8  contact_8_61
timestamp 1624494425
transform 1 0 1720 0 1 1382
box 0 0 64 64
use contact_7  contact_7_60
timestamp 1624494425
transform 1 0 1723 0 1 -33
box 0 0 58 66
use contact_7  contact_7_61
timestamp 1624494425
transform 1 0 1723 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_29
timestamp 1624494425
transform 1 0 2336 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_29
timestamp 1624494425
transform 1 0 2699 0 1 271
box 0 0 66 74
use contact_9  contact_9_90
timestamp 1624494425
transform 1 0 2887 0 1 -37
box 0 0 66 74
use contact_9  contact_9_91
timestamp 1624494425
transform 1 0 2887 0 1 1377
box 0 0 66 74
use contact_8  contact_8_58
timestamp 1624494425
transform 1 0 2888 0 1 -32
box 0 0 64 64
use contact_8  contact_8_59
timestamp 1624494425
transform 1 0 2888 0 1 1382
box 0 0 64 64
use contact_7  contact_7_58
timestamp 1624494425
transform 1 0 2891 0 1 -33
box 0 0 58 66
use contact_7  contact_7_59
timestamp 1624494425
transform 1 0 2891 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_28
timestamp 1624494425
transform 1 0 3504 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_28
timestamp 1624494425
transform 1 0 3867 0 1 271
box 0 0 66 74
use contact_9  contact_9_88
timestamp 1624494425
transform 1 0 4055 0 1 -37
box 0 0 66 74
use contact_9  contact_9_89
timestamp 1624494425
transform 1 0 4055 0 1 1377
box 0 0 66 74
use contact_8  contact_8_56
timestamp 1624494425
transform 1 0 4056 0 1 -32
box 0 0 64 64
use contact_8  contact_8_57
timestamp 1624494425
transform 1 0 4056 0 1 1382
box 0 0 64 64
use contact_7  contact_7_56
timestamp 1624494425
transform 1 0 4059 0 1 -33
box 0 0 58 66
use contact_7  contact_7_57
timestamp 1624494425
transform 1 0 4059 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_27
timestamp 1624494425
transform 1 0 4672 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_27
timestamp 1624494425
transform 1 0 5035 0 1 271
box 0 0 66 74
use contact_9  contact_9_86
timestamp 1624494425
transform 1 0 5223 0 1 -37
box 0 0 66 74
use contact_9  contact_9_87
timestamp 1624494425
transform 1 0 5223 0 1 1377
box 0 0 66 74
use contact_8  contact_8_54
timestamp 1624494425
transform 1 0 5224 0 1 -32
box 0 0 64 64
use contact_8  contact_8_55
timestamp 1624494425
transform 1 0 5224 0 1 1382
box 0 0 64 64
use contact_7  contact_7_54
timestamp 1624494425
transform 1 0 5227 0 1 -33
box 0 0 58 66
use contact_7  contact_7_55
timestamp 1624494425
transform 1 0 5227 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_26
timestamp 1624494425
transform 1 0 5840 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_25
timestamp 1624494425
transform 1 0 7371 0 1 271
box 0 0 66 74
use contact_9  contact_9_26
timestamp 1624494425
transform 1 0 6203 0 1 271
box 0 0 66 74
use contact_9  contact_9_84
timestamp 1624494425
transform 1 0 6391 0 1 -37
box 0 0 66 74
use contact_9  contact_9_85
timestamp 1624494425
transform 1 0 6391 0 1 1377
box 0 0 66 74
use contact_8  contact_8_52
timestamp 1624494425
transform 1 0 6392 0 1 -32
box 0 0 64 64
use contact_8  contact_8_53
timestamp 1624494425
transform 1 0 6392 0 1 1382
box 0 0 64 64
use contact_7  contact_7_52
timestamp 1624494425
transform 1 0 6395 0 1 -33
box 0 0 58 66
use contact_7  contact_7_53
timestamp 1624494425
transform 1 0 6395 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_25
timestamp 1624494425
transform 1 0 7008 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_24
timestamp 1624494425
transform 1 0 8539 0 1 271
box 0 0 66 74
use contact_9  contact_9_82
timestamp 1624494425
transform 1 0 7559 0 1 -37
box 0 0 66 74
use contact_9  contact_9_83
timestamp 1624494425
transform 1 0 7559 0 1 1377
box 0 0 66 74
use contact_8  contact_8_50
timestamp 1624494425
transform 1 0 7560 0 1 -32
box 0 0 64 64
use contact_8  contact_8_51
timestamp 1624494425
transform 1 0 7560 0 1 1382
box 0 0 64 64
use contact_7  contact_7_50
timestamp 1624494425
transform 1 0 7563 0 1 -33
box 0 0 58 66
use contact_7  contact_7_51
timestamp 1624494425
transform 1 0 7563 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_24
timestamp 1624494425
transform 1 0 8176 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_23
timestamp 1624494425
transform 1 0 9707 0 1 271
box 0 0 66 74
use contact_9  contact_9_80
timestamp 1624494425
transform 1 0 8727 0 1 -37
box 0 0 66 74
use contact_9  contact_9_81
timestamp 1624494425
transform 1 0 8727 0 1 1377
box 0 0 66 74
use contact_8  contact_8_48
timestamp 1624494425
transform 1 0 8728 0 1 -32
box 0 0 64 64
use contact_8  contact_8_49
timestamp 1624494425
transform 1 0 8728 0 1 1382
box 0 0 64 64
use contact_7  contact_7_48
timestamp 1624494425
transform 1 0 8731 0 1 -33
box 0 0 58 66
use contact_7  contact_7_49
timestamp 1624494425
transform 1 0 8731 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_23
timestamp 1624494425
transform 1 0 9344 0 1 0
box -36 -43 1204 1467
use contact_7  contact_7_46
timestamp 1624494425
transform 1 0 9899 0 1 -33
box 0 0 58 66
use contact_7  contact_7_44
timestamp 1624494425
transform 1 0 11067 0 1 -33
box 0 0 58 66
use contact_8  contact_8_46
timestamp 1624494425
transform 1 0 9896 0 1 -32
box 0 0 64 64
use contact_8  contact_8_44
timestamp 1624494425
transform 1 0 11064 0 1 -32
box 0 0 64 64
use contact_9  contact_9_78
timestamp 1624494425
transform 1 0 9895 0 1 -37
box 0 0 66 74
use contact_9  contact_9_76
timestamp 1624494425
transform 1 0 11063 0 1 -37
box 0 0 66 74
use contact_9  contact_9_22
timestamp 1624494425
transform 1 0 10875 0 1 271
box 0 0 66 74
use contact_7  contact_7_47
timestamp 1624494425
transform 1 0 9899 0 1 1381
box 0 0 58 66
use contact_7  contact_7_45
timestamp 1624494425
transform 1 0 11067 0 1 1381
box 0 0 58 66
use contact_8  contact_8_47
timestamp 1624494425
transform 1 0 9896 0 1 1382
box 0 0 64 64
use contact_8  contact_8_45
timestamp 1624494425
transform 1 0 11064 0 1 1382
box 0 0 64 64
use contact_9  contact_9_79
timestamp 1624494425
transform 1 0 9895 0 1 1377
box 0 0 66 74
use contact_9  contact_9_77
timestamp 1624494425
transform 1 0 11063 0 1 1377
box 0 0 66 74
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_22
timestamp 1624494425
transform 1 0 10512 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_21
timestamp 1624494425
transform 1 0 12043 0 1 271
box 0 0 66 74
use contact_9  contact_9_74
timestamp 1624494425
transform 1 0 12231 0 1 -37
box 0 0 66 74
use contact_9  contact_9_75
timestamp 1624494425
transform 1 0 12231 0 1 1377
box 0 0 66 74
use contact_8  contact_8_42
timestamp 1624494425
transform 1 0 12232 0 1 -32
box 0 0 64 64
use contact_8  contact_8_43
timestamp 1624494425
transform 1 0 12232 0 1 1382
box 0 0 64 64
use contact_7  contact_7_42
timestamp 1624494425
transform 1 0 12235 0 1 -33
box 0 0 58 66
use contact_7  contact_7_43
timestamp 1624494425
transform 1 0 12235 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_21
timestamp 1624494425
transform 1 0 11680 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_20
timestamp 1624494425
transform 1 0 13211 0 1 271
box 0 0 66 74
use contact_9  contact_9_72
timestamp 1624494425
transform 1 0 13399 0 1 -37
box 0 0 66 74
use contact_9  contact_9_73
timestamp 1624494425
transform 1 0 13399 0 1 1377
box 0 0 66 74
use contact_8  contact_8_40
timestamp 1624494425
transform 1 0 13400 0 1 -32
box 0 0 64 64
use contact_8  contact_8_41
timestamp 1624494425
transform 1 0 13400 0 1 1382
box 0 0 64 64
use contact_7  contact_7_40
timestamp 1624494425
transform 1 0 13403 0 1 -33
box 0 0 58 66
use contact_7  contact_7_41
timestamp 1624494425
transform 1 0 13403 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_20
timestamp 1624494425
transform 1 0 12848 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_19
timestamp 1624494425
transform 1 0 14379 0 1 271
box 0 0 66 74
use contact_9  contact_9_70
timestamp 1624494425
transform 1 0 14567 0 1 -37
box 0 0 66 74
use contact_9  contact_9_71
timestamp 1624494425
transform 1 0 14567 0 1 1377
box 0 0 66 74
use contact_8  contact_8_38
timestamp 1624494425
transform 1 0 14568 0 1 -32
box 0 0 64 64
use contact_8  contact_8_39
timestamp 1624494425
transform 1 0 14568 0 1 1382
box 0 0 64 64
use contact_7  contact_7_38
timestamp 1624494425
transform 1 0 14571 0 1 -33
box 0 0 58 66
use contact_7  contact_7_39
timestamp 1624494425
transform 1 0 14571 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_19
timestamp 1624494425
transform 1 0 14016 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_18
timestamp 1624494425
transform 1 0 15547 0 1 271
box 0 0 66 74
use contact_9  contact_9_68
timestamp 1624494425
transform 1 0 15735 0 1 -37
box 0 0 66 74
use contact_9  contact_9_69
timestamp 1624494425
transform 1 0 15735 0 1 1377
box 0 0 66 74
use contact_8  contact_8_36
timestamp 1624494425
transform 1 0 15736 0 1 -32
box 0 0 64 64
use contact_8  contact_8_37
timestamp 1624494425
transform 1 0 15736 0 1 1382
box 0 0 64 64
use contact_7  contact_7_36
timestamp 1624494425
transform 1 0 15739 0 1 -33
box 0 0 58 66
use contact_7  contact_7_37
timestamp 1624494425
transform 1 0 15739 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_18
timestamp 1624494425
transform 1 0 15184 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_17
timestamp 1624494425
transform 1 0 16715 0 1 271
box 0 0 66 74
use contact_9  contact_9_66
timestamp 1624494425
transform 1 0 16903 0 1 -37
box 0 0 66 74
use contact_9  contact_9_67
timestamp 1624494425
transform 1 0 16903 0 1 1377
box 0 0 66 74
use contact_8  contact_8_34
timestamp 1624494425
transform 1 0 16904 0 1 -32
box 0 0 64 64
use contact_8  contact_8_35
timestamp 1624494425
transform 1 0 16904 0 1 1382
box 0 0 64 64
use contact_7  contact_7_34
timestamp 1624494425
transform 1 0 16907 0 1 -33
box 0 0 58 66
use contact_7  contact_7_35
timestamp 1624494425
transform 1 0 16907 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_17
timestamp 1624494425
transform 1 0 16352 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_16
timestamp 1624494425
transform 1 0 17883 0 1 271
box 0 0 66 74
use contact_9  contact_9_64
timestamp 1624494425
transform 1 0 18071 0 1 -37
box 0 0 66 74
use contact_9  contact_9_65
timestamp 1624494425
transform 1 0 18071 0 1 1377
box 0 0 66 74
use contact_8  contact_8_32
timestamp 1624494425
transform 1 0 18072 0 1 -32
box 0 0 64 64
use contact_8  contact_8_33
timestamp 1624494425
transform 1 0 18072 0 1 1382
box 0 0 64 64
use contact_7  contact_7_32
timestamp 1624494425
transform 1 0 18075 0 1 -33
box 0 0 58 66
use contact_7  contact_7_33
timestamp 1624494425
transform 1 0 18075 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_16
timestamp 1624494425
transform 1 0 17520 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_15
timestamp 1624494425
transform 1 0 19051 0 1 271
box 0 0 66 74
use contact_9  contact_9_62
timestamp 1624494425
transform 1 0 19239 0 1 -37
box 0 0 66 74
use contact_9  contact_9_63
timestamp 1624494425
transform 1 0 19239 0 1 1377
box 0 0 66 74
use contact_8  contact_8_30
timestamp 1624494425
transform 1 0 19240 0 1 -32
box 0 0 64 64
use contact_8  contact_8_31
timestamp 1624494425
transform 1 0 19240 0 1 1382
box 0 0 64 64
use contact_7  contact_7_30
timestamp 1624494425
transform 1 0 19243 0 1 -33
box 0 0 58 66
use contact_7  contact_7_31
timestamp 1624494425
transform 1 0 19243 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_15
timestamp 1624494425
transform 1 0 18688 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_14
timestamp 1624494425
transform 1 0 20219 0 1 271
box 0 0 66 74
use contact_9  contact_9_60
timestamp 1624494425
transform 1 0 20407 0 1 -37
box 0 0 66 74
use contact_9  contact_9_61
timestamp 1624494425
transform 1 0 20407 0 1 1377
box 0 0 66 74
use contact_8  contact_8_28
timestamp 1624494425
transform 1 0 20408 0 1 -32
box 0 0 64 64
use contact_8  contact_8_29
timestamp 1624494425
transform 1 0 20408 0 1 1382
box 0 0 64 64
use contact_7  contact_7_28
timestamp 1624494425
transform 1 0 20411 0 1 -33
box 0 0 58 66
use contact_7  contact_7_29
timestamp 1624494425
transform 1 0 20411 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_13
timestamp 1624494425
transform 1 0 21024 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_14
timestamp 1624494425
transform 1 0 19856 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_13
timestamp 1624494425
transform 1 0 21387 0 1 271
box 0 0 66 74
use contact_9  contact_9_58
timestamp 1624494425
transform 1 0 21575 0 1 -37
box 0 0 66 74
use contact_9  contact_9_59
timestamp 1624494425
transform 1 0 21575 0 1 1377
box 0 0 66 74
use contact_8  contact_8_26
timestamp 1624494425
transform 1 0 21576 0 1 -32
box 0 0 64 64
use contact_8  contact_8_27
timestamp 1624494425
transform 1 0 21576 0 1 1382
box 0 0 64 64
use contact_7  contact_7_26
timestamp 1624494425
transform 1 0 21579 0 1 -33
box 0 0 58 66
use contact_7  contact_7_27
timestamp 1624494425
transform 1 0 21579 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_12
timestamp 1624494425
transform 1 0 22192 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_12
timestamp 1624494425
transform 1 0 22555 0 1 271
box 0 0 66 74
use contact_9  contact_9_56
timestamp 1624494425
transform 1 0 22743 0 1 -37
box 0 0 66 74
use contact_9  contact_9_57
timestamp 1624494425
transform 1 0 22743 0 1 1377
box 0 0 66 74
use contact_8  contact_8_24
timestamp 1624494425
transform 1 0 22744 0 1 -32
box 0 0 64 64
use contact_8  contact_8_25
timestamp 1624494425
transform 1 0 22744 0 1 1382
box 0 0 64 64
use contact_7  contact_7_24
timestamp 1624494425
transform 1 0 22747 0 1 -33
box 0 0 58 66
use contact_7  contact_7_25
timestamp 1624494425
transform 1 0 22747 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_11
timestamp 1624494425
transform 1 0 23360 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_11
timestamp 1624494425
transform 1 0 23723 0 1 271
box 0 0 66 74
use contact_9  contact_9_54
timestamp 1624494425
transform 1 0 23911 0 1 -37
box 0 0 66 74
use contact_9  contact_9_55
timestamp 1624494425
transform 1 0 23911 0 1 1377
box 0 0 66 74
use contact_8  contact_8_22
timestamp 1624494425
transform 1 0 23912 0 1 -32
box 0 0 64 64
use contact_8  contact_8_23
timestamp 1624494425
transform 1 0 23912 0 1 1382
box 0 0 64 64
use contact_7  contact_7_22
timestamp 1624494425
transform 1 0 23915 0 1 -33
box 0 0 58 66
use contact_7  contact_7_23
timestamp 1624494425
transform 1 0 23915 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_10
timestamp 1624494425
transform 1 0 24528 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_10
timestamp 1624494425
transform 1 0 24891 0 1 271
box 0 0 66 74
use contact_9  contact_9_52
timestamp 1624494425
transform 1 0 25079 0 1 -37
box 0 0 66 74
use contact_9  contact_9_53
timestamp 1624494425
transform 1 0 25079 0 1 1377
box 0 0 66 74
use contact_8  contact_8_20
timestamp 1624494425
transform 1 0 25080 0 1 -32
box 0 0 64 64
use contact_8  contact_8_21
timestamp 1624494425
transform 1 0 25080 0 1 1382
box 0 0 64 64
use contact_7  contact_7_20
timestamp 1624494425
transform 1 0 25083 0 1 -33
box 0 0 58 66
use contact_7  contact_7_21
timestamp 1624494425
transform 1 0 25083 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_9
timestamp 1624494425
transform 1 0 25696 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_8
timestamp 1624494425
transform 1 0 27227 0 1 271
box 0 0 66 74
use contact_9  contact_9_9
timestamp 1624494425
transform 1 0 26059 0 1 271
box 0 0 66 74
use contact_9  contact_9_50
timestamp 1624494425
transform 1 0 26247 0 1 -37
box 0 0 66 74
use contact_9  contact_9_51
timestamp 1624494425
transform 1 0 26247 0 1 1377
box 0 0 66 74
use contact_8  contact_8_18
timestamp 1624494425
transform 1 0 26248 0 1 -32
box 0 0 64 64
use contact_8  contact_8_19
timestamp 1624494425
transform 1 0 26248 0 1 1382
box 0 0 64 64
use contact_7  contact_7_18
timestamp 1624494425
transform 1 0 26251 0 1 -33
box 0 0 58 66
use contact_7  contact_7_19
timestamp 1624494425
transform 1 0 26251 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_8
timestamp 1624494425
transform 1 0 26864 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_7
timestamp 1624494425
transform 1 0 28395 0 1 271
box 0 0 66 74
use contact_9  contact_9_48
timestamp 1624494425
transform 1 0 27415 0 1 -37
box 0 0 66 74
use contact_9  contact_9_49
timestamp 1624494425
transform 1 0 27415 0 1 1377
box 0 0 66 74
use contact_8  contact_8_16
timestamp 1624494425
transform 1 0 27416 0 1 -32
box 0 0 64 64
use contact_8  contact_8_17
timestamp 1624494425
transform 1 0 27416 0 1 1382
box 0 0 64 64
use contact_7  contact_7_16
timestamp 1624494425
transform 1 0 27419 0 1 -33
box 0 0 58 66
use contact_7  contact_7_17
timestamp 1624494425
transform 1 0 27419 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_7
timestamp 1624494425
transform 1 0 28032 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_6
timestamp 1624494425
transform 1 0 29563 0 1 271
box 0 0 66 74
use contact_9  contact_9_46
timestamp 1624494425
transform 1 0 28583 0 1 -37
box 0 0 66 74
use contact_9  contact_9_47
timestamp 1624494425
transform 1 0 28583 0 1 1377
box 0 0 66 74
use contact_8  contact_8_14
timestamp 1624494425
transform 1 0 28584 0 1 -32
box 0 0 64 64
use contact_8  contact_8_15
timestamp 1624494425
transform 1 0 28584 0 1 1382
box 0 0 64 64
use contact_7  contact_7_14
timestamp 1624494425
transform 1 0 28587 0 1 -33
box 0 0 58 66
use contact_7  contact_7_15
timestamp 1624494425
transform 1 0 28587 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_6
timestamp 1624494425
transform 1 0 29200 0 1 0
box -36 -43 1204 1467
use contact_7  contact_7_12
timestamp 1624494425
transform 1 0 29755 0 1 -33
box 0 0 58 66
use contact_7  contact_7_10
timestamp 1624494425
transform 1 0 30923 0 1 -33
box 0 0 58 66
use contact_8  contact_8_12
timestamp 1624494425
transform 1 0 29752 0 1 -32
box 0 0 64 64
use contact_8  contact_8_10
timestamp 1624494425
transform 1 0 30920 0 1 -32
box 0 0 64 64
use contact_9  contact_9_44
timestamp 1624494425
transform 1 0 29751 0 1 -37
box 0 0 66 74
use contact_9  contact_9_42
timestamp 1624494425
transform 1 0 30919 0 1 -37
box 0 0 66 74
use contact_9  contact_9_5
timestamp 1624494425
transform 1 0 30731 0 1 271
box 0 0 66 74
use contact_7  contact_7_13
timestamp 1624494425
transform 1 0 29755 0 1 1381
box 0 0 58 66
use contact_7  contact_7_11
timestamp 1624494425
transform 1 0 30923 0 1 1381
box 0 0 58 66
use contact_8  contact_8_13
timestamp 1624494425
transform 1 0 29752 0 1 1382
box 0 0 64 64
use contact_8  contact_8_11
timestamp 1624494425
transform 1 0 30920 0 1 1382
box 0 0 64 64
use contact_9  contact_9_45
timestamp 1624494425
transform 1 0 29751 0 1 1377
box 0 0 66 74
use contact_9  contact_9_43
timestamp 1624494425
transform 1 0 30919 0 1 1377
box 0 0 66 74
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_5
timestamp 1624494425
transform 1 0 30368 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_4
timestamp 1624494425
transform 1 0 31899 0 1 271
box 0 0 66 74
use contact_9  contact_9_40
timestamp 1624494425
transform 1 0 32087 0 1 -37
box 0 0 66 74
use contact_9  contact_9_41
timestamp 1624494425
transform 1 0 32087 0 1 1377
box 0 0 66 74
use contact_8  contact_8_8
timestamp 1624494425
transform 1 0 32088 0 1 -32
box 0 0 64 64
use contact_8  contact_8_9
timestamp 1624494425
transform 1 0 32088 0 1 1382
box 0 0 64 64
use contact_7  contact_7_8
timestamp 1624494425
transform 1 0 32091 0 1 -33
box 0 0 58 66
use contact_7  contact_7_9
timestamp 1624494425
transform 1 0 32091 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_4
timestamp 1624494425
transform 1 0 31536 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_3
timestamp 1624494425
transform 1 0 33067 0 1 271
box 0 0 66 74
use contact_9  contact_9_38
timestamp 1624494425
transform 1 0 33255 0 1 -37
box 0 0 66 74
use contact_9  contact_9_39
timestamp 1624494425
transform 1 0 33255 0 1 1377
box 0 0 66 74
use contact_8  contact_8_6
timestamp 1624494425
transform 1 0 33256 0 1 -32
box 0 0 64 64
use contact_8  contact_8_7
timestamp 1624494425
transform 1 0 33256 0 1 1382
box 0 0 64 64
use contact_7  contact_7_6
timestamp 1624494425
transform 1 0 33259 0 1 -33
box 0 0 58 66
use contact_7  contact_7_7
timestamp 1624494425
transform 1 0 33259 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_3
timestamp 1624494425
transform 1 0 32704 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_2
timestamp 1624494425
transform 1 0 34235 0 1 271
box 0 0 66 74
use contact_9  contact_9_36
timestamp 1624494425
transform 1 0 34423 0 1 -37
box 0 0 66 74
use contact_9  contact_9_37
timestamp 1624494425
transform 1 0 34423 0 1 1377
box 0 0 66 74
use contact_8  contact_8_4
timestamp 1624494425
transform 1 0 34424 0 1 -32
box 0 0 64 64
use contact_8  contact_8_5
timestamp 1624494425
transform 1 0 34424 0 1 1382
box 0 0 64 64
use contact_7  contact_7_4
timestamp 1624494425
transform 1 0 34427 0 1 -33
box 0 0 58 66
use contact_7  contact_7_5
timestamp 1624494425
transform 1 0 34427 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_2
timestamp 1624494425
transform 1 0 33872 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_1
timestamp 1624494425
transform 1 0 35403 0 1 271
box 0 0 66 74
use contact_9  contact_9_34
timestamp 1624494425
transform 1 0 35591 0 1 -37
box 0 0 66 74
use contact_9  contact_9_35
timestamp 1624494425
transform 1 0 35591 0 1 1377
box 0 0 66 74
use contact_8  contact_8_2
timestamp 1624494425
transform 1 0 35592 0 1 -32
box 0 0 64 64
use contact_8  contact_8_3
timestamp 1624494425
transform 1 0 35592 0 1 1382
box 0 0 64 64
use contact_7  contact_7_2
timestamp 1624494425
transform 1 0 35595 0 1 -33
box 0 0 58 66
use contact_7  contact_7_3
timestamp 1624494425
transform 1 0 35595 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_1
timestamp 1624494425
transform 1 0 35040 0 1 0
box -36 -43 1204 1467
use contact_9  contact_9_0
timestamp 1624494425
transform 1 0 36571 0 1 271
box 0 0 66 74
use contact_9  contact_9_32
timestamp 1624494425
transform 1 0 36759 0 1 -37
box 0 0 66 74
use contact_9  contact_9_33
timestamp 1624494425
transform 1 0 36759 0 1 1377
box 0 0 66 74
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 36760 0 1 -32
box 0 0 64 64
use contact_8  contact_8_1
timestamp 1624494425
transform 1 0 36760 0 1 1382
box 0 0 64 64
use contact_7  contact_7_0
timestamp 1624494425
transform 1 0 36763 0 1 -33
box 0 0 58 66
use contact_7  contact_7_1
timestamp 1624494425
transform 1 0 36763 0 1 1381
box 0 0 58 66
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_0
timestamp 1624494425
transform 1 0 36208 0 1 0
box -36 -43 1204 1467
<< labels >>
rlabel metal3 s 9879 1365 9977 1463 4 vdd
rlabel metal3 s 12215 1365 12313 1463 4 vdd
rlabel metal3 s 2871 1365 2969 1463 4 vdd
rlabel metal3 s 19223 1365 19321 1463 4 vdd
rlabel metal3 s 34407 1365 34505 1463 4 vdd
rlabel metal3 s 5207 1365 5305 1463 4 vdd
rlabel metal3 s 22727 1365 22825 1463 4 vdd
rlabel metal3 s 36743 1365 36841 1463 4 vdd
rlabel metal3 s 21559 1365 21657 1463 4 vdd
rlabel metal3 s 1703 1365 1801 1463 4 vdd
rlabel metal3 s 535 1365 633 1463 4 vdd
rlabel metal3 s 13383 1365 13481 1463 4 vdd
rlabel metal3 s 11047 1365 11145 1463 4 vdd
rlabel metal3 s 14551 1365 14649 1463 4 vdd
rlabel metal3 s 25063 1365 25161 1463 4 vdd
rlabel metal3 s 30903 1365 31001 1463 4 vdd
rlabel metal3 s 28567 1365 28665 1463 4 vdd
rlabel metal3 s 29735 1365 29833 1463 4 vdd
rlabel metal3 s 15719 1365 15817 1463 4 vdd
rlabel metal3 s 16887 1365 16985 1463 4 vdd
rlabel metal3 s 7543 1365 7641 1463 4 vdd
rlabel metal3 s 23895 1365 23993 1463 4 vdd
rlabel metal3 s 27399 1365 27497 1463 4 vdd
rlabel metal3 s 4039 1365 4137 1463 4 vdd
rlabel metal3 s 33239 1365 33337 1463 4 vdd
rlabel metal3 s 32071 1365 32169 1463 4 vdd
rlabel metal3 s 20391 1365 20489 1463 4 vdd
rlabel metal3 s 18055 1365 18153 1463 4 vdd
rlabel metal3 s 6375 1365 6473 1463 4 vdd
rlabel metal3 s 8711 1365 8809 1463 4 vdd
rlabel metal3 s 26231 1365 26329 1463 4 vdd
rlabel metal3 s 35575 1365 35673 1463 4 vdd
rlabel metal3 s 34407 -49 34505 49 4 gnd
rlabel metal3 s 12215 -49 12313 49 4 gnd
rlabel metal3 s 30903 -49 31001 49 4 gnd
rlabel metal3 s 25063 -49 25161 49 4 gnd
rlabel metal3 s 23895 -49 23993 49 4 gnd
rlabel metal3 s 8711 -49 8809 49 4 gnd
rlabel metal3 s 19223 -49 19321 49 4 gnd
rlabel metal3 s 27399 -49 27497 49 4 gnd
rlabel metal3 s 16887 -49 16985 49 4 gnd
rlabel metal3 s 21559 -49 21657 49 4 gnd
rlabel metal3 s 35575 -49 35673 49 4 gnd
rlabel metal3 s 15719 -49 15817 49 4 gnd
rlabel metal3 s 26231 -49 26329 49 4 gnd
rlabel metal3 s 13383 -49 13481 49 4 gnd
rlabel metal3 s 6375 -49 6473 49 4 gnd
rlabel metal3 s 5207 -49 5305 49 4 gnd
rlabel metal3 s 20391 -49 20489 49 4 gnd
rlabel metal3 s 1703 -49 1801 49 4 gnd
rlabel metal3 s 7543 -49 7641 49 4 gnd
rlabel metal3 s 4039 -49 4137 49 4 gnd
rlabel metal3 s 36743 -49 36841 49 4 gnd
rlabel metal3 s 33239 -49 33337 49 4 gnd
rlabel metal3 s 14551 -49 14649 49 4 gnd
rlabel metal3 s 11047 -49 11145 49 4 gnd
rlabel metal3 s 535 -49 633 49 4 gnd
rlabel metal3 s 9879 -49 9977 49 4 gnd
rlabel metal3 s 2871 -49 2969 49 4 gnd
rlabel metal3 s 28567 -49 28665 49 4 gnd
rlabel metal3 s 32071 -49 32169 49 4 gnd
rlabel metal3 s 18055 -49 18153 49 4 gnd
rlabel metal3 s 22727 -49 22825 49 4 gnd
rlabel metal3 s 29735 -49 29833 49 4 gnd
rlabel metal2 s 137 538 203 590 4 din_0
rlabel metal2 s 1082 609 1148 661 4 dout_0
rlabel metal2 s 1305 538 1371 590 4 din_1
rlabel metal2 s 2250 609 2316 661 4 dout_1
rlabel metal2 s 2473 538 2539 590 4 din_2
rlabel metal2 s 3418 609 3484 661 4 dout_2
rlabel metal2 s 3641 538 3707 590 4 din_3
rlabel metal2 s 4586 609 4652 661 4 dout_3
rlabel metal2 s 4809 538 4875 590 4 din_4
rlabel metal2 s 5754 609 5820 661 4 dout_4
rlabel metal2 s 5977 538 6043 590 4 din_5
rlabel metal2 s 6922 609 6988 661 4 dout_5
rlabel metal2 s 7145 538 7211 590 4 din_6
rlabel metal2 s 8090 609 8156 661 4 dout_6
rlabel metal2 s 8313 538 8379 590 4 din_7
rlabel metal2 s 9258 609 9324 661 4 dout_7
rlabel metal2 s 9481 538 9547 590 4 din_8
rlabel metal2 s 10426 609 10492 661 4 dout_8
rlabel metal2 s 10649 538 10715 590 4 din_9
rlabel metal2 s 11594 609 11660 661 4 dout_9
rlabel metal2 s 11817 538 11883 590 4 din_10
rlabel metal2 s 12762 609 12828 661 4 dout_10
rlabel metal2 s 12985 538 13051 590 4 din_11
rlabel metal2 s 13930 609 13996 661 4 dout_11
rlabel metal2 s 14153 538 14219 590 4 din_12
rlabel metal2 s 15098 609 15164 661 4 dout_12
rlabel metal2 s 15321 538 15387 590 4 din_13
rlabel metal2 s 16266 609 16332 661 4 dout_13
rlabel metal2 s 16489 538 16555 590 4 din_14
rlabel metal2 s 17434 609 17500 661 4 dout_14
rlabel metal2 s 17657 538 17723 590 4 din_15
rlabel metal2 s 18602 609 18668 661 4 dout_15
rlabel metal2 s 18825 538 18891 590 4 din_16
rlabel metal2 s 19770 609 19836 661 4 dout_16
rlabel metal2 s 19993 538 20059 590 4 din_17
rlabel metal2 s 20938 609 21004 661 4 dout_17
rlabel metal2 s 21161 538 21227 590 4 din_18
rlabel metal2 s 22106 609 22172 661 4 dout_18
rlabel metal2 s 22329 538 22395 590 4 din_19
rlabel metal2 s 23274 609 23340 661 4 dout_19
rlabel metal2 s 23497 538 23563 590 4 din_20
rlabel metal2 s 24442 609 24508 661 4 dout_20
rlabel metal2 s 24665 538 24731 590 4 din_21
rlabel metal2 s 25610 609 25676 661 4 dout_21
rlabel metal2 s 25833 538 25899 590 4 din_22
rlabel metal2 s 26778 609 26844 661 4 dout_22
rlabel metal2 s 27001 538 27067 590 4 din_23
rlabel metal2 s 27946 609 28012 661 4 dout_23
rlabel metal2 s 28169 538 28235 590 4 din_24
rlabel metal2 s 29114 609 29180 661 4 dout_24
rlabel metal2 s 29337 538 29403 590 4 din_25
rlabel metal2 s 30282 609 30348 661 4 dout_25
rlabel metal2 s 30505 538 30571 590 4 din_26
rlabel metal2 s 31450 609 31516 661 4 dout_26
rlabel metal2 s 31673 538 31739 590 4 din_27
rlabel metal2 s 32618 609 32684 661 4 dout_27
rlabel metal2 s 32841 538 32907 590 4 din_28
rlabel metal2 s 33786 609 33852 661 4 dout_28
rlabel metal2 s 34009 538 34075 590 4 din_29
rlabel metal2 s 34954 609 35020 661 4 dout_29
rlabel metal2 s 35177 538 35243 590 4 din_30
rlabel metal2 s 36122 609 36188 661 4 dout_30
rlabel metal2 s 36345 538 36411 590 4 din_31
rlabel metal2 s 37290 609 37356 661 4 dout_31
rlabel metal3 s 0 278 37376 338 4 clk
<< properties >>
string FIXED_BBOX 0 0 37376 1414
<< end >>
