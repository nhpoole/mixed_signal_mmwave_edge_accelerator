magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< nwell >>
rect -54 -54 420 390
<< scpmos >>
rect 60 0 90 336
rect 168 0 198 336
rect 276 0 306 336
<< pdiff >>
rect 0 0 60 336
rect 90 0 168 336
rect 198 0 276 336
rect 306 0 366 336
<< poly >>
rect 60 336 90 362
rect 168 336 198 362
rect 276 336 306 362
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 60 -56 306 -26
<< locali >>
rect 8 135 42 201
rect 112 101 146 168
rect 220 135 254 201
rect 324 101 358 168
rect 112 67 358 101
use contact_12  contact_12_0
timestamp 1624494425
transform 1 0 316 0 1 135
box -59 -51 109 117
use contact_12  contact_12_1
timestamp 1624494425
transform 1 0 212 0 1 135
box -59 -51 109 117
use contact_12  contact_12_2
timestamp 1624494425
transform 1 0 104 0 1 135
box -59 -51 109 117
use contact_12  contact_12_3
timestamp 1624494425
transform 1 0 0 0 1 135
box -59 -51 109 117
<< labels >>
rlabel poly s 183 -41 183 -41 4 G
rlabel locali s 25 168 25 168 4 S
rlabel locali s 237 168 237 168 4 S
rlabel locali s 235 84 235 84 4 D
<< properties >>
string FIXED_BBOX -54 -56 420 390
<< end >>
