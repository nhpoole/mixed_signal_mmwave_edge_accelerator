magic
tech sky130A
magscale 1 2
timestamp 1622257752
<< nwell >>
rect -941 -419 941 419
<< pmoshvt >>
rect -745 -200 -545 200
rect -487 -200 -287 200
rect -229 -200 -29 200
rect 29 -200 229 200
rect 287 -200 487 200
rect 545 -200 745 200
<< pdiff >>
rect -803 188 -745 200
rect -803 -188 -791 188
rect -757 -188 -745 188
rect -803 -200 -745 -188
rect -545 188 -487 200
rect -545 -188 -533 188
rect -499 -188 -487 188
rect -545 -200 -487 -188
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
rect 487 188 545 200
rect 487 -188 499 188
rect 533 -188 545 188
rect 487 -200 545 -188
rect 745 188 803 200
rect 745 -188 757 188
rect 791 -188 803 188
rect 745 -200 803 -188
<< pdiffc >>
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
<< nsubdiff >>
rect -905 349 -809 383
rect 809 349 905 383
rect -905 287 -871 349
rect 871 287 905 349
rect -905 -349 -871 -287
rect 871 -349 905 -287
rect -905 -383 -809 -349
rect 809 -383 905 -349
<< nsubdiffcont >>
rect -809 349 809 383
rect -905 -287 -871 287
rect 871 -287 905 287
rect -809 -383 809 -349
<< poly >>
rect -711 281 -579 297
rect -711 264 -695 281
rect -745 247 -695 264
rect -595 264 -579 281
rect -453 281 -321 297
rect -453 264 -437 281
rect -595 247 -545 264
rect -745 200 -545 247
rect -487 247 -437 264
rect -337 264 -321 281
rect -195 281 -63 297
rect -195 264 -179 281
rect -337 247 -287 264
rect -487 200 -287 247
rect -229 247 -179 264
rect -79 264 -63 281
rect 63 281 195 297
rect 63 264 79 281
rect -79 247 -29 264
rect -229 200 -29 247
rect 29 247 79 264
rect 179 264 195 281
rect 321 281 453 297
rect 321 264 337 281
rect 179 247 229 264
rect 29 200 229 247
rect 287 247 337 264
rect 437 264 453 281
rect 579 281 711 297
rect 579 264 595 281
rect 437 247 487 264
rect 287 200 487 247
rect 545 247 595 264
rect 695 264 711 281
rect 695 247 745 264
rect 545 200 745 247
rect -745 -247 -545 -200
rect -745 -264 -695 -247
rect -711 -281 -695 -264
rect -595 -264 -545 -247
rect -487 -247 -287 -200
rect -487 -264 -437 -247
rect -595 -281 -579 -264
rect -711 -297 -579 -281
rect -453 -281 -437 -264
rect -337 -264 -287 -247
rect -229 -247 -29 -200
rect -229 -264 -179 -247
rect -337 -281 -321 -264
rect -453 -297 -321 -281
rect -195 -281 -179 -264
rect -79 -264 -29 -247
rect 29 -247 229 -200
rect 29 -264 79 -247
rect -79 -281 -63 -264
rect -195 -297 -63 -281
rect 63 -281 79 -264
rect 179 -264 229 -247
rect 287 -247 487 -200
rect 287 -264 337 -247
rect 179 -281 195 -264
rect 63 -297 195 -281
rect 321 -281 337 -264
rect 437 -264 487 -247
rect 545 -247 745 -200
rect 545 -264 595 -247
rect 437 -281 453 -264
rect 321 -297 453 -281
rect 579 -281 595 -264
rect 695 -264 745 -247
rect 695 -281 711 -264
rect 579 -297 711 -281
<< polycont >>
rect -695 247 -595 281
rect -437 247 -337 281
rect -179 247 -79 281
rect 79 247 179 281
rect 337 247 437 281
rect 595 247 695 281
rect -695 -281 -595 -247
rect -437 -281 -337 -247
rect -179 -281 -79 -247
rect 79 -281 179 -247
rect 337 -281 437 -247
rect 595 -281 695 -247
<< locali >>
rect -905 349 -809 383
rect 809 349 905 383
rect -905 287 -871 349
rect 871 287 905 349
rect -711 247 -695 281
rect -595 247 -579 281
rect -453 247 -437 281
rect -337 247 -321 281
rect -195 247 -179 281
rect -79 247 -63 281
rect 63 247 79 281
rect 179 247 195 281
rect 321 247 337 281
rect 437 247 453 281
rect 579 247 595 281
rect 695 247 711 281
rect -791 188 -757 204
rect -791 -204 -757 -188
rect -533 188 -499 204
rect -533 -204 -499 -188
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect 499 188 533 204
rect 499 -204 533 -188
rect 757 188 791 204
rect 757 -204 791 -188
rect -711 -281 -695 -247
rect -595 -281 -579 -247
rect -453 -281 -437 -247
rect -337 -281 -321 -247
rect -195 -281 -179 -247
rect -79 -281 -63 -247
rect 63 -281 79 -247
rect 179 -281 195 -247
rect 321 -281 337 -247
rect 437 -281 453 -247
rect 579 -281 595 -247
rect 695 -281 711 -247
rect -905 -349 -871 -287
rect 871 -349 905 -287
rect -905 -383 -809 -349
rect 809 -383 905 -349
<< viali >>
rect -687 247 -603 281
rect -429 247 -345 281
rect -171 247 -87 281
rect 87 247 171 281
rect 345 247 429 281
rect 603 247 687 281
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect -687 -281 -603 -247
rect -429 -281 -345 -247
rect -171 -281 -87 -247
rect 87 -281 171 -247
rect 345 -281 429 -247
rect 603 -281 687 -247
<< metal1 >>
rect -699 281 -591 287
rect -699 247 -687 281
rect -603 247 -591 281
rect -699 241 -591 247
rect -441 281 -333 287
rect -441 247 -429 281
rect -345 247 -333 281
rect -441 241 -333 247
rect -183 281 -75 287
rect -183 247 -171 281
rect -87 247 -75 281
rect -183 241 -75 247
rect 75 281 183 287
rect 75 247 87 281
rect 171 247 183 281
rect 75 241 183 247
rect 333 281 441 287
rect 333 247 345 281
rect 429 247 441 281
rect 333 241 441 247
rect 591 281 699 287
rect 591 247 603 281
rect 687 247 699 281
rect 591 241 699 247
rect -797 188 -751 200
rect -797 -188 -791 188
rect -757 -188 -751 188
rect -797 -200 -751 -188
rect -539 188 -493 200
rect -539 -188 -533 188
rect -499 -188 -493 188
rect -539 -200 -493 -188
rect -281 188 -235 200
rect -281 -188 -275 188
rect -241 -188 -235 188
rect -281 -200 -235 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 235 188 281 200
rect 235 -188 241 188
rect 275 -188 281 188
rect 235 -200 281 -188
rect 493 188 539 200
rect 493 -188 499 188
rect 533 -188 539 188
rect 493 -200 539 -188
rect 751 188 797 200
rect 751 -188 757 188
rect 791 -188 797 188
rect 751 -200 797 -188
rect -699 -247 -591 -241
rect -699 -281 -687 -247
rect -603 -281 -591 -247
rect -699 -287 -591 -281
rect -441 -247 -333 -241
rect -441 -281 -429 -247
rect -345 -281 -333 -247
rect -441 -287 -333 -281
rect -183 -247 -75 -241
rect -183 -281 -171 -247
rect -87 -281 -75 -247
rect -183 -287 -75 -281
rect 75 -247 183 -241
rect 75 -281 87 -247
rect 171 -281 183 -247
rect 75 -287 183 -281
rect 333 -247 441 -241
rect 333 -281 345 -247
rect 429 -281 441 -247
rect 333 -287 441 -281
rect 591 -247 699 -241
rect 591 -281 603 -247
rect 687 -281 699 -247
rect 591 -287 699 -281
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_hvt
string FIXED_BBOX -888 -366 888 366
string parameters w 2 l 1 m 1 nf 6 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
