magic
tech sky130A
timestamp 1626065694
<< checkpaint >>
rect -798 -654 798 654
<< metal1 >>
rect -168 13 168 24
rect -168 -13 -157 13
rect -131 -13 -125 13
rect -99 -13 -93 13
rect -67 -13 -61 13
rect -35 -13 -29 13
rect -3 -13 3 13
rect 29 -13 35 13
rect 61 -13 67 13
rect 93 -13 99 13
rect 125 -13 131 13
rect 157 -13 168 13
rect -168 -24 168 -13
<< via1 >>
rect -157 -13 -131 13
rect -125 -13 -99 13
rect -93 -13 -67 13
rect -61 -13 -35 13
rect -29 -13 -3 13
rect 3 -13 29 13
rect 35 -13 61 13
rect 67 -13 93 13
rect 99 -13 125 13
rect 131 -13 157 13
<< metal2 >>
rect -168 13 168 24
rect -168 -13 -157 13
rect -131 -13 -125 13
rect -99 -13 -93 13
rect -67 -13 -61 13
rect -35 -13 -29 13
rect -3 -13 3 13
rect 29 -13 35 13
rect 61 -13 67 13
rect 93 -13 99 13
rect 125 -13 131 13
rect 157 -13 168 13
rect -168 -24 168 -13
<< end >>
