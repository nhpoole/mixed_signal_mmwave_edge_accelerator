magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect 72925 56100 77802 60376
<< nwell >>
rect 74185 58186 76094 59026
<< locali >>
rect 74267 58956 74288 58990
rect 74322 58956 74360 58990
rect 74394 58956 74432 58990
rect 74466 58956 74487 58990
rect 75759 58956 75771 58990
rect 75805 58956 75843 58990
rect 75877 58956 75915 58990
rect 75949 58956 75961 58990
rect 74219 58875 74257 58892
rect 74219 58841 74221 58875
rect 74255 58841 74257 58875
rect 74219 58803 74257 58841
rect 74219 58769 74221 58803
rect 74255 58769 74257 58803
rect 74219 58731 74257 58769
rect 74219 58697 74221 58731
rect 74255 58697 74257 58731
rect 74219 58659 74257 58697
rect 74219 58625 74221 58659
rect 74255 58625 74257 58659
rect 74219 58587 74257 58625
rect 74219 58553 74221 58587
rect 74255 58553 74257 58587
rect 74219 58515 74257 58553
rect 74219 58481 74221 58515
rect 74255 58481 74257 58515
rect 74219 58443 74257 58481
rect 74219 58409 74221 58443
rect 74255 58409 74257 58443
rect 74219 58371 74257 58409
rect 74219 58337 74221 58371
rect 74255 58337 74257 58371
rect 74219 58320 74257 58337
rect 75995 58875 76031 58894
rect 75995 58841 75996 58875
rect 76030 58841 76031 58875
rect 75995 58803 76031 58841
rect 75995 58769 75996 58803
rect 76030 58769 76031 58803
rect 75995 58731 76031 58769
rect 75995 58697 75996 58731
rect 76030 58697 76031 58731
rect 75995 58659 76031 58697
rect 75995 58625 75996 58659
rect 76030 58625 76031 58659
rect 75995 58587 76031 58625
rect 75995 58553 75996 58587
rect 76030 58553 76031 58587
rect 75995 58515 76031 58553
rect 75995 58481 75996 58515
rect 76030 58481 76031 58515
rect 75995 58443 76031 58481
rect 75995 58409 75996 58443
rect 76030 58409 76031 58443
rect 75995 58371 76031 58409
rect 75995 58337 75996 58371
rect 76030 58337 76031 58371
rect 75995 58318 76031 58337
rect 74267 58222 74288 58256
rect 74322 58222 74360 58256
rect 74394 58222 74432 58256
rect 74466 58222 74487 58256
rect 75759 58224 75771 58258
rect 75805 58224 75843 58258
rect 75877 58224 75915 58258
rect 75949 58224 75961 58258
rect 76268 58183 76314 58186
rect 76164 58157 76212 58164
rect 76164 58123 76171 58157
rect 76205 58123 76212 58157
rect 76268 58149 76274 58183
rect 76308 58149 76314 58183
rect 76268 58146 76314 58149
rect 76164 58116 76212 58123
rect 75763 58058 75961 58060
rect 74291 58056 74499 58058
rect 74291 58022 74306 58056
rect 74340 58022 74378 58056
rect 74412 58022 74450 58056
rect 74484 58022 74499 58056
rect 75763 58024 75773 58058
rect 75807 58024 75845 58058
rect 75879 58024 75917 58058
rect 75951 58024 75961 58058
rect 75763 58022 75961 58024
rect 74291 58020 74499 58022
rect 74219 57943 74255 57960
rect 74219 57909 74220 57943
rect 74254 57909 74255 57943
rect 74219 57871 74255 57909
rect 74219 57837 74220 57871
rect 74254 57837 74255 57871
rect 74219 57799 74255 57837
rect 74219 57765 74220 57799
rect 74254 57765 74255 57799
rect 74219 57727 74255 57765
rect 74219 57693 74220 57727
rect 74254 57693 74255 57727
rect 74219 57655 74255 57693
rect 74219 57621 74220 57655
rect 74254 57621 74255 57655
rect 74219 57604 74255 57621
rect 75995 57943 76033 57960
rect 75995 57909 75997 57943
rect 76031 57909 76033 57943
rect 75995 57871 76033 57909
rect 75995 57837 75997 57871
rect 76031 57837 76033 57871
rect 75995 57799 76033 57837
rect 75995 57765 75997 57799
rect 76031 57765 76033 57799
rect 75995 57727 76033 57765
rect 75995 57693 75997 57727
rect 76031 57693 76033 57727
rect 75995 57655 76033 57693
rect 75995 57621 75997 57655
rect 76031 57621 76033 57655
rect 75995 57604 76033 57621
rect 74289 57543 74497 57544
rect 74289 57509 74304 57543
rect 74338 57509 74376 57543
rect 74410 57509 74448 57543
rect 74482 57509 74497 57543
rect 74289 57508 74497 57509
rect 75761 57541 75963 57542
rect 75761 57507 75773 57541
rect 75807 57507 75845 57541
rect 75879 57507 75917 57541
rect 75951 57507 75963 57541
rect 75761 57506 75963 57507
<< viali >>
rect 74288 58956 74322 58990
rect 74360 58956 74394 58990
rect 74432 58956 74466 58990
rect 75771 58956 75805 58990
rect 75843 58956 75877 58990
rect 75915 58956 75949 58990
rect 74221 58841 74255 58875
rect 74221 58769 74255 58803
rect 74221 58697 74255 58731
rect 74221 58625 74255 58659
rect 74221 58553 74255 58587
rect 74221 58481 74255 58515
rect 74221 58409 74255 58443
rect 74221 58337 74255 58371
rect 75996 58841 76030 58875
rect 75996 58769 76030 58803
rect 75996 58697 76030 58731
rect 75996 58625 76030 58659
rect 75996 58553 76030 58587
rect 75996 58481 76030 58515
rect 75996 58409 76030 58443
rect 75996 58337 76030 58371
rect 74288 58222 74322 58256
rect 74360 58222 74394 58256
rect 74432 58222 74466 58256
rect 75771 58224 75805 58258
rect 75843 58224 75877 58258
rect 75915 58224 75949 58258
rect 76171 58123 76205 58157
rect 76274 58149 76308 58183
rect 74306 58022 74340 58056
rect 74378 58022 74412 58056
rect 74450 58022 74484 58056
rect 75773 58024 75807 58058
rect 75845 58024 75879 58058
rect 75917 58024 75951 58058
rect 74220 57909 74254 57943
rect 74220 57837 74254 57871
rect 74220 57765 74254 57799
rect 74220 57693 74254 57727
rect 74220 57621 74254 57655
rect 75997 57909 76031 57943
rect 75997 57837 76031 57871
rect 75997 57765 76031 57799
rect 75997 57693 76031 57727
rect 75997 57621 76031 57655
rect 74304 57509 74338 57543
rect 74376 57509 74410 57543
rect 74448 57509 74482 57543
rect 75773 57507 75807 57541
rect 75845 57507 75879 57541
rect 75917 57507 75951 57541
<< metal1 >>
rect 74208 59056 76044 59116
rect 74208 58990 74513 59056
rect 74208 58956 74288 58990
rect 74322 58956 74360 58990
rect 74394 58956 74432 58990
rect 74466 58956 74513 58990
rect 74208 58942 74513 58956
rect 74208 58875 74269 58942
rect 74208 58862 74221 58875
rect 74209 58841 74221 58862
rect 74255 58841 74269 58875
rect 74209 58803 74269 58841
rect 74209 58769 74221 58803
rect 74255 58769 74269 58803
rect 74209 58731 74269 58769
rect 74209 58697 74221 58731
rect 74255 58697 74269 58731
rect 74209 58659 74269 58697
rect 74209 58634 74221 58659
rect 74208 58625 74221 58634
rect 74255 58634 74269 58659
rect 74319 58634 74379 58942
rect 74453 58851 74513 58942
rect 74709 59008 74769 59009
rect 75485 59008 75545 59014
rect 74709 59004 75545 59008
rect 74709 58952 75489 59004
rect 75541 58952 75545 59004
rect 74709 58948 75545 58952
rect 74709 58853 74769 58948
rect 74967 58851 75027 58948
rect 75225 58853 75285 58948
rect 75485 58853 75545 58948
rect 75741 58990 76044 59056
rect 75741 58956 75771 58990
rect 75805 58956 75843 58990
rect 75877 58956 75915 58990
rect 75949 58956 76044 58990
rect 75741 58942 76044 58956
rect 75741 58851 75801 58942
rect 74255 58625 74379 58634
rect 74208 58587 74379 58625
rect 74208 58574 74221 58587
rect 74209 58553 74221 58574
rect 74255 58574 74379 58587
rect 75869 58636 75929 58942
rect 75983 58878 76044 58942
rect 75983 58875 76043 58878
rect 75983 58841 75996 58875
rect 76030 58841 76043 58875
rect 75983 58803 76043 58841
rect 75983 58769 75996 58803
rect 76030 58769 76043 58803
rect 75983 58731 76043 58769
rect 75983 58697 75996 58731
rect 76030 58697 76043 58731
rect 75983 58659 76043 58697
rect 75983 58636 75996 58659
rect 75869 58625 75996 58636
rect 76030 58625 76043 58659
rect 75869 58587 76043 58625
rect 75869 58576 75996 58587
rect 74255 58553 74269 58574
rect 74209 58515 74269 58553
rect 74209 58481 74221 58515
rect 74255 58481 74269 58515
rect 74209 58443 74269 58481
rect 75983 58553 75996 58576
rect 76030 58553 76043 58587
rect 75983 58518 76043 58553
rect 75983 58515 76144 58518
rect 75983 58481 75996 58515
rect 76030 58481 76144 58515
rect 74209 58409 74221 58443
rect 74255 58409 74269 58443
rect 74209 58371 74269 58409
rect 74209 58337 74221 58371
rect 74255 58337 74269 58371
rect 74209 58270 74269 58337
rect 74321 58270 74381 58452
rect 74449 58270 74509 58358
rect 74208 58256 74509 58270
rect 74208 58222 74288 58256
rect 74322 58222 74360 58256
rect 74394 58222 74432 58256
rect 74466 58222 74509 58256
rect 74208 58210 74509 58222
rect 74579 58093 74639 58463
rect 74837 58242 74897 58438
rect 74831 58238 74903 58242
rect 74831 58186 74841 58238
rect 74893 58186 74903 58238
rect 74831 58182 74903 58186
rect 74573 58089 74645 58093
rect 74207 58056 74511 58068
rect 74207 58022 74306 58056
rect 74340 58022 74378 58056
rect 74412 58022 74450 58056
rect 74484 58022 74511 58056
rect 74573 58037 74583 58089
rect 74635 58037 74645 58089
rect 74573 58033 74645 58037
rect 74207 58008 74511 58022
rect 74207 57943 74267 58008
rect 74207 57909 74220 57943
rect 74254 57909 74267 57943
rect 74207 57871 74267 57909
rect 74207 57837 74220 57871
rect 74254 57837 74267 57871
rect 74207 57799 74267 57837
rect 74321 57820 74381 58008
rect 74451 57920 74511 58008
rect 74579 57833 74639 58033
rect 74837 57900 74897 58182
rect 75095 58093 75155 58461
rect 75355 58242 75415 58456
rect 75349 58238 75421 58242
rect 75349 58186 75359 58238
rect 75411 58186 75421 58238
rect 75349 58182 75421 58186
rect 75089 58089 75161 58093
rect 75089 58037 75099 58089
rect 75151 58037 75161 58089
rect 75089 58033 75161 58037
rect 74837 57834 74899 57900
rect 74207 57765 74220 57799
rect 74254 57765 74267 57799
rect 74207 57727 74267 57765
rect 74207 57693 74220 57727
rect 74254 57693 74267 57727
rect 74207 57655 74267 57693
rect 74207 57621 74220 57655
rect 74254 57621 74267 57655
rect 74207 57555 74267 57621
rect 74323 57555 74383 57733
rect 74839 57654 74899 57834
rect 75095 57714 75155 58033
rect 75355 57654 75415 58182
rect 75613 58089 75673 58461
rect 75737 58270 75797 58358
rect 75871 58270 75931 58448
rect 75983 58443 76144 58481
rect 75983 58409 75996 58443
rect 76030 58422 76144 58443
rect 76030 58409 76043 58422
rect 75983 58371 76043 58409
rect 75983 58337 75996 58371
rect 76030 58337 76043 58371
rect 75983 58270 76043 58337
rect 75737 58258 76043 58270
rect 75737 58224 75771 58258
rect 75805 58224 75843 58258
rect 75877 58224 75915 58258
rect 75949 58224 76043 58258
rect 75737 58210 76043 58224
rect 76476 58192 76536 58198
rect 76256 58188 76536 58192
rect 76256 58183 76480 58188
rect 76158 58170 76218 58176
rect 76152 58166 76224 58170
rect 76152 58114 76162 58166
rect 76214 58114 76224 58166
rect 76256 58149 76274 58183
rect 76308 58149 76480 58183
rect 76256 58136 76480 58149
rect 76532 58136 76536 58188
rect 76256 58132 76536 58136
rect 76476 58126 76536 58132
rect 76152 58110 76224 58114
rect 76158 58104 76218 58110
rect 75613 58037 75617 58089
rect 75669 58037 75673 58089
rect 75613 57831 75673 58037
rect 75743 58058 76045 58070
rect 75743 58024 75773 58058
rect 75807 58024 75845 58058
rect 75879 58024 75917 58058
rect 75951 58024 76045 58058
rect 75743 58010 76045 58024
rect 75743 57922 75803 58010
rect 75871 57824 75931 58010
rect 75985 57974 76045 58010
rect 75985 57943 76136 57974
rect 75985 57909 75997 57943
rect 76031 57909 76136 57943
rect 75985 57878 76136 57909
rect 75985 57871 76045 57878
rect 75985 57837 75997 57871
rect 76031 57837 76045 57871
rect 75985 57799 76045 57837
rect 75985 57765 75997 57799
rect 76031 57765 76045 57799
rect 75985 57727 76045 57765
rect 74451 57555 74511 57644
rect 74207 57543 74511 57555
rect 74207 57509 74304 57543
rect 74338 57509 74376 57543
rect 74410 57509 74448 57543
rect 74482 57509 74511 57543
rect 74207 57438 74511 57509
rect 74709 57545 74769 57645
rect 74969 57545 75029 57645
rect 75227 57545 75287 57643
rect 75483 57545 75543 57643
rect 75741 57555 75801 57646
rect 75869 57555 75929 57727
rect 75985 57693 75997 57727
rect 76031 57693 76045 57727
rect 75985 57655 76045 57693
rect 75985 57621 75997 57655
rect 76031 57621 76045 57655
rect 75985 57555 76045 57621
rect 74709 57541 75549 57545
rect 74709 57489 75487 57541
rect 75539 57489 75549 57541
rect 74709 57485 75549 57489
rect 75741 57541 76045 57555
rect 75741 57507 75773 57541
rect 75807 57507 75845 57541
rect 75879 57507 75917 57541
rect 75951 57507 76045 57541
rect 74208 57420 74511 57438
rect 75741 57420 76045 57507
rect 74208 57360 76046 57420
<< via1 >>
rect 75489 58952 75541 59004
rect 74841 58186 74893 58238
rect 74583 58037 74635 58089
rect 75359 58186 75411 58238
rect 75099 58037 75151 58089
rect 76162 58157 76214 58166
rect 76162 58123 76171 58157
rect 76171 58123 76205 58157
rect 76205 58123 76214 58157
rect 76162 58114 76214 58123
rect 76480 58136 76532 58188
rect 75617 58037 75669 58089
rect 75487 57489 75539 57541
<< metal2 >>
rect 75479 59004 76144 59008
rect 75479 58952 75489 59004
rect 75541 58952 76144 59004
rect 75479 58948 76144 58952
rect 74837 58242 74897 58248
rect 75355 58242 75415 58248
rect 74837 58238 75415 58242
rect 74837 58186 74841 58238
rect 74893 58186 75359 58238
rect 75411 58186 75415 58238
rect 74837 58182 75415 58186
rect 74837 58176 74897 58182
rect 75355 58176 75415 58182
rect 76084 58170 76144 58948
rect 76470 58188 76542 58192
rect 76084 58166 76224 58170
rect 76084 58114 76162 58166
rect 76214 58114 76224 58166
rect 76470 58136 76480 58188
rect 76532 58136 76542 58188
rect 76470 58132 76542 58136
rect 76084 58110 76224 58114
rect 74579 58093 74639 58099
rect 75095 58093 75155 58099
rect 74568 58089 75679 58093
rect 74568 58037 74583 58089
rect 74635 58037 75099 58089
rect 75151 58037 75617 58089
rect 75669 58037 75679 58089
rect 74568 58033 75679 58037
rect 74579 58027 74639 58033
rect 75095 58027 75155 58033
rect 75483 57545 75543 57551
rect 76476 57546 76536 58132
rect 75990 57545 76536 57546
rect 75483 57541 76536 57545
rect 75483 57489 75487 57541
rect 75539 57489 76536 57541
rect 75483 57486 76536 57489
rect 75483 57485 76094 57486
rect 75483 57479 75543 57485
use sky130_fd_pr__pfet_01v8_hvt_SCHXZ7  sky130_fd_pr__pfet_01v8_hvt_SCHXZ7_0
timestamp 1626486988
transform 1 0 75126 0 1 58606
box -941 -419 941 419
use sky130_fd_pr__nfet_01v8_N6QVV6  sky130_fd_pr__nfet_01v8_N6QVV6_0
timestamp 1626486988
transform 1 0 75126 0 1 57782
box -931 -300 931 300
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1626486988
transform -1 0 76381 0 1 57926
box -38 -48 314 592
<< labels >>
flabel metal1 s 76416 58154 76424 58160 1 FreeSans 600 0 0 0 tx
flabel metal1 s 74598 58134 74608 58142 1 FreeSans 600 0 0 0 out
flabel metal1 s 74860 58140 74870 58148 1 FreeSans 600 0 0 0 in
flabel metal1 s 75114 59082 75124 59092 1 FreeSans 600 0 0 0 VDD
flabel metal1 s 75112 57392 75120 57398 1 FreeSans 600 0 0 0 VSS
flabel metal2 s 76114 58656 76124 58664 1 FreeSans 600 0 0 0 txb
<< end >>
