magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< pwell >>
rect -26 -26 4712 426
<< scnmos >>
rect 60 0 90 400
rect 168 0 198 400
rect 276 0 306 400
rect 384 0 414 400
rect 492 0 522 400
rect 600 0 630 400
rect 708 0 738 400
rect 816 0 846 400
rect 924 0 954 400
rect 1032 0 1062 400
rect 1140 0 1170 400
rect 1248 0 1278 400
rect 1356 0 1386 400
rect 1464 0 1494 400
rect 1572 0 1602 400
rect 1680 0 1710 400
rect 1788 0 1818 400
rect 1896 0 1926 400
rect 2004 0 2034 400
rect 2112 0 2142 400
rect 2220 0 2250 400
rect 2328 0 2358 400
rect 2436 0 2466 400
rect 2544 0 2574 400
rect 2652 0 2682 400
rect 2760 0 2790 400
rect 2868 0 2898 400
rect 2976 0 3006 400
rect 3084 0 3114 400
rect 3192 0 3222 400
rect 3300 0 3330 400
rect 3408 0 3438 400
rect 3516 0 3546 400
rect 3624 0 3654 400
rect 3732 0 3762 400
rect 3840 0 3870 400
rect 3948 0 3978 400
rect 4056 0 4086 400
rect 4164 0 4194 400
rect 4272 0 4302 400
rect 4380 0 4410 400
rect 4488 0 4518 400
rect 4596 0 4626 400
<< ndiff >>
rect 0 0 60 400
rect 90 0 168 400
rect 198 0 276 400
rect 306 0 384 400
rect 414 0 492 400
rect 522 0 600 400
rect 630 0 708 400
rect 738 0 816 400
rect 846 0 924 400
rect 954 0 1032 400
rect 1062 0 1140 400
rect 1170 0 1248 400
rect 1278 0 1356 400
rect 1386 0 1464 400
rect 1494 0 1572 400
rect 1602 0 1680 400
rect 1710 0 1788 400
rect 1818 0 1896 400
rect 1926 0 2004 400
rect 2034 0 2112 400
rect 2142 0 2220 400
rect 2250 0 2328 400
rect 2358 0 2436 400
rect 2466 0 2544 400
rect 2574 0 2652 400
rect 2682 0 2760 400
rect 2790 0 2868 400
rect 2898 0 2976 400
rect 3006 0 3084 400
rect 3114 0 3192 400
rect 3222 0 3300 400
rect 3330 0 3408 400
rect 3438 0 3516 400
rect 3546 0 3624 400
rect 3654 0 3732 400
rect 3762 0 3840 400
rect 3870 0 3948 400
rect 3978 0 4056 400
rect 4086 0 4164 400
rect 4194 0 4272 400
rect 4302 0 4380 400
rect 4410 0 4488 400
rect 4518 0 4596 400
rect 4626 0 4686 400
<< poly >>
rect 60 426 4626 456
rect 60 400 90 426
rect 168 400 198 426
rect 276 400 306 426
rect 384 400 414 426
rect 492 400 522 426
rect 600 400 630 426
rect 708 400 738 426
rect 816 400 846 426
rect 924 400 954 426
rect 1032 400 1062 426
rect 1140 400 1170 426
rect 1248 400 1278 426
rect 1356 400 1386 426
rect 1464 400 1494 426
rect 1572 400 1602 426
rect 1680 400 1710 426
rect 1788 400 1818 426
rect 1896 400 1926 426
rect 2004 400 2034 426
rect 2112 400 2142 426
rect 2220 400 2250 426
rect 2328 400 2358 426
rect 2436 400 2466 426
rect 2544 400 2574 426
rect 2652 400 2682 426
rect 2760 400 2790 426
rect 2868 400 2898 426
rect 2976 400 3006 426
rect 3084 400 3114 426
rect 3192 400 3222 426
rect 3300 400 3330 426
rect 3408 400 3438 426
rect 3516 400 3546 426
rect 3624 400 3654 426
rect 3732 400 3762 426
rect 3840 400 3870 426
rect 3948 400 3978 426
rect 4056 400 4086 426
rect 4164 400 4194 426
rect 4272 400 4302 426
rect 4380 400 4410 426
rect 4488 400 4518 426
rect 4596 400 4626 426
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
rect 1032 -26 1062 0
rect 1140 -26 1170 0
rect 1248 -26 1278 0
rect 1356 -26 1386 0
rect 1464 -26 1494 0
rect 1572 -26 1602 0
rect 1680 -26 1710 0
rect 1788 -26 1818 0
rect 1896 -26 1926 0
rect 2004 -26 2034 0
rect 2112 -26 2142 0
rect 2220 -26 2250 0
rect 2328 -26 2358 0
rect 2436 -26 2466 0
rect 2544 -26 2574 0
rect 2652 -26 2682 0
rect 2760 -26 2790 0
rect 2868 -26 2898 0
rect 2976 -26 3006 0
rect 3084 -26 3114 0
rect 3192 -26 3222 0
rect 3300 -26 3330 0
rect 3408 -26 3438 0
rect 3516 -26 3546 0
rect 3624 -26 3654 0
rect 3732 -26 3762 0
rect 3840 -26 3870 0
rect 3948 -26 3978 0
rect 4056 -26 4086 0
rect 4164 -26 4194 0
rect 4272 -26 4302 0
rect 4380 -26 4410 0
rect 4488 -26 4518 0
rect 4596 -26 4626 0
<< locali >>
rect 112 267 4678 301
rect 8 167 42 233
rect 112 200 146 267
rect 220 167 254 233
rect 328 200 362 267
rect 436 167 470 233
rect 544 200 578 267
rect 652 167 686 233
rect 760 200 794 267
rect 868 167 902 233
rect 976 200 1010 267
rect 1084 167 1118 233
rect 1192 200 1226 267
rect 1300 167 1334 233
rect 1408 200 1442 267
rect 1516 167 1550 233
rect 1624 200 1658 267
rect 1732 167 1766 233
rect 1840 200 1874 267
rect 1948 167 1982 233
rect 2056 200 2090 267
rect 2164 167 2198 233
rect 2272 200 2306 267
rect 2380 167 2414 233
rect 2488 200 2522 267
rect 2596 167 2630 233
rect 2704 200 2738 267
rect 2812 167 2846 233
rect 2920 200 2954 267
rect 3028 167 3062 233
rect 3136 200 3170 267
rect 3244 167 3278 233
rect 3352 200 3386 267
rect 3460 167 3494 233
rect 3568 200 3602 267
rect 3676 167 3710 233
rect 3784 200 3818 267
rect 3892 167 3926 233
rect 4000 200 4034 267
rect 4108 167 4142 233
rect 4216 200 4250 267
rect 4324 167 4358 233
rect 4432 200 4466 267
rect 4540 167 4574 233
rect 4644 200 4678 267
use contact_11  contact_11_42
timestamp 1624494425
transform 1 0 104 0 1 167
box -26 -22 76 88
use contact_11  contact_11_43
timestamp 1624494425
transform 1 0 0 0 1 167
box -26 -22 76 88
use contact_11  contact_11_41
timestamp 1624494425
transform 1 0 212 0 1 167
box -26 -22 76 88
use contact_11  contact_11_40
timestamp 1624494425
transform 1 0 320 0 1 167
box -26 -22 76 88
use contact_11  contact_11_39
timestamp 1624494425
transform 1 0 428 0 1 167
box -26 -22 76 88
use contact_11  contact_11_38
timestamp 1624494425
transform 1 0 536 0 1 167
box -26 -22 76 88
use contact_11  contact_11_37
timestamp 1624494425
transform 1 0 644 0 1 167
box -26 -22 76 88
use contact_11  contact_11_36
timestamp 1624494425
transform 1 0 752 0 1 167
box -26 -22 76 88
use contact_11  contact_11_35
timestamp 1624494425
transform 1 0 860 0 1 167
box -26 -22 76 88
use contact_11  contact_11_34
timestamp 1624494425
transform 1 0 968 0 1 167
box -26 -22 76 88
use contact_11  contact_11_33
timestamp 1624494425
transform 1 0 1076 0 1 167
box -26 -22 76 88
use contact_11  contact_11_32
timestamp 1624494425
transform 1 0 1184 0 1 167
box -26 -22 76 88
use contact_11  contact_11_31
timestamp 1624494425
transform 1 0 1292 0 1 167
box -26 -22 76 88
use contact_11  contact_11_30
timestamp 1624494425
transform 1 0 1400 0 1 167
box -26 -22 76 88
use contact_11  contact_11_29
timestamp 1624494425
transform 1 0 1508 0 1 167
box -26 -22 76 88
use contact_11  contact_11_28
timestamp 1624494425
transform 1 0 1616 0 1 167
box -26 -22 76 88
use contact_11  contact_11_27
timestamp 1624494425
transform 1 0 1724 0 1 167
box -26 -22 76 88
use contact_11  contact_11_26
timestamp 1624494425
transform 1 0 1832 0 1 167
box -26 -22 76 88
use contact_11  contact_11_25
timestamp 1624494425
transform 1 0 1940 0 1 167
box -26 -22 76 88
use contact_11  contact_11_24
timestamp 1624494425
transform 1 0 2048 0 1 167
box -26 -22 76 88
use contact_11  contact_11_23
timestamp 1624494425
transform 1 0 2156 0 1 167
box -26 -22 76 88
use contact_11  contact_11_22
timestamp 1624494425
transform 1 0 2264 0 1 167
box -26 -22 76 88
use contact_11  contact_11_21
timestamp 1624494425
transform 1 0 2372 0 1 167
box -26 -22 76 88
use contact_11  contact_11_20
timestamp 1624494425
transform 1 0 2480 0 1 167
box -26 -22 76 88
use contact_11  contact_11_19
timestamp 1624494425
transform 1 0 2588 0 1 167
box -26 -22 76 88
use contact_11  contact_11_18
timestamp 1624494425
transform 1 0 2696 0 1 167
box -26 -22 76 88
use contact_11  contact_11_17
timestamp 1624494425
transform 1 0 2804 0 1 167
box -26 -22 76 88
use contact_11  contact_11_16
timestamp 1624494425
transform 1 0 2912 0 1 167
box -26 -22 76 88
use contact_11  contact_11_15
timestamp 1624494425
transform 1 0 3020 0 1 167
box -26 -22 76 88
use contact_11  contact_11_14
timestamp 1624494425
transform 1 0 3128 0 1 167
box -26 -22 76 88
use contact_11  contact_11_13
timestamp 1624494425
transform 1 0 3236 0 1 167
box -26 -22 76 88
use contact_11  contact_11_12
timestamp 1624494425
transform 1 0 3344 0 1 167
box -26 -22 76 88
use contact_11  contact_11_11
timestamp 1624494425
transform 1 0 3452 0 1 167
box -26 -22 76 88
use contact_11  contact_11_10
timestamp 1624494425
transform 1 0 3560 0 1 167
box -26 -22 76 88
use contact_11  contact_11_9
timestamp 1624494425
transform 1 0 3668 0 1 167
box -26 -22 76 88
use contact_11  contact_11_8
timestamp 1624494425
transform 1 0 3776 0 1 167
box -26 -22 76 88
use contact_11  contact_11_7
timestamp 1624494425
transform 1 0 3884 0 1 167
box -26 -22 76 88
use contact_11  contact_11_6
timestamp 1624494425
transform 1 0 3992 0 1 167
box -26 -22 76 88
use contact_11  contact_11_5
timestamp 1624494425
transform 1 0 4100 0 1 167
box -26 -22 76 88
use contact_11  contact_11_4
timestamp 1624494425
transform 1 0 4208 0 1 167
box -26 -22 76 88
use contact_11  contact_11_3
timestamp 1624494425
transform 1 0 4316 0 1 167
box -26 -22 76 88
use contact_11  contact_11_2
timestamp 1624494425
transform 1 0 4424 0 1 167
box -26 -22 76 88
use contact_11  contact_11_1
timestamp 1624494425
transform 1 0 4532 0 1 167
box -26 -22 76 88
use contact_11  contact_11_0
timestamp 1624494425
transform 1 0 4636 0 1 167
box -26 -22 76 88
<< labels >>
rlabel poly s 2343 441 2343 441 4 G
rlabel locali s 669 200 669 200 4 S
rlabel locali s 1965 200 1965 200 4 S
rlabel locali s 2829 200 2829 200 4 S
rlabel locali s 3261 200 3261 200 4 S
rlabel locali s 2397 200 2397 200 4 S
rlabel locali s 4557 200 4557 200 4 S
rlabel locali s 3045 200 3045 200 4 S
rlabel locali s 1749 200 1749 200 4 S
rlabel locali s 1533 200 1533 200 4 S
rlabel locali s 453 200 453 200 4 S
rlabel locali s 1101 200 1101 200 4 S
rlabel locali s 3909 200 3909 200 4 S
rlabel locali s 237 200 237 200 4 S
rlabel locali s 4125 200 4125 200 4 S
rlabel locali s 4341 200 4341 200 4 S
rlabel locali s 885 200 885 200 4 S
rlabel locali s 3693 200 3693 200 4 S
rlabel locali s 3477 200 3477 200 4 S
rlabel locali s 2613 200 2613 200 4 S
rlabel locali s 25 200 25 200 4 S
rlabel locali s 2181 200 2181 200 4 S
rlabel locali s 1317 200 1317 200 4 S
rlabel locali s 2395 284 2395 284 4 D
<< properties >>
string FIXED_BBOX -25 -26 4711 456
<< end >>
