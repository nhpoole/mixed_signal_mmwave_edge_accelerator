magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< error_s >>
rect 1168 2149 1204 2152
rect 1422 679 1458 2149
<< locali >>
rect 3642 9881 12502 9915
rect 3642 8467 12502 8501
rect 3806 7350 3840 7832
rect 3621 7316 3840 7350
rect 6388 7053 12502 7087
rect 5956 5639 12502 5673
rect 4668 4225 12502 4259
rect 4668 2811 12502 2845
rect 3603 2541 3788 2575
rect 3603 2176 3637 2541
rect 3470 2142 3637 2176
rect 5036 1397 12502 1431
rect 12070 -17 12502 17
<< metal1 >>
rect 12470 11286 12534 11338
rect 2700 10629 3355 10657
rect 9818 10579 9882 10631
rect 12470 9872 12534 9924
rect 2616 9139 3355 9167
rect 3438 9127 3502 9179
rect 12470 8458 12534 8510
rect 2784 8200 3403 8228
rect 2616 7952 3503 7980
rect 8018 7751 8082 7803
rect 12470 7044 12534 7096
rect 5000 6337 5064 6389
rect 2700 6160 3636 6188
rect 2532 6036 3503 6064
rect 2868 5912 3370 5940
rect 12470 5630 12534 5682
rect 2616 5372 3370 5400
rect 2700 5248 3503 5276
rect 2952 5124 3636 5152
rect 4784 4923 4848 4975
rect 1553 4308 2616 4336
rect 12470 4216 12534 4268
rect 383 4148 3036 4176
rect 4142 3493 4206 3545
rect 3120 3332 3503 3360
rect 3036 3084 3403 3112
rect 12470 2802 12534 2854
rect 3839 2284 3903 2336
rect 3036 2145 3355 2173
rect 4510 2111 4574 2163
rect 12470 1388 12534 1440
rect 3323 643 3387 695
rect 9600 681 9664 733
rect 12470 -26 12534 26
<< metal2 >>
rect -57 17699 -29 17727
rect 1539 4322 1567 6401
rect 369 2828 397 4162
rect 137 2238 203 2290
rect 137 538 203 590
rect 2518 0 2546 11352
rect 2602 0 2630 11352
rect 2686 0 2714 11352
rect 2770 0 2798 11352
rect 2854 0 2882 11352
rect 2938 0 2966 11352
rect 3022 0 3050 11352
rect 3106 0 3134 11352
rect 12474 11288 12530 11336
rect 9850 10591 12586 10619
rect 12474 9874 12530 9922
rect 3456 8587 3484 9153
rect 12474 8460 12530 8508
rect 8050 7763 12586 7791
rect 12474 7046 12530 7094
rect 5032 6349 12586 6377
rect 12474 5632 12530 5680
rect 4816 4935 12586 4963
rect 12474 4218 12530 4266
rect 4146 3495 4202 3543
rect 12474 2804 12530 2852
rect 3843 2286 3899 2334
rect 4528 1571 4556 2137
rect 12474 1390 12530 1438
rect 9632 707 12586 721
rect 9618 693 12586 707
rect 3341 655 3369 683
rect 9618 141 9646 693
rect 12474 -24 12530 24
<< metal3 >>
rect 607 18333 705 18431
rect 1343 18333 1441 18431
rect 607 16919 705 17017
rect 1343 16919 1441 17017
rect 607 15505 705 15603
rect 1343 15505 1441 15603
rect 607 14091 705 14189
rect 1343 14091 1441 14189
rect 607 12677 705 12775
rect 1343 12677 1441 12775
rect 607 11263 705 11361
rect 1343 11263 1441 11361
rect 12453 11263 12551 11361
rect 607 9849 705 9947
rect 1343 9849 1441 9947
rect 12453 9849 12551 9947
rect 2532 8557 3470 8617
rect 607 8435 705 8533
rect 1343 8435 1441 8533
rect 12453 8435 12551 8533
rect 607 7021 705 7119
rect 1343 7021 1441 7119
rect 12453 7021 12551 7119
rect 607 5607 705 5705
rect 1343 5607 1441 5705
rect 12453 5607 12551 5705
rect 12453 4193 12551 4291
rect 2784 3489 4174 3549
rect -49 2779 49 2877
rect 12453 2779 12551 2877
rect 2342 2295 2952 2355
rect 3120 2280 3871 2340
rect 1836 1913 2868 1973
rect 2700 1541 4542 1601
rect -49 1365 49 1463
rect 12453 1365 12551 1463
rect 1836 855 3120 915
rect 3036 111 9632 171
rect -49 -49 49 49
rect 12453 -49 12551 49
use dff_buf_array  dff_buf_array_0
timestamp 1624494425
transform 1 0 0 0 1 0
box -49 -49 2554 2877
use contact_9  contact_9_21
timestamp 1624494425
transform 1 0 1803 0 1 848
box 0 0 66 74
use contact_9  contact_9_20
timestamp 1624494425
transform 1 0 1803 0 1 1906
box 0 0 66 74
use contact_9  contact_9_19
timestamp 1624494425
transform 1 0 2309 0 1 2288
box 0 0 66 74
use contact_31  contact_31_9
timestamp 1624494425
transform 1 0 2835 0 1 1906
box 0 0 66 74
use contact_31  contact_31_8
timestamp 1624494425
transform 1 0 2919 0 1 2288
box 0 0 66 74
use contact_31  contact_31_1
timestamp 1624494425
transform 1 0 2667 0 1 1534
box 0 0 66 74
use pinv_1  pinv_1_1
timestamp 1624494425
transform 1 0 3274 0 -1 2828
box -36 -17 404 1471
use contact_7  contact_7_26
timestamp 1624494425
transform 1 0 3326 0 1 636
box 0 0 58 66
use contact_7  contact_7_23
timestamp 1624494425
transform 1 0 3326 0 1 2126
box 0 0 58 66
use contact_8  contact_8_26
timestamp 1624494425
transform 1 0 3323 0 1 637
box 0 0 64 64
use contact_8  contact_8_23
timestamp 1624494425
transform 1 0 3004 0 1 2127
box 0 0 64 64
use contact_31  contact_31_10
timestamp 1624494425
transform 1 0 3087 0 1 848
box 0 0 66 74
use contact_31  contact_31_4
timestamp 1624494425
transform 1 0 3003 0 1 104
box 0 0 66 74
use contact_31  contact_31_3
timestamp 1624494425
transform 1 0 3087 0 1 2273
box 0 0 66 74
use contact_31  contact_31_2
timestamp 1624494425
transform 1 0 4509 0 1 1534
box 0 0 66 74
use contact_9  contact_9_17
timestamp 1624494425
transform 1 0 3838 0 1 2273
box 0 0 66 74
use contact_9  contact_9_18
timestamp 1624494425
transform 1 0 3838 0 1 2273
box 0 0 66 74
use contact_8  contact_8_20
timestamp 1624494425
transform 1 0 4510 0 1 2105
box 0 0 64 64
use contact_8  contact_8_21
timestamp 1624494425
transform 1 0 3839 0 1 2278
box 0 0 64 64
use contact_8  contact_8_22
timestamp 1624494425
transform 1 0 3839 0 1 2278
box 0 0 64 64
use contact_7  contact_7_20
timestamp 1624494425
transform 1 0 4513 0 1 2104
box 0 0 58 66
use contact_7  contact_7_21
timestamp 1624494425
transform 1 0 3842 0 1 2277
box 0 0 58 66
use contact_7  contact_7_22
timestamp 1624494425
transform 1 0 3842 0 1 2277
box 0 0 58 66
use pand2_1  pand2_1_0
timestamp 1624494425
transform 1 0 3274 0 1 2828
box -36 -17 1430 1471
use pand2_1  pand2_1_1
timestamp 1624494425
transform 1 0 3642 0 -1 2828
box -36 -17 1430 1471
use contact_7  contact_7_25
timestamp 1624494425
transform 1 0 9603 0 1 674
box 0 0 58 66
use contact_7  contact_7_24
timestamp 1624494425
transform 1 0 9603 0 1 674
box 0 0 58 66
use contact_8  contact_8_25
timestamp 1624494425
transform 1 0 9600 0 1 675
box 0 0 64 64
use contact_8  contact_8_24
timestamp 1624494425
transform 1 0 9600 0 1 675
box 0 0 64 64
use contact_31  contact_31_5
timestamp 1624494425
transform 1 0 9599 0 1 104
box 0 0 66 74
use contact_7  contact_7_14
timestamp 1624494425
transform 1 0 12473 0 1 -33
box 0 0 58 66
use contact_8  contact_8_14
timestamp 1624494425
transform 1 0 12470 0 1 -32
box 0 0 64 64
use contact_9  contact_9_14
timestamp 1624494425
transform 1 0 12469 0 1 -37
box 0 0 66 74
use contact_7  contact_7_15
timestamp 1624494425
transform 1 0 12473 0 1 1381
box 0 0 58 66
use contact_7  contact_7_13
timestamp 1624494425
transform 1 0 12473 0 1 1381
box 0 0 58 66
use contact_8  contact_8_15
timestamp 1624494425
transform 1 0 12470 0 1 1382
box 0 0 64 64
use contact_8  contact_8_13
timestamp 1624494425
transform 1 0 12470 0 1 1382
box 0 0 64 64
use contact_9  contact_9_15
timestamp 1624494425
transform 1 0 12469 0 1 1377
box 0 0 66 74
use contact_9  contact_9_13
timestamp 1624494425
transform 1 0 12469 0 1 1377
box 0 0 66 74
use contact_7  contact_7_12
timestamp 1624494425
transform 1 0 12473 0 1 2795
box 0 0 58 66
use contact_7  contact_7_10
timestamp 1624494425
transform 1 0 12473 0 1 2795
box 0 0 58 66
use contact_8  contact_8_12
timestamp 1624494425
transform 1 0 12470 0 1 2796
box 0 0 64 64
use contact_8  contact_8_10
timestamp 1624494425
transform 1 0 12470 0 1 2796
box 0 0 64 64
use contact_9  contact_9_12
timestamp 1624494425
transform 1 0 12469 0 1 2791
box 0 0 66 74
use contact_9  contact_9_10
timestamp 1624494425
transform 1 0 12469 0 1 2791
box 0 0 66 74
use pdriver_2  pdriver_2_0
timestamp 1624494425
transform 1 0 3274 0 1 0
box -36 -17 8832 1471
use contact_31  contact_31_0
timestamp 1624494425
transform 1 0 2751 0 1 3482
box 0 0 66 74
use contact_8  contact_8_19
timestamp 1624494425
transform 1 0 3004 0 1 3066
box 0 0 64 64
use contact_8  contact_8_18
timestamp 1624494425
transform 1 0 3088 0 1 3314
box 0 0 64 64
use contact_8  contact_8_45
timestamp 1624494425
transform 1 0 351 0 1 4130
box 0 0 64 64
use contact_8  contact_8_31
timestamp 1624494425
transform 1 0 1521 0 1 4290
box 0 0 64 64
use contact_8  contact_8_30
timestamp 1624494425
transform 1 0 2584 0 1 4290
box 0 0 64 64
use contact_8  contact_8_44
timestamp 1624494425
transform 1 0 3004 0 1 4130
box 0 0 64 64
use contact_8  contact_8_35
timestamp 1624494425
transform 1 0 2584 0 1 5354
box 0 0 64 64
use contact_8  contact_8_34
timestamp 1624494425
transform 1 0 2668 0 1 5230
box 0 0 64 64
use contact_8  contact_8_33
timestamp 1624494425
transform 1 0 2920 0 1 5106
box 0 0 64 64
use contact_7  contact_7_19
timestamp 1624494425
transform 1 0 3374 0 1 3065
box 0 0 58 66
use contact_7  contact_7_18
timestamp 1624494425
transform 1 0 3474 0 1 3313
box 0 0 58 66
use contact_7  contact_7_17
timestamp 1624494425
transform 1 0 4145 0 1 3486
box 0 0 58 66
use contact_7  contact_7_16
timestamp 1624494425
transform 1 0 4145 0 1 3486
box 0 0 58 66
use contact_8  contact_8_17
timestamp 1624494425
transform 1 0 4142 0 1 3487
box 0 0 64 64
use contact_8  contact_8_16
timestamp 1624494425
transform 1 0 4142 0 1 3487
box 0 0 64 64
use contact_9  contact_9_16
timestamp 1624494425
transform 1 0 4141 0 1 3482
box 0 0 66 74
use contact_7  contact_7_33
timestamp 1624494425
transform 1 0 3341 0 1 5353
box 0 0 58 66
use contact_7  contact_7_32
timestamp 1624494425
transform 1 0 3474 0 1 5229
box 0 0 58 66
use contact_7  contact_7_31
timestamp 1624494425
transform 1 0 3607 0 1 5105
box 0 0 58 66
use contact_7  contact_7_30
timestamp 1624494425
transform 1 0 4787 0 1 4916
box 0 0 58 66
use contact_8  contact_8_32
timestamp 1624494425
transform 1 0 4784 0 1 4917
box 0 0 64 64
use pand3_0  pand3_0_0
timestamp 1624494425
transform 1 0 3274 0 -1 5656
box -36 -17 2718 1471
use pand3  pand3_0
timestamp 1624494425
transform 1 0 3274 0 1 5656
box -36 -17 3150 1471
use contact_7  contact_7_11
timestamp 1624494425
transform 1 0 12473 0 1 4209
box 0 0 58 66
use contact_7  contact_7_9
timestamp 1624494425
transform 1 0 12473 0 1 4209
box 0 0 58 66
use contact_8  contact_8_11
timestamp 1624494425
transform 1 0 12470 0 1 4210
box 0 0 64 64
use contact_8  contact_8_9
timestamp 1624494425
transform 1 0 12470 0 1 4210
box 0 0 64 64
use contact_9  contact_9_11
timestamp 1624494425
transform 1 0 12469 0 1 4205
box 0 0 66 74
use contact_9  contact_9_9
timestamp 1624494425
transform 1 0 12469 0 1 4205
box 0 0 66 74
use contact_7  contact_7_8
timestamp 1624494425
transform 1 0 12473 0 1 5623
box 0 0 58 66
use contact_7  contact_7_6
timestamp 1624494425
transform 1 0 12473 0 1 5623
box 0 0 58 66
use contact_8  contact_8_8
timestamp 1624494425
transform 1 0 12470 0 1 5624
box 0 0 64 64
use contact_8  contact_8_6
timestamp 1624494425
transform 1 0 12470 0 1 5624
box 0 0 64 64
use contact_9  contact_9_8
timestamp 1624494425
transform 1 0 12469 0 1 5619
box 0 0 66 74
use contact_9  contact_9_6
timestamp 1624494425
transform 1 0 12469 0 1 5619
box 0 0 66 74
use contact_8  contact_8_39
timestamp 1624494425
transform 1 0 2836 0 1 5894
box 0 0 64 64
use contact_8  contact_8_38
timestamp 1624494425
transform 1 0 2500 0 1 6018
box 0 0 64 64
use contact_8  contact_8_37
timestamp 1624494425
transform 1 0 2668 0 1 6142
box 0 0 64 64
use contact_8  contact_8_29
timestamp 1624494425
transform 1 0 2752 0 1 8182
box 0 0 64 64
use contact_8  contact_8_28
timestamp 1624494425
transform 1 0 2584 0 1 7934
box 0 0 64 64
use contact_31  contact_31_6
timestamp 1624494425
transform 1 0 2499 0 1 8550
box 0 0 66 74
use contact_7  contact_7_29
timestamp 1624494425
transform 1 0 3374 0 1 8181
box 0 0 58 66
use contact_7  contact_7_37
timestamp 1624494425
transform 1 0 3341 0 1 5893
box 0 0 58 66
use pinv_1  pinv_1_0
timestamp 1624494425
transform 1 0 3274 0 1 8484
box -36 -17 404 1471
use pnand2_1  pnand2_1_0
timestamp 1624494425
transform 1 0 3274 0 -1 8484
box -36 -17 504 1471
use contact_31  contact_31_7
timestamp 1624494425
transform 1 0 3437 0 1 8550
box 0 0 66 74
use contact_7  contact_7_28
timestamp 1624494425
transform 1 0 3474 0 1 7933
box 0 0 58 66
use contact_7  contact_7_35
timestamp 1624494425
transform 1 0 3607 0 1 6141
box 0 0 58 66
use contact_7  contact_7_36
timestamp 1624494425
transform 1 0 3474 0 1 6017
box 0 0 58 66
use contact_8  contact_8_36
timestamp 1624494425
transform 1 0 5000 0 1 6331
box 0 0 64 64
use contact_7  contact_7_34
timestamp 1624494425
transform 1 0 5003 0 1 6330
box 0 0 58 66
use pdriver_6  pdriver_6_0
timestamp 1624494425
transform 1 0 3742 0 -1 8484
box -36 -17 5808 1471
use contact_8  contact_8_27
timestamp 1624494425
transform 1 0 8018 0 1 7745
box 0 0 64 64
use contact_7  contact_7_27
timestamp 1624494425
transform 1 0 8021 0 1 7744
box 0 0 58 66
use contact_7  contact_7_7
timestamp 1624494425
transform 1 0 12473 0 1 7037
box 0 0 58 66
use contact_7  contact_7_5
timestamp 1624494425
transform 1 0 12473 0 1 7037
box 0 0 58 66
use contact_8  contact_8_7
timestamp 1624494425
transform 1 0 12470 0 1 7038
box 0 0 64 64
use contact_8  contact_8_5
timestamp 1624494425
transform 1 0 12470 0 1 7038
box 0 0 64 64
use contact_9  contact_9_7
timestamp 1624494425
transform 1 0 12469 0 1 7033
box 0 0 66 74
use contact_9  contact_9_5
timestamp 1624494425
transform 1 0 12469 0 1 7033
box 0 0 66 74
use contact_7  contact_7_4
timestamp 1624494425
transform 1 0 12473 0 1 8451
box 0 0 58 66
use contact_7  contact_7_2
timestamp 1624494425
transform 1 0 12473 0 1 8451
box 0 0 58 66
use contact_8  contact_8_4
timestamp 1624494425
transform 1 0 12470 0 1 8452
box 0 0 64 64
use contact_8  contact_8_2
timestamp 1624494425
transform 1 0 12470 0 1 8452
box 0 0 64 64
use contact_9  contact_9_4
timestamp 1624494425
transform 1 0 12469 0 1 8447
box 0 0 66 74
use contact_9  contact_9_2
timestamp 1624494425
transform 1 0 12469 0 1 8447
box 0 0 66 74
use contact_7  contact_7_39
timestamp 1624494425
transform 1 0 3441 0 1 9120
box 0 0 58 66
use contact_7  contact_7_38
timestamp 1624494425
transform 1 0 3326 0 1 9120
box 0 0 58 66
use contact_8  contact_8_41
timestamp 1624494425
transform 1 0 3438 0 1 9121
box 0 0 64 64
use contact_8  contact_8_40
timestamp 1624494425
transform 1 0 2584 0 1 9121
box 0 0 64 64
use contact_9  contact_9_1
timestamp 1624494425
transform 1 0 12469 0 1 9861
box 0 0 66 74
use contact_9  contact_9_3
timestamp 1624494425
transform 1 0 12469 0 1 9861
box 0 0 66 74
use contact_8  contact_8_1
timestamp 1624494425
transform 1 0 12470 0 1 9866
box 0 0 64 64
use contact_8  contact_8_3
timestamp 1624494425
transform 1 0 12470 0 1 9866
box 0 0 64 64
use contact_7  contact_7_1
timestamp 1624494425
transform 1 0 12473 0 1 9865
box 0 0 58 66
use contact_7  contact_7_3
timestamp 1624494425
transform 1 0 12473 0 1 9865
box 0 0 58 66
use contact_8  contact_8_42
timestamp 1624494425
transform 1 0 9818 0 1 10573
box 0 0 64 64
use contact_8  contact_8_43
timestamp 1624494425
transform 1 0 2668 0 1 10611
box 0 0 64 64
use contact_7  contact_7_40
timestamp 1624494425
transform 1 0 9821 0 1 10572
box 0 0 58 66
use contact_7  contact_7_41
timestamp 1624494425
transform 1 0 3326 0 1 10610
box 0 0 58 66
use pdriver_3  pdriver_3_0
timestamp 1624494425
transform 1 0 3274 0 -1 11312
box -36 -17 9264 1471
use contact_7  contact_7_0
timestamp 1624494425
transform 1 0 12473 0 1 11279
box 0 0 58 66
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 12470 0 1 11280
box 0 0 64 64
use contact_9  contact_9_0
timestamp 1624494425
transform 1 0 12469 0 1 11275
box 0 0 66 74
use delay_chain  delay_chain_0
timestamp 1624494425
transform 1 0 0 0 -1 18382
box -75 -49 1876 12783
<< labels >>
rlabel metal2 s 137 538 203 590 4 csb
rlabel metal2 s 137 2238 203 2290 4 web
rlabel metal2 s 9850 10591 12586 10619 4 wl_en
rlabel metal2 s 5032 6349 12586 6377 4 w_en
rlabel metal2 s 4816 4935 12586 4963 4 s_en
rlabel metal2 s -57 17699 -29 17727 4 rbl_bl
rlabel metal2 s 8050 7763 12586 7791 4 p_en_bar
rlabel metal2 s 3341 655 3369 683 4 clk
rlabel metal2 s 9632 693 12586 721 4 clk_buf
rlabel metal3 s 1343 5607 1441 5705 4 vdd
rlabel metal3 s 12453 9849 12551 9947 4 vdd
rlabel metal3 s 12453 7021 12551 7119 4 vdd
rlabel metal3 s 607 8435 705 8533 4 vdd
rlabel metal3 s 607 16919 705 17017 4 vdd
rlabel metal3 s 1343 16919 1441 17017 4 vdd
rlabel metal3 s 607 11263 705 11361 4 vdd
rlabel metal3 s 607 14091 705 14189 4 vdd
rlabel metal3 s 1343 14091 1441 14189 4 vdd
rlabel metal3 s 1343 11263 1441 11361 4 vdd
rlabel metal3 s -49 1365 49 1463 4 vdd
rlabel metal3 s 12453 4193 12551 4291 4 vdd
rlabel metal3 s 1343 8435 1441 8533 4 vdd
rlabel metal3 s 12453 1365 12551 1463 4 vdd
rlabel metal3 s 607 5607 705 5705 4 vdd
rlabel metal3 s 1343 7021 1441 7119 4 gnd
rlabel metal3 s 12453 2779 12551 2877 4 gnd
rlabel metal3 s 1343 15505 1441 15603 4 gnd
rlabel metal3 s 607 9849 705 9947 4 gnd
rlabel metal3 s 1343 9849 1441 9947 4 gnd
rlabel metal3 s 12453 8435 12551 8533 4 gnd
rlabel metal3 s 12453 5607 12551 5705 4 gnd
rlabel metal3 s 12453 -49 12551 49 4 gnd
rlabel metal3 s 12453 11263 12551 11361 4 gnd
rlabel metal3 s 1343 18333 1441 18431 4 gnd
rlabel metal3 s 607 15505 705 15603 4 gnd
rlabel metal3 s 607 7021 705 7119 4 gnd
rlabel metal3 s -49 2779 49 2877 4 gnd
rlabel metal3 s 607 18333 705 18431 4 gnd
rlabel metal3 s 607 12677 705 12775 4 gnd
rlabel metal3 s 1343 12677 1441 12775 4 gnd
rlabel metal3 s -49 -49 49 49 4 gnd
<< properties >>
string FIXED_BBOX 0 0 12586 18542
<< end >>
