magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -2405 -1448 2405 1448
<< pwell >>
rect -1145 -126 1145 126
<< nmoslvt >>
rect -1061 -100 -901 100
rect -843 -100 -683 100
rect -625 -100 -465 100
rect -407 -100 -247 100
rect -189 -100 -29 100
rect 29 -100 189 100
rect 247 -100 407 100
rect 465 -100 625 100
rect 683 -100 843 100
rect 901 -100 1061 100
<< ndiff >>
rect -1119 85 -1061 100
rect -1119 51 -1107 85
rect -1073 51 -1061 85
rect -1119 17 -1061 51
rect -1119 -17 -1107 17
rect -1073 -17 -1061 17
rect -1119 -51 -1061 -17
rect -1119 -85 -1107 -51
rect -1073 -85 -1061 -51
rect -1119 -100 -1061 -85
rect -901 85 -843 100
rect -901 51 -889 85
rect -855 51 -843 85
rect -901 17 -843 51
rect -901 -17 -889 17
rect -855 -17 -843 17
rect -901 -51 -843 -17
rect -901 -85 -889 -51
rect -855 -85 -843 -51
rect -901 -100 -843 -85
rect -683 85 -625 100
rect -683 51 -671 85
rect -637 51 -625 85
rect -683 17 -625 51
rect -683 -17 -671 17
rect -637 -17 -625 17
rect -683 -51 -625 -17
rect -683 -85 -671 -51
rect -637 -85 -625 -51
rect -683 -100 -625 -85
rect -465 85 -407 100
rect -465 51 -453 85
rect -419 51 -407 85
rect -465 17 -407 51
rect -465 -17 -453 17
rect -419 -17 -407 17
rect -465 -51 -407 -17
rect -465 -85 -453 -51
rect -419 -85 -407 -51
rect -465 -100 -407 -85
rect -247 85 -189 100
rect -247 51 -235 85
rect -201 51 -189 85
rect -247 17 -189 51
rect -247 -17 -235 17
rect -201 -17 -189 17
rect -247 -51 -189 -17
rect -247 -85 -235 -51
rect -201 -85 -189 -51
rect -247 -100 -189 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 189 85 247 100
rect 189 51 201 85
rect 235 51 247 85
rect 189 17 247 51
rect 189 -17 201 17
rect 235 -17 247 17
rect 189 -51 247 -17
rect 189 -85 201 -51
rect 235 -85 247 -51
rect 189 -100 247 -85
rect 407 85 465 100
rect 407 51 419 85
rect 453 51 465 85
rect 407 17 465 51
rect 407 -17 419 17
rect 453 -17 465 17
rect 407 -51 465 -17
rect 407 -85 419 -51
rect 453 -85 465 -51
rect 407 -100 465 -85
rect 625 85 683 100
rect 625 51 637 85
rect 671 51 683 85
rect 625 17 683 51
rect 625 -17 637 17
rect 671 -17 683 17
rect 625 -51 683 -17
rect 625 -85 637 -51
rect 671 -85 683 -51
rect 625 -100 683 -85
rect 843 85 901 100
rect 843 51 855 85
rect 889 51 901 85
rect 843 17 901 51
rect 843 -17 855 17
rect 889 -17 901 17
rect 843 -51 901 -17
rect 843 -85 855 -51
rect 889 -85 901 -51
rect 843 -100 901 -85
rect 1061 85 1119 100
rect 1061 51 1073 85
rect 1107 51 1119 85
rect 1061 17 1119 51
rect 1061 -17 1073 17
rect 1107 -17 1119 17
rect 1061 -51 1119 -17
rect 1061 -85 1073 -51
rect 1107 -85 1119 -51
rect 1061 -100 1119 -85
<< ndiffc >>
rect -1107 51 -1073 85
rect -1107 -17 -1073 17
rect -1107 -85 -1073 -51
rect -889 51 -855 85
rect -889 -17 -855 17
rect -889 -85 -855 -51
rect -671 51 -637 85
rect -671 -17 -637 17
rect -671 -85 -637 -51
rect -453 51 -419 85
rect -453 -17 -419 17
rect -453 -85 -419 -51
rect -235 51 -201 85
rect -235 -17 -201 17
rect -235 -85 -201 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 201 51 235 85
rect 201 -17 235 17
rect 201 -85 235 -51
rect 419 51 453 85
rect 419 -17 453 17
rect 419 -85 453 -51
rect 637 51 671 85
rect 637 -17 671 17
rect 637 -85 671 -51
rect 855 51 889 85
rect 855 -17 889 17
rect 855 -85 889 -51
rect 1073 51 1107 85
rect 1073 -17 1107 17
rect 1073 -85 1107 -51
<< poly >>
rect -1035 172 -927 188
rect -1035 155 -998 172
rect -1061 138 -998 155
rect -964 155 -927 172
rect -817 172 -709 188
rect -817 155 -780 172
rect -964 138 -901 155
rect -1061 100 -901 138
rect -843 138 -780 155
rect -746 155 -709 172
rect -599 172 -491 188
rect -599 155 -562 172
rect -746 138 -683 155
rect -843 100 -683 138
rect -625 138 -562 155
rect -528 155 -491 172
rect -381 172 -273 188
rect -381 155 -344 172
rect -528 138 -465 155
rect -625 100 -465 138
rect -407 138 -344 155
rect -310 155 -273 172
rect -163 172 -55 188
rect -163 155 -126 172
rect -310 138 -247 155
rect -407 100 -247 138
rect -189 138 -126 155
rect -92 155 -55 172
rect 55 172 163 188
rect 55 155 92 172
rect -92 138 -29 155
rect -189 100 -29 138
rect 29 138 92 155
rect 126 155 163 172
rect 273 172 381 188
rect 273 155 310 172
rect 126 138 189 155
rect 29 100 189 138
rect 247 138 310 155
rect 344 155 381 172
rect 491 172 599 188
rect 491 155 528 172
rect 344 138 407 155
rect 247 100 407 138
rect 465 138 528 155
rect 562 155 599 172
rect 709 172 817 188
rect 709 155 746 172
rect 562 138 625 155
rect 465 100 625 138
rect 683 138 746 155
rect 780 155 817 172
rect 927 172 1035 188
rect 927 155 964 172
rect 780 138 843 155
rect 683 100 843 138
rect 901 138 964 155
rect 998 155 1035 172
rect 998 138 1061 155
rect 901 100 1061 138
rect -1061 -138 -901 -100
rect -1061 -155 -998 -138
rect -1035 -172 -998 -155
rect -964 -155 -901 -138
rect -843 -138 -683 -100
rect -843 -155 -780 -138
rect -964 -172 -927 -155
rect -1035 -188 -927 -172
rect -817 -172 -780 -155
rect -746 -155 -683 -138
rect -625 -138 -465 -100
rect -625 -155 -562 -138
rect -746 -172 -709 -155
rect -817 -188 -709 -172
rect -599 -172 -562 -155
rect -528 -155 -465 -138
rect -407 -138 -247 -100
rect -407 -155 -344 -138
rect -528 -172 -491 -155
rect -599 -188 -491 -172
rect -381 -172 -344 -155
rect -310 -155 -247 -138
rect -189 -138 -29 -100
rect -189 -155 -126 -138
rect -310 -172 -273 -155
rect -381 -188 -273 -172
rect -163 -172 -126 -155
rect -92 -155 -29 -138
rect 29 -138 189 -100
rect 29 -155 92 -138
rect -92 -172 -55 -155
rect -163 -188 -55 -172
rect 55 -172 92 -155
rect 126 -155 189 -138
rect 247 -138 407 -100
rect 247 -155 310 -138
rect 126 -172 163 -155
rect 55 -188 163 -172
rect 273 -172 310 -155
rect 344 -155 407 -138
rect 465 -138 625 -100
rect 465 -155 528 -138
rect 344 -172 381 -155
rect 273 -188 381 -172
rect 491 -172 528 -155
rect 562 -155 625 -138
rect 683 -138 843 -100
rect 683 -155 746 -138
rect 562 -172 599 -155
rect 491 -188 599 -172
rect 709 -172 746 -155
rect 780 -155 843 -138
rect 901 -138 1061 -100
rect 901 -155 964 -138
rect 780 -172 817 -155
rect 709 -188 817 -172
rect 927 -172 964 -155
rect 998 -155 1061 -138
rect 998 -172 1035 -155
rect 927 -188 1035 -172
<< polycont >>
rect -998 138 -964 172
rect -780 138 -746 172
rect -562 138 -528 172
rect -344 138 -310 172
rect -126 138 -92 172
rect 92 138 126 172
rect 310 138 344 172
rect 528 138 562 172
rect 746 138 780 172
rect 964 138 998 172
rect -998 -172 -964 -138
rect -780 -172 -746 -138
rect -562 -172 -528 -138
rect -344 -172 -310 -138
rect -126 -172 -92 -138
rect 92 -172 126 -138
rect 310 -172 344 -138
rect 528 -172 562 -138
rect 746 -172 780 -138
rect 964 -172 998 -138
<< locali >>
rect -1035 138 -998 172
rect -964 138 -927 172
rect -817 138 -780 172
rect -746 138 -709 172
rect -599 138 -562 172
rect -528 138 -491 172
rect -381 138 -344 172
rect -310 138 -273 172
rect -163 138 -126 172
rect -92 138 -55 172
rect 55 138 92 172
rect 126 138 163 172
rect 273 138 310 172
rect 344 138 381 172
rect 491 138 528 172
rect 562 138 599 172
rect 709 138 746 172
rect 780 138 817 172
rect 927 138 964 172
rect 998 138 1035 172
rect -1107 85 -1073 104
rect -1107 17 -1073 19
rect -1107 -19 -1073 -17
rect -1107 -104 -1073 -85
rect -889 85 -855 104
rect -889 17 -855 19
rect -889 -19 -855 -17
rect -889 -104 -855 -85
rect -671 85 -637 104
rect -671 17 -637 19
rect -671 -19 -637 -17
rect -671 -104 -637 -85
rect -453 85 -419 104
rect -453 17 -419 19
rect -453 -19 -419 -17
rect -453 -104 -419 -85
rect -235 85 -201 104
rect -235 17 -201 19
rect -235 -19 -201 -17
rect -235 -104 -201 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 201 85 235 104
rect 201 17 235 19
rect 201 -19 235 -17
rect 201 -104 235 -85
rect 419 85 453 104
rect 419 17 453 19
rect 419 -19 453 -17
rect 419 -104 453 -85
rect 637 85 671 104
rect 637 17 671 19
rect 637 -19 671 -17
rect 637 -104 671 -85
rect 855 85 889 104
rect 855 17 889 19
rect 855 -19 889 -17
rect 855 -104 889 -85
rect 1073 85 1107 104
rect 1073 17 1107 19
rect 1073 -19 1107 -17
rect 1073 -104 1107 -85
rect -1035 -172 -998 -138
rect -964 -172 -927 -138
rect -817 -172 -780 -138
rect -746 -172 -709 -138
rect -599 -172 -562 -138
rect -528 -172 -491 -138
rect -381 -172 -344 -138
rect -310 -172 -273 -138
rect -163 -172 -126 -138
rect -92 -172 -55 -138
rect 55 -172 92 -138
rect 126 -172 163 -138
rect 273 -172 310 -138
rect 344 -172 381 -138
rect 491 -172 528 -138
rect 562 -172 599 -138
rect 709 -172 746 -138
rect 780 -172 817 -138
rect 927 -172 964 -138
rect 998 -172 1035 -138
<< viali >>
rect -998 138 -964 172
rect -780 138 -746 172
rect -562 138 -528 172
rect -344 138 -310 172
rect -126 138 -92 172
rect 92 138 126 172
rect 310 138 344 172
rect 528 138 562 172
rect 746 138 780 172
rect 964 138 998 172
rect -1107 51 -1073 53
rect -1107 19 -1073 51
rect -1107 -51 -1073 -19
rect -1107 -53 -1073 -51
rect -889 51 -855 53
rect -889 19 -855 51
rect -889 -51 -855 -19
rect -889 -53 -855 -51
rect -671 51 -637 53
rect -671 19 -637 51
rect -671 -51 -637 -19
rect -671 -53 -637 -51
rect -453 51 -419 53
rect -453 19 -419 51
rect -453 -51 -419 -19
rect -453 -53 -419 -51
rect -235 51 -201 53
rect -235 19 -201 51
rect -235 -51 -201 -19
rect -235 -53 -201 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 201 51 235 53
rect 201 19 235 51
rect 201 -51 235 -19
rect 201 -53 235 -51
rect 419 51 453 53
rect 419 19 453 51
rect 419 -51 453 -19
rect 419 -53 453 -51
rect 637 51 671 53
rect 637 19 671 51
rect 637 -51 671 -19
rect 637 -53 671 -51
rect 855 51 889 53
rect 855 19 889 51
rect 855 -51 889 -19
rect 855 -53 889 -51
rect 1073 51 1107 53
rect 1073 19 1107 51
rect 1073 -51 1107 -19
rect 1073 -53 1107 -51
rect -998 -172 -964 -138
rect -780 -172 -746 -138
rect -562 -172 -528 -138
rect -344 -172 -310 -138
rect -126 -172 -92 -138
rect 92 -172 126 -138
rect 310 -172 344 -138
rect 528 -172 562 -138
rect 746 -172 780 -138
rect 964 -172 998 -138
<< metal1 >>
rect -1025 172 -937 178
rect -1025 138 -998 172
rect -964 138 -937 172
rect -1025 132 -937 138
rect -807 172 -719 178
rect -807 138 -780 172
rect -746 138 -719 172
rect -807 132 -719 138
rect -589 172 -501 178
rect -589 138 -562 172
rect -528 138 -501 172
rect -589 132 -501 138
rect -371 172 -283 178
rect -371 138 -344 172
rect -310 138 -283 172
rect -371 132 -283 138
rect -153 172 -65 178
rect -153 138 -126 172
rect -92 138 -65 172
rect -153 132 -65 138
rect 65 172 153 178
rect 65 138 92 172
rect 126 138 153 172
rect 65 132 153 138
rect 283 172 371 178
rect 283 138 310 172
rect 344 138 371 172
rect 283 132 371 138
rect 501 172 589 178
rect 501 138 528 172
rect 562 138 589 172
rect 501 132 589 138
rect 719 172 807 178
rect 719 138 746 172
rect 780 138 807 172
rect 719 132 807 138
rect 937 172 1025 178
rect 937 138 964 172
rect 998 138 1025 172
rect 937 132 1025 138
rect -1113 53 -1067 100
rect -1113 19 -1107 53
rect -1073 19 -1067 53
rect -1113 -19 -1067 19
rect -1113 -53 -1107 -19
rect -1073 -53 -1067 -19
rect -1113 -100 -1067 -53
rect -895 53 -849 100
rect -895 19 -889 53
rect -855 19 -849 53
rect -895 -19 -849 19
rect -895 -53 -889 -19
rect -855 -53 -849 -19
rect -895 -100 -849 -53
rect -677 53 -631 100
rect -677 19 -671 53
rect -637 19 -631 53
rect -677 -19 -631 19
rect -677 -53 -671 -19
rect -637 -53 -631 -19
rect -677 -100 -631 -53
rect -459 53 -413 100
rect -459 19 -453 53
rect -419 19 -413 53
rect -459 -19 -413 19
rect -459 -53 -453 -19
rect -419 -53 -413 -19
rect -459 -100 -413 -53
rect -241 53 -195 100
rect -241 19 -235 53
rect -201 19 -195 53
rect -241 -19 -195 19
rect -241 -53 -235 -19
rect -201 -53 -195 -19
rect -241 -100 -195 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 195 53 241 100
rect 195 19 201 53
rect 235 19 241 53
rect 195 -19 241 19
rect 195 -53 201 -19
rect 235 -53 241 -19
rect 195 -100 241 -53
rect 413 53 459 100
rect 413 19 419 53
rect 453 19 459 53
rect 413 -19 459 19
rect 413 -53 419 -19
rect 453 -53 459 -19
rect 413 -100 459 -53
rect 631 53 677 100
rect 631 19 637 53
rect 671 19 677 53
rect 631 -19 677 19
rect 631 -53 637 -19
rect 671 -53 677 -19
rect 631 -100 677 -53
rect 849 53 895 100
rect 849 19 855 53
rect 889 19 895 53
rect 849 -19 895 19
rect 849 -53 855 -19
rect 889 -53 895 -19
rect 849 -100 895 -53
rect 1067 53 1113 100
rect 1067 19 1073 53
rect 1107 19 1113 53
rect 1067 -19 1113 19
rect 1067 -53 1073 -19
rect 1107 -53 1113 -19
rect 1067 -100 1113 -53
rect -1025 -138 -937 -132
rect -1025 -172 -998 -138
rect -964 -172 -937 -138
rect -1025 -178 -937 -172
rect -807 -138 -719 -132
rect -807 -172 -780 -138
rect -746 -172 -719 -138
rect -807 -178 -719 -172
rect -589 -138 -501 -132
rect -589 -172 -562 -138
rect -528 -172 -501 -138
rect -589 -178 -501 -172
rect -371 -138 -283 -132
rect -371 -172 -344 -138
rect -310 -172 -283 -138
rect -371 -178 -283 -172
rect -153 -138 -65 -132
rect -153 -172 -126 -138
rect -92 -172 -65 -138
rect -153 -178 -65 -172
rect 65 -138 153 -132
rect 65 -172 92 -138
rect 126 -172 153 -138
rect 65 -178 153 -172
rect 283 -138 371 -132
rect 283 -172 310 -138
rect 344 -172 371 -138
rect 283 -178 371 -172
rect 501 -138 589 -132
rect 501 -172 528 -138
rect 562 -172 589 -138
rect 501 -178 589 -172
rect 719 -138 807 -132
rect 719 -172 746 -138
rect 780 -172 807 -138
rect 719 -178 807 -172
rect 937 -138 1025 -132
rect 937 -172 964 -138
rect 998 -172 1025 -138
rect 937 -178 1025 -172
<< end >>
