magic
tech sky130A
magscale 1 2
timestamp 1623983327
<< metal1 >>
rect -100 30 100 87
rect -100 -87 100 -30
<< rmetal1 >>
rect -100 -30 100 30
<< properties >>
string gencell sky130_fd_pr__res_generic_m1
string parameters w 1 l 0.30 m 1 nx 1 wmin 0.14 lmin 0.14 rho 0.125 val 37.5m dummy 0 dw 0.0 term 0.0 roverlap 0
string library sky130
<< end >>
