magic
tech sky130A
magscale 1 2
timestamp 1621481787
<< metal4 >>
rect -1151 -900 657 900
<< mimcap2 >>
rect -1051 760 549 800
rect -1051 -760 -1011 760
rect 509 -760 549 760
rect -1051 -800 549 -760
<< mimcap2contact >>
rect -1011 -760 509 760
<< metal5 >>
rect -1035 760 533 784
rect -1035 -760 -1011 760
rect 509 -760 533 760
rect -1035 -784 533 -760
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -1151 -900 649 900
string parameters w 8.00 l 8.00 val 134.08 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
