magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -3860 -5120 8260 4000
<< nwell >>
rect -2562 -664 6962 2702
<< pwell >>
rect -2548 -1644 6948 -1492
rect -2548 -3656 -2396 -1644
rect 6796 -3656 6948 -1644
rect -2548 -3808 6948 -3656
<< psubdiff >>
rect -2522 -1551 6922 -1518
rect -2522 -1585 -2339 -1551
rect -2305 -1585 -2271 -1551
rect -2237 -1585 -2203 -1551
rect -2169 -1585 -2135 -1551
rect -2101 -1585 -2067 -1551
rect -2033 -1585 -1999 -1551
rect -1965 -1585 -1931 -1551
rect -1897 -1585 -1863 -1551
rect -1829 -1585 -1795 -1551
rect -1761 -1585 -1727 -1551
rect -1693 -1585 -1659 -1551
rect -1625 -1585 -1591 -1551
rect -1557 -1585 -1523 -1551
rect -1489 -1585 -1455 -1551
rect -1421 -1585 -1387 -1551
rect -1353 -1585 -1319 -1551
rect -1285 -1585 -1251 -1551
rect -1217 -1585 -1183 -1551
rect -1149 -1585 -1115 -1551
rect -1081 -1585 -1047 -1551
rect -1013 -1585 -979 -1551
rect -945 -1585 -911 -1551
rect -877 -1585 -843 -1551
rect -809 -1585 -775 -1551
rect -741 -1585 -707 -1551
rect -673 -1585 -639 -1551
rect -605 -1585 -571 -1551
rect -537 -1585 -503 -1551
rect -469 -1585 -435 -1551
rect -401 -1585 -367 -1551
rect -333 -1585 -299 -1551
rect -265 -1585 -231 -1551
rect -197 -1585 -163 -1551
rect -129 -1585 -95 -1551
rect -61 -1585 -27 -1551
rect 7 -1585 41 -1551
rect 75 -1585 109 -1551
rect 143 -1585 177 -1551
rect 211 -1585 245 -1551
rect 279 -1585 313 -1551
rect 347 -1585 381 -1551
rect 415 -1585 449 -1551
rect 483 -1585 517 -1551
rect 551 -1585 585 -1551
rect 619 -1585 653 -1551
rect 687 -1585 721 -1551
rect 755 -1585 789 -1551
rect 823 -1585 857 -1551
rect 891 -1585 925 -1551
rect 959 -1585 993 -1551
rect 1027 -1585 1061 -1551
rect 1095 -1585 1129 -1551
rect 1163 -1585 1197 -1551
rect 1231 -1585 1265 -1551
rect 1299 -1585 1333 -1551
rect 1367 -1585 1401 -1551
rect 1435 -1585 1469 -1551
rect 1503 -1585 1537 -1551
rect 1571 -1585 1605 -1551
rect 1639 -1585 1673 -1551
rect 1707 -1585 1741 -1551
rect 1775 -1585 1809 -1551
rect 1843 -1585 1877 -1551
rect 1911 -1585 1945 -1551
rect 1979 -1585 2013 -1551
rect 2047 -1585 2081 -1551
rect 2115 -1585 2149 -1551
rect 2183 -1585 2217 -1551
rect 2251 -1585 2285 -1551
rect 2319 -1585 2353 -1551
rect 2387 -1585 2421 -1551
rect 2455 -1585 2489 -1551
rect 2523 -1585 2557 -1551
rect 2591 -1585 2625 -1551
rect 2659 -1585 2693 -1551
rect 2727 -1585 2761 -1551
rect 2795 -1585 2829 -1551
rect 2863 -1585 2897 -1551
rect 2931 -1585 2965 -1551
rect 2999 -1585 3033 -1551
rect 3067 -1585 3101 -1551
rect 3135 -1585 3169 -1551
rect 3203 -1585 3237 -1551
rect 3271 -1585 3305 -1551
rect 3339 -1585 3373 -1551
rect 3407 -1585 3441 -1551
rect 3475 -1585 3509 -1551
rect 3543 -1585 3577 -1551
rect 3611 -1585 3645 -1551
rect 3679 -1585 3713 -1551
rect 3747 -1585 3781 -1551
rect 3815 -1585 3849 -1551
rect 3883 -1585 3917 -1551
rect 3951 -1585 3985 -1551
rect 4019 -1585 4053 -1551
rect 4087 -1585 4121 -1551
rect 4155 -1585 4189 -1551
rect 4223 -1585 4257 -1551
rect 4291 -1585 4325 -1551
rect 4359 -1585 4393 -1551
rect 4427 -1585 4461 -1551
rect 4495 -1585 4529 -1551
rect 4563 -1585 4597 -1551
rect 4631 -1585 4665 -1551
rect 4699 -1585 4733 -1551
rect 4767 -1585 4801 -1551
rect 4835 -1585 4869 -1551
rect 4903 -1585 4937 -1551
rect 4971 -1585 5005 -1551
rect 5039 -1585 5073 -1551
rect 5107 -1585 5141 -1551
rect 5175 -1585 5209 -1551
rect 5243 -1585 5277 -1551
rect 5311 -1585 5345 -1551
rect 5379 -1585 5413 -1551
rect 5447 -1585 5481 -1551
rect 5515 -1585 5549 -1551
rect 5583 -1585 5617 -1551
rect 5651 -1585 5685 -1551
rect 5719 -1585 5753 -1551
rect 5787 -1585 5821 -1551
rect 5855 -1585 5889 -1551
rect 5923 -1585 5957 -1551
rect 5991 -1585 6025 -1551
rect 6059 -1585 6093 -1551
rect 6127 -1585 6161 -1551
rect 6195 -1585 6229 -1551
rect 6263 -1585 6297 -1551
rect 6331 -1585 6365 -1551
rect 6399 -1585 6433 -1551
rect 6467 -1585 6501 -1551
rect 6535 -1585 6569 -1551
rect 6603 -1585 6637 -1551
rect 6671 -1585 6705 -1551
rect 6739 -1585 6922 -1551
rect -2522 -1618 6922 -1585
rect -2522 -1681 -2422 -1618
rect -2522 -1715 -2489 -1681
rect -2455 -1715 -2422 -1681
rect -2522 -1749 -2422 -1715
rect -2522 -1783 -2489 -1749
rect -2455 -1783 -2422 -1749
rect -2522 -1817 -2422 -1783
rect -2522 -1851 -2489 -1817
rect -2455 -1851 -2422 -1817
rect -2522 -1885 -2422 -1851
rect -2522 -1919 -2489 -1885
rect -2455 -1919 -2422 -1885
rect -2522 -1953 -2422 -1919
rect -2522 -1987 -2489 -1953
rect -2455 -1987 -2422 -1953
rect -2522 -2021 -2422 -1987
rect -2522 -2055 -2489 -2021
rect -2455 -2055 -2422 -2021
rect -2522 -2089 -2422 -2055
rect -2522 -2123 -2489 -2089
rect -2455 -2123 -2422 -2089
rect -2522 -2157 -2422 -2123
rect -2522 -2191 -2489 -2157
rect -2455 -2191 -2422 -2157
rect -2522 -2225 -2422 -2191
rect -2522 -2259 -2489 -2225
rect -2455 -2259 -2422 -2225
rect -2522 -2293 -2422 -2259
rect -2522 -2327 -2489 -2293
rect -2455 -2327 -2422 -2293
rect -2522 -2361 -2422 -2327
rect -2522 -2395 -2489 -2361
rect -2455 -2395 -2422 -2361
rect -2522 -2429 -2422 -2395
rect -2522 -2463 -2489 -2429
rect -2455 -2463 -2422 -2429
rect -2522 -2497 -2422 -2463
rect -2522 -2531 -2489 -2497
rect -2455 -2531 -2422 -2497
rect -2522 -2565 -2422 -2531
rect -2522 -2599 -2489 -2565
rect -2455 -2599 -2422 -2565
rect -2522 -2633 -2422 -2599
rect -2522 -2667 -2489 -2633
rect -2455 -2667 -2422 -2633
rect -2522 -2701 -2422 -2667
rect -2522 -2735 -2489 -2701
rect -2455 -2735 -2422 -2701
rect -2522 -2769 -2422 -2735
rect -2522 -2803 -2489 -2769
rect -2455 -2803 -2422 -2769
rect -2522 -2837 -2422 -2803
rect -2522 -2871 -2489 -2837
rect -2455 -2871 -2422 -2837
rect -2522 -2905 -2422 -2871
rect -2522 -2939 -2489 -2905
rect -2455 -2939 -2422 -2905
rect -2522 -2973 -2422 -2939
rect -2522 -3007 -2489 -2973
rect -2455 -3007 -2422 -2973
rect -2522 -3041 -2422 -3007
rect -2522 -3075 -2489 -3041
rect -2455 -3075 -2422 -3041
rect -2522 -3109 -2422 -3075
rect -2522 -3143 -2489 -3109
rect -2455 -3143 -2422 -3109
rect -2522 -3177 -2422 -3143
rect -2522 -3211 -2489 -3177
rect -2455 -3211 -2422 -3177
rect -2522 -3245 -2422 -3211
rect -2522 -3279 -2489 -3245
rect -2455 -3279 -2422 -3245
rect -2522 -3313 -2422 -3279
rect -2522 -3347 -2489 -3313
rect -2455 -3347 -2422 -3313
rect -2522 -3381 -2422 -3347
rect -2522 -3415 -2489 -3381
rect -2455 -3415 -2422 -3381
rect -2522 -3449 -2422 -3415
rect -2522 -3483 -2489 -3449
rect -2455 -3483 -2422 -3449
rect -2522 -3517 -2422 -3483
rect -2522 -3551 -2489 -3517
rect -2455 -3551 -2422 -3517
rect -2522 -3585 -2422 -3551
rect -2522 -3619 -2489 -3585
rect -2455 -3619 -2422 -3585
rect -2522 -3682 -2422 -3619
rect 6822 -1681 6922 -1618
rect 6822 -1715 6855 -1681
rect 6889 -1715 6922 -1681
rect 6822 -1749 6922 -1715
rect 6822 -1783 6855 -1749
rect 6889 -1783 6922 -1749
rect 6822 -1817 6922 -1783
rect 6822 -1851 6855 -1817
rect 6889 -1851 6922 -1817
rect 6822 -1885 6922 -1851
rect 6822 -1919 6855 -1885
rect 6889 -1919 6922 -1885
rect 6822 -1953 6922 -1919
rect 6822 -1987 6855 -1953
rect 6889 -1987 6922 -1953
rect 6822 -2021 6922 -1987
rect 6822 -2055 6855 -2021
rect 6889 -2055 6922 -2021
rect 6822 -2089 6922 -2055
rect 6822 -2123 6855 -2089
rect 6889 -2123 6922 -2089
rect 6822 -2157 6922 -2123
rect 6822 -2191 6855 -2157
rect 6889 -2191 6922 -2157
rect 6822 -2225 6922 -2191
rect 6822 -2259 6855 -2225
rect 6889 -2259 6922 -2225
rect 6822 -2293 6922 -2259
rect 6822 -2327 6855 -2293
rect 6889 -2327 6922 -2293
rect 6822 -2361 6922 -2327
rect 6822 -2395 6855 -2361
rect 6889 -2395 6922 -2361
rect 6822 -2429 6922 -2395
rect 6822 -2463 6855 -2429
rect 6889 -2463 6922 -2429
rect 6822 -2497 6922 -2463
rect 6822 -2531 6855 -2497
rect 6889 -2531 6922 -2497
rect 6822 -2565 6922 -2531
rect 6822 -2599 6855 -2565
rect 6889 -2599 6922 -2565
rect 6822 -2633 6922 -2599
rect 6822 -2667 6855 -2633
rect 6889 -2667 6922 -2633
rect 6822 -2701 6922 -2667
rect 6822 -2735 6855 -2701
rect 6889 -2735 6922 -2701
rect 6822 -2769 6922 -2735
rect 6822 -2803 6855 -2769
rect 6889 -2803 6922 -2769
rect 6822 -2837 6922 -2803
rect 6822 -2871 6855 -2837
rect 6889 -2871 6922 -2837
rect 6822 -2905 6922 -2871
rect 6822 -2939 6855 -2905
rect 6889 -2939 6922 -2905
rect 6822 -2973 6922 -2939
rect 6822 -3007 6855 -2973
rect 6889 -3007 6922 -2973
rect 6822 -3041 6922 -3007
rect 6822 -3075 6855 -3041
rect 6889 -3075 6922 -3041
rect 6822 -3109 6922 -3075
rect 6822 -3143 6855 -3109
rect 6889 -3143 6922 -3109
rect 6822 -3177 6922 -3143
rect 6822 -3211 6855 -3177
rect 6889 -3211 6922 -3177
rect 6822 -3245 6922 -3211
rect 6822 -3279 6855 -3245
rect 6889 -3279 6922 -3245
rect 6822 -3313 6922 -3279
rect 6822 -3347 6855 -3313
rect 6889 -3347 6922 -3313
rect 6822 -3381 6922 -3347
rect 6822 -3415 6855 -3381
rect 6889 -3415 6922 -3381
rect 6822 -3449 6922 -3415
rect 6822 -3483 6855 -3449
rect 6889 -3483 6922 -3449
rect 6822 -3517 6922 -3483
rect 6822 -3551 6855 -3517
rect 6889 -3551 6922 -3517
rect 6822 -3585 6922 -3551
rect 6822 -3619 6855 -3585
rect 6889 -3619 6922 -3585
rect 6822 -3682 6922 -3619
rect -2522 -3715 6922 -3682
rect -2522 -3749 -2339 -3715
rect -2305 -3749 -2271 -3715
rect -2237 -3749 -2203 -3715
rect -2169 -3749 -2135 -3715
rect -2101 -3749 -2067 -3715
rect -2033 -3749 -1999 -3715
rect -1965 -3749 -1931 -3715
rect -1897 -3749 -1863 -3715
rect -1829 -3749 -1795 -3715
rect -1761 -3749 -1727 -3715
rect -1693 -3749 -1659 -3715
rect -1625 -3749 -1591 -3715
rect -1557 -3749 -1523 -3715
rect -1489 -3749 -1455 -3715
rect -1421 -3749 -1387 -3715
rect -1353 -3749 -1319 -3715
rect -1285 -3749 -1251 -3715
rect -1217 -3749 -1183 -3715
rect -1149 -3749 -1115 -3715
rect -1081 -3749 -1047 -3715
rect -1013 -3749 -979 -3715
rect -945 -3749 -911 -3715
rect -877 -3749 -843 -3715
rect -809 -3749 -775 -3715
rect -741 -3749 -707 -3715
rect -673 -3749 -639 -3715
rect -605 -3749 -571 -3715
rect -537 -3749 -503 -3715
rect -469 -3749 -435 -3715
rect -401 -3749 -367 -3715
rect -333 -3749 -299 -3715
rect -265 -3749 -231 -3715
rect -197 -3749 -163 -3715
rect -129 -3749 -95 -3715
rect -61 -3749 -27 -3715
rect 7 -3749 41 -3715
rect 75 -3749 109 -3715
rect 143 -3749 177 -3715
rect 211 -3749 245 -3715
rect 279 -3749 313 -3715
rect 347 -3749 381 -3715
rect 415 -3749 449 -3715
rect 483 -3749 517 -3715
rect 551 -3749 585 -3715
rect 619 -3749 653 -3715
rect 687 -3749 721 -3715
rect 755 -3749 789 -3715
rect 823 -3749 857 -3715
rect 891 -3749 925 -3715
rect 959 -3749 993 -3715
rect 1027 -3749 1061 -3715
rect 1095 -3749 1129 -3715
rect 1163 -3749 1197 -3715
rect 1231 -3749 1265 -3715
rect 1299 -3749 1333 -3715
rect 1367 -3749 1401 -3715
rect 1435 -3749 1469 -3715
rect 1503 -3749 1537 -3715
rect 1571 -3749 1605 -3715
rect 1639 -3749 1673 -3715
rect 1707 -3749 1741 -3715
rect 1775 -3749 1809 -3715
rect 1843 -3749 1877 -3715
rect 1911 -3749 1945 -3715
rect 1979 -3749 2013 -3715
rect 2047 -3749 2081 -3715
rect 2115 -3749 2149 -3715
rect 2183 -3749 2217 -3715
rect 2251 -3749 2285 -3715
rect 2319 -3749 2353 -3715
rect 2387 -3749 2421 -3715
rect 2455 -3749 2489 -3715
rect 2523 -3749 2557 -3715
rect 2591 -3749 2625 -3715
rect 2659 -3749 2693 -3715
rect 2727 -3749 2761 -3715
rect 2795 -3749 2829 -3715
rect 2863 -3749 2897 -3715
rect 2931 -3749 2965 -3715
rect 2999 -3749 3033 -3715
rect 3067 -3749 3101 -3715
rect 3135 -3749 3169 -3715
rect 3203 -3749 3237 -3715
rect 3271 -3749 3305 -3715
rect 3339 -3749 3373 -3715
rect 3407 -3749 3441 -3715
rect 3475 -3749 3509 -3715
rect 3543 -3749 3577 -3715
rect 3611 -3749 3645 -3715
rect 3679 -3749 3713 -3715
rect 3747 -3749 3781 -3715
rect 3815 -3749 3849 -3715
rect 3883 -3749 3917 -3715
rect 3951 -3749 3985 -3715
rect 4019 -3749 4053 -3715
rect 4087 -3749 4121 -3715
rect 4155 -3749 4189 -3715
rect 4223 -3749 4257 -3715
rect 4291 -3749 4325 -3715
rect 4359 -3749 4393 -3715
rect 4427 -3749 4461 -3715
rect 4495 -3749 4529 -3715
rect 4563 -3749 4597 -3715
rect 4631 -3749 4665 -3715
rect 4699 -3749 4733 -3715
rect 4767 -3749 4801 -3715
rect 4835 -3749 4869 -3715
rect 4903 -3749 4937 -3715
rect 4971 -3749 5005 -3715
rect 5039 -3749 5073 -3715
rect 5107 -3749 5141 -3715
rect 5175 -3749 5209 -3715
rect 5243 -3749 5277 -3715
rect 5311 -3749 5345 -3715
rect 5379 -3749 5413 -3715
rect 5447 -3749 5481 -3715
rect 5515 -3749 5549 -3715
rect 5583 -3749 5617 -3715
rect 5651 -3749 5685 -3715
rect 5719 -3749 5753 -3715
rect 5787 -3749 5821 -3715
rect 5855 -3749 5889 -3715
rect 5923 -3749 5957 -3715
rect 5991 -3749 6025 -3715
rect 6059 -3749 6093 -3715
rect 6127 -3749 6161 -3715
rect 6195 -3749 6229 -3715
rect 6263 -3749 6297 -3715
rect 6331 -3749 6365 -3715
rect 6399 -3749 6433 -3715
rect 6467 -3749 6501 -3715
rect 6535 -3749 6569 -3715
rect 6603 -3749 6637 -3715
rect 6671 -3749 6705 -3715
rect 6739 -3749 6922 -3715
rect -2522 -3782 6922 -3749
<< nsubdiff >>
rect -2522 2629 6922 2662
rect -2522 2595 -2339 2629
rect -2305 2595 -2271 2629
rect -2237 2595 -2203 2629
rect -2169 2595 -2135 2629
rect -2101 2595 -2067 2629
rect -2033 2595 -1999 2629
rect -1965 2595 -1931 2629
rect -1897 2595 -1863 2629
rect -1829 2595 -1795 2629
rect -1761 2595 -1727 2629
rect -1693 2595 -1659 2629
rect -1625 2595 -1591 2629
rect -1557 2595 -1523 2629
rect -1489 2595 -1455 2629
rect -1421 2595 -1387 2629
rect -1353 2595 -1319 2629
rect -1285 2595 -1251 2629
rect -1217 2595 -1183 2629
rect -1149 2595 -1115 2629
rect -1081 2595 -1047 2629
rect -1013 2595 -979 2629
rect -945 2595 -911 2629
rect -877 2595 -843 2629
rect -809 2595 -775 2629
rect -741 2595 -707 2629
rect -673 2595 -639 2629
rect -605 2595 -571 2629
rect -537 2595 -503 2629
rect -469 2595 -435 2629
rect -401 2595 -367 2629
rect -333 2595 -299 2629
rect -265 2595 -231 2629
rect -197 2595 -163 2629
rect -129 2595 -95 2629
rect -61 2595 -27 2629
rect 7 2595 41 2629
rect 75 2595 109 2629
rect 143 2595 177 2629
rect 211 2595 245 2629
rect 279 2595 313 2629
rect 347 2595 381 2629
rect 415 2595 449 2629
rect 483 2595 517 2629
rect 551 2595 585 2629
rect 619 2595 653 2629
rect 687 2595 721 2629
rect 755 2595 789 2629
rect 823 2595 857 2629
rect 891 2595 925 2629
rect 959 2595 993 2629
rect 1027 2595 1061 2629
rect 1095 2595 1129 2629
rect 1163 2595 1197 2629
rect 1231 2595 1265 2629
rect 1299 2595 1333 2629
rect 1367 2595 1401 2629
rect 1435 2595 1469 2629
rect 1503 2595 1537 2629
rect 1571 2595 1605 2629
rect 1639 2595 1673 2629
rect 1707 2595 1741 2629
rect 1775 2595 1809 2629
rect 1843 2595 1877 2629
rect 1911 2595 1945 2629
rect 1979 2595 2013 2629
rect 2047 2595 2081 2629
rect 2115 2595 2149 2629
rect 2183 2595 2217 2629
rect 2251 2595 2285 2629
rect 2319 2595 2353 2629
rect 2387 2595 2421 2629
rect 2455 2595 2489 2629
rect 2523 2595 2557 2629
rect 2591 2595 2625 2629
rect 2659 2595 2693 2629
rect 2727 2595 2761 2629
rect 2795 2595 2829 2629
rect 2863 2595 2897 2629
rect 2931 2595 2965 2629
rect 2999 2595 3033 2629
rect 3067 2595 3101 2629
rect 3135 2595 3169 2629
rect 3203 2595 3237 2629
rect 3271 2595 3305 2629
rect 3339 2595 3373 2629
rect 3407 2595 3441 2629
rect 3475 2595 3509 2629
rect 3543 2595 3577 2629
rect 3611 2595 3645 2629
rect 3679 2595 3713 2629
rect 3747 2595 3781 2629
rect 3815 2595 3849 2629
rect 3883 2595 3917 2629
rect 3951 2595 3985 2629
rect 4019 2595 4053 2629
rect 4087 2595 4121 2629
rect 4155 2595 4189 2629
rect 4223 2595 4257 2629
rect 4291 2595 4325 2629
rect 4359 2595 4393 2629
rect 4427 2595 4461 2629
rect 4495 2595 4529 2629
rect 4563 2595 4597 2629
rect 4631 2595 4665 2629
rect 4699 2595 4733 2629
rect 4767 2595 4801 2629
rect 4835 2595 4869 2629
rect 4903 2595 4937 2629
rect 4971 2595 5005 2629
rect 5039 2595 5073 2629
rect 5107 2595 5141 2629
rect 5175 2595 5209 2629
rect 5243 2595 5277 2629
rect 5311 2595 5345 2629
rect 5379 2595 5413 2629
rect 5447 2595 5481 2629
rect 5515 2595 5549 2629
rect 5583 2595 5617 2629
rect 5651 2595 5685 2629
rect 5719 2595 5753 2629
rect 5787 2595 5821 2629
rect 5855 2595 5889 2629
rect 5923 2595 5957 2629
rect 5991 2595 6025 2629
rect 6059 2595 6093 2629
rect 6127 2595 6161 2629
rect 6195 2595 6229 2629
rect 6263 2595 6297 2629
rect 6331 2595 6365 2629
rect 6399 2595 6433 2629
rect 6467 2595 6501 2629
rect 6535 2595 6569 2629
rect 6603 2595 6637 2629
rect 6671 2595 6705 2629
rect 6739 2595 6922 2629
rect -2522 2562 6922 2595
rect -2522 2479 -2422 2562
rect -2522 2445 -2489 2479
rect -2455 2445 -2422 2479
rect -2522 2411 -2422 2445
rect -2522 2377 -2489 2411
rect -2455 2377 -2422 2411
rect -2522 2343 -2422 2377
rect -2522 2309 -2489 2343
rect -2455 2309 -2422 2343
rect -2522 2275 -2422 2309
rect -2522 2241 -2489 2275
rect -2455 2241 -2422 2275
rect -2522 2207 -2422 2241
rect -2522 2173 -2489 2207
rect -2455 2173 -2422 2207
rect -2522 2139 -2422 2173
rect -2522 2105 -2489 2139
rect -2455 2105 -2422 2139
rect -2522 2071 -2422 2105
rect -2522 2037 -2489 2071
rect -2455 2037 -2422 2071
rect -2522 2003 -2422 2037
rect -2522 1969 -2489 2003
rect -2455 1969 -2422 2003
rect -2522 1935 -2422 1969
rect -2522 1901 -2489 1935
rect -2455 1901 -2422 1935
rect -2522 1867 -2422 1901
rect -2522 1833 -2489 1867
rect -2455 1833 -2422 1867
rect -2522 1799 -2422 1833
rect -2522 1765 -2489 1799
rect -2455 1765 -2422 1799
rect -2522 1731 -2422 1765
rect -2522 1697 -2489 1731
rect -2455 1697 -2422 1731
rect -2522 1663 -2422 1697
rect -2522 1629 -2489 1663
rect -2455 1629 -2422 1663
rect -2522 1595 -2422 1629
rect -2522 1561 -2489 1595
rect -2455 1561 -2422 1595
rect -2522 1527 -2422 1561
rect -2522 1493 -2489 1527
rect -2455 1493 -2422 1527
rect -2522 1459 -2422 1493
rect -2522 1425 -2489 1459
rect -2455 1425 -2422 1459
rect -2522 1391 -2422 1425
rect -2522 1357 -2489 1391
rect -2455 1357 -2422 1391
rect -2522 1323 -2422 1357
rect -2522 1289 -2489 1323
rect -2455 1289 -2422 1323
rect -2522 1255 -2422 1289
rect -2522 1221 -2489 1255
rect -2455 1221 -2422 1255
rect -2522 1187 -2422 1221
rect -2522 1153 -2489 1187
rect -2455 1153 -2422 1187
rect -2522 1119 -2422 1153
rect -2522 1085 -2489 1119
rect -2455 1085 -2422 1119
rect -2522 1051 -2422 1085
rect -2522 1017 -2489 1051
rect -2455 1017 -2422 1051
rect -2522 983 -2422 1017
rect -2522 949 -2489 983
rect -2455 949 -2422 983
rect -2522 915 -2422 949
rect -2522 881 -2489 915
rect -2455 881 -2422 915
rect -2522 847 -2422 881
rect -2522 813 -2489 847
rect -2455 813 -2422 847
rect -2522 779 -2422 813
rect -2522 745 -2489 779
rect -2455 745 -2422 779
rect -2522 711 -2422 745
rect -2522 677 -2489 711
rect -2455 677 -2422 711
rect -2522 643 -2422 677
rect -2522 609 -2489 643
rect -2455 609 -2422 643
rect -2522 575 -2422 609
rect -2522 541 -2489 575
rect -2455 541 -2422 575
rect -2522 458 -2422 541
rect 6822 2479 6922 2562
rect 6822 2445 6855 2479
rect 6889 2445 6922 2479
rect 6822 2411 6922 2445
rect 6822 2377 6855 2411
rect 6889 2377 6922 2411
rect 6822 2343 6922 2377
rect 6822 2309 6855 2343
rect 6889 2309 6922 2343
rect 6822 2275 6922 2309
rect 6822 2241 6855 2275
rect 6889 2241 6922 2275
rect 6822 2207 6922 2241
rect 6822 2173 6855 2207
rect 6889 2173 6922 2207
rect 6822 2139 6922 2173
rect 6822 2105 6855 2139
rect 6889 2105 6922 2139
rect 6822 2071 6922 2105
rect 6822 2037 6855 2071
rect 6889 2037 6922 2071
rect 6822 2003 6922 2037
rect 6822 1969 6855 2003
rect 6889 1969 6922 2003
rect 6822 1935 6922 1969
rect 6822 1901 6855 1935
rect 6889 1901 6922 1935
rect 6822 1867 6922 1901
rect 6822 1833 6855 1867
rect 6889 1833 6922 1867
rect 6822 1799 6922 1833
rect 6822 1765 6855 1799
rect 6889 1765 6922 1799
rect 6822 1731 6922 1765
rect 6822 1697 6855 1731
rect 6889 1697 6922 1731
rect 6822 1663 6922 1697
rect 6822 1629 6855 1663
rect 6889 1629 6922 1663
rect 6822 1595 6922 1629
rect 6822 1561 6855 1595
rect 6889 1561 6922 1595
rect 6822 1527 6922 1561
rect 6822 1493 6855 1527
rect 6889 1493 6922 1527
rect 6822 1459 6922 1493
rect 6822 1425 6855 1459
rect 6889 1425 6922 1459
rect 6822 1391 6922 1425
rect 6822 1357 6855 1391
rect 6889 1357 6922 1391
rect 6822 1323 6922 1357
rect 6822 1289 6855 1323
rect 6889 1289 6922 1323
rect 6822 1255 6922 1289
rect 6822 1221 6855 1255
rect 6889 1221 6922 1255
rect 6822 1187 6922 1221
rect 6822 1153 6855 1187
rect 6889 1153 6922 1187
rect 6822 1119 6922 1153
rect 6822 1085 6855 1119
rect 6889 1085 6922 1119
rect 6822 1051 6922 1085
rect 6822 1017 6855 1051
rect 6889 1017 6922 1051
rect 6822 983 6922 1017
rect 6822 949 6855 983
rect 6889 949 6922 983
rect 6822 915 6922 949
rect 6822 881 6855 915
rect 6889 881 6922 915
rect 6822 847 6922 881
rect 6822 813 6855 847
rect 6889 813 6922 847
rect 6822 779 6922 813
rect 6822 745 6855 779
rect 6889 745 6922 779
rect 6822 711 6922 745
rect 6822 677 6855 711
rect 6889 677 6922 711
rect 6822 643 6922 677
rect 6822 609 6855 643
rect 6889 609 6922 643
rect 6822 575 6922 609
rect 6822 541 6855 575
rect 6889 541 6922 575
rect 6822 458 6922 541
rect -2522 425 6922 458
rect -2522 391 -2339 425
rect -2305 391 -2271 425
rect -2237 391 -2203 425
rect -2169 391 -2135 425
rect -2101 391 -2067 425
rect -2033 391 -1999 425
rect -1965 391 -1931 425
rect -1897 391 -1863 425
rect -1829 391 -1795 425
rect -1761 391 -1727 425
rect -1693 391 -1659 425
rect -1625 391 -1591 425
rect -1557 391 -1523 425
rect -1489 391 -1455 425
rect -1421 391 -1387 425
rect -1353 391 -1319 425
rect -1285 391 -1251 425
rect -1217 391 -1183 425
rect -1149 391 -1115 425
rect -1081 391 -1047 425
rect -1013 391 -979 425
rect -945 391 -911 425
rect -877 391 -843 425
rect -809 391 -775 425
rect -741 391 -707 425
rect -673 391 -639 425
rect -605 391 -571 425
rect -537 391 -503 425
rect -469 391 -435 425
rect -401 391 -367 425
rect -333 391 -299 425
rect -265 391 -231 425
rect -197 391 -163 425
rect -129 391 -95 425
rect -61 391 -27 425
rect 7 391 41 425
rect 75 391 109 425
rect 143 391 177 425
rect 211 391 245 425
rect 279 391 313 425
rect 347 391 381 425
rect 415 391 449 425
rect 483 391 517 425
rect 551 391 585 425
rect 619 391 653 425
rect 687 391 721 425
rect 755 391 789 425
rect 823 391 857 425
rect 891 391 925 425
rect 959 391 993 425
rect 1027 391 1061 425
rect 1095 391 1129 425
rect 1163 391 1197 425
rect 1231 391 1265 425
rect 1299 391 1333 425
rect 1367 391 1401 425
rect 1435 391 1469 425
rect 1503 391 1537 425
rect 1571 391 1605 425
rect 1639 391 1673 425
rect 1707 391 1741 425
rect 1775 391 1809 425
rect 1843 391 1877 425
rect 1911 391 1945 425
rect 1979 391 2013 425
rect 2047 391 2081 425
rect 2115 391 2149 425
rect 2183 391 2217 425
rect 2251 391 2285 425
rect 2319 391 2353 425
rect 2387 391 2421 425
rect 2455 391 2489 425
rect 2523 391 2557 425
rect 2591 391 2625 425
rect 2659 391 2693 425
rect 2727 391 2761 425
rect 2795 391 2829 425
rect 2863 391 2897 425
rect 2931 391 2965 425
rect 2999 391 3033 425
rect 3067 391 3101 425
rect 3135 391 3169 425
rect 3203 391 3237 425
rect 3271 391 3305 425
rect 3339 391 3373 425
rect 3407 391 3441 425
rect 3475 391 3509 425
rect 3543 391 3577 425
rect 3611 391 3645 425
rect 3679 391 3713 425
rect 3747 391 3781 425
rect 3815 391 3849 425
rect 3883 391 3917 425
rect 3951 391 3985 425
rect 4019 391 4053 425
rect 4087 391 4121 425
rect 4155 391 4189 425
rect 4223 391 4257 425
rect 4291 391 4325 425
rect 4359 391 4393 425
rect 4427 391 4461 425
rect 4495 391 4529 425
rect 4563 391 4597 425
rect 4631 391 4665 425
rect 4699 391 4733 425
rect 4767 391 4801 425
rect 4835 391 4869 425
rect 4903 391 4937 425
rect 4971 391 5005 425
rect 5039 391 5073 425
rect 5107 391 5141 425
rect 5175 391 5209 425
rect 5243 391 5277 425
rect 5311 391 5345 425
rect 5379 391 5413 425
rect 5447 391 5481 425
rect 5515 391 5549 425
rect 5583 391 5617 425
rect 5651 391 5685 425
rect 5719 391 5753 425
rect 5787 391 5821 425
rect 5855 391 5889 425
rect 5923 391 5957 425
rect 5991 391 6025 425
rect 6059 391 6093 425
rect 6127 391 6161 425
rect 6195 391 6229 425
rect 6263 391 6297 425
rect 6331 391 6365 425
rect 6399 391 6433 425
rect 6467 391 6501 425
rect 6535 391 6569 425
rect 6603 391 6637 425
rect 6671 391 6705 425
rect 6739 391 6922 425
rect -2522 358 6922 391
<< psubdiffcont >>
rect -2339 -1585 -2305 -1551
rect -2271 -1585 -2237 -1551
rect -2203 -1585 -2169 -1551
rect -2135 -1585 -2101 -1551
rect -2067 -1585 -2033 -1551
rect -1999 -1585 -1965 -1551
rect -1931 -1585 -1897 -1551
rect -1863 -1585 -1829 -1551
rect -1795 -1585 -1761 -1551
rect -1727 -1585 -1693 -1551
rect -1659 -1585 -1625 -1551
rect -1591 -1585 -1557 -1551
rect -1523 -1585 -1489 -1551
rect -1455 -1585 -1421 -1551
rect -1387 -1585 -1353 -1551
rect -1319 -1585 -1285 -1551
rect -1251 -1585 -1217 -1551
rect -1183 -1585 -1149 -1551
rect -1115 -1585 -1081 -1551
rect -1047 -1585 -1013 -1551
rect -979 -1585 -945 -1551
rect -911 -1585 -877 -1551
rect -843 -1585 -809 -1551
rect -775 -1585 -741 -1551
rect -707 -1585 -673 -1551
rect -639 -1585 -605 -1551
rect -571 -1585 -537 -1551
rect -503 -1585 -469 -1551
rect -435 -1585 -401 -1551
rect -367 -1585 -333 -1551
rect -299 -1585 -265 -1551
rect -231 -1585 -197 -1551
rect -163 -1585 -129 -1551
rect -95 -1585 -61 -1551
rect -27 -1585 7 -1551
rect 41 -1585 75 -1551
rect 109 -1585 143 -1551
rect 177 -1585 211 -1551
rect 245 -1585 279 -1551
rect 313 -1585 347 -1551
rect 381 -1585 415 -1551
rect 449 -1585 483 -1551
rect 517 -1585 551 -1551
rect 585 -1585 619 -1551
rect 653 -1585 687 -1551
rect 721 -1585 755 -1551
rect 789 -1585 823 -1551
rect 857 -1585 891 -1551
rect 925 -1585 959 -1551
rect 993 -1585 1027 -1551
rect 1061 -1585 1095 -1551
rect 1129 -1585 1163 -1551
rect 1197 -1585 1231 -1551
rect 1265 -1585 1299 -1551
rect 1333 -1585 1367 -1551
rect 1401 -1585 1435 -1551
rect 1469 -1585 1503 -1551
rect 1537 -1585 1571 -1551
rect 1605 -1585 1639 -1551
rect 1673 -1585 1707 -1551
rect 1741 -1585 1775 -1551
rect 1809 -1585 1843 -1551
rect 1877 -1585 1911 -1551
rect 1945 -1585 1979 -1551
rect 2013 -1585 2047 -1551
rect 2081 -1585 2115 -1551
rect 2149 -1585 2183 -1551
rect 2217 -1585 2251 -1551
rect 2285 -1585 2319 -1551
rect 2353 -1585 2387 -1551
rect 2421 -1585 2455 -1551
rect 2489 -1585 2523 -1551
rect 2557 -1585 2591 -1551
rect 2625 -1585 2659 -1551
rect 2693 -1585 2727 -1551
rect 2761 -1585 2795 -1551
rect 2829 -1585 2863 -1551
rect 2897 -1585 2931 -1551
rect 2965 -1585 2999 -1551
rect 3033 -1585 3067 -1551
rect 3101 -1585 3135 -1551
rect 3169 -1585 3203 -1551
rect 3237 -1585 3271 -1551
rect 3305 -1585 3339 -1551
rect 3373 -1585 3407 -1551
rect 3441 -1585 3475 -1551
rect 3509 -1585 3543 -1551
rect 3577 -1585 3611 -1551
rect 3645 -1585 3679 -1551
rect 3713 -1585 3747 -1551
rect 3781 -1585 3815 -1551
rect 3849 -1585 3883 -1551
rect 3917 -1585 3951 -1551
rect 3985 -1585 4019 -1551
rect 4053 -1585 4087 -1551
rect 4121 -1585 4155 -1551
rect 4189 -1585 4223 -1551
rect 4257 -1585 4291 -1551
rect 4325 -1585 4359 -1551
rect 4393 -1585 4427 -1551
rect 4461 -1585 4495 -1551
rect 4529 -1585 4563 -1551
rect 4597 -1585 4631 -1551
rect 4665 -1585 4699 -1551
rect 4733 -1585 4767 -1551
rect 4801 -1585 4835 -1551
rect 4869 -1585 4903 -1551
rect 4937 -1585 4971 -1551
rect 5005 -1585 5039 -1551
rect 5073 -1585 5107 -1551
rect 5141 -1585 5175 -1551
rect 5209 -1585 5243 -1551
rect 5277 -1585 5311 -1551
rect 5345 -1585 5379 -1551
rect 5413 -1585 5447 -1551
rect 5481 -1585 5515 -1551
rect 5549 -1585 5583 -1551
rect 5617 -1585 5651 -1551
rect 5685 -1585 5719 -1551
rect 5753 -1585 5787 -1551
rect 5821 -1585 5855 -1551
rect 5889 -1585 5923 -1551
rect 5957 -1585 5991 -1551
rect 6025 -1585 6059 -1551
rect 6093 -1585 6127 -1551
rect 6161 -1585 6195 -1551
rect 6229 -1585 6263 -1551
rect 6297 -1585 6331 -1551
rect 6365 -1585 6399 -1551
rect 6433 -1585 6467 -1551
rect 6501 -1585 6535 -1551
rect 6569 -1585 6603 -1551
rect 6637 -1585 6671 -1551
rect 6705 -1585 6739 -1551
rect -2489 -1715 -2455 -1681
rect -2489 -1783 -2455 -1749
rect -2489 -1851 -2455 -1817
rect -2489 -1919 -2455 -1885
rect -2489 -1987 -2455 -1953
rect -2489 -2055 -2455 -2021
rect -2489 -2123 -2455 -2089
rect -2489 -2191 -2455 -2157
rect -2489 -2259 -2455 -2225
rect -2489 -2327 -2455 -2293
rect -2489 -2395 -2455 -2361
rect -2489 -2463 -2455 -2429
rect -2489 -2531 -2455 -2497
rect -2489 -2599 -2455 -2565
rect -2489 -2667 -2455 -2633
rect -2489 -2735 -2455 -2701
rect -2489 -2803 -2455 -2769
rect -2489 -2871 -2455 -2837
rect -2489 -2939 -2455 -2905
rect -2489 -3007 -2455 -2973
rect -2489 -3075 -2455 -3041
rect -2489 -3143 -2455 -3109
rect -2489 -3211 -2455 -3177
rect -2489 -3279 -2455 -3245
rect -2489 -3347 -2455 -3313
rect -2489 -3415 -2455 -3381
rect -2489 -3483 -2455 -3449
rect -2489 -3551 -2455 -3517
rect -2489 -3619 -2455 -3585
rect 6855 -1715 6889 -1681
rect 6855 -1783 6889 -1749
rect 6855 -1851 6889 -1817
rect 6855 -1919 6889 -1885
rect 6855 -1987 6889 -1953
rect 6855 -2055 6889 -2021
rect 6855 -2123 6889 -2089
rect 6855 -2191 6889 -2157
rect 6855 -2259 6889 -2225
rect 6855 -2327 6889 -2293
rect 6855 -2395 6889 -2361
rect 6855 -2463 6889 -2429
rect 6855 -2531 6889 -2497
rect 6855 -2599 6889 -2565
rect 6855 -2667 6889 -2633
rect 6855 -2735 6889 -2701
rect 6855 -2803 6889 -2769
rect 6855 -2871 6889 -2837
rect 6855 -2939 6889 -2905
rect 6855 -3007 6889 -2973
rect 6855 -3075 6889 -3041
rect 6855 -3143 6889 -3109
rect 6855 -3211 6889 -3177
rect 6855 -3279 6889 -3245
rect 6855 -3347 6889 -3313
rect 6855 -3415 6889 -3381
rect 6855 -3483 6889 -3449
rect 6855 -3551 6889 -3517
rect 6855 -3619 6889 -3585
rect -2339 -3749 -2305 -3715
rect -2271 -3749 -2237 -3715
rect -2203 -3749 -2169 -3715
rect -2135 -3749 -2101 -3715
rect -2067 -3749 -2033 -3715
rect -1999 -3749 -1965 -3715
rect -1931 -3749 -1897 -3715
rect -1863 -3749 -1829 -3715
rect -1795 -3749 -1761 -3715
rect -1727 -3749 -1693 -3715
rect -1659 -3749 -1625 -3715
rect -1591 -3749 -1557 -3715
rect -1523 -3749 -1489 -3715
rect -1455 -3749 -1421 -3715
rect -1387 -3749 -1353 -3715
rect -1319 -3749 -1285 -3715
rect -1251 -3749 -1217 -3715
rect -1183 -3749 -1149 -3715
rect -1115 -3749 -1081 -3715
rect -1047 -3749 -1013 -3715
rect -979 -3749 -945 -3715
rect -911 -3749 -877 -3715
rect -843 -3749 -809 -3715
rect -775 -3749 -741 -3715
rect -707 -3749 -673 -3715
rect -639 -3749 -605 -3715
rect -571 -3749 -537 -3715
rect -503 -3749 -469 -3715
rect -435 -3749 -401 -3715
rect -367 -3749 -333 -3715
rect -299 -3749 -265 -3715
rect -231 -3749 -197 -3715
rect -163 -3749 -129 -3715
rect -95 -3749 -61 -3715
rect -27 -3749 7 -3715
rect 41 -3749 75 -3715
rect 109 -3749 143 -3715
rect 177 -3749 211 -3715
rect 245 -3749 279 -3715
rect 313 -3749 347 -3715
rect 381 -3749 415 -3715
rect 449 -3749 483 -3715
rect 517 -3749 551 -3715
rect 585 -3749 619 -3715
rect 653 -3749 687 -3715
rect 721 -3749 755 -3715
rect 789 -3749 823 -3715
rect 857 -3749 891 -3715
rect 925 -3749 959 -3715
rect 993 -3749 1027 -3715
rect 1061 -3749 1095 -3715
rect 1129 -3749 1163 -3715
rect 1197 -3749 1231 -3715
rect 1265 -3749 1299 -3715
rect 1333 -3749 1367 -3715
rect 1401 -3749 1435 -3715
rect 1469 -3749 1503 -3715
rect 1537 -3749 1571 -3715
rect 1605 -3749 1639 -3715
rect 1673 -3749 1707 -3715
rect 1741 -3749 1775 -3715
rect 1809 -3749 1843 -3715
rect 1877 -3749 1911 -3715
rect 1945 -3749 1979 -3715
rect 2013 -3749 2047 -3715
rect 2081 -3749 2115 -3715
rect 2149 -3749 2183 -3715
rect 2217 -3749 2251 -3715
rect 2285 -3749 2319 -3715
rect 2353 -3749 2387 -3715
rect 2421 -3749 2455 -3715
rect 2489 -3749 2523 -3715
rect 2557 -3749 2591 -3715
rect 2625 -3749 2659 -3715
rect 2693 -3749 2727 -3715
rect 2761 -3749 2795 -3715
rect 2829 -3749 2863 -3715
rect 2897 -3749 2931 -3715
rect 2965 -3749 2999 -3715
rect 3033 -3749 3067 -3715
rect 3101 -3749 3135 -3715
rect 3169 -3749 3203 -3715
rect 3237 -3749 3271 -3715
rect 3305 -3749 3339 -3715
rect 3373 -3749 3407 -3715
rect 3441 -3749 3475 -3715
rect 3509 -3749 3543 -3715
rect 3577 -3749 3611 -3715
rect 3645 -3749 3679 -3715
rect 3713 -3749 3747 -3715
rect 3781 -3749 3815 -3715
rect 3849 -3749 3883 -3715
rect 3917 -3749 3951 -3715
rect 3985 -3749 4019 -3715
rect 4053 -3749 4087 -3715
rect 4121 -3749 4155 -3715
rect 4189 -3749 4223 -3715
rect 4257 -3749 4291 -3715
rect 4325 -3749 4359 -3715
rect 4393 -3749 4427 -3715
rect 4461 -3749 4495 -3715
rect 4529 -3749 4563 -3715
rect 4597 -3749 4631 -3715
rect 4665 -3749 4699 -3715
rect 4733 -3749 4767 -3715
rect 4801 -3749 4835 -3715
rect 4869 -3749 4903 -3715
rect 4937 -3749 4971 -3715
rect 5005 -3749 5039 -3715
rect 5073 -3749 5107 -3715
rect 5141 -3749 5175 -3715
rect 5209 -3749 5243 -3715
rect 5277 -3749 5311 -3715
rect 5345 -3749 5379 -3715
rect 5413 -3749 5447 -3715
rect 5481 -3749 5515 -3715
rect 5549 -3749 5583 -3715
rect 5617 -3749 5651 -3715
rect 5685 -3749 5719 -3715
rect 5753 -3749 5787 -3715
rect 5821 -3749 5855 -3715
rect 5889 -3749 5923 -3715
rect 5957 -3749 5991 -3715
rect 6025 -3749 6059 -3715
rect 6093 -3749 6127 -3715
rect 6161 -3749 6195 -3715
rect 6229 -3749 6263 -3715
rect 6297 -3749 6331 -3715
rect 6365 -3749 6399 -3715
rect 6433 -3749 6467 -3715
rect 6501 -3749 6535 -3715
rect 6569 -3749 6603 -3715
rect 6637 -3749 6671 -3715
rect 6705 -3749 6739 -3715
<< nsubdiffcont >>
rect -2339 2595 -2305 2629
rect -2271 2595 -2237 2629
rect -2203 2595 -2169 2629
rect -2135 2595 -2101 2629
rect -2067 2595 -2033 2629
rect -1999 2595 -1965 2629
rect -1931 2595 -1897 2629
rect -1863 2595 -1829 2629
rect -1795 2595 -1761 2629
rect -1727 2595 -1693 2629
rect -1659 2595 -1625 2629
rect -1591 2595 -1557 2629
rect -1523 2595 -1489 2629
rect -1455 2595 -1421 2629
rect -1387 2595 -1353 2629
rect -1319 2595 -1285 2629
rect -1251 2595 -1217 2629
rect -1183 2595 -1149 2629
rect -1115 2595 -1081 2629
rect -1047 2595 -1013 2629
rect -979 2595 -945 2629
rect -911 2595 -877 2629
rect -843 2595 -809 2629
rect -775 2595 -741 2629
rect -707 2595 -673 2629
rect -639 2595 -605 2629
rect -571 2595 -537 2629
rect -503 2595 -469 2629
rect -435 2595 -401 2629
rect -367 2595 -333 2629
rect -299 2595 -265 2629
rect -231 2595 -197 2629
rect -163 2595 -129 2629
rect -95 2595 -61 2629
rect -27 2595 7 2629
rect 41 2595 75 2629
rect 109 2595 143 2629
rect 177 2595 211 2629
rect 245 2595 279 2629
rect 313 2595 347 2629
rect 381 2595 415 2629
rect 449 2595 483 2629
rect 517 2595 551 2629
rect 585 2595 619 2629
rect 653 2595 687 2629
rect 721 2595 755 2629
rect 789 2595 823 2629
rect 857 2595 891 2629
rect 925 2595 959 2629
rect 993 2595 1027 2629
rect 1061 2595 1095 2629
rect 1129 2595 1163 2629
rect 1197 2595 1231 2629
rect 1265 2595 1299 2629
rect 1333 2595 1367 2629
rect 1401 2595 1435 2629
rect 1469 2595 1503 2629
rect 1537 2595 1571 2629
rect 1605 2595 1639 2629
rect 1673 2595 1707 2629
rect 1741 2595 1775 2629
rect 1809 2595 1843 2629
rect 1877 2595 1911 2629
rect 1945 2595 1979 2629
rect 2013 2595 2047 2629
rect 2081 2595 2115 2629
rect 2149 2595 2183 2629
rect 2217 2595 2251 2629
rect 2285 2595 2319 2629
rect 2353 2595 2387 2629
rect 2421 2595 2455 2629
rect 2489 2595 2523 2629
rect 2557 2595 2591 2629
rect 2625 2595 2659 2629
rect 2693 2595 2727 2629
rect 2761 2595 2795 2629
rect 2829 2595 2863 2629
rect 2897 2595 2931 2629
rect 2965 2595 2999 2629
rect 3033 2595 3067 2629
rect 3101 2595 3135 2629
rect 3169 2595 3203 2629
rect 3237 2595 3271 2629
rect 3305 2595 3339 2629
rect 3373 2595 3407 2629
rect 3441 2595 3475 2629
rect 3509 2595 3543 2629
rect 3577 2595 3611 2629
rect 3645 2595 3679 2629
rect 3713 2595 3747 2629
rect 3781 2595 3815 2629
rect 3849 2595 3883 2629
rect 3917 2595 3951 2629
rect 3985 2595 4019 2629
rect 4053 2595 4087 2629
rect 4121 2595 4155 2629
rect 4189 2595 4223 2629
rect 4257 2595 4291 2629
rect 4325 2595 4359 2629
rect 4393 2595 4427 2629
rect 4461 2595 4495 2629
rect 4529 2595 4563 2629
rect 4597 2595 4631 2629
rect 4665 2595 4699 2629
rect 4733 2595 4767 2629
rect 4801 2595 4835 2629
rect 4869 2595 4903 2629
rect 4937 2595 4971 2629
rect 5005 2595 5039 2629
rect 5073 2595 5107 2629
rect 5141 2595 5175 2629
rect 5209 2595 5243 2629
rect 5277 2595 5311 2629
rect 5345 2595 5379 2629
rect 5413 2595 5447 2629
rect 5481 2595 5515 2629
rect 5549 2595 5583 2629
rect 5617 2595 5651 2629
rect 5685 2595 5719 2629
rect 5753 2595 5787 2629
rect 5821 2595 5855 2629
rect 5889 2595 5923 2629
rect 5957 2595 5991 2629
rect 6025 2595 6059 2629
rect 6093 2595 6127 2629
rect 6161 2595 6195 2629
rect 6229 2595 6263 2629
rect 6297 2595 6331 2629
rect 6365 2595 6399 2629
rect 6433 2595 6467 2629
rect 6501 2595 6535 2629
rect 6569 2595 6603 2629
rect 6637 2595 6671 2629
rect 6705 2595 6739 2629
rect -2489 2445 -2455 2479
rect -2489 2377 -2455 2411
rect -2489 2309 -2455 2343
rect -2489 2241 -2455 2275
rect -2489 2173 -2455 2207
rect -2489 2105 -2455 2139
rect -2489 2037 -2455 2071
rect -2489 1969 -2455 2003
rect -2489 1901 -2455 1935
rect -2489 1833 -2455 1867
rect -2489 1765 -2455 1799
rect -2489 1697 -2455 1731
rect -2489 1629 -2455 1663
rect -2489 1561 -2455 1595
rect -2489 1493 -2455 1527
rect -2489 1425 -2455 1459
rect -2489 1357 -2455 1391
rect -2489 1289 -2455 1323
rect -2489 1221 -2455 1255
rect -2489 1153 -2455 1187
rect -2489 1085 -2455 1119
rect -2489 1017 -2455 1051
rect -2489 949 -2455 983
rect -2489 881 -2455 915
rect -2489 813 -2455 847
rect -2489 745 -2455 779
rect -2489 677 -2455 711
rect -2489 609 -2455 643
rect -2489 541 -2455 575
rect 6855 2445 6889 2479
rect 6855 2377 6889 2411
rect 6855 2309 6889 2343
rect 6855 2241 6889 2275
rect 6855 2173 6889 2207
rect 6855 2105 6889 2139
rect 6855 2037 6889 2071
rect 6855 1969 6889 2003
rect 6855 1901 6889 1935
rect 6855 1833 6889 1867
rect 6855 1765 6889 1799
rect 6855 1697 6889 1731
rect 6855 1629 6889 1663
rect 6855 1561 6889 1595
rect 6855 1493 6889 1527
rect 6855 1425 6889 1459
rect 6855 1357 6889 1391
rect 6855 1289 6889 1323
rect 6855 1221 6889 1255
rect 6855 1153 6889 1187
rect 6855 1085 6889 1119
rect 6855 1017 6889 1051
rect 6855 949 6889 983
rect 6855 881 6889 915
rect 6855 813 6889 847
rect 6855 745 6889 779
rect 6855 677 6889 711
rect 6855 609 6889 643
rect 6855 541 6889 575
rect -2339 391 -2305 425
rect -2271 391 -2237 425
rect -2203 391 -2169 425
rect -2135 391 -2101 425
rect -2067 391 -2033 425
rect -1999 391 -1965 425
rect -1931 391 -1897 425
rect -1863 391 -1829 425
rect -1795 391 -1761 425
rect -1727 391 -1693 425
rect -1659 391 -1625 425
rect -1591 391 -1557 425
rect -1523 391 -1489 425
rect -1455 391 -1421 425
rect -1387 391 -1353 425
rect -1319 391 -1285 425
rect -1251 391 -1217 425
rect -1183 391 -1149 425
rect -1115 391 -1081 425
rect -1047 391 -1013 425
rect -979 391 -945 425
rect -911 391 -877 425
rect -843 391 -809 425
rect -775 391 -741 425
rect -707 391 -673 425
rect -639 391 -605 425
rect -571 391 -537 425
rect -503 391 -469 425
rect -435 391 -401 425
rect -367 391 -333 425
rect -299 391 -265 425
rect -231 391 -197 425
rect -163 391 -129 425
rect -95 391 -61 425
rect -27 391 7 425
rect 41 391 75 425
rect 109 391 143 425
rect 177 391 211 425
rect 245 391 279 425
rect 313 391 347 425
rect 381 391 415 425
rect 449 391 483 425
rect 517 391 551 425
rect 585 391 619 425
rect 653 391 687 425
rect 721 391 755 425
rect 789 391 823 425
rect 857 391 891 425
rect 925 391 959 425
rect 993 391 1027 425
rect 1061 391 1095 425
rect 1129 391 1163 425
rect 1197 391 1231 425
rect 1265 391 1299 425
rect 1333 391 1367 425
rect 1401 391 1435 425
rect 1469 391 1503 425
rect 1537 391 1571 425
rect 1605 391 1639 425
rect 1673 391 1707 425
rect 1741 391 1775 425
rect 1809 391 1843 425
rect 1877 391 1911 425
rect 1945 391 1979 425
rect 2013 391 2047 425
rect 2081 391 2115 425
rect 2149 391 2183 425
rect 2217 391 2251 425
rect 2285 391 2319 425
rect 2353 391 2387 425
rect 2421 391 2455 425
rect 2489 391 2523 425
rect 2557 391 2591 425
rect 2625 391 2659 425
rect 2693 391 2727 425
rect 2761 391 2795 425
rect 2829 391 2863 425
rect 2897 391 2931 425
rect 2965 391 2999 425
rect 3033 391 3067 425
rect 3101 391 3135 425
rect 3169 391 3203 425
rect 3237 391 3271 425
rect 3305 391 3339 425
rect 3373 391 3407 425
rect 3441 391 3475 425
rect 3509 391 3543 425
rect 3577 391 3611 425
rect 3645 391 3679 425
rect 3713 391 3747 425
rect 3781 391 3815 425
rect 3849 391 3883 425
rect 3917 391 3951 425
rect 3985 391 4019 425
rect 4053 391 4087 425
rect 4121 391 4155 425
rect 4189 391 4223 425
rect 4257 391 4291 425
rect 4325 391 4359 425
rect 4393 391 4427 425
rect 4461 391 4495 425
rect 4529 391 4563 425
rect 4597 391 4631 425
rect 4665 391 4699 425
rect 4733 391 4767 425
rect 4801 391 4835 425
rect 4869 391 4903 425
rect 4937 391 4971 425
rect 5005 391 5039 425
rect 5073 391 5107 425
rect 5141 391 5175 425
rect 5209 391 5243 425
rect 5277 391 5311 425
rect 5345 391 5379 425
rect 5413 391 5447 425
rect 5481 391 5515 425
rect 5549 391 5583 425
rect 5617 391 5651 425
rect 5685 391 5719 425
rect 5753 391 5787 425
rect 5821 391 5855 425
rect 5889 391 5923 425
rect 5957 391 5991 425
rect 6025 391 6059 425
rect 6093 391 6127 425
rect 6161 391 6195 425
rect 6229 391 6263 425
rect 6297 391 6331 425
rect 6365 391 6399 425
rect 6433 391 6467 425
rect 6501 391 6535 425
rect 6569 391 6603 425
rect 6637 391 6671 425
rect 6705 391 6739 425
<< locali >>
rect -2522 2629 6922 2662
rect -2522 2595 -2389 2629
rect -2355 2595 -2339 2629
rect -2283 2595 -2271 2629
rect -2211 2595 -2203 2629
rect -2139 2595 -2135 2629
rect -2033 2595 -2029 2629
rect -1965 2595 -1957 2629
rect -1897 2595 -1885 2629
rect -1829 2595 -1813 2629
rect -1761 2595 -1741 2629
rect -1693 2595 -1669 2629
rect -1625 2595 -1597 2629
rect -1557 2595 -1525 2629
rect -1489 2595 -1455 2629
rect -1419 2595 -1387 2629
rect -1347 2595 -1319 2629
rect -1275 2595 -1251 2629
rect -1203 2595 -1183 2629
rect -1131 2595 -1115 2629
rect -1059 2595 -1047 2629
rect -987 2595 -979 2629
rect -915 2595 -911 2629
rect -809 2595 -805 2629
rect -741 2595 -733 2629
rect -673 2595 -661 2629
rect -605 2595 -589 2629
rect -537 2595 -517 2629
rect -469 2595 -445 2629
rect -401 2595 -373 2629
rect -333 2595 -301 2629
rect -265 2595 -231 2629
rect -195 2595 -163 2629
rect -123 2595 -95 2629
rect -51 2595 -27 2629
rect 21 2595 41 2629
rect 93 2595 109 2629
rect 165 2595 177 2629
rect 237 2595 245 2629
rect 309 2595 313 2629
rect 415 2595 419 2629
rect 483 2595 491 2629
rect 551 2595 563 2629
rect 619 2595 635 2629
rect 687 2595 707 2629
rect 755 2595 779 2629
rect 823 2595 851 2629
rect 891 2595 923 2629
rect 959 2595 993 2629
rect 1029 2595 1061 2629
rect 1101 2595 1129 2629
rect 1173 2595 1197 2629
rect 1245 2595 1265 2629
rect 1317 2595 1333 2629
rect 1389 2595 1401 2629
rect 1461 2595 1469 2629
rect 1533 2595 1537 2629
rect 1639 2595 1643 2629
rect 1707 2595 1715 2629
rect 1775 2595 1787 2629
rect 1843 2595 1859 2629
rect 1911 2595 1931 2629
rect 1979 2595 2003 2629
rect 2047 2595 2075 2629
rect 2115 2595 2147 2629
rect 2183 2595 2217 2629
rect 2253 2595 2285 2629
rect 2325 2595 2353 2629
rect 2397 2595 2421 2629
rect 2469 2595 2489 2629
rect 2541 2595 2557 2629
rect 2613 2595 2625 2629
rect 2685 2595 2693 2629
rect 2757 2595 2761 2629
rect 2863 2595 2867 2629
rect 2931 2595 2939 2629
rect 2999 2595 3011 2629
rect 3067 2595 3083 2629
rect 3135 2595 3155 2629
rect 3203 2595 3227 2629
rect 3271 2595 3299 2629
rect 3339 2595 3371 2629
rect 3407 2595 3441 2629
rect 3477 2595 3509 2629
rect 3549 2595 3577 2629
rect 3621 2595 3645 2629
rect 3693 2595 3713 2629
rect 3765 2595 3781 2629
rect 3837 2595 3849 2629
rect 3909 2595 3917 2629
rect 3981 2595 3985 2629
rect 4087 2595 4091 2629
rect 4155 2595 4163 2629
rect 4223 2595 4235 2629
rect 4291 2595 4307 2629
rect 4359 2595 4379 2629
rect 4427 2595 4451 2629
rect 4495 2595 4523 2629
rect 4563 2595 4595 2629
rect 4631 2595 4665 2629
rect 4701 2595 4733 2629
rect 4773 2595 4801 2629
rect 4845 2595 4869 2629
rect 4917 2595 4937 2629
rect 4989 2595 5005 2629
rect 5061 2595 5073 2629
rect 5133 2595 5141 2629
rect 5205 2595 5209 2629
rect 5311 2595 5315 2629
rect 5379 2595 5387 2629
rect 5447 2595 5459 2629
rect 5515 2595 5531 2629
rect 5583 2595 5603 2629
rect 5651 2595 5675 2629
rect 5719 2595 5747 2629
rect 5787 2595 5819 2629
rect 5855 2595 5889 2629
rect 5925 2595 5957 2629
rect 5997 2595 6025 2629
rect 6069 2595 6093 2629
rect 6141 2595 6161 2629
rect 6213 2595 6229 2629
rect 6285 2595 6297 2629
rect 6357 2595 6365 2629
rect 6429 2595 6433 2629
rect 6535 2595 6539 2629
rect 6603 2595 6611 2629
rect 6671 2595 6683 2629
rect 6739 2595 6755 2629
rect 6789 2595 6922 2629
rect -2522 2562 6922 2595
rect -2522 2479 -2422 2562
rect -2522 2445 -2489 2479
rect -2455 2445 -2422 2479
rect -2522 2427 -2422 2445
rect -2522 2377 -2489 2427
rect -2455 2377 -2422 2427
rect -2522 2355 -2422 2377
rect -2522 2309 -2489 2355
rect -2455 2309 -2422 2355
rect -2522 2283 -2422 2309
rect -2522 2241 -2489 2283
rect -2455 2241 -2422 2283
rect -2522 2211 -2422 2241
rect -2522 2173 -2489 2211
rect -2455 2173 -2422 2211
rect -2522 2139 -2422 2173
rect -2522 2105 -2489 2139
rect -2455 2105 -2422 2139
rect -2522 2071 -2422 2105
rect -2522 2033 -2489 2071
rect -2455 2033 -2422 2071
rect -2522 2003 -2422 2033
rect -2522 1961 -2489 2003
rect -2455 1961 -2422 2003
rect -2522 1935 -2422 1961
rect -2522 1889 -2489 1935
rect -2455 1889 -2422 1935
rect -2522 1867 -2422 1889
rect -2522 1817 -2489 1867
rect -2455 1817 -2422 1867
rect -2522 1799 -2422 1817
rect -2522 1745 -2489 1799
rect -2455 1745 -2422 1799
rect -2522 1731 -2422 1745
rect -2522 1673 -2489 1731
rect -2455 1673 -2422 1731
rect -2522 1663 -2422 1673
rect -2522 1601 -2489 1663
rect -2455 1601 -2422 1663
rect -2522 1595 -2422 1601
rect -2522 1529 -2489 1595
rect -2455 1529 -2422 1595
rect -2522 1527 -2422 1529
rect -2522 1493 -2489 1527
rect -2455 1493 -2422 1527
rect -2522 1491 -2422 1493
rect -2522 1425 -2489 1491
rect -2455 1425 -2422 1491
rect -2522 1419 -2422 1425
rect -2522 1357 -2489 1419
rect -2455 1357 -2422 1419
rect -2522 1347 -2422 1357
rect -2522 1289 -2489 1347
rect -2455 1289 -2422 1347
rect -2522 1275 -2422 1289
rect -2522 1221 -2489 1275
rect -2455 1221 -2422 1275
rect -2522 1203 -2422 1221
rect -2522 1153 -2489 1203
rect -2455 1153 -2422 1203
rect -2522 1131 -2422 1153
rect -2522 1085 -2489 1131
rect -2455 1085 -2422 1131
rect -2522 1059 -2422 1085
rect -2522 1017 -2489 1059
rect -2455 1017 -2422 1059
rect -2522 987 -2422 1017
rect -2522 949 -2489 987
rect -2455 949 -2422 987
rect -2522 915 -2422 949
rect -2522 881 -2489 915
rect -2455 881 -2422 915
rect -2522 847 -2422 881
rect -2522 809 -2489 847
rect -2455 809 -2422 847
rect -2522 779 -2422 809
rect -2522 737 -2489 779
rect -2455 737 -2422 779
rect -2522 711 -2422 737
rect -2522 665 -2489 711
rect -2455 665 -2422 711
rect -2522 643 -2422 665
rect -2522 593 -2489 643
rect -2455 593 -2422 643
rect -2522 575 -2422 593
rect -2522 541 -2489 575
rect -2455 541 -2422 575
rect -2522 458 -2422 541
rect 6822 2479 6922 2562
rect 6822 2445 6855 2479
rect 6889 2445 6922 2479
rect 6822 2427 6922 2445
rect 6822 2377 6855 2427
rect 6889 2377 6922 2427
rect 6822 2355 6922 2377
rect 6822 2309 6855 2355
rect 6889 2309 6922 2355
rect 6822 2283 6922 2309
rect 6822 2241 6855 2283
rect 6889 2241 6922 2283
rect 6822 2211 6922 2241
rect 6822 2173 6855 2211
rect 6889 2173 6922 2211
rect 6822 2139 6922 2173
rect 6822 2105 6855 2139
rect 6889 2105 6922 2139
rect 6822 2071 6922 2105
rect 6822 2033 6855 2071
rect 6889 2033 6922 2071
rect 6822 2003 6922 2033
rect 6822 1961 6855 2003
rect 6889 1961 6922 2003
rect 6822 1935 6922 1961
rect 6822 1889 6855 1935
rect 6889 1889 6922 1935
rect 6822 1867 6922 1889
rect 6822 1817 6855 1867
rect 6889 1817 6922 1867
rect 6822 1799 6922 1817
rect 6822 1745 6855 1799
rect 6889 1745 6922 1799
rect 6822 1731 6922 1745
rect 6822 1673 6855 1731
rect 6889 1673 6922 1731
rect 6822 1663 6922 1673
rect 6822 1601 6855 1663
rect 6889 1601 6922 1663
rect 6822 1595 6922 1601
rect 6822 1529 6855 1595
rect 6889 1529 6922 1595
rect 6822 1527 6922 1529
rect 6822 1493 6855 1527
rect 6889 1493 6922 1527
rect 6822 1491 6922 1493
rect 6822 1425 6855 1491
rect 6889 1425 6922 1491
rect 6822 1419 6922 1425
rect 6822 1357 6855 1419
rect 6889 1357 6922 1419
rect 6822 1347 6922 1357
rect 6822 1289 6855 1347
rect 6889 1289 6922 1347
rect 6822 1275 6922 1289
rect 6822 1221 6855 1275
rect 6889 1221 6922 1275
rect 6822 1203 6922 1221
rect 6822 1153 6855 1203
rect 6889 1153 6922 1203
rect 6822 1131 6922 1153
rect 6822 1085 6855 1131
rect 6889 1085 6922 1131
rect 6822 1059 6922 1085
rect 6822 1017 6855 1059
rect 6889 1017 6922 1059
rect 6822 987 6922 1017
rect 6822 949 6855 987
rect 6889 949 6922 987
rect 6822 915 6922 949
rect 6822 881 6855 915
rect 6889 881 6922 915
rect 6822 847 6922 881
rect 6822 809 6855 847
rect 6889 809 6922 847
rect 6822 779 6922 809
rect 6822 737 6855 779
rect 6889 737 6922 779
rect 6822 711 6922 737
rect 6822 665 6855 711
rect 6889 665 6922 711
rect 6822 643 6922 665
rect 6822 593 6855 643
rect 6889 593 6922 643
rect 6822 575 6922 593
rect 6822 541 6855 575
rect 6889 541 6922 575
rect 6822 458 6922 541
rect -2522 425 6922 458
rect -2522 391 -2389 425
rect -2355 391 -2339 425
rect -2283 391 -2271 425
rect -2211 391 -2203 425
rect -2139 391 -2135 425
rect -2033 391 -2029 425
rect -1965 391 -1957 425
rect -1897 391 -1885 425
rect -1829 391 -1813 425
rect -1761 391 -1741 425
rect -1693 391 -1669 425
rect -1625 391 -1597 425
rect -1557 391 -1525 425
rect -1489 391 -1455 425
rect -1419 391 -1387 425
rect -1347 391 -1319 425
rect -1275 391 -1251 425
rect -1203 391 -1183 425
rect -1131 391 -1115 425
rect -1059 391 -1047 425
rect -987 391 -979 425
rect -915 391 -911 425
rect -809 391 -805 425
rect -741 391 -733 425
rect -673 391 -661 425
rect -605 391 -589 425
rect -537 391 -517 425
rect -469 391 -445 425
rect -401 391 -373 425
rect -333 391 -301 425
rect -265 391 -231 425
rect -195 391 -163 425
rect -123 391 -95 425
rect -51 391 -27 425
rect 21 391 41 425
rect 93 391 109 425
rect 165 391 177 425
rect 237 391 245 425
rect 309 391 313 425
rect 415 391 419 425
rect 483 391 491 425
rect 551 391 563 425
rect 619 391 635 425
rect 687 391 707 425
rect 755 391 779 425
rect 823 391 851 425
rect 891 391 923 425
rect 959 391 993 425
rect 1029 391 1061 425
rect 1101 391 1129 425
rect 1173 391 1197 425
rect 1245 391 1265 425
rect 1317 391 1333 425
rect 1389 391 1401 425
rect 1461 391 1469 425
rect 1533 391 1537 425
rect 1639 391 1643 425
rect 1707 391 1715 425
rect 1775 391 1787 425
rect 1843 391 1859 425
rect 1911 391 1931 425
rect 1979 391 2003 425
rect 2047 391 2075 425
rect 2115 391 2147 425
rect 2183 391 2217 425
rect 2253 391 2285 425
rect 2325 391 2353 425
rect 2397 391 2421 425
rect 2469 391 2489 425
rect 2541 391 2557 425
rect 2613 391 2625 425
rect 2685 391 2693 425
rect 2757 391 2761 425
rect 2863 391 2867 425
rect 2931 391 2939 425
rect 2999 391 3011 425
rect 3067 391 3083 425
rect 3135 391 3155 425
rect 3203 391 3227 425
rect 3271 391 3299 425
rect 3339 391 3371 425
rect 3407 391 3441 425
rect 3477 391 3509 425
rect 3549 391 3577 425
rect 3621 391 3645 425
rect 3693 391 3713 425
rect 3765 391 3781 425
rect 3837 391 3849 425
rect 3909 391 3917 425
rect 3981 391 3985 425
rect 4087 391 4091 425
rect 4155 391 4163 425
rect 4223 391 4235 425
rect 4291 391 4307 425
rect 4359 391 4379 425
rect 4427 391 4451 425
rect 4495 391 4523 425
rect 4563 391 4595 425
rect 4631 391 4665 425
rect 4701 391 4733 425
rect 4773 391 4801 425
rect 4845 391 4869 425
rect 4917 391 4937 425
rect 4989 391 5005 425
rect 5061 391 5073 425
rect 5133 391 5141 425
rect 5205 391 5209 425
rect 5311 391 5315 425
rect 5379 391 5387 425
rect 5447 391 5459 425
rect 5515 391 5531 425
rect 5583 391 5603 425
rect 5651 391 5675 425
rect 5719 391 5747 425
rect 5787 391 5819 425
rect 5855 391 5889 425
rect 5925 391 5957 425
rect 5997 391 6025 425
rect 6069 391 6093 425
rect 6141 391 6161 425
rect 6213 391 6229 425
rect 6285 391 6297 425
rect 6357 391 6365 425
rect 6429 391 6433 425
rect 6535 391 6539 425
rect 6603 391 6611 425
rect 6671 391 6683 425
rect 6739 391 6755 425
rect 6789 391 6922 425
rect -2522 358 6922 391
rect 3274 27 3308 46
rect 3274 -45 3308 -7
rect 3274 -117 3308 -79
rect 3274 -189 3308 -151
rect 3274 -261 3308 -223
rect 3274 -333 3308 -295
rect 3274 -405 3308 -367
rect -1782 -445 -1736 -442
rect -1782 -479 -1776 -445
rect -1742 -479 -1736 -445
rect 2674 -453 2714 -450
rect -1782 -482 -1736 -479
rect 208 -477 256 -470
rect 208 -511 215 -477
rect 249 -511 256 -477
rect 2674 -487 2677 -453
rect 2711 -487 2714 -453
rect 2674 -490 2714 -487
rect 3274 -477 3308 -439
rect 208 -518 256 -511
rect 3274 -530 3308 -511
rect 5050 26 5086 44
rect 5050 -8 5051 26
rect 5085 -8 5086 26
rect 5050 -46 5086 -8
rect 5050 -80 5051 -46
rect 5085 -80 5086 -46
rect 5050 -118 5086 -80
rect 5050 -152 5051 -118
rect 5085 -152 5086 -118
rect 5050 -190 5086 -152
rect 5050 -224 5051 -190
rect 5085 -224 5086 -190
rect 5050 -262 5086 -224
rect 5050 -296 5051 -262
rect 5085 -296 5086 -262
rect 5050 -334 5086 -296
rect 5050 -368 5051 -334
rect 5085 -368 5086 -334
rect 5050 -406 5086 -368
rect 5050 -440 5051 -406
rect 5085 -440 5086 -406
rect 5050 -478 5086 -440
rect 5050 -512 5051 -478
rect 5085 -512 5086 -478
rect 5050 -530 5086 -512
rect 5170 26 5206 44
rect 5170 -8 5171 26
rect 5205 -8 5206 26
rect 5170 -46 5206 -8
rect 5170 -80 5171 -46
rect 5205 -80 5206 -46
rect 5170 -118 5206 -80
rect 5170 -152 5171 -118
rect 5205 -152 5206 -118
rect 5170 -190 5206 -152
rect 5170 -224 5171 -190
rect 5205 -224 5206 -190
rect 5170 -262 5206 -224
rect 5170 -296 5171 -262
rect 5205 -296 5206 -262
rect 5170 -334 5206 -296
rect 5170 -368 5171 -334
rect 5205 -368 5206 -334
rect 5170 -406 5206 -368
rect 5170 -440 5171 -406
rect 5205 -440 5206 -406
rect 5170 -478 5206 -440
rect 5170 -512 5171 -478
rect 5205 -512 5206 -478
rect 5170 -530 5206 -512
rect 6172 26 6208 44
rect 6172 -8 6173 26
rect 6207 -8 6208 26
rect 6172 -46 6208 -8
rect 6172 -80 6173 -46
rect 6207 -80 6208 -46
rect 6172 -118 6208 -80
rect 6172 -152 6173 -118
rect 6207 -152 6208 -118
rect 6172 -190 6208 -152
rect 6172 -224 6173 -190
rect 6207 -224 6208 -190
rect 6172 -262 6208 -224
rect 6172 -296 6173 -262
rect 6207 -296 6208 -262
rect 6172 -334 6208 -296
rect 6172 -368 6173 -334
rect 6207 -368 6208 -334
rect 6172 -406 6208 -368
rect 6172 -440 6173 -406
rect 6207 -440 6208 -406
rect 6172 -478 6208 -440
rect 6172 -512 6173 -478
rect 6207 -512 6208 -478
rect 6172 -530 6208 -512
rect 442 -570 490 -562
rect 442 -574 492 -570
rect 442 -608 451 -574
rect 485 -608 492 -574
rect 442 -610 492 -608
rect 444 -612 492 -610
rect 2934 -655 2982 -648
rect -2044 -673 -1996 -666
rect -2044 -707 -2037 -673
rect -2003 -707 -1996 -673
rect -2044 -714 -1996 -707
rect -320 -675 -272 -668
rect -320 -709 -313 -675
rect -279 -709 -272 -675
rect 118 -671 166 -668
rect 118 -705 125 -671
rect 159 -705 166 -671
rect 118 -708 166 -705
rect 352 -672 400 -668
rect 352 -706 359 -672
rect 393 -706 400 -672
rect -320 -716 -272 -709
rect 352 -710 400 -706
rect 526 -672 574 -668
rect 526 -706 533 -672
rect 567 -706 574 -672
rect 526 -710 574 -706
rect 764 -671 812 -668
rect 764 -705 771 -671
rect 805 -705 812 -671
rect 764 -708 812 -705
rect 1204 -675 1252 -668
rect 1204 -709 1211 -675
rect 1245 -709 1252 -675
rect 2934 -689 2941 -655
rect 2975 -689 2982 -655
rect 2934 -696 2982 -689
rect 1204 -716 1252 -709
rect 676 -787 724 -780
rect 676 -821 683 -787
rect 717 -821 724 -787
rect 676 -828 724 -821
rect 3276 -869 3310 -852
rect 3276 -941 3310 -903
rect 3276 -1013 3310 -975
rect 3276 -1085 3310 -1047
rect 3276 -1157 3310 -1119
rect 3276 -1208 3310 -1191
rect 5052 -870 5086 -854
rect 5052 -942 5086 -904
rect 5052 -1014 5086 -976
rect 5052 -1086 5086 -1048
rect 5052 -1158 5086 -1120
rect 5052 -1208 5086 -1192
rect 5172 -870 5206 -854
rect 5172 -942 5206 -904
rect 5172 -1014 5206 -976
rect 5172 -1086 5206 -1048
rect 5172 -1158 5206 -1120
rect 5172 -1208 5206 -1192
rect 6174 -869 6208 -852
rect 6174 -941 6208 -903
rect 6174 -1013 6208 -975
rect 6174 -1085 6208 -1047
rect 6174 -1157 6208 -1119
rect 6174 -1208 6208 -1191
rect -2522 -1551 6922 -1518
rect -2522 -1585 -2389 -1551
rect -2355 -1585 -2339 -1551
rect -2283 -1585 -2271 -1551
rect -2211 -1585 -2203 -1551
rect -2139 -1585 -2135 -1551
rect -2033 -1585 -2029 -1551
rect -1965 -1585 -1957 -1551
rect -1897 -1585 -1885 -1551
rect -1829 -1585 -1813 -1551
rect -1761 -1585 -1741 -1551
rect -1693 -1585 -1669 -1551
rect -1625 -1585 -1597 -1551
rect -1557 -1585 -1525 -1551
rect -1489 -1585 -1455 -1551
rect -1419 -1585 -1387 -1551
rect -1347 -1585 -1319 -1551
rect -1275 -1585 -1251 -1551
rect -1203 -1585 -1183 -1551
rect -1131 -1585 -1115 -1551
rect -1059 -1585 -1047 -1551
rect -987 -1585 -979 -1551
rect -915 -1585 -911 -1551
rect -809 -1585 -805 -1551
rect -741 -1585 -733 -1551
rect -673 -1585 -661 -1551
rect -605 -1585 -589 -1551
rect -537 -1585 -517 -1551
rect -469 -1585 -445 -1551
rect -401 -1585 -373 -1551
rect -333 -1585 -301 -1551
rect -265 -1585 -231 -1551
rect -195 -1585 -163 -1551
rect -123 -1585 -95 -1551
rect -51 -1585 -27 -1551
rect 21 -1585 41 -1551
rect 93 -1585 109 -1551
rect 165 -1585 177 -1551
rect 237 -1585 245 -1551
rect 309 -1585 313 -1551
rect 415 -1585 419 -1551
rect 483 -1585 491 -1551
rect 551 -1585 563 -1551
rect 619 -1585 635 -1551
rect 687 -1585 707 -1551
rect 755 -1585 779 -1551
rect 823 -1585 851 -1551
rect 891 -1585 923 -1551
rect 959 -1585 993 -1551
rect 1029 -1585 1061 -1551
rect 1101 -1585 1129 -1551
rect 1173 -1585 1197 -1551
rect 1245 -1585 1265 -1551
rect 1317 -1585 1333 -1551
rect 1389 -1585 1401 -1551
rect 1461 -1585 1469 -1551
rect 1533 -1585 1537 -1551
rect 1639 -1585 1643 -1551
rect 1707 -1585 1715 -1551
rect 1775 -1585 1787 -1551
rect 1843 -1585 1859 -1551
rect 1911 -1585 1931 -1551
rect 1979 -1585 2003 -1551
rect 2047 -1585 2075 -1551
rect 2115 -1585 2147 -1551
rect 2183 -1585 2217 -1551
rect 2253 -1585 2285 -1551
rect 2325 -1585 2353 -1551
rect 2397 -1585 2421 -1551
rect 2469 -1585 2489 -1551
rect 2541 -1585 2557 -1551
rect 2613 -1585 2625 -1551
rect 2685 -1585 2693 -1551
rect 2757 -1585 2761 -1551
rect 2863 -1585 2867 -1551
rect 2931 -1585 2939 -1551
rect 2999 -1585 3011 -1551
rect 3067 -1585 3083 -1551
rect 3135 -1585 3155 -1551
rect 3203 -1585 3227 -1551
rect 3271 -1585 3299 -1551
rect 3339 -1585 3371 -1551
rect 3407 -1585 3441 -1551
rect 3477 -1585 3509 -1551
rect 3549 -1585 3577 -1551
rect 3621 -1585 3645 -1551
rect 3693 -1585 3713 -1551
rect 3765 -1585 3781 -1551
rect 3837 -1585 3849 -1551
rect 3909 -1585 3917 -1551
rect 3981 -1585 3985 -1551
rect 4087 -1585 4091 -1551
rect 4155 -1585 4163 -1551
rect 4223 -1585 4235 -1551
rect 4291 -1585 4307 -1551
rect 4359 -1585 4379 -1551
rect 4427 -1585 4451 -1551
rect 4495 -1585 4523 -1551
rect 4563 -1585 4595 -1551
rect 4631 -1585 4665 -1551
rect 4701 -1585 4733 -1551
rect 4773 -1585 4801 -1551
rect 4845 -1585 4869 -1551
rect 4917 -1585 4937 -1551
rect 4989 -1585 5005 -1551
rect 5061 -1585 5073 -1551
rect 5133 -1585 5141 -1551
rect 5205 -1585 5209 -1551
rect 5311 -1585 5315 -1551
rect 5379 -1585 5387 -1551
rect 5447 -1585 5459 -1551
rect 5515 -1585 5531 -1551
rect 5583 -1585 5603 -1551
rect 5651 -1585 5675 -1551
rect 5719 -1585 5747 -1551
rect 5787 -1585 5819 -1551
rect 5855 -1585 5889 -1551
rect 5925 -1585 5957 -1551
rect 5997 -1585 6025 -1551
rect 6069 -1585 6093 -1551
rect 6141 -1585 6161 -1551
rect 6213 -1585 6229 -1551
rect 6285 -1585 6297 -1551
rect 6357 -1585 6365 -1551
rect 6429 -1585 6433 -1551
rect 6535 -1585 6539 -1551
rect 6603 -1585 6611 -1551
rect 6671 -1585 6683 -1551
rect 6739 -1585 6755 -1551
rect 6789 -1585 6922 -1551
rect -2522 -1618 6922 -1585
rect -2522 -1681 -2422 -1618
rect -2522 -1715 -2489 -1681
rect -2455 -1715 -2422 -1681
rect -2522 -1733 -2422 -1715
rect -2522 -1783 -2489 -1733
rect -2455 -1783 -2422 -1733
rect -2522 -1805 -2422 -1783
rect -2522 -1851 -2489 -1805
rect -2455 -1851 -2422 -1805
rect -2522 -1877 -2422 -1851
rect -2522 -1919 -2489 -1877
rect -2455 -1919 -2422 -1877
rect -2522 -1949 -2422 -1919
rect -2522 -1987 -2489 -1949
rect -2455 -1987 -2422 -1949
rect -2522 -2021 -2422 -1987
rect -2522 -2055 -2489 -2021
rect -2455 -2055 -2422 -2021
rect -2522 -2089 -2422 -2055
rect -2522 -2127 -2489 -2089
rect -2455 -2127 -2422 -2089
rect -2522 -2157 -2422 -2127
rect -2522 -2199 -2489 -2157
rect -2455 -2199 -2422 -2157
rect -2522 -2225 -2422 -2199
rect -2522 -2271 -2489 -2225
rect -2455 -2271 -2422 -2225
rect -2522 -2293 -2422 -2271
rect -2522 -2343 -2489 -2293
rect -2455 -2343 -2422 -2293
rect -2522 -2361 -2422 -2343
rect -2522 -2415 -2489 -2361
rect -2455 -2415 -2422 -2361
rect -2522 -2429 -2422 -2415
rect -2522 -2487 -2489 -2429
rect -2455 -2487 -2422 -2429
rect -2522 -2497 -2422 -2487
rect -2522 -2559 -2489 -2497
rect -2455 -2559 -2422 -2497
rect -2522 -2565 -2422 -2559
rect -2522 -2631 -2489 -2565
rect -2455 -2631 -2422 -2565
rect -2522 -2633 -2422 -2631
rect -2522 -2667 -2489 -2633
rect -2455 -2667 -2422 -2633
rect -2522 -2669 -2422 -2667
rect -2522 -2735 -2489 -2669
rect -2455 -2735 -2422 -2669
rect -2522 -2741 -2422 -2735
rect -2522 -2803 -2489 -2741
rect -2455 -2803 -2422 -2741
rect -2522 -2813 -2422 -2803
rect -2522 -2871 -2489 -2813
rect -2455 -2871 -2422 -2813
rect -2522 -2885 -2422 -2871
rect -2522 -2939 -2489 -2885
rect -2455 -2939 -2422 -2885
rect -2522 -2957 -2422 -2939
rect -2522 -3007 -2489 -2957
rect -2455 -3007 -2422 -2957
rect -2522 -3029 -2422 -3007
rect -2522 -3075 -2489 -3029
rect -2455 -3075 -2422 -3029
rect -2522 -3101 -2422 -3075
rect -2522 -3143 -2489 -3101
rect -2455 -3143 -2422 -3101
rect -2522 -3173 -2422 -3143
rect -2522 -3211 -2489 -3173
rect -2455 -3211 -2422 -3173
rect -2522 -3245 -2422 -3211
rect -2522 -3279 -2489 -3245
rect -2455 -3279 -2422 -3245
rect -2522 -3313 -2422 -3279
rect -2522 -3351 -2489 -3313
rect -2455 -3351 -2422 -3313
rect -2522 -3381 -2422 -3351
rect -2522 -3423 -2489 -3381
rect -2455 -3423 -2422 -3381
rect -2522 -3449 -2422 -3423
rect -2522 -3495 -2489 -3449
rect -2455 -3495 -2422 -3449
rect -2522 -3517 -2422 -3495
rect -2522 -3567 -2489 -3517
rect -2455 -3567 -2422 -3517
rect -2522 -3585 -2422 -3567
rect -2522 -3619 -2489 -3585
rect -2455 -3619 -2422 -3585
rect -2522 -3682 -2422 -3619
rect 6822 -1681 6922 -1618
rect 6822 -1715 6855 -1681
rect 6889 -1715 6922 -1681
rect 6822 -1733 6922 -1715
rect 6822 -1783 6855 -1733
rect 6889 -1783 6922 -1733
rect 6822 -1805 6922 -1783
rect 6822 -1851 6855 -1805
rect 6889 -1851 6922 -1805
rect 6822 -1877 6922 -1851
rect 6822 -1919 6855 -1877
rect 6889 -1919 6922 -1877
rect 6822 -1949 6922 -1919
rect 6822 -1987 6855 -1949
rect 6889 -1987 6922 -1949
rect 6822 -2021 6922 -1987
rect 6822 -2055 6855 -2021
rect 6889 -2055 6922 -2021
rect 6822 -2089 6922 -2055
rect 6822 -2127 6855 -2089
rect 6889 -2127 6922 -2089
rect 6822 -2157 6922 -2127
rect 6822 -2199 6855 -2157
rect 6889 -2199 6922 -2157
rect 6822 -2225 6922 -2199
rect 6822 -2271 6855 -2225
rect 6889 -2271 6922 -2225
rect 6822 -2293 6922 -2271
rect 6822 -2343 6855 -2293
rect 6889 -2343 6922 -2293
rect 6822 -2361 6922 -2343
rect 6822 -2415 6855 -2361
rect 6889 -2415 6922 -2361
rect 6822 -2429 6922 -2415
rect 6822 -2487 6855 -2429
rect 6889 -2487 6922 -2429
rect 6822 -2497 6922 -2487
rect 6822 -2559 6855 -2497
rect 6889 -2559 6922 -2497
rect 6822 -2565 6922 -2559
rect 6822 -2631 6855 -2565
rect 6889 -2631 6922 -2565
rect 6822 -2633 6922 -2631
rect 6822 -2667 6855 -2633
rect 6889 -2667 6922 -2633
rect 6822 -2669 6922 -2667
rect 6822 -2735 6855 -2669
rect 6889 -2735 6922 -2669
rect 6822 -2741 6922 -2735
rect 6822 -2803 6855 -2741
rect 6889 -2803 6922 -2741
rect 6822 -2813 6922 -2803
rect 6822 -2871 6855 -2813
rect 6889 -2871 6922 -2813
rect 6822 -2885 6922 -2871
rect 6822 -2939 6855 -2885
rect 6889 -2939 6922 -2885
rect 6822 -2957 6922 -2939
rect 6822 -3007 6855 -2957
rect 6889 -3007 6922 -2957
rect 6822 -3029 6922 -3007
rect 6822 -3075 6855 -3029
rect 6889 -3075 6922 -3029
rect 6822 -3101 6922 -3075
rect 6822 -3143 6855 -3101
rect 6889 -3143 6922 -3101
rect 6822 -3173 6922 -3143
rect 6822 -3211 6855 -3173
rect 6889 -3211 6922 -3173
rect 6822 -3245 6922 -3211
rect 6822 -3279 6855 -3245
rect 6889 -3279 6922 -3245
rect 6822 -3313 6922 -3279
rect 6822 -3351 6855 -3313
rect 6889 -3351 6922 -3313
rect 6822 -3381 6922 -3351
rect 6822 -3423 6855 -3381
rect 6889 -3423 6922 -3381
rect 6822 -3449 6922 -3423
rect 6822 -3495 6855 -3449
rect 6889 -3495 6922 -3449
rect 6822 -3517 6922 -3495
rect 6822 -3567 6855 -3517
rect 6889 -3567 6922 -3517
rect 6822 -3585 6922 -3567
rect 6822 -3619 6855 -3585
rect 6889 -3619 6922 -3585
rect 6822 -3682 6922 -3619
rect -2522 -3715 6922 -3682
rect -2522 -3749 -2389 -3715
rect -2355 -3749 -2339 -3715
rect -2283 -3749 -2271 -3715
rect -2211 -3749 -2203 -3715
rect -2139 -3749 -2135 -3715
rect -2033 -3749 -2029 -3715
rect -1965 -3749 -1957 -3715
rect -1897 -3749 -1885 -3715
rect -1829 -3749 -1813 -3715
rect -1761 -3749 -1741 -3715
rect -1693 -3749 -1669 -3715
rect -1625 -3749 -1597 -3715
rect -1557 -3749 -1525 -3715
rect -1489 -3749 -1455 -3715
rect -1419 -3749 -1387 -3715
rect -1347 -3749 -1319 -3715
rect -1275 -3749 -1251 -3715
rect -1203 -3749 -1183 -3715
rect -1131 -3749 -1115 -3715
rect -1059 -3749 -1047 -3715
rect -987 -3749 -979 -3715
rect -915 -3749 -911 -3715
rect -809 -3749 -805 -3715
rect -741 -3749 -733 -3715
rect -673 -3749 -661 -3715
rect -605 -3749 -589 -3715
rect -537 -3749 -517 -3715
rect -469 -3749 -445 -3715
rect -401 -3749 -373 -3715
rect -333 -3749 -301 -3715
rect -265 -3749 -231 -3715
rect -195 -3749 -163 -3715
rect -123 -3749 -95 -3715
rect -51 -3749 -27 -3715
rect 21 -3749 41 -3715
rect 93 -3749 109 -3715
rect 165 -3749 177 -3715
rect 237 -3749 245 -3715
rect 309 -3749 313 -3715
rect 415 -3749 419 -3715
rect 483 -3749 491 -3715
rect 551 -3749 563 -3715
rect 619 -3749 635 -3715
rect 687 -3749 707 -3715
rect 755 -3749 779 -3715
rect 823 -3749 851 -3715
rect 891 -3749 923 -3715
rect 959 -3749 993 -3715
rect 1029 -3749 1061 -3715
rect 1101 -3749 1129 -3715
rect 1173 -3749 1197 -3715
rect 1245 -3749 1265 -3715
rect 1317 -3749 1333 -3715
rect 1389 -3749 1401 -3715
rect 1461 -3749 1469 -3715
rect 1533 -3749 1537 -3715
rect 1639 -3749 1643 -3715
rect 1707 -3749 1715 -3715
rect 1775 -3749 1787 -3715
rect 1843 -3749 1859 -3715
rect 1911 -3749 1931 -3715
rect 1979 -3749 2003 -3715
rect 2047 -3749 2075 -3715
rect 2115 -3749 2147 -3715
rect 2183 -3749 2217 -3715
rect 2253 -3749 2285 -3715
rect 2325 -3749 2353 -3715
rect 2397 -3749 2421 -3715
rect 2469 -3749 2489 -3715
rect 2541 -3749 2557 -3715
rect 2613 -3749 2625 -3715
rect 2685 -3749 2693 -3715
rect 2757 -3749 2761 -3715
rect 2863 -3749 2867 -3715
rect 2931 -3749 2939 -3715
rect 2999 -3749 3011 -3715
rect 3067 -3749 3083 -3715
rect 3135 -3749 3155 -3715
rect 3203 -3749 3227 -3715
rect 3271 -3749 3299 -3715
rect 3339 -3749 3371 -3715
rect 3407 -3749 3441 -3715
rect 3477 -3749 3509 -3715
rect 3549 -3749 3577 -3715
rect 3621 -3749 3645 -3715
rect 3693 -3749 3713 -3715
rect 3765 -3749 3781 -3715
rect 3837 -3749 3849 -3715
rect 3909 -3749 3917 -3715
rect 3981 -3749 3985 -3715
rect 4087 -3749 4091 -3715
rect 4155 -3749 4163 -3715
rect 4223 -3749 4235 -3715
rect 4291 -3749 4307 -3715
rect 4359 -3749 4379 -3715
rect 4427 -3749 4451 -3715
rect 4495 -3749 4523 -3715
rect 4563 -3749 4595 -3715
rect 4631 -3749 4665 -3715
rect 4701 -3749 4733 -3715
rect 4773 -3749 4801 -3715
rect 4845 -3749 4869 -3715
rect 4917 -3749 4937 -3715
rect 4989 -3749 5005 -3715
rect 5061 -3749 5073 -3715
rect 5133 -3749 5141 -3715
rect 5205 -3749 5209 -3715
rect 5311 -3749 5315 -3715
rect 5379 -3749 5387 -3715
rect 5447 -3749 5459 -3715
rect 5515 -3749 5531 -3715
rect 5583 -3749 5603 -3715
rect 5651 -3749 5675 -3715
rect 5719 -3749 5747 -3715
rect 5787 -3749 5819 -3715
rect 5855 -3749 5889 -3715
rect 5925 -3749 5957 -3715
rect 5997 -3749 6025 -3715
rect 6069 -3749 6093 -3715
rect 6141 -3749 6161 -3715
rect 6213 -3749 6229 -3715
rect 6285 -3749 6297 -3715
rect 6357 -3749 6365 -3715
rect 6429 -3749 6433 -3715
rect 6535 -3749 6539 -3715
rect 6603 -3749 6611 -3715
rect 6671 -3749 6683 -3715
rect 6739 -3749 6755 -3715
rect 6789 -3749 6922 -3715
rect -2522 -3782 6922 -3749
<< viali >>
rect -2389 2595 -2355 2629
rect -2317 2595 -2305 2629
rect -2305 2595 -2283 2629
rect -2245 2595 -2237 2629
rect -2237 2595 -2211 2629
rect -2173 2595 -2169 2629
rect -2169 2595 -2139 2629
rect -2101 2595 -2067 2629
rect -2029 2595 -1999 2629
rect -1999 2595 -1995 2629
rect -1957 2595 -1931 2629
rect -1931 2595 -1923 2629
rect -1885 2595 -1863 2629
rect -1863 2595 -1851 2629
rect -1813 2595 -1795 2629
rect -1795 2595 -1779 2629
rect -1741 2595 -1727 2629
rect -1727 2595 -1707 2629
rect -1669 2595 -1659 2629
rect -1659 2595 -1635 2629
rect -1597 2595 -1591 2629
rect -1591 2595 -1563 2629
rect -1525 2595 -1523 2629
rect -1523 2595 -1491 2629
rect -1453 2595 -1421 2629
rect -1421 2595 -1419 2629
rect -1381 2595 -1353 2629
rect -1353 2595 -1347 2629
rect -1309 2595 -1285 2629
rect -1285 2595 -1275 2629
rect -1237 2595 -1217 2629
rect -1217 2595 -1203 2629
rect -1165 2595 -1149 2629
rect -1149 2595 -1131 2629
rect -1093 2595 -1081 2629
rect -1081 2595 -1059 2629
rect -1021 2595 -1013 2629
rect -1013 2595 -987 2629
rect -949 2595 -945 2629
rect -945 2595 -915 2629
rect -877 2595 -843 2629
rect -805 2595 -775 2629
rect -775 2595 -771 2629
rect -733 2595 -707 2629
rect -707 2595 -699 2629
rect -661 2595 -639 2629
rect -639 2595 -627 2629
rect -589 2595 -571 2629
rect -571 2595 -555 2629
rect -517 2595 -503 2629
rect -503 2595 -483 2629
rect -445 2595 -435 2629
rect -435 2595 -411 2629
rect -373 2595 -367 2629
rect -367 2595 -339 2629
rect -301 2595 -299 2629
rect -299 2595 -267 2629
rect -229 2595 -197 2629
rect -197 2595 -195 2629
rect -157 2595 -129 2629
rect -129 2595 -123 2629
rect -85 2595 -61 2629
rect -61 2595 -51 2629
rect -13 2595 7 2629
rect 7 2595 21 2629
rect 59 2595 75 2629
rect 75 2595 93 2629
rect 131 2595 143 2629
rect 143 2595 165 2629
rect 203 2595 211 2629
rect 211 2595 237 2629
rect 275 2595 279 2629
rect 279 2595 309 2629
rect 347 2595 381 2629
rect 419 2595 449 2629
rect 449 2595 453 2629
rect 491 2595 517 2629
rect 517 2595 525 2629
rect 563 2595 585 2629
rect 585 2595 597 2629
rect 635 2595 653 2629
rect 653 2595 669 2629
rect 707 2595 721 2629
rect 721 2595 741 2629
rect 779 2595 789 2629
rect 789 2595 813 2629
rect 851 2595 857 2629
rect 857 2595 885 2629
rect 923 2595 925 2629
rect 925 2595 957 2629
rect 995 2595 1027 2629
rect 1027 2595 1029 2629
rect 1067 2595 1095 2629
rect 1095 2595 1101 2629
rect 1139 2595 1163 2629
rect 1163 2595 1173 2629
rect 1211 2595 1231 2629
rect 1231 2595 1245 2629
rect 1283 2595 1299 2629
rect 1299 2595 1317 2629
rect 1355 2595 1367 2629
rect 1367 2595 1389 2629
rect 1427 2595 1435 2629
rect 1435 2595 1461 2629
rect 1499 2595 1503 2629
rect 1503 2595 1533 2629
rect 1571 2595 1605 2629
rect 1643 2595 1673 2629
rect 1673 2595 1677 2629
rect 1715 2595 1741 2629
rect 1741 2595 1749 2629
rect 1787 2595 1809 2629
rect 1809 2595 1821 2629
rect 1859 2595 1877 2629
rect 1877 2595 1893 2629
rect 1931 2595 1945 2629
rect 1945 2595 1965 2629
rect 2003 2595 2013 2629
rect 2013 2595 2037 2629
rect 2075 2595 2081 2629
rect 2081 2595 2109 2629
rect 2147 2595 2149 2629
rect 2149 2595 2181 2629
rect 2219 2595 2251 2629
rect 2251 2595 2253 2629
rect 2291 2595 2319 2629
rect 2319 2595 2325 2629
rect 2363 2595 2387 2629
rect 2387 2595 2397 2629
rect 2435 2595 2455 2629
rect 2455 2595 2469 2629
rect 2507 2595 2523 2629
rect 2523 2595 2541 2629
rect 2579 2595 2591 2629
rect 2591 2595 2613 2629
rect 2651 2595 2659 2629
rect 2659 2595 2685 2629
rect 2723 2595 2727 2629
rect 2727 2595 2757 2629
rect 2795 2595 2829 2629
rect 2867 2595 2897 2629
rect 2897 2595 2901 2629
rect 2939 2595 2965 2629
rect 2965 2595 2973 2629
rect 3011 2595 3033 2629
rect 3033 2595 3045 2629
rect 3083 2595 3101 2629
rect 3101 2595 3117 2629
rect 3155 2595 3169 2629
rect 3169 2595 3189 2629
rect 3227 2595 3237 2629
rect 3237 2595 3261 2629
rect 3299 2595 3305 2629
rect 3305 2595 3333 2629
rect 3371 2595 3373 2629
rect 3373 2595 3405 2629
rect 3443 2595 3475 2629
rect 3475 2595 3477 2629
rect 3515 2595 3543 2629
rect 3543 2595 3549 2629
rect 3587 2595 3611 2629
rect 3611 2595 3621 2629
rect 3659 2595 3679 2629
rect 3679 2595 3693 2629
rect 3731 2595 3747 2629
rect 3747 2595 3765 2629
rect 3803 2595 3815 2629
rect 3815 2595 3837 2629
rect 3875 2595 3883 2629
rect 3883 2595 3909 2629
rect 3947 2595 3951 2629
rect 3951 2595 3981 2629
rect 4019 2595 4053 2629
rect 4091 2595 4121 2629
rect 4121 2595 4125 2629
rect 4163 2595 4189 2629
rect 4189 2595 4197 2629
rect 4235 2595 4257 2629
rect 4257 2595 4269 2629
rect 4307 2595 4325 2629
rect 4325 2595 4341 2629
rect 4379 2595 4393 2629
rect 4393 2595 4413 2629
rect 4451 2595 4461 2629
rect 4461 2595 4485 2629
rect 4523 2595 4529 2629
rect 4529 2595 4557 2629
rect 4595 2595 4597 2629
rect 4597 2595 4629 2629
rect 4667 2595 4699 2629
rect 4699 2595 4701 2629
rect 4739 2595 4767 2629
rect 4767 2595 4773 2629
rect 4811 2595 4835 2629
rect 4835 2595 4845 2629
rect 4883 2595 4903 2629
rect 4903 2595 4917 2629
rect 4955 2595 4971 2629
rect 4971 2595 4989 2629
rect 5027 2595 5039 2629
rect 5039 2595 5061 2629
rect 5099 2595 5107 2629
rect 5107 2595 5133 2629
rect 5171 2595 5175 2629
rect 5175 2595 5205 2629
rect 5243 2595 5277 2629
rect 5315 2595 5345 2629
rect 5345 2595 5349 2629
rect 5387 2595 5413 2629
rect 5413 2595 5421 2629
rect 5459 2595 5481 2629
rect 5481 2595 5493 2629
rect 5531 2595 5549 2629
rect 5549 2595 5565 2629
rect 5603 2595 5617 2629
rect 5617 2595 5637 2629
rect 5675 2595 5685 2629
rect 5685 2595 5709 2629
rect 5747 2595 5753 2629
rect 5753 2595 5781 2629
rect 5819 2595 5821 2629
rect 5821 2595 5853 2629
rect 5891 2595 5923 2629
rect 5923 2595 5925 2629
rect 5963 2595 5991 2629
rect 5991 2595 5997 2629
rect 6035 2595 6059 2629
rect 6059 2595 6069 2629
rect 6107 2595 6127 2629
rect 6127 2595 6141 2629
rect 6179 2595 6195 2629
rect 6195 2595 6213 2629
rect 6251 2595 6263 2629
rect 6263 2595 6285 2629
rect 6323 2595 6331 2629
rect 6331 2595 6357 2629
rect 6395 2595 6399 2629
rect 6399 2595 6429 2629
rect 6467 2595 6501 2629
rect 6539 2595 6569 2629
rect 6569 2595 6573 2629
rect 6611 2595 6637 2629
rect 6637 2595 6645 2629
rect 6683 2595 6705 2629
rect 6705 2595 6717 2629
rect 6755 2595 6789 2629
rect -2489 2411 -2455 2427
rect -2489 2393 -2455 2411
rect -2489 2343 -2455 2355
rect -2489 2321 -2455 2343
rect -2489 2275 -2455 2283
rect -2489 2249 -2455 2275
rect -2489 2207 -2455 2211
rect -2489 2177 -2455 2207
rect -2489 2105 -2455 2139
rect -2489 2037 -2455 2067
rect -2489 2033 -2455 2037
rect -2489 1969 -2455 1995
rect -2489 1961 -2455 1969
rect -2489 1901 -2455 1923
rect -2489 1889 -2455 1901
rect -2489 1833 -2455 1851
rect -2489 1817 -2455 1833
rect -2489 1765 -2455 1779
rect -2489 1745 -2455 1765
rect -2489 1697 -2455 1707
rect -2489 1673 -2455 1697
rect -2489 1629 -2455 1635
rect -2489 1601 -2455 1629
rect -2489 1561 -2455 1563
rect -2489 1529 -2455 1561
rect -2489 1459 -2455 1491
rect -2489 1457 -2455 1459
rect -2489 1391 -2455 1419
rect -2489 1385 -2455 1391
rect -2489 1323 -2455 1347
rect -2489 1313 -2455 1323
rect -2489 1255 -2455 1275
rect -2489 1241 -2455 1255
rect -2489 1187 -2455 1203
rect -2489 1169 -2455 1187
rect -2489 1119 -2455 1131
rect -2489 1097 -2455 1119
rect -2489 1051 -2455 1059
rect -2489 1025 -2455 1051
rect -2489 983 -2455 987
rect -2489 953 -2455 983
rect -2489 881 -2455 915
rect -2489 813 -2455 843
rect -2489 809 -2455 813
rect -2489 745 -2455 771
rect -2489 737 -2455 745
rect -2489 677 -2455 699
rect -2489 665 -2455 677
rect -2489 609 -2455 627
rect -2489 593 -2455 609
rect 6855 2411 6889 2427
rect 6855 2393 6889 2411
rect 6855 2343 6889 2355
rect 6855 2321 6889 2343
rect 6855 2275 6889 2283
rect 6855 2249 6889 2275
rect 6855 2207 6889 2211
rect 6855 2177 6889 2207
rect 6855 2105 6889 2139
rect 6855 2037 6889 2067
rect 6855 2033 6889 2037
rect 6855 1969 6889 1995
rect 6855 1961 6889 1969
rect 6855 1901 6889 1923
rect 6855 1889 6889 1901
rect 6855 1833 6889 1851
rect 6855 1817 6889 1833
rect 6855 1765 6889 1779
rect 6855 1745 6889 1765
rect 6855 1697 6889 1707
rect 6855 1673 6889 1697
rect 6855 1629 6889 1635
rect 6855 1601 6889 1629
rect 6855 1561 6889 1563
rect 6855 1529 6889 1561
rect 6855 1459 6889 1491
rect 6855 1457 6889 1459
rect 6855 1391 6889 1419
rect 6855 1385 6889 1391
rect 6855 1323 6889 1347
rect 6855 1313 6889 1323
rect 6855 1255 6889 1275
rect 6855 1241 6889 1255
rect 6855 1187 6889 1203
rect 6855 1169 6889 1187
rect 6855 1119 6889 1131
rect 6855 1097 6889 1119
rect 6855 1051 6889 1059
rect 6855 1025 6889 1051
rect 6855 983 6889 987
rect 6855 953 6889 983
rect 6855 881 6889 915
rect 6855 813 6889 843
rect 6855 809 6889 813
rect 6855 745 6889 771
rect 6855 737 6889 745
rect 6855 677 6889 699
rect 6855 665 6889 677
rect 6855 609 6889 627
rect 6855 593 6889 609
rect -2389 391 -2355 425
rect -2317 391 -2305 425
rect -2305 391 -2283 425
rect -2245 391 -2237 425
rect -2237 391 -2211 425
rect -2173 391 -2169 425
rect -2169 391 -2139 425
rect -2101 391 -2067 425
rect -2029 391 -1999 425
rect -1999 391 -1995 425
rect -1957 391 -1931 425
rect -1931 391 -1923 425
rect -1885 391 -1863 425
rect -1863 391 -1851 425
rect -1813 391 -1795 425
rect -1795 391 -1779 425
rect -1741 391 -1727 425
rect -1727 391 -1707 425
rect -1669 391 -1659 425
rect -1659 391 -1635 425
rect -1597 391 -1591 425
rect -1591 391 -1563 425
rect -1525 391 -1523 425
rect -1523 391 -1491 425
rect -1453 391 -1421 425
rect -1421 391 -1419 425
rect -1381 391 -1353 425
rect -1353 391 -1347 425
rect -1309 391 -1285 425
rect -1285 391 -1275 425
rect -1237 391 -1217 425
rect -1217 391 -1203 425
rect -1165 391 -1149 425
rect -1149 391 -1131 425
rect -1093 391 -1081 425
rect -1081 391 -1059 425
rect -1021 391 -1013 425
rect -1013 391 -987 425
rect -949 391 -945 425
rect -945 391 -915 425
rect -877 391 -843 425
rect -805 391 -775 425
rect -775 391 -771 425
rect -733 391 -707 425
rect -707 391 -699 425
rect -661 391 -639 425
rect -639 391 -627 425
rect -589 391 -571 425
rect -571 391 -555 425
rect -517 391 -503 425
rect -503 391 -483 425
rect -445 391 -435 425
rect -435 391 -411 425
rect -373 391 -367 425
rect -367 391 -339 425
rect -301 391 -299 425
rect -299 391 -267 425
rect -229 391 -197 425
rect -197 391 -195 425
rect -157 391 -129 425
rect -129 391 -123 425
rect -85 391 -61 425
rect -61 391 -51 425
rect -13 391 7 425
rect 7 391 21 425
rect 59 391 75 425
rect 75 391 93 425
rect 131 391 143 425
rect 143 391 165 425
rect 203 391 211 425
rect 211 391 237 425
rect 275 391 279 425
rect 279 391 309 425
rect 347 391 381 425
rect 419 391 449 425
rect 449 391 453 425
rect 491 391 517 425
rect 517 391 525 425
rect 563 391 585 425
rect 585 391 597 425
rect 635 391 653 425
rect 653 391 669 425
rect 707 391 721 425
rect 721 391 741 425
rect 779 391 789 425
rect 789 391 813 425
rect 851 391 857 425
rect 857 391 885 425
rect 923 391 925 425
rect 925 391 957 425
rect 995 391 1027 425
rect 1027 391 1029 425
rect 1067 391 1095 425
rect 1095 391 1101 425
rect 1139 391 1163 425
rect 1163 391 1173 425
rect 1211 391 1231 425
rect 1231 391 1245 425
rect 1283 391 1299 425
rect 1299 391 1317 425
rect 1355 391 1367 425
rect 1367 391 1389 425
rect 1427 391 1435 425
rect 1435 391 1461 425
rect 1499 391 1503 425
rect 1503 391 1533 425
rect 1571 391 1605 425
rect 1643 391 1673 425
rect 1673 391 1677 425
rect 1715 391 1741 425
rect 1741 391 1749 425
rect 1787 391 1809 425
rect 1809 391 1821 425
rect 1859 391 1877 425
rect 1877 391 1893 425
rect 1931 391 1945 425
rect 1945 391 1965 425
rect 2003 391 2013 425
rect 2013 391 2037 425
rect 2075 391 2081 425
rect 2081 391 2109 425
rect 2147 391 2149 425
rect 2149 391 2181 425
rect 2219 391 2251 425
rect 2251 391 2253 425
rect 2291 391 2319 425
rect 2319 391 2325 425
rect 2363 391 2387 425
rect 2387 391 2397 425
rect 2435 391 2455 425
rect 2455 391 2469 425
rect 2507 391 2523 425
rect 2523 391 2541 425
rect 2579 391 2591 425
rect 2591 391 2613 425
rect 2651 391 2659 425
rect 2659 391 2685 425
rect 2723 391 2727 425
rect 2727 391 2757 425
rect 2795 391 2829 425
rect 2867 391 2897 425
rect 2897 391 2901 425
rect 2939 391 2965 425
rect 2965 391 2973 425
rect 3011 391 3033 425
rect 3033 391 3045 425
rect 3083 391 3101 425
rect 3101 391 3117 425
rect 3155 391 3169 425
rect 3169 391 3189 425
rect 3227 391 3237 425
rect 3237 391 3261 425
rect 3299 391 3305 425
rect 3305 391 3333 425
rect 3371 391 3373 425
rect 3373 391 3405 425
rect 3443 391 3475 425
rect 3475 391 3477 425
rect 3515 391 3543 425
rect 3543 391 3549 425
rect 3587 391 3611 425
rect 3611 391 3621 425
rect 3659 391 3679 425
rect 3679 391 3693 425
rect 3731 391 3747 425
rect 3747 391 3765 425
rect 3803 391 3815 425
rect 3815 391 3837 425
rect 3875 391 3883 425
rect 3883 391 3909 425
rect 3947 391 3951 425
rect 3951 391 3981 425
rect 4019 391 4053 425
rect 4091 391 4121 425
rect 4121 391 4125 425
rect 4163 391 4189 425
rect 4189 391 4197 425
rect 4235 391 4257 425
rect 4257 391 4269 425
rect 4307 391 4325 425
rect 4325 391 4341 425
rect 4379 391 4393 425
rect 4393 391 4413 425
rect 4451 391 4461 425
rect 4461 391 4485 425
rect 4523 391 4529 425
rect 4529 391 4557 425
rect 4595 391 4597 425
rect 4597 391 4629 425
rect 4667 391 4699 425
rect 4699 391 4701 425
rect 4739 391 4767 425
rect 4767 391 4773 425
rect 4811 391 4835 425
rect 4835 391 4845 425
rect 4883 391 4903 425
rect 4903 391 4917 425
rect 4955 391 4971 425
rect 4971 391 4989 425
rect 5027 391 5039 425
rect 5039 391 5061 425
rect 5099 391 5107 425
rect 5107 391 5133 425
rect 5171 391 5175 425
rect 5175 391 5205 425
rect 5243 391 5277 425
rect 5315 391 5345 425
rect 5345 391 5349 425
rect 5387 391 5413 425
rect 5413 391 5421 425
rect 5459 391 5481 425
rect 5481 391 5493 425
rect 5531 391 5549 425
rect 5549 391 5565 425
rect 5603 391 5617 425
rect 5617 391 5637 425
rect 5675 391 5685 425
rect 5685 391 5709 425
rect 5747 391 5753 425
rect 5753 391 5781 425
rect 5819 391 5821 425
rect 5821 391 5853 425
rect 5891 391 5923 425
rect 5923 391 5925 425
rect 5963 391 5991 425
rect 5991 391 5997 425
rect 6035 391 6059 425
rect 6059 391 6069 425
rect 6107 391 6127 425
rect 6127 391 6141 425
rect 6179 391 6195 425
rect 6195 391 6213 425
rect 6251 391 6263 425
rect 6263 391 6285 425
rect 6323 391 6331 425
rect 6331 391 6357 425
rect 6395 391 6399 425
rect 6399 391 6429 425
rect 6467 391 6501 425
rect 6539 391 6569 425
rect 6569 391 6573 425
rect 6611 391 6637 425
rect 6637 391 6645 425
rect 6683 391 6705 425
rect 6705 391 6717 425
rect 6755 391 6789 425
rect 3274 -7 3308 27
rect 3274 -79 3308 -45
rect 3274 -151 3308 -117
rect 3274 -223 3308 -189
rect 3274 -295 3308 -261
rect 3274 -367 3308 -333
rect 3274 -439 3308 -405
rect -1776 -479 -1742 -445
rect 215 -511 249 -477
rect 2677 -487 2711 -453
rect 3274 -511 3308 -477
rect 5051 -8 5085 26
rect 5051 -80 5085 -46
rect 5051 -152 5085 -118
rect 5051 -224 5085 -190
rect 5051 -296 5085 -262
rect 5051 -368 5085 -334
rect 5051 -440 5085 -406
rect 5051 -512 5085 -478
rect 5171 -8 5205 26
rect 5171 -80 5205 -46
rect 5171 -152 5205 -118
rect 5171 -224 5205 -190
rect 5171 -296 5205 -262
rect 5171 -368 5205 -334
rect 5171 -440 5205 -406
rect 5171 -512 5205 -478
rect 6173 -8 6207 26
rect 6173 -80 6207 -46
rect 6173 -152 6207 -118
rect 6173 -224 6207 -190
rect 6173 -296 6207 -262
rect 6173 -368 6207 -334
rect 6173 -440 6207 -406
rect 6173 -512 6207 -478
rect 451 -608 485 -574
rect -2037 -707 -2003 -673
rect -313 -709 -279 -675
rect 125 -705 159 -671
rect 359 -706 393 -672
rect 533 -706 567 -672
rect 771 -705 805 -671
rect 1211 -709 1245 -675
rect 2941 -689 2975 -655
rect 683 -821 717 -787
rect 3276 -903 3310 -869
rect 3276 -975 3310 -941
rect 3276 -1047 3310 -1013
rect 3276 -1119 3310 -1085
rect 3276 -1191 3310 -1157
rect 5052 -904 5086 -870
rect 5052 -976 5086 -942
rect 5052 -1048 5086 -1014
rect 5052 -1120 5086 -1086
rect 5052 -1192 5086 -1158
rect 5172 -904 5206 -870
rect 5172 -976 5206 -942
rect 5172 -1048 5206 -1014
rect 5172 -1120 5206 -1086
rect 5172 -1192 5206 -1158
rect 6174 -903 6208 -869
rect 6174 -975 6208 -941
rect 6174 -1047 6208 -1013
rect 6174 -1119 6208 -1085
rect 6174 -1191 6208 -1157
rect -2389 -1585 -2355 -1551
rect -2317 -1585 -2305 -1551
rect -2305 -1585 -2283 -1551
rect -2245 -1585 -2237 -1551
rect -2237 -1585 -2211 -1551
rect -2173 -1585 -2169 -1551
rect -2169 -1585 -2139 -1551
rect -2101 -1585 -2067 -1551
rect -2029 -1585 -1999 -1551
rect -1999 -1585 -1995 -1551
rect -1957 -1585 -1931 -1551
rect -1931 -1585 -1923 -1551
rect -1885 -1585 -1863 -1551
rect -1863 -1585 -1851 -1551
rect -1813 -1585 -1795 -1551
rect -1795 -1585 -1779 -1551
rect -1741 -1585 -1727 -1551
rect -1727 -1585 -1707 -1551
rect -1669 -1585 -1659 -1551
rect -1659 -1585 -1635 -1551
rect -1597 -1585 -1591 -1551
rect -1591 -1585 -1563 -1551
rect -1525 -1585 -1523 -1551
rect -1523 -1585 -1491 -1551
rect -1453 -1585 -1421 -1551
rect -1421 -1585 -1419 -1551
rect -1381 -1585 -1353 -1551
rect -1353 -1585 -1347 -1551
rect -1309 -1585 -1285 -1551
rect -1285 -1585 -1275 -1551
rect -1237 -1585 -1217 -1551
rect -1217 -1585 -1203 -1551
rect -1165 -1585 -1149 -1551
rect -1149 -1585 -1131 -1551
rect -1093 -1585 -1081 -1551
rect -1081 -1585 -1059 -1551
rect -1021 -1585 -1013 -1551
rect -1013 -1585 -987 -1551
rect -949 -1585 -945 -1551
rect -945 -1585 -915 -1551
rect -877 -1585 -843 -1551
rect -805 -1585 -775 -1551
rect -775 -1585 -771 -1551
rect -733 -1585 -707 -1551
rect -707 -1585 -699 -1551
rect -661 -1585 -639 -1551
rect -639 -1585 -627 -1551
rect -589 -1585 -571 -1551
rect -571 -1585 -555 -1551
rect -517 -1585 -503 -1551
rect -503 -1585 -483 -1551
rect -445 -1585 -435 -1551
rect -435 -1585 -411 -1551
rect -373 -1585 -367 -1551
rect -367 -1585 -339 -1551
rect -301 -1585 -299 -1551
rect -299 -1585 -267 -1551
rect -229 -1585 -197 -1551
rect -197 -1585 -195 -1551
rect -157 -1585 -129 -1551
rect -129 -1585 -123 -1551
rect -85 -1585 -61 -1551
rect -61 -1585 -51 -1551
rect -13 -1585 7 -1551
rect 7 -1585 21 -1551
rect 59 -1585 75 -1551
rect 75 -1585 93 -1551
rect 131 -1585 143 -1551
rect 143 -1585 165 -1551
rect 203 -1585 211 -1551
rect 211 -1585 237 -1551
rect 275 -1585 279 -1551
rect 279 -1585 309 -1551
rect 347 -1585 381 -1551
rect 419 -1585 449 -1551
rect 449 -1585 453 -1551
rect 491 -1585 517 -1551
rect 517 -1585 525 -1551
rect 563 -1585 585 -1551
rect 585 -1585 597 -1551
rect 635 -1585 653 -1551
rect 653 -1585 669 -1551
rect 707 -1585 721 -1551
rect 721 -1585 741 -1551
rect 779 -1585 789 -1551
rect 789 -1585 813 -1551
rect 851 -1585 857 -1551
rect 857 -1585 885 -1551
rect 923 -1585 925 -1551
rect 925 -1585 957 -1551
rect 995 -1585 1027 -1551
rect 1027 -1585 1029 -1551
rect 1067 -1585 1095 -1551
rect 1095 -1585 1101 -1551
rect 1139 -1585 1163 -1551
rect 1163 -1585 1173 -1551
rect 1211 -1585 1231 -1551
rect 1231 -1585 1245 -1551
rect 1283 -1585 1299 -1551
rect 1299 -1585 1317 -1551
rect 1355 -1585 1367 -1551
rect 1367 -1585 1389 -1551
rect 1427 -1585 1435 -1551
rect 1435 -1585 1461 -1551
rect 1499 -1585 1503 -1551
rect 1503 -1585 1533 -1551
rect 1571 -1585 1605 -1551
rect 1643 -1585 1673 -1551
rect 1673 -1585 1677 -1551
rect 1715 -1585 1741 -1551
rect 1741 -1585 1749 -1551
rect 1787 -1585 1809 -1551
rect 1809 -1585 1821 -1551
rect 1859 -1585 1877 -1551
rect 1877 -1585 1893 -1551
rect 1931 -1585 1945 -1551
rect 1945 -1585 1965 -1551
rect 2003 -1585 2013 -1551
rect 2013 -1585 2037 -1551
rect 2075 -1585 2081 -1551
rect 2081 -1585 2109 -1551
rect 2147 -1585 2149 -1551
rect 2149 -1585 2181 -1551
rect 2219 -1585 2251 -1551
rect 2251 -1585 2253 -1551
rect 2291 -1585 2319 -1551
rect 2319 -1585 2325 -1551
rect 2363 -1585 2387 -1551
rect 2387 -1585 2397 -1551
rect 2435 -1585 2455 -1551
rect 2455 -1585 2469 -1551
rect 2507 -1585 2523 -1551
rect 2523 -1585 2541 -1551
rect 2579 -1585 2591 -1551
rect 2591 -1585 2613 -1551
rect 2651 -1585 2659 -1551
rect 2659 -1585 2685 -1551
rect 2723 -1585 2727 -1551
rect 2727 -1585 2757 -1551
rect 2795 -1585 2829 -1551
rect 2867 -1585 2897 -1551
rect 2897 -1585 2901 -1551
rect 2939 -1585 2965 -1551
rect 2965 -1585 2973 -1551
rect 3011 -1585 3033 -1551
rect 3033 -1585 3045 -1551
rect 3083 -1585 3101 -1551
rect 3101 -1585 3117 -1551
rect 3155 -1585 3169 -1551
rect 3169 -1585 3189 -1551
rect 3227 -1585 3237 -1551
rect 3237 -1585 3261 -1551
rect 3299 -1585 3305 -1551
rect 3305 -1585 3333 -1551
rect 3371 -1585 3373 -1551
rect 3373 -1585 3405 -1551
rect 3443 -1585 3475 -1551
rect 3475 -1585 3477 -1551
rect 3515 -1585 3543 -1551
rect 3543 -1585 3549 -1551
rect 3587 -1585 3611 -1551
rect 3611 -1585 3621 -1551
rect 3659 -1585 3679 -1551
rect 3679 -1585 3693 -1551
rect 3731 -1585 3747 -1551
rect 3747 -1585 3765 -1551
rect 3803 -1585 3815 -1551
rect 3815 -1585 3837 -1551
rect 3875 -1585 3883 -1551
rect 3883 -1585 3909 -1551
rect 3947 -1585 3951 -1551
rect 3951 -1585 3981 -1551
rect 4019 -1585 4053 -1551
rect 4091 -1585 4121 -1551
rect 4121 -1585 4125 -1551
rect 4163 -1585 4189 -1551
rect 4189 -1585 4197 -1551
rect 4235 -1585 4257 -1551
rect 4257 -1585 4269 -1551
rect 4307 -1585 4325 -1551
rect 4325 -1585 4341 -1551
rect 4379 -1585 4393 -1551
rect 4393 -1585 4413 -1551
rect 4451 -1585 4461 -1551
rect 4461 -1585 4485 -1551
rect 4523 -1585 4529 -1551
rect 4529 -1585 4557 -1551
rect 4595 -1585 4597 -1551
rect 4597 -1585 4629 -1551
rect 4667 -1585 4699 -1551
rect 4699 -1585 4701 -1551
rect 4739 -1585 4767 -1551
rect 4767 -1585 4773 -1551
rect 4811 -1585 4835 -1551
rect 4835 -1585 4845 -1551
rect 4883 -1585 4903 -1551
rect 4903 -1585 4917 -1551
rect 4955 -1585 4971 -1551
rect 4971 -1585 4989 -1551
rect 5027 -1585 5039 -1551
rect 5039 -1585 5061 -1551
rect 5099 -1585 5107 -1551
rect 5107 -1585 5133 -1551
rect 5171 -1585 5175 -1551
rect 5175 -1585 5205 -1551
rect 5243 -1585 5277 -1551
rect 5315 -1585 5345 -1551
rect 5345 -1585 5349 -1551
rect 5387 -1585 5413 -1551
rect 5413 -1585 5421 -1551
rect 5459 -1585 5481 -1551
rect 5481 -1585 5493 -1551
rect 5531 -1585 5549 -1551
rect 5549 -1585 5565 -1551
rect 5603 -1585 5617 -1551
rect 5617 -1585 5637 -1551
rect 5675 -1585 5685 -1551
rect 5685 -1585 5709 -1551
rect 5747 -1585 5753 -1551
rect 5753 -1585 5781 -1551
rect 5819 -1585 5821 -1551
rect 5821 -1585 5853 -1551
rect 5891 -1585 5923 -1551
rect 5923 -1585 5925 -1551
rect 5963 -1585 5991 -1551
rect 5991 -1585 5997 -1551
rect 6035 -1585 6059 -1551
rect 6059 -1585 6069 -1551
rect 6107 -1585 6127 -1551
rect 6127 -1585 6141 -1551
rect 6179 -1585 6195 -1551
rect 6195 -1585 6213 -1551
rect 6251 -1585 6263 -1551
rect 6263 -1585 6285 -1551
rect 6323 -1585 6331 -1551
rect 6331 -1585 6357 -1551
rect 6395 -1585 6399 -1551
rect 6399 -1585 6429 -1551
rect 6467 -1585 6501 -1551
rect 6539 -1585 6569 -1551
rect 6569 -1585 6573 -1551
rect 6611 -1585 6637 -1551
rect 6637 -1585 6645 -1551
rect 6683 -1585 6705 -1551
rect 6705 -1585 6717 -1551
rect 6755 -1585 6789 -1551
rect -2489 -1749 -2455 -1733
rect -2489 -1767 -2455 -1749
rect -2489 -1817 -2455 -1805
rect -2489 -1839 -2455 -1817
rect -2489 -1885 -2455 -1877
rect -2489 -1911 -2455 -1885
rect -2489 -1953 -2455 -1949
rect -2489 -1983 -2455 -1953
rect -2489 -2055 -2455 -2021
rect -2489 -2123 -2455 -2093
rect -2489 -2127 -2455 -2123
rect -2489 -2191 -2455 -2165
rect -2489 -2199 -2455 -2191
rect -2489 -2259 -2455 -2237
rect -2489 -2271 -2455 -2259
rect -2489 -2327 -2455 -2309
rect -2489 -2343 -2455 -2327
rect -2489 -2395 -2455 -2381
rect -2489 -2415 -2455 -2395
rect -2489 -2463 -2455 -2453
rect -2489 -2487 -2455 -2463
rect -2489 -2531 -2455 -2525
rect -2489 -2559 -2455 -2531
rect -2489 -2599 -2455 -2597
rect -2489 -2631 -2455 -2599
rect -2489 -2701 -2455 -2669
rect -2489 -2703 -2455 -2701
rect -2489 -2769 -2455 -2741
rect -2489 -2775 -2455 -2769
rect -2489 -2837 -2455 -2813
rect -2489 -2847 -2455 -2837
rect -2489 -2905 -2455 -2885
rect -2489 -2919 -2455 -2905
rect -2489 -2973 -2455 -2957
rect -2489 -2991 -2455 -2973
rect -2489 -3041 -2455 -3029
rect -2489 -3063 -2455 -3041
rect -2489 -3109 -2455 -3101
rect -2489 -3135 -2455 -3109
rect -2489 -3177 -2455 -3173
rect -2489 -3207 -2455 -3177
rect -2489 -3279 -2455 -3245
rect -2489 -3347 -2455 -3317
rect -2489 -3351 -2455 -3347
rect -2489 -3415 -2455 -3389
rect -2489 -3423 -2455 -3415
rect -2489 -3483 -2455 -3461
rect -2489 -3495 -2455 -3483
rect -2489 -3551 -2455 -3533
rect -2489 -3567 -2455 -3551
rect 6855 -1749 6889 -1733
rect 6855 -1767 6889 -1749
rect 6855 -1817 6889 -1805
rect 6855 -1839 6889 -1817
rect 6855 -1885 6889 -1877
rect 6855 -1911 6889 -1885
rect 6855 -1953 6889 -1949
rect 6855 -1983 6889 -1953
rect 6855 -2055 6889 -2021
rect 6855 -2123 6889 -2093
rect 6855 -2127 6889 -2123
rect 6855 -2191 6889 -2165
rect 6855 -2199 6889 -2191
rect 6855 -2259 6889 -2237
rect 6855 -2271 6889 -2259
rect 6855 -2327 6889 -2309
rect 6855 -2343 6889 -2327
rect 6855 -2395 6889 -2381
rect 6855 -2415 6889 -2395
rect 6855 -2463 6889 -2453
rect 6855 -2487 6889 -2463
rect 6855 -2531 6889 -2525
rect 6855 -2559 6889 -2531
rect 6855 -2599 6889 -2597
rect 6855 -2631 6889 -2599
rect 6855 -2701 6889 -2669
rect 6855 -2703 6889 -2701
rect 6855 -2769 6889 -2741
rect 6855 -2775 6889 -2769
rect 6855 -2837 6889 -2813
rect 6855 -2847 6889 -2837
rect 6855 -2905 6889 -2885
rect 6855 -2919 6889 -2905
rect 6855 -2973 6889 -2957
rect 6855 -2991 6889 -2973
rect 6855 -3041 6889 -3029
rect 6855 -3063 6889 -3041
rect 6855 -3109 6889 -3101
rect 6855 -3135 6889 -3109
rect 6855 -3177 6889 -3173
rect 6855 -3207 6889 -3177
rect 6855 -3279 6889 -3245
rect 6855 -3347 6889 -3317
rect 6855 -3351 6889 -3347
rect 6855 -3415 6889 -3389
rect 6855 -3423 6889 -3415
rect 6855 -3483 6889 -3461
rect 6855 -3495 6889 -3483
rect 6855 -3551 6889 -3533
rect 6855 -3567 6889 -3551
rect -2389 -3749 -2355 -3715
rect -2317 -3749 -2305 -3715
rect -2305 -3749 -2283 -3715
rect -2245 -3749 -2237 -3715
rect -2237 -3749 -2211 -3715
rect -2173 -3749 -2169 -3715
rect -2169 -3749 -2139 -3715
rect -2101 -3749 -2067 -3715
rect -2029 -3749 -1999 -3715
rect -1999 -3749 -1995 -3715
rect -1957 -3749 -1931 -3715
rect -1931 -3749 -1923 -3715
rect -1885 -3749 -1863 -3715
rect -1863 -3749 -1851 -3715
rect -1813 -3749 -1795 -3715
rect -1795 -3749 -1779 -3715
rect -1741 -3749 -1727 -3715
rect -1727 -3749 -1707 -3715
rect -1669 -3749 -1659 -3715
rect -1659 -3749 -1635 -3715
rect -1597 -3749 -1591 -3715
rect -1591 -3749 -1563 -3715
rect -1525 -3749 -1523 -3715
rect -1523 -3749 -1491 -3715
rect -1453 -3749 -1421 -3715
rect -1421 -3749 -1419 -3715
rect -1381 -3749 -1353 -3715
rect -1353 -3749 -1347 -3715
rect -1309 -3749 -1285 -3715
rect -1285 -3749 -1275 -3715
rect -1237 -3749 -1217 -3715
rect -1217 -3749 -1203 -3715
rect -1165 -3749 -1149 -3715
rect -1149 -3749 -1131 -3715
rect -1093 -3749 -1081 -3715
rect -1081 -3749 -1059 -3715
rect -1021 -3749 -1013 -3715
rect -1013 -3749 -987 -3715
rect -949 -3749 -945 -3715
rect -945 -3749 -915 -3715
rect -877 -3749 -843 -3715
rect -805 -3749 -775 -3715
rect -775 -3749 -771 -3715
rect -733 -3749 -707 -3715
rect -707 -3749 -699 -3715
rect -661 -3749 -639 -3715
rect -639 -3749 -627 -3715
rect -589 -3749 -571 -3715
rect -571 -3749 -555 -3715
rect -517 -3749 -503 -3715
rect -503 -3749 -483 -3715
rect -445 -3749 -435 -3715
rect -435 -3749 -411 -3715
rect -373 -3749 -367 -3715
rect -367 -3749 -339 -3715
rect -301 -3749 -299 -3715
rect -299 -3749 -267 -3715
rect -229 -3749 -197 -3715
rect -197 -3749 -195 -3715
rect -157 -3749 -129 -3715
rect -129 -3749 -123 -3715
rect -85 -3749 -61 -3715
rect -61 -3749 -51 -3715
rect -13 -3749 7 -3715
rect 7 -3749 21 -3715
rect 59 -3749 75 -3715
rect 75 -3749 93 -3715
rect 131 -3749 143 -3715
rect 143 -3749 165 -3715
rect 203 -3749 211 -3715
rect 211 -3749 237 -3715
rect 275 -3749 279 -3715
rect 279 -3749 309 -3715
rect 347 -3749 381 -3715
rect 419 -3749 449 -3715
rect 449 -3749 453 -3715
rect 491 -3749 517 -3715
rect 517 -3749 525 -3715
rect 563 -3749 585 -3715
rect 585 -3749 597 -3715
rect 635 -3749 653 -3715
rect 653 -3749 669 -3715
rect 707 -3749 721 -3715
rect 721 -3749 741 -3715
rect 779 -3749 789 -3715
rect 789 -3749 813 -3715
rect 851 -3749 857 -3715
rect 857 -3749 885 -3715
rect 923 -3749 925 -3715
rect 925 -3749 957 -3715
rect 995 -3749 1027 -3715
rect 1027 -3749 1029 -3715
rect 1067 -3749 1095 -3715
rect 1095 -3749 1101 -3715
rect 1139 -3749 1163 -3715
rect 1163 -3749 1173 -3715
rect 1211 -3749 1231 -3715
rect 1231 -3749 1245 -3715
rect 1283 -3749 1299 -3715
rect 1299 -3749 1317 -3715
rect 1355 -3749 1367 -3715
rect 1367 -3749 1389 -3715
rect 1427 -3749 1435 -3715
rect 1435 -3749 1461 -3715
rect 1499 -3749 1503 -3715
rect 1503 -3749 1533 -3715
rect 1571 -3749 1605 -3715
rect 1643 -3749 1673 -3715
rect 1673 -3749 1677 -3715
rect 1715 -3749 1741 -3715
rect 1741 -3749 1749 -3715
rect 1787 -3749 1809 -3715
rect 1809 -3749 1821 -3715
rect 1859 -3749 1877 -3715
rect 1877 -3749 1893 -3715
rect 1931 -3749 1945 -3715
rect 1945 -3749 1965 -3715
rect 2003 -3749 2013 -3715
rect 2013 -3749 2037 -3715
rect 2075 -3749 2081 -3715
rect 2081 -3749 2109 -3715
rect 2147 -3749 2149 -3715
rect 2149 -3749 2181 -3715
rect 2219 -3749 2251 -3715
rect 2251 -3749 2253 -3715
rect 2291 -3749 2319 -3715
rect 2319 -3749 2325 -3715
rect 2363 -3749 2387 -3715
rect 2387 -3749 2397 -3715
rect 2435 -3749 2455 -3715
rect 2455 -3749 2469 -3715
rect 2507 -3749 2523 -3715
rect 2523 -3749 2541 -3715
rect 2579 -3749 2591 -3715
rect 2591 -3749 2613 -3715
rect 2651 -3749 2659 -3715
rect 2659 -3749 2685 -3715
rect 2723 -3749 2727 -3715
rect 2727 -3749 2757 -3715
rect 2795 -3749 2829 -3715
rect 2867 -3749 2897 -3715
rect 2897 -3749 2901 -3715
rect 2939 -3749 2965 -3715
rect 2965 -3749 2973 -3715
rect 3011 -3749 3033 -3715
rect 3033 -3749 3045 -3715
rect 3083 -3749 3101 -3715
rect 3101 -3749 3117 -3715
rect 3155 -3749 3169 -3715
rect 3169 -3749 3189 -3715
rect 3227 -3749 3237 -3715
rect 3237 -3749 3261 -3715
rect 3299 -3749 3305 -3715
rect 3305 -3749 3333 -3715
rect 3371 -3749 3373 -3715
rect 3373 -3749 3405 -3715
rect 3443 -3749 3475 -3715
rect 3475 -3749 3477 -3715
rect 3515 -3749 3543 -3715
rect 3543 -3749 3549 -3715
rect 3587 -3749 3611 -3715
rect 3611 -3749 3621 -3715
rect 3659 -3749 3679 -3715
rect 3679 -3749 3693 -3715
rect 3731 -3749 3747 -3715
rect 3747 -3749 3765 -3715
rect 3803 -3749 3815 -3715
rect 3815 -3749 3837 -3715
rect 3875 -3749 3883 -3715
rect 3883 -3749 3909 -3715
rect 3947 -3749 3951 -3715
rect 3951 -3749 3981 -3715
rect 4019 -3749 4053 -3715
rect 4091 -3749 4121 -3715
rect 4121 -3749 4125 -3715
rect 4163 -3749 4189 -3715
rect 4189 -3749 4197 -3715
rect 4235 -3749 4257 -3715
rect 4257 -3749 4269 -3715
rect 4307 -3749 4325 -3715
rect 4325 -3749 4341 -3715
rect 4379 -3749 4393 -3715
rect 4393 -3749 4413 -3715
rect 4451 -3749 4461 -3715
rect 4461 -3749 4485 -3715
rect 4523 -3749 4529 -3715
rect 4529 -3749 4557 -3715
rect 4595 -3749 4597 -3715
rect 4597 -3749 4629 -3715
rect 4667 -3749 4699 -3715
rect 4699 -3749 4701 -3715
rect 4739 -3749 4767 -3715
rect 4767 -3749 4773 -3715
rect 4811 -3749 4835 -3715
rect 4835 -3749 4845 -3715
rect 4883 -3749 4903 -3715
rect 4903 -3749 4917 -3715
rect 4955 -3749 4971 -3715
rect 4971 -3749 4989 -3715
rect 5027 -3749 5039 -3715
rect 5039 -3749 5061 -3715
rect 5099 -3749 5107 -3715
rect 5107 -3749 5133 -3715
rect 5171 -3749 5175 -3715
rect 5175 -3749 5205 -3715
rect 5243 -3749 5277 -3715
rect 5315 -3749 5345 -3715
rect 5345 -3749 5349 -3715
rect 5387 -3749 5413 -3715
rect 5413 -3749 5421 -3715
rect 5459 -3749 5481 -3715
rect 5481 -3749 5493 -3715
rect 5531 -3749 5549 -3715
rect 5549 -3749 5565 -3715
rect 5603 -3749 5617 -3715
rect 5617 -3749 5637 -3715
rect 5675 -3749 5685 -3715
rect 5685 -3749 5709 -3715
rect 5747 -3749 5753 -3715
rect 5753 -3749 5781 -3715
rect 5819 -3749 5821 -3715
rect 5821 -3749 5853 -3715
rect 5891 -3749 5923 -3715
rect 5923 -3749 5925 -3715
rect 5963 -3749 5991 -3715
rect 5991 -3749 5997 -3715
rect 6035 -3749 6059 -3715
rect 6059 -3749 6069 -3715
rect 6107 -3749 6127 -3715
rect 6127 -3749 6141 -3715
rect 6179 -3749 6195 -3715
rect 6195 -3749 6213 -3715
rect 6251 -3749 6263 -3715
rect 6263 -3749 6285 -3715
rect 6323 -3749 6331 -3715
rect 6331 -3749 6357 -3715
rect 6395 -3749 6399 -3715
rect 6399 -3749 6429 -3715
rect 6467 -3749 6501 -3715
rect 6539 -3749 6569 -3715
rect 6569 -3749 6573 -3715
rect 6611 -3749 6637 -3715
rect 6637 -3749 6645 -3715
rect 6683 -3749 6705 -3715
rect 6705 -3749 6717 -3715
rect 6755 -3749 6789 -3715
<< metal1 >>
rect -2528 2629 6928 2668
rect -2528 2595 -2389 2629
rect -2355 2595 -2317 2629
rect -2283 2595 -2245 2629
rect -2211 2595 -2173 2629
rect -2139 2595 -2101 2629
rect -2067 2595 -2029 2629
rect -1995 2595 -1957 2629
rect -1923 2595 -1885 2629
rect -1851 2595 -1813 2629
rect -1779 2595 -1741 2629
rect -1707 2595 -1669 2629
rect -1635 2595 -1597 2629
rect -1563 2595 -1525 2629
rect -1491 2595 -1453 2629
rect -1419 2595 -1381 2629
rect -1347 2595 -1309 2629
rect -1275 2595 -1237 2629
rect -1203 2595 -1165 2629
rect -1131 2595 -1093 2629
rect -1059 2595 -1021 2629
rect -987 2595 -949 2629
rect -915 2595 -877 2629
rect -843 2595 -805 2629
rect -771 2595 -733 2629
rect -699 2595 -661 2629
rect -627 2595 -589 2629
rect -555 2595 -517 2629
rect -483 2595 -445 2629
rect -411 2595 -373 2629
rect -339 2595 -301 2629
rect -267 2595 -229 2629
rect -195 2595 -157 2629
rect -123 2595 -85 2629
rect -51 2595 -13 2629
rect 21 2595 59 2629
rect 93 2595 131 2629
rect 165 2595 203 2629
rect 237 2595 275 2629
rect 309 2595 347 2629
rect 381 2595 419 2629
rect 453 2595 491 2629
rect 525 2595 563 2629
rect 597 2595 635 2629
rect 669 2595 707 2629
rect 741 2595 779 2629
rect 813 2595 851 2629
rect 885 2595 923 2629
rect 957 2595 995 2629
rect 1029 2595 1067 2629
rect 1101 2595 1139 2629
rect 1173 2595 1211 2629
rect 1245 2595 1283 2629
rect 1317 2595 1355 2629
rect 1389 2595 1427 2629
rect 1461 2595 1499 2629
rect 1533 2595 1571 2629
rect 1605 2595 1643 2629
rect 1677 2595 1715 2629
rect 1749 2595 1787 2629
rect 1821 2595 1859 2629
rect 1893 2595 1931 2629
rect 1965 2595 2003 2629
rect 2037 2595 2075 2629
rect 2109 2595 2147 2629
rect 2181 2595 2219 2629
rect 2253 2595 2291 2629
rect 2325 2595 2363 2629
rect 2397 2595 2435 2629
rect 2469 2595 2507 2629
rect 2541 2595 2579 2629
rect 2613 2595 2651 2629
rect 2685 2595 2723 2629
rect 2757 2595 2795 2629
rect 2829 2595 2867 2629
rect 2901 2595 2939 2629
rect 2973 2595 3011 2629
rect 3045 2595 3083 2629
rect 3117 2595 3155 2629
rect 3189 2595 3227 2629
rect 3261 2595 3299 2629
rect 3333 2595 3371 2629
rect 3405 2595 3443 2629
rect 3477 2595 3515 2629
rect 3549 2595 3587 2629
rect 3621 2595 3659 2629
rect 3693 2595 3731 2629
rect 3765 2595 3803 2629
rect 3837 2595 3875 2629
rect 3909 2595 3947 2629
rect 3981 2595 4019 2629
rect 4053 2595 4091 2629
rect 4125 2595 4163 2629
rect 4197 2595 4235 2629
rect 4269 2595 4307 2629
rect 4341 2595 4379 2629
rect 4413 2595 4451 2629
rect 4485 2595 4523 2629
rect 4557 2595 4595 2629
rect 4629 2595 4667 2629
rect 4701 2595 4739 2629
rect 4773 2595 4811 2629
rect 4845 2595 4883 2629
rect 4917 2595 4955 2629
rect 4989 2595 5027 2629
rect 5061 2595 5099 2629
rect 5133 2595 5171 2629
rect 5205 2595 5243 2629
rect 5277 2595 5315 2629
rect 5349 2595 5387 2629
rect 5421 2595 5459 2629
rect 5493 2595 5531 2629
rect 5565 2595 5603 2629
rect 5637 2595 5675 2629
rect 5709 2595 5747 2629
rect 5781 2595 5819 2629
rect 5853 2595 5891 2629
rect 5925 2595 5963 2629
rect 5997 2595 6035 2629
rect 6069 2595 6107 2629
rect 6141 2595 6179 2629
rect 6213 2595 6251 2629
rect 6285 2595 6323 2629
rect 6357 2595 6395 2629
rect 6429 2595 6467 2629
rect 6501 2595 6539 2629
rect 6573 2595 6611 2629
rect 6645 2595 6683 2629
rect 6717 2595 6755 2629
rect 6789 2595 6928 2629
rect -2528 2556 6928 2595
rect -2528 2528 -1806 2556
rect -2528 2427 -2398 2528
rect -2528 2393 -2489 2427
rect -2455 2393 -2398 2427
rect -2528 2355 -2398 2393
rect -2528 2321 -2489 2355
rect -2455 2321 -2398 2355
rect -2528 2284 -2398 2321
rect -1834 2284 -1806 2528
rect -2528 2283 -1806 2284
rect -2528 2249 -2489 2283
rect -2455 2256 -1806 2283
rect 6206 2528 6928 2556
rect 6206 2284 6234 2528
rect 6798 2427 6928 2528
rect 6798 2393 6855 2427
rect 6889 2393 6928 2427
rect 6798 2355 6928 2393
rect 6798 2321 6855 2355
rect 6889 2321 6928 2355
rect 6798 2284 6928 2321
rect 6206 2283 6928 2284
rect 6206 2256 6855 2283
rect -2455 2249 -2416 2256
rect -2528 2211 -2416 2249
rect -2528 2177 -2489 2211
rect -2455 2177 -2416 2211
rect -2528 2139 -2416 2177
rect 6816 2249 6855 2256
rect 6889 2249 6928 2283
rect 6816 2211 6928 2249
rect 6816 2177 6855 2211
rect 6889 2177 6928 2211
rect -2528 2105 -2489 2139
rect -2455 2105 -2416 2139
rect -2528 2067 -2416 2105
rect -2528 2033 -2489 2067
rect -2455 2033 -2416 2067
rect -2528 1995 -2416 2033
rect -2528 1961 -2489 1995
rect -2455 1961 -2416 1995
rect -2340 2111 6730 2174
rect -2340 2059 -2278 2111
rect -2226 2059 -2214 2111
rect -2162 2059 -2150 2111
rect -2098 2059 -2086 2111
rect -2034 2059 -2022 2111
rect -1970 2059 -1958 2111
rect -1906 2059 -1894 2111
rect -1842 2059 -1830 2111
rect -1778 2059 -1766 2111
rect -1714 2059 -1702 2111
rect -1650 2059 -1638 2111
rect -1586 2059 -1574 2111
rect -1522 2059 -1510 2111
rect -1458 2059 -1446 2111
rect -1394 2059 -1382 2111
rect -1330 2059 -1318 2111
rect -1266 2059 -1254 2111
rect -1202 2059 -1190 2111
rect -1138 2059 -1126 2111
rect -1074 2059 -1062 2111
rect -1010 2059 -998 2111
rect -946 2059 -934 2111
rect -882 2059 -870 2111
rect -818 2059 -806 2111
rect -754 2059 -742 2111
rect -690 2059 -678 2111
rect -626 2059 -614 2111
rect -562 2059 -550 2111
rect -498 2059 -486 2111
rect -434 2059 -422 2111
rect -370 2059 -358 2111
rect -306 2059 -294 2111
rect -242 2059 -230 2111
rect -178 2059 -166 2111
rect -114 2059 -102 2111
rect -50 2059 -38 2111
rect 14 2059 26 2111
rect 78 2059 90 2111
rect 142 2059 154 2111
rect 206 2059 218 2111
rect 270 2059 282 2111
rect 334 2059 346 2111
rect 398 2059 410 2111
rect 462 2059 474 2111
rect 526 2059 538 2111
rect 590 2059 602 2111
rect 654 2059 666 2111
rect 718 2059 730 2111
rect 782 2059 794 2111
rect 846 2059 858 2111
rect 910 2059 922 2111
rect 974 2059 986 2111
rect 1038 2059 1050 2111
rect 1102 2059 1114 2111
rect 1166 2059 1178 2111
rect 1230 2059 1242 2111
rect 1294 2059 1306 2111
rect 1358 2059 1370 2111
rect 1422 2059 1434 2111
rect 1486 2059 1498 2111
rect 1550 2059 1562 2111
rect 1614 2059 1626 2111
rect 1678 2059 1690 2111
rect 1742 2059 1754 2111
rect 1806 2059 1818 2111
rect 1870 2059 1882 2111
rect 1934 2059 1946 2111
rect 1998 2059 2010 2111
rect 2062 2059 2074 2111
rect 2126 2059 2138 2111
rect 2190 2059 2202 2111
rect 2254 2059 2266 2111
rect 2318 2059 2330 2111
rect 2382 2059 2394 2111
rect 2446 2059 2458 2111
rect 2510 2059 2522 2111
rect 2574 2059 2586 2111
rect 2638 2059 2650 2111
rect 2702 2059 2714 2111
rect 2766 2059 2778 2111
rect 2830 2059 2842 2111
rect 2894 2059 2906 2111
rect 2958 2059 2970 2111
rect 3022 2059 3034 2111
rect 3086 2059 3098 2111
rect 3150 2059 3162 2111
rect 3214 2059 3226 2111
rect 3278 2059 3290 2111
rect 3342 2059 3354 2111
rect 3406 2059 3418 2111
rect 3470 2059 3482 2111
rect 3534 2059 3546 2111
rect 3598 2059 3610 2111
rect 3662 2059 3674 2111
rect 3726 2059 3738 2111
rect 3790 2059 3802 2111
rect 3854 2059 3866 2111
rect 3918 2059 3930 2111
rect 3982 2059 3994 2111
rect 4046 2059 4058 2111
rect 4110 2059 4122 2111
rect 4174 2059 4186 2111
rect 4238 2059 4250 2111
rect 4302 2059 4314 2111
rect 4366 2059 4378 2111
rect 4430 2059 4442 2111
rect 4494 2059 4506 2111
rect 4558 2059 4570 2111
rect 4622 2059 4634 2111
rect 4686 2059 4698 2111
rect 4750 2059 4762 2111
rect 4814 2059 4826 2111
rect 4878 2059 4890 2111
rect 4942 2059 4954 2111
rect 5006 2059 5018 2111
rect 5070 2059 5082 2111
rect 5134 2059 5146 2111
rect 5198 2059 5210 2111
rect 5262 2059 5274 2111
rect 5326 2059 5338 2111
rect 5390 2059 5402 2111
rect 5454 2059 5466 2111
rect 5518 2059 5530 2111
rect 5582 2059 5594 2111
rect 5646 2059 5658 2111
rect 5710 2059 5722 2111
rect 5774 2059 5786 2111
rect 5838 2059 5850 2111
rect 5902 2059 5914 2111
rect 5966 2059 5978 2111
rect 6030 2059 6042 2111
rect 6094 2059 6106 2111
rect 6158 2059 6170 2111
rect 6222 2059 6234 2111
rect 6286 2059 6298 2111
rect 6350 2059 6362 2111
rect 6414 2059 6426 2111
rect 6478 2059 6490 2111
rect 6542 2059 6554 2111
rect 6606 2059 6618 2111
rect 6670 2059 6730 2111
rect -2340 1992 6730 2059
rect 6816 2139 6928 2177
rect 6816 2105 6855 2139
rect 6889 2105 6928 2139
rect 6816 2067 6928 2105
rect 6816 2033 6855 2067
rect 6889 2033 6928 2067
rect 6816 1995 6928 2033
rect -2528 1923 -2416 1961
rect -2528 1889 -2489 1923
rect -2455 1889 -2416 1923
rect -2528 1851 -2416 1889
rect -2528 1817 -2489 1851
rect -2455 1817 -2416 1851
rect -2528 1779 -2416 1817
rect -2528 1745 -2489 1779
rect -2455 1745 -2416 1779
rect -2304 1830 -2232 1834
rect -2304 1778 -2294 1830
rect -2242 1778 -2232 1830
rect -2304 1774 -2232 1778
rect -2146 1806 -2086 1992
rect -1724 1806 -1664 1992
rect -2528 1707 -2416 1745
rect -2528 1673 -2489 1707
rect -2455 1673 -2416 1707
rect -2528 1635 -2416 1673
rect -2528 1601 -2489 1635
rect -2455 1601 -2416 1635
rect -2528 1563 -2416 1601
rect -2528 1529 -2489 1563
rect -2455 1529 -2416 1563
rect -2528 1491 -2416 1529
rect -2528 1457 -2489 1491
rect -2455 1457 -2416 1491
rect -2528 1419 -2416 1457
rect -2528 1385 -2489 1419
rect -2455 1385 -2416 1419
rect -2528 1347 -2416 1385
rect -2528 1313 -2489 1347
rect -2455 1313 -2416 1347
rect -2528 1275 -2416 1313
rect -2528 1241 -2489 1275
rect -2455 1241 -2416 1275
rect -2528 1203 -2416 1241
rect -2528 1169 -2489 1203
rect -2455 1169 -2416 1203
rect -2528 1131 -2416 1169
rect -2528 1097 -2489 1131
rect -2455 1097 -2416 1131
rect -2528 1059 -2416 1097
rect -2528 1025 -2489 1059
rect -2455 1025 -2416 1059
rect -2528 987 -2416 1025
rect -2528 953 -2489 987
rect -2455 953 -2416 987
rect -2528 915 -2416 953
rect -2528 881 -2489 915
rect -2455 881 -2416 915
rect -2528 843 -2416 881
rect -2528 809 -2489 843
rect -2455 809 -2416 843
rect -2528 771 -2416 809
rect -2528 737 -2489 771
rect -2455 737 -2416 771
rect -2528 699 -2416 737
rect -2528 665 -2489 699
rect -2455 665 -2416 699
rect -2528 627 -2416 665
rect -2298 636 -2238 1774
rect -2146 1746 -1664 1806
rect -1296 1830 -1224 1834
rect -1296 1778 -1286 1830
rect -1234 1778 -1224 1830
rect -1296 1774 -1224 1778
rect -432 1828 -372 1992
rect 1286 1828 1346 1992
rect 3002 1832 3062 1992
rect 4716 1832 4776 1992
rect -2146 1228 -2086 1746
rect -1724 1642 -1664 1746
rect -1290 1536 -1230 1774
rect -432 1768 1346 1828
rect 2134 1824 2206 1828
rect 2134 1772 2144 1824
rect 2196 1772 2206 1824
rect 2134 1768 2206 1772
rect 3002 1772 4776 1832
rect -1722 1228 -1662 1348
rect -856 1228 -796 1353
rect -2146 1168 -1662 1228
rect -1296 1224 -1224 1228
rect -1296 1172 -1286 1224
rect -1234 1172 -1224 1224
rect -1296 1168 -1224 1172
rect -862 1224 -790 1228
rect -862 1172 -852 1224
rect -800 1172 -790 1224
rect -862 1168 -790 1172
rect -2146 648 -2086 1168
rect -1722 1042 -1662 1168
rect -1290 942 -1230 1168
rect -856 1042 -796 1168
rect -432 946 -372 1768
rect -6 1228 54 1348
rect 426 1228 486 1470
rect 856 1228 916 1350
rect -12 1224 60 1228
rect -12 1172 -2 1224
rect 50 1172 60 1224
rect -12 1168 60 1172
rect 420 1224 492 1228
rect 420 1172 430 1224
rect 482 1172 492 1224
rect 420 1168 492 1172
rect 850 1224 922 1228
rect 850 1172 860 1224
rect 912 1172 922 1224
rect 850 1168 922 1172
rect -6 1050 54 1168
rect 856 1050 916 1168
rect 1286 930 1346 1768
rect 2140 1530 2200 1768
rect 1712 1228 1772 1348
rect 2564 1228 2624 1350
rect 1706 1224 1778 1228
rect 1706 1172 1716 1224
rect 1768 1172 1778 1224
rect 1706 1168 1778 1172
rect 2138 1224 2210 1228
rect 2138 1172 2148 1224
rect 2200 1172 2210 1224
rect 2138 1168 2210 1172
rect 2558 1224 2630 1228
rect 2558 1172 2568 1224
rect 2620 1172 2630 1224
rect 2558 1168 2630 1172
rect 1712 1044 1772 1168
rect 2144 938 2204 1168
rect 2564 1044 2624 1168
rect 3002 934 3062 1772
rect 3426 1228 3486 1348
rect 3860 1228 3920 1470
rect 4296 1228 4356 1346
rect 3420 1224 3492 1228
rect 3420 1172 3430 1224
rect 3482 1172 3492 1224
rect 3420 1168 3492 1172
rect 3854 1224 3926 1228
rect 3854 1172 3864 1224
rect 3916 1172 3926 1224
rect 3854 1168 3926 1172
rect 4290 1224 4362 1228
rect 4290 1172 4300 1224
rect 4352 1172 4362 1224
rect 4290 1168 4362 1172
rect 3426 1048 3486 1168
rect 4296 1048 4356 1168
rect 4716 940 4776 1772
rect 5568 1824 5640 1828
rect 5568 1772 5578 1824
rect 5630 1772 5640 1824
rect 5568 1768 5640 1772
rect 6000 1820 6060 1992
rect 6432 1820 6492 1992
rect 6816 1961 6855 1995
rect 6889 1961 6928 1995
rect 6816 1923 6928 1961
rect 6816 1889 6855 1923
rect 6889 1889 6928 1923
rect 6816 1851 6928 1889
rect 5574 1554 5634 1768
rect 6000 1760 6492 1820
rect 6588 1824 6660 1828
rect 6588 1772 6598 1824
rect 6650 1772 6660 1824
rect 6588 1768 6660 1772
rect 6816 1817 6855 1851
rect 6889 1817 6928 1851
rect 6816 1779 6928 1817
rect 6000 1644 6060 1760
rect 5136 1228 5196 1348
rect 5130 1224 5202 1228
rect 5130 1172 5140 1224
rect 5192 1172 5202 1224
rect 5130 1168 5202 1172
rect 5570 1224 5642 1228
rect 5570 1172 5580 1224
rect 5632 1172 5642 1224
rect 5570 1168 5642 1172
rect 6000 1226 6060 1350
rect 6432 1226 6492 1760
rect 5136 1048 5196 1168
rect 5576 938 5636 1168
rect 6000 1166 6492 1226
rect 6000 1044 6060 1166
rect -1726 648 -1666 748
rect -2528 593 -2489 627
rect -2455 593 -2416 627
rect -2528 464 -2416 593
rect -2304 632 -2232 636
rect -2304 580 -2294 632
rect -2242 580 -2232 632
rect -2304 576 -2232 580
rect -2146 588 -1666 648
rect 426 636 486 854
rect 3856 636 3916 858
rect 5996 644 6056 750
rect 6432 644 6492 1166
rect -2146 464 -2086 588
rect -1726 464 -1666 588
rect 420 632 492 636
rect 420 580 430 632
rect 482 580 492 632
rect 420 576 492 580
rect 3850 632 3922 636
rect 3850 580 3860 632
rect 3912 580 3922 632
rect 3850 576 3922 580
rect 5996 584 6494 644
rect 6594 636 6654 1768
rect 6816 1745 6855 1779
rect 6889 1745 6928 1779
rect 6816 1707 6928 1745
rect 6816 1673 6855 1707
rect 6889 1673 6928 1707
rect 6816 1635 6928 1673
rect 6816 1601 6855 1635
rect 6889 1601 6928 1635
rect 6816 1563 6928 1601
rect 6816 1529 6855 1563
rect 6889 1529 6928 1563
rect 6816 1491 6928 1529
rect 6816 1457 6855 1491
rect 6889 1457 6928 1491
rect 6816 1419 6928 1457
rect 6816 1385 6855 1419
rect 6889 1385 6928 1419
rect 6816 1347 6928 1385
rect 6816 1313 6855 1347
rect 6889 1313 6928 1347
rect 6816 1275 6928 1313
rect 6816 1241 6855 1275
rect 6889 1241 6928 1275
rect 6816 1203 6928 1241
rect 6816 1169 6855 1203
rect 6889 1169 6928 1203
rect 6816 1131 6928 1169
rect 6816 1097 6855 1131
rect 6889 1097 6928 1131
rect 6816 1059 6928 1097
rect 6816 1025 6855 1059
rect 6889 1025 6928 1059
rect 6816 987 6928 1025
rect 6816 953 6855 987
rect 6889 953 6928 987
rect 6816 915 6928 953
rect 6816 881 6855 915
rect 6889 881 6928 915
rect 6816 843 6928 881
rect 6816 809 6855 843
rect 6889 809 6928 843
rect 6816 771 6928 809
rect 6816 737 6855 771
rect 6889 737 6928 771
rect 6816 699 6928 737
rect 6816 665 6855 699
rect 6889 665 6928 699
rect 6588 632 6660 636
rect 5996 464 6056 584
rect 6432 464 6492 584
rect 6588 580 6598 632
rect 6650 580 6660 632
rect 6588 576 6660 580
rect 6816 627 6928 665
rect 6816 593 6855 627
rect 6889 593 6928 627
rect 6816 464 6928 593
rect -2528 425 6928 464
rect -2528 391 -2389 425
rect -2355 391 -2317 425
rect -2283 391 -2245 425
rect -2211 391 -2173 425
rect -2139 391 -2101 425
rect -2067 391 -2029 425
rect -1995 391 -1957 425
rect -1923 391 -1885 425
rect -1851 391 -1813 425
rect -1779 391 -1741 425
rect -1707 391 -1669 425
rect -1635 391 -1597 425
rect -1563 391 -1525 425
rect -1491 391 -1453 425
rect -1419 391 -1381 425
rect -1347 391 -1309 425
rect -1275 391 -1237 425
rect -1203 391 -1165 425
rect -1131 391 -1093 425
rect -1059 391 -1021 425
rect -987 391 -949 425
rect -915 391 -877 425
rect -843 391 -805 425
rect -771 391 -733 425
rect -699 391 -661 425
rect -627 391 -589 425
rect -555 391 -517 425
rect -483 391 -445 425
rect -411 391 -373 425
rect -339 391 -301 425
rect -267 391 -229 425
rect -195 391 -157 425
rect -123 391 -85 425
rect -51 391 -13 425
rect 21 391 59 425
rect 93 391 131 425
rect 165 391 203 425
rect 237 391 275 425
rect 309 391 347 425
rect 381 391 419 425
rect 453 391 491 425
rect 525 391 563 425
rect 597 391 635 425
rect 669 391 707 425
rect 741 391 779 425
rect 813 391 851 425
rect 885 391 923 425
rect 957 391 995 425
rect 1029 391 1067 425
rect 1101 391 1139 425
rect 1173 391 1211 425
rect 1245 391 1283 425
rect 1317 391 1355 425
rect 1389 391 1427 425
rect 1461 391 1499 425
rect 1533 391 1571 425
rect 1605 391 1643 425
rect 1677 391 1715 425
rect 1749 391 1787 425
rect 1821 391 1859 425
rect 1893 391 1931 425
rect 1965 391 2003 425
rect 2037 391 2075 425
rect 2109 391 2147 425
rect 2181 391 2219 425
rect 2253 391 2291 425
rect 2325 391 2363 425
rect 2397 391 2435 425
rect 2469 391 2507 425
rect 2541 391 2579 425
rect 2613 391 2651 425
rect 2685 391 2723 425
rect 2757 391 2795 425
rect 2829 391 2867 425
rect 2901 391 2939 425
rect 2973 391 3011 425
rect 3045 391 3083 425
rect 3117 391 3155 425
rect 3189 391 3227 425
rect 3261 391 3299 425
rect 3333 391 3371 425
rect 3405 391 3443 425
rect 3477 391 3515 425
rect 3549 391 3587 425
rect 3621 391 3659 425
rect 3693 391 3731 425
rect 3765 391 3803 425
rect 3837 391 3875 425
rect 3909 391 3947 425
rect 3981 391 4019 425
rect 4053 391 4091 425
rect 4125 391 4163 425
rect 4197 391 4235 425
rect 4269 391 4307 425
rect 4341 391 4379 425
rect 4413 391 4451 425
rect 4485 391 4523 425
rect 4557 391 4595 425
rect 4629 391 4667 425
rect 4701 391 4739 425
rect 4773 391 4811 425
rect 4845 391 4883 425
rect 4917 391 4955 425
rect 4989 391 5027 425
rect 5061 391 5099 425
rect 5133 391 5171 425
rect 5205 391 5243 425
rect 5277 391 5315 425
rect 5349 391 5387 425
rect 5421 391 5459 425
rect 5493 391 5531 425
rect 5565 391 5603 425
rect 5637 391 5675 425
rect 5709 391 5747 425
rect 5781 391 5819 425
rect 5853 391 5891 425
rect 5925 391 5963 425
rect 5997 391 6035 425
rect 6069 391 6107 425
rect 6141 391 6179 425
rect 6213 391 6251 425
rect 6285 391 6323 425
rect 6357 391 6395 425
rect 6429 391 6467 425
rect 6501 391 6539 425
rect 6573 391 6611 425
rect 6645 391 6683 425
rect 6717 391 6755 425
rect 6789 391 6928 425
rect -2528 352 6928 391
rect -2066 -428 -1822 352
rect -1794 -445 -1728 -370
rect -1066 -428 -822 352
rect -66 -428 178 352
rect 934 -428 1178 352
rect 1934 -428 2178 352
rect 2660 -424 2724 -376
rect -1794 -479 -1776 -445
rect -1742 -479 -1728 -445
rect 2660 -453 2726 -424
rect 2750 -428 2994 352
rect 3260 156 3324 352
rect 3376 156 3436 352
rect 3510 156 3570 352
rect 3634 156 3694 352
rect 3260 96 3694 156
rect 3260 27 3324 96
rect 3260 -7 3274 27
rect 3308 -7 3324 27
rect 3260 -45 3324 -7
rect 3260 -79 3274 -45
rect 3308 -79 3324 -45
rect 3376 -72 3436 96
rect 3510 10 3570 96
rect 3260 -117 3324 -79
rect 3634 -94 3694 96
rect 4022 156 4082 352
rect 4152 156 4212 352
rect 4280 156 4340 352
rect 4798 164 4858 352
rect 4928 164 4988 352
rect 4022 96 4340 156
rect 4534 154 4606 158
rect 4534 102 4544 154
rect 4596 102 4606 154
rect 4534 98 4606 102
rect 4662 152 4734 156
rect 4662 100 4672 152
rect 4724 100 4734 152
rect 4022 10 4082 96
rect 4152 -84 4212 96
rect 4280 8 4340 96
rect 4540 7 4600 98
rect 4662 96 4734 100
rect 4798 104 4988 164
rect 4668 -96 4728 96
rect 4798 7 4858 104
rect 4928 -107 4988 104
rect 5034 159 5224 352
rect 5274 159 5334 352
rect 5404 159 5464 352
rect 5656 296 5728 300
rect 5656 244 5666 296
rect 5718 244 5728 296
rect 5656 240 5728 244
rect 5034 99 5464 159
rect 5034 26 5224 99
rect 5034 -8 5051 26
rect 5085 -8 5171 26
rect 5205 -8 5224 26
rect 5034 -46 5224 -8
rect 5034 -80 5051 -46
rect 5085 -80 5171 -46
rect 5205 -80 5224 -46
rect 3260 -151 3274 -117
rect 3308 -151 3324 -117
rect 3260 -189 3324 -151
rect 3260 -223 3274 -189
rect 3308 -223 3324 -189
rect 3260 -261 3324 -223
rect 3260 -295 3274 -261
rect 3308 -295 3324 -261
rect 3260 -333 3324 -295
rect 3260 -367 3274 -333
rect 3308 -367 3324 -333
rect 3260 -405 3324 -367
rect 5034 -118 5224 -80
rect 5274 -98 5334 99
rect 5404 2 5464 99
rect 5526 152 5598 156
rect 5526 100 5536 152
rect 5588 100 5598 152
rect 5526 96 5598 100
rect 5532 -92 5592 96
rect 5662 -2 5722 240
rect 5920 164 5980 352
rect 6044 164 6104 352
rect 6158 164 6222 352
rect 5920 104 6222 164
rect 5920 2 5980 104
rect 6044 -84 6104 104
rect 6158 26 6222 104
rect 6158 -8 6173 26
rect 6207 -8 6222 26
rect 6158 -46 6222 -8
rect 6158 -80 6173 -46
rect 6207 -80 6222 -46
rect 5034 -152 5051 -118
rect 5085 -152 5171 -118
rect 5205 -152 5224 -118
rect 5034 -190 5224 -152
rect 5034 -224 5051 -190
rect 5085 -224 5171 -190
rect 5205 -224 5224 -190
rect 5034 -262 5224 -224
rect 5034 -296 5051 -262
rect 5085 -296 5171 -262
rect 5205 -296 5224 -262
rect 5034 -334 5224 -296
rect 5034 -368 5051 -334
rect 5085 -368 5171 -334
rect 5205 -368 5224 -334
rect 202 -464 262 -458
rect -1794 -496 -1728 -479
rect 196 -468 268 -464
rect 196 -520 206 -468
rect 258 -520 268 -468
rect 2660 -487 2677 -453
rect 2711 -487 2726 -453
rect 2660 -502 2726 -487
rect 3260 -439 3274 -405
rect 3308 -439 3324 -405
rect 3260 -477 3324 -439
rect 196 -524 268 -520
rect 3260 -511 3274 -477
rect 3308 -511 3324 -477
rect 202 -530 262 -524
rect 3260 -540 3324 -511
rect -660 -574 1586 -564
rect 3764 -574 3824 -488
rect 3892 -574 3952 -384
rect -660 -608 451 -574
rect 485 -608 1586 -574
rect -660 -624 1586 -608
rect -2292 -673 -1984 -660
rect -2292 -707 -2037 -673
rect -2003 -707 -1984 -673
rect -2292 -720 -1984 -707
rect -660 -768 -600 -624
rect 436 -626 496 -624
rect 348 -662 408 -656
rect 840 -662 900 -656
rect -332 -666 412 -662
rect -332 -671 352 -666
rect -332 -675 125 -671
rect -332 -709 -313 -675
rect -279 -705 125 -675
rect 159 -705 352 -671
rect -279 -709 352 -705
rect -332 -718 352 -709
rect 404 -718 412 -666
rect -332 -722 412 -718
rect 514 -666 1264 -662
rect 514 -671 844 -666
rect 514 -672 771 -671
rect 514 -706 533 -672
rect 567 -705 771 -672
rect 805 -705 844 -671
rect 567 -706 844 -705
rect 514 -718 844 -706
rect 896 -675 1264 -666
rect 896 -709 1211 -675
rect 1245 -709 1264 -675
rect 896 -718 1264 -709
rect 514 -722 1264 -718
rect 348 -728 408 -722
rect 840 -728 900 -722
rect 1526 -766 1586 -624
rect 3632 -634 3952 -574
rect 2922 -655 3104 -642
rect 2922 -689 2941 -655
rect 2975 -689 3104 -655
rect 2922 -702 3104 -689
rect 670 -774 730 -768
rect 664 -778 736 -774
rect 664 -830 674 -778
rect 726 -830 736 -778
rect 664 -834 736 -830
rect 670 -840 730 -834
rect 3262 -869 3326 -840
rect 3262 -903 3276 -869
rect 3310 -903 3326 -869
rect 3262 -941 3326 -903
rect -2066 -1512 -1822 -942
rect -1066 -1512 -822 -942
rect -66 -1512 178 -942
rect 934 -1512 1178 -942
rect 1934 -1512 2178 -942
rect 2752 -1512 2996 -942
rect 3262 -975 3276 -941
rect 3310 -975 3326 -941
rect 3262 -1013 3326 -975
rect 3632 -982 3692 -634
rect 4410 -744 4470 -398
rect 5034 -406 5224 -368
rect 6158 -118 6222 -80
rect 6158 -152 6173 -118
rect 6207 -152 6222 -118
rect 6158 -190 6222 -152
rect 6158 -224 6173 -190
rect 6207 -224 6222 -190
rect 6158 -262 6222 -224
rect 6158 -296 6173 -262
rect 6207 -296 6222 -262
rect 6158 -334 6222 -296
rect 6158 -368 6173 -334
rect 6207 -368 6222 -334
rect 6158 -406 6222 -368
rect 5034 -440 5051 -406
rect 5085 -440 5171 -406
rect 5205 -440 5224 -406
rect 5034 -478 5224 -440
rect 5034 -512 5051 -478
rect 5085 -512 5171 -478
rect 5205 -512 5224 -478
rect 5034 -544 5224 -512
rect 4410 -804 4598 -744
rect 4410 -982 4470 -804
rect 4538 -894 4598 -804
rect 5032 -870 5226 -832
rect 5032 -904 5052 -870
rect 5086 -904 5172 -870
rect 5206 -904 5226 -870
rect 5032 -942 5226 -904
rect 5032 -976 5052 -942
rect 5086 -976 5172 -942
rect 5206 -976 5226 -942
rect 5788 -970 5848 -406
rect 6158 -440 6173 -406
rect 6207 -440 6222 -406
rect 6158 -478 6222 -440
rect 6158 -512 6173 -478
rect 6207 -512 6222 -478
rect 6158 -542 6222 -512
rect 6158 -869 6226 -834
rect 6158 -903 6174 -869
rect 6208 -903 6226 -869
rect 6158 -941 6226 -903
rect 3262 -1047 3276 -1013
rect 3310 -1047 3326 -1013
rect 3262 -1085 3326 -1047
rect 5032 -1014 5226 -976
rect 5032 -1048 5052 -1014
rect 5086 -1048 5172 -1014
rect 5206 -1048 5226 -1014
rect 3262 -1119 3276 -1085
rect 3310 -1119 3326 -1085
rect 3262 -1157 3326 -1119
rect 3262 -1191 3276 -1157
rect 3310 -1191 3326 -1157
rect 3262 -1258 3326 -1191
rect 3376 -1258 3436 -1072
rect 3510 -1258 3570 -1172
rect 3262 -1318 3570 -1258
rect 3262 -1512 3326 -1318
rect 3376 -1512 3436 -1318
rect 3510 -1512 3570 -1318
rect 3754 -1394 3814 -1172
rect 3748 -1398 3820 -1394
rect 3892 -1396 3952 -1086
rect 4022 -1260 4082 -1170
rect 4150 -1260 4210 -1082
rect 4280 -1260 4340 -1172
rect 4022 -1320 4340 -1260
rect 3748 -1450 3758 -1398
rect 3810 -1450 3820 -1398
rect 3748 -1454 3820 -1450
rect 3886 -1400 3958 -1396
rect 3886 -1452 3896 -1400
rect 3948 -1452 3958 -1400
rect 3886 -1456 3958 -1452
rect 4022 -1512 4082 -1320
rect 4150 -1512 4210 -1320
rect 4280 -1512 4340 -1320
rect 4666 -1272 4726 -1080
rect 4794 -1272 4854 -1172
rect 4922 -1272 4982 -1080
rect 5032 -1086 5226 -1048
rect 6158 -975 6174 -941
rect 6208 -975 6226 -941
rect 6158 -1013 6226 -975
rect 6158 -1047 6174 -1013
rect 6208 -1047 6226 -1013
rect 5032 -1120 5052 -1086
rect 5086 -1120 5172 -1086
rect 5206 -1120 5226 -1086
rect 5032 -1158 5226 -1120
rect 5032 -1192 5052 -1158
rect 5086 -1192 5172 -1158
rect 5206 -1192 5226 -1158
rect 5032 -1270 5226 -1192
rect 5274 -1270 5334 -1082
rect 6158 -1085 6226 -1047
rect 5402 -1270 5462 -1166
rect 5530 -1182 5590 -1088
rect 5530 -1248 5592 -1182
rect 5032 -1272 5462 -1270
rect 4666 -1330 5462 -1272
rect 4666 -1332 5226 -1330
rect 5032 -1512 5226 -1332
rect 5532 -1396 5592 -1248
rect 5666 -1274 5726 -1167
rect 5660 -1278 5732 -1274
rect 5660 -1330 5670 -1278
rect 5722 -1330 5732 -1278
rect 5660 -1334 5732 -1330
rect 5916 -1276 5976 -1166
rect 6048 -1276 6108 -1094
rect 6158 -1119 6174 -1085
rect 6208 -1119 6226 -1085
rect 6158 -1157 6226 -1119
rect 6158 -1191 6174 -1157
rect 6208 -1191 6226 -1157
rect 6158 -1276 6226 -1191
rect 5532 -1448 5536 -1396
rect 5588 -1448 5592 -1396
rect 5532 -1458 5592 -1448
rect 5916 -1336 6226 -1276
rect 5916 -1512 5976 -1336
rect 6048 -1512 6108 -1336
rect 6158 -1512 6226 -1336
rect -2528 -1551 6928 -1512
rect -2528 -1585 -2389 -1551
rect -2355 -1585 -2317 -1551
rect -2283 -1585 -2245 -1551
rect -2211 -1585 -2173 -1551
rect -2139 -1585 -2101 -1551
rect -2067 -1585 -2029 -1551
rect -1995 -1585 -1957 -1551
rect -1923 -1585 -1885 -1551
rect -1851 -1585 -1813 -1551
rect -1779 -1585 -1741 -1551
rect -1707 -1585 -1669 -1551
rect -1635 -1585 -1597 -1551
rect -1563 -1585 -1525 -1551
rect -1491 -1585 -1453 -1551
rect -1419 -1585 -1381 -1551
rect -1347 -1585 -1309 -1551
rect -1275 -1585 -1237 -1551
rect -1203 -1585 -1165 -1551
rect -1131 -1585 -1093 -1551
rect -1059 -1585 -1021 -1551
rect -987 -1585 -949 -1551
rect -915 -1585 -877 -1551
rect -843 -1585 -805 -1551
rect -771 -1585 -733 -1551
rect -699 -1585 -661 -1551
rect -627 -1585 -589 -1551
rect -555 -1585 -517 -1551
rect -483 -1585 -445 -1551
rect -411 -1585 -373 -1551
rect -339 -1585 -301 -1551
rect -267 -1585 -229 -1551
rect -195 -1585 -157 -1551
rect -123 -1585 -85 -1551
rect -51 -1585 -13 -1551
rect 21 -1585 59 -1551
rect 93 -1585 131 -1551
rect 165 -1585 203 -1551
rect 237 -1585 275 -1551
rect 309 -1585 347 -1551
rect 381 -1585 419 -1551
rect 453 -1585 491 -1551
rect 525 -1585 563 -1551
rect 597 -1585 635 -1551
rect 669 -1585 707 -1551
rect 741 -1585 779 -1551
rect 813 -1585 851 -1551
rect 885 -1585 923 -1551
rect 957 -1585 995 -1551
rect 1029 -1585 1067 -1551
rect 1101 -1585 1139 -1551
rect 1173 -1585 1211 -1551
rect 1245 -1585 1283 -1551
rect 1317 -1585 1355 -1551
rect 1389 -1585 1427 -1551
rect 1461 -1585 1499 -1551
rect 1533 -1585 1571 -1551
rect 1605 -1585 1643 -1551
rect 1677 -1585 1715 -1551
rect 1749 -1585 1787 -1551
rect 1821 -1585 1859 -1551
rect 1893 -1585 1931 -1551
rect 1965 -1585 2003 -1551
rect 2037 -1585 2075 -1551
rect 2109 -1585 2147 -1551
rect 2181 -1585 2219 -1551
rect 2253 -1585 2291 -1551
rect 2325 -1585 2363 -1551
rect 2397 -1585 2435 -1551
rect 2469 -1585 2507 -1551
rect 2541 -1585 2579 -1551
rect 2613 -1585 2651 -1551
rect 2685 -1585 2723 -1551
rect 2757 -1585 2795 -1551
rect 2829 -1585 2867 -1551
rect 2901 -1585 2939 -1551
rect 2973 -1585 3011 -1551
rect 3045 -1585 3083 -1551
rect 3117 -1585 3155 -1551
rect 3189 -1585 3227 -1551
rect 3261 -1585 3299 -1551
rect 3333 -1585 3371 -1551
rect 3405 -1585 3443 -1551
rect 3477 -1585 3515 -1551
rect 3549 -1585 3587 -1551
rect 3621 -1585 3659 -1551
rect 3693 -1585 3731 -1551
rect 3765 -1585 3803 -1551
rect 3837 -1585 3875 -1551
rect 3909 -1585 3947 -1551
rect 3981 -1585 4019 -1551
rect 4053 -1585 4091 -1551
rect 4125 -1585 4163 -1551
rect 4197 -1585 4235 -1551
rect 4269 -1585 4307 -1551
rect 4341 -1585 4379 -1551
rect 4413 -1585 4451 -1551
rect 4485 -1585 4523 -1551
rect 4557 -1585 4595 -1551
rect 4629 -1585 4667 -1551
rect 4701 -1585 4739 -1551
rect 4773 -1585 4811 -1551
rect 4845 -1585 4883 -1551
rect 4917 -1585 4955 -1551
rect 4989 -1585 5027 -1551
rect 5061 -1585 5099 -1551
rect 5133 -1585 5171 -1551
rect 5205 -1585 5243 -1551
rect 5277 -1585 5315 -1551
rect 5349 -1585 5387 -1551
rect 5421 -1585 5459 -1551
rect 5493 -1585 5531 -1551
rect 5565 -1585 5603 -1551
rect 5637 -1585 5675 -1551
rect 5709 -1585 5747 -1551
rect 5781 -1585 5819 -1551
rect 5853 -1585 5891 -1551
rect 5925 -1585 5963 -1551
rect 5997 -1585 6035 -1551
rect 6069 -1585 6107 -1551
rect 6141 -1585 6179 -1551
rect 6213 -1585 6251 -1551
rect 6285 -1585 6323 -1551
rect 6357 -1585 6395 -1551
rect 6429 -1585 6467 -1551
rect 6501 -1585 6539 -1551
rect 6573 -1585 6611 -1551
rect 6645 -1585 6683 -1551
rect 6717 -1585 6755 -1551
rect 6789 -1585 6928 -1551
rect -2528 -1624 6928 -1585
rect -2528 -1733 -2416 -1624
rect 3892 -1674 3952 -1670
rect 5532 -1674 5592 -1668
rect 3892 -1676 5592 -1674
rect -2528 -1767 -2489 -1733
rect -2455 -1767 -2416 -1733
rect -2528 -1805 -2416 -1767
rect 2526 -1678 5592 -1676
rect 2526 -1680 5536 -1678
rect 2526 -1732 3896 -1680
rect 3948 -1730 5536 -1680
rect 5588 -1730 5592 -1678
rect 3948 -1732 5592 -1730
rect 2526 -1734 5592 -1732
rect 2526 -1736 3952 -1734
rect -2528 -1839 -2489 -1805
rect -2455 -1839 -2416 -1805
rect -2528 -1877 -2416 -1839
rect -2528 -1911 -2489 -1877
rect -2455 -1911 -2416 -1877
rect -2528 -1949 -2416 -1911
rect -2528 -1983 -2489 -1949
rect -2455 -1983 -2416 -1949
rect -2528 -2021 -2416 -1983
rect -2528 -2055 -2489 -2021
rect -2455 -2055 -2416 -2021
rect -2528 -2093 -2416 -2055
rect -2528 -2127 -2489 -2093
rect -2455 -2127 -2416 -2093
rect -2528 -2165 -2416 -2127
rect -2528 -2199 -2489 -2165
rect -2455 -2199 -2416 -2165
rect -2528 -2237 -2416 -2199
rect -2528 -2271 -2489 -2237
rect -2455 -2271 -2416 -2237
rect -2528 -2309 -2416 -2271
rect -2528 -2343 -2489 -2309
rect -2455 -2343 -2416 -2309
rect -2528 -2381 -2416 -2343
rect -2528 -2415 -2489 -2381
rect -2455 -2415 -2416 -2381
rect -2528 -2453 -2416 -2415
rect -2528 -2487 -2489 -2453
rect -2455 -2487 -2416 -2453
rect -2528 -2525 -2416 -2487
rect -2528 -2559 -2489 -2525
rect -2455 -2559 -2416 -2525
rect -2528 -2597 -2416 -2559
rect -2528 -2631 -2489 -2597
rect -2455 -2631 -2416 -2597
rect -2528 -2669 -2416 -2631
rect -2528 -2703 -2489 -2669
rect -2455 -2703 -2416 -2669
rect -2528 -2741 -2416 -2703
rect -2528 -2775 -2489 -2741
rect -2455 -2775 -2416 -2741
rect -2528 -2813 -2416 -2775
rect -2528 -2847 -2489 -2813
rect -2455 -2847 -2416 -2813
rect -2528 -2885 -2416 -2847
rect -2528 -2919 -2489 -2885
rect -2455 -2919 -2416 -2885
rect -2528 -2957 -2416 -2919
rect -2528 -2991 -2489 -2957
rect -2455 -2991 -2416 -2957
rect -2528 -3029 -2416 -2991
rect -2528 -3063 -2489 -3029
rect -2455 -3063 -2416 -3029
rect -2528 -3101 -2416 -3063
rect -1764 -1792 18 -1788
rect -1764 -1844 -44 -1792
rect 8 -1844 18 -1792
rect -1764 -1848 18 -1844
rect 1664 -1792 1736 -1788
rect 1664 -1844 1674 -1792
rect 1726 -1844 1736 -1792
rect 1664 -1848 1736 -1844
rect -1764 -2344 -1704 -1848
rect -1340 -1946 -1280 -1848
rect -48 -2042 12 -1848
rect 1670 -2032 1730 -1848
rect 2526 -2026 2586 -1736
rect 3892 -1742 3952 -1736
rect 5532 -1740 5592 -1734
rect 6816 -1733 6928 -1624
rect 6816 -1767 6855 -1733
rect 6889 -1767 6928 -1733
rect 2944 -1792 3016 -1788
rect 2944 -1844 2954 -1792
rect 3006 -1844 3016 -1792
rect 2944 -1848 3016 -1844
rect 3382 -1792 3454 -1788
rect 3382 -1844 3392 -1792
rect 3444 -1844 3454 -1792
rect 3382 -1848 3454 -1844
rect 5092 -1792 6018 -1788
rect 5092 -1844 5102 -1792
rect 5154 -1844 6018 -1792
rect 5092 -1848 6018 -1844
rect 2950 -1948 3010 -1848
rect 3388 -2036 3448 -1848
rect 5098 -2046 5158 -1848
rect 5518 -1946 5578 -1848
rect -1348 -2344 -1288 -2224
rect -908 -2340 -848 -2124
rect -476 -2340 -416 -2224
rect 378 -2340 438 -2218
rect 810 -2340 870 -2134
rect 1230 -2340 1290 -2218
rect 2094 -2340 2154 -2226
rect 3818 -2340 3878 -2226
rect 4244 -2340 4304 -2122
rect 4666 -2340 4726 -2226
rect 5516 -2336 5576 -2222
rect 5958 -2336 6018 -1848
rect -1764 -2404 -1288 -2344
rect -914 -2344 -842 -2340
rect -914 -2396 -904 -2344
rect -852 -2396 -842 -2344
rect -914 -2400 -842 -2396
rect -482 -2344 -410 -2340
rect -482 -2396 -472 -2344
rect -420 -2396 -410 -2344
rect -482 -2400 -410 -2396
rect -58 -2344 14 -2340
rect -58 -2396 -48 -2344
rect 4 -2396 14 -2344
rect -58 -2400 14 -2396
rect 372 -2344 444 -2340
rect 372 -2396 382 -2344
rect 434 -2396 444 -2344
rect 372 -2400 444 -2396
rect 804 -2344 876 -2340
rect 804 -2396 814 -2344
rect 866 -2396 876 -2344
rect 804 -2400 876 -2396
rect 1224 -2344 1296 -2340
rect 1224 -2396 1234 -2344
rect 1286 -2396 1296 -2344
rect 1224 -2400 1296 -2396
rect 2088 -2344 2160 -2340
rect 2088 -2396 2098 -2344
rect 2150 -2396 2160 -2344
rect 2088 -2400 2160 -2396
rect 2944 -2344 3016 -2340
rect 2944 -2396 2954 -2344
rect 3006 -2396 3016 -2344
rect 2944 -2400 3016 -2396
rect 3378 -2344 3450 -2340
rect 3378 -2396 3388 -2344
rect 3440 -2396 3450 -2344
rect 3378 -2400 3450 -2396
rect 3812 -2344 3884 -2340
rect 3812 -2396 3822 -2344
rect 3874 -2396 3884 -2344
rect 3812 -2400 3884 -2396
rect 4238 -2344 4310 -2340
rect 4238 -2396 4248 -2344
rect 4300 -2396 4310 -2344
rect 4238 -2400 4310 -2396
rect 4660 -2344 4732 -2340
rect 4660 -2396 4670 -2344
rect 4722 -2396 4732 -2344
rect 4660 -2400 4732 -2396
rect 5094 -2344 5166 -2340
rect 5094 -2396 5104 -2344
rect 5156 -2396 5166 -2344
rect 5094 -2400 5166 -2396
rect 5516 -2396 6018 -2336
rect -1764 -2892 -1704 -2404
rect -1348 -2526 -1288 -2404
rect -908 -2406 -848 -2400
rect -476 -2530 -416 -2400
rect -52 -2626 8 -2400
rect 378 -2522 438 -2400
rect 2094 -2526 2154 -2400
rect 2950 -2526 3010 -2400
rect 3384 -2636 3444 -2400
rect 3818 -2530 3878 -2400
rect 4666 -2522 4726 -2400
rect 5100 -2618 5160 -2400
rect 5516 -2526 5576 -2396
rect -1340 -2892 -1280 -2800
rect -906 -2892 -846 -2722
rect -1764 -2952 -846 -2892
rect -1764 -3082 -1704 -2952
rect -1340 -3082 -1280 -2952
rect -906 -3082 -846 -2952
rect 808 -2906 868 -2700
rect 1234 -2906 1294 -2804
rect 1670 -2904 1730 -2696
rect 808 -2966 1294 -2906
rect 1664 -2908 1736 -2904
rect 1664 -2960 1674 -2908
rect 1726 -2960 1736 -2908
rect 1664 -2964 1736 -2960
rect 808 -3082 868 -2966
rect 1234 -3082 1294 -2966
rect 2526 -3082 2586 -2736
rect 4242 -3082 4302 -2700
rect 5516 -2904 5576 -2800
rect 5958 -2904 6018 -2396
rect 5516 -2964 6018 -2904
rect 5516 -3082 5576 -2964
rect 5958 -3082 6018 -2964
rect 6816 -1805 6928 -1767
rect 6816 -1839 6855 -1805
rect 6889 -1839 6928 -1805
rect 6816 -1877 6928 -1839
rect 6816 -1911 6855 -1877
rect 6889 -1911 6928 -1877
rect 6816 -1949 6928 -1911
rect 6816 -1983 6855 -1949
rect 6889 -1983 6928 -1949
rect 6816 -2021 6928 -1983
rect 6816 -2055 6855 -2021
rect 6889 -2055 6928 -2021
rect 6816 -2093 6928 -2055
rect 6816 -2127 6855 -2093
rect 6889 -2127 6928 -2093
rect 6816 -2165 6928 -2127
rect 6816 -2199 6855 -2165
rect 6889 -2199 6928 -2165
rect 6816 -2237 6928 -2199
rect 6816 -2271 6855 -2237
rect 6889 -2271 6928 -2237
rect 6816 -2309 6928 -2271
rect 6816 -2343 6855 -2309
rect 6889 -2343 6928 -2309
rect 6816 -2381 6928 -2343
rect 6816 -2415 6855 -2381
rect 6889 -2415 6928 -2381
rect 6816 -2453 6928 -2415
rect 6816 -2487 6855 -2453
rect 6889 -2487 6928 -2453
rect 6816 -2525 6928 -2487
rect 6816 -2559 6855 -2525
rect 6889 -2559 6928 -2525
rect 6816 -2597 6928 -2559
rect 6816 -2631 6855 -2597
rect 6889 -2631 6928 -2597
rect 6816 -2669 6928 -2631
rect 6816 -2703 6855 -2669
rect 6889 -2703 6928 -2669
rect 6816 -2741 6928 -2703
rect 6816 -2775 6855 -2741
rect 6889 -2775 6928 -2741
rect 6816 -2813 6928 -2775
rect 6816 -2847 6855 -2813
rect 6889 -2847 6928 -2813
rect 6816 -2885 6928 -2847
rect 6816 -2919 6855 -2885
rect 6889 -2919 6928 -2885
rect 6816 -2957 6928 -2919
rect 6816 -2991 6855 -2957
rect 6889 -2991 6928 -2957
rect 6816 -3029 6928 -2991
rect 6816 -3063 6855 -3029
rect 6889 -3063 6928 -3029
rect -2528 -3135 -2489 -3101
rect -2455 -3135 -2416 -3101
rect -2528 -3173 -2416 -3135
rect -2528 -3207 -2489 -3173
rect -2455 -3207 -2416 -3173
rect -2528 -3245 -2416 -3207
rect -2528 -3279 -2489 -3245
rect -2455 -3279 -2416 -3245
rect -2528 -3317 -2416 -3279
rect -1820 -3136 6120 -3082
rect -1820 -3252 -1781 -3136
rect 6079 -3252 6120 -3136
rect -1820 -3296 6120 -3252
rect 6816 -3101 6928 -3063
rect 6816 -3135 6855 -3101
rect 6889 -3135 6928 -3101
rect 6816 -3173 6928 -3135
rect 6816 -3207 6855 -3173
rect 6889 -3207 6928 -3173
rect 6816 -3245 6928 -3207
rect 6816 -3279 6855 -3245
rect 6889 -3279 6928 -3245
rect -2528 -3351 -2489 -3317
rect -2455 -3351 -2416 -3317
rect -2528 -3376 -2416 -3351
rect 6816 -3317 6928 -3279
rect 6816 -3351 6855 -3317
rect 6889 -3351 6928 -3317
rect 6816 -3376 6928 -3351
rect -2528 -3389 -1806 -3376
rect -2528 -3423 -2489 -3389
rect -2455 -3404 -1806 -3389
rect -2455 -3423 -2398 -3404
rect -2528 -3461 -2398 -3423
rect -2528 -3495 -2489 -3461
rect -2455 -3495 -2398 -3461
rect -2528 -3533 -2398 -3495
rect -2528 -3567 -2489 -3533
rect -2455 -3567 -2398 -3533
rect -2528 -3648 -2398 -3567
rect -1834 -3648 -1806 -3404
rect -2528 -3676 -1806 -3648
rect 6206 -3389 6928 -3376
rect 6206 -3404 6855 -3389
rect 6206 -3648 6234 -3404
rect 6798 -3423 6855 -3404
rect 6889 -3423 6928 -3389
rect 6798 -3461 6928 -3423
rect 6798 -3495 6855 -3461
rect 6889 -3495 6928 -3461
rect 6798 -3533 6928 -3495
rect 6798 -3567 6855 -3533
rect 6889 -3567 6928 -3533
rect 6798 -3648 6928 -3567
rect 6206 -3676 6928 -3648
rect -2528 -3715 6928 -3676
rect -2528 -3749 -2389 -3715
rect -2355 -3749 -2317 -3715
rect -2283 -3749 -2245 -3715
rect -2211 -3749 -2173 -3715
rect -2139 -3749 -2101 -3715
rect -2067 -3749 -2029 -3715
rect -1995 -3749 -1957 -3715
rect -1923 -3749 -1885 -3715
rect -1851 -3749 -1813 -3715
rect -1779 -3749 -1741 -3715
rect -1707 -3749 -1669 -3715
rect -1635 -3749 -1597 -3715
rect -1563 -3749 -1525 -3715
rect -1491 -3749 -1453 -3715
rect -1419 -3749 -1381 -3715
rect -1347 -3749 -1309 -3715
rect -1275 -3749 -1237 -3715
rect -1203 -3749 -1165 -3715
rect -1131 -3749 -1093 -3715
rect -1059 -3749 -1021 -3715
rect -987 -3749 -949 -3715
rect -915 -3749 -877 -3715
rect -843 -3749 -805 -3715
rect -771 -3749 -733 -3715
rect -699 -3749 -661 -3715
rect -627 -3749 -589 -3715
rect -555 -3749 -517 -3715
rect -483 -3749 -445 -3715
rect -411 -3749 -373 -3715
rect -339 -3749 -301 -3715
rect -267 -3749 -229 -3715
rect -195 -3749 -157 -3715
rect -123 -3749 -85 -3715
rect -51 -3749 -13 -3715
rect 21 -3749 59 -3715
rect 93 -3749 131 -3715
rect 165 -3749 203 -3715
rect 237 -3749 275 -3715
rect 309 -3749 347 -3715
rect 381 -3749 419 -3715
rect 453 -3749 491 -3715
rect 525 -3749 563 -3715
rect 597 -3749 635 -3715
rect 669 -3749 707 -3715
rect 741 -3749 779 -3715
rect 813 -3749 851 -3715
rect 885 -3749 923 -3715
rect 957 -3749 995 -3715
rect 1029 -3749 1067 -3715
rect 1101 -3749 1139 -3715
rect 1173 -3749 1211 -3715
rect 1245 -3749 1283 -3715
rect 1317 -3749 1355 -3715
rect 1389 -3749 1427 -3715
rect 1461 -3749 1499 -3715
rect 1533 -3749 1571 -3715
rect 1605 -3749 1643 -3715
rect 1677 -3749 1715 -3715
rect 1749 -3749 1787 -3715
rect 1821 -3749 1859 -3715
rect 1893 -3749 1931 -3715
rect 1965 -3749 2003 -3715
rect 2037 -3749 2075 -3715
rect 2109 -3749 2147 -3715
rect 2181 -3749 2219 -3715
rect 2253 -3749 2291 -3715
rect 2325 -3749 2363 -3715
rect 2397 -3749 2435 -3715
rect 2469 -3749 2507 -3715
rect 2541 -3749 2579 -3715
rect 2613 -3749 2651 -3715
rect 2685 -3749 2723 -3715
rect 2757 -3749 2795 -3715
rect 2829 -3749 2867 -3715
rect 2901 -3749 2939 -3715
rect 2973 -3749 3011 -3715
rect 3045 -3749 3083 -3715
rect 3117 -3749 3155 -3715
rect 3189 -3749 3227 -3715
rect 3261 -3749 3299 -3715
rect 3333 -3749 3371 -3715
rect 3405 -3749 3443 -3715
rect 3477 -3749 3515 -3715
rect 3549 -3749 3587 -3715
rect 3621 -3749 3659 -3715
rect 3693 -3749 3731 -3715
rect 3765 -3749 3803 -3715
rect 3837 -3749 3875 -3715
rect 3909 -3749 3947 -3715
rect 3981 -3749 4019 -3715
rect 4053 -3749 4091 -3715
rect 4125 -3749 4163 -3715
rect 4197 -3749 4235 -3715
rect 4269 -3749 4307 -3715
rect 4341 -3749 4379 -3715
rect 4413 -3749 4451 -3715
rect 4485 -3749 4523 -3715
rect 4557 -3749 4595 -3715
rect 4629 -3749 4667 -3715
rect 4701 -3749 4739 -3715
rect 4773 -3749 4811 -3715
rect 4845 -3749 4883 -3715
rect 4917 -3749 4955 -3715
rect 4989 -3749 5027 -3715
rect 5061 -3749 5099 -3715
rect 5133 -3749 5171 -3715
rect 5205 -3749 5243 -3715
rect 5277 -3749 5315 -3715
rect 5349 -3749 5387 -3715
rect 5421 -3749 5459 -3715
rect 5493 -3749 5531 -3715
rect 5565 -3749 5603 -3715
rect 5637 -3749 5675 -3715
rect 5709 -3749 5747 -3715
rect 5781 -3749 5819 -3715
rect 5853 -3749 5891 -3715
rect 5925 -3749 5963 -3715
rect 5997 -3749 6035 -3715
rect 6069 -3749 6107 -3715
rect 6141 -3749 6179 -3715
rect 6213 -3749 6251 -3715
rect 6285 -3749 6323 -3715
rect 6357 -3749 6395 -3715
rect 6429 -3749 6467 -3715
rect 6501 -3749 6539 -3715
rect 6573 -3749 6611 -3715
rect 6645 -3749 6683 -3715
rect 6717 -3749 6755 -3715
rect 6789 -3749 6928 -3715
rect -2528 -3788 6928 -3749
<< via1 >>
rect -2398 2284 -1834 2528
rect 6234 2284 6798 2528
rect -2278 2059 -2226 2111
rect -2214 2059 -2162 2111
rect -2150 2059 -2098 2111
rect -2086 2059 -2034 2111
rect -2022 2059 -1970 2111
rect -1958 2059 -1906 2111
rect -1894 2059 -1842 2111
rect -1830 2059 -1778 2111
rect -1766 2059 -1714 2111
rect -1702 2059 -1650 2111
rect -1638 2059 -1586 2111
rect -1574 2059 -1522 2111
rect -1510 2059 -1458 2111
rect -1446 2059 -1394 2111
rect -1382 2059 -1330 2111
rect -1318 2059 -1266 2111
rect -1254 2059 -1202 2111
rect -1190 2059 -1138 2111
rect -1126 2059 -1074 2111
rect -1062 2059 -1010 2111
rect -998 2059 -946 2111
rect -934 2059 -882 2111
rect -870 2059 -818 2111
rect -806 2059 -754 2111
rect -742 2059 -690 2111
rect -678 2059 -626 2111
rect -614 2059 -562 2111
rect -550 2059 -498 2111
rect -486 2059 -434 2111
rect -422 2059 -370 2111
rect -358 2059 -306 2111
rect -294 2059 -242 2111
rect -230 2059 -178 2111
rect -166 2059 -114 2111
rect -102 2059 -50 2111
rect -38 2059 14 2111
rect 26 2059 78 2111
rect 90 2059 142 2111
rect 154 2059 206 2111
rect 218 2059 270 2111
rect 282 2059 334 2111
rect 346 2059 398 2111
rect 410 2059 462 2111
rect 474 2059 526 2111
rect 538 2059 590 2111
rect 602 2059 654 2111
rect 666 2059 718 2111
rect 730 2059 782 2111
rect 794 2059 846 2111
rect 858 2059 910 2111
rect 922 2059 974 2111
rect 986 2059 1038 2111
rect 1050 2059 1102 2111
rect 1114 2059 1166 2111
rect 1178 2059 1230 2111
rect 1242 2059 1294 2111
rect 1306 2059 1358 2111
rect 1370 2059 1422 2111
rect 1434 2059 1486 2111
rect 1498 2059 1550 2111
rect 1562 2059 1614 2111
rect 1626 2059 1678 2111
rect 1690 2059 1742 2111
rect 1754 2059 1806 2111
rect 1818 2059 1870 2111
rect 1882 2059 1934 2111
rect 1946 2059 1998 2111
rect 2010 2059 2062 2111
rect 2074 2059 2126 2111
rect 2138 2059 2190 2111
rect 2202 2059 2254 2111
rect 2266 2059 2318 2111
rect 2330 2059 2382 2111
rect 2394 2059 2446 2111
rect 2458 2059 2510 2111
rect 2522 2059 2574 2111
rect 2586 2059 2638 2111
rect 2650 2059 2702 2111
rect 2714 2059 2766 2111
rect 2778 2059 2830 2111
rect 2842 2059 2894 2111
rect 2906 2059 2958 2111
rect 2970 2059 3022 2111
rect 3034 2059 3086 2111
rect 3098 2059 3150 2111
rect 3162 2059 3214 2111
rect 3226 2059 3278 2111
rect 3290 2059 3342 2111
rect 3354 2059 3406 2111
rect 3418 2059 3470 2111
rect 3482 2059 3534 2111
rect 3546 2059 3598 2111
rect 3610 2059 3662 2111
rect 3674 2059 3726 2111
rect 3738 2059 3790 2111
rect 3802 2059 3854 2111
rect 3866 2059 3918 2111
rect 3930 2059 3982 2111
rect 3994 2059 4046 2111
rect 4058 2059 4110 2111
rect 4122 2059 4174 2111
rect 4186 2059 4238 2111
rect 4250 2059 4302 2111
rect 4314 2059 4366 2111
rect 4378 2059 4430 2111
rect 4442 2059 4494 2111
rect 4506 2059 4558 2111
rect 4570 2059 4622 2111
rect 4634 2059 4686 2111
rect 4698 2059 4750 2111
rect 4762 2059 4814 2111
rect 4826 2059 4878 2111
rect 4890 2059 4942 2111
rect 4954 2059 5006 2111
rect 5018 2059 5070 2111
rect 5082 2059 5134 2111
rect 5146 2059 5198 2111
rect 5210 2059 5262 2111
rect 5274 2059 5326 2111
rect 5338 2059 5390 2111
rect 5402 2059 5454 2111
rect 5466 2059 5518 2111
rect 5530 2059 5582 2111
rect 5594 2059 5646 2111
rect 5658 2059 5710 2111
rect 5722 2059 5774 2111
rect 5786 2059 5838 2111
rect 5850 2059 5902 2111
rect 5914 2059 5966 2111
rect 5978 2059 6030 2111
rect 6042 2059 6094 2111
rect 6106 2059 6158 2111
rect 6170 2059 6222 2111
rect 6234 2059 6286 2111
rect 6298 2059 6350 2111
rect 6362 2059 6414 2111
rect 6426 2059 6478 2111
rect 6490 2059 6542 2111
rect 6554 2059 6606 2111
rect 6618 2059 6670 2111
rect -2294 1778 -2242 1830
rect -1286 1778 -1234 1830
rect 2144 1772 2196 1824
rect -1286 1172 -1234 1224
rect -852 1172 -800 1224
rect -2 1172 50 1224
rect 430 1172 482 1224
rect 860 1172 912 1224
rect 1716 1172 1768 1224
rect 2148 1172 2200 1224
rect 2568 1172 2620 1224
rect 3430 1172 3482 1224
rect 3864 1172 3916 1224
rect 4300 1172 4352 1224
rect 5578 1772 5630 1824
rect 6598 1772 6650 1824
rect 5140 1172 5192 1224
rect 5580 1172 5632 1224
rect -2294 580 -2242 632
rect 430 580 482 632
rect 3860 580 3912 632
rect 6598 580 6650 632
rect 4544 102 4596 154
rect 4672 100 4724 152
rect 5666 244 5718 296
rect 5536 100 5588 152
rect 206 -477 258 -468
rect 206 -511 215 -477
rect 215 -511 249 -477
rect 249 -511 258 -477
rect 206 -520 258 -511
rect 352 -672 404 -666
rect 352 -706 359 -672
rect 359 -706 393 -672
rect 393 -706 404 -672
rect 352 -718 404 -706
rect 844 -718 896 -666
rect 674 -787 726 -778
rect 674 -821 683 -787
rect 683 -821 717 -787
rect 717 -821 726 -787
rect 674 -830 726 -821
rect 3758 -1450 3810 -1398
rect 3896 -1452 3948 -1400
rect 5670 -1330 5722 -1278
rect 5536 -1448 5588 -1396
rect 3896 -1732 3948 -1680
rect 5536 -1730 5588 -1678
rect -44 -1844 8 -1792
rect 1674 -1844 1726 -1792
rect 2954 -1844 3006 -1792
rect 3392 -1844 3444 -1792
rect 5102 -1844 5154 -1792
rect -904 -2396 -852 -2344
rect -472 -2396 -420 -2344
rect -48 -2396 4 -2344
rect 382 -2396 434 -2344
rect 814 -2396 866 -2344
rect 1234 -2396 1286 -2344
rect 2098 -2396 2150 -2344
rect 2954 -2396 3006 -2344
rect 3388 -2396 3440 -2344
rect 3822 -2396 3874 -2344
rect 4248 -2396 4300 -2344
rect 4670 -2396 4722 -2344
rect 5104 -2396 5156 -2344
rect 1674 -2960 1726 -2908
rect -1781 -3252 6079 -3136
rect -2398 -3648 -1834 -3404
rect 6234 -3648 6798 -3404
<< metal2 >>
rect -2416 2554 -1816 2566
rect -2416 2528 -2384 2554
rect -1848 2528 -1816 2554
rect -2416 2284 -2398 2528
rect -1834 2284 -1816 2528
rect -2416 2258 -2384 2284
rect -1848 2258 -1816 2284
rect -2416 2246 -1816 2258
rect 6216 2554 6816 2566
rect 6216 2528 6248 2554
rect 6784 2528 6816 2554
rect 6216 2284 6234 2528
rect 6798 2284 6816 2528
rect 6216 2258 6248 2284
rect 6784 2258 6816 2284
rect 6216 2246 6816 2258
rect -2340 2113 6730 2174
rect -2340 2111 -2272 2113
rect -2216 2111 -2192 2113
rect -2136 2111 -2112 2113
rect -2056 2111 -2032 2113
rect -1976 2111 -1952 2113
rect -1896 2111 -1872 2113
rect -1816 2111 -1792 2113
rect -1736 2111 -1712 2113
rect -1656 2111 -1632 2113
rect -1576 2111 -1552 2113
rect -1496 2111 -1472 2113
rect -1416 2111 -1392 2113
rect -1336 2111 -1312 2113
rect -1256 2111 -1232 2113
rect -1176 2111 -1152 2113
rect -1096 2111 -1072 2113
rect -1016 2111 -992 2113
rect -936 2111 -912 2113
rect -856 2111 -832 2113
rect -776 2111 -752 2113
rect -696 2111 -672 2113
rect -616 2111 -592 2113
rect -536 2111 -512 2113
rect -456 2111 -432 2113
rect -376 2111 -352 2113
rect -296 2111 -272 2113
rect -216 2111 -192 2113
rect -136 2111 -112 2113
rect -56 2111 -32 2113
rect 24 2111 48 2113
rect 104 2111 128 2113
rect 184 2111 208 2113
rect 264 2111 288 2113
rect 344 2111 368 2113
rect 424 2111 448 2113
rect 504 2111 528 2113
rect 584 2111 608 2113
rect 664 2111 688 2113
rect 744 2111 768 2113
rect 824 2111 848 2113
rect 904 2111 928 2113
rect 984 2111 1008 2113
rect 1064 2111 1088 2113
rect 1144 2111 1168 2113
rect 1224 2111 1248 2113
rect 1304 2111 1328 2113
rect 1384 2111 1408 2113
rect 1464 2111 1488 2113
rect 1544 2111 1568 2113
rect 1624 2111 1648 2113
rect 1704 2111 1728 2113
rect 1784 2111 1808 2113
rect 1864 2111 1888 2113
rect 1944 2111 1968 2113
rect 2024 2111 2048 2113
rect 2104 2111 2128 2113
rect 2184 2111 2208 2113
rect 2264 2111 2288 2113
rect 2344 2111 2368 2113
rect 2424 2111 2448 2113
rect 2504 2111 2528 2113
rect 2584 2111 2608 2113
rect 2664 2111 2688 2113
rect 2744 2111 2768 2113
rect 2824 2111 2848 2113
rect 2904 2111 2928 2113
rect 2984 2111 3008 2113
rect 3064 2111 3088 2113
rect 3144 2111 3168 2113
rect 3224 2111 3248 2113
rect 3304 2111 3328 2113
rect 3384 2111 3408 2113
rect 3464 2111 3488 2113
rect 3544 2111 3568 2113
rect 3624 2111 3648 2113
rect 3704 2111 3728 2113
rect 3784 2111 3808 2113
rect 3864 2111 3888 2113
rect 3944 2111 3968 2113
rect 4024 2111 4048 2113
rect 4104 2111 4128 2113
rect 4184 2111 4208 2113
rect 4264 2111 4288 2113
rect 4344 2111 4368 2113
rect 4424 2111 4448 2113
rect 4504 2111 4528 2113
rect 4584 2111 4608 2113
rect 4664 2111 4688 2113
rect 4744 2111 4768 2113
rect 4824 2111 4848 2113
rect 4904 2111 4928 2113
rect 4984 2111 5008 2113
rect 5064 2111 5088 2113
rect 5144 2111 5168 2113
rect 5224 2111 5248 2113
rect 5304 2111 5328 2113
rect 5384 2111 5408 2113
rect 5464 2111 5488 2113
rect 5544 2111 5568 2113
rect 5624 2111 5648 2113
rect 5704 2111 5728 2113
rect 5784 2111 5808 2113
rect 5864 2111 5888 2113
rect 5944 2111 5968 2113
rect 6024 2111 6048 2113
rect 6104 2111 6128 2113
rect 6184 2111 6208 2113
rect 6264 2111 6288 2113
rect 6344 2111 6368 2113
rect 6424 2111 6448 2113
rect 6504 2111 6528 2113
rect 6584 2111 6608 2113
rect 6664 2111 6730 2113
rect -2340 2059 -2278 2111
rect -2216 2059 -2214 2111
rect -2034 2059 -2032 2111
rect -1970 2059 -1958 2111
rect -1896 2059 -1894 2111
rect -1714 2059 -1712 2111
rect -1650 2059 -1638 2111
rect -1576 2059 -1574 2111
rect -1394 2059 -1392 2111
rect -1330 2059 -1318 2111
rect -1256 2059 -1254 2111
rect -1074 2059 -1072 2111
rect -1010 2059 -998 2111
rect -936 2059 -934 2111
rect -754 2059 -752 2111
rect -690 2059 -678 2111
rect -616 2059 -614 2111
rect -434 2059 -432 2111
rect -370 2059 -358 2111
rect -296 2059 -294 2111
rect -114 2059 -112 2111
rect -50 2059 -38 2111
rect 24 2059 26 2111
rect 206 2059 208 2111
rect 270 2059 282 2111
rect 344 2059 346 2111
rect 526 2059 528 2111
rect 590 2059 602 2111
rect 664 2059 666 2111
rect 846 2059 848 2111
rect 910 2059 922 2111
rect 984 2059 986 2111
rect 1166 2059 1168 2111
rect 1230 2059 1242 2111
rect 1304 2059 1306 2111
rect 1486 2059 1488 2111
rect 1550 2059 1562 2111
rect 1624 2059 1626 2111
rect 1806 2059 1808 2111
rect 1870 2059 1882 2111
rect 1944 2059 1946 2111
rect 2126 2059 2128 2111
rect 2190 2059 2202 2111
rect 2264 2059 2266 2111
rect 2446 2059 2448 2111
rect 2510 2059 2522 2111
rect 2584 2059 2586 2111
rect 2766 2059 2768 2111
rect 2830 2059 2842 2111
rect 2904 2059 2906 2111
rect 3086 2059 3088 2111
rect 3150 2059 3162 2111
rect 3224 2059 3226 2111
rect 3406 2059 3408 2111
rect 3470 2059 3482 2111
rect 3544 2059 3546 2111
rect 3726 2059 3728 2111
rect 3790 2059 3802 2111
rect 3864 2059 3866 2111
rect 4046 2059 4048 2111
rect 4110 2059 4122 2111
rect 4184 2059 4186 2111
rect 4366 2059 4368 2111
rect 4430 2059 4442 2111
rect 4504 2059 4506 2111
rect 4686 2059 4688 2111
rect 4750 2059 4762 2111
rect 4824 2059 4826 2111
rect 5006 2059 5008 2111
rect 5070 2059 5082 2111
rect 5144 2059 5146 2111
rect 5326 2059 5328 2111
rect 5390 2059 5402 2111
rect 5464 2059 5466 2111
rect 5646 2059 5648 2111
rect 5710 2059 5722 2111
rect 5784 2059 5786 2111
rect 5966 2059 5968 2111
rect 6030 2059 6042 2111
rect 6104 2059 6106 2111
rect 6286 2059 6288 2111
rect 6350 2059 6362 2111
rect 6424 2059 6426 2111
rect 6606 2059 6608 2111
rect 6670 2059 6730 2111
rect -2340 2057 -2272 2059
rect -2216 2057 -2192 2059
rect -2136 2057 -2112 2059
rect -2056 2057 -2032 2059
rect -1976 2057 -1952 2059
rect -1896 2057 -1872 2059
rect -1816 2057 -1792 2059
rect -1736 2057 -1712 2059
rect -1656 2057 -1632 2059
rect -1576 2057 -1552 2059
rect -1496 2057 -1472 2059
rect -1416 2057 -1392 2059
rect -1336 2057 -1312 2059
rect -1256 2057 -1232 2059
rect -1176 2057 -1152 2059
rect -1096 2057 -1072 2059
rect -1016 2057 -992 2059
rect -936 2057 -912 2059
rect -856 2057 -832 2059
rect -776 2057 -752 2059
rect -696 2057 -672 2059
rect -616 2057 -592 2059
rect -536 2057 -512 2059
rect -456 2057 -432 2059
rect -376 2057 -352 2059
rect -296 2057 -272 2059
rect -216 2057 -192 2059
rect -136 2057 -112 2059
rect -56 2057 -32 2059
rect 24 2057 48 2059
rect 104 2057 128 2059
rect 184 2057 208 2059
rect 264 2057 288 2059
rect 344 2057 368 2059
rect 424 2057 448 2059
rect 504 2057 528 2059
rect 584 2057 608 2059
rect 664 2057 688 2059
rect 744 2057 768 2059
rect 824 2057 848 2059
rect 904 2057 928 2059
rect 984 2057 1008 2059
rect 1064 2057 1088 2059
rect 1144 2057 1168 2059
rect 1224 2057 1248 2059
rect 1304 2057 1328 2059
rect 1384 2057 1408 2059
rect 1464 2057 1488 2059
rect 1544 2057 1568 2059
rect 1624 2057 1648 2059
rect 1704 2057 1728 2059
rect 1784 2057 1808 2059
rect 1864 2057 1888 2059
rect 1944 2057 1968 2059
rect 2024 2057 2048 2059
rect 2104 2057 2128 2059
rect 2184 2057 2208 2059
rect 2264 2057 2288 2059
rect 2344 2057 2368 2059
rect 2424 2057 2448 2059
rect 2504 2057 2528 2059
rect 2584 2057 2608 2059
rect 2664 2057 2688 2059
rect 2744 2057 2768 2059
rect 2824 2057 2848 2059
rect 2904 2057 2928 2059
rect 2984 2057 3008 2059
rect 3064 2057 3088 2059
rect 3144 2057 3168 2059
rect 3224 2057 3248 2059
rect 3304 2057 3328 2059
rect 3384 2057 3408 2059
rect 3464 2057 3488 2059
rect 3544 2057 3568 2059
rect 3624 2057 3648 2059
rect 3704 2057 3728 2059
rect 3784 2057 3808 2059
rect 3864 2057 3888 2059
rect 3944 2057 3968 2059
rect 4024 2057 4048 2059
rect 4104 2057 4128 2059
rect 4184 2057 4208 2059
rect 4264 2057 4288 2059
rect 4344 2057 4368 2059
rect 4424 2057 4448 2059
rect 4504 2057 4528 2059
rect 4584 2057 4608 2059
rect 4664 2057 4688 2059
rect 4744 2057 4768 2059
rect 4824 2057 4848 2059
rect 4904 2057 4928 2059
rect 4984 2057 5008 2059
rect 5064 2057 5088 2059
rect 5144 2057 5168 2059
rect 5224 2057 5248 2059
rect 5304 2057 5328 2059
rect 5384 2057 5408 2059
rect 5464 2057 5488 2059
rect 5544 2057 5568 2059
rect 5624 2057 5648 2059
rect 5704 2057 5728 2059
rect 5784 2057 5808 2059
rect 5864 2057 5888 2059
rect 5944 2057 5968 2059
rect 6024 2057 6048 2059
rect 6104 2057 6128 2059
rect 6184 2057 6208 2059
rect 6264 2057 6288 2059
rect 6344 2057 6368 2059
rect 6424 2057 6448 2059
rect 6504 2057 6528 2059
rect 6584 2057 6608 2059
rect 6664 2057 6730 2059
rect -2340 1992 6730 2057
rect -2298 1834 -2238 1840
rect -1290 1834 -1230 1840
rect -2298 1830 -1230 1834
rect -2298 1778 -2294 1830
rect -2242 1778 -1286 1830
rect -1234 1778 -1230 1830
rect -2298 1774 -1230 1778
rect -2298 1768 -2238 1774
rect -1290 1768 -1230 1774
rect 2140 1828 2200 1834
rect 5574 1828 5634 1834
rect 6594 1828 6654 1834
rect 2140 1824 6654 1828
rect 2140 1772 2144 1824
rect 2196 1772 5578 1824
rect 5630 1772 6598 1824
rect 6650 1772 6654 1824
rect 2140 1768 6654 1772
rect 2140 1762 2200 1768
rect 5574 1762 5634 1768
rect 6594 1762 6654 1768
rect -1290 1228 -1230 1234
rect -856 1228 -796 1234
rect -6 1228 54 1234
rect 426 1228 486 1234
rect 856 1228 916 1234
rect 1712 1228 1772 1234
rect 2144 1228 2204 1234
rect 2564 1228 2624 1234
rect 3426 1228 3486 1234
rect 3860 1228 3920 1234
rect 4296 1228 4356 1234
rect 5136 1228 5196 1234
rect 5576 1228 5636 1234
rect -1290 1224 6776 1228
rect -1290 1172 -1286 1224
rect -1234 1172 -852 1224
rect -800 1172 -2 1224
rect 50 1172 430 1224
rect 482 1172 860 1224
rect 912 1172 1716 1224
rect 1768 1172 2148 1224
rect 2200 1172 2568 1224
rect 2620 1172 3430 1224
rect 3482 1172 3864 1224
rect 3916 1172 4300 1224
rect 4352 1172 5140 1224
rect 5192 1172 5580 1224
rect 5632 1172 6776 1224
rect -1290 1168 6776 1172
rect -1290 1162 -1230 1168
rect -856 1162 -796 1168
rect -6 1162 54 1168
rect 426 1162 486 1168
rect 856 1162 916 1168
rect 1712 1162 1772 1168
rect 2144 1162 2204 1168
rect 2564 1162 2624 1168
rect 3426 1162 3486 1168
rect 3860 1162 3920 1168
rect 4296 1162 4356 1168
rect 5136 1162 5196 1168
rect 5576 1162 5636 1168
rect -2298 636 -2238 642
rect 426 636 486 642
rect 3856 636 3916 642
rect 6594 636 6654 642
rect -2298 632 6654 636
rect -2298 580 -2294 632
rect -2242 580 430 632
rect 482 580 3860 632
rect 3912 580 6598 632
rect 6650 580 6654 632
rect -2298 576 6654 580
rect -2298 570 -2238 576
rect 426 570 486 576
rect 3856 570 3916 576
rect 5662 300 5722 306
rect 202 296 5722 300
rect 202 244 5666 296
rect 5718 244 5722 296
rect 202 240 5722 244
rect 202 -464 262 240
rect 5662 234 5722 240
rect 4540 158 4600 164
rect 348 154 4600 158
rect 348 102 4544 154
rect 4596 102 4600 154
rect 348 98 4600 102
rect 196 -468 268 -464
rect 196 -520 206 -468
rect 258 -520 268 -468
rect 196 -524 268 -520
rect 348 -662 408 98
rect 4540 92 4600 98
rect 4668 156 4728 162
rect 5532 156 5592 162
rect 5802 156 5862 576
rect 6594 570 6654 576
rect 4668 152 5862 156
rect 4668 100 4672 152
rect 4724 100 5536 152
rect 5588 100 5862 152
rect 4668 96 5862 100
rect 4668 90 4728 96
rect 5532 90 5592 96
rect 6716 32 6776 1168
rect 6378 -28 6776 32
rect 342 -666 414 -662
rect 342 -718 352 -666
rect 404 -718 414 -666
rect 342 -722 414 -718
rect 834 -666 906 -662
rect 834 -718 844 -666
rect 896 -718 906 -666
rect 834 -722 906 -718
rect 664 -778 736 -774
rect 664 -830 674 -778
rect 726 -830 736 -778
rect 664 -834 736 -830
rect 670 -1394 730 -834
rect 840 -1050 900 -722
rect 840 -1110 3214 -1050
rect 3154 -1274 3214 -1110
rect 5666 -1274 5726 -1268
rect 3154 -1278 5726 -1274
rect 3154 -1330 5670 -1278
rect 5722 -1330 5726 -1278
rect 3154 -1334 5726 -1330
rect 5666 -1340 5726 -1334
rect 3754 -1394 3814 -1388
rect 670 -1398 3814 -1394
rect 670 -1450 3758 -1398
rect 3810 -1450 3814 -1398
rect 670 -1454 3814 -1450
rect 3754 -1460 3814 -1454
rect 3892 -1400 3952 -1390
rect 3892 -1452 3896 -1400
rect 3948 -1452 3952 -1400
rect 5526 -1396 5598 -1392
rect 5526 -1448 5536 -1396
rect 5588 -1448 5598 -1396
rect 5526 -1452 5598 -1448
rect 3892 -1676 3952 -1452
rect 5532 -1674 5592 -1452
rect 3886 -1680 3958 -1676
rect 3886 -1732 3896 -1680
rect 3948 -1732 3958 -1680
rect 3886 -1736 3958 -1732
rect 5526 -1678 5598 -1674
rect 5526 -1730 5536 -1678
rect 5588 -1730 5598 -1678
rect 5526 -1734 5598 -1730
rect -48 -1788 12 -1782
rect 1670 -1788 1730 -1782
rect 2950 -1788 3010 -1782
rect 3388 -1788 3448 -1782
rect 5098 -1788 5158 -1782
rect -48 -1792 5158 -1788
rect -48 -1844 -44 -1792
rect 8 -1844 1674 -1792
rect 1726 -1844 2954 -1792
rect 3006 -1844 3392 -1792
rect 3444 -1844 5102 -1792
rect 5154 -1844 5158 -1792
rect -48 -1848 5158 -1844
rect -48 -1854 12 -1848
rect 1670 -1854 1730 -1848
rect 2950 -1854 3010 -1848
rect 3388 -1854 3448 -1848
rect 5098 -1854 5158 -1848
rect -908 -2340 -848 -2334
rect -476 -2340 -416 -2334
rect -52 -2340 8 -2334
rect 378 -2340 438 -2334
rect 810 -2340 870 -2334
rect 1230 -2340 1290 -2334
rect 2094 -2340 2154 -2334
rect 2950 -2340 3010 -2334
rect 3384 -2340 3444 -2334
rect 3818 -2340 3878 -2334
rect 4244 -2340 4304 -2334
rect 4666 -2340 4726 -2334
rect 5100 -2340 5160 -2334
rect -908 -2344 5160 -2340
rect -908 -2396 -904 -2344
rect -852 -2396 -472 -2344
rect -420 -2396 -48 -2344
rect 4 -2396 382 -2344
rect 434 -2396 814 -2344
rect 866 -2396 1234 -2344
rect 1286 -2396 2098 -2344
rect 2150 -2396 2954 -2344
rect 3006 -2396 3388 -2344
rect 3440 -2396 3822 -2344
rect 3874 -2396 4248 -2344
rect 4300 -2396 4670 -2344
rect 4722 -2396 5104 -2344
rect 5156 -2396 5160 -2344
rect -908 -2400 5160 -2396
rect -908 -2406 -848 -2400
rect -476 -2406 -416 -2400
rect -52 -2406 8 -2400
rect 378 -2406 438 -2400
rect 810 -2406 870 -2400
rect 1230 -2406 1290 -2400
rect 2094 -2406 2154 -2400
rect 2950 -2406 3010 -2400
rect 3384 -2406 3444 -2400
rect 3818 -2406 3878 -2400
rect 4244 -2406 4304 -2400
rect 4666 -2406 4726 -2400
rect 5100 -2406 5160 -2400
rect 1670 -2904 1730 -2898
rect 6378 -2904 6438 -28
rect 1670 -2908 6438 -2904
rect 1670 -2960 1674 -2908
rect 1726 -2960 6438 -2908
rect 1670 -2964 6438 -2960
rect 1670 -2970 1730 -2964
rect -1820 -3126 6120 -3082
rect -1820 -3136 -1759 -3126
rect 6057 -3136 6120 -3126
rect -1820 -3252 -1781 -3136
rect 6079 -3252 6120 -3136
rect -1820 -3262 -1759 -3252
rect 6057 -3262 6120 -3252
rect -1820 -3296 6120 -3262
rect -2416 -3378 -1816 -3366
rect -2416 -3404 -2384 -3378
rect -1848 -3404 -1816 -3378
rect -2416 -3648 -2398 -3404
rect -1834 -3648 -1816 -3404
rect -2416 -3674 -2384 -3648
rect -1848 -3674 -1816 -3648
rect -2416 -3686 -1816 -3674
rect 6216 -3378 6816 -3366
rect 6216 -3404 6248 -3378
rect 6784 -3404 6816 -3378
rect 6216 -3648 6234 -3404
rect 6798 -3648 6816 -3404
rect 6216 -3674 6248 -3648
rect 6784 -3674 6816 -3648
rect 6216 -3686 6816 -3674
<< via2 >>
rect -2384 2528 -1848 2554
rect -2384 2284 -1848 2528
rect -2384 2258 -1848 2284
rect 6248 2528 6784 2554
rect 6248 2284 6784 2528
rect 6248 2258 6784 2284
rect -2272 2111 -2216 2113
rect -2192 2111 -2136 2113
rect -2112 2111 -2056 2113
rect -2032 2111 -1976 2113
rect -1952 2111 -1896 2113
rect -1872 2111 -1816 2113
rect -1792 2111 -1736 2113
rect -1712 2111 -1656 2113
rect -1632 2111 -1576 2113
rect -1552 2111 -1496 2113
rect -1472 2111 -1416 2113
rect -1392 2111 -1336 2113
rect -1312 2111 -1256 2113
rect -1232 2111 -1176 2113
rect -1152 2111 -1096 2113
rect -1072 2111 -1016 2113
rect -992 2111 -936 2113
rect -912 2111 -856 2113
rect -832 2111 -776 2113
rect -752 2111 -696 2113
rect -672 2111 -616 2113
rect -592 2111 -536 2113
rect -512 2111 -456 2113
rect -432 2111 -376 2113
rect -352 2111 -296 2113
rect -272 2111 -216 2113
rect -192 2111 -136 2113
rect -112 2111 -56 2113
rect -32 2111 24 2113
rect 48 2111 104 2113
rect 128 2111 184 2113
rect 208 2111 264 2113
rect 288 2111 344 2113
rect 368 2111 424 2113
rect 448 2111 504 2113
rect 528 2111 584 2113
rect 608 2111 664 2113
rect 688 2111 744 2113
rect 768 2111 824 2113
rect 848 2111 904 2113
rect 928 2111 984 2113
rect 1008 2111 1064 2113
rect 1088 2111 1144 2113
rect 1168 2111 1224 2113
rect 1248 2111 1304 2113
rect 1328 2111 1384 2113
rect 1408 2111 1464 2113
rect 1488 2111 1544 2113
rect 1568 2111 1624 2113
rect 1648 2111 1704 2113
rect 1728 2111 1784 2113
rect 1808 2111 1864 2113
rect 1888 2111 1944 2113
rect 1968 2111 2024 2113
rect 2048 2111 2104 2113
rect 2128 2111 2184 2113
rect 2208 2111 2264 2113
rect 2288 2111 2344 2113
rect 2368 2111 2424 2113
rect 2448 2111 2504 2113
rect 2528 2111 2584 2113
rect 2608 2111 2664 2113
rect 2688 2111 2744 2113
rect 2768 2111 2824 2113
rect 2848 2111 2904 2113
rect 2928 2111 2984 2113
rect 3008 2111 3064 2113
rect 3088 2111 3144 2113
rect 3168 2111 3224 2113
rect 3248 2111 3304 2113
rect 3328 2111 3384 2113
rect 3408 2111 3464 2113
rect 3488 2111 3544 2113
rect 3568 2111 3624 2113
rect 3648 2111 3704 2113
rect 3728 2111 3784 2113
rect 3808 2111 3864 2113
rect 3888 2111 3944 2113
rect 3968 2111 4024 2113
rect 4048 2111 4104 2113
rect 4128 2111 4184 2113
rect 4208 2111 4264 2113
rect 4288 2111 4344 2113
rect 4368 2111 4424 2113
rect 4448 2111 4504 2113
rect 4528 2111 4584 2113
rect 4608 2111 4664 2113
rect 4688 2111 4744 2113
rect 4768 2111 4824 2113
rect 4848 2111 4904 2113
rect 4928 2111 4984 2113
rect 5008 2111 5064 2113
rect 5088 2111 5144 2113
rect 5168 2111 5224 2113
rect 5248 2111 5304 2113
rect 5328 2111 5384 2113
rect 5408 2111 5464 2113
rect 5488 2111 5544 2113
rect 5568 2111 5624 2113
rect 5648 2111 5704 2113
rect 5728 2111 5784 2113
rect 5808 2111 5864 2113
rect 5888 2111 5944 2113
rect 5968 2111 6024 2113
rect 6048 2111 6104 2113
rect 6128 2111 6184 2113
rect 6208 2111 6264 2113
rect 6288 2111 6344 2113
rect 6368 2111 6424 2113
rect 6448 2111 6504 2113
rect 6528 2111 6584 2113
rect 6608 2111 6664 2113
rect -2272 2059 -2226 2111
rect -2226 2059 -2216 2111
rect -2192 2059 -2162 2111
rect -2162 2059 -2150 2111
rect -2150 2059 -2136 2111
rect -2112 2059 -2098 2111
rect -2098 2059 -2086 2111
rect -2086 2059 -2056 2111
rect -2032 2059 -2022 2111
rect -2022 2059 -1976 2111
rect -1952 2059 -1906 2111
rect -1906 2059 -1896 2111
rect -1872 2059 -1842 2111
rect -1842 2059 -1830 2111
rect -1830 2059 -1816 2111
rect -1792 2059 -1778 2111
rect -1778 2059 -1766 2111
rect -1766 2059 -1736 2111
rect -1712 2059 -1702 2111
rect -1702 2059 -1656 2111
rect -1632 2059 -1586 2111
rect -1586 2059 -1576 2111
rect -1552 2059 -1522 2111
rect -1522 2059 -1510 2111
rect -1510 2059 -1496 2111
rect -1472 2059 -1458 2111
rect -1458 2059 -1446 2111
rect -1446 2059 -1416 2111
rect -1392 2059 -1382 2111
rect -1382 2059 -1336 2111
rect -1312 2059 -1266 2111
rect -1266 2059 -1256 2111
rect -1232 2059 -1202 2111
rect -1202 2059 -1190 2111
rect -1190 2059 -1176 2111
rect -1152 2059 -1138 2111
rect -1138 2059 -1126 2111
rect -1126 2059 -1096 2111
rect -1072 2059 -1062 2111
rect -1062 2059 -1016 2111
rect -992 2059 -946 2111
rect -946 2059 -936 2111
rect -912 2059 -882 2111
rect -882 2059 -870 2111
rect -870 2059 -856 2111
rect -832 2059 -818 2111
rect -818 2059 -806 2111
rect -806 2059 -776 2111
rect -752 2059 -742 2111
rect -742 2059 -696 2111
rect -672 2059 -626 2111
rect -626 2059 -616 2111
rect -592 2059 -562 2111
rect -562 2059 -550 2111
rect -550 2059 -536 2111
rect -512 2059 -498 2111
rect -498 2059 -486 2111
rect -486 2059 -456 2111
rect -432 2059 -422 2111
rect -422 2059 -376 2111
rect -352 2059 -306 2111
rect -306 2059 -296 2111
rect -272 2059 -242 2111
rect -242 2059 -230 2111
rect -230 2059 -216 2111
rect -192 2059 -178 2111
rect -178 2059 -166 2111
rect -166 2059 -136 2111
rect -112 2059 -102 2111
rect -102 2059 -56 2111
rect -32 2059 14 2111
rect 14 2059 24 2111
rect 48 2059 78 2111
rect 78 2059 90 2111
rect 90 2059 104 2111
rect 128 2059 142 2111
rect 142 2059 154 2111
rect 154 2059 184 2111
rect 208 2059 218 2111
rect 218 2059 264 2111
rect 288 2059 334 2111
rect 334 2059 344 2111
rect 368 2059 398 2111
rect 398 2059 410 2111
rect 410 2059 424 2111
rect 448 2059 462 2111
rect 462 2059 474 2111
rect 474 2059 504 2111
rect 528 2059 538 2111
rect 538 2059 584 2111
rect 608 2059 654 2111
rect 654 2059 664 2111
rect 688 2059 718 2111
rect 718 2059 730 2111
rect 730 2059 744 2111
rect 768 2059 782 2111
rect 782 2059 794 2111
rect 794 2059 824 2111
rect 848 2059 858 2111
rect 858 2059 904 2111
rect 928 2059 974 2111
rect 974 2059 984 2111
rect 1008 2059 1038 2111
rect 1038 2059 1050 2111
rect 1050 2059 1064 2111
rect 1088 2059 1102 2111
rect 1102 2059 1114 2111
rect 1114 2059 1144 2111
rect 1168 2059 1178 2111
rect 1178 2059 1224 2111
rect 1248 2059 1294 2111
rect 1294 2059 1304 2111
rect 1328 2059 1358 2111
rect 1358 2059 1370 2111
rect 1370 2059 1384 2111
rect 1408 2059 1422 2111
rect 1422 2059 1434 2111
rect 1434 2059 1464 2111
rect 1488 2059 1498 2111
rect 1498 2059 1544 2111
rect 1568 2059 1614 2111
rect 1614 2059 1624 2111
rect 1648 2059 1678 2111
rect 1678 2059 1690 2111
rect 1690 2059 1704 2111
rect 1728 2059 1742 2111
rect 1742 2059 1754 2111
rect 1754 2059 1784 2111
rect 1808 2059 1818 2111
rect 1818 2059 1864 2111
rect 1888 2059 1934 2111
rect 1934 2059 1944 2111
rect 1968 2059 1998 2111
rect 1998 2059 2010 2111
rect 2010 2059 2024 2111
rect 2048 2059 2062 2111
rect 2062 2059 2074 2111
rect 2074 2059 2104 2111
rect 2128 2059 2138 2111
rect 2138 2059 2184 2111
rect 2208 2059 2254 2111
rect 2254 2059 2264 2111
rect 2288 2059 2318 2111
rect 2318 2059 2330 2111
rect 2330 2059 2344 2111
rect 2368 2059 2382 2111
rect 2382 2059 2394 2111
rect 2394 2059 2424 2111
rect 2448 2059 2458 2111
rect 2458 2059 2504 2111
rect 2528 2059 2574 2111
rect 2574 2059 2584 2111
rect 2608 2059 2638 2111
rect 2638 2059 2650 2111
rect 2650 2059 2664 2111
rect 2688 2059 2702 2111
rect 2702 2059 2714 2111
rect 2714 2059 2744 2111
rect 2768 2059 2778 2111
rect 2778 2059 2824 2111
rect 2848 2059 2894 2111
rect 2894 2059 2904 2111
rect 2928 2059 2958 2111
rect 2958 2059 2970 2111
rect 2970 2059 2984 2111
rect 3008 2059 3022 2111
rect 3022 2059 3034 2111
rect 3034 2059 3064 2111
rect 3088 2059 3098 2111
rect 3098 2059 3144 2111
rect 3168 2059 3214 2111
rect 3214 2059 3224 2111
rect 3248 2059 3278 2111
rect 3278 2059 3290 2111
rect 3290 2059 3304 2111
rect 3328 2059 3342 2111
rect 3342 2059 3354 2111
rect 3354 2059 3384 2111
rect 3408 2059 3418 2111
rect 3418 2059 3464 2111
rect 3488 2059 3534 2111
rect 3534 2059 3544 2111
rect 3568 2059 3598 2111
rect 3598 2059 3610 2111
rect 3610 2059 3624 2111
rect 3648 2059 3662 2111
rect 3662 2059 3674 2111
rect 3674 2059 3704 2111
rect 3728 2059 3738 2111
rect 3738 2059 3784 2111
rect 3808 2059 3854 2111
rect 3854 2059 3864 2111
rect 3888 2059 3918 2111
rect 3918 2059 3930 2111
rect 3930 2059 3944 2111
rect 3968 2059 3982 2111
rect 3982 2059 3994 2111
rect 3994 2059 4024 2111
rect 4048 2059 4058 2111
rect 4058 2059 4104 2111
rect 4128 2059 4174 2111
rect 4174 2059 4184 2111
rect 4208 2059 4238 2111
rect 4238 2059 4250 2111
rect 4250 2059 4264 2111
rect 4288 2059 4302 2111
rect 4302 2059 4314 2111
rect 4314 2059 4344 2111
rect 4368 2059 4378 2111
rect 4378 2059 4424 2111
rect 4448 2059 4494 2111
rect 4494 2059 4504 2111
rect 4528 2059 4558 2111
rect 4558 2059 4570 2111
rect 4570 2059 4584 2111
rect 4608 2059 4622 2111
rect 4622 2059 4634 2111
rect 4634 2059 4664 2111
rect 4688 2059 4698 2111
rect 4698 2059 4744 2111
rect 4768 2059 4814 2111
rect 4814 2059 4824 2111
rect 4848 2059 4878 2111
rect 4878 2059 4890 2111
rect 4890 2059 4904 2111
rect 4928 2059 4942 2111
rect 4942 2059 4954 2111
rect 4954 2059 4984 2111
rect 5008 2059 5018 2111
rect 5018 2059 5064 2111
rect 5088 2059 5134 2111
rect 5134 2059 5144 2111
rect 5168 2059 5198 2111
rect 5198 2059 5210 2111
rect 5210 2059 5224 2111
rect 5248 2059 5262 2111
rect 5262 2059 5274 2111
rect 5274 2059 5304 2111
rect 5328 2059 5338 2111
rect 5338 2059 5384 2111
rect 5408 2059 5454 2111
rect 5454 2059 5464 2111
rect 5488 2059 5518 2111
rect 5518 2059 5530 2111
rect 5530 2059 5544 2111
rect 5568 2059 5582 2111
rect 5582 2059 5594 2111
rect 5594 2059 5624 2111
rect 5648 2059 5658 2111
rect 5658 2059 5704 2111
rect 5728 2059 5774 2111
rect 5774 2059 5784 2111
rect 5808 2059 5838 2111
rect 5838 2059 5850 2111
rect 5850 2059 5864 2111
rect 5888 2059 5902 2111
rect 5902 2059 5914 2111
rect 5914 2059 5944 2111
rect 5968 2059 5978 2111
rect 5978 2059 6024 2111
rect 6048 2059 6094 2111
rect 6094 2059 6104 2111
rect 6128 2059 6158 2111
rect 6158 2059 6170 2111
rect 6170 2059 6184 2111
rect 6208 2059 6222 2111
rect 6222 2059 6234 2111
rect 6234 2059 6264 2111
rect 6288 2059 6298 2111
rect 6298 2059 6344 2111
rect 6368 2059 6414 2111
rect 6414 2059 6424 2111
rect 6448 2059 6478 2111
rect 6478 2059 6490 2111
rect 6490 2059 6504 2111
rect 6528 2059 6542 2111
rect 6542 2059 6554 2111
rect 6554 2059 6584 2111
rect 6608 2059 6618 2111
rect 6618 2059 6664 2111
rect -2272 2057 -2216 2059
rect -2192 2057 -2136 2059
rect -2112 2057 -2056 2059
rect -2032 2057 -1976 2059
rect -1952 2057 -1896 2059
rect -1872 2057 -1816 2059
rect -1792 2057 -1736 2059
rect -1712 2057 -1656 2059
rect -1632 2057 -1576 2059
rect -1552 2057 -1496 2059
rect -1472 2057 -1416 2059
rect -1392 2057 -1336 2059
rect -1312 2057 -1256 2059
rect -1232 2057 -1176 2059
rect -1152 2057 -1096 2059
rect -1072 2057 -1016 2059
rect -992 2057 -936 2059
rect -912 2057 -856 2059
rect -832 2057 -776 2059
rect -752 2057 -696 2059
rect -672 2057 -616 2059
rect -592 2057 -536 2059
rect -512 2057 -456 2059
rect -432 2057 -376 2059
rect -352 2057 -296 2059
rect -272 2057 -216 2059
rect -192 2057 -136 2059
rect -112 2057 -56 2059
rect -32 2057 24 2059
rect 48 2057 104 2059
rect 128 2057 184 2059
rect 208 2057 264 2059
rect 288 2057 344 2059
rect 368 2057 424 2059
rect 448 2057 504 2059
rect 528 2057 584 2059
rect 608 2057 664 2059
rect 688 2057 744 2059
rect 768 2057 824 2059
rect 848 2057 904 2059
rect 928 2057 984 2059
rect 1008 2057 1064 2059
rect 1088 2057 1144 2059
rect 1168 2057 1224 2059
rect 1248 2057 1304 2059
rect 1328 2057 1384 2059
rect 1408 2057 1464 2059
rect 1488 2057 1544 2059
rect 1568 2057 1624 2059
rect 1648 2057 1704 2059
rect 1728 2057 1784 2059
rect 1808 2057 1864 2059
rect 1888 2057 1944 2059
rect 1968 2057 2024 2059
rect 2048 2057 2104 2059
rect 2128 2057 2184 2059
rect 2208 2057 2264 2059
rect 2288 2057 2344 2059
rect 2368 2057 2424 2059
rect 2448 2057 2504 2059
rect 2528 2057 2584 2059
rect 2608 2057 2664 2059
rect 2688 2057 2744 2059
rect 2768 2057 2824 2059
rect 2848 2057 2904 2059
rect 2928 2057 2984 2059
rect 3008 2057 3064 2059
rect 3088 2057 3144 2059
rect 3168 2057 3224 2059
rect 3248 2057 3304 2059
rect 3328 2057 3384 2059
rect 3408 2057 3464 2059
rect 3488 2057 3544 2059
rect 3568 2057 3624 2059
rect 3648 2057 3704 2059
rect 3728 2057 3784 2059
rect 3808 2057 3864 2059
rect 3888 2057 3944 2059
rect 3968 2057 4024 2059
rect 4048 2057 4104 2059
rect 4128 2057 4184 2059
rect 4208 2057 4264 2059
rect 4288 2057 4344 2059
rect 4368 2057 4424 2059
rect 4448 2057 4504 2059
rect 4528 2057 4584 2059
rect 4608 2057 4664 2059
rect 4688 2057 4744 2059
rect 4768 2057 4824 2059
rect 4848 2057 4904 2059
rect 4928 2057 4984 2059
rect 5008 2057 5064 2059
rect 5088 2057 5144 2059
rect 5168 2057 5224 2059
rect 5248 2057 5304 2059
rect 5328 2057 5384 2059
rect 5408 2057 5464 2059
rect 5488 2057 5544 2059
rect 5568 2057 5624 2059
rect 5648 2057 5704 2059
rect 5728 2057 5784 2059
rect 5808 2057 5864 2059
rect 5888 2057 5944 2059
rect 5968 2057 6024 2059
rect 6048 2057 6104 2059
rect 6128 2057 6184 2059
rect 6208 2057 6264 2059
rect 6288 2057 6344 2059
rect 6368 2057 6424 2059
rect 6448 2057 6504 2059
rect 6528 2057 6584 2059
rect 6608 2057 6664 2059
rect -1759 -3136 6057 -3126
rect -1759 -3252 6057 -3136
rect -1759 -3262 6057 -3252
rect -2384 -3404 -1848 -3378
rect -2384 -3648 -1848 -3404
rect -2384 -3674 -1848 -3648
rect 6248 -3404 6784 -3378
rect 6248 -3648 6784 -3404
rect 6248 -3674 6784 -3648
<< metal3 >>
rect -2426 2554 -1806 2561
rect -2426 2518 -2384 2554
rect -1848 2518 -1806 2554
rect -2426 2294 -2388 2518
rect -1844 2294 -1806 2518
rect -2426 2258 -2384 2294
rect -1848 2258 -1806 2294
rect -2426 2251 -1806 2258
rect 6206 2554 6826 2561
rect 6206 2518 6248 2554
rect 6784 2518 6826 2554
rect 6206 2294 6244 2518
rect 6788 2294 6826 2518
rect 6206 2258 6248 2294
rect 6784 2258 6826 2294
rect 6206 2251 6826 2258
rect -2340 2117 6730 2174
rect -2340 2053 -2276 2117
rect -2212 2053 -2196 2117
rect -2132 2053 -2116 2117
rect -2052 2053 -2036 2117
rect -1972 2053 -1956 2117
rect -1892 2053 -1876 2117
rect -1812 2053 -1796 2117
rect -1732 2053 -1716 2117
rect -1652 2053 -1636 2117
rect -1572 2053 -1556 2117
rect -1492 2053 -1476 2117
rect -1412 2053 -1396 2117
rect -1332 2053 -1316 2117
rect -1252 2053 -1236 2117
rect -1172 2053 -1156 2117
rect -1092 2053 -1076 2117
rect -1012 2053 -996 2117
rect -932 2053 -916 2117
rect -852 2053 -836 2117
rect -772 2053 -756 2117
rect -692 2053 -676 2117
rect -612 2053 -596 2117
rect -532 2053 -516 2117
rect -452 2053 -436 2117
rect -372 2053 -356 2117
rect -292 2053 -276 2117
rect -212 2053 -196 2117
rect -132 2053 -116 2117
rect -52 2053 -36 2117
rect 28 2053 44 2117
rect 108 2053 124 2117
rect 188 2053 204 2117
rect 268 2053 284 2117
rect 348 2053 364 2117
rect 428 2053 444 2117
rect 508 2053 524 2117
rect 588 2053 604 2117
rect 668 2053 684 2117
rect 748 2053 764 2117
rect 828 2053 844 2117
rect 908 2053 924 2117
rect 988 2053 1004 2117
rect 1068 2053 1084 2117
rect 1148 2053 1164 2117
rect 1228 2053 1244 2117
rect 1308 2053 1324 2117
rect 1388 2053 1404 2117
rect 1468 2053 1484 2117
rect 1548 2053 1564 2117
rect 1628 2053 1644 2117
rect 1708 2053 1724 2117
rect 1788 2053 1804 2117
rect 1868 2053 1884 2117
rect 1948 2053 1964 2117
rect 2028 2053 2044 2117
rect 2108 2053 2124 2117
rect 2188 2053 2204 2117
rect 2268 2053 2284 2117
rect 2348 2053 2364 2117
rect 2428 2053 2444 2117
rect 2508 2053 2524 2117
rect 2588 2053 2604 2117
rect 2668 2053 2684 2117
rect 2748 2053 2764 2117
rect 2828 2053 2844 2117
rect 2908 2053 2924 2117
rect 2988 2053 3004 2117
rect 3068 2053 3084 2117
rect 3148 2053 3164 2117
rect 3228 2053 3244 2117
rect 3308 2053 3324 2117
rect 3388 2053 3404 2117
rect 3468 2053 3484 2117
rect 3548 2053 3564 2117
rect 3628 2053 3644 2117
rect 3708 2053 3724 2117
rect 3788 2053 3804 2117
rect 3868 2053 3884 2117
rect 3948 2053 3964 2117
rect 4028 2053 4044 2117
rect 4108 2053 4124 2117
rect 4188 2053 4204 2117
rect 4268 2053 4284 2117
rect 4348 2053 4364 2117
rect 4428 2053 4444 2117
rect 4508 2053 4524 2117
rect 4588 2053 4604 2117
rect 4668 2053 4684 2117
rect 4748 2053 4764 2117
rect 4828 2053 4844 2117
rect 4908 2053 4924 2117
rect 4988 2053 5004 2117
rect 5068 2053 5084 2117
rect 5148 2053 5164 2117
rect 5228 2053 5244 2117
rect 5308 2053 5324 2117
rect 5388 2053 5404 2117
rect 5468 2053 5484 2117
rect 5548 2053 5564 2117
rect 5628 2053 5644 2117
rect 5708 2053 5724 2117
rect 5788 2053 5804 2117
rect 5868 2053 5884 2117
rect 5948 2053 5964 2117
rect 6028 2053 6044 2117
rect 6108 2053 6124 2117
rect 6188 2053 6204 2117
rect 6268 2053 6284 2117
rect 6348 2053 6364 2117
rect 6428 2053 6444 2117
rect 6508 2053 6524 2117
rect 6588 2053 6604 2117
rect 6668 2053 6730 2117
rect -2340 1992 6730 2053
rect -1820 -3122 6120 -3082
rect -1820 -3266 -1763 -3122
rect 6061 -3266 6120 -3122
rect -1820 -3296 6120 -3266
rect -2426 -3378 -1806 -3371
rect -2426 -3414 -2384 -3378
rect -1848 -3414 -1806 -3378
rect -2426 -3638 -2388 -3414
rect -1844 -3638 -1806 -3414
rect -2426 -3674 -2384 -3638
rect -1848 -3674 -1806 -3638
rect -2426 -3681 -1806 -3674
rect 6206 -3378 6826 -3371
rect 6206 -3414 6248 -3378
rect 6784 -3414 6826 -3378
rect 6206 -3638 6244 -3414
rect 6788 -3638 6826 -3414
rect 6206 -3674 6248 -3638
rect 6784 -3674 6826 -3638
rect 6206 -3681 6826 -3674
<< via3 >>
rect -2388 2294 -2384 2518
rect -2384 2294 -1848 2518
rect -1848 2294 -1844 2518
rect 6244 2294 6248 2518
rect 6248 2294 6784 2518
rect 6784 2294 6788 2518
rect -2276 2113 -2212 2117
rect -2276 2057 -2272 2113
rect -2272 2057 -2216 2113
rect -2216 2057 -2212 2113
rect -2276 2053 -2212 2057
rect -2196 2113 -2132 2117
rect -2196 2057 -2192 2113
rect -2192 2057 -2136 2113
rect -2136 2057 -2132 2113
rect -2196 2053 -2132 2057
rect -2116 2113 -2052 2117
rect -2116 2057 -2112 2113
rect -2112 2057 -2056 2113
rect -2056 2057 -2052 2113
rect -2116 2053 -2052 2057
rect -2036 2113 -1972 2117
rect -2036 2057 -2032 2113
rect -2032 2057 -1976 2113
rect -1976 2057 -1972 2113
rect -2036 2053 -1972 2057
rect -1956 2113 -1892 2117
rect -1956 2057 -1952 2113
rect -1952 2057 -1896 2113
rect -1896 2057 -1892 2113
rect -1956 2053 -1892 2057
rect -1876 2113 -1812 2117
rect -1876 2057 -1872 2113
rect -1872 2057 -1816 2113
rect -1816 2057 -1812 2113
rect -1876 2053 -1812 2057
rect -1796 2113 -1732 2117
rect -1796 2057 -1792 2113
rect -1792 2057 -1736 2113
rect -1736 2057 -1732 2113
rect -1796 2053 -1732 2057
rect -1716 2113 -1652 2117
rect -1716 2057 -1712 2113
rect -1712 2057 -1656 2113
rect -1656 2057 -1652 2113
rect -1716 2053 -1652 2057
rect -1636 2113 -1572 2117
rect -1636 2057 -1632 2113
rect -1632 2057 -1576 2113
rect -1576 2057 -1572 2113
rect -1636 2053 -1572 2057
rect -1556 2113 -1492 2117
rect -1556 2057 -1552 2113
rect -1552 2057 -1496 2113
rect -1496 2057 -1492 2113
rect -1556 2053 -1492 2057
rect -1476 2113 -1412 2117
rect -1476 2057 -1472 2113
rect -1472 2057 -1416 2113
rect -1416 2057 -1412 2113
rect -1476 2053 -1412 2057
rect -1396 2113 -1332 2117
rect -1396 2057 -1392 2113
rect -1392 2057 -1336 2113
rect -1336 2057 -1332 2113
rect -1396 2053 -1332 2057
rect -1316 2113 -1252 2117
rect -1316 2057 -1312 2113
rect -1312 2057 -1256 2113
rect -1256 2057 -1252 2113
rect -1316 2053 -1252 2057
rect -1236 2113 -1172 2117
rect -1236 2057 -1232 2113
rect -1232 2057 -1176 2113
rect -1176 2057 -1172 2113
rect -1236 2053 -1172 2057
rect -1156 2113 -1092 2117
rect -1156 2057 -1152 2113
rect -1152 2057 -1096 2113
rect -1096 2057 -1092 2113
rect -1156 2053 -1092 2057
rect -1076 2113 -1012 2117
rect -1076 2057 -1072 2113
rect -1072 2057 -1016 2113
rect -1016 2057 -1012 2113
rect -1076 2053 -1012 2057
rect -996 2113 -932 2117
rect -996 2057 -992 2113
rect -992 2057 -936 2113
rect -936 2057 -932 2113
rect -996 2053 -932 2057
rect -916 2113 -852 2117
rect -916 2057 -912 2113
rect -912 2057 -856 2113
rect -856 2057 -852 2113
rect -916 2053 -852 2057
rect -836 2113 -772 2117
rect -836 2057 -832 2113
rect -832 2057 -776 2113
rect -776 2057 -772 2113
rect -836 2053 -772 2057
rect -756 2113 -692 2117
rect -756 2057 -752 2113
rect -752 2057 -696 2113
rect -696 2057 -692 2113
rect -756 2053 -692 2057
rect -676 2113 -612 2117
rect -676 2057 -672 2113
rect -672 2057 -616 2113
rect -616 2057 -612 2113
rect -676 2053 -612 2057
rect -596 2113 -532 2117
rect -596 2057 -592 2113
rect -592 2057 -536 2113
rect -536 2057 -532 2113
rect -596 2053 -532 2057
rect -516 2113 -452 2117
rect -516 2057 -512 2113
rect -512 2057 -456 2113
rect -456 2057 -452 2113
rect -516 2053 -452 2057
rect -436 2113 -372 2117
rect -436 2057 -432 2113
rect -432 2057 -376 2113
rect -376 2057 -372 2113
rect -436 2053 -372 2057
rect -356 2113 -292 2117
rect -356 2057 -352 2113
rect -352 2057 -296 2113
rect -296 2057 -292 2113
rect -356 2053 -292 2057
rect -276 2113 -212 2117
rect -276 2057 -272 2113
rect -272 2057 -216 2113
rect -216 2057 -212 2113
rect -276 2053 -212 2057
rect -196 2113 -132 2117
rect -196 2057 -192 2113
rect -192 2057 -136 2113
rect -136 2057 -132 2113
rect -196 2053 -132 2057
rect -116 2113 -52 2117
rect -116 2057 -112 2113
rect -112 2057 -56 2113
rect -56 2057 -52 2113
rect -116 2053 -52 2057
rect -36 2113 28 2117
rect -36 2057 -32 2113
rect -32 2057 24 2113
rect 24 2057 28 2113
rect -36 2053 28 2057
rect 44 2113 108 2117
rect 44 2057 48 2113
rect 48 2057 104 2113
rect 104 2057 108 2113
rect 44 2053 108 2057
rect 124 2113 188 2117
rect 124 2057 128 2113
rect 128 2057 184 2113
rect 184 2057 188 2113
rect 124 2053 188 2057
rect 204 2113 268 2117
rect 204 2057 208 2113
rect 208 2057 264 2113
rect 264 2057 268 2113
rect 204 2053 268 2057
rect 284 2113 348 2117
rect 284 2057 288 2113
rect 288 2057 344 2113
rect 344 2057 348 2113
rect 284 2053 348 2057
rect 364 2113 428 2117
rect 364 2057 368 2113
rect 368 2057 424 2113
rect 424 2057 428 2113
rect 364 2053 428 2057
rect 444 2113 508 2117
rect 444 2057 448 2113
rect 448 2057 504 2113
rect 504 2057 508 2113
rect 444 2053 508 2057
rect 524 2113 588 2117
rect 524 2057 528 2113
rect 528 2057 584 2113
rect 584 2057 588 2113
rect 524 2053 588 2057
rect 604 2113 668 2117
rect 604 2057 608 2113
rect 608 2057 664 2113
rect 664 2057 668 2113
rect 604 2053 668 2057
rect 684 2113 748 2117
rect 684 2057 688 2113
rect 688 2057 744 2113
rect 744 2057 748 2113
rect 684 2053 748 2057
rect 764 2113 828 2117
rect 764 2057 768 2113
rect 768 2057 824 2113
rect 824 2057 828 2113
rect 764 2053 828 2057
rect 844 2113 908 2117
rect 844 2057 848 2113
rect 848 2057 904 2113
rect 904 2057 908 2113
rect 844 2053 908 2057
rect 924 2113 988 2117
rect 924 2057 928 2113
rect 928 2057 984 2113
rect 984 2057 988 2113
rect 924 2053 988 2057
rect 1004 2113 1068 2117
rect 1004 2057 1008 2113
rect 1008 2057 1064 2113
rect 1064 2057 1068 2113
rect 1004 2053 1068 2057
rect 1084 2113 1148 2117
rect 1084 2057 1088 2113
rect 1088 2057 1144 2113
rect 1144 2057 1148 2113
rect 1084 2053 1148 2057
rect 1164 2113 1228 2117
rect 1164 2057 1168 2113
rect 1168 2057 1224 2113
rect 1224 2057 1228 2113
rect 1164 2053 1228 2057
rect 1244 2113 1308 2117
rect 1244 2057 1248 2113
rect 1248 2057 1304 2113
rect 1304 2057 1308 2113
rect 1244 2053 1308 2057
rect 1324 2113 1388 2117
rect 1324 2057 1328 2113
rect 1328 2057 1384 2113
rect 1384 2057 1388 2113
rect 1324 2053 1388 2057
rect 1404 2113 1468 2117
rect 1404 2057 1408 2113
rect 1408 2057 1464 2113
rect 1464 2057 1468 2113
rect 1404 2053 1468 2057
rect 1484 2113 1548 2117
rect 1484 2057 1488 2113
rect 1488 2057 1544 2113
rect 1544 2057 1548 2113
rect 1484 2053 1548 2057
rect 1564 2113 1628 2117
rect 1564 2057 1568 2113
rect 1568 2057 1624 2113
rect 1624 2057 1628 2113
rect 1564 2053 1628 2057
rect 1644 2113 1708 2117
rect 1644 2057 1648 2113
rect 1648 2057 1704 2113
rect 1704 2057 1708 2113
rect 1644 2053 1708 2057
rect 1724 2113 1788 2117
rect 1724 2057 1728 2113
rect 1728 2057 1784 2113
rect 1784 2057 1788 2113
rect 1724 2053 1788 2057
rect 1804 2113 1868 2117
rect 1804 2057 1808 2113
rect 1808 2057 1864 2113
rect 1864 2057 1868 2113
rect 1804 2053 1868 2057
rect 1884 2113 1948 2117
rect 1884 2057 1888 2113
rect 1888 2057 1944 2113
rect 1944 2057 1948 2113
rect 1884 2053 1948 2057
rect 1964 2113 2028 2117
rect 1964 2057 1968 2113
rect 1968 2057 2024 2113
rect 2024 2057 2028 2113
rect 1964 2053 2028 2057
rect 2044 2113 2108 2117
rect 2044 2057 2048 2113
rect 2048 2057 2104 2113
rect 2104 2057 2108 2113
rect 2044 2053 2108 2057
rect 2124 2113 2188 2117
rect 2124 2057 2128 2113
rect 2128 2057 2184 2113
rect 2184 2057 2188 2113
rect 2124 2053 2188 2057
rect 2204 2113 2268 2117
rect 2204 2057 2208 2113
rect 2208 2057 2264 2113
rect 2264 2057 2268 2113
rect 2204 2053 2268 2057
rect 2284 2113 2348 2117
rect 2284 2057 2288 2113
rect 2288 2057 2344 2113
rect 2344 2057 2348 2113
rect 2284 2053 2348 2057
rect 2364 2113 2428 2117
rect 2364 2057 2368 2113
rect 2368 2057 2424 2113
rect 2424 2057 2428 2113
rect 2364 2053 2428 2057
rect 2444 2113 2508 2117
rect 2444 2057 2448 2113
rect 2448 2057 2504 2113
rect 2504 2057 2508 2113
rect 2444 2053 2508 2057
rect 2524 2113 2588 2117
rect 2524 2057 2528 2113
rect 2528 2057 2584 2113
rect 2584 2057 2588 2113
rect 2524 2053 2588 2057
rect 2604 2113 2668 2117
rect 2604 2057 2608 2113
rect 2608 2057 2664 2113
rect 2664 2057 2668 2113
rect 2604 2053 2668 2057
rect 2684 2113 2748 2117
rect 2684 2057 2688 2113
rect 2688 2057 2744 2113
rect 2744 2057 2748 2113
rect 2684 2053 2748 2057
rect 2764 2113 2828 2117
rect 2764 2057 2768 2113
rect 2768 2057 2824 2113
rect 2824 2057 2828 2113
rect 2764 2053 2828 2057
rect 2844 2113 2908 2117
rect 2844 2057 2848 2113
rect 2848 2057 2904 2113
rect 2904 2057 2908 2113
rect 2844 2053 2908 2057
rect 2924 2113 2988 2117
rect 2924 2057 2928 2113
rect 2928 2057 2984 2113
rect 2984 2057 2988 2113
rect 2924 2053 2988 2057
rect 3004 2113 3068 2117
rect 3004 2057 3008 2113
rect 3008 2057 3064 2113
rect 3064 2057 3068 2113
rect 3004 2053 3068 2057
rect 3084 2113 3148 2117
rect 3084 2057 3088 2113
rect 3088 2057 3144 2113
rect 3144 2057 3148 2113
rect 3084 2053 3148 2057
rect 3164 2113 3228 2117
rect 3164 2057 3168 2113
rect 3168 2057 3224 2113
rect 3224 2057 3228 2113
rect 3164 2053 3228 2057
rect 3244 2113 3308 2117
rect 3244 2057 3248 2113
rect 3248 2057 3304 2113
rect 3304 2057 3308 2113
rect 3244 2053 3308 2057
rect 3324 2113 3388 2117
rect 3324 2057 3328 2113
rect 3328 2057 3384 2113
rect 3384 2057 3388 2113
rect 3324 2053 3388 2057
rect 3404 2113 3468 2117
rect 3404 2057 3408 2113
rect 3408 2057 3464 2113
rect 3464 2057 3468 2113
rect 3404 2053 3468 2057
rect 3484 2113 3548 2117
rect 3484 2057 3488 2113
rect 3488 2057 3544 2113
rect 3544 2057 3548 2113
rect 3484 2053 3548 2057
rect 3564 2113 3628 2117
rect 3564 2057 3568 2113
rect 3568 2057 3624 2113
rect 3624 2057 3628 2113
rect 3564 2053 3628 2057
rect 3644 2113 3708 2117
rect 3644 2057 3648 2113
rect 3648 2057 3704 2113
rect 3704 2057 3708 2113
rect 3644 2053 3708 2057
rect 3724 2113 3788 2117
rect 3724 2057 3728 2113
rect 3728 2057 3784 2113
rect 3784 2057 3788 2113
rect 3724 2053 3788 2057
rect 3804 2113 3868 2117
rect 3804 2057 3808 2113
rect 3808 2057 3864 2113
rect 3864 2057 3868 2113
rect 3804 2053 3868 2057
rect 3884 2113 3948 2117
rect 3884 2057 3888 2113
rect 3888 2057 3944 2113
rect 3944 2057 3948 2113
rect 3884 2053 3948 2057
rect 3964 2113 4028 2117
rect 3964 2057 3968 2113
rect 3968 2057 4024 2113
rect 4024 2057 4028 2113
rect 3964 2053 4028 2057
rect 4044 2113 4108 2117
rect 4044 2057 4048 2113
rect 4048 2057 4104 2113
rect 4104 2057 4108 2113
rect 4044 2053 4108 2057
rect 4124 2113 4188 2117
rect 4124 2057 4128 2113
rect 4128 2057 4184 2113
rect 4184 2057 4188 2113
rect 4124 2053 4188 2057
rect 4204 2113 4268 2117
rect 4204 2057 4208 2113
rect 4208 2057 4264 2113
rect 4264 2057 4268 2113
rect 4204 2053 4268 2057
rect 4284 2113 4348 2117
rect 4284 2057 4288 2113
rect 4288 2057 4344 2113
rect 4344 2057 4348 2113
rect 4284 2053 4348 2057
rect 4364 2113 4428 2117
rect 4364 2057 4368 2113
rect 4368 2057 4424 2113
rect 4424 2057 4428 2113
rect 4364 2053 4428 2057
rect 4444 2113 4508 2117
rect 4444 2057 4448 2113
rect 4448 2057 4504 2113
rect 4504 2057 4508 2113
rect 4444 2053 4508 2057
rect 4524 2113 4588 2117
rect 4524 2057 4528 2113
rect 4528 2057 4584 2113
rect 4584 2057 4588 2113
rect 4524 2053 4588 2057
rect 4604 2113 4668 2117
rect 4604 2057 4608 2113
rect 4608 2057 4664 2113
rect 4664 2057 4668 2113
rect 4604 2053 4668 2057
rect 4684 2113 4748 2117
rect 4684 2057 4688 2113
rect 4688 2057 4744 2113
rect 4744 2057 4748 2113
rect 4684 2053 4748 2057
rect 4764 2113 4828 2117
rect 4764 2057 4768 2113
rect 4768 2057 4824 2113
rect 4824 2057 4828 2113
rect 4764 2053 4828 2057
rect 4844 2113 4908 2117
rect 4844 2057 4848 2113
rect 4848 2057 4904 2113
rect 4904 2057 4908 2113
rect 4844 2053 4908 2057
rect 4924 2113 4988 2117
rect 4924 2057 4928 2113
rect 4928 2057 4984 2113
rect 4984 2057 4988 2113
rect 4924 2053 4988 2057
rect 5004 2113 5068 2117
rect 5004 2057 5008 2113
rect 5008 2057 5064 2113
rect 5064 2057 5068 2113
rect 5004 2053 5068 2057
rect 5084 2113 5148 2117
rect 5084 2057 5088 2113
rect 5088 2057 5144 2113
rect 5144 2057 5148 2113
rect 5084 2053 5148 2057
rect 5164 2113 5228 2117
rect 5164 2057 5168 2113
rect 5168 2057 5224 2113
rect 5224 2057 5228 2113
rect 5164 2053 5228 2057
rect 5244 2113 5308 2117
rect 5244 2057 5248 2113
rect 5248 2057 5304 2113
rect 5304 2057 5308 2113
rect 5244 2053 5308 2057
rect 5324 2113 5388 2117
rect 5324 2057 5328 2113
rect 5328 2057 5384 2113
rect 5384 2057 5388 2113
rect 5324 2053 5388 2057
rect 5404 2113 5468 2117
rect 5404 2057 5408 2113
rect 5408 2057 5464 2113
rect 5464 2057 5468 2113
rect 5404 2053 5468 2057
rect 5484 2113 5548 2117
rect 5484 2057 5488 2113
rect 5488 2057 5544 2113
rect 5544 2057 5548 2113
rect 5484 2053 5548 2057
rect 5564 2113 5628 2117
rect 5564 2057 5568 2113
rect 5568 2057 5624 2113
rect 5624 2057 5628 2113
rect 5564 2053 5628 2057
rect 5644 2113 5708 2117
rect 5644 2057 5648 2113
rect 5648 2057 5704 2113
rect 5704 2057 5708 2113
rect 5644 2053 5708 2057
rect 5724 2113 5788 2117
rect 5724 2057 5728 2113
rect 5728 2057 5784 2113
rect 5784 2057 5788 2113
rect 5724 2053 5788 2057
rect 5804 2113 5868 2117
rect 5804 2057 5808 2113
rect 5808 2057 5864 2113
rect 5864 2057 5868 2113
rect 5804 2053 5868 2057
rect 5884 2113 5948 2117
rect 5884 2057 5888 2113
rect 5888 2057 5944 2113
rect 5944 2057 5948 2113
rect 5884 2053 5948 2057
rect 5964 2113 6028 2117
rect 5964 2057 5968 2113
rect 5968 2057 6024 2113
rect 6024 2057 6028 2113
rect 5964 2053 6028 2057
rect 6044 2113 6108 2117
rect 6044 2057 6048 2113
rect 6048 2057 6104 2113
rect 6104 2057 6108 2113
rect 6044 2053 6108 2057
rect 6124 2113 6188 2117
rect 6124 2057 6128 2113
rect 6128 2057 6184 2113
rect 6184 2057 6188 2113
rect 6124 2053 6188 2057
rect 6204 2113 6268 2117
rect 6204 2057 6208 2113
rect 6208 2057 6264 2113
rect 6264 2057 6268 2113
rect 6204 2053 6268 2057
rect 6284 2113 6348 2117
rect 6284 2057 6288 2113
rect 6288 2057 6344 2113
rect 6344 2057 6348 2113
rect 6284 2053 6348 2057
rect 6364 2113 6428 2117
rect 6364 2057 6368 2113
rect 6368 2057 6424 2113
rect 6424 2057 6428 2113
rect 6364 2053 6428 2057
rect 6444 2113 6508 2117
rect 6444 2057 6448 2113
rect 6448 2057 6504 2113
rect 6504 2057 6508 2113
rect 6444 2053 6508 2057
rect 6524 2113 6588 2117
rect 6524 2057 6528 2113
rect 6528 2057 6584 2113
rect 6584 2057 6588 2113
rect 6524 2053 6588 2057
rect 6604 2113 6668 2117
rect 6604 2057 6608 2113
rect 6608 2057 6664 2113
rect 6664 2057 6668 2113
rect 6604 2053 6668 2057
rect -1763 -3126 6061 -3122
rect -1763 -3262 -1759 -3126
rect -1759 -3262 6057 -3126
rect 6057 -3262 6061 -3126
rect -1763 -3266 6061 -3262
rect -2388 -3638 -2384 -3414
rect -2384 -3638 -1848 -3414
rect -1848 -3638 -1844 -3414
rect 6244 -3638 6248 -3414
rect 6248 -3638 6784 -3414
rect 6784 -3638 6788 -3414
<< metal4 >>
rect -2600 2518 7000 2740
rect -2600 2294 -2388 2518
rect -1844 2294 6244 2518
rect 6788 2294 7000 2518
rect -2600 2117 7000 2294
rect -2600 2053 -2276 2117
rect -2212 2053 -2196 2117
rect -2132 2053 -2116 2117
rect -2052 2053 -2036 2117
rect -1972 2053 -1956 2117
rect -1892 2053 -1876 2117
rect -1812 2053 -1796 2117
rect -1732 2053 -1716 2117
rect -1652 2053 -1636 2117
rect -1572 2053 -1556 2117
rect -1492 2053 -1476 2117
rect -1412 2053 -1396 2117
rect -1332 2053 -1316 2117
rect -1252 2053 -1236 2117
rect -1172 2053 -1156 2117
rect -1092 2053 -1076 2117
rect -1012 2053 -996 2117
rect -932 2053 -916 2117
rect -852 2053 -836 2117
rect -772 2053 -756 2117
rect -692 2053 -676 2117
rect -612 2053 -596 2117
rect -532 2053 -516 2117
rect -452 2053 -436 2117
rect -372 2053 -356 2117
rect -292 2053 -276 2117
rect -212 2053 -196 2117
rect -132 2053 -116 2117
rect -52 2053 -36 2117
rect 28 2053 44 2117
rect 108 2053 124 2117
rect 188 2053 204 2117
rect 268 2053 284 2117
rect 348 2053 364 2117
rect 428 2053 444 2117
rect 508 2053 524 2117
rect 588 2053 604 2117
rect 668 2053 684 2117
rect 748 2053 764 2117
rect 828 2053 844 2117
rect 908 2053 924 2117
rect 988 2053 1004 2117
rect 1068 2053 1084 2117
rect 1148 2053 1164 2117
rect 1228 2053 1244 2117
rect 1308 2053 1324 2117
rect 1388 2053 1404 2117
rect 1468 2053 1484 2117
rect 1548 2053 1564 2117
rect 1628 2053 1644 2117
rect 1708 2053 1724 2117
rect 1788 2053 1804 2117
rect 1868 2053 1884 2117
rect 1948 2053 1964 2117
rect 2028 2053 2044 2117
rect 2108 2053 2124 2117
rect 2188 2053 2204 2117
rect 2268 2053 2284 2117
rect 2348 2053 2364 2117
rect 2428 2053 2444 2117
rect 2508 2053 2524 2117
rect 2588 2053 2604 2117
rect 2668 2053 2684 2117
rect 2748 2053 2764 2117
rect 2828 2053 2844 2117
rect 2908 2053 2924 2117
rect 2988 2053 3004 2117
rect 3068 2053 3084 2117
rect 3148 2053 3164 2117
rect 3228 2053 3244 2117
rect 3308 2053 3324 2117
rect 3388 2053 3404 2117
rect 3468 2053 3484 2117
rect 3548 2053 3564 2117
rect 3628 2053 3644 2117
rect 3708 2053 3724 2117
rect 3788 2053 3804 2117
rect 3868 2053 3884 2117
rect 3948 2053 3964 2117
rect 4028 2053 4044 2117
rect 4108 2053 4124 2117
rect 4188 2053 4204 2117
rect 4268 2053 4284 2117
rect 4348 2053 4364 2117
rect 4428 2053 4444 2117
rect 4508 2053 4524 2117
rect 4588 2053 4604 2117
rect 4668 2053 4684 2117
rect 4748 2053 4764 2117
rect 4828 2053 4844 2117
rect 4908 2053 4924 2117
rect 4988 2053 5004 2117
rect 5068 2053 5084 2117
rect 5148 2053 5164 2117
rect 5228 2053 5244 2117
rect 5308 2053 5324 2117
rect 5388 2053 5404 2117
rect 5468 2053 5484 2117
rect 5548 2053 5564 2117
rect 5628 2053 5644 2117
rect 5708 2053 5724 2117
rect 5788 2053 5804 2117
rect 5868 2053 5884 2117
rect 5948 2053 5964 2117
rect 6028 2053 6044 2117
rect 6108 2053 6124 2117
rect 6188 2053 6204 2117
rect 6268 2053 6284 2117
rect 6348 2053 6364 2117
rect 6428 2053 6444 2117
rect 6508 2053 6524 2117
rect 6588 2053 6604 2117
rect 6668 2053 7000 2117
rect -2600 1940 7000 2053
rect -2600 -3122 7000 -3060
rect -2600 -3266 -1763 -3122
rect 6061 -3266 7000 -3122
rect -2600 -3414 7000 -3266
rect -2600 -3638 -2388 -3414
rect -1844 -3638 6244 -3414
rect 6788 -3638 7000 -3414
rect -2600 -3860 7000 -3638
use sky130_fd_pr__nfet_01v8_58Q5WU  sky130_fd_pr__nfet_01v8_58Q5WU_0
timestamp 1626486988
transform 1 0 2128 0 1 -2666
box -3916 -188 3916 188
use sky130_fd_pr__nfet_01v8_58Q5WU  sky130_fd_pr__nfet_01v8_58Q5WU_1
timestamp 1626486988
transform 1 0 2128 0 1 -2084
box -3916 -188 3916 188
use sky130_fd_pr__nfet_01v8_N6QVV6  sky130_fd_pr__nfet_01v8_N6QVV6_0
timestamp 1626486988
transform 1 0 4180 0 1 -1031
box -931 -300 931 300
use sky130_fd_pr__nfet_01v8_lvt_V7QMZR  sky130_fd_pr__nfet_01v8_lvt_V7QMZR_0
timestamp 1626486988
transform 1 0 5689 0 1 -1031
box -544 -300 544 300
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1626486988
transform -1 0 880 0 1 -924
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1626486988
transform 1 0 52 0 1 -924
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0
timestamp 1626486988
transform -1 0 604 0 1 -924
box -38 -48 314 592
use sky130_fd_pr__pfet_01v8_SCHXZ7  sky130_fd_pr__pfet_01v8_SCHXZ7_0
timestamp 1626486988
transform 1 0 4180 0 1 -244
box -941 -419 941 419
use sky130_fd_pr__pfet_01v8_lvt_HJ2CZP  sky130_fd_pr__pfet_01v8_lvt_HJ2CZP_0
timestamp 1626486988
transform 1 0 5689 0 1 -244
box -554 -419 554 419
use sky130_fd_sc_hd__dfrbp_1  sky130_fd_sc_hd__dfrbp_1_0
timestamp 1626486988
transform 1 0 -2064 0 1 -924
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  sky130_fd_sc_hd__dfrbp_1_1
timestamp 1626486988
transform -1 0 2996 0 1 -924
box -38 -48 2154 592
use sky130_fd_pr__pfet_01v8_2Q5KMA  sky130_fd_pr__pfet_01v8_2Q5KMA_0
timestamp 1626486988
transform 1 0 2173 0 1 1496
box -4355 -200 4355 200
use sky130_fd_pr__pfet_01v8_2Q5KMA  sky130_fd_pr__pfet_01v8_2Q5KMA_1
timestamp 1626486988
transform 1 0 2173 0 1 896
box -4355 -200 4355 200
<< labels >>
flabel metal1 s 2548 -1880 2560 -1874 1 FreeSans 600 0 0 0 vswitchl
flabel metal2 s 1694 -2378 1704 -2366 1 FreeSans 600 0 0 0 ibiasn
flabel metal1 s 3656 -862 3666 -854 1 FreeSans 600 0 0 0 vpdiode
flabel metal1 s 5552 -1226 5564 -1208 1 FreeSans 600 0 0 0 vswitchl
flabel metal2 s 4962 114 4976 132 1 FreeSans 600 0 0 0 vswitchh
flabel metal2 s 1104 596 1120 610 1 FreeSans 600 0 0 0 vswitchh
flabel metal1 s 5812 -840 5822 -830 1 FreeSans 600 0 0 0 vcp
flabel metal1 s 620 -692 624 -688 1 FreeSans 600 0 0 0 vQB
flabel metal1 s 294 -700 300 -692 1 FreeSans 600 0 0 0 vQA
flabel metal1 s -2200 -692 -2194 -688 1 FreeSans 600 0 0 0 vsig_in
flabel metal1 s 3070 -680 3078 -676 1 FreeSans 600 0 0 0 vin_div
flabel metal1 s 300 -592 304 -588 1 FreeSans 600 0 0 0 vRSTN
flabel metal2 s 944 -1420 952 -1412 1 FreeSans 600 0 0 0 VQBb
flabel metal2 s 220 -146 228 -138 1 FreeSans 600 0 0 0 vQAb
flabel metal2 s 1582 1194 1598 1204 1 FreeSans 600 0 0 0 vpbias
flabel metal2 s 2204 -2944 2214 -2936 1 FreeSans 600 0 0 0 vpbias
flabel metal4 s 886 2206 898 2222 1 FreeSans 600 0 0 0 VDD
flabel metal4 s 1252 -3422 1278 -3396 1 FreeSans 600 0 0 0 VSS
flabel metal1 s 4436 -580 4442 -570 1 FreeSans 600 0 0 0 vndiode
<< properties >>
string FIXED_BBOX -2472 -3732 6872 -1668
<< end >>
