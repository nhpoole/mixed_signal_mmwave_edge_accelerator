magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< metal2 >>
rect 0 101759 28 101807
rect 0 101539 28 101587
rect 0 101443 28 101491
rect 0 101223 28 101271
rect 0 100969 28 101017
rect 0 100749 28 100797
rect 0 100653 28 100701
rect 0 100433 28 100481
rect 0 100179 28 100227
rect 0 99959 28 100007
rect 0 99863 28 99911
rect 0 99643 28 99691
rect 0 99389 28 99437
rect 0 99169 28 99217
rect 0 99073 28 99121
rect 0 98853 28 98901
rect 0 98599 28 98647
rect 0 98379 28 98427
rect 0 98283 28 98331
rect 0 98063 28 98111
rect 0 97809 28 97857
rect 0 97589 28 97637
rect 0 97493 28 97541
rect 0 97273 28 97321
rect 0 97019 28 97067
rect 0 96799 28 96847
rect 0 96703 28 96751
rect 0 96483 28 96531
rect 0 96229 28 96277
rect 0 96009 28 96057
rect 0 95913 28 95961
rect 0 95693 28 95741
rect 0 95439 28 95487
rect 0 95219 28 95267
rect 0 95123 28 95171
rect 0 94903 28 94951
rect 0 94649 28 94697
rect 0 94429 28 94477
rect 0 94333 28 94381
rect 0 94113 28 94161
rect 0 93859 28 93907
rect 0 93639 28 93687
rect 0 93543 28 93591
rect 0 93323 28 93371
rect 0 93069 28 93117
rect 0 92849 28 92897
rect 0 92753 28 92801
rect 0 92533 28 92581
rect 0 92279 28 92327
rect 0 92059 28 92107
rect 0 91963 28 92011
rect 0 91743 28 91791
rect 0 91489 28 91537
rect 0 91269 28 91317
rect 0 91173 28 91221
rect 0 90953 28 91001
rect 0 90699 28 90747
rect 0 90479 28 90527
rect 0 90383 28 90431
rect 0 90163 28 90211
rect 0 89909 28 89957
rect 0 89689 28 89737
rect 0 89593 28 89641
rect 0 89373 28 89421
rect 0 89119 28 89167
rect 0 88899 28 88947
rect 0 88803 28 88851
rect 0 88583 28 88631
rect 0 88329 28 88377
rect 0 88109 28 88157
rect 0 88013 28 88061
rect 0 87793 28 87841
rect 0 87539 28 87587
rect 0 87319 28 87367
rect 0 87223 28 87271
rect 0 87003 28 87051
rect 0 86749 28 86797
rect 0 86529 28 86577
rect 0 86433 28 86481
rect 0 86213 28 86261
rect 0 85959 28 86007
rect 0 85739 28 85787
rect 0 85643 28 85691
rect 0 85423 28 85471
rect 0 85169 28 85217
rect 0 84949 28 84997
rect 0 84853 28 84901
rect 0 84633 28 84681
rect 0 84379 28 84427
rect 0 84159 28 84207
rect 0 84063 28 84111
rect 0 83843 28 83891
rect 0 83589 28 83637
rect 0 83369 28 83417
rect 0 83273 28 83321
rect 0 83053 28 83101
rect 0 82799 28 82847
rect 0 82579 28 82627
rect 0 82483 28 82531
rect 0 82263 28 82311
rect 0 82009 28 82057
rect 0 81789 28 81837
rect 0 81693 28 81741
rect 0 81473 28 81521
rect 0 81219 28 81267
rect 0 80999 28 81047
rect 0 80903 28 80951
rect 0 80683 28 80731
rect 0 80429 28 80477
rect 0 80209 28 80257
rect 0 80113 28 80161
rect 0 79893 28 79941
rect 0 79639 28 79687
rect 0 79419 28 79467
rect 0 79323 28 79371
rect 0 79103 28 79151
rect 0 78849 28 78897
rect 0 78629 28 78677
rect 0 78533 28 78581
rect 0 78313 28 78361
rect 0 78059 28 78107
rect 0 77839 28 77887
rect 0 77743 28 77791
rect 0 77523 28 77571
rect 0 77269 28 77317
rect 0 77049 28 77097
rect 0 76953 28 77001
rect 0 76733 28 76781
rect 0 76479 28 76527
rect 0 76259 28 76307
rect 0 76163 28 76211
rect 0 75943 28 75991
rect 0 75689 28 75737
rect 0 75469 28 75517
rect 0 75373 28 75421
rect 0 75153 28 75201
rect 0 74899 28 74947
rect 0 74679 28 74727
rect 0 74583 28 74631
rect 0 74363 28 74411
rect 0 74109 28 74157
rect 0 73889 28 73937
rect 0 73793 28 73841
rect 0 73573 28 73621
rect 0 73319 28 73367
rect 0 73099 28 73147
rect 0 73003 28 73051
rect 0 72783 28 72831
rect 0 72529 28 72577
rect 0 72309 28 72357
rect 0 72213 28 72261
rect 0 71993 28 72041
rect 0 71739 28 71787
rect 0 71519 28 71567
rect 0 71423 28 71471
rect 0 71203 28 71251
rect 0 70949 28 70997
rect 0 70729 28 70777
rect 0 70633 28 70681
rect 0 70413 28 70461
rect 0 70159 28 70207
rect 0 69939 28 69987
rect 0 69843 28 69891
rect 0 69623 28 69671
rect 0 69369 28 69417
rect 0 69149 28 69197
rect 0 69053 28 69101
rect 0 68833 28 68881
rect 0 68579 28 68627
rect 0 68359 28 68407
rect 0 68263 28 68311
rect 0 68043 28 68091
rect 0 67789 28 67837
rect 0 67569 28 67617
rect 0 67473 28 67521
rect 0 67253 28 67301
rect 0 66999 28 67047
rect 0 66779 28 66827
rect 0 66683 28 66731
rect 0 66463 28 66511
rect 0 66209 28 66257
rect 0 65989 28 66037
rect 0 65893 28 65941
rect 0 65673 28 65721
rect 0 65419 28 65467
rect 0 65199 28 65247
rect 0 65103 28 65151
rect 0 64883 28 64931
rect 0 64629 28 64677
rect 0 64409 28 64457
rect 0 64313 28 64361
rect 0 64093 28 64141
rect 0 63839 28 63887
rect 0 63619 28 63667
rect 0 63523 28 63571
rect 0 63303 28 63351
rect 0 63049 28 63097
rect 0 62829 28 62877
rect 0 62733 28 62781
rect 0 62513 28 62561
rect 0 62259 28 62307
rect 0 62039 28 62087
rect 0 61943 28 61991
rect 0 61723 28 61771
rect 0 61469 28 61517
rect 0 61249 28 61297
rect 0 61153 28 61201
rect 0 60933 28 60981
rect 0 60679 28 60727
rect 0 60459 28 60507
rect 0 60363 28 60411
rect 0 60143 28 60191
rect 0 59889 28 59937
rect 0 59669 28 59717
rect 0 59573 28 59621
rect 0 59353 28 59401
rect 0 59099 28 59147
rect 0 58879 28 58927
rect 0 58783 28 58831
rect 0 58563 28 58611
rect 0 58309 28 58357
rect 0 58089 28 58137
rect 0 57993 28 58041
rect 0 57773 28 57821
rect 0 57519 28 57567
rect 0 57299 28 57347
rect 0 57203 28 57251
rect 0 56983 28 57031
rect 0 56729 28 56777
rect 0 56509 28 56557
rect 0 56413 28 56461
rect 0 56193 28 56241
rect 0 55939 28 55987
rect 0 55719 28 55767
rect 0 55623 28 55671
rect 0 55403 28 55451
rect 0 55149 28 55197
rect 0 54929 28 54977
rect 0 54833 28 54881
rect 0 54613 28 54661
rect 0 54359 28 54407
rect 0 54139 28 54187
rect 0 54043 28 54091
rect 0 53823 28 53871
rect 0 53569 28 53617
rect 0 53349 28 53397
rect 0 53253 28 53301
rect 0 53033 28 53081
rect 0 52779 28 52827
rect 0 52559 28 52607
rect 0 52463 28 52511
rect 0 52243 28 52291
rect 0 51989 28 52037
rect 0 51769 28 51817
rect 0 51673 28 51721
rect 0 51453 28 51501
rect 0 51199 28 51247
rect 0 50979 28 51027
rect 0 50883 28 50931
rect 0 50663 28 50711
rect 0 50409 28 50457
rect 0 50189 28 50237
rect 0 50093 28 50141
rect 0 49873 28 49921
rect 0 49619 28 49667
rect 0 49399 28 49447
rect 0 49303 28 49351
rect 0 49083 28 49131
rect 0 48829 28 48877
rect 0 48609 28 48657
rect 0 48513 28 48561
rect 0 48293 28 48341
rect 0 48039 28 48087
rect 0 47819 28 47867
rect 0 47723 28 47771
rect 0 47503 28 47551
rect 0 47249 28 47297
rect 0 47029 28 47077
rect 0 46933 28 46981
rect 0 46713 28 46761
rect 0 46459 28 46507
rect 0 46239 28 46287
rect 0 46143 28 46191
rect 0 45923 28 45971
rect 0 45669 28 45717
rect 0 45449 28 45497
rect 0 45353 28 45401
rect 0 45133 28 45181
rect 0 44879 28 44927
rect 0 44659 28 44707
rect 0 44563 28 44611
rect 0 44343 28 44391
rect 0 44089 28 44137
rect 0 43869 28 43917
rect 0 43773 28 43821
rect 0 43553 28 43601
rect 0 43299 28 43347
rect 0 43079 28 43127
rect 0 42983 28 43031
rect 0 42763 28 42811
rect 0 42509 28 42557
rect 0 42289 28 42337
rect 0 42193 28 42241
rect 0 41973 28 42021
rect 0 41719 28 41767
rect 0 41499 28 41547
rect 0 41403 28 41451
rect 0 41183 28 41231
rect 0 40929 28 40977
rect 0 40709 28 40757
rect 0 40613 28 40661
rect 0 40393 28 40441
rect 0 40139 28 40187
rect 0 39919 28 39967
rect 0 39823 28 39871
rect 0 39603 28 39651
rect 0 39349 28 39397
rect 0 39129 28 39177
rect 0 39033 28 39081
rect 0 38813 28 38861
rect 0 38559 28 38607
rect 0 38339 28 38387
rect 0 38243 28 38291
rect 0 38023 28 38071
rect 0 37769 28 37817
rect 0 37549 28 37597
rect 0 37453 28 37501
rect 0 37233 28 37281
rect 0 36979 28 37027
rect 0 36759 28 36807
rect 0 36663 28 36711
rect 0 36443 28 36491
rect 0 36189 28 36237
rect 0 35969 28 36017
rect 0 35873 28 35921
rect 0 35653 28 35701
rect 0 35399 28 35447
rect 0 35179 28 35227
rect 0 35083 28 35131
rect 0 34863 28 34911
rect 0 34609 28 34657
rect 0 34389 28 34437
rect 0 34293 28 34341
rect 0 34073 28 34121
rect 0 33819 28 33867
rect 0 33599 28 33647
rect 0 33503 28 33551
rect 0 33283 28 33331
rect 0 33029 28 33077
rect 0 32809 28 32857
rect 0 32713 28 32761
rect 0 32493 28 32541
rect 0 32239 28 32287
rect 0 32019 28 32067
rect 0 31923 28 31971
rect 0 31703 28 31751
rect 0 31449 28 31497
rect 0 31229 28 31277
rect 0 31133 28 31181
rect 0 30913 28 30961
rect 0 30659 28 30707
rect 0 30439 28 30487
rect 0 30343 28 30391
rect 0 30123 28 30171
rect 0 29869 28 29917
rect 0 29649 28 29697
rect 0 29553 28 29601
rect 0 29333 28 29381
rect 0 29079 28 29127
rect 0 28859 28 28907
rect 0 28763 28 28811
rect 0 28543 28 28591
rect 0 28289 28 28337
rect 0 28069 28 28117
rect 0 27973 28 28021
rect 0 27753 28 27801
rect 0 27499 28 27547
rect 0 27279 28 27327
rect 0 27183 28 27231
rect 0 26963 28 27011
rect 0 26709 28 26757
rect 0 26489 28 26537
rect 0 26393 28 26441
rect 0 26173 28 26221
rect 0 25919 28 25967
rect 0 25699 28 25747
rect 0 25603 28 25651
rect 0 25383 28 25431
rect 0 25129 28 25177
rect 0 24909 28 24957
rect 0 24813 28 24861
rect 0 24593 28 24641
rect 0 24339 28 24387
rect 0 24119 28 24167
rect 0 24023 28 24071
rect 0 23803 28 23851
rect 0 23549 28 23597
rect 0 23329 28 23377
rect 0 23233 28 23281
rect 0 23013 28 23061
rect 0 22759 28 22807
rect 0 22539 28 22587
rect 0 22443 28 22491
rect 0 22223 28 22271
rect 0 21969 28 22017
rect 0 21749 28 21797
rect 0 21653 28 21701
rect 0 21433 28 21481
rect 0 21179 28 21227
rect 0 20959 28 21007
rect 0 20863 28 20911
rect 0 20643 28 20691
rect 0 20389 28 20437
rect 0 20169 28 20217
rect 0 20073 28 20121
rect 0 19853 28 19901
rect 0 19599 28 19647
rect 0 19379 28 19427
rect 0 19283 28 19331
rect 0 19063 28 19111
rect 0 18809 28 18857
rect 0 18589 28 18637
rect 0 18493 28 18541
rect 0 18273 28 18321
rect 0 18019 28 18067
rect 0 17799 28 17847
rect 0 17703 28 17751
rect 0 17483 28 17531
rect 0 17229 28 17277
rect 0 17009 28 17057
rect 0 16913 28 16961
rect 0 16693 28 16741
rect 0 16439 28 16487
rect 0 16219 28 16267
rect 0 16123 28 16171
rect 0 15903 28 15951
rect 0 15649 28 15697
rect 0 15429 28 15477
rect 0 15333 28 15381
rect 0 15113 28 15161
rect 0 14859 28 14907
rect 0 14639 28 14687
rect 0 14543 28 14591
rect 0 14323 28 14371
rect 0 14069 28 14117
rect 0 13849 28 13897
rect 0 13753 28 13801
rect 0 13533 28 13581
rect 0 13279 28 13327
rect 0 13059 28 13107
rect 0 12963 28 13011
rect 0 12743 28 12791
rect 0 12489 28 12537
rect 0 12269 28 12317
rect 0 12173 28 12221
rect 0 11953 28 12001
rect 0 11699 28 11747
rect 0 11479 28 11527
rect 0 11383 28 11431
rect 0 11163 28 11211
rect 0 10909 28 10957
rect 0 10689 28 10737
rect 0 10593 28 10641
rect 0 10373 28 10421
rect 0 10119 28 10167
rect 0 9899 28 9947
rect 0 9803 28 9851
rect 0 9583 28 9631
rect 0 9329 28 9377
rect 0 9109 28 9157
rect 0 9013 28 9061
rect 0 8793 28 8841
rect 0 8539 28 8587
rect 0 8319 28 8367
rect 0 8223 28 8271
rect 0 8003 28 8051
rect 0 7749 28 7797
rect 0 7529 28 7577
rect 0 7433 28 7481
rect 0 7213 28 7261
rect 0 6959 28 7007
rect 0 6739 28 6787
rect 0 6643 28 6691
rect 0 6423 28 6471
rect 0 6169 28 6217
rect 0 5949 28 5997
rect 0 5853 28 5901
rect 0 5633 28 5681
rect 0 5379 28 5427
rect 0 5159 28 5207
rect 0 5063 28 5111
rect 0 4843 28 4891
rect 0 4589 28 4637
rect 0 4369 28 4417
rect 0 4273 28 4321
rect 0 4053 28 4101
rect 0 3799 28 3847
rect 0 3579 28 3627
rect 0 3483 28 3531
rect 0 3263 28 3311
rect 0 3009 28 3057
rect 0 2789 28 2837
rect 0 2693 28 2741
rect 0 2473 28 2521
rect 0 2219 28 2267
rect 0 1999 28 2047
rect 0 1903 28 1951
rect 0 1683 28 1731
rect 0 1429 28 1477
rect 0 1209 28 1257
rect 0 1113 28 1161
rect 0 893 28 941
<< metal3 >>
rect 335 101861 433 101959
rect 335 101624 433 101722
rect 335 101308 433 101406
rect 335 101071 433 101169
rect 335 100834 433 100932
rect 335 100518 433 100616
rect 335 100281 433 100379
rect 335 100044 433 100142
rect 335 99728 433 99826
rect 335 99491 433 99589
rect 335 99254 433 99352
rect 335 98938 433 99036
rect 335 98701 433 98799
rect 335 98464 433 98562
rect 335 98148 433 98246
rect 335 97911 433 98009
rect 335 97674 433 97772
rect 335 97358 433 97456
rect 335 97121 433 97219
rect 335 96884 433 96982
rect 335 96568 433 96666
rect 335 96331 433 96429
rect 335 96094 433 96192
rect 335 95778 433 95876
rect 335 95541 433 95639
rect 335 95304 433 95402
rect 335 94988 433 95086
rect 335 94751 433 94849
rect 335 94514 433 94612
rect 335 94198 433 94296
rect 335 93961 433 94059
rect 335 93724 433 93822
rect 335 93408 433 93506
rect 335 93171 433 93269
rect 335 92934 433 93032
rect 335 92618 433 92716
rect 335 92381 433 92479
rect 335 92144 433 92242
rect 335 91828 433 91926
rect 335 91591 433 91689
rect 335 91354 433 91452
rect 335 91038 433 91136
rect 335 90801 433 90899
rect 335 90564 433 90662
rect 335 90248 433 90346
rect 335 90011 433 90109
rect 335 89774 433 89872
rect 335 89458 433 89556
rect 335 89221 433 89319
rect 335 88984 433 89082
rect 335 88668 433 88766
rect 335 88431 433 88529
rect 335 88194 433 88292
rect 335 87878 433 87976
rect 335 87641 433 87739
rect 335 87404 433 87502
rect 335 87088 433 87186
rect 335 86851 433 86949
rect 335 86614 433 86712
rect 335 86298 433 86396
rect 335 86061 433 86159
rect 335 85824 433 85922
rect 335 85508 433 85606
rect 335 85271 433 85369
rect 335 85034 433 85132
rect 335 84718 433 84816
rect 335 84481 433 84579
rect 335 84244 433 84342
rect 335 83928 433 84026
rect 335 83691 433 83789
rect 335 83454 433 83552
rect 335 83138 433 83236
rect 335 82901 433 82999
rect 335 82664 433 82762
rect 335 82348 433 82446
rect 335 82111 433 82209
rect 335 81874 433 81972
rect 335 81558 433 81656
rect 335 81321 433 81419
rect 335 81084 433 81182
rect 335 80768 433 80866
rect 335 80531 433 80629
rect 335 80294 433 80392
rect 335 79978 433 80076
rect 335 79741 433 79839
rect 335 79504 433 79602
rect 335 79188 433 79286
rect 335 78951 433 79049
rect 335 78714 433 78812
rect 335 78398 433 78496
rect 335 78161 433 78259
rect 335 77924 433 78022
rect 335 77608 433 77706
rect 335 77371 433 77469
rect 335 77134 433 77232
rect 335 76818 433 76916
rect 335 76581 433 76679
rect 335 76344 433 76442
rect 335 76028 433 76126
rect 335 75791 433 75889
rect 335 75554 433 75652
rect 335 75238 433 75336
rect 335 75001 433 75099
rect 335 74764 433 74862
rect 335 74448 433 74546
rect 335 74211 433 74309
rect 335 73974 433 74072
rect 335 73658 433 73756
rect 335 73421 433 73519
rect 335 73184 433 73282
rect 335 72868 433 72966
rect 335 72631 433 72729
rect 335 72394 433 72492
rect 335 72078 433 72176
rect 335 71841 433 71939
rect 335 71604 433 71702
rect 335 71288 433 71386
rect 335 71051 433 71149
rect 335 70814 433 70912
rect 335 70498 433 70596
rect 335 70261 433 70359
rect 335 70024 433 70122
rect 335 69708 433 69806
rect 335 69471 433 69569
rect 335 69234 433 69332
rect 335 68918 433 69016
rect 335 68681 433 68779
rect 335 68444 433 68542
rect 335 68128 433 68226
rect 335 67891 433 67989
rect 335 67654 433 67752
rect 335 67338 433 67436
rect 335 67101 433 67199
rect 335 66864 433 66962
rect 335 66548 433 66646
rect 335 66311 433 66409
rect 335 66074 433 66172
rect 335 65758 433 65856
rect 335 65521 433 65619
rect 335 65284 433 65382
rect 335 64968 433 65066
rect 335 64731 433 64829
rect 335 64494 433 64592
rect 335 64178 433 64276
rect 335 63941 433 64039
rect 335 63704 433 63802
rect 335 63388 433 63486
rect 335 63151 433 63249
rect 335 62914 433 63012
rect 335 62598 433 62696
rect 335 62361 433 62459
rect 335 62124 433 62222
rect 335 61808 433 61906
rect 335 61571 433 61669
rect 335 61334 433 61432
rect 335 61018 433 61116
rect 335 60781 433 60879
rect 335 60544 433 60642
rect 335 60228 433 60326
rect 335 59991 433 60089
rect 335 59754 433 59852
rect 335 59438 433 59536
rect 335 59201 433 59299
rect 335 58964 433 59062
rect 335 58648 433 58746
rect 335 58411 433 58509
rect 335 58174 433 58272
rect 335 57858 433 57956
rect 335 57621 433 57719
rect 335 57384 433 57482
rect 335 57068 433 57166
rect 335 56831 433 56929
rect 335 56594 433 56692
rect 335 56278 433 56376
rect 335 56041 433 56139
rect 335 55804 433 55902
rect 335 55488 433 55586
rect 335 55251 433 55349
rect 335 55014 433 55112
rect 335 54698 433 54796
rect 335 54461 433 54559
rect 335 54224 433 54322
rect 335 53908 433 54006
rect 335 53671 433 53769
rect 335 53434 433 53532
rect 335 53118 433 53216
rect 335 52881 433 52979
rect 335 52644 433 52742
rect 335 52328 433 52426
rect 335 52091 433 52189
rect 335 51854 433 51952
rect 335 51538 433 51636
rect 335 51301 433 51399
rect 335 51064 433 51162
rect 335 50748 433 50846
rect 335 50511 433 50609
rect 335 50274 433 50372
rect 335 49958 433 50056
rect 335 49721 433 49819
rect 335 49484 433 49582
rect 335 49168 433 49266
rect 335 48931 433 49029
rect 335 48694 433 48792
rect 335 48378 433 48476
rect 335 48141 433 48239
rect 335 47904 433 48002
rect 335 47588 433 47686
rect 335 47351 433 47449
rect 335 47114 433 47212
rect 335 46798 433 46896
rect 335 46561 433 46659
rect 335 46324 433 46422
rect 335 46008 433 46106
rect 335 45771 433 45869
rect 335 45534 433 45632
rect 335 45218 433 45316
rect 335 44981 433 45079
rect 335 44744 433 44842
rect 335 44428 433 44526
rect 335 44191 433 44289
rect 335 43954 433 44052
rect 335 43638 433 43736
rect 335 43401 433 43499
rect 335 43164 433 43262
rect 335 42848 433 42946
rect 335 42611 433 42709
rect 335 42374 433 42472
rect 335 42058 433 42156
rect 335 41821 433 41919
rect 335 41584 433 41682
rect 335 41268 433 41366
rect 335 41031 433 41129
rect 335 40794 433 40892
rect 335 40478 433 40576
rect 335 40241 433 40339
rect 335 40004 433 40102
rect 335 39688 433 39786
rect 335 39451 433 39549
rect 335 39214 433 39312
rect 335 38898 433 38996
rect 335 38661 433 38759
rect 335 38424 433 38522
rect 335 38108 433 38206
rect 335 37871 433 37969
rect 335 37634 433 37732
rect 335 37318 433 37416
rect 335 37081 433 37179
rect 335 36844 433 36942
rect 335 36528 433 36626
rect 335 36291 433 36389
rect 335 36054 433 36152
rect 335 35738 433 35836
rect 335 35501 433 35599
rect 335 35264 433 35362
rect 335 34948 433 35046
rect 335 34711 433 34809
rect 335 34474 433 34572
rect 335 34158 433 34256
rect 335 33921 433 34019
rect 335 33684 433 33782
rect 335 33368 433 33466
rect 335 33131 433 33229
rect 335 32894 433 32992
rect 335 32578 433 32676
rect 335 32341 433 32439
rect 335 32104 433 32202
rect 335 31788 433 31886
rect 335 31551 433 31649
rect 335 31314 433 31412
rect 335 30998 433 31096
rect 335 30761 433 30859
rect 335 30524 433 30622
rect 335 30208 433 30306
rect 335 29971 433 30069
rect 335 29734 433 29832
rect 335 29418 433 29516
rect 335 29181 433 29279
rect 335 28944 433 29042
rect 335 28628 433 28726
rect 335 28391 433 28489
rect 335 28154 433 28252
rect 335 27838 433 27936
rect 335 27601 433 27699
rect 335 27364 433 27462
rect 335 27048 433 27146
rect 335 26811 433 26909
rect 335 26574 433 26672
rect 335 26258 433 26356
rect 335 26021 433 26119
rect 335 25784 433 25882
rect 335 25468 433 25566
rect 335 25231 433 25329
rect 335 24994 433 25092
rect 335 24678 433 24776
rect 335 24441 433 24539
rect 335 24204 433 24302
rect 335 23888 433 23986
rect 335 23651 433 23749
rect 335 23414 433 23512
rect 335 23098 433 23196
rect 335 22861 433 22959
rect 335 22624 433 22722
rect 335 22308 433 22406
rect 335 22071 433 22169
rect 335 21834 433 21932
rect 335 21518 433 21616
rect 335 21281 433 21379
rect 335 21044 433 21142
rect 335 20728 433 20826
rect 335 20491 433 20589
rect 335 20254 433 20352
rect 335 19938 433 20036
rect 335 19701 433 19799
rect 335 19464 433 19562
rect 335 19148 433 19246
rect 335 18911 433 19009
rect 335 18674 433 18772
rect 335 18358 433 18456
rect 335 18121 433 18219
rect 335 17884 433 17982
rect 335 17568 433 17666
rect 335 17331 433 17429
rect 335 17094 433 17192
rect 335 16778 433 16876
rect 335 16541 433 16639
rect 335 16304 433 16402
rect 335 15988 433 16086
rect 335 15751 433 15849
rect 335 15514 433 15612
rect 335 15198 433 15296
rect 335 14961 433 15059
rect 335 14724 433 14822
rect 335 14408 433 14506
rect 335 14171 433 14269
rect 335 13934 433 14032
rect 335 13618 433 13716
rect 335 13381 433 13479
rect 335 13144 433 13242
rect 335 12828 433 12926
rect 335 12591 433 12689
rect 335 12354 433 12452
rect 335 12038 433 12136
rect 335 11801 433 11899
rect 335 11564 433 11662
rect 335 11248 433 11346
rect 335 11011 433 11109
rect 335 10774 433 10872
rect 335 10458 433 10556
rect 335 10221 433 10319
rect 335 9984 433 10082
rect 335 9668 433 9766
rect 335 9431 433 9529
rect 335 9194 433 9292
rect 335 8878 433 8976
rect 335 8641 433 8739
rect 335 8404 433 8502
rect 335 8088 433 8186
rect 335 7851 433 7949
rect 335 7614 433 7712
rect 335 7298 433 7396
rect 335 7061 433 7159
rect 335 6824 433 6922
rect 335 6508 433 6606
rect 335 6271 433 6369
rect 335 6034 433 6132
rect 335 5718 433 5816
rect 335 5481 433 5579
rect 335 5244 433 5342
rect 335 4928 433 5026
rect 335 4691 433 4789
rect 335 4454 433 4552
rect 335 4138 433 4236
rect 335 3901 433 3999
rect 335 3664 433 3762
rect 335 3348 433 3446
rect 335 3111 433 3209
rect 335 2874 433 2972
rect 335 2558 433 2656
rect 335 2321 433 2419
rect 335 2084 433 2182
rect 335 1768 433 1866
rect 335 1531 433 1629
rect 335 1294 433 1392
rect 335 978 433 1076
rect 335 741 433 839
use contact_9  contact_9_510
timestamp 1624494425
transform 1 0 351 0 1 753
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_256
timestamp 1624494425
transform -1 0 624 0 1 790
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_257
timestamp 1624494425
transform -1 0 624 0 -1 790
box -42 -55 624 371
use contact_9  contact_9_511
timestamp 1624494425
transform 1 0 351 0 1 990
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_255
timestamp 1624494425
transform -1 0 624 0 -1 1580
box -42 -55 624 371
use contact_9  contact_9_509
timestamp 1624494425
transform 1 0 351 0 1 1306
box 0 0 66 74
use contact_9  contact_9_508
timestamp 1624494425
transform 1 0 351 0 1 1543
box 0 0 66 74
use contact_9  contact_9_506
timestamp 1624494425
transform 1 0 351 0 1 1543
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_254
timestamp 1624494425
transform -1 0 624 0 1 1580
box -42 -55 624 371
use contact_9  contact_9_507
timestamp 1624494425
transform 1 0 351 0 1 1780
box 0 0 66 74
use contact_9  contact_9_505
timestamp 1624494425
transform 1 0 351 0 1 2096
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_253
timestamp 1624494425
transform -1 0 624 0 -1 2370
box -42 -55 624 371
use contact_9  contact_9_504
timestamp 1624494425
transform 1 0 351 0 1 2333
box 0 0 66 74
use contact_9  contact_9_502
timestamp 1624494425
transform 1 0 351 0 1 2333
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_252
timestamp 1624494425
transform -1 0 624 0 1 2370
box -42 -55 624 371
use contact_9  contact_9_503
timestamp 1624494425
transform 1 0 351 0 1 2570
box 0 0 66 74
use contact_9  contact_9_501
timestamp 1624494425
transform 1 0 351 0 1 2886
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_251
timestamp 1624494425
transform -1 0 624 0 -1 3160
box -42 -55 624 371
use contact_9  contact_9_500
timestamp 1624494425
transform 1 0 351 0 1 3123
box 0 0 66 74
use contact_9  contact_9_499
timestamp 1624494425
transform 1 0 351 0 1 3360
box 0 0 66 74
use contact_9  contact_9_498
timestamp 1624494425
transform 1 0 351 0 1 3123
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_250
timestamp 1624494425
transform -1 0 624 0 1 3160
box -42 -55 624 371
use contact_9  contact_9_497
timestamp 1624494425
transform 1 0 351 0 1 3676
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_249
timestamp 1624494425
transform -1 0 624 0 -1 3950
box -42 -55 624 371
use contact_9  contact_9_496
timestamp 1624494425
transform 1 0 351 0 1 3913
box 0 0 66 74
use contact_9  contact_9_495
timestamp 1624494425
transform 1 0 351 0 1 4150
box 0 0 66 74
use contact_9  contact_9_494
timestamp 1624494425
transform 1 0 351 0 1 3913
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_248
timestamp 1624494425
transform -1 0 624 0 1 3950
box -42 -55 624 371
use contact_9  contact_9_493
timestamp 1624494425
transform 1 0 351 0 1 4466
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_246
timestamp 1624494425
transform -1 0 624 0 1 4740
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_247
timestamp 1624494425
transform -1 0 624 0 -1 4740
box -42 -55 624 371
use contact_9  contact_9_492
timestamp 1624494425
transform 1 0 351 0 1 4703
box 0 0 66 74
use contact_9  contact_9_491
timestamp 1624494425
transform 1 0 351 0 1 4940
box 0 0 66 74
use contact_9  contact_9_490
timestamp 1624494425
transform 1 0 351 0 1 4703
box 0 0 66 74
use contact_9  contact_9_489
timestamp 1624494425
transform 1 0 351 0 1 5256
box 0 0 66 74
use contact_9  contact_9_488
timestamp 1624494425
transform 1 0 351 0 1 5493
box 0 0 66 74
use contact_9  contact_9_486
timestamp 1624494425
transform 1 0 351 0 1 5493
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_244
timestamp 1624494425
transform -1 0 624 0 1 5530
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_245
timestamp 1624494425
transform -1 0 624 0 -1 5530
box -42 -55 624 371
use contact_9  contact_9_487
timestamp 1624494425
transform 1 0 351 0 1 5730
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_243
timestamp 1624494425
transform -1 0 624 0 -1 6320
box -42 -55 624 371
use contact_9  contact_9_485
timestamp 1624494425
transform 1 0 351 0 1 6046
box 0 0 66 74
use contact_9  contact_9_484
timestamp 1624494425
transform 1 0 351 0 1 6283
box 0 0 66 74
use contact_9  contact_9_482
timestamp 1624494425
transform 1 0 351 0 1 6283
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_242
timestamp 1624494425
transform -1 0 624 0 1 6320
box -42 -55 624 371
use contact_9  contact_9_483
timestamp 1624494425
transform 1 0 351 0 1 6520
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_241
timestamp 1624494425
transform -1 0 624 0 -1 7110
box -42 -55 624 371
use contact_9  contact_9_481
timestamp 1624494425
transform 1 0 351 0 1 6836
box 0 0 66 74
use contact_9  contact_9_480
timestamp 1624494425
transform 1 0 351 0 1 7073
box 0 0 66 74
use contact_9  contact_9_478
timestamp 1624494425
transform 1 0 351 0 1 7073
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_240
timestamp 1624494425
transform -1 0 624 0 1 7110
box -42 -55 624 371
use contact_9  contact_9_479
timestamp 1624494425
transform 1 0 351 0 1 7310
box 0 0 66 74
use contact_9  contact_9_477
timestamp 1624494425
transform 1 0 351 0 1 7626
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_239
timestamp 1624494425
transform -1 0 624 0 -1 7900
box -42 -55 624 371
use contact_9  contact_9_476
timestamp 1624494425
transform 1 0 351 0 1 7863
box 0 0 66 74
use contact_9  contact_9_475
timestamp 1624494425
transform 1 0 351 0 1 8100
box 0 0 66 74
use contact_9  contact_9_474
timestamp 1624494425
transform 1 0 351 0 1 7863
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_238
timestamp 1624494425
transform -1 0 624 0 1 7900
box -42 -55 624 371
use contact_9  contact_9_473
timestamp 1624494425
transform 1 0 351 0 1 8416
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_237
timestamp 1624494425
transform -1 0 624 0 -1 8690
box -42 -55 624 371
use contact_9  contact_9_472
timestamp 1624494425
transform 1 0 351 0 1 8653
box 0 0 66 74
use contact_9  contact_9_471
timestamp 1624494425
transform 1 0 351 0 1 8890
box 0 0 66 74
use contact_9  contact_9_470
timestamp 1624494425
transform 1 0 351 0 1 8653
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_236
timestamp 1624494425
transform -1 0 624 0 1 8690
box -42 -55 624 371
use contact_9  contact_9_469
timestamp 1624494425
transform 1 0 351 0 1 9206
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_235
timestamp 1624494425
transform -1 0 624 0 -1 9480
box -42 -55 624 371
use contact_9  contact_9_468
timestamp 1624494425
transform 1 0 351 0 1 9443
box 0 0 66 74
use contact_9  contact_9_467
timestamp 1624494425
transform 1 0 351 0 1 9680
box 0 0 66 74
use contact_9  contact_9_466
timestamp 1624494425
transform 1 0 351 0 1 9443
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_234
timestamp 1624494425
transform -1 0 624 0 1 9480
box -42 -55 624 371
use contact_9  contact_9_465
timestamp 1624494425
transform 1 0 351 0 1 9996
box 0 0 66 74
use contact_9  contact_9_464
timestamp 1624494425
transform 1 0 351 0 1 10233
box 0 0 66 74
use contact_9  contact_9_462
timestamp 1624494425
transform 1 0 351 0 1 10233
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_232
timestamp 1624494425
transform -1 0 624 0 1 10270
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_233
timestamp 1624494425
transform -1 0 624 0 -1 10270
box -42 -55 624 371
use contact_9  contact_9_463
timestamp 1624494425
transform 1 0 351 0 1 10470
box 0 0 66 74
use contact_9  contact_9_461
timestamp 1624494425
transform 1 0 351 0 1 10786
box 0 0 66 74
use contact_9  contact_9_460
timestamp 1624494425
transform 1 0 351 0 1 11023
box 0 0 66 74
use contact_9  contact_9_458
timestamp 1624494425
transform 1 0 351 0 1 11023
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_230
timestamp 1624494425
transform -1 0 624 0 1 11060
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_231
timestamp 1624494425
transform -1 0 624 0 -1 11060
box -42 -55 624 371
use contact_9  contact_9_459
timestamp 1624494425
transform 1 0 351 0 1 11260
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_229
timestamp 1624494425
transform -1 0 624 0 -1 11850
box -42 -55 624 371
use contact_9  contact_9_457
timestamp 1624494425
transform 1 0 351 0 1 11576
box 0 0 66 74
use contact_9  contact_9_456
timestamp 1624494425
transform 1 0 351 0 1 11813
box 0 0 66 74
use contact_9  contact_9_454
timestamp 1624494425
transform 1 0 351 0 1 11813
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_228
timestamp 1624494425
transform -1 0 624 0 1 11850
box -42 -55 624 371
use contact_9  contact_9_455
timestamp 1624494425
transform 1 0 351 0 1 12050
box 0 0 66 74
use contact_9  contact_9_453
timestamp 1624494425
transform 1 0 351 0 1 12366
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_227
timestamp 1624494425
transform -1 0 624 0 -1 12640
box -42 -55 624 371
use contact_9  contact_9_452
timestamp 1624494425
transform 1 0 351 0 1 12603
box 0 0 66 74
use contact_9  contact_9_450
timestamp 1624494425
transform 1 0 351 0 1 12603
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_226
timestamp 1624494425
transform -1 0 624 0 1 12640
box -42 -55 624 371
use contact_9  contact_9_451
timestamp 1624494425
transform 1 0 351 0 1 12840
box 0 0 66 74
use contact_9  contact_9_449
timestamp 1624494425
transform 1 0 351 0 1 13156
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_225
timestamp 1624494425
transform -1 0 624 0 -1 13430
box -42 -55 624 371
use contact_9  contact_9_448
timestamp 1624494425
transform 1 0 351 0 1 13393
box 0 0 66 74
use contact_9  contact_9_447
timestamp 1624494425
transform 1 0 351 0 1 13630
box 0 0 66 74
use contact_9  contact_9_446
timestamp 1624494425
transform 1 0 351 0 1 13393
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_224
timestamp 1624494425
transform -1 0 624 0 1 13430
box -42 -55 624 371
use contact_9  contact_9_445
timestamp 1624494425
transform 1 0 351 0 1 13946
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_223
timestamp 1624494425
transform -1 0 624 0 -1 14220
box -42 -55 624 371
use contact_9  contact_9_444
timestamp 1624494425
transform 1 0 351 0 1 14183
box 0 0 66 74
use contact_9  contact_9_443
timestamp 1624494425
transform 1 0 351 0 1 14420
box 0 0 66 74
use contact_9  contact_9_442
timestamp 1624494425
transform 1 0 351 0 1 14183
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_222
timestamp 1624494425
transform -1 0 624 0 1 14220
box -42 -55 624 371
use contact_9  contact_9_441
timestamp 1624494425
transform 1 0 351 0 1 14736
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_221
timestamp 1624494425
transform -1 0 624 0 -1 15010
box -42 -55 624 371
use contact_9  contact_9_440
timestamp 1624494425
transform 1 0 351 0 1 14973
box 0 0 66 74
use contact_9  contact_9_439
timestamp 1624494425
transform 1 0 351 0 1 15210
box 0 0 66 74
use contact_9  contact_9_438
timestamp 1624494425
transform 1 0 351 0 1 14973
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_220
timestamp 1624494425
transform -1 0 624 0 1 15010
box -42 -55 624 371
use contact_9  contact_9_437
timestamp 1624494425
transform 1 0 351 0 1 15526
box 0 0 66 74
use contact_9  contact_9_436
timestamp 1624494425
transform 1 0 351 0 1 15763
box 0 0 66 74
use contact_9  contact_9_434
timestamp 1624494425
transform 1 0 351 0 1 15763
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_218
timestamp 1624494425
transform -1 0 624 0 1 15800
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_219
timestamp 1624494425
transform -1 0 624 0 -1 15800
box -42 -55 624 371
use contact_9  contact_9_435
timestamp 1624494425
transform 1 0 351 0 1 16000
box 0 0 66 74
use contact_9  contact_9_433
timestamp 1624494425
transform 1 0 351 0 1 16316
box 0 0 66 74
use contact_9  contact_9_432
timestamp 1624494425
transform 1 0 351 0 1 16553
box 0 0 66 74
use contact_9  contact_9_430
timestamp 1624494425
transform 1 0 351 0 1 16553
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_216
timestamp 1624494425
transform -1 0 624 0 1 16590
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_217
timestamp 1624494425
transform -1 0 624 0 -1 16590
box -42 -55 624 371
use contact_9  contact_9_431
timestamp 1624494425
transform 1 0 351 0 1 16790
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_215
timestamp 1624494425
transform -1 0 624 0 -1 17380
box -42 -55 624 371
use contact_9  contact_9_429
timestamp 1624494425
transform 1 0 351 0 1 17106
box 0 0 66 74
use contact_9  contact_9_428
timestamp 1624494425
transform 1 0 351 0 1 17343
box 0 0 66 74
use contact_9  contact_9_426
timestamp 1624494425
transform 1 0 351 0 1 17343
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_214
timestamp 1624494425
transform -1 0 624 0 1 17380
box -42 -55 624 371
use contact_9  contact_9_427
timestamp 1624494425
transform 1 0 351 0 1 17580
box 0 0 66 74
use contact_9  contact_9_425
timestamp 1624494425
transform 1 0 351 0 1 17896
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_213
timestamp 1624494425
transform -1 0 624 0 -1 18170
box -42 -55 624 371
use contact_9  contact_9_424
timestamp 1624494425
transform 1 0 351 0 1 18133
box 0 0 66 74
use contact_9  contact_9_422
timestamp 1624494425
transform 1 0 351 0 1 18133
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_212
timestamp 1624494425
transform -1 0 624 0 1 18170
box -42 -55 624 371
use contact_9  contact_9_423
timestamp 1624494425
transform 1 0 351 0 1 18370
box 0 0 66 74
use contact_9  contact_9_421
timestamp 1624494425
transform 1 0 351 0 1 18686
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_211
timestamp 1624494425
transform -1 0 624 0 -1 18960
box -42 -55 624 371
use contact_9  contact_9_420
timestamp 1624494425
transform 1 0 351 0 1 18923
box 0 0 66 74
use contact_9  contact_9_419
timestamp 1624494425
transform 1 0 351 0 1 19160
box 0 0 66 74
use contact_9  contact_9_418
timestamp 1624494425
transform 1 0 351 0 1 18923
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_210
timestamp 1624494425
transform -1 0 624 0 1 18960
box -42 -55 624 371
use contact_9  contact_9_417
timestamp 1624494425
transform 1 0 351 0 1 19476
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_209
timestamp 1624494425
transform -1 0 624 0 -1 19750
box -42 -55 624 371
use contact_9  contact_9_416
timestamp 1624494425
transform 1 0 351 0 1 19713
box 0 0 66 74
use contact_9  contact_9_415
timestamp 1624494425
transform 1 0 351 0 1 19950
box 0 0 66 74
use contact_9  contact_9_414
timestamp 1624494425
transform 1 0 351 0 1 19713
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_208
timestamp 1624494425
transform -1 0 624 0 1 19750
box -42 -55 624 371
use contact_9  contact_9_413
timestamp 1624494425
transform 1 0 351 0 1 20266
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_206
timestamp 1624494425
transform -1 0 624 0 1 20540
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_207
timestamp 1624494425
transform -1 0 624 0 -1 20540
box -42 -55 624 371
use contact_9  contact_9_412
timestamp 1624494425
transform 1 0 351 0 1 20503
box 0 0 66 74
use contact_9  contact_9_411
timestamp 1624494425
transform 1 0 351 0 1 20740
box 0 0 66 74
use contact_9  contact_9_410
timestamp 1624494425
transform 1 0 351 0 1 20503
box 0 0 66 74
use contact_9  contact_9_409
timestamp 1624494425
transform 1 0 351 0 1 21056
box 0 0 66 74
use contact_9  contact_9_408
timestamp 1624494425
transform 1 0 351 0 1 21293
box 0 0 66 74
use contact_9  contact_9_406
timestamp 1624494425
transform 1 0 351 0 1 21293
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_204
timestamp 1624494425
transform -1 0 624 0 1 21330
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_205
timestamp 1624494425
transform -1 0 624 0 -1 21330
box -42 -55 624 371
use contact_9  contact_9_407
timestamp 1624494425
transform 1 0 351 0 1 21530
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_203
timestamp 1624494425
transform -1 0 624 0 -1 22120
box -42 -55 624 371
use contact_9  contact_9_405
timestamp 1624494425
transform 1 0 351 0 1 21846
box 0 0 66 74
use contact_9  contact_9_404
timestamp 1624494425
transform 1 0 351 0 1 22083
box 0 0 66 74
use contact_9  contact_9_402
timestamp 1624494425
transform 1 0 351 0 1 22083
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_202
timestamp 1624494425
transform -1 0 624 0 1 22120
box -42 -55 624 371
use contact_9  contact_9_403
timestamp 1624494425
transform 1 0 351 0 1 22320
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_201
timestamp 1624494425
transform -1 0 624 0 -1 22910
box -42 -55 624 371
use contact_9  contact_9_401
timestamp 1624494425
transform 1 0 351 0 1 22636
box 0 0 66 74
use contact_9  contact_9_400
timestamp 1624494425
transform 1 0 351 0 1 22873
box 0 0 66 74
use contact_9  contact_9_398
timestamp 1624494425
transform 1 0 351 0 1 22873
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_200
timestamp 1624494425
transform -1 0 624 0 1 22910
box -42 -55 624 371
use contact_9  contact_9_399
timestamp 1624494425
transform 1 0 351 0 1 23110
box 0 0 66 74
use contact_9  contact_9_397
timestamp 1624494425
transform 1 0 351 0 1 23426
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_199
timestamp 1624494425
transform -1 0 624 0 -1 23700
box -42 -55 624 371
use contact_9  contact_9_396
timestamp 1624494425
transform 1 0 351 0 1 23663
box 0 0 66 74
use contact_9  contact_9_395
timestamp 1624494425
transform 1 0 351 0 1 23900
box 0 0 66 74
use contact_9  contact_9_394
timestamp 1624494425
transform 1 0 351 0 1 23663
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_198
timestamp 1624494425
transform -1 0 624 0 1 23700
box -42 -55 624 371
use contact_9  contact_9_393
timestamp 1624494425
transform 1 0 351 0 1 24216
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_197
timestamp 1624494425
transform -1 0 624 0 -1 24490
box -42 -55 624 371
use contact_9  contact_9_392
timestamp 1624494425
transform 1 0 351 0 1 24453
box 0 0 66 74
use contact_9  contact_9_391
timestamp 1624494425
transform 1 0 351 0 1 24690
box 0 0 66 74
use contact_9  contact_9_390
timestamp 1624494425
transform 1 0 351 0 1 24453
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_196
timestamp 1624494425
transform -1 0 624 0 1 24490
box -42 -55 624 371
use contact_9  contact_9_389
timestamp 1624494425
transform 1 0 351 0 1 25006
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_195
timestamp 1624494425
transform -1 0 624 0 -1 25280
box -42 -55 624 371
use contact_9  contact_9_388
timestamp 1624494425
transform 1 0 351 0 1 25243
box 0 0 66 74
use contact_9  contact_9_387
timestamp 1624494425
transform 1 0 351 0 1 25480
box 0 0 66 74
use contact_9  contact_9_386
timestamp 1624494425
transform 1 0 351 0 1 25243
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_194
timestamp 1624494425
transform -1 0 624 0 1 25280
box -42 -55 624 371
use contact_9  contact_9_385
timestamp 1624494425
transform 1 0 351 0 1 25796
box 0 0 66 74
use contact_9  contact_9_384
timestamp 1624494425
transform 1 0 351 0 1 26033
box 0 0 66 74
use contact_9  contact_9_382
timestamp 1624494425
transform 1 0 351 0 1 26033
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_192
timestamp 1624494425
transform -1 0 624 0 1 26070
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_193
timestamp 1624494425
transform -1 0 624 0 -1 26070
box -42 -55 624 371
use contact_9  contact_9_383
timestamp 1624494425
transform 1 0 351 0 1 26270
box 0 0 66 74
use contact_9  contact_9_381
timestamp 1624494425
transform 1 0 351 0 1 26586
box 0 0 66 74
use contact_9  contact_9_380
timestamp 1624494425
transform 1 0 351 0 1 26823
box 0 0 66 74
use contact_9  contact_9_378
timestamp 1624494425
transform 1 0 351 0 1 26823
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_190
timestamp 1624494425
transform -1 0 624 0 1 26860
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_191
timestamp 1624494425
transform -1 0 624 0 -1 26860
box -42 -55 624 371
use contact_9  contact_9_379
timestamp 1624494425
transform 1 0 351 0 1 27060
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_189
timestamp 1624494425
transform -1 0 624 0 -1 27650
box -42 -55 624 371
use contact_9  contact_9_377
timestamp 1624494425
transform 1 0 351 0 1 27376
box 0 0 66 74
use contact_9  contact_9_376
timestamp 1624494425
transform 1 0 351 0 1 27613
box 0 0 66 74
use contact_9  contact_9_374
timestamp 1624494425
transform 1 0 351 0 1 27613
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_188
timestamp 1624494425
transform -1 0 624 0 1 27650
box -42 -55 624 371
use contact_9  contact_9_375
timestamp 1624494425
transform 1 0 351 0 1 27850
box 0 0 66 74
use contact_9  contact_9_373
timestamp 1624494425
transform 1 0 351 0 1 28166
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_187
timestamp 1624494425
transform -1 0 624 0 -1 28440
box -42 -55 624 371
use contact_9  contact_9_372
timestamp 1624494425
transform 1 0 351 0 1 28403
box 0 0 66 74
use contact_9  contact_9_370
timestamp 1624494425
transform 1 0 351 0 1 28403
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_186
timestamp 1624494425
transform -1 0 624 0 1 28440
box -42 -55 624 371
use contact_9  contact_9_371
timestamp 1624494425
transform 1 0 351 0 1 28640
box 0 0 66 74
use contact_9  contact_9_369
timestamp 1624494425
transform 1 0 351 0 1 28956
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_185
timestamp 1624494425
transform -1 0 624 0 -1 29230
box -42 -55 624 371
use contact_9  contact_9_368
timestamp 1624494425
transform 1 0 351 0 1 29193
box 0 0 66 74
use contact_9  contact_9_367
timestamp 1624494425
transform 1 0 351 0 1 29430
box 0 0 66 74
use contact_9  contact_9_366
timestamp 1624494425
transform 1 0 351 0 1 29193
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_184
timestamp 1624494425
transform -1 0 624 0 1 29230
box -42 -55 624 371
use contact_9  contact_9_365
timestamp 1624494425
transform 1 0 351 0 1 29746
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_183
timestamp 1624494425
transform -1 0 624 0 -1 30020
box -42 -55 624 371
use contact_9  contact_9_364
timestamp 1624494425
transform 1 0 351 0 1 29983
box 0 0 66 74
use contact_9  contact_9_363
timestamp 1624494425
transform 1 0 351 0 1 30220
box 0 0 66 74
use contact_9  contact_9_362
timestamp 1624494425
transform 1 0 351 0 1 29983
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_182
timestamp 1624494425
transform -1 0 624 0 1 30020
box -42 -55 624 371
use contact_9  contact_9_361
timestamp 1624494425
transform 1 0 351 0 1 30536
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_181
timestamp 1624494425
transform -1 0 624 0 -1 30810
box -42 -55 624 371
use contact_9  contact_9_360
timestamp 1624494425
transform 1 0 351 0 1 30773
box 0 0 66 74
use contact_9  contact_9_359
timestamp 1624494425
transform 1 0 351 0 1 31010
box 0 0 66 74
use contact_9  contact_9_358
timestamp 1624494425
transform 1 0 351 0 1 30773
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_180
timestamp 1624494425
transform -1 0 624 0 1 30810
box -42 -55 624 371
use contact_9  contact_9_357
timestamp 1624494425
transform 1 0 351 0 1 31326
box 0 0 66 74
use contact_9  contact_9_356
timestamp 1624494425
transform 1 0 351 0 1 31563
box 0 0 66 74
use contact_9  contact_9_354
timestamp 1624494425
transform 1 0 351 0 1 31563
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_178
timestamp 1624494425
transform -1 0 624 0 1 31600
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_179
timestamp 1624494425
transform -1 0 624 0 -1 31600
box -42 -55 624 371
use contact_9  contact_9_355
timestamp 1624494425
transform 1 0 351 0 1 31800
box 0 0 66 74
use contact_9  contact_9_353
timestamp 1624494425
transform 1 0 351 0 1 32116
box 0 0 66 74
use contact_9  contact_9_352
timestamp 1624494425
transform 1 0 351 0 1 32353
box 0 0 66 74
use contact_9  contact_9_350
timestamp 1624494425
transform 1 0 351 0 1 32353
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_176
timestamp 1624494425
transform -1 0 624 0 1 32390
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_177
timestamp 1624494425
transform -1 0 624 0 -1 32390
box -42 -55 624 371
use contact_9  contact_9_351
timestamp 1624494425
transform 1 0 351 0 1 32590
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_175
timestamp 1624494425
transform -1 0 624 0 -1 33180
box -42 -55 624 371
use contact_9  contact_9_349
timestamp 1624494425
transform 1 0 351 0 1 32906
box 0 0 66 74
use contact_9  contact_9_348
timestamp 1624494425
transform 1 0 351 0 1 33143
box 0 0 66 74
use contact_9  contact_9_346
timestamp 1624494425
transform 1 0 351 0 1 33143
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_174
timestamp 1624494425
transform -1 0 624 0 1 33180
box -42 -55 624 371
use contact_9  contact_9_347
timestamp 1624494425
transform 1 0 351 0 1 33380
box 0 0 66 74
use contact_9  contact_9_345
timestamp 1624494425
transform 1 0 351 0 1 33696
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_173
timestamp 1624494425
transform -1 0 624 0 -1 33970
box -42 -55 624 371
use contact_9  contact_9_344
timestamp 1624494425
transform 1 0 351 0 1 33933
box 0 0 66 74
use contact_9  contact_9_342
timestamp 1624494425
transform 1 0 351 0 1 33933
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_172
timestamp 1624494425
transform -1 0 624 0 1 33970
box -42 -55 624 371
use contact_9  contact_9_343
timestamp 1624494425
transform 1 0 351 0 1 34170
box 0 0 66 74
use contact_9  contact_9_341
timestamp 1624494425
transform 1 0 351 0 1 34486
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_171
timestamp 1624494425
transform -1 0 624 0 -1 34760
box -42 -55 624 371
use contact_9  contact_9_340
timestamp 1624494425
transform 1 0 351 0 1 34723
box 0 0 66 74
use contact_9  contact_9_339
timestamp 1624494425
transform 1 0 351 0 1 34960
box 0 0 66 74
use contact_9  contact_9_338
timestamp 1624494425
transform 1 0 351 0 1 34723
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_170
timestamp 1624494425
transform -1 0 624 0 1 34760
box -42 -55 624 371
use contact_9  contact_9_337
timestamp 1624494425
transform 1 0 351 0 1 35276
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_169
timestamp 1624494425
transform -1 0 624 0 -1 35550
box -42 -55 624 371
use contact_9  contact_9_336
timestamp 1624494425
transform 1 0 351 0 1 35513
box 0 0 66 74
use contact_9  contact_9_335
timestamp 1624494425
transform 1 0 351 0 1 35750
box 0 0 66 74
use contact_9  contact_9_334
timestamp 1624494425
transform 1 0 351 0 1 35513
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_168
timestamp 1624494425
transform -1 0 624 0 1 35550
box -42 -55 624 371
use contact_9  contact_9_333
timestamp 1624494425
transform 1 0 351 0 1 36066
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_166
timestamp 1624494425
transform -1 0 624 0 1 36340
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_167
timestamp 1624494425
transform -1 0 624 0 -1 36340
box -42 -55 624 371
use contact_9  contact_9_332
timestamp 1624494425
transform 1 0 351 0 1 36303
box 0 0 66 74
use contact_9  contact_9_331
timestamp 1624494425
transform 1 0 351 0 1 36540
box 0 0 66 74
use contact_9  contact_9_330
timestamp 1624494425
transform 1 0 351 0 1 36303
box 0 0 66 74
use contact_9  contact_9_329
timestamp 1624494425
transform 1 0 351 0 1 36856
box 0 0 66 74
use contact_9  contact_9_328
timestamp 1624494425
transform 1 0 351 0 1 37093
box 0 0 66 74
use contact_9  contact_9_326
timestamp 1624494425
transform 1 0 351 0 1 37093
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_164
timestamp 1624494425
transform -1 0 624 0 1 37130
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_165
timestamp 1624494425
transform -1 0 624 0 -1 37130
box -42 -55 624 371
use contact_9  contact_9_327
timestamp 1624494425
transform 1 0 351 0 1 37330
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_163
timestamp 1624494425
transform -1 0 624 0 -1 37920
box -42 -55 624 371
use contact_9  contact_9_325
timestamp 1624494425
transform 1 0 351 0 1 37646
box 0 0 66 74
use contact_9  contact_9_324
timestamp 1624494425
transform 1 0 351 0 1 37883
box 0 0 66 74
use contact_9  contact_9_322
timestamp 1624494425
transform 1 0 351 0 1 37883
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_162
timestamp 1624494425
transform -1 0 624 0 1 37920
box -42 -55 624 371
use contact_9  contact_9_323
timestamp 1624494425
transform 1 0 351 0 1 38120
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_161
timestamp 1624494425
transform -1 0 624 0 -1 38710
box -42 -55 624 371
use contact_9  contact_9_321
timestamp 1624494425
transform 1 0 351 0 1 38436
box 0 0 66 74
use contact_9  contact_9_320
timestamp 1624494425
transform 1 0 351 0 1 38673
box 0 0 66 74
use contact_9  contact_9_318
timestamp 1624494425
transform 1 0 351 0 1 38673
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_160
timestamp 1624494425
transform -1 0 624 0 1 38710
box -42 -55 624 371
use contact_9  contact_9_319
timestamp 1624494425
transform 1 0 351 0 1 38910
box 0 0 66 74
use contact_9  contact_9_317
timestamp 1624494425
transform 1 0 351 0 1 39226
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_159
timestamp 1624494425
transform -1 0 624 0 -1 39500
box -42 -55 624 371
use contact_9  contact_9_316
timestamp 1624494425
transform 1 0 351 0 1 39463
box 0 0 66 74
use contact_9  contact_9_315
timestamp 1624494425
transform 1 0 351 0 1 39700
box 0 0 66 74
use contact_9  contact_9_314
timestamp 1624494425
transform 1 0 351 0 1 39463
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_158
timestamp 1624494425
transform -1 0 624 0 1 39500
box -42 -55 624 371
use contact_9  contact_9_313
timestamp 1624494425
transform 1 0 351 0 1 40016
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_157
timestamp 1624494425
transform -1 0 624 0 -1 40290
box -42 -55 624 371
use contact_9  contact_9_312
timestamp 1624494425
transform 1 0 351 0 1 40253
box 0 0 66 74
use contact_9  contact_9_311
timestamp 1624494425
transform 1 0 351 0 1 40490
box 0 0 66 74
use contact_9  contact_9_310
timestamp 1624494425
transform 1 0 351 0 1 40253
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_156
timestamp 1624494425
transform -1 0 624 0 1 40290
box -42 -55 624 371
use contact_9  contact_9_309
timestamp 1624494425
transform 1 0 351 0 1 40806
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_155
timestamp 1624494425
transform -1 0 624 0 -1 41080
box -42 -55 624 371
use contact_9  contact_9_308
timestamp 1624494425
transform 1 0 351 0 1 41043
box 0 0 66 74
use contact_9  contact_9_307
timestamp 1624494425
transform 1 0 351 0 1 41280
box 0 0 66 74
use contact_9  contact_9_306
timestamp 1624494425
transform 1 0 351 0 1 41043
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_154
timestamp 1624494425
transform -1 0 624 0 1 41080
box -42 -55 624 371
use contact_9  contact_9_305
timestamp 1624494425
transform 1 0 351 0 1 41596
box 0 0 66 74
use contact_9  contact_9_304
timestamp 1624494425
transform 1 0 351 0 1 41833
box 0 0 66 74
use contact_9  contact_9_302
timestamp 1624494425
transform 1 0 351 0 1 41833
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_152
timestamp 1624494425
transform -1 0 624 0 1 41870
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_153
timestamp 1624494425
transform -1 0 624 0 -1 41870
box -42 -55 624 371
use contact_9  contact_9_303
timestamp 1624494425
transform 1 0 351 0 1 42070
box 0 0 66 74
use contact_9  contact_9_301
timestamp 1624494425
transform 1 0 351 0 1 42386
box 0 0 66 74
use contact_9  contact_9_300
timestamp 1624494425
transform 1 0 351 0 1 42623
box 0 0 66 74
use contact_9  contact_9_298
timestamp 1624494425
transform 1 0 351 0 1 42623
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_150
timestamp 1624494425
transform -1 0 624 0 1 42660
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_151
timestamp 1624494425
transform -1 0 624 0 -1 42660
box -42 -55 624 371
use contact_9  contact_9_299
timestamp 1624494425
transform 1 0 351 0 1 42860
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_149
timestamp 1624494425
transform -1 0 624 0 -1 43450
box -42 -55 624 371
use contact_9  contact_9_297
timestamp 1624494425
transform 1 0 351 0 1 43176
box 0 0 66 74
use contact_9  contact_9_296
timestamp 1624494425
transform 1 0 351 0 1 43413
box 0 0 66 74
use contact_9  contact_9_294
timestamp 1624494425
transform 1 0 351 0 1 43413
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_148
timestamp 1624494425
transform -1 0 624 0 1 43450
box -42 -55 624 371
use contact_9  contact_9_295
timestamp 1624494425
transform 1 0 351 0 1 43650
box 0 0 66 74
use contact_9  contact_9_293
timestamp 1624494425
transform 1 0 351 0 1 43966
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_147
timestamp 1624494425
transform -1 0 624 0 -1 44240
box -42 -55 624 371
use contact_9  contact_9_292
timestamp 1624494425
transform 1 0 351 0 1 44203
box 0 0 66 74
use contact_9  contact_9_290
timestamp 1624494425
transform 1 0 351 0 1 44203
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_146
timestamp 1624494425
transform -1 0 624 0 1 44240
box -42 -55 624 371
use contact_9  contact_9_291
timestamp 1624494425
transform 1 0 351 0 1 44440
box 0 0 66 74
use contact_9  contact_9_289
timestamp 1624494425
transform 1 0 351 0 1 44756
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_145
timestamp 1624494425
transform -1 0 624 0 -1 45030
box -42 -55 624 371
use contact_9  contact_9_288
timestamp 1624494425
transform 1 0 351 0 1 44993
box 0 0 66 74
use contact_9  contact_9_287
timestamp 1624494425
transform 1 0 351 0 1 45230
box 0 0 66 74
use contact_9  contact_9_286
timestamp 1624494425
transform 1 0 351 0 1 44993
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_144
timestamp 1624494425
transform -1 0 624 0 1 45030
box -42 -55 624 371
use contact_9  contact_9_285
timestamp 1624494425
transform 1 0 351 0 1 45546
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_143
timestamp 1624494425
transform -1 0 624 0 -1 45820
box -42 -55 624 371
use contact_9  contact_9_284
timestamp 1624494425
transform 1 0 351 0 1 45783
box 0 0 66 74
use contact_9  contact_9_283
timestamp 1624494425
transform 1 0 351 0 1 46020
box 0 0 66 74
use contact_9  contact_9_282
timestamp 1624494425
transform 1 0 351 0 1 45783
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_142
timestamp 1624494425
transform -1 0 624 0 1 45820
box -42 -55 624 371
use contact_9  contact_9_281
timestamp 1624494425
transform 1 0 351 0 1 46336
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_141
timestamp 1624494425
transform -1 0 624 0 -1 46610
box -42 -55 624 371
use contact_9  contact_9_280
timestamp 1624494425
transform 1 0 351 0 1 46573
box 0 0 66 74
use contact_9  contact_9_279
timestamp 1624494425
transform 1 0 351 0 1 46810
box 0 0 66 74
use contact_9  contact_9_278
timestamp 1624494425
transform 1 0 351 0 1 46573
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_140
timestamp 1624494425
transform -1 0 624 0 1 46610
box -42 -55 624 371
use contact_9  contact_9_277
timestamp 1624494425
transform 1 0 351 0 1 47126
box 0 0 66 74
use contact_9  contact_9_276
timestamp 1624494425
transform 1 0 351 0 1 47363
box 0 0 66 74
use contact_9  contact_9_274
timestamp 1624494425
transform 1 0 351 0 1 47363
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_138
timestamp 1624494425
transform -1 0 624 0 1 47400
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_139
timestamp 1624494425
transform -1 0 624 0 -1 47400
box -42 -55 624 371
use contact_9  contact_9_275
timestamp 1624494425
transform 1 0 351 0 1 47600
box 0 0 66 74
use contact_9  contact_9_273
timestamp 1624494425
transform 1 0 351 0 1 47916
box 0 0 66 74
use contact_9  contact_9_272
timestamp 1624494425
transform 1 0 351 0 1 48153
box 0 0 66 74
use contact_9  contact_9_270
timestamp 1624494425
transform 1 0 351 0 1 48153
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_136
timestamp 1624494425
transform -1 0 624 0 1 48190
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_137
timestamp 1624494425
transform -1 0 624 0 -1 48190
box -42 -55 624 371
use contact_9  contact_9_271
timestamp 1624494425
transform 1 0 351 0 1 48390
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_135
timestamp 1624494425
transform -1 0 624 0 -1 48980
box -42 -55 624 371
use contact_9  contact_9_269
timestamp 1624494425
transform 1 0 351 0 1 48706
box 0 0 66 74
use contact_9  contact_9_268
timestamp 1624494425
transform 1 0 351 0 1 48943
box 0 0 66 74
use contact_9  contact_9_266
timestamp 1624494425
transform 1 0 351 0 1 48943
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_134
timestamp 1624494425
transform -1 0 624 0 1 48980
box -42 -55 624 371
use contact_9  contact_9_267
timestamp 1624494425
transform 1 0 351 0 1 49180
box 0 0 66 74
use contact_9  contact_9_265
timestamp 1624494425
transform 1 0 351 0 1 49496
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_133
timestamp 1624494425
transform -1 0 624 0 -1 49770
box -42 -55 624 371
use contact_9  contact_9_264
timestamp 1624494425
transform 1 0 351 0 1 49733
box 0 0 66 74
use contact_9  contact_9_262
timestamp 1624494425
transform 1 0 351 0 1 49733
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_132
timestamp 1624494425
transform -1 0 624 0 1 49770
box -42 -55 624 371
use contact_9  contact_9_263
timestamp 1624494425
transform 1 0 351 0 1 49970
box 0 0 66 74
use contact_9  contact_9_261
timestamp 1624494425
transform 1 0 351 0 1 50286
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_131
timestamp 1624494425
transform -1 0 624 0 -1 50560
box -42 -55 624 371
use contact_9  contact_9_260
timestamp 1624494425
transform 1 0 351 0 1 50523
box 0 0 66 74
use contact_9  contact_9_259
timestamp 1624494425
transform 1 0 351 0 1 50760
box 0 0 66 74
use contact_9  contact_9_258
timestamp 1624494425
transform 1 0 351 0 1 50523
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_130
timestamp 1624494425
transform -1 0 624 0 1 50560
box -42 -55 624 371
use contact_9  contact_9_257
timestamp 1624494425
transform 1 0 351 0 1 51076
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_129
timestamp 1624494425
transform -1 0 624 0 -1 51350
box -42 -55 624 371
use contact_9  contact_9_256
timestamp 1624494425
transform 1 0 351 0 1 51313
box 0 0 66 74
use contact_9  contact_9_255
timestamp 1624494425
transform 1 0 351 0 1 51550
box 0 0 66 74
use contact_9  contact_9_254
timestamp 1624494425
transform 1 0 351 0 1 51313
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_128
timestamp 1624494425
transform -1 0 624 0 1 51350
box -42 -55 624 371
use contact_9  contact_9_253
timestamp 1624494425
transform 1 0 351 0 1 51866
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_126
timestamp 1624494425
transform -1 0 624 0 1 52140
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_127
timestamp 1624494425
transform -1 0 624 0 -1 52140
box -42 -55 624 371
use contact_9  contact_9_252
timestamp 1624494425
transform 1 0 351 0 1 52103
box 0 0 66 74
use contact_9  contact_9_251
timestamp 1624494425
transform 1 0 351 0 1 52340
box 0 0 66 74
use contact_9  contact_9_250
timestamp 1624494425
transform 1 0 351 0 1 52103
box 0 0 66 74
use contact_9  contact_9_249
timestamp 1624494425
transform 1 0 351 0 1 52656
box 0 0 66 74
use contact_9  contact_9_248
timestamp 1624494425
transform 1 0 351 0 1 52893
box 0 0 66 74
use contact_9  contact_9_246
timestamp 1624494425
transform 1 0 351 0 1 52893
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_124
timestamp 1624494425
transform -1 0 624 0 1 52930
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_125
timestamp 1624494425
transform -1 0 624 0 -1 52930
box -42 -55 624 371
use contact_9  contact_9_247
timestamp 1624494425
transform 1 0 351 0 1 53130
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_123
timestamp 1624494425
transform -1 0 624 0 -1 53720
box -42 -55 624 371
use contact_9  contact_9_245
timestamp 1624494425
transform 1 0 351 0 1 53446
box 0 0 66 74
use contact_9  contact_9_244
timestamp 1624494425
transform 1 0 351 0 1 53683
box 0 0 66 74
use contact_9  contact_9_242
timestamp 1624494425
transform 1 0 351 0 1 53683
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_122
timestamp 1624494425
transform -1 0 624 0 1 53720
box -42 -55 624 371
use contact_9  contact_9_243
timestamp 1624494425
transform 1 0 351 0 1 53920
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_121
timestamp 1624494425
transform -1 0 624 0 -1 54510
box -42 -55 624 371
use contact_9  contact_9_241
timestamp 1624494425
transform 1 0 351 0 1 54236
box 0 0 66 74
use contact_9  contact_9_240
timestamp 1624494425
transform 1 0 351 0 1 54473
box 0 0 66 74
use contact_9  contact_9_238
timestamp 1624494425
transform 1 0 351 0 1 54473
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_120
timestamp 1624494425
transform -1 0 624 0 1 54510
box -42 -55 624 371
use contact_9  contact_9_239
timestamp 1624494425
transform 1 0 351 0 1 54710
box 0 0 66 74
use contact_9  contact_9_237
timestamp 1624494425
transform 1 0 351 0 1 55026
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_119
timestamp 1624494425
transform -1 0 624 0 -1 55300
box -42 -55 624 371
use contact_9  contact_9_236
timestamp 1624494425
transform 1 0 351 0 1 55263
box 0 0 66 74
use contact_9  contact_9_235
timestamp 1624494425
transform 1 0 351 0 1 55500
box 0 0 66 74
use contact_9  contact_9_234
timestamp 1624494425
transform 1 0 351 0 1 55263
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_118
timestamp 1624494425
transform -1 0 624 0 1 55300
box -42 -55 624 371
use contact_9  contact_9_233
timestamp 1624494425
transform 1 0 351 0 1 55816
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_117
timestamp 1624494425
transform -1 0 624 0 -1 56090
box -42 -55 624 371
use contact_9  contact_9_232
timestamp 1624494425
transform 1 0 351 0 1 56053
box 0 0 66 74
use contact_9  contact_9_231
timestamp 1624494425
transform 1 0 351 0 1 56290
box 0 0 66 74
use contact_9  contact_9_230
timestamp 1624494425
transform 1 0 351 0 1 56053
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_116
timestamp 1624494425
transform -1 0 624 0 1 56090
box -42 -55 624 371
use contact_9  contact_9_229
timestamp 1624494425
transform 1 0 351 0 1 56606
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_115
timestamp 1624494425
transform -1 0 624 0 -1 56880
box -42 -55 624 371
use contact_9  contact_9_228
timestamp 1624494425
transform 1 0 351 0 1 56843
box 0 0 66 74
use contact_9  contact_9_227
timestamp 1624494425
transform 1 0 351 0 1 57080
box 0 0 66 74
use contact_9  contact_9_226
timestamp 1624494425
transform 1 0 351 0 1 56843
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_114
timestamp 1624494425
transform -1 0 624 0 1 56880
box -42 -55 624 371
use contact_9  contact_9_225
timestamp 1624494425
transform 1 0 351 0 1 57396
box 0 0 66 74
use contact_9  contact_9_224
timestamp 1624494425
transform 1 0 351 0 1 57633
box 0 0 66 74
use contact_9  contact_9_222
timestamp 1624494425
transform 1 0 351 0 1 57633
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_112
timestamp 1624494425
transform -1 0 624 0 1 57670
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_113
timestamp 1624494425
transform -1 0 624 0 -1 57670
box -42 -55 624 371
use contact_9  contact_9_223
timestamp 1624494425
transform 1 0 351 0 1 57870
box 0 0 66 74
use contact_9  contact_9_221
timestamp 1624494425
transform 1 0 351 0 1 58186
box 0 0 66 74
use contact_9  contact_9_220
timestamp 1624494425
transform 1 0 351 0 1 58423
box 0 0 66 74
use contact_9  contact_9_218
timestamp 1624494425
transform 1 0 351 0 1 58423
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_110
timestamp 1624494425
transform -1 0 624 0 1 58460
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_111
timestamp 1624494425
transform -1 0 624 0 -1 58460
box -42 -55 624 371
use contact_9  contact_9_219
timestamp 1624494425
transform 1 0 351 0 1 58660
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_109
timestamp 1624494425
transform -1 0 624 0 -1 59250
box -42 -55 624 371
use contact_9  contact_9_217
timestamp 1624494425
transform 1 0 351 0 1 58976
box 0 0 66 74
use contact_9  contact_9_216
timestamp 1624494425
transform 1 0 351 0 1 59213
box 0 0 66 74
use contact_9  contact_9_214
timestamp 1624494425
transform 1 0 351 0 1 59213
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_108
timestamp 1624494425
transform -1 0 624 0 1 59250
box -42 -55 624 371
use contact_9  contact_9_215
timestamp 1624494425
transform 1 0 351 0 1 59450
box 0 0 66 74
use contact_9  contact_9_213
timestamp 1624494425
transform 1 0 351 0 1 59766
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_107
timestamp 1624494425
transform -1 0 624 0 -1 60040
box -42 -55 624 371
use contact_9  contact_9_212
timestamp 1624494425
transform 1 0 351 0 1 60003
box 0 0 66 74
use contact_9  contact_9_210
timestamp 1624494425
transform 1 0 351 0 1 60003
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_106
timestamp 1624494425
transform -1 0 624 0 1 60040
box -42 -55 624 371
use contact_9  contact_9_211
timestamp 1624494425
transform 1 0 351 0 1 60240
box 0 0 66 74
use contact_9  contact_9_209
timestamp 1624494425
transform 1 0 351 0 1 60556
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_105
timestamp 1624494425
transform -1 0 624 0 -1 60830
box -42 -55 624 371
use contact_9  contact_9_208
timestamp 1624494425
transform 1 0 351 0 1 60793
box 0 0 66 74
use contact_9  contact_9_207
timestamp 1624494425
transform 1 0 351 0 1 61030
box 0 0 66 74
use contact_9  contact_9_206
timestamp 1624494425
transform 1 0 351 0 1 60793
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_104
timestamp 1624494425
transform -1 0 624 0 1 60830
box -42 -55 624 371
use contact_9  contact_9_205
timestamp 1624494425
transform 1 0 351 0 1 61346
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_103
timestamp 1624494425
transform -1 0 624 0 -1 61620
box -42 -55 624 371
use contact_9  contact_9_204
timestamp 1624494425
transform 1 0 351 0 1 61583
box 0 0 66 74
use contact_9  contact_9_203
timestamp 1624494425
transform 1 0 351 0 1 61820
box 0 0 66 74
use contact_9  contact_9_202
timestamp 1624494425
transform 1 0 351 0 1 61583
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_102
timestamp 1624494425
transform -1 0 624 0 1 61620
box -42 -55 624 371
use contact_9  contact_9_201
timestamp 1624494425
transform 1 0 351 0 1 62136
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_101
timestamp 1624494425
transform -1 0 624 0 -1 62410
box -42 -55 624 371
use contact_9  contact_9_200
timestamp 1624494425
transform 1 0 351 0 1 62373
box 0 0 66 74
use contact_9  contact_9_199
timestamp 1624494425
transform 1 0 351 0 1 62610
box 0 0 66 74
use contact_9  contact_9_198
timestamp 1624494425
transform 1 0 351 0 1 62373
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_100
timestamp 1624494425
transform -1 0 624 0 1 62410
box -42 -55 624 371
use contact_9  contact_9_197
timestamp 1624494425
transform 1 0 351 0 1 62926
box 0 0 66 74
use contact_9  contact_9_196
timestamp 1624494425
transform 1 0 351 0 1 63163
box 0 0 66 74
use contact_9  contact_9_194
timestamp 1624494425
transform 1 0 351 0 1 63163
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_98
timestamp 1624494425
transform -1 0 624 0 1 63200
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_99
timestamp 1624494425
transform -1 0 624 0 -1 63200
box -42 -55 624 371
use contact_9  contact_9_195
timestamp 1624494425
transform 1 0 351 0 1 63400
box 0 0 66 74
use contact_9  contact_9_193
timestamp 1624494425
transform 1 0 351 0 1 63716
box 0 0 66 74
use contact_9  contact_9_192
timestamp 1624494425
transform 1 0 351 0 1 63953
box 0 0 66 74
use contact_9  contact_9_190
timestamp 1624494425
transform 1 0 351 0 1 63953
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_96
timestamp 1624494425
transform -1 0 624 0 1 63990
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_97
timestamp 1624494425
transform -1 0 624 0 -1 63990
box -42 -55 624 371
use contact_9  contact_9_191
timestamp 1624494425
transform 1 0 351 0 1 64190
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_95
timestamp 1624494425
transform -1 0 624 0 -1 64780
box -42 -55 624 371
use contact_9  contact_9_189
timestamp 1624494425
transform 1 0 351 0 1 64506
box 0 0 66 74
use contact_9  contact_9_188
timestamp 1624494425
transform 1 0 351 0 1 64743
box 0 0 66 74
use contact_9  contact_9_186
timestamp 1624494425
transform 1 0 351 0 1 64743
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_94
timestamp 1624494425
transform -1 0 624 0 1 64780
box -42 -55 624 371
use contact_9  contact_9_187
timestamp 1624494425
transform 1 0 351 0 1 64980
box 0 0 66 74
use contact_9  contact_9_185
timestamp 1624494425
transform 1 0 351 0 1 65296
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_93
timestamp 1624494425
transform -1 0 624 0 -1 65570
box -42 -55 624 371
use contact_9  contact_9_184
timestamp 1624494425
transform 1 0 351 0 1 65533
box 0 0 66 74
use contact_9  contact_9_182
timestamp 1624494425
transform 1 0 351 0 1 65533
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_92
timestamp 1624494425
transform -1 0 624 0 1 65570
box -42 -55 624 371
use contact_9  contact_9_183
timestamp 1624494425
transform 1 0 351 0 1 65770
box 0 0 66 74
use contact_9  contact_9_181
timestamp 1624494425
transform 1 0 351 0 1 66086
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_91
timestamp 1624494425
transform -1 0 624 0 -1 66360
box -42 -55 624 371
use contact_9  contact_9_180
timestamp 1624494425
transform 1 0 351 0 1 66323
box 0 0 66 74
use contact_9  contact_9_179
timestamp 1624494425
transform 1 0 351 0 1 66560
box 0 0 66 74
use contact_9  contact_9_178
timestamp 1624494425
transform 1 0 351 0 1 66323
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_90
timestamp 1624494425
transform -1 0 624 0 1 66360
box -42 -55 624 371
use contact_9  contact_9_177
timestamp 1624494425
transform 1 0 351 0 1 66876
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_89
timestamp 1624494425
transform -1 0 624 0 -1 67150
box -42 -55 624 371
use contact_9  contact_9_176
timestamp 1624494425
transform 1 0 351 0 1 67113
box 0 0 66 74
use contact_9  contact_9_175
timestamp 1624494425
transform 1 0 351 0 1 67350
box 0 0 66 74
use contact_9  contact_9_174
timestamp 1624494425
transform 1 0 351 0 1 67113
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_88
timestamp 1624494425
transform -1 0 624 0 1 67150
box -42 -55 624 371
use contact_9  contact_9_173
timestamp 1624494425
transform 1 0 351 0 1 67666
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_87
timestamp 1624494425
transform -1 0 624 0 -1 67940
box -42 -55 624 371
use contact_9  contact_9_172
timestamp 1624494425
transform 1 0 351 0 1 67903
box 0 0 66 74
use contact_9  contact_9_171
timestamp 1624494425
transform 1 0 351 0 1 68140
box 0 0 66 74
use contact_9  contact_9_170
timestamp 1624494425
transform 1 0 351 0 1 67903
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_86
timestamp 1624494425
transform -1 0 624 0 1 67940
box -42 -55 624 371
use contact_9  contact_9_169
timestamp 1624494425
transform 1 0 351 0 1 68456
box 0 0 66 74
use contact_9  contact_9_168
timestamp 1624494425
transform 1 0 351 0 1 68693
box 0 0 66 74
use contact_9  contact_9_166
timestamp 1624494425
transform 1 0 351 0 1 68693
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_84
timestamp 1624494425
transform -1 0 624 0 1 68730
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_85
timestamp 1624494425
transform -1 0 624 0 -1 68730
box -42 -55 624 371
use contact_9  contact_9_167
timestamp 1624494425
transform 1 0 351 0 1 68930
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_83
timestamp 1624494425
transform -1 0 624 0 -1 69520
box -42 -55 624 371
use contact_9  contact_9_165
timestamp 1624494425
transform 1 0 351 0 1 69246
box 0 0 66 74
use contact_9  contact_9_164
timestamp 1624494425
transform 1 0 351 0 1 69483
box 0 0 66 74
use contact_9  contact_9_162
timestamp 1624494425
transform 1 0 351 0 1 69483
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_82
timestamp 1624494425
transform -1 0 624 0 1 69520
box -42 -55 624 371
use contact_9  contact_9_163
timestamp 1624494425
transform 1 0 351 0 1 69720
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_81
timestamp 1624494425
transform -1 0 624 0 -1 70310
box -42 -55 624 371
use contact_9  contact_9_161
timestamp 1624494425
transform 1 0 351 0 1 70036
box 0 0 66 74
use contact_9  contact_9_160
timestamp 1624494425
transform 1 0 351 0 1 70273
box 0 0 66 74
use contact_9  contact_9_158
timestamp 1624494425
transform 1 0 351 0 1 70273
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_80
timestamp 1624494425
transform -1 0 624 0 1 70310
box -42 -55 624 371
use contact_9  contact_9_159
timestamp 1624494425
transform 1 0 351 0 1 70510
box 0 0 66 74
use contact_9  contact_9_157
timestamp 1624494425
transform 1 0 351 0 1 70826
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_79
timestamp 1624494425
transform -1 0 624 0 -1 71100
box -42 -55 624 371
use contact_9  contact_9_156
timestamp 1624494425
transform 1 0 351 0 1 71063
box 0 0 66 74
use contact_9  contact_9_155
timestamp 1624494425
transform 1 0 351 0 1 71300
box 0 0 66 74
use contact_9  contact_9_154
timestamp 1624494425
transform 1 0 351 0 1 71063
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_78
timestamp 1624494425
transform -1 0 624 0 1 71100
box -42 -55 624 371
use contact_9  contact_9_153
timestamp 1624494425
transform 1 0 351 0 1 71616
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_77
timestamp 1624494425
transform -1 0 624 0 -1 71890
box -42 -55 624 371
use contact_9  contact_9_152
timestamp 1624494425
transform 1 0 351 0 1 71853
box 0 0 66 74
use contact_9  contact_9_151
timestamp 1624494425
transform 1 0 351 0 1 72090
box 0 0 66 74
use contact_9  contact_9_150
timestamp 1624494425
transform 1 0 351 0 1 71853
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_76
timestamp 1624494425
transform -1 0 624 0 1 71890
box -42 -55 624 371
use contact_9  contact_9_149
timestamp 1624494425
transform 1 0 351 0 1 72406
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_75
timestamp 1624494425
transform -1 0 624 0 -1 72680
box -42 -55 624 371
use contact_9  contact_9_148
timestamp 1624494425
transform 1 0 351 0 1 72643
box 0 0 66 74
use contact_9  contact_9_147
timestamp 1624494425
transform 1 0 351 0 1 72880
box 0 0 66 74
use contact_9  contact_9_146
timestamp 1624494425
transform 1 0 351 0 1 72643
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_74
timestamp 1624494425
transform -1 0 624 0 1 72680
box -42 -55 624 371
use contact_9  contact_9_145
timestamp 1624494425
transform 1 0 351 0 1 73196
box 0 0 66 74
use contact_9  contact_9_144
timestamp 1624494425
transform 1 0 351 0 1 73433
box 0 0 66 74
use contact_9  contact_9_142
timestamp 1624494425
transform 1 0 351 0 1 73433
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_72
timestamp 1624494425
transform -1 0 624 0 1 73470
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_73
timestamp 1624494425
transform -1 0 624 0 -1 73470
box -42 -55 624 371
use contact_9  contact_9_143
timestamp 1624494425
transform 1 0 351 0 1 73670
box 0 0 66 74
use contact_9  contact_9_141
timestamp 1624494425
transform 1 0 351 0 1 73986
box 0 0 66 74
use contact_9  contact_9_140
timestamp 1624494425
transform 1 0 351 0 1 74223
box 0 0 66 74
use contact_9  contact_9_138
timestamp 1624494425
transform 1 0 351 0 1 74223
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_70
timestamp 1624494425
transform -1 0 624 0 1 74260
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_71
timestamp 1624494425
transform -1 0 624 0 -1 74260
box -42 -55 624 371
use contact_9  contact_9_139
timestamp 1624494425
transform 1 0 351 0 1 74460
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_69
timestamp 1624494425
transform -1 0 624 0 -1 75050
box -42 -55 624 371
use contact_9  contact_9_137
timestamp 1624494425
transform 1 0 351 0 1 74776
box 0 0 66 74
use contact_9  contact_9_136
timestamp 1624494425
transform 1 0 351 0 1 75013
box 0 0 66 74
use contact_9  contact_9_134
timestamp 1624494425
transform 1 0 351 0 1 75013
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_68
timestamp 1624494425
transform -1 0 624 0 1 75050
box -42 -55 624 371
use contact_9  contact_9_135
timestamp 1624494425
transform 1 0 351 0 1 75250
box 0 0 66 74
use contact_9  contact_9_133
timestamp 1624494425
transform 1 0 351 0 1 75566
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_67
timestamp 1624494425
transform -1 0 624 0 -1 75840
box -42 -55 624 371
use contact_9  contact_9_132
timestamp 1624494425
transform 1 0 351 0 1 75803
box 0 0 66 74
use contact_9  contact_9_130
timestamp 1624494425
transform 1 0 351 0 1 75803
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_66
timestamp 1624494425
transform -1 0 624 0 1 75840
box -42 -55 624 371
use contact_9  contact_9_131
timestamp 1624494425
transform 1 0 351 0 1 76040
box 0 0 66 74
use contact_9  contact_9_129
timestamp 1624494425
transform 1 0 351 0 1 76356
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_65
timestamp 1624494425
transform -1 0 624 0 -1 76630
box -42 -55 624 371
use contact_9  contact_9_128
timestamp 1624494425
transform 1 0 351 0 1 76593
box 0 0 66 74
use contact_9  contact_9_127
timestamp 1624494425
transform 1 0 351 0 1 76830
box 0 0 66 74
use contact_9  contact_9_126
timestamp 1624494425
transform 1 0 351 0 1 76593
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_64
timestamp 1624494425
transform -1 0 624 0 1 76630
box -42 -55 624 371
use contact_9  contact_9_125
timestamp 1624494425
transform 1 0 351 0 1 77146
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_63
timestamp 1624494425
transform -1 0 624 0 -1 77420
box -42 -55 624 371
use contact_9  contact_9_124
timestamp 1624494425
transform 1 0 351 0 1 77383
box 0 0 66 74
use contact_9  contact_9_123
timestamp 1624494425
transform 1 0 351 0 1 77620
box 0 0 66 74
use contact_9  contact_9_122
timestamp 1624494425
transform 1 0 351 0 1 77383
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_62
timestamp 1624494425
transform -1 0 624 0 1 77420
box -42 -55 624 371
use contact_9  contact_9_121
timestamp 1624494425
transform 1 0 351 0 1 77936
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_61
timestamp 1624494425
transform -1 0 624 0 -1 78210
box -42 -55 624 371
use contact_9  contact_9_120
timestamp 1624494425
transform 1 0 351 0 1 78173
box 0 0 66 74
use contact_9  contact_9_119
timestamp 1624494425
transform 1 0 351 0 1 78410
box 0 0 66 74
use contact_9  contact_9_118
timestamp 1624494425
transform 1 0 351 0 1 78173
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_60
timestamp 1624494425
transform -1 0 624 0 1 78210
box -42 -55 624 371
use contact_9  contact_9_117
timestamp 1624494425
transform 1 0 351 0 1 78726
box 0 0 66 74
use contact_9  contact_9_116
timestamp 1624494425
transform 1 0 351 0 1 78963
box 0 0 66 74
use contact_9  contact_9_114
timestamp 1624494425
transform 1 0 351 0 1 78963
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_58
timestamp 1624494425
transform -1 0 624 0 1 79000
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_59
timestamp 1624494425
transform -1 0 624 0 -1 79000
box -42 -55 624 371
use contact_9  contact_9_115
timestamp 1624494425
transform 1 0 351 0 1 79200
box 0 0 66 74
use contact_9  contact_9_113
timestamp 1624494425
transform 1 0 351 0 1 79516
box 0 0 66 74
use contact_9  contact_9_112
timestamp 1624494425
transform 1 0 351 0 1 79753
box 0 0 66 74
use contact_9  contact_9_110
timestamp 1624494425
transform 1 0 351 0 1 79753
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_56
timestamp 1624494425
transform -1 0 624 0 1 79790
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_57
timestamp 1624494425
transform -1 0 624 0 -1 79790
box -42 -55 624 371
use contact_9  contact_9_111
timestamp 1624494425
transform 1 0 351 0 1 79990
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_55
timestamp 1624494425
transform -1 0 624 0 -1 80580
box -42 -55 624 371
use contact_9  contact_9_109
timestamp 1624494425
transform 1 0 351 0 1 80306
box 0 0 66 74
use contact_9  contact_9_108
timestamp 1624494425
transform 1 0 351 0 1 80543
box 0 0 66 74
use contact_9  contact_9_106
timestamp 1624494425
transform 1 0 351 0 1 80543
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_54
timestamp 1624494425
transform -1 0 624 0 1 80580
box -42 -55 624 371
use contact_9  contact_9_107
timestamp 1624494425
transform 1 0 351 0 1 80780
box 0 0 66 74
use contact_9  contact_9_105
timestamp 1624494425
transform 1 0 351 0 1 81096
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_53
timestamp 1624494425
transform -1 0 624 0 -1 81370
box -42 -55 624 371
use contact_9  contact_9_104
timestamp 1624494425
transform 1 0 351 0 1 81333
box 0 0 66 74
use contact_9  contact_9_102
timestamp 1624494425
transform 1 0 351 0 1 81333
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_52
timestamp 1624494425
transform -1 0 624 0 1 81370
box -42 -55 624 371
use contact_9  contact_9_103
timestamp 1624494425
transform 1 0 351 0 1 81570
box 0 0 66 74
use contact_9  contact_9_101
timestamp 1624494425
transform 1 0 351 0 1 81886
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_51
timestamp 1624494425
transform -1 0 624 0 -1 82160
box -42 -55 624 371
use contact_9  contact_9_100
timestamp 1624494425
transform 1 0 351 0 1 82123
box 0 0 66 74
use contact_9  contact_9_99
timestamp 1624494425
transform 1 0 351 0 1 82360
box 0 0 66 74
use contact_9  contact_9_98
timestamp 1624494425
transform 1 0 351 0 1 82123
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_50
timestamp 1624494425
transform -1 0 624 0 1 82160
box -42 -55 624 371
use contact_9  contact_9_97
timestamp 1624494425
transform 1 0 351 0 1 82676
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_49
timestamp 1624494425
transform -1 0 624 0 -1 82950
box -42 -55 624 371
use contact_9  contact_9_96
timestamp 1624494425
transform 1 0 351 0 1 82913
box 0 0 66 74
use contact_9  contact_9_95
timestamp 1624494425
transform 1 0 351 0 1 83150
box 0 0 66 74
use contact_9  contact_9_94
timestamp 1624494425
transform 1 0 351 0 1 82913
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_48
timestamp 1624494425
transform -1 0 624 0 1 82950
box -42 -55 624 371
use contact_9  contact_9_93
timestamp 1624494425
transform 1 0 351 0 1 83466
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_47
timestamp 1624494425
transform -1 0 624 0 -1 83740
box -42 -55 624 371
use contact_9  contact_9_92
timestamp 1624494425
transform 1 0 351 0 1 83703
box 0 0 66 74
use contact_9  contact_9_91
timestamp 1624494425
transform 1 0 351 0 1 83940
box 0 0 66 74
use contact_9  contact_9_90
timestamp 1624494425
transform 1 0 351 0 1 83703
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_46
timestamp 1624494425
transform -1 0 624 0 1 83740
box -42 -55 624 371
use contact_9  contact_9_89
timestamp 1624494425
transform 1 0 351 0 1 84256
box 0 0 66 74
use contact_9  contact_9_88
timestamp 1624494425
transform 1 0 351 0 1 84493
box 0 0 66 74
use contact_9  contact_9_86
timestamp 1624494425
transform 1 0 351 0 1 84493
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_44
timestamp 1624494425
transform -1 0 624 0 1 84530
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_45
timestamp 1624494425
transform -1 0 624 0 -1 84530
box -42 -55 624 371
use contact_9  contact_9_87
timestamp 1624494425
transform 1 0 351 0 1 84730
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_43
timestamp 1624494425
transform -1 0 624 0 -1 85320
box -42 -55 624 371
use contact_9  contact_9_85
timestamp 1624494425
transform 1 0 351 0 1 85046
box 0 0 66 74
use contact_9  contact_9_84
timestamp 1624494425
transform 1 0 351 0 1 85283
box 0 0 66 74
use contact_9  contact_9_82
timestamp 1624494425
transform 1 0 351 0 1 85283
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_42
timestamp 1624494425
transform -1 0 624 0 1 85320
box -42 -55 624 371
use contact_9  contact_9_83
timestamp 1624494425
transform 1 0 351 0 1 85520
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_41
timestamp 1624494425
transform -1 0 624 0 -1 86110
box -42 -55 624 371
use contact_9  contact_9_81
timestamp 1624494425
transform 1 0 351 0 1 85836
box 0 0 66 74
use contact_9  contact_9_80
timestamp 1624494425
transform 1 0 351 0 1 86073
box 0 0 66 74
use contact_9  contact_9_78
timestamp 1624494425
transform 1 0 351 0 1 86073
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_40
timestamp 1624494425
transform -1 0 624 0 1 86110
box -42 -55 624 371
use contact_9  contact_9_79
timestamp 1624494425
transform 1 0 351 0 1 86310
box 0 0 66 74
use contact_9  contact_9_77
timestamp 1624494425
transform 1 0 351 0 1 86626
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_39
timestamp 1624494425
transform -1 0 624 0 -1 86900
box -42 -55 624 371
use contact_9  contact_9_76
timestamp 1624494425
transform 1 0 351 0 1 86863
box 0 0 66 74
use contact_9  contact_9_74
timestamp 1624494425
transform 1 0 351 0 1 86863
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_38
timestamp 1624494425
transform -1 0 624 0 1 86900
box -42 -55 624 371
use contact_9  contact_9_75
timestamp 1624494425
transform 1 0 351 0 1 87100
box 0 0 66 74
use contact_9  contact_9_73
timestamp 1624494425
transform 1 0 351 0 1 87416
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_37
timestamp 1624494425
transform -1 0 624 0 -1 87690
box -42 -55 624 371
use contact_9  contact_9_72
timestamp 1624494425
transform 1 0 351 0 1 87653
box 0 0 66 74
use contact_9  contact_9_71
timestamp 1624494425
transform 1 0 351 0 1 87890
box 0 0 66 74
use contact_9  contact_9_70
timestamp 1624494425
transform 1 0 351 0 1 87653
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_36
timestamp 1624494425
transform -1 0 624 0 1 87690
box -42 -55 624 371
use contact_9  contact_9_69
timestamp 1624494425
transform 1 0 351 0 1 88206
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_35
timestamp 1624494425
transform -1 0 624 0 -1 88480
box -42 -55 624 371
use contact_9  contact_9_68
timestamp 1624494425
transform 1 0 351 0 1 88443
box 0 0 66 74
use contact_9  contact_9_67
timestamp 1624494425
transform 1 0 351 0 1 88680
box 0 0 66 74
use contact_9  contact_9_66
timestamp 1624494425
transform 1 0 351 0 1 88443
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_34
timestamp 1624494425
transform -1 0 624 0 1 88480
box -42 -55 624 371
use contact_9  contact_9_65
timestamp 1624494425
transform 1 0 351 0 1 88996
box 0 0 66 74
use contact_9  contact_9_64
timestamp 1624494425
transform 1 0 351 0 1 89233
box 0 0 66 74
use contact_9  contact_9_62
timestamp 1624494425
transform 1 0 351 0 1 89233
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_32
timestamp 1624494425
transform -1 0 624 0 1 89270
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_33
timestamp 1624494425
transform -1 0 624 0 -1 89270
box -42 -55 624 371
use contact_9  contact_9_63
timestamp 1624494425
transform 1 0 351 0 1 89470
box 0 0 66 74
use contact_9  contact_9_61
timestamp 1624494425
transform 1 0 351 0 1 89786
box 0 0 66 74
use contact_9  contact_9_60
timestamp 1624494425
transform 1 0 351 0 1 90023
box 0 0 66 74
use contact_9  contact_9_58
timestamp 1624494425
transform 1 0 351 0 1 90023
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_30
timestamp 1624494425
transform -1 0 624 0 1 90060
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_31
timestamp 1624494425
transform -1 0 624 0 -1 90060
box -42 -55 624 371
use contact_9  contact_9_59
timestamp 1624494425
transform 1 0 351 0 1 90260
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_29
timestamp 1624494425
transform -1 0 624 0 -1 90850
box -42 -55 624 371
use contact_9  contact_9_57
timestamp 1624494425
transform 1 0 351 0 1 90576
box 0 0 66 74
use contact_9  contact_9_56
timestamp 1624494425
transform 1 0 351 0 1 90813
box 0 0 66 74
use contact_9  contact_9_54
timestamp 1624494425
transform 1 0 351 0 1 90813
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_28
timestamp 1624494425
transform -1 0 624 0 1 90850
box -42 -55 624 371
use contact_9  contact_9_55
timestamp 1624494425
transform 1 0 351 0 1 91050
box 0 0 66 74
use contact_9  contact_9_53
timestamp 1624494425
transform 1 0 351 0 1 91366
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_27
timestamp 1624494425
transform -1 0 624 0 -1 91640
box -42 -55 624 371
use contact_9  contact_9_52
timestamp 1624494425
transform 1 0 351 0 1 91603
box 0 0 66 74
use contact_9  contact_9_50
timestamp 1624494425
transform 1 0 351 0 1 91603
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_26
timestamp 1624494425
transform -1 0 624 0 1 91640
box -42 -55 624 371
use contact_9  contact_9_51
timestamp 1624494425
transform 1 0 351 0 1 91840
box 0 0 66 74
use contact_9  contact_9_49
timestamp 1624494425
transform 1 0 351 0 1 92156
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_25
timestamp 1624494425
transform -1 0 624 0 -1 92430
box -42 -55 624 371
use contact_9  contact_9_48
timestamp 1624494425
transform 1 0 351 0 1 92393
box 0 0 66 74
use contact_9  contact_9_47
timestamp 1624494425
transform 1 0 351 0 1 92630
box 0 0 66 74
use contact_9  contact_9_46
timestamp 1624494425
transform 1 0 351 0 1 92393
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_24
timestamp 1624494425
transform -1 0 624 0 1 92430
box -42 -55 624 371
use contact_9  contact_9_45
timestamp 1624494425
transform 1 0 351 0 1 92946
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_23
timestamp 1624494425
transform -1 0 624 0 -1 93220
box -42 -55 624 371
use contact_9  contact_9_44
timestamp 1624494425
transform 1 0 351 0 1 93183
box 0 0 66 74
use contact_9  contact_9_43
timestamp 1624494425
transform 1 0 351 0 1 93420
box 0 0 66 74
use contact_9  contact_9_42
timestamp 1624494425
transform 1 0 351 0 1 93183
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_22
timestamp 1624494425
transform -1 0 624 0 1 93220
box -42 -55 624 371
use contact_9  contact_9_41
timestamp 1624494425
transform 1 0 351 0 1 93736
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_21
timestamp 1624494425
transform -1 0 624 0 -1 94010
box -42 -55 624 371
use contact_9  contact_9_40
timestamp 1624494425
transform 1 0 351 0 1 93973
box 0 0 66 74
use contact_9  contact_9_39
timestamp 1624494425
transform 1 0 351 0 1 94210
box 0 0 66 74
use contact_9  contact_9_38
timestamp 1624494425
transform 1 0 351 0 1 93973
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_20
timestamp 1624494425
transform -1 0 624 0 1 94010
box -42 -55 624 371
use contact_9  contact_9_37
timestamp 1624494425
transform 1 0 351 0 1 94526
box 0 0 66 74
use contact_9  contact_9_36
timestamp 1624494425
transform 1 0 351 0 1 94763
box 0 0 66 74
use contact_9  contact_9_34
timestamp 1624494425
transform 1 0 351 0 1 94763
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_18
timestamp 1624494425
transform -1 0 624 0 1 94800
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_19
timestamp 1624494425
transform -1 0 624 0 -1 94800
box -42 -55 624 371
use contact_9  contact_9_35
timestamp 1624494425
transform 1 0 351 0 1 95000
box 0 0 66 74
use contact_9  contact_9_33
timestamp 1624494425
transform 1 0 351 0 1 95316
box 0 0 66 74
use contact_9  contact_9_32
timestamp 1624494425
transform 1 0 351 0 1 95553
box 0 0 66 74
use contact_9  contact_9_30
timestamp 1624494425
transform 1 0 351 0 1 95553
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_16
timestamp 1624494425
transform -1 0 624 0 1 95590
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_17
timestamp 1624494425
transform -1 0 624 0 -1 95590
box -42 -55 624 371
use contact_9  contact_9_31
timestamp 1624494425
transform 1 0 351 0 1 95790
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_15
timestamp 1624494425
transform -1 0 624 0 -1 96380
box -42 -55 624 371
use contact_9  contact_9_29
timestamp 1624494425
transform 1 0 351 0 1 96106
box 0 0 66 74
use contact_9  contact_9_28
timestamp 1624494425
transform 1 0 351 0 1 96343
box 0 0 66 74
use contact_9  contact_9_26
timestamp 1624494425
transform 1 0 351 0 1 96343
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_14
timestamp 1624494425
transform -1 0 624 0 1 96380
box -42 -55 624 371
use contact_9  contact_9_27
timestamp 1624494425
transform 1 0 351 0 1 96580
box 0 0 66 74
use contact_9  contact_9_25
timestamp 1624494425
transform 1 0 351 0 1 96896
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_13
timestamp 1624494425
transform -1 0 624 0 -1 97170
box -42 -55 624 371
use contact_9  contact_9_24
timestamp 1624494425
transform 1 0 351 0 1 97133
box 0 0 66 74
use contact_9  contact_9_22
timestamp 1624494425
transform 1 0 351 0 1 97133
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_12
timestamp 1624494425
transform -1 0 624 0 1 97170
box -42 -55 624 371
use contact_9  contact_9_23
timestamp 1624494425
transform 1 0 351 0 1 97370
box 0 0 66 74
use contact_9  contact_9_21
timestamp 1624494425
transform 1 0 351 0 1 97686
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_11
timestamp 1624494425
transform -1 0 624 0 -1 97960
box -42 -55 624 371
use contact_9  contact_9_20
timestamp 1624494425
transform 1 0 351 0 1 97923
box 0 0 66 74
use contact_9  contact_9_19
timestamp 1624494425
transform 1 0 351 0 1 98160
box 0 0 66 74
use contact_9  contact_9_18
timestamp 1624494425
transform 1 0 351 0 1 97923
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_10
timestamp 1624494425
transform -1 0 624 0 1 97960
box -42 -55 624 371
use contact_9  contact_9_17
timestamp 1624494425
transform 1 0 351 0 1 98476
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_9
timestamp 1624494425
transform -1 0 624 0 -1 98750
box -42 -55 624 371
use contact_9  contact_9_16
timestamp 1624494425
transform 1 0 351 0 1 98713
box 0 0 66 74
use contact_9  contact_9_15
timestamp 1624494425
transform 1 0 351 0 1 98950
box 0 0 66 74
use contact_9  contact_9_14
timestamp 1624494425
transform 1 0 351 0 1 98713
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_8
timestamp 1624494425
transform -1 0 624 0 1 98750
box -42 -55 624 371
use contact_9  contact_9_13
timestamp 1624494425
transform 1 0 351 0 1 99266
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_7
timestamp 1624494425
transform -1 0 624 0 -1 99540
box -42 -55 624 371
use contact_9  contact_9_12
timestamp 1624494425
transform 1 0 351 0 1 99503
box 0 0 66 74
use contact_9  contact_9_11
timestamp 1624494425
transform 1 0 351 0 1 99740
box 0 0 66 74
use contact_9  contact_9_10
timestamp 1624494425
transform 1 0 351 0 1 99503
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_6
timestamp 1624494425
transform -1 0 624 0 1 99540
box -42 -55 624 371
use contact_9  contact_9_9
timestamp 1624494425
transform 1 0 351 0 1 100056
box 0 0 66 74
use contact_9  contact_9_8
timestamp 1624494425
transform 1 0 351 0 1 100293
box 0 0 66 74
use contact_9  contact_9_6
timestamp 1624494425
transform 1 0 351 0 1 100293
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_4
timestamp 1624494425
transform -1 0 624 0 1 100330
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_5
timestamp 1624494425
transform -1 0 624 0 -1 100330
box -42 -55 624 371
use contact_9  contact_9_7
timestamp 1624494425
transform 1 0 351 0 1 100530
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_3
timestamp 1624494425
transform -1 0 624 0 -1 101120
box -42 -55 624 371
use contact_9  contact_9_5
timestamp 1624494425
transform 1 0 351 0 1 100846
box 0 0 66 74
use contact_9  contact_9_4
timestamp 1624494425
transform 1 0 351 0 1 101083
box 0 0 66 74
use contact_9  contact_9_2
timestamp 1624494425
transform 1 0 351 0 1 101083
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_2
timestamp 1624494425
transform -1 0 624 0 1 101120
box -42 -55 624 371
use contact_9  contact_9_3
timestamp 1624494425
transform 1 0 351 0 1 101320
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_1
timestamp 1624494425
transform -1 0 624 0 -1 101910
box -42 -55 624 371
use contact_9  contact_9_1
timestamp 1624494425
transform 1 0 351 0 1 101636
box 0 0 66 74
use contact_9  contact_9_0
timestamp 1624494425
transform 1 0 351 0 1 101873
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_row  sky130_fd_bd_sram__openram_dp_cell_cap_row_0
timestamp 1624494425
transform -1 0 624 0 1 101910
box -42 -55 624 371
<< labels >>
rlabel metal2 s 0 1113 28 1161 4 wl0_1
rlabel metal2 s 0 893 28 941 4 wl1_1
rlabel metal2 s 0 1209 28 1257 4 wl0_2
rlabel metal2 s 0 1429 28 1477 4 wl1_2
rlabel metal2 s 0 1903 28 1951 4 wl0_3
rlabel metal2 s 0 1683 28 1731 4 wl1_3
rlabel metal2 s 0 1999 28 2047 4 wl0_4
rlabel metal2 s 0 2219 28 2267 4 wl1_4
rlabel metal2 s 0 2693 28 2741 4 wl0_5
rlabel metal2 s 0 2473 28 2521 4 wl1_5
rlabel metal2 s 0 2789 28 2837 4 wl0_6
rlabel metal2 s 0 3009 28 3057 4 wl1_6
rlabel metal2 s 0 3483 28 3531 4 wl0_7
rlabel metal2 s 0 3263 28 3311 4 wl1_7
rlabel metal2 s 0 3579 28 3627 4 wl0_8
rlabel metal2 s 0 3799 28 3847 4 wl1_8
rlabel metal2 s 0 4273 28 4321 4 wl0_9
rlabel metal2 s 0 4053 28 4101 4 wl1_9
rlabel metal2 s 0 4369 28 4417 4 wl0_10
rlabel metal2 s 0 4589 28 4637 4 wl1_10
rlabel metal2 s 0 5063 28 5111 4 wl0_11
rlabel metal2 s 0 4843 28 4891 4 wl1_11
rlabel metal2 s 0 5159 28 5207 4 wl0_12
rlabel metal2 s 0 5379 28 5427 4 wl1_12
rlabel metal2 s 0 5853 28 5901 4 wl0_13
rlabel metal2 s 0 5633 28 5681 4 wl1_13
rlabel metal2 s 0 5949 28 5997 4 wl0_14
rlabel metal2 s 0 6169 28 6217 4 wl1_14
rlabel metal2 s 0 6643 28 6691 4 wl0_15
rlabel metal2 s 0 6423 28 6471 4 wl1_15
rlabel metal2 s 0 6739 28 6787 4 wl0_16
rlabel metal2 s 0 6959 28 7007 4 wl1_16
rlabel metal2 s 0 7433 28 7481 4 wl0_17
rlabel metal2 s 0 7213 28 7261 4 wl1_17
rlabel metal2 s 0 7529 28 7577 4 wl0_18
rlabel metal2 s 0 7749 28 7797 4 wl1_18
rlabel metal2 s 0 8223 28 8271 4 wl0_19
rlabel metal2 s 0 8003 28 8051 4 wl1_19
rlabel metal2 s 0 8319 28 8367 4 wl0_20
rlabel metal2 s 0 8539 28 8587 4 wl1_20
rlabel metal2 s 0 9013 28 9061 4 wl0_21
rlabel metal2 s 0 8793 28 8841 4 wl1_21
rlabel metal2 s 0 9109 28 9157 4 wl0_22
rlabel metal2 s 0 9329 28 9377 4 wl1_22
rlabel metal2 s 0 9803 28 9851 4 wl0_23
rlabel metal2 s 0 9583 28 9631 4 wl1_23
rlabel metal2 s 0 9899 28 9947 4 wl0_24
rlabel metal2 s 0 10119 28 10167 4 wl1_24
rlabel metal2 s 0 10593 28 10641 4 wl0_25
rlabel metal2 s 0 10373 28 10421 4 wl1_25
rlabel metal2 s 0 10689 28 10737 4 wl0_26
rlabel metal2 s 0 10909 28 10957 4 wl1_26
rlabel metal2 s 0 11383 28 11431 4 wl0_27
rlabel metal2 s 0 11163 28 11211 4 wl1_27
rlabel metal2 s 0 11479 28 11527 4 wl0_28
rlabel metal2 s 0 11699 28 11747 4 wl1_28
rlabel metal2 s 0 12173 28 12221 4 wl0_29
rlabel metal2 s 0 11953 28 12001 4 wl1_29
rlabel metal2 s 0 12269 28 12317 4 wl0_30
rlabel metal2 s 0 12489 28 12537 4 wl1_30
rlabel metal2 s 0 12963 28 13011 4 wl0_31
rlabel metal2 s 0 12743 28 12791 4 wl1_31
rlabel metal2 s 0 13059 28 13107 4 wl0_32
rlabel metal2 s 0 13279 28 13327 4 wl1_32
rlabel metal2 s 0 13753 28 13801 4 wl0_33
rlabel metal2 s 0 13533 28 13581 4 wl1_33
rlabel metal2 s 0 13849 28 13897 4 wl0_34
rlabel metal2 s 0 14069 28 14117 4 wl1_34
rlabel metal2 s 0 14543 28 14591 4 wl0_35
rlabel metal2 s 0 14323 28 14371 4 wl1_35
rlabel metal2 s 0 14639 28 14687 4 wl0_36
rlabel metal2 s 0 14859 28 14907 4 wl1_36
rlabel metal2 s 0 15333 28 15381 4 wl0_37
rlabel metal2 s 0 15113 28 15161 4 wl1_37
rlabel metal2 s 0 15429 28 15477 4 wl0_38
rlabel metal2 s 0 15649 28 15697 4 wl1_38
rlabel metal2 s 0 16123 28 16171 4 wl0_39
rlabel metal2 s 0 15903 28 15951 4 wl1_39
rlabel metal2 s 0 16219 28 16267 4 wl0_40
rlabel metal2 s 0 16439 28 16487 4 wl1_40
rlabel metal2 s 0 16913 28 16961 4 wl0_41
rlabel metal2 s 0 16693 28 16741 4 wl1_41
rlabel metal2 s 0 17009 28 17057 4 wl0_42
rlabel metal2 s 0 17229 28 17277 4 wl1_42
rlabel metal2 s 0 17703 28 17751 4 wl0_43
rlabel metal2 s 0 17483 28 17531 4 wl1_43
rlabel metal2 s 0 17799 28 17847 4 wl0_44
rlabel metal2 s 0 18019 28 18067 4 wl1_44
rlabel metal2 s 0 18493 28 18541 4 wl0_45
rlabel metal2 s 0 18273 28 18321 4 wl1_45
rlabel metal2 s 0 18589 28 18637 4 wl0_46
rlabel metal2 s 0 18809 28 18857 4 wl1_46
rlabel metal2 s 0 19283 28 19331 4 wl0_47
rlabel metal2 s 0 19063 28 19111 4 wl1_47
rlabel metal2 s 0 19379 28 19427 4 wl0_48
rlabel metal2 s 0 19599 28 19647 4 wl1_48
rlabel metal2 s 0 20073 28 20121 4 wl0_49
rlabel metal2 s 0 19853 28 19901 4 wl1_49
rlabel metal2 s 0 20169 28 20217 4 wl0_50
rlabel metal2 s 0 20389 28 20437 4 wl1_50
rlabel metal2 s 0 20863 28 20911 4 wl0_51
rlabel metal2 s 0 20643 28 20691 4 wl1_51
rlabel metal2 s 0 20959 28 21007 4 wl0_52
rlabel metal2 s 0 21179 28 21227 4 wl1_52
rlabel metal2 s 0 21653 28 21701 4 wl0_53
rlabel metal2 s 0 21433 28 21481 4 wl1_53
rlabel metal2 s 0 21749 28 21797 4 wl0_54
rlabel metal2 s 0 21969 28 22017 4 wl1_54
rlabel metal2 s 0 22443 28 22491 4 wl0_55
rlabel metal2 s 0 22223 28 22271 4 wl1_55
rlabel metal2 s 0 22539 28 22587 4 wl0_56
rlabel metal2 s 0 22759 28 22807 4 wl1_56
rlabel metal2 s 0 23233 28 23281 4 wl0_57
rlabel metal2 s 0 23013 28 23061 4 wl1_57
rlabel metal2 s 0 23329 28 23377 4 wl0_58
rlabel metal2 s 0 23549 28 23597 4 wl1_58
rlabel metal2 s 0 24023 28 24071 4 wl0_59
rlabel metal2 s 0 23803 28 23851 4 wl1_59
rlabel metal2 s 0 24119 28 24167 4 wl0_60
rlabel metal2 s 0 24339 28 24387 4 wl1_60
rlabel metal2 s 0 24813 28 24861 4 wl0_61
rlabel metal2 s 0 24593 28 24641 4 wl1_61
rlabel metal2 s 0 24909 28 24957 4 wl0_62
rlabel metal2 s 0 25129 28 25177 4 wl1_62
rlabel metal2 s 0 25603 28 25651 4 wl0_63
rlabel metal2 s 0 25383 28 25431 4 wl1_63
rlabel metal2 s 0 25699 28 25747 4 wl0_64
rlabel metal2 s 0 25919 28 25967 4 wl1_64
rlabel metal2 s 0 26393 28 26441 4 wl0_65
rlabel metal2 s 0 26173 28 26221 4 wl1_65
rlabel metal2 s 0 26489 28 26537 4 wl0_66
rlabel metal2 s 0 26709 28 26757 4 wl1_66
rlabel metal2 s 0 27183 28 27231 4 wl0_67
rlabel metal2 s 0 26963 28 27011 4 wl1_67
rlabel metal2 s 0 27279 28 27327 4 wl0_68
rlabel metal2 s 0 27499 28 27547 4 wl1_68
rlabel metal2 s 0 27973 28 28021 4 wl0_69
rlabel metal2 s 0 27753 28 27801 4 wl1_69
rlabel metal2 s 0 28069 28 28117 4 wl0_70
rlabel metal2 s 0 28289 28 28337 4 wl1_70
rlabel metal2 s 0 28763 28 28811 4 wl0_71
rlabel metal2 s 0 28543 28 28591 4 wl1_71
rlabel metal2 s 0 28859 28 28907 4 wl0_72
rlabel metal2 s 0 29079 28 29127 4 wl1_72
rlabel metal2 s 0 29553 28 29601 4 wl0_73
rlabel metal2 s 0 29333 28 29381 4 wl1_73
rlabel metal2 s 0 29649 28 29697 4 wl0_74
rlabel metal2 s 0 29869 28 29917 4 wl1_74
rlabel metal2 s 0 30343 28 30391 4 wl0_75
rlabel metal2 s 0 30123 28 30171 4 wl1_75
rlabel metal2 s 0 30439 28 30487 4 wl0_76
rlabel metal2 s 0 30659 28 30707 4 wl1_76
rlabel metal2 s 0 31133 28 31181 4 wl0_77
rlabel metal2 s 0 30913 28 30961 4 wl1_77
rlabel metal2 s 0 31229 28 31277 4 wl0_78
rlabel metal2 s 0 31449 28 31497 4 wl1_78
rlabel metal2 s 0 31923 28 31971 4 wl0_79
rlabel metal2 s 0 31703 28 31751 4 wl1_79
rlabel metal2 s 0 32019 28 32067 4 wl0_80
rlabel metal2 s 0 32239 28 32287 4 wl1_80
rlabel metal2 s 0 32713 28 32761 4 wl0_81
rlabel metal2 s 0 32493 28 32541 4 wl1_81
rlabel metal2 s 0 32809 28 32857 4 wl0_82
rlabel metal2 s 0 33029 28 33077 4 wl1_82
rlabel metal2 s 0 33503 28 33551 4 wl0_83
rlabel metal2 s 0 33283 28 33331 4 wl1_83
rlabel metal2 s 0 33599 28 33647 4 wl0_84
rlabel metal2 s 0 33819 28 33867 4 wl1_84
rlabel metal2 s 0 34293 28 34341 4 wl0_85
rlabel metal2 s 0 34073 28 34121 4 wl1_85
rlabel metal2 s 0 34389 28 34437 4 wl0_86
rlabel metal2 s 0 34609 28 34657 4 wl1_86
rlabel metal2 s 0 35083 28 35131 4 wl0_87
rlabel metal2 s 0 34863 28 34911 4 wl1_87
rlabel metal2 s 0 35179 28 35227 4 wl0_88
rlabel metal2 s 0 35399 28 35447 4 wl1_88
rlabel metal2 s 0 35873 28 35921 4 wl0_89
rlabel metal2 s 0 35653 28 35701 4 wl1_89
rlabel metal2 s 0 35969 28 36017 4 wl0_90
rlabel metal2 s 0 36189 28 36237 4 wl1_90
rlabel metal2 s 0 36663 28 36711 4 wl0_91
rlabel metal2 s 0 36443 28 36491 4 wl1_91
rlabel metal2 s 0 36759 28 36807 4 wl0_92
rlabel metal2 s 0 36979 28 37027 4 wl1_92
rlabel metal2 s 0 37453 28 37501 4 wl0_93
rlabel metal2 s 0 37233 28 37281 4 wl1_93
rlabel metal2 s 0 37549 28 37597 4 wl0_94
rlabel metal2 s 0 37769 28 37817 4 wl1_94
rlabel metal2 s 0 38243 28 38291 4 wl0_95
rlabel metal2 s 0 38023 28 38071 4 wl1_95
rlabel metal2 s 0 38339 28 38387 4 wl0_96
rlabel metal2 s 0 38559 28 38607 4 wl1_96
rlabel metal2 s 0 39033 28 39081 4 wl0_97
rlabel metal2 s 0 38813 28 38861 4 wl1_97
rlabel metal2 s 0 39129 28 39177 4 wl0_98
rlabel metal2 s 0 39349 28 39397 4 wl1_98
rlabel metal2 s 0 39823 28 39871 4 wl0_99
rlabel metal2 s 0 39603 28 39651 4 wl1_99
rlabel metal2 s 0 39919 28 39967 4 wl0_100
rlabel metal2 s 0 40139 28 40187 4 wl1_100
rlabel metal2 s 0 40613 28 40661 4 wl0_101
rlabel metal2 s 0 40393 28 40441 4 wl1_101
rlabel metal2 s 0 40709 28 40757 4 wl0_102
rlabel metal2 s 0 40929 28 40977 4 wl1_102
rlabel metal2 s 0 41403 28 41451 4 wl0_103
rlabel metal2 s 0 41183 28 41231 4 wl1_103
rlabel metal2 s 0 41499 28 41547 4 wl0_104
rlabel metal2 s 0 41719 28 41767 4 wl1_104
rlabel metal2 s 0 42193 28 42241 4 wl0_105
rlabel metal2 s 0 41973 28 42021 4 wl1_105
rlabel metal2 s 0 42289 28 42337 4 wl0_106
rlabel metal2 s 0 42509 28 42557 4 wl1_106
rlabel metal2 s 0 42983 28 43031 4 wl0_107
rlabel metal2 s 0 42763 28 42811 4 wl1_107
rlabel metal2 s 0 43079 28 43127 4 wl0_108
rlabel metal2 s 0 43299 28 43347 4 wl1_108
rlabel metal2 s 0 43773 28 43821 4 wl0_109
rlabel metal2 s 0 43553 28 43601 4 wl1_109
rlabel metal2 s 0 43869 28 43917 4 wl0_110
rlabel metal2 s 0 44089 28 44137 4 wl1_110
rlabel metal2 s 0 44563 28 44611 4 wl0_111
rlabel metal2 s 0 44343 28 44391 4 wl1_111
rlabel metal2 s 0 44659 28 44707 4 wl0_112
rlabel metal2 s 0 44879 28 44927 4 wl1_112
rlabel metal2 s 0 45353 28 45401 4 wl0_113
rlabel metal2 s 0 45133 28 45181 4 wl1_113
rlabel metal2 s 0 45449 28 45497 4 wl0_114
rlabel metal2 s 0 45669 28 45717 4 wl1_114
rlabel metal2 s 0 46143 28 46191 4 wl0_115
rlabel metal2 s 0 45923 28 45971 4 wl1_115
rlabel metal2 s 0 46239 28 46287 4 wl0_116
rlabel metal2 s 0 46459 28 46507 4 wl1_116
rlabel metal2 s 0 46933 28 46981 4 wl0_117
rlabel metal2 s 0 46713 28 46761 4 wl1_117
rlabel metal2 s 0 47029 28 47077 4 wl0_118
rlabel metal2 s 0 47249 28 47297 4 wl1_118
rlabel metal2 s 0 47723 28 47771 4 wl0_119
rlabel metal2 s 0 47503 28 47551 4 wl1_119
rlabel metal2 s 0 47819 28 47867 4 wl0_120
rlabel metal2 s 0 48039 28 48087 4 wl1_120
rlabel metal2 s 0 48513 28 48561 4 wl0_121
rlabel metal2 s 0 48293 28 48341 4 wl1_121
rlabel metal2 s 0 48609 28 48657 4 wl0_122
rlabel metal2 s 0 48829 28 48877 4 wl1_122
rlabel metal2 s 0 49303 28 49351 4 wl0_123
rlabel metal2 s 0 49083 28 49131 4 wl1_123
rlabel metal2 s 0 49399 28 49447 4 wl0_124
rlabel metal2 s 0 49619 28 49667 4 wl1_124
rlabel metal2 s 0 50093 28 50141 4 wl0_125
rlabel metal2 s 0 49873 28 49921 4 wl1_125
rlabel metal2 s 0 50189 28 50237 4 wl0_126
rlabel metal2 s 0 50409 28 50457 4 wl1_126
rlabel metal2 s 0 50883 28 50931 4 wl0_127
rlabel metal2 s 0 50663 28 50711 4 wl1_127
rlabel metal2 s 0 50979 28 51027 4 wl0_128
rlabel metal2 s 0 51199 28 51247 4 wl1_128
rlabel metal2 s 0 51673 28 51721 4 wl0_129
rlabel metal2 s 0 51453 28 51501 4 wl1_129
rlabel metal2 s 0 51769 28 51817 4 wl0_130
rlabel metal2 s 0 51989 28 52037 4 wl1_130
rlabel metal2 s 0 52463 28 52511 4 wl0_131
rlabel metal2 s 0 52243 28 52291 4 wl1_131
rlabel metal2 s 0 52559 28 52607 4 wl0_132
rlabel metal2 s 0 52779 28 52827 4 wl1_132
rlabel metal2 s 0 53253 28 53301 4 wl0_133
rlabel metal2 s 0 53033 28 53081 4 wl1_133
rlabel metal2 s 0 53349 28 53397 4 wl0_134
rlabel metal2 s 0 53569 28 53617 4 wl1_134
rlabel metal2 s 0 54043 28 54091 4 wl0_135
rlabel metal2 s 0 53823 28 53871 4 wl1_135
rlabel metal2 s 0 54139 28 54187 4 wl0_136
rlabel metal2 s 0 54359 28 54407 4 wl1_136
rlabel metal2 s 0 54833 28 54881 4 wl0_137
rlabel metal2 s 0 54613 28 54661 4 wl1_137
rlabel metal2 s 0 54929 28 54977 4 wl0_138
rlabel metal2 s 0 55149 28 55197 4 wl1_138
rlabel metal2 s 0 55623 28 55671 4 wl0_139
rlabel metal2 s 0 55403 28 55451 4 wl1_139
rlabel metal2 s 0 55719 28 55767 4 wl0_140
rlabel metal2 s 0 55939 28 55987 4 wl1_140
rlabel metal2 s 0 56413 28 56461 4 wl0_141
rlabel metal2 s 0 56193 28 56241 4 wl1_141
rlabel metal2 s 0 56509 28 56557 4 wl0_142
rlabel metal2 s 0 56729 28 56777 4 wl1_142
rlabel metal2 s 0 57203 28 57251 4 wl0_143
rlabel metal2 s 0 56983 28 57031 4 wl1_143
rlabel metal2 s 0 57299 28 57347 4 wl0_144
rlabel metal2 s 0 57519 28 57567 4 wl1_144
rlabel metal2 s 0 57993 28 58041 4 wl0_145
rlabel metal2 s 0 57773 28 57821 4 wl1_145
rlabel metal2 s 0 58089 28 58137 4 wl0_146
rlabel metal2 s 0 58309 28 58357 4 wl1_146
rlabel metal2 s 0 58783 28 58831 4 wl0_147
rlabel metal2 s 0 58563 28 58611 4 wl1_147
rlabel metal2 s 0 58879 28 58927 4 wl0_148
rlabel metal2 s 0 59099 28 59147 4 wl1_148
rlabel metal2 s 0 59573 28 59621 4 wl0_149
rlabel metal2 s 0 59353 28 59401 4 wl1_149
rlabel metal2 s 0 59669 28 59717 4 wl0_150
rlabel metal2 s 0 59889 28 59937 4 wl1_150
rlabel metal2 s 0 60363 28 60411 4 wl0_151
rlabel metal2 s 0 60143 28 60191 4 wl1_151
rlabel metal2 s 0 60459 28 60507 4 wl0_152
rlabel metal2 s 0 60679 28 60727 4 wl1_152
rlabel metal2 s 0 61153 28 61201 4 wl0_153
rlabel metal2 s 0 60933 28 60981 4 wl1_153
rlabel metal2 s 0 61249 28 61297 4 wl0_154
rlabel metal2 s 0 61469 28 61517 4 wl1_154
rlabel metal2 s 0 61943 28 61991 4 wl0_155
rlabel metal2 s 0 61723 28 61771 4 wl1_155
rlabel metal2 s 0 62039 28 62087 4 wl0_156
rlabel metal2 s 0 62259 28 62307 4 wl1_156
rlabel metal2 s 0 62733 28 62781 4 wl0_157
rlabel metal2 s 0 62513 28 62561 4 wl1_157
rlabel metal2 s 0 62829 28 62877 4 wl0_158
rlabel metal2 s 0 63049 28 63097 4 wl1_158
rlabel metal2 s 0 63523 28 63571 4 wl0_159
rlabel metal2 s 0 63303 28 63351 4 wl1_159
rlabel metal2 s 0 63619 28 63667 4 wl0_160
rlabel metal2 s 0 63839 28 63887 4 wl1_160
rlabel metal2 s 0 64313 28 64361 4 wl0_161
rlabel metal2 s 0 64093 28 64141 4 wl1_161
rlabel metal2 s 0 64409 28 64457 4 wl0_162
rlabel metal2 s 0 64629 28 64677 4 wl1_162
rlabel metal2 s 0 65103 28 65151 4 wl0_163
rlabel metal2 s 0 64883 28 64931 4 wl1_163
rlabel metal2 s 0 65199 28 65247 4 wl0_164
rlabel metal2 s 0 65419 28 65467 4 wl1_164
rlabel metal2 s 0 65893 28 65941 4 wl0_165
rlabel metal2 s 0 65673 28 65721 4 wl1_165
rlabel metal2 s 0 65989 28 66037 4 wl0_166
rlabel metal2 s 0 66209 28 66257 4 wl1_166
rlabel metal2 s 0 66683 28 66731 4 wl0_167
rlabel metal2 s 0 66463 28 66511 4 wl1_167
rlabel metal2 s 0 66779 28 66827 4 wl0_168
rlabel metal2 s 0 66999 28 67047 4 wl1_168
rlabel metal2 s 0 67473 28 67521 4 wl0_169
rlabel metal2 s 0 67253 28 67301 4 wl1_169
rlabel metal2 s 0 67569 28 67617 4 wl0_170
rlabel metal2 s 0 67789 28 67837 4 wl1_170
rlabel metal2 s 0 68263 28 68311 4 wl0_171
rlabel metal2 s 0 68043 28 68091 4 wl1_171
rlabel metal2 s 0 68359 28 68407 4 wl0_172
rlabel metal2 s 0 68579 28 68627 4 wl1_172
rlabel metal2 s 0 69053 28 69101 4 wl0_173
rlabel metal2 s 0 68833 28 68881 4 wl1_173
rlabel metal2 s 0 69149 28 69197 4 wl0_174
rlabel metal2 s 0 69369 28 69417 4 wl1_174
rlabel metal2 s 0 69843 28 69891 4 wl0_175
rlabel metal2 s 0 69623 28 69671 4 wl1_175
rlabel metal2 s 0 69939 28 69987 4 wl0_176
rlabel metal2 s 0 70159 28 70207 4 wl1_176
rlabel metal2 s 0 70633 28 70681 4 wl0_177
rlabel metal2 s 0 70413 28 70461 4 wl1_177
rlabel metal2 s 0 70729 28 70777 4 wl0_178
rlabel metal2 s 0 70949 28 70997 4 wl1_178
rlabel metal2 s 0 71423 28 71471 4 wl0_179
rlabel metal2 s 0 71203 28 71251 4 wl1_179
rlabel metal2 s 0 71519 28 71567 4 wl0_180
rlabel metal2 s 0 71739 28 71787 4 wl1_180
rlabel metal2 s 0 72213 28 72261 4 wl0_181
rlabel metal2 s 0 71993 28 72041 4 wl1_181
rlabel metal2 s 0 72309 28 72357 4 wl0_182
rlabel metal2 s 0 72529 28 72577 4 wl1_182
rlabel metal2 s 0 73003 28 73051 4 wl0_183
rlabel metal2 s 0 72783 28 72831 4 wl1_183
rlabel metal2 s 0 73099 28 73147 4 wl0_184
rlabel metal2 s 0 73319 28 73367 4 wl1_184
rlabel metal2 s 0 73793 28 73841 4 wl0_185
rlabel metal2 s 0 73573 28 73621 4 wl1_185
rlabel metal2 s 0 73889 28 73937 4 wl0_186
rlabel metal2 s 0 74109 28 74157 4 wl1_186
rlabel metal2 s 0 74583 28 74631 4 wl0_187
rlabel metal2 s 0 74363 28 74411 4 wl1_187
rlabel metal2 s 0 74679 28 74727 4 wl0_188
rlabel metal2 s 0 74899 28 74947 4 wl1_188
rlabel metal2 s 0 75373 28 75421 4 wl0_189
rlabel metal2 s 0 75153 28 75201 4 wl1_189
rlabel metal2 s 0 75469 28 75517 4 wl0_190
rlabel metal2 s 0 75689 28 75737 4 wl1_190
rlabel metal2 s 0 76163 28 76211 4 wl0_191
rlabel metal2 s 0 75943 28 75991 4 wl1_191
rlabel metal2 s 0 76259 28 76307 4 wl0_192
rlabel metal2 s 0 76479 28 76527 4 wl1_192
rlabel metal2 s 0 76953 28 77001 4 wl0_193
rlabel metal2 s 0 76733 28 76781 4 wl1_193
rlabel metal2 s 0 77049 28 77097 4 wl0_194
rlabel metal2 s 0 77269 28 77317 4 wl1_194
rlabel metal2 s 0 77743 28 77791 4 wl0_195
rlabel metal2 s 0 77523 28 77571 4 wl1_195
rlabel metal2 s 0 77839 28 77887 4 wl0_196
rlabel metal2 s 0 78059 28 78107 4 wl1_196
rlabel metal2 s 0 78533 28 78581 4 wl0_197
rlabel metal2 s 0 78313 28 78361 4 wl1_197
rlabel metal2 s 0 78629 28 78677 4 wl0_198
rlabel metal2 s 0 78849 28 78897 4 wl1_198
rlabel metal2 s 0 79323 28 79371 4 wl0_199
rlabel metal2 s 0 79103 28 79151 4 wl1_199
rlabel metal2 s 0 79419 28 79467 4 wl0_200
rlabel metal2 s 0 79639 28 79687 4 wl1_200
rlabel metal2 s 0 80113 28 80161 4 wl0_201
rlabel metal2 s 0 79893 28 79941 4 wl1_201
rlabel metal2 s 0 80209 28 80257 4 wl0_202
rlabel metal2 s 0 80429 28 80477 4 wl1_202
rlabel metal2 s 0 80903 28 80951 4 wl0_203
rlabel metal2 s 0 80683 28 80731 4 wl1_203
rlabel metal2 s 0 80999 28 81047 4 wl0_204
rlabel metal2 s 0 81219 28 81267 4 wl1_204
rlabel metal2 s 0 81693 28 81741 4 wl0_205
rlabel metal2 s 0 81473 28 81521 4 wl1_205
rlabel metal2 s 0 81789 28 81837 4 wl0_206
rlabel metal2 s 0 82009 28 82057 4 wl1_206
rlabel metal2 s 0 82483 28 82531 4 wl0_207
rlabel metal2 s 0 82263 28 82311 4 wl1_207
rlabel metal2 s 0 82579 28 82627 4 wl0_208
rlabel metal2 s 0 82799 28 82847 4 wl1_208
rlabel metal2 s 0 83273 28 83321 4 wl0_209
rlabel metal2 s 0 83053 28 83101 4 wl1_209
rlabel metal2 s 0 83369 28 83417 4 wl0_210
rlabel metal2 s 0 83589 28 83637 4 wl1_210
rlabel metal2 s 0 84063 28 84111 4 wl0_211
rlabel metal2 s 0 83843 28 83891 4 wl1_211
rlabel metal2 s 0 84159 28 84207 4 wl0_212
rlabel metal2 s 0 84379 28 84427 4 wl1_212
rlabel metal2 s 0 84853 28 84901 4 wl0_213
rlabel metal2 s 0 84633 28 84681 4 wl1_213
rlabel metal2 s 0 84949 28 84997 4 wl0_214
rlabel metal2 s 0 85169 28 85217 4 wl1_214
rlabel metal2 s 0 85643 28 85691 4 wl0_215
rlabel metal2 s 0 85423 28 85471 4 wl1_215
rlabel metal2 s 0 85739 28 85787 4 wl0_216
rlabel metal2 s 0 85959 28 86007 4 wl1_216
rlabel metal2 s 0 86433 28 86481 4 wl0_217
rlabel metal2 s 0 86213 28 86261 4 wl1_217
rlabel metal2 s 0 86529 28 86577 4 wl0_218
rlabel metal2 s 0 86749 28 86797 4 wl1_218
rlabel metal2 s 0 87223 28 87271 4 wl0_219
rlabel metal2 s 0 87003 28 87051 4 wl1_219
rlabel metal2 s 0 87319 28 87367 4 wl0_220
rlabel metal2 s 0 87539 28 87587 4 wl1_220
rlabel metal2 s 0 88013 28 88061 4 wl0_221
rlabel metal2 s 0 87793 28 87841 4 wl1_221
rlabel metal2 s 0 88109 28 88157 4 wl0_222
rlabel metal2 s 0 88329 28 88377 4 wl1_222
rlabel metal2 s 0 88803 28 88851 4 wl0_223
rlabel metal2 s 0 88583 28 88631 4 wl1_223
rlabel metal2 s 0 88899 28 88947 4 wl0_224
rlabel metal2 s 0 89119 28 89167 4 wl1_224
rlabel metal2 s 0 89593 28 89641 4 wl0_225
rlabel metal2 s 0 89373 28 89421 4 wl1_225
rlabel metal2 s 0 89689 28 89737 4 wl0_226
rlabel metal2 s 0 89909 28 89957 4 wl1_226
rlabel metal2 s 0 90383 28 90431 4 wl0_227
rlabel metal2 s 0 90163 28 90211 4 wl1_227
rlabel metal2 s 0 90479 28 90527 4 wl0_228
rlabel metal2 s 0 90699 28 90747 4 wl1_228
rlabel metal2 s 0 91173 28 91221 4 wl0_229
rlabel metal2 s 0 90953 28 91001 4 wl1_229
rlabel metal2 s 0 91269 28 91317 4 wl0_230
rlabel metal2 s 0 91489 28 91537 4 wl1_230
rlabel metal2 s 0 91963 28 92011 4 wl0_231
rlabel metal2 s 0 91743 28 91791 4 wl1_231
rlabel metal2 s 0 92059 28 92107 4 wl0_232
rlabel metal2 s 0 92279 28 92327 4 wl1_232
rlabel metal2 s 0 92753 28 92801 4 wl0_233
rlabel metal2 s 0 92533 28 92581 4 wl1_233
rlabel metal2 s 0 92849 28 92897 4 wl0_234
rlabel metal2 s 0 93069 28 93117 4 wl1_234
rlabel metal2 s 0 93543 28 93591 4 wl0_235
rlabel metal2 s 0 93323 28 93371 4 wl1_235
rlabel metal2 s 0 93639 28 93687 4 wl0_236
rlabel metal2 s 0 93859 28 93907 4 wl1_236
rlabel metal2 s 0 94333 28 94381 4 wl0_237
rlabel metal2 s 0 94113 28 94161 4 wl1_237
rlabel metal2 s 0 94429 28 94477 4 wl0_238
rlabel metal2 s 0 94649 28 94697 4 wl1_238
rlabel metal2 s 0 95123 28 95171 4 wl0_239
rlabel metal2 s 0 94903 28 94951 4 wl1_239
rlabel metal2 s 0 95219 28 95267 4 wl0_240
rlabel metal2 s 0 95439 28 95487 4 wl1_240
rlabel metal2 s 0 95913 28 95961 4 wl0_241
rlabel metal2 s 0 95693 28 95741 4 wl1_241
rlabel metal2 s 0 96009 28 96057 4 wl0_242
rlabel metal2 s 0 96229 28 96277 4 wl1_242
rlabel metal2 s 0 96703 28 96751 4 wl0_243
rlabel metal2 s 0 96483 28 96531 4 wl1_243
rlabel metal2 s 0 96799 28 96847 4 wl0_244
rlabel metal2 s 0 97019 28 97067 4 wl1_244
rlabel metal2 s 0 97493 28 97541 4 wl0_245
rlabel metal2 s 0 97273 28 97321 4 wl1_245
rlabel metal2 s 0 97589 28 97637 4 wl0_246
rlabel metal2 s 0 97809 28 97857 4 wl1_246
rlabel metal2 s 0 98283 28 98331 4 wl0_247
rlabel metal2 s 0 98063 28 98111 4 wl1_247
rlabel metal2 s 0 98379 28 98427 4 wl0_248
rlabel metal2 s 0 98599 28 98647 4 wl1_248
rlabel metal2 s 0 99073 28 99121 4 wl0_249
rlabel metal2 s 0 98853 28 98901 4 wl1_249
rlabel metal2 s 0 99169 28 99217 4 wl0_250
rlabel metal2 s 0 99389 28 99437 4 wl1_250
rlabel metal2 s 0 99863 28 99911 4 wl0_251
rlabel metal2 s 0 99643 28 99691 4 wl1_251
rlabel metal2 s 0 99959 28 100007 4 wl0_252
rlabel metal2 s 0 100179 28 100227 4 wl1_252
rlabel metal2 s 0 100653 28 100701 4 wl0_253
rlabel metal2 s 0 100433 28 100481 4 wl1_253
rlabel metal2 s 0 100749 28 100797 4 wl0_254
rlabel metal2 s 0 100969 28 101017 4 wl1_254
rlabel metal2 s 0 101443 28 101491 4 wl0_255
rlabel metal2 s 0 101223 28 101271 4 wl1_255
rlabel metal2 s 0 101539 28 101587 4 wl0_256
rlabel metal2 s 0 101759 28 101807 4 wl1_256
rlabel metal3 s 335 24994 433 25092 4 gnd
rlabel metal3 s 335 45534 433 45632 4 gnd
rlabel metal3 s 335 9194 433 9292 4 gnd
rlabel metal3 s 335 47114 433 47212 4 gnd
rlabel metal3 s 335 68918 433 69016 4 gnd
rlabel metal3 s 335 83928 433 84026 4 gnd
rlabel metal3 s 335 66074 433 66172 4 gnd
rlabel metal3 s 335 65284 433 65382 4 gnd
rlabel metal3 s 335 60544 433 60642 4 gnd
rlabel metal3 s 335 68444 433 68542 4 gnd
rlabel metal3 s 335 81321 433 81419 4 gnd
rlabel metal3 s 335 8878 433 8976 4 gnd
rlabel metal3 s 335 73421 433 73519 4 gnd
rlabel metal3 s 335 18358 433 18456 4 gnd
rlabel metal3 s 335 97121 433 97219 4 gnd
rlabel metal3 s 335 19148 433 19246 4 gnd
rlabel metal3 s 335 64968 433 65066 4 gnd
rlabel metal3 s 335 6824 433 6922 4 gnd
rlabel metal3 s 335 16304 433 16402 4 gnd
rlabel metal3 s 335 20254 433 20352 4 gnd
rlabel metal3 s 335 28944 433 29042 4 gnd
rlabel metal3 s 335 66864 433 66962 4 gnd
rlabel metal3 s 335 22861 433 22959 4 gnd
rlabel metal3 s 335 48694 433 48792 4 gnd
rlabel metal3 s 335 46798 433 46896 4 gnd
rlabel metal3 s 335 83691 433 83789 4 gnd
rlabel metal3 s 335 98701 433 98799 4 gnd
rlabel metal3 s 335 10221 433 10319 4 gnd
rlabel metal3 s 335 63704 433 63802 4 gnd
rlabel metal3 s 335 49168 433 49266 4 gnd
rlabel metal3 s 335 61334 433 61432 4 gnd
rlabel metal3 s 335 38661 433 38759 4 gnd
rlabel metal3 s 335 49484 433 49582 4 gnd
rlabel metal3 s 335 28628 433 28726 4 gnd
rlabel metal3 s 335 14408 433 14506 4 gnd
rlabel metal3 s 335 72394 433 72492 4 gnd
rlabel metal3 s 335 92934 433 93032 4 gnd
rlabel metal3 s 335 32578 433 32676 4 gnd
rlabel metal3 s 335 83138 433 83236 4 gnd
rlabel metal3 s 335 10774 433 10872 4 gnd
rlabel metal3 s 335 39688 433 39786 4 gnd
rlabel metal3 s 335 40794 433 40892 4 gnd
rlabel metal3 s 335 74448 433 74546 4 gnd
rlabel metal3 s 335 3111 433 3209 4 gnd
rlabel metal3 s 335 7061 433 7159 4 gnd
rlabel metal3 s 335 97674 433 97772 4 gnd
rlabel metal3 s 335 76028 433 76126 4 gnd
rlabel metal3 s 335 18674 433 18772 4 gnd
rlabel metal3 s 335 80531 433 80629 4 gnd
rlabel metal3 s 335 57384 433 57482 4 gnd
rlabel metal3 s 335 67101 433 67199 4 gnd
rlabel metal3 s 335 86061 433 86159 4 gnd
rlabel metal3 s 335 81874 433 81972 4 gnd
rlabel metal3 s 335 1294 433 1392 4 gnd
rlabel metal3 s 335 16541 433 16639 4 gnd
rlabel metal3 s 335 75791 433 75889 4 gnd
rlabel metal3 s 335 96568 433 96666 4 gnd
rlabel metal3 s 335 54224 433 54322 4 gnd
rlabel metal3 s 335 50274 433 50372 4 gnd
rlabel metal3 s 335 61808 433 61906 4 gnd
rlabel metal3 s 335 77924 433 78022 4 gnd
rlabel metal3 s 335 32894 433 32992 4 gnd
rlabel metal3 s 335 14171 433 14269 4 gnd
rlabel metal3 s 335 93171 433 93269 4 gnd
rlabel metal3 s 335 31788 433 31886 4 gnd
rlabel metal3 s 335 52881 433 52979 4 gnd
rlabel metal3 s 335 34158 433 34256 4 gnd
rlabel metal3 s 335 98148 433 98246 4 gnd
rlabel metal3 s 335 13934 433 14032 4 gnd
rlabel metal3 s 335 94988 433 95086 4 gnd
rlabel metal3 s 335 34474 433 34572 4 gnd
rlabel metal3 s 335 88984 433 89082 4 gnd
rlabel metal3 s 335 67891 433 67989 4 gnd
rlabel metal3 s 335 21834 433 21932 4 gnd
rlabel metal3 s 335 64731 433 64829 4 gnd
rlabel metal3 s 335 82348 433 82446 4 gnd
rlabel metal3 s 335 82664 433 82762 4 gnd
rlabel metal3 s 335 2321 433 2419 4 gnd
rlabel metal3 s 335 21044 433 21142 4 gnd
rlabel metal3 s 335 66548 433 66646 4 gnd
rlabel metal3 s 335 28154 433 28252 4 gnd
rlabel metal3 s 335 88431 433 88529 4 gnd
rlabel metal3 s 335 34711 433 34809 4 gnd
rlabel metal3 s 335 9431 433 9529 4 gnd
rlabel metal3 s 335 75001 433 75099 4 gnd
rlabel metal3 s 335 70498 433 70596 4 gnd
rlabel metal3 s 335 65521 433 65619 4 gnd
rlabel metal3 s 335 59438 433 59536 4 gnd
rlabel metal3 s 335 50748 433 50846 4 gnd
rlabel metal3 s 335 57621 433 57719 4 gnd
rlabel metal3 s 335 81558 433 81656 4 gnd
rlabel metal3 s 335 12354 433 12452 4 gnd
rlabel metal3 s 335 51854 433 51952 4 gnd
rlabel metal3 s 335 69234 433 69332 4 gnd
rlabel metal3 s 335 53118 433 53216 4 gnd
rlabel metal3 s 335 41268 433 41366 4 gnd
rlabel metal3 s 335 56278 433 56376 4 gnd
rlabel metal3 s 335 18121 433 18219 4 gnd
rlabel metal3 s 335 57858 433 57956 4 gnd
rlabel metal3 s 335 40241 433 40339 4 gnd
rlabel metal3 s 335 40004 433 40102 4 gnd
rlabel metal3 s 335 68681 433 68779 4 gnd
rlabel metal3 s 335 88194 433 88292 4 gnd
rlabel metal3 s 335 22624 433 22722 4 gnd
rlabel metal3 s 335 58174 433 58272 4 gnd
rlabel metal3 s 335 3901 433 3999 4 gnd
rlabel metal3 s 335 13618 433 13716 4 gnd
rlabel metal3 s 335 5481 433 5579 4 gnd
rlabel metal3 s 335 24204 433 24302 4 gnd
rlabel metal3 s 335 62914 433 63012 4 gnd
rlabel metal3 s 335 3664 433 3762 4 gnd
rlabel metal3 s 335 87641 433 87739 4 gnd
rlabel metal3 s 335 6271 433 6369 4 gnd
rlabel metal3 s 335 42058 433 42156 4 gnd
rlabel metal3 s 335 25468 433 25566 4 gnd
rlabel metal3 s 335 48378 433 48476 4 gnd
rlabel metal3 s 335 99491 433 99589 4 gnd
rlabel metal3 s 335 37634 433 37732 4 gnd
rlabel metal3 s 335 19938 433 20036 4 gnd
rlabel metal3 s 335 65758 433 65856 4 gnd
rlabel metal3 s 335 64494 433 64592 4 gnd
rlabel metal3 s 335 98464 433 98562 4 gnd
rlabel metal3 s 335 12038 433 12136 4 gnd
rlabel metal3 s 335 47904 433 48002 4 gnd
rlabel metal3 s 335 6508 433 6606 4 gnd
rlabel metal3 s 335 47351 433 47449 4 gnd
rlabel metal3 s 335 27838 433 27936 4 gnd
rlabel metal3 s 335 26811 433 26909 4 gnd
rlabel metal3 s 335 7851 433 7949 4 gnd
rlabel metal3 s 335 5718 433 5816 4 gnd
rlabel metal3 s 335 978 433 1076 4 gnd
rlabel metal3 s 335 90801 433 90899 4 gnd
rlabel metal3 s 335 59754 433 59852 4 gnd
rlabel metal3 s 335 25231 433 25329 4 gnd
rlabel metal3 s 335 14961 433 15059 4 gnd
rlabel metal3 s 335 53434 433 53532 4 gnd
rlabel metal3 s 335 18911 433 19009 4 gnd
rlabel metal3 s 335 23888 433 23986 4 gnd
rlabel metal3 s 335 15988 433 16086 4 gnd
rlabel metal3 s 335 25784 433 25882 4 gnd
rlabel metal3 s 335 49958 433 50056 4 gnd
rlabel metal3 s 335 3348 433 3446 4 gnd
rlabel metal3 s 335 45771 433 45869 4 gnd
rlabel metal3 s 335 100281 433 100379 4 gnd
rlabel metal3 s 335 52091 433 52189 4 gnd
rlabel metal3 s 335 86851 433 86949 4 gnd
rlabel metal3 s 335 13144 433 13242 4 gnd
rlabel metal3 s 335 75238 433 75336 4 gnd
rlabel metal3 s 335 41031 433 41129 4 gnd
rlabel metal3 s 335 87878 433 87976 4 gnd
rlabel metal3 s 335 11011 433 11109 4 gnd
rlabel metal3 s 335 46561 433 46659 4 gnd
rlabel metal3 s 335 68128 433 68226 4 gnd
rlabel metal3 s 335 60781 433 60879 4 gnd
rlabel metal3 s 335 94198 433 94296 4 gnd
rlabel metal3 s 335 19701 433 19799 4 gnd
rlabel metal3 s 335 17568 433 17666 4 gnd
rlabel metal3 s 335 38898 433 38996 4 gnd
rlabel metal3 s 335 44981 433 45079 4 gnd
rlabel metal3 s 335 1768 433 1866 4 gnd
rlabel metal3 s 335 56041 433 56139 4 gnd
rlabel metal3 s 335 80294 433 80392 4 gnd
rlabel metal3 s 335 50511 433 50609 4 gnd
rlabel metal3 s 335 26021 433 26119 4 gnd
rlabel metal3 s 335 31314 433 31412 4 gnd
rlabel metal3 s 335 33921 433 34019 4 gnd
rlabel metal3 s 335 92381 433 92479 4 gnd
rlabel metal3 s 335 85508 433 85606 4 gnd
rlabel metal3 s 335 101861 433 101959 4 gnd
rlabel metal3 s 335 5244 433 5342 4 gnd
rlabel metal3 s 335 35264 433 35362 4 gnd
rlabel metal3 s 335 66311 433 66409 4 gnd
rlabel metal3 s 335 95541 433 95639 4 gnd
rlabel metal3 s 335 87404 433 87502 4 gnd
rlabel metal3 s 335 7298 433 7396 4 gnd
rlabel metal3 s 335 37871 433 37969 4 gnd
rlabel metal3 s 335 14724 433 14822 4 gnd
rlabel metal3 s 335 27364 433 27462 4 gnd
rlabel metal3 s 335 97358 433 97456 4 gnd
rlabel metal3 s 335 2084 433 2182 4 gnd
rlabel metal3 s 335 6034 433 6132 4 gnd
rlabel metal3 s 335 45218 433 45316 4 gnd
rlabel metal3 s 335 83454 433 83552 4 gnd
rlabel metal3 s 335 35738 433 35836 4 gnd
rlabel metal3 s 335 43164 433 43262 4 gnd
rlabel metal3 s 335 59991 433 60089 4 gnd
rlabel metal3 s 335 78161 433 78259 4 gnd
rlabel metal3 s 335 42848 433 42946 4 gnd
rlabel metal3 s 335 64178 433 64276 4 gnd
rlabel metal3 s 335 42374 433 42472 4 gnd
rlabel metal3 s 335 46008 433 46106 4 gnd
rlabel metal3 s 335 72868 433 72966 4 gnd
rlabel metal3 s 335 89458 433 89556 4 gnd
rlabel metal3 s 335 1531 433 1629 4 gnd
rlabel metal3 s 335 72078 433 72176 4 gnd
rlabel metal3 s 335 2874 433 2972 4 gnd
rlabel metal3 s 335 52328 433 52426 4 gnd
rlabel metal3 s 335 17331 433 17429 4 gnd
rlabel metal3 s 335 34948 433 35046 4 gnd
rlabel metal3 s 335 86614 433 86712 4 gnd
rlabel metal3 s 335 81084 433 81182 4 gnd
rlabel metal3 s 335 100518 433 100616 4 gnd
rlabel metal3 s 335 741 433 839 4 gnd
rlabel metal3 s 335 29181 433 29279 4 gnd
rlabel metal3 s 335 22308 433 22406 4 gnd
rlabel metal3 s 335 93724 433 93822 4 gnd
rlabel metal3 s 335 20491 433 20589 4 gnd
rlabel metal3 s 335 55251 433 55349 4 gnd
rlabel metal3 s 335 21281 433 21379 4 gnd
rlabel metal3 s 335 77371 433 77469 4 gnd
rlabel metal3 s 335 24678 433 24776 4 gnd
rlabel metal3 s 335 37318 433 37416 4 gnd
rlabel metal3 s 335 7614 433 7712 4 gnd
rlabel metal3 s 335 28391 433 28489 4 gnd
rlabel metal3 s 335 93961 433 94059 4 gnd
rlabel metal3 s 335 63388 433 63486 4 gnd
rlabel metal3 s 335 99728 433 99826 4 gnd
rlabel metal3 s 335 9668 433 9766 4 gnd
rlabel metal3 s 335 55488 433 55586 4 gnd
rlabel metal3 s 335 80768 433 80866 4 gnd
rlabel metal3 s 335 43401 433 43499 4 gnd
rlabel metal3 s 335 95778 433 95876 4 gnd
rlabel metal3 s 335 51301 433 51399 4 gnd
rlabel metal3 s 335 11564 433 11662 4 gnd
rlabel metal3 s 335 8641 433 8739 4 gnd
rlabel metal3 s 335 26258 433 26356 4 gnd
rlabel metal3 s 335 30761 433 30859 4 gnd
rlabel metal3 s 335 77608 433 77706 4 gnd
rlabel metal3 s 335 92144 433 92242 4 gnd
rlabel metal3 s 335 67654 433 67752 4 gnd
rlabel metal3 s 335 85824 433 85922 4 gnd
rlabel metal3 s 335 29418 433 29516 4 gnd
rlabel metal3 s 335 32341 433 32439 4 gnd
rlabel metal3 s 335 43638 433 43736 4 gnd
rlabel metal3 s 335 33684 433 33782 4 gnd
rlabel metal3 s 335 71604 433 71702 4 gnd
rlabel metal3 s 335 41584 433 41682 4 gnd
rlabel metal3 s 335 63941 433 64039 4 gnd
rlabel metal3 s 335 13381 433 13479 4 gnd
rlabel metal3 s 335 44191 433 44289 4 gnd
rlabel metal3 s 335 47588 433 47686 4 gnd
rlabel metal3 s 335 30524 433 30622 4 gnd
rlabel metal3 s 335 11248 433 11346 4 gnd
rlabel metal3 s 335 62598 433 62696 4 gnd
rlabel metal3 s 335 37081 433 37179 4 gnd
rlabel metal3 s 335 27048 433 27146 4 gnd
rlabel metal3 s 335 38108 433 38206 4 gnd
rlabel metal3 s 335 101308 433 101406 4 gnd
rlabel metal3 s 335 36844 433 36942 4 gnd
rlabel metal3 s 335 60228 433 60326 4 gnd
rlabel metal3 s 335 36054 433 36152 4 gnd
rlabel metal3 s 335 54461 433 54559 4 gnd
rlabel metal3 s 335 63151 433 63249 4 gnd
rlabel metal3 s 335 46324 433 46422 4 gnd
rlabel metal3 s 335 76818 433 76916 4 gnd
rlabel metal3 s 335 78398 433 78496 4 gnd
rlabel metal3 s 335 55804 433 55902 4 gnd
rlabel metal3 s 335 67338 433 67436 4 gnd
rlabel metal3 s 335 78714 433 78812 4 gnd
rlabel metal3 s 335 79188 433 79286 4 gnd
rlabel metal3 s 335 23651 433 23749 4 gnd
rlabel metal3 s 335 23098 433 23196 4 gnd
rlabel metal3 s 335 48141 433 48239 4 gnd
rlabel metal3 s 335 9984 433 10082 4 gnd
rlabel metal3 s 335 55014 433 55112 4 gnd
rlabel metal3 s 335 53671 433 53769 4 gnd
rlabel metal3 s 335 48931 433 49029 4 gnd
rlabel metal3 s 335 101624 433 101722 4 gnd
rlabel metal3 s 335 84481 433 84579 4 gnd
rlabel metal3 s 335 36291 433 36389 4 gnd
rlabel metal3 s 335 70261 433 70359 4 gnd
rlabel metal3 s 335 72631 433 72729 4 gnd
rlabel metal3 s 335 53908 433 54006 4 gnd
rlabel metal3 s 335 88668 433 88766 4 gnd
rlabel metal3 s 335 16778 433 16876 4 gnd
rlabel metal3 s 335 58964 433 59062 4 gnd
rlabel metal3 s 335 56594 433 56692 4 gnd
rlabel metal3 s 335 24441 433 24539 4 gnd
rlabel metal3 s 335 84244 433 84342 4 gnd
rlabel metal3 s 335 76581 433 76679 4 gnd
rlabel metal3 s 335 27601 433 27699 4 gnd
rlabel metal3 s 335 33131 433 33229 4 gnd
rlabel metal3 s 335 59201 433 59299 4 gnd
rlabel metal3 s 335 58411 433 58509 4 gnd
rlabel metal3 s 335 91591 433 91689 4 gnd
rlabel metal3 s 335 89774 433 89872 4 gnd
rlabel metal3 s 335 91038 433 91136 4 gnd
rlabel metal3 s 335 4138 433 4236 4 gnd
rlabel metal3 s 335 15198 433 15296 4 gnd
rlabel metal3 s 335 33368 433 33466 4 gnd
rlabel metal3 s 335 44744 433 44842 4 gnd
rlabel metal3 s 335 84718 433 84816 4 gnd
rlabel metal3 s 335 70814 433 70912 4 gnd
rlabel metal3 s 335 23414 433 23512 4 gnd
rlabel metal3 s 335 29971 433 30069 4 gnd
rlabel metal3 s 335 96094 433 96192 4 gnd
rlabel metal3 s 335 32104 433 32202 4 gnd
rlabel metal3 s 335 79741 433 79839 4 gnd
rlabel metal3 s 335 79504 433 79602 4 gnd
rlabel metal3 s 335 17094 433 17192 4 gnd
rlabel metal3 s 335 61018 433 61116 4 gnd
rlabel metal3 s 335 17884 433 17982 4 gnd
rlabel metal3 s 335 79978 433 80076 4 gnd
rlabel metal3 s 335 92618 433 92716 4 gnd
rlabel metal3 s 335 38424 433 38522 4 gnd
rlabel metal3 s 335 58648 433 58746 4 gnd
rlabel metal3 s 335 49721 433 49819 4 gnd
rlabel metal3 s 335 71841 433 71939 4 gnd
rlabel metal3 s 335 99254 433 99352 4 gnd
rlabel metal3 s 335 12828 433 12926 4 gnd
rlabel metal3 s 335 41821 433 41919 4 gnd
rlabel metal3 s 335 82901 433 82999 4 gnd
rlabel metal3 s 335 95304 433 95402 4 gnd
rlabel metal3 s 335 74764 433 74862 4 gnd
rlabel metal3 s 335 22071 433 22169 4 gnd
rlabel metal3 s 335 96331 433 96429 4 gnd
rlabel metal3 s 335 76344 433 76442 4 gnd
rlabel metal3 s 335 29734 433 29832 4 gnd
rlabel metal3 s 335 85034 433 85132 4 gnd
rlabel metal3 s 335 31551 433 31649 4 gnd
rlabel metal3 s 335 70024 433 70122 4 gnd
rlabel metal3 s 335 100044 433 100142 4 gnd
rlabel metal3 s 335 71288 433 71386 4 gnd
rlabel metal3 s 335 4691 433 4789 4 gnd
rlabel metal3 s 335 86298 433 86396 4 gnd
rlabel metal3 s 335 89221 433 89319 4 gnd
rlabel metal3 s 335 96884 433 96982 4 gnd
rlabel metal3 s 335 4928 433 5026 4 gnd
rlabel metal3 s 335 94514 433 94612 4 gnd
rlabel metal3 s 335 15751 433 15849 4 gnd
rlabel metal3 s 335 52644 433 52742 4 gnd
rlabel metal3 s 335 77134 433 77232 4 gnd
rlabel metal3 s 335 94751 433 94849 4 gnd
rlabel metal3 s 335 21518 433 21616 4 gnd
rlabel metal3 s 335 69471 433 69569 4 gnd
rlabel metal3 s 335 51064 433 51162 4 gnd
rlabel metal3 s 335 40478 433 40576 4 gnd
rlabel metal3 s 335 85271 433 85369 4 gnd
rlabel metal3 s 335 2558 433 2656 4 gnd
rlabel metal3 s 335 56831 433 56929 4 gnd
rlabel metal3 s 335 62361 433 62459 4 gnd
rlabel metal3 s 335 12591 433 12689 4 gnd
rlabel metal3 s 335 42611 433 42709 4 gnd
rlabel metal3 s 335 43954 433 44052 4 gnd
rlabel metal3 s 335 98938 433 99036 4 gnd
rlabel metal3 s 335 69708 433 69806 4 gnd
rlabel metal3 s 335 10458 433 10556 4 gnd
rlabel metal3 s 335 97911 433 98009 4 gnd
rlabel metal3 s 335 19464 433 19562 4 gnd
rlabel metal3 s 335 90248 433 90346 4 gnd
rlabel metal3 s 335 39451 433 39549 4 gnd
rlabel metal3 s 335 73658 433 73756 4 gnd
rlabel metal3 s 335 100834 433 100932 4 gnd
rlabel metal3 s 335 91354 433 91452 4 gnd
rlabel metal3 s 335 78951 433 79049 4 gnd
rlabel metal3 s 335 54698 433 54796 4 gnd
rlabel metal3 s 335 82111 433 82209 4 gnd
rlabel metal3 s 335 20728 433 20826 4 gnd
rlabel metal3 s 335 71051 433 71149 4 gnd
rlabel metal3 s 335 44428 433 44526 4 gnd
rlabel metal3 s 335 36528 433 36626 4 gnd
rlabel metal3 s 335 73184 433 73282 4 gnd
rlabel metal3 s 335 57068 433 57166 4 gnd
rlabel metal3 s 335 74211 433 74309 4 gnd
rlabel metal3 s 335 39214 433 39312 4 gnd
rlabel metal3 s 335 90011 433 90109 4 gnd
rlabel metal3 s 335 4454 433 4552 4 gnd
rlabel metal3 s 335 8404 433 8502 4 gnd
rlabel metal3 s 335 30998 433 31096 4 gnd
rlabel metal3 s 335 75554 433 75652 4 gnd
rlabel metal3 s 335 91828 433 91926 4 gnd
rlabel metal3 s 335 73974 433 74072 4 gnd
rlabel metal3 s 335 35501 433 35599 4 gnd
rlabel metal3 s 335 93408 433 93506 4 gnd
rlabel metal3 s 335 30208 433 30306 4 gnd
rlabel metal3 s 335 87088 433 87186 4 gnd
rlabel metal3 s 335 26574 433 26672 4 gnd
rlabel metal3 s 335 101071 433 101169 4 gnd
rlabel metal3 s 335 62124 433 62222 4 gnd
rlabel metal3 s 335 51538 433 51636 4 gnd
rlabel metal3 s 335 11801 433 11899 4 gnd
rlabel metal3 s 335 90564 433 90662 4 gnd
rlabel metal3 s 335 8088 433 8186 4 gnd
rlabel metal3 s 335 61571 433 61669 4 gnd
rlabel metal3 s 335 15514 433 15612 4 gnd
<< properties >>
string FIXED_BBOX 0 0 624 102305
<< end >>
