* NGSPICE file created from low_freq_pll_flat.ext - technology: sky130A

.subckt low_freq_pll_flat VDD VSS vsigin ibiasn vcp
X0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_34309_6805# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=4.23972e+13p ps=4.1226e+08u w=650000u l=150000u
X1 VSS a_31186_5717# a_31144_6121# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+11p ps=1.53e+06u w=420000u l=150000u
X2 cs_ring_osc_0/cs_ring_osc_stage_3/vin cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_17431_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X3 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N a_29107_13961# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=1.60678e+14p ps=1.23322e+09u w=1e+06u l=150000u
X4 a_26616_1344# cs_ring_osc_0/vpbias a_27074_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X5 a_11056_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/vin a_10598_n20414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X6 a_26208_9468# cs_ring_osc_0/cs_ring_osc_stage_5/vout a_25750_9468# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X7 cs_ring_osc_0/cs_ring_osc_stage_0/voutcs cs_ring_osc_0/vosc a_12430_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X8 a_20446_n5874# vcp a_19988_n5874# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X9 VDD freq_div_0/sky130_fd_sc_hd__inv_4_10/A freq_div_0/sky130_fd_sc_hd__inv_4_10/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X10 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X11 VSS VSS cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X12 cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X13 pfd_cp_lpf_0/vRSTN pfd_cp_lpf_0/vQA a_29765_13961# VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X14 a_33716_7741# a_33443_7375# a_33631_7375# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X15 a_13614_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/voutcs cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X16 freq_div_0/sky130_fd_sc_hd__inv_4_0/A freq_div_0/sky130_fd_sc_hd__inv_1_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X17 VSS a_31611_7643# a_31569_7375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X18 a_25599_n921# cs_ring_osc_0/cs_ring_osc_stage_5/vin a_25141_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X19 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q a_31611_7893# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20 a_14698_6217# cs_ring_osc_0/vpbias a_15156_6217# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X21 a_9683_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/vin cs_ring_osc_0/cs_ring_osc_stage_2/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=4.06e+12p ps=2.916e+07u w=6e+06u l=2e+06u
X22 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q a_33277_6287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X23 a_11972_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/vin a_11514_n20414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X24 VSS VSS cs_ring_osc_0/cs_ring_osc_stage_4/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=2e+06u
X25 a_16056_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_15598_n20414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X26 VSS freq_div_0/sky130_fd_sc_hd__inv_4_3/A freq_div_0/sky130_fd_sc_hd__inv_4_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X27 cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X28 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X29 a_26056_n21082# vcp a_25598_n21082# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X30 cs_ring_osc_0/cs_ring_osc_stage_5/vin VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=2e+06u
X31 VSS freq_div_0/vout a_27287_13961# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X32 cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X33 a_28613_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs cs_ring_osc_0/cs_ring_osc_stage_5/vin VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=2e+06u
X34 a_31079_14103# vsigin VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X35 freq_div_0/sky130_fd_sc_hd__inv_4_10/A freq_div_0/sky130_fd_sc_hd__inv_1_10/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X36 VDD a_34309_5717# a_34225_5743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.764e+11p ps=1.68e+06u w=420000u l=150000u
X37 VSS freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_30579_5749# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X38 a_29682_n2414# cs_ring_osc_0/cs_ring_osc_stage_5/voutcs VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X39 a_21362_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/vin a_20904_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X40 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X41 VSS VDD a_31798_14327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X42 a_31018_8829# a_30745_8463# a_30933_8463# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X43 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q a_31611_6805# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X44 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X45 a_33716_7919# a_33443_7925# a_33631_7919# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X46 cs_ring_osc_0/cs_ring_osc_stage_1/csinvn cs_ring_osc_0/cs_ring_osc_stage_1/vin a_21362_n6542# VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=2e+06u
X47 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X48 cs_ring_osc_0/cs_ring_osc_stage_4/csinvp cs_ring_osc_0/vpbias a_32138_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.06e+12p pd=2.916e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X49 VDD VDD pfd_cp_lpf_0/vpbias VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.29e+07u w=1e+06u l=4e+06u
X50 VDD a_30294_13935# pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X51 a_31166_14327# a_31040_14229# a_30762_14213# VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X52 a_15599_n921# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_15141_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X53 a_16972_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_16514_n20414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X54 a_31443_8829# a_30745_8463# a_31186_8575# VSS sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=1.978e+11p ps=1.99e+06u w=360000u l=150000u
X55 VSS a_31611_7893# a_32042_7919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X56 VDD a_33884_7487# a_33811_7741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X57 a_27074_1344# cs_ring_osc_0/vpbias a_26616_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X58 a_26972_n21082# vcp a_26514_n21082# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X59 VDD freq_div_0/sky130_fd_sc_hd__inv_4_5/A freq_div_0/sky130_fd_sc_hd__inv_4_5/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X60 a_25242_1344# cs_ring_osc_0/vpbias a_25700_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X61 a_27990_n16656# cs_ring_osc_0/vpbias cs_ring_osc_0/cs_ring_osc_stage_3/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=4.06e+12p ps=2.916e+07u w=8e+06u l=2e+06u
X62 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X63 a_36361_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/vin a_35903_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X64 VDD a_28543_13935# a_28530_14327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X65 a_31018_7741# a_30745_7375# a_30933_7375# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X66 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X67 a_33716_6831# a_33443_6837# a_33631_6831# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X68 pfd_cp_lpf_0/vpbias ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=4e+06u
X69 a_33811_7741# a_33277_7375# a_33716_7741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X70 freq_div_0/sky130_fd_sc_hd__inv_1_5/A a_32042_5743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X71 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X72 a_16988_6217# cs_ring_osc_0/vpbias a_16530_6217# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X73 freq_div_0/sky130_fd_sc_hd__inv_4_0/Y freq_div_0/sky130_fd_sc_hd__inv_4_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X74 a_15140_n2414# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_14682_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X75 VSS ibiasn ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.74e+12p ps=1.548e+07u w=1e+06u l=4e+06u
X76 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X77 a_11158_1344# cs_ring_osc_0/vpbias a_11616_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X78 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X79 a_33884_7893# a_33716_7919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.978e+11p pd=1.99e+06u as=0p ps=0u w=640000u l=150000u
X80 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X81 a_29529_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_29071_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X82 VDD a_33884_7893# a_33811_7919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X83 a_34141_7919# a_33443_7925# a_33884_7893# VSS sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=0p ps=0u w=360000u l=150000u
X84 VSS VSS cs_ring_osc_0/cs_ring_osc_stage_1/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X85 cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X86 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X87 a_27074_n16656# cs_ring_osc_0/vpbias a_27532_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X88 a_20445_n9035# cs_ring_osc_0/cs_ring_osc_stage_1/vin a_19987_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X89 VDD a_31611_6555# a_32042_6609# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X90 a_31018_7919# a_30745_7925# a_30933_7919# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X91 a_34072_n5874# vcp a_33614_n5874# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X92 a_26972_n2414# cs_ring_osc_0/cs_ring_osc_stage_5/vin a_26514_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X93 a_33811_7919# a_33277_7925# a_33716_7919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X94 VSS freq_div_0/sky130_fd_sc_hd__inv_4_7/A freq_div_0/sky130_fd_sc_hd__inv_4_7/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X95 freq_div_0/sky130_fd_sc_hd__inv_1_10/A a_34740_5743# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X96 a_34530_n5874# vcp a_34072_n5874# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X97 VSS vcp a_12430_n21082# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X98 a_30762_14213# a_31079_14103# a_31037_13961# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=360000u l=150000u
X99 a_27430_n2414# cs_ring_osc_0/cs_ring_osc_stage_5/vin a_26972_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X100 VSS a_31611_7643# a_32042_7697# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X101 VDD a_33884_6805# a_33811_6831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X102 a_27125_7037# cs_ring_osc_0/cs_ring_osc_stage_5/vout a_26667_7037# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X103 VDD VDD cs_ring_osc_0/cs_ring_osc_stage_4/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X104 a_31018_6831# a_30745_6837# a_30933_6831# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X105 a_31222_n11700# cs_ring_osc_0/vpbias a_30764_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X106 a_27708_13961# VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X107 VDD a_31079_14103# a_31040_14229# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X108 a_10598_n2414# cs_ring_osc_0/vosc a_10140_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X109 a_14848_n11700# cs_ring_osc_0/vpbias a_14390_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X110 a_33811_6831# a_33277_6837# a_33716_6831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X111 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X112 VSS VSS cs_ring_osc_0/cs_ring_osc_stage_3/voutcs VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X113 a_26973_n921# cs_ring_osc_0/cs_ring_osc_stage_5/vin a_26515_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X114 a_16056_n2414# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_15598_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X115 a_16514_n2414# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_16056_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X116 VDD cs_ring_osc_0/vpbias a_25242_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X117 VDD pfd_cp_lpf_0/vpbias pfd_cp_lpf_0/vswitchh VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.61e+12p ps=2.206e+07u w=1e+06u l=4e+06u
X118 a_26666_9468# cs_ring_osc_0/cs_ring_osc_stage_5/vout a_26208_9468# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X119 a_31186_7893# a_31018_7919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.978e+11p pd=1.99e+06u as=0p ps=0u w=640000u l=150000u
X120 a_11158_n16656# cs_ring_osc_0/vpbias a_11616_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X121 VDD a_31443_8829# a_31611_8731# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X122 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X123 a_28021_14203# a_27803_13961# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X124 a_31443_7919# a_30745_7925# a_31186_7893# VSS sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=0p ps=0u w=360000u l=150000u
X125 a_34225_7741# a_33443_7375# a_34141_7741# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X126 a_12990_1344# cs_ring_osc_0/vpbias a_12532_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X127 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X128 VDD pfd_cp_lpf_0/vpbias pfd_cp_lpf_0/vswitchh VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X129 a_34988_n5874# vcp a_34530_n5874# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X130 cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X131 a_15764_n11700# cs_ring_osc_0/vpbias a_15306_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X132 a_31018_8829# a_30579_8463# a_30933_8463# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=1.626e+11p ps=1.66e+06u w=360000u l=150000u
X133 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs cs_ring_osc_0/cs_ring_osc_stage_5/vin a_27430_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X134 a_35446_n5874# vcp a_34988_n5874# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X135 cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X136 VSS freq_div_0/sky130_fd_sc_hd__inv_4_3/A freq_div_0/sky130_fd_sc_hd__inv_4_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X137 cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X138 a_9682_n21082# vcp cs_ring_osc_0/cs_ring_osc_stage_2/csinvn VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=5.8e+11p ps=5.16e+06u w=1e+06u l=2e+06u
X139 a_26515_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/vin a_26057_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X140 a_28614_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X141 a_17446_9468# vcp a_16988_9468# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X142 a_10242_n16656# cs_ring_osc_0/vpbias a_10700_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X143 VSS ibiasn ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X144 freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_34309_7643# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X145 a_16973_n921# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_16515_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X146 a_31144_8463# a_30745_8463# a_31018_8829# VSS sky130_fd_pr__nfet_01v8 ad=1.392e+11p pd=1.53e+06u as=0p ps=0u w=360000u l=150000u
X147 VSS a_31443_8829# a_31611_8731# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X148 freq_div_0/sky130_fd_sc_hd__inv_1_3/A a_32042_7697# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X149 a_31527_8829# a_30745_8463# a_31443_8829# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X150 a_34225_7919# a_33443_7925# a_34141_7919# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X151 a_16680_n11700# cs_ring_osc_0/vpbias a_16222_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X152 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X153 a_34071_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/vin a_33613_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X154 VSS VSS cs_ring_osc_0/cs_ring_osc_stage_0/voutcs VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X155 a_20904_n5874# vcp a_20446_n5874# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X156 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X157 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X158 a_27431_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/vin a_26973_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X159 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X160 a_36362_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/vin a_35904_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X161 a_16530_6217# cs_ring_osc_0/vpbias a_16988_6217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X162 VSS a_31186_8575# a_31144_8463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X163 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_33277_7925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X164 a_31527_7741# a_30745_7375# a_31443_7741# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X165 freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_34309_7643# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X166 VDD a_31186_6399# a_31113_6653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X167 VDD cs_ring_osc_0/vpbias a_10242_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X168 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X169 cs_ring_osc_0/cs_ring_osc_stage_4/csinvn cs_ring_osc_0/cs_ring_osc_stage_4/vin a_36362_n6542# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X170 a_34225_6831# a_33443_6837# a_34141_6831# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X171 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y freq_div_0/sky130_fd_sc_hd__inv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X172 cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X173 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X174 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q a_30579_6837# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X175 a_33443_7375# a_33277_7375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X176 a_33443_7925# a_33277_7925# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X177 a_31113_6653# a_30579_6287# a_31018_6653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X178 freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q a_31611_7643# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X179 VSS a_34309_5717# a_34267_6121# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X180 a_20446_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/vin a_19988_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X181 a_24682_n2414# cs_ring_osc_0/cs_ring_osc_stage_5/vin cs_ring_osc_0/cs_ring_osc_stage_5/csinvn VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=5.8e+11p ps=5.16e+06u w=1e+06u l=2e+06u
X182 cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X183 a_31527_7919# a_30745_7925# a_31443_7919# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X184 a_25242_1344# cs_ring_osc_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X185 a_30140_n2414# cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_29682_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X186 a_33443_5749# a_33277_5749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X187 a_34987_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/vin a_34529_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X188 VSS a_33884_6805# a_33842_7209# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+11p ps=1.53e+06u w=420000u l=150000u
X189 a_30745_8463# a_30579_8463# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X190 a_31018_7919# a_30579_7925# a_30933_7919# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=1.626e+11p ps=1.66e+06u w=360000u l=150000u
X191 VDD a_34309_5717# a_34740_5743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X192 a_35445_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/vin a_34987_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=2e+06u
X193 VSS VSS cs_ring_osc_0/cs_ring_osc_stage_4/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X194 VSS freq_div_0/vin a_30579_8463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X195 freq_div_0/sky130_fd_sc_hd__inv_4_9/A freq_div_0/sky130_fd_sc_hd__inv_1_9/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X196 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X197 a_31361_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_30903_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X198 a_15156_6217# cs_ring_osc_0/vpbias a_14698_6217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X199 a_27583_7037# cs_ring_osc_0/cs_ring_osc_stage_5/vout a_27125_7037# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=2e+06u
X200 freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q a_31611_7643# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X201 a_33716_6653# a_33277_6287# a_33631_6287# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=1.626e+11p ps=1.66e+06u w=360000u l=150000u
X202 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X203 VSS ibiasn ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X204 cs_ring_osc_0/vosc cs_ring_osc_0/cs_ring_osc_stage_5/vout a_27582_9468# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X205 a_31527_6831# a_30745_6837# a_31443_6831# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X206 VDD a_31186_5717# a_31113_5743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X207 a_12990_1344# cs_ring_osc_0/vpbias cs_ring_osc_0/cs_ring_osc_stage_0/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.06e+12p ps=2.916e+07u w=8e+06u l=2e+06u
X208 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X209 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y freq_div_0/sky130_fd_sc_hd__inv_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X210 cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X211 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X212 cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X213 a_31144_8297# a_30745_7925# a_31018_7919# VSS sky130_fd_pr__nfet_01v8 ad=1.392e+11p pd=1.53e+06u as=0p ps=0u w=360000u l=150000u
X214 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X215 a_30745_7375# a_30579_7375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X216 pfd_cp_lpf_0/vndiode pfd_cp_lpf_0/vndiode VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X217 a_30745_7925# a_30579_7925# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X218 a_31113_5743# a_30579_5749# a_31018_5743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X219 a_11514_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/vin a_11056_n20414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X220 a_33443_7375# a_33277_7375# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X221 a_33842_6287# a_33443_6287# a_33716_6653# VSS sky130_fd_pr__nfet_01v8 ad=1.392e+11p pd=1.53e+06u as=0p ps=0u w=360000u l=150000u
X222 VSS a_31611_5717# a_31569_6121# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X223 a_25598_n2414# cs_ring_osc_0/cs_ring_osc_stage_5/vin a_25140_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X224 a_18820_9468# vcp a_18362_9468# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X225 a_20903_n9035# cs_ring_osc_0/cs_ring_osc_stage_1/vin a_20445_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=2e+06u
X226 a_33631_6831# freq_div_0/sky130_fd_sc_hd__inv_4_8/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.626e+11p pd=1.66e+06u as=0p ps=0u w=420000u l=150000u
X227 VDD freq_div_0/sky130_fd_sc_hd__inv_4_9/A freq_div_0/sky130_fd_sc_hd__inv_4_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X228 a_30745_5749# a_30579_5749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X229 pfd_cp_lpf_0/vswitchh VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X230 VSS a_33884_6399# a_33842_6287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X231 a_25700_n16656# cs_ring_osc_0/vpbias a_26158_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X232 a_28530_14327# a_27453_13961# a_28368_13961# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X233 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X234 a_12430_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/vin a_11972_n20414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X235 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X236 VSS ibiasn ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X237 a_16514_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_16056_n20414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X238 VDD pfd_cp_lpf_0/vQA pfd_cp_lpf_0/vQAb VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X239 cs_ring_osc_0/cs_ring_osc_stage_5/csinvp cs_ring_osc_0/vpbias a_27990_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.06e+12p pd=2.916e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X240 a_25141_n921# cs_ring_osc_0/cs_ring_osc_stage_5/vin a_24683_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X241 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X242 a_26514_n21082# vcp a_26056_n21082# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X243 cs_ring_osc_0/cs_ring_osc_stage_0/csinvn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=2e+06u
X244 a_24834_9468# cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X245 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X246 cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X247 freq_div_0/sky130_fd_sc_hd__inv_1_9/A a_34740_6609# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X248 a_11056_n2414# cs_ring_osc_0/vosc a_10598_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X249 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X250 a_34072_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/vin a_33614_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X251 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X252 a_11514_n2414# cs_ring_osc_0/vosc a_11056_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X253 a_34530_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/vin a_34072_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X254 VDD freq_div_0/sky130_fd_sc_hd__inv_4_6/A freq_div_0/sky130_fd_sc_hd__inv_4_6/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X255 freq_div_0/sky130_fd_sc_hd__inv_4_3/A freq_div_0/sky130_fd_sc_hd__inv_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X256 a_25599_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/vin a_25141_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X257 a_29848_n11700# cs_ring_osc_0/vpbias a_30306_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X258 a_30745_7375# a_30579_7375# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X259 a_17430_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_16972_n20414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X260 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y freq_div_0/sky130_fd_sc_hd__inv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X261 a_27430_n21082# vcp a_26972_n21082# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X262 cs_ring_osc_0/cs_ring_osc_stage_1/csinvp cs_ring_osc_0/cs_ring_osc_stage_1/vin a_21361_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.06e+12p pd=2.916e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X263 cs_ring_osc_0/vpbias VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X264 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X265 a_25700_1344# cs_ring_osc_0/vpbias a_26158_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X266 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X267 cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X268 a_30933_6831# freq_div_0/sky130_fd_sc_hd__inv_4_2/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.626e+11p pd=1.66e+06u as=0p ps=0u w=420000u l=150000u
X269 VDD freq_div_0/sky130_fd_sc_hd__inv_4_4/A freq_div_0/sky130_fd_sc_hd__inv_4_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X270 a_33631_6287# freq_div_0/sky130_fd_sc_hd__inv_4_9/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X271 a_15141_n921# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_14683_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X272 VSS VSS cs_ring_osc_0/cs_ring_osc_stage_5/voutcs VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X273 a_35904_n5874# vcp a_35446_n5874# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X274 VDD a_34309_7643# a_34740_7697# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X275 VDD freq_div_0/sky130_fd_sc_hd__inv_4_8/A freq_div_0/sky130_fd_sc_hd__inv_4_8/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X276 VDD cs_ring_osc_0/vpbias a_29390_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X277 a_28543_13935# a_28368_13961# a_28722_13961# VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X278 a_33884_7487# a_33716_7741# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X279 a_33884_7487# a_33716_7741# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.978e+11p pd=1.99e+06u as=0p ps=0u w=640000u l=150000u
X280 a_15306_n11700# cs_ring_osc_0/vpbias a_15764_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X281 a_33884_5717# a_33716_5743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X282 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X283 a_34141_6653# a_33277_6287# a_33884_6399# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=2.19e+11p ps=2.15e+06u w=420000u l=150000u
X284 a_9682_n3082# vcp cs_ring_osc_0/cs_ring_osc_stage_0/csinvn VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X285 a_34988_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/vin a_34530_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X286 cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X287 a_35446_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/vin a_34988_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X288 VSS cs_ring_osc_0/vosc2 freq_div_0/vin VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X289 VDD cs_ring_osc_0/vpbias a_14240_6217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X290 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X291 VDD VDD pfd_cp_lpf_0/vswitchh VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X292 VSS a_30391_13935# pfd_cp_lpf_0/vQA VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X293 VDD freq_div_0/sky130_fd_sc_hd__inv_4_1/A freq_div_0/sky130_fd_sc_hd__inv_4_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X294 VSS a_31611_5717# a_32042_5743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X295 a_31362_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_30904_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X296 cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X297 a_24682_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/vin cs_ring_osc_0/cs_ring_osc_stage_3/csinvn VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=5.8e+11p ps=5.16e+06u w=1e+06u l=2e+06u
X298 VSS cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_31362_n6542# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X299 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y freq_div_0/sky130_fd_sc_hd__inv_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X300 cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X301 a_29683_n921# cs_ring_osc_0/cs_ring_osc_stage_5/voutcs VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=2e+06u
X302 VSS a_31235_14198# a_31166_14327# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X303 a_30933_6287# freq_div_0/sky130_fd_sc_hd__inv_4_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.626e+11p pd=1.66e+06u as=0p ps=0u w=420000u l=150000u
X304 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X305 cs_ring_osc_0/cs_ring_osc_stage_4/vin cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_32431_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X306 VDD freq_div_0/sky130_fd_sc_hd__inv_4_2/A freq_div_0/sky130_fd_sc_hd__inv_4_2/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X307 VDD a_34141_5743# a_34309_5717# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X308 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X309 cs_ring_osc_0/cs_ring_osc_stage_3/csinvp VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X310 a_12532_n16656# cs_ring_osc_0/vpbias a_12990_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X311 freq_div_0/sky130_fd_sc_hd__inv_4_10/Y freq_div_0/sky130_fd_sc_hd__inv_4_10/A VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X312 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X313 cs_ring_osc_0/vosc2 cs_ring_osc_0/vosc VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X314 a_31186_7487# a_31018_7741# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X315 a_31186_7487# a_31018_7741# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.978e+11p pd=1.99e+06u as=0p ps=0u w=640000u l=150000u
X316 VDD freq_div_0/sky130_fd_sc_hd__inv_4_9/A freq_div_0/sky130_fd_sc_hd__inv_4_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X317 a_20904_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/vin a_20446_n6542# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X318 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X319 a_29682_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/voutcs VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X320 a_14390_n11700# cs_ring_osc_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X321 a_33716_6831# a_33277_6837# a_33631_6831# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=0p ps=0u w=360000u l=150000u
X322 a_31186_5717# a_31018_5743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X323 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X324 a_25140_n2414# cs_ring_osc_0/cs_ring_osc_stage_5/vin a_24682_n2414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X325 a_31569_8463# a_30579_8463# a_31443_8829# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X326 a_31443_6653# a_30579_6287# a_31186_6399# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=2.19e+11p ps=2.15e+06u w=420000u l=150000u
X327 a_34141_5743# a_33277_5749# a_33884_5717# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X328 a_27074_1344# cs_ring_osc_0/vpbias a_27532_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X329 VSS freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_33277_6837# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X330 a_25141_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/vin a_24683_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X331 a_11616_n16656# cs_ring_osc_0/vpbias a_12074_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X332 a_25751_7037# cs_ring_osc_0/cs_ring_osc_stage_5/vout a_25293_7037# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X333 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X334 a_10242_n16656# cs_ring_osc_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X335 a_30445_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_29987_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X336 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X337 a_31056_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_30598_n20414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X338 a_10598_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/vin a_10140_n20414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X339 a_28477_13961# a_27287_13961# a_28368_13961# VSS sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X340 a_35903_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/vin a_35445_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X341 a_31235_14198# a_31040_14229# a_31545_13961# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=2.802e+11p ps=2.2e+06u w=360000u l=150000u
X342 a_33842_7209# a_33443_6837# a_33716_6831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X343 a_16988_9468# vcp a_16530_9468# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X344 a_33716_5743# a_33277_5749# a_33631_5743# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=1.626e+11p ps=1.66e+06u w=360000u l=150000u
X345 a_15156_6217# cs_ring_osc_0/vpbias a_15614_6217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X346 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X347 cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X348 cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X349 VDD freq_div_0/sky130_fd_sc_hd__inv_4_6/A freq_div_0/sky130_fd_sc_hd__inv_4_6/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X350 VDD a_34309_7643# a_34225_7741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X351 VDD a_31443_5743# a_31611_5717# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X352 cs_ring_osc_0/cs_ring_osc_stage_0/csinvp VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X353 a_30141_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_29683_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X354 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y freq_div_0/sky130_fd_sc_hd__inv_4_5/A VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X355 a_31972_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_31514_n20414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X356 pfd_cp_lpf_0/vswitchl pfd_cp_lpf_0/vQB vcp VSS sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X357 a_34267_8297# a_33277_7925# a_34141_7919# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X358 a_33842_6121# a_33443_5749# a_33716_5743# VSS sky130_fd_pr__nfet_01v8 ad=1.392e+11p pd=1.53e+06u as=0p ps=0u w=360000u l=150000u
X359 a_15598_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_15140_n20414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X360 VDD a_31611_6555# a_31527_6653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.764e+11p ps=1.68e+06u w=420000u l=150000u
X361 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X362 a_25598_n21082# vcp a_25140_n21082# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X363 VDD pfd_cp_lpf_0/vpbias pfd_cp_lpf_0/vpbias VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X364 VDD freq_div_0/sky130_fd_sc_hd__inv_4_4/A freq_div_0/sky130_fd_sc_hd__inv_4_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X365 a_26056_n2414# cs_ring_osc_0/cs_ring_osc_stage_5/vin a_25598_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X366 a_33614_n5874# vcp VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X367 a_10700_n16656# cs_ring_osc_0/vpbias a_10242_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X368 VDD freq_div_0/sky130_fd_sc_hd__inv_4_8/A freq_div_0/sky130_fd_sc_hd__inv_4_8/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X369 a_26514_n2414# cs_ring_osc_0/cs_ring_osc_stage_5/vin a_26056_n2414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X370 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X371 a_11057_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/vin a_10599_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X372 a_31443_5743# a_30579_5749# a_31186_5717# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X373 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X374 freq_div_0/sky130_fd_sc_hd__inv_1_4/A a_32042_6609# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X375 a_26616_1344# cs_ring_osc_0/vpbias a_26158_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X376 VSS a_31611_8731# a_31569_8463# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X377 freq_div_0/sky130_fd_sc_hd__inv_4_6/A freq_div_0/sky130_fd_sc_hd__inv_1_6/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X378 VDD a_34309_7893# a_34225_7919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X379 VSS freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q a_33277_6287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X380 cs_ring_osc_0/cs_ring_osc_stage_4/csinvp cs_ring_osc_0/cs_ring_osc_stage_4/vin a_36361_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X381 freq_div_0/vin cs_ring_osc_0/vosc2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X382 a_28368_13961# a_27453_13961# a_28021_14203# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X383 a_31235_14198# a_31079_14103# a_31380_14327# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=3.402e+11p ps=3.3e+06u w=420000u l=150000u
X384 VSS freq_div_0/sky130_fd_sc_hd__inv_4_0/A freq_div_0/sky130_fd_sc_hd__inv_4_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X385 cs_ring_osc_0/cs_ring_osc_stage_3/csinvp cs_ring_osc_0/vpbias a_27990_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X386 a_11973_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/vin a_11515_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X387 a_28543_13935# pfd_cp_lpf_0/vRSTN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X388 VDD pfd_cp_lpf_0/vRSTN a_31380_14327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X389 cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X390 a_16057_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_15599_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X391 VDD freq_div_0/sky130_fd_sc_hd__inv_4_1/A freq_div_0/sky130_fd_sc_hd__inv_4_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X392 freq_div_0/sky130_fd_sc_hd__inv_4_8/A freq_div_0/sky130_fd_sc_hd__inv_1_8/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X393 VDD a_34309_6805# a_34225_6831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X394 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q a_30579_6287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X395 cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X396 a_31079_14103# vsigin VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X397 a_31569_8297# a_30579_7925# a_31443_7919# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X398 freq_div_0/sky130_fd_sc_hd__inv_1_1/A a_32042_7919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X399 VDD a_31611_5717# a_31527_5743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.764e+11p ps=1.68e+06u w=420000u l=150000u
X400 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X401 freq_div_0/sky130_fd_sc_hd__inv_4_5/A freq_div_0/sky130_fd_sc_hd__inv_1_5/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X402 a_30294_13935# a_30391_13935# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X403 VDD freq_div_0/sky130_fd_sc_hd__inv_4_2/A freq_div_0/sky130_fd_sc_hd__inv_4_2/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X404 freq_div_0/sky130_fd_sc_hd__inv_4_10/Y freq_div_0/sky130_fd_sc_hd__inv_4_10/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X405 a_16973_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_16515_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X406 vcp VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X407 VDD VDD cs_ring_osc_0/cs_ring_osc_stage_5/vout VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X408 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X409 pfd_cp_lpf_0/VQBb pfd_cp_lpf_0/vQB VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X410 a_33443_5749# a_33277_5749# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X411 cs_ring_osc_0/cs_ring_osc_stage_3/csinvn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X412 freq_div_0/sky130_fd_sc_hd__inv_1_2/A a_32042_6831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X413 a_26158_n16656# cs_ring_osc_0/vpbias a_26616_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X414 pfd_cp_lpf_0/vRSTN pfd_cp_lpf_0/vQB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X415 freq_div_0/sky130_fd_sc_hd__inv_1_6/A a_34740_7919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X416 a_26515_n921# cs_ring_osc_0/cs_ring_osc_stage_5/vin a_26057_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X417 cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X418 a_30764_n11700# cs_ring_osc_0/vpbias a_30306_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X419 cs_ring_osc_0/cs_ring_osc_stage_4/voutcs VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=2e+06u
X420 a_18362_9468# vcp a_17904_9468# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X421 a_10140_n3082# vcp a_9682_n3082# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X422 cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X423 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X424 a_33613_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/vin cs_ring_osc_0/cs_ring_osc_stage_4/voutcs VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X425 a_30446_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_29988_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X426 a_15140_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_14682_n20414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X427 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X428 a_25140_n21082# vcp a_24682_n21082# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X429 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs cs_ring_osc_0/cs_ring_osc_stage_3/vin a_27430_n20414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X430 a_35904_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/vin a_35446_n6542# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X431 a_11972_n3082# vcp a_11514_n3082# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X432 a_25242_n16656# cs_ring_osc_0/vpbias a_25700_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X433 VSS VSS pfd_cp_lpf_0/vpbias VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X434 a_12532_1344# cs_ring_osc_0/vpbias a_12074_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X435 a_32431_n921# cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_31973_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X436 a_12430_n3082# vcp a_11972_n3082# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X437 freq_div_0/sky130_fd_sc_hd__inv_1_8/A a_34740_6831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X438 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X439 a_31680_n11700# cs_ring_osc_0/vpbias a_31222_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=0p ps=0u w=8e+06u l=2e+06u
X440 VSS a_31611_8731# a_32042_8785# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X441 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y freq_div_0/sky130_fd_sc_hd__inv_4_5/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X442 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X443 a_30745_5749# a_30579_5749# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X444 a_9683_n921# cs_ring_osc_0/vosc cs_ring_osc_0/cs_ring_osc_stage_0/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=2e+06u
X445 a_16515_n921# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_16057_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X446 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X447 VDD pfd_cp_lpf_0/vpbias pfd_cp_lpf_0/vpbias VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X448 VSS a_31079_14103# a_31040_14229# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X449 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X450 a_28722_13961# pfd_cp_lpf_0/vRSTN VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X451 a_31380_14327# a_31166_14327# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X452 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X453 a_29390_n11700# cs_ring_osc_0/vpbias a_29848_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X454 VDD VDD cs_ring_osc_0/cs_ring_osc_stage_3/voutcs VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X455 a_15764_n11700# cs_ring_osc_0/vpbias a_16222_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X456 a_34529_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/vin a_34071_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X457 a_30294_13935# a_30391_13935# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X458 VSS a_28543_13935# a_28477_13961# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X459 VDD VDD cs_ring_osc_0/cs_ring_osc_stage_0/voutcs VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X460 freq_div_0/sky130_fd_sc_hd__inv_4_9/Y freq_div_0/sky130_fd_sc_hd__inv_4_9/A VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X461 a_11056_n21082# vcp a_10598_n21082# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X462 VSS vcp a_12430_n3082# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X463 cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X464 cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X465 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X466 a_16988_6217# cs_ring_osc_0/vpbias cs_ring_osc_0/vpbias VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.32e+12p ps=1.658e+07u w=8e+06u l=2e+06u
X467 freq_div_0/sky130_fd_sc_hd__inv_4_10/A freq_div_0/sky130_fd_sc_hd__inv_1_10/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X468 a_30903_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_30445_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X469 VSS a_34141_5743# a_34309_5717# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X470 a_31972_n2414# cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_31514_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X471 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X472 a_31166_14327# a_31079_14103# a_30762_14213# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X473 VSS freq_div_0/sky130_fd_sc_hd__inv_4_0/A freq_div_0/sky130_fd_sc_hd__inv_4_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X474 VSS a_34309_6805# a_34740_6831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X475 a_32430_n2414# cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_31972_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X476 freq_div_0/sky130_fd_sc_hd__inv_1_0/A a_32042_8785# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X477 a_11972_n21082# vcp a_11514_n21082# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X478 pfd_cp_lpf_0/vndiode pfd_cp_lpf_0/vQA pfd_cp_lpf_0/vswitchh VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=1e+06u
X479 VDD a_31186_8575# a_31113_8829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X480 a_12431_n921# cs_ring_osc_0/vosc a_11973_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X481 pfd_cp_lpf_0/vpbias pfd_cp_lpf_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X482 a_12990_n16656# cs_ring_osc_0/vpbias cs_ring_osc_0/cs_ring_osc_stage_2/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X483 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X484 a_33631_6287# freq_div_0/sky130_fd_sc_hd__inv_4_9/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X485 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs cs_ring_osc_0/cs_ring_osc_stage_5/vin a_27431_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X486 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X487 VSS cs_ring_osc_0/vosc2 freq_div_0/vin VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X488 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X489 a_31113_8829# a_30579_8463# a_31018_8829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X490 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X491 cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X492 freq_div_0/sky130_fd_sc_hd__inv_4_4/Y freq_div_0/sky130_fd_sc_hd__inv_4_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X493 VDD a_31186_7487# a_31113_7741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X494 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X495 VDD cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_31361_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X496 cs_ring_osc_0/cs_ring_osc_stage_5/vout cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_32430_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X497 a_12074_n16656# cs_ring_osc_0/vpbias a_12532_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X498 VSS a_31443_5743# a_31611_5717# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X499 cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X500 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_30579_7925# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X501 cs_ring_osc_0/cs_ring_osc_stage_4/voutcs VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X502 VSS a_34309_6555# a_34740_6609# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X503 freq_div_0/sky130_fd_sc_hd__inv_1_10/A a_34740_5743# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X504 a_31113_7741# a_30579_7375# a_31018_7741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X505 a_33614_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/vin cs_ring_osc_0/cs_ring_osc_stage_4/voutcs VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X506 VDD a_34309_7893# a_34740_7919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X507 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_31611_8731# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X508 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X509 cs_ring_osc_0/cs_ring_osc_stage_1/vin cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_17431_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X510 pfd_cp_lpf_0/vQB a_28543_13935# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X511 a_27532_1344# cs_ring_osc_0/vpbias a_27990_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X512 VSS ibiasn ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X513 a_25293_7037# cs_ring_osc_0/cs_ring_osc_stage_5/vout a_24835_7037# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X514 VDD a_31186_7893# a_31113_7919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X515 a_31514_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_31056_n20414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X516 a_33443_6837# a_33277_6837# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X517 VSS a_33884_7893# a_33842_8297# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+11p ps=1.53e+06u w=420000u l=150000u
X518 a_30933_6287# freq_div_0/sky130_fd_sc_hd__inv_4_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X519 a_33631_5743# freq_div_0/sky130_fd_sc_hd__inv_4_10/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X520 VSS VSS cs_ring_osc_0/cs_ring_osc_stage_2/voutcs VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X521 VDD a_34309_6805# a_34740_6831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X522 a_15614_6217# cs_ring_osc_0/vpbias a_16072_6217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.64e+12p ps=3.316e+07u w=8e+06u l=2e+06u
X523 a_31113_7919# a_30579_7925# a_31018_7919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X524 freq_div_0/sky130_fd_sc_hd__inv_4_7/A freq_div_0/sky130_fd_sc_hd__inv_1_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X525 a_34141_6653# a_33443_6287# a_33884_6399# VSS sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=1.978e+11p ps=1.99e+06u w=360000u l=150000u
X526 a_26972_n3082# vcp a_26514_n3082# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X527 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X528 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_31611_8731# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X529 a_33716_7741# a_33277_7375# a_33631_7375# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=1.626e+11p ps=1.66e+06u w=360000u l=150000u
X530 a_27430_n3082# vcp a_26972_n3082# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X531 VDD a_31186_6805# a_31113_6831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X532 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X533 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X534 freq_div_0/sky130_fd_sc_hd__inv_4_0/Y freq_div_0/sky130_fd_sc_hd__inv_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X535 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X536 freq_div_0/sky130_fd_sc_hd__inv_4_4/A freq_div_0/sky130_fd_sc_hd__inv_1_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X537 a_30599_n921# cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_30141_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X538 a_32430_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_31972_n20414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X539 a_26158_n16656# cs_ring_osc_0/vpbias a_25700_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X540 a_31113_6831# a_30579_6837# a_31018_6831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X541 freq_div_0/sky130_fd_sc_hd__inv_4_9/Y freq_div_0/sky130_fd_sc_hd__inv_4_9/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X542 a_10598_n3082# vcp a_10140_n3082# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X543 VSS VSS cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X544 cs_ring_osc_0/cs_ring_osc_stage_2/csinvn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X545 a_33842_7375# a_33443_7375# a_33716_7741# VSS sky130_fd_pr__nfet_01v8 ad=1.392e+11p pd=1.53e+06u as=0p ps=0u w=360000u l=150000u
X546 a_10700_1344# cs_ring_osc_0/vpbias a_10242_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=0p ps=0u w=8e+06u l=2e+06u
X547 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X548 a_11515_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/vin a_11057_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X549 a_30904_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_30446_n6542# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X550 VDD freq_div_0/sky130_fd_sc_hd__inv_4_7/A freq_div_0/sky130_fd_sc_hd__inv_4_7/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X551 cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X552 a_33631_7919# freq_div_0/sky130_fd_sc_hd__inv_4_6/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.626e+11p pd=1.66e+06u as=0p ps=0u w=420000u l=150000u
X553 a_26158_1344# cs_ring_osc_0/vpbias a_25700_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X554 a_27074_n16656# cs_ring_osc_0/vpbias a_26616_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X555 a_30306_n11700# cs_ring_osc_0/vpbias a_30764_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X556 a_30745_6837# a_30579_6837# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X557 a_26158_1344# cs_ring_osc_0/vpbias a_26616_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X558 VSS VSS pfd_cp_lpf_0/vndiode VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X559 a_30306_n11700# cs_ring_osc_0/vpbias a_29848_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X560 ibiasn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X561 VSS a_33884_7487# a_33842_7375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X562 a_30933_5743# freq_div_0/sky130_fd_sc_hd__inv_4_5/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X563 VSS vcp a_27430_n3082# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X564 a_10140_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/vin a_9682_n20414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X565 a_31443_6653# a_30745_6287# a_31186_6399# VSS sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=1.978e+11p ps=1.99e+06u w=360000u l=150000u
X566 a_28065_13961# a_28021_14203# a_27899_13961# VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X567 cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X568 a_12431_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/vin a_11973_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=2e+06u
X569 VDD VDD cs_ring_osc_0/vosc VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X570 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X571 a_16515_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_16057_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X572 freq_div_0/sky130_fd_sc_hd__inv_1_7/A a_34740_7697# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X573 cs_ring_osc_0/cs_ring_osc_stage_5/csinvn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X574 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X575 cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X576 a_27990_n16656# cs_ring_osc_0/vpbias a_27532_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X577 a_27803_13961# a_27453_13961# a_27708_13961# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X578 a_11616_1344# cs_ring_osc_0/vpbias a_12074_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X579 a_27803_13961# a_27287_13961# a_27708_13961# VSS sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=0p ps=0u w=360000u l=150000u
X580 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N a_29107_13961# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X581 freq_div_0/sky130_fd_sc_hd__inv_4_0/A freq_div_0/sky130_fd_sc_hd__inv_1_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X582 freq_div_0/sky130_fd_sc_hd__inv_4_4/Y freq_div_0/sky130_fd_sc_hd__inv_4_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X583 a_30745_8463# a_30579_8463# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X584 a_30391_13935# a_30762_14213# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X585 a_30598_n2414# cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_30140_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X586 VSS ibiasn pfd_cp_lpf_0/vswitchl VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X587 a_33884_5717# a_33716_5743# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.978e+11p pd=1.99e+06u as=0p ps=0u w=640000u l=150000u
X588 a_17431_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_16973_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X589 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X590 VDD a_34141_6653# a_34309_6555# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X591 a_10599_n921# cs_ring_osc_0/vosc a_10141_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X592 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X593 a_30933_7919# freq_div_0/sky130_fd_sc_hd__inv_4_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X594 a_33884_7893# a_33716_7919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X595 VDD freq_div_0/sky130_fd_sc_hd__inv_4_3/A freq_div_0/sky130_fd_sc_hd__inv_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X596 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X597 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X598 cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X599 ibiasn ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X600 a_33631_7375# freq_div_0/sky130_fd_sc_hd__inv_4_7/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X601 a_26209_7037# cs_ring_osc_0/cs_ring_osc_stage_5/vout a_25751_7037# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=2e+06u
X602 VDD a_28368_13961# a_28543_13935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X603 a_33884_6805# a_33716_6831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X604 a_26057_n921# cs_ring_osc_0/cs_ring_osc_stage_5/vin a_25599_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X605 a_34141_7741# a_33277_7375# a_33884_7487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X606 VSS a_34141_6653# a_34309_6555# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X607 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X608 a_31798_14327# a_31040_14229# a_31235_14198# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X609 a_17138_n11700# cs_ring_osc_0/vpbias a_16680_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=4.64e+12p pd=3.316e+07u as=0p ps=0u w=8e+06u l=2e+06u
X610 VSS pfd_cp_lpf_0/vRSTN a_28065_13961# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X611 a_24682_n3082# vcp cs_ring_osc_0/cs_ring_osc_stage_5/csinvn VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X612 VSS a_30294_13935# pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X613 VDD a_34141_7919# a_34309_7893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X614 freq_div_0/sky130_fd_sc_hd__inv_4_6/Y freq_div_0/sky130_fd_sc_hd__inv_4_6/A VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X615 a_12074_1344# cs_ring_osc_0/vpbias a_11616_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X616 a_31973_n921# cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_31515_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X617 cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X618 freq_div_0/sky130_fd_sc_hd__inv_4_0/Y freq_div_0/sky130_fd_sc_hd__inv_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X619 VSS a_31186_6805# a_31144_7209# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+11p ps=1.53e+06u w=420000u l=150000u
X620 a_31186_5717# a_31018_5743# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.978e+11p pd=1.99e+06u as=0p ps=0u w=640000u l=150000u
X621 VDD a_31443_6653# a_31611_6555# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X622 VDD a_31611_5717# a_32042_5743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X623 a_24683_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/vin cs_ring_osc_0/cs_ring_osc_stage_3/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X624 a_31186_7893# a_31018_7919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X625 cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X626 a_30933_7375# freq_div_0/sky130_fd_sc_hd__inv_4_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.626e+11p pd=1.66e+06u as=0p ps=0u w=420000u l=150000u
X627 a_30598_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_30140_n20414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X628 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X629 a_17138_n11700# cs_ring_osc_0/vpbias cs_ring_osc_0/cs_ring_osc_stage_1/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X630 a_31443_8829# a_30579_8463# a_31186_8575# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.19e+11p ps=2.15e+06u w=420000u l=150000u
X631 a_34141_7919# a_33277_7925# a_33884_7893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X632 VDD a_34141_6831# a_34309_6805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X633 a_31018_6653# a_30579_6287# a_30933_6287# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=0p ps=0u w=360000u l=150000u
X634 a_16057_n921# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_15599_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X635 VSS VSS cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X636 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X637 VDD pfd_cp_lpf_0/vQA pfd_cp_lpf_0/vRSTN VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X638 freq_div_0/sky130_fd_sc_hd__inv_4_8/Y freq_div_0/sky130_fd_sc_hd__inv_4_8/A VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X639 a_31186_8575# a_31018_8829# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X640 VDD cs_ring_osc_0/vpbias a_25242_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X641 a_31186_8575# a_31018_8829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X642 VDD freq_div_0/sky130_fd_sc_hd__inv_4_7/A freq_div_0/sky130_fd_sc_hd__inv_4_7/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X643 a_34141_6831# a_33443_6837# a_33884_6805# VSS sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=1.978e+11p ps=1.99e+06u w=360000u l=150000u
X644 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X645 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X646 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X647 a_31186_6805# a_31018_6831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X648 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X649 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X650 a_11514_n21082# vcp a_11056_n21082# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X651 a_29683_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/voutcs VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X652 a_31443_7741# a_30579_7375# a_31186_7487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X653 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_33277_7375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X654 a_31144_6287# a_30745_6287# a_31018_6653# VSS sky130_fd_pr__nfet_01v8 ad=1.392e+11p pd=1.53e+06u as=0p ps=0u w=360000u l=150000u
X655 VSS a_31443_6653# a_31611_6555# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X656 a_25598_n3082# vcp a_25140_n3082# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X657 a_16222_n11700# cs_ring_osc_0/vpbias a_16680_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X658 VSS freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_33277_7925# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X659 a_34141_6831# a_33277_6837# a_33884_6805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X660 a_19072_n5874# vcp a_18614_n5874# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X661 VDD a_31443_7919# a_31611_7893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X662 ibiasn ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X663 a_19530_n5874# vcp a_19072_n5874# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X664 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y freq_div_0/sky130_fd_sc_hd__inv_4_1/A VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X665 a_34141_5743# a_33443_5749# a_33884_5717# VSS sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=0p ps=0u w=360000u l=150000u
X666 a_31057_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_30599_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X667 a_10599_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/vin a_10141_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X668 VDD a_31611_8731# a_31527_8829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X669 VSS freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q a_30579_6837# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X670 VSS a_31186_6399# a_31144_6287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X671 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q a_33277_5749# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X672 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X673 a_12430_n21082# vcp a_11972_n21082# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X674 VDD a_31443_6831# a_31611_6805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X675 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X676 freq_div_0/vin cs_ring_osc_0/vosc2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X677 a_31443_7919# a_30579_7925# a_31186_7893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X678 a_11973_n921# cs_ring_osc_0/vosc a_11515_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X679 cs_ring_osc_0/cs_ring_osc_stage_0/csinvn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X680 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X681 VDD pfd_cp_lpf_0/vpbias pfd_cp_lpf_0/vswitchh VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X682 freq_div_0/sky130_fd_sc_hd__inv_4_2/Y freq_div_0/sky130_fd_sc_hd__inv_4_2/A VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X683 a_16530_6217# cs_ring_osc_0/vpbias a_16072_6217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X684 VDD a_31611_7643# a_31527_7741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X685 a_31443_6831# a_30745_6837# a_31186_6805# VSS sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=1.978e+11p ps=1.99e+06u w=360000u l=150000u
X686 a_11056_n3082# vcp a_10598_n3082# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X687 a_31973_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_31515_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X688 VDD freq_div_0/sky130_fd_sc_hd__inv_4_3/A freq_div_0/sky130_fd_sc_hd__inv_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X689 a_11514_n3082# vcp a_11056_n3082# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X690 a_15599_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_15141_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X691 VDD cs_ring_osc_0/vpbias a_14390_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X692 cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X693 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X694 a_31443_6831# a_30579_6837# a_31186_6805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X695 a_19988_n5874# vcp a_19530_n5874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X696 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X697 freq_div_0/sky130_fd_sc_hd__inv_1_3/A a_32042_7697# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X698 freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q a_34309_5717# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X699 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X700 a_26667_7037# cs_ring_osc_0/cs_ring_osc_stage_5/vout a_26209_7037# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X701 VSS freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_33277_7375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X702 VSS freq_div_0/sky130_fd_sc_hd__inv_4_10/A freq_div_0/sky130_fd_sc_hd__inv_4_10/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X703 VSS VSS pfd_cp_lpf_0/vswitchl VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X704 a_27124_9468# cs_ring_osc_0/cs_ring_osc_stage_5/vout a_26666_9468# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X705 a_31443_5743# a_30745_5749# a_31186_5717# VSS sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=0p ps=0u w=360000u l=150000u
X706 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X707 VDD a_31611_7643# a_32042_7697# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X708 cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X709 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X710 freq_div_0/sky130_fd_sc_hd__inv_4_1/A freq_div_0/sky130_fd_sc_hd__inv_1_1/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X711 VDD a_31611_7893# a_31527_7919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X712 VSS freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q a_30579_6287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X713 cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X714 pfd_cp_lpf_0/vswitchh pfd_cp_lpf_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X715 freq_div_0/sky130_fd_sc_hd__inv_4_6/Y freq_div_0/sky130_fd_sc_hd__inv_4_6/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X716 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X717 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X718 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X719 pfd_cp_lpf_0/vpbias VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X720 a_17904_9468# vcp a_17446_9468# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X721 freq_div_0/sky130_fd_sc_hd__inv_4_10/Y freq_div_0/sky130_fd_sc_hd__inv_4_10/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X722 a_19071_n9035# cs_ring_osc_0/cs_ring_osc_stage_1/vin a_18613_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X723 pfd_cp_lpf_0/vswitchl VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X724 VDD a_31611_6805# a_31527_6831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X725 freq_div_0/sky130_fd_sc_hd__inv_4_2/A freq_div_0/sky130_fd_sc_hd__inv_1_2/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X726 a_31056_n2414# cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_30598_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X727 a_31514_n2414# cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_31056_n2414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X728 a_14682_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X729 pfd_cp_lpf_0/vpdiode pfd_cp_lpf_0/VQBb pfd_cp_lpf_0/vswitchl VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X730 freq_div_0/sky130_fd_sc_hd__inv_4_8/Y freq_div_0/sky130_fd_sc_hd__inv_4_8/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X731 freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q a_31611_5717# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X732 a_24682_n21082# vcp cs_ring_osc_0/cs_ring_osc_stage_3/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X733 a_33443_6287# a_33277_6287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X734 VSS freq_div_0/sky130_fd_sc_hd__inv_4_5/A freq_div_0/sky130_fd_sc_hd__inv_4_5/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X735 cs_ring_osc_0/cs_ring_osc_stage_5/csinvp VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X736 a_26616_n16656# cs_ring_osc_0/vpbias a_26158_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X737 a_30764_n11700# cs_ring_osc_0/vpbias a_31222_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X738 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X739 a_27990_1344# cs_ring_osc_0/vpbias a_27532_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X740 pfd_cp_lpf_0/vswitchh pfd_cp_lpf_0/vQAb vcp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X741 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X742 cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X743 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X744 freq_div_0/sky130_fd_sc_hd__inv_4_9/A freq_div_0/sky130_fd_sc_hd__inv_1_9/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X745 a_31798_14327# a_31079_14103# a_31235_14198# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X746 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y freq_div_0/sky130_fd_sc_hd__inv_4_1/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X747 a_31018_6831# a_30579_6837# a_30933_6831# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=0p ps=0u w=360000u l=150000u
X748 VSS a_33884_5717# a_33842_6121# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X749 cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X750 cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X751 a_25140_n3082# vcp a_24682_n3082# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X752 a_27532_n16656# cs_ring_osc_0/vpbias a_27074_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X753 a_19987_n9035# cs_ring_osc_0/cs_ring_osc_stage_1/vin a_19529_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X754 VDD cs_ring_osc_0/vosc2 freq_div_0/vin VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X755 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y freq_div_0/sky130_fd_sc_hd__inv_4_5/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X756 a_15141_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_14683_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X757 a_10242_1344# cs_ring_osc_0/vpbias a_10700_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X758 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs cs_ring_osc_0/cs_ring_osc_stage_3/vin a_27431_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X759 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X760 a_16361_n9035# cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_15903_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X761 a_10598_n21082# vcp a_10140_n21082# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X762 a_31144_7209# a_30745_6837# a_31018_6831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X763 freq_div_0/sky130_fd_sc_hd__inv_4_2/Y freq_div_0/sky130_fd_sc_hd__inv_4_2/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X764 a_30745_6287# a_30579_6287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X765 a_31018_5743# a_30579_5749# a_30933_5743# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=1.626e+11p ps=1.66e+06u w=360000u l=150000u
X766 freq_div_0/sky130_fd_sc_hd__inv_4_6/A freq_div_0/sky130_fd_sc_hd__inv_1_6/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X767 cs_ring_osc_0/vosc cs_ring_osc_0/cs_ring_osc_stage_5/vout a_27583_7037# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X768 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X769 pfd_cp_lpf_0/vswitchl VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X770 VSS a_34141_7919# a_34309_7893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X771 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X772 a_26056_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/vin a_25598_n20414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X773 a_31144_6121# a_30745_5749# a_31018_5743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X774 a_33631_5743# freq_div_0/sky130_fd_sc_hd__inv_4_10/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X775 VSS freq_div_0/sky130_fd_sc_hd__inv_4_10/A freq_div_0/sky130_fd_sc_hd__inv_4_10/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X776 cs_ring_osc_0/cs_ring_osc_stage_2/csinvp cs_ring_osc_0/vpbias a_12990_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X777 vcp VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X778 VSS vcp a_18820_9468# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X779 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y freq_div_0/sky130_fd_sc_hd__inv_4_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X780 a_34267_6287# a_33277_6287# a_34141_6653# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X781 a_26056_n3082# vcp a_25598_n3082# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X782 VSS a_34309_6805# a_34267_7209# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X783 freq_div_0/sky130_fd_sc_hd__inv_4_8/A freq_div_0/sky130_fd_sc_hd__inv_1_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X784 a_26514_n3082# vcp a_26056_n3082# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X785 cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X786 a_14698_6217# cs_ring_osc_0/vpbias a_14240_6217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X787 freq_div_0/sky130_fd_sc_hd__inv_1_9/A a_34740_6609# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X788 a_27582_9468# cs_ring_osc_0/cs_ring_osc_stage_5/vout a_27124_9468# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X789 VSS a_34141_6831# a_34309_6805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X790 cs_ring_osc_0/cs_ring_osc_stage_0/csinvp cs_ring_osc_0/vpbias a_12990_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X791 cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X792 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X793 VDD pfd_cp_lpf_0/vpbias pfd_cp_lpf_0/vswitchh VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X794 VSS a_34309_7893# a_34740_7919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X795 a_26972_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/vin a_26514_n20414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X796 VSS pfd_cp_lpf_0/vQA pfd_cp_lpf_0/vQAb VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X797 freq_div_0/sky130_fd_sc_hd__inv_4_5/A freq_div_0/sky130_fd_sc_hd__inv_1_5/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X798 freq_div_0/sky130_fd_sc_hd__inv_4_10/Y freq_div_0/sky130_fd_sc_hd__inv_4_10/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X799 VSS a_28543_13935# a_29107_13961# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X800 a_19072_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/vin a_18614_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X801 a_19530_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/vin a_19072_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X802 VSS a_31443_7919# a_31611_7893# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X803 a_27990_1344# cs_ring_osc_0/vpbias cs_ring_osc_0/cs_ring_osc_stage_5/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X804 a_24835_7037# cs_ring_osc_0/cs_ring_osc_stage_5/vout VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X805 a_33631_7375# freq_div_0/sky130_fd_sc_hd__inv_4_7/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X806 VDD pfd_cp_lpf_0/vRSTN a_30391_13935# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X807 freq_div_0/sky130_fd_sc_hd__inv_1_6/A a_34740_7919# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X808 a_30933_5743# freq_div_0/sky130_fd_sc_hd__inv_4_5/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X809 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X810 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X811 a_27453_13961# a_27287_13961# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X812 VSS freq_div_0/sky130_fd_sc_hd__inv_4_5/A freq_div_0/sky130_fd_sc_hd__inv_4_5/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X813 VDD VDD pfd_cp_lpf_0/vndiode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X814 a_27911_14327# a_27287_13961# a_27803_13961# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X815 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y freq_div_0/sky130_fd_sc_hd__inv_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X816 VDD a_34309_6555# a_34740_6609# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X817 cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X818 a_31569_6287# a_30579_6287# a_31443_6653# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X819 a_16680_n11700# cs_ring_osc_0/vpbias a_17138_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X820 VSS a_31611_6805# a_31569_7209# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X821 VSS VSS cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X822 VSS a_34309_6555# a_34267_6287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X823 freq_div_0/sky130_fd_sc_hd__inv_1_5/A a_32042_5743# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X824 a_24683_n921# cs_ring_osc_0/cs_ring_osc_stage_5/vin cs_ring_osc_0/cs_ring_osc_stage_5/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X825 cs_ring_osc_0/cs_ring_osc_stage_2/voutcs cs_ring_osc_0/cs_ring_osc_stage_2/vin a_12430_n20414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X826 VSS a_31443_6831# a_31611_6805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X827 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X828 VSS a_34309_7643# a_34740_7697# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X829 freq_div_0/sky130_fd_sc_hd__inv_1_8/A a_34740_6831# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X830 a_30933_8463# freq_div_0/sky130_fd_sc_hd__inv_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X831 a_33631_7919# freq_div_0/sky130_fd_sc_hd__inv_4_6/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X832 VSS freq_div_0/sky130_fd_sc_hd__inv_4_9/A freq_div_0/sky130_fd_sc_hd__inv_4_9/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X833 a_19988_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/vin a_19530_n6542# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X834 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y freq_div_0/sky130_fd_sc_hd__inv_4_5/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X835 cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X836 a_14071_n9035# cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_13613_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X837 a_33443_7925# a_33277_7925# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X838 freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q a_34309_5717# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X839 a_16362_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_15904_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X840 cs_ring_osc_0/cs_ring_osc_stage_3/vin cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_17430_n20414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X841 a_30933_7375# freq_div_0/sky130_fd_sc_hd__inv_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X842 VSS cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_16362_n6542# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X843 VSS vcp a_27430_n21082# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X844 a_31515_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_31057_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X845 a_33631_6831# freq_div_0/sky130_fd_sc_hd__inv_4_8/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X846 a_14683_n921# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X847 a_14390_n11700# cs_ring_osc_0/vpbias a_14848_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X848 a_34141_7741# a_33443_7375# a_33884_7487# VSS sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=0p ps=0u w=360000u l=150000u
X849 VDD VDD cs_ring_osc_0/cs_ring_osc_stage_2/voutcs VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X850 pfd_cp_lpf_0/vpbias pfd_cp_lpf_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X851 VDD a_28543_13935# a_29107_13961# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X852 a_33716_6653# a_33443_6287# a_33631_6287# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X853 VSS a_31611_6555# a_31569_6287# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X854 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X855 a_29848_n11700# cs_ring_osc_0/vpbias a_29390_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X856 freq_div_0/sky130_fd_sc_hd__inv_4_3/A freq_div_0/sky130_fd_sc_hd__inv_1_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X857 a_9682_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/vin cs_ring_osc_0/cs_ring_osc_stage_2/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X858 a_32431_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_31973_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X859 a_16072_6217# cs_ring_osc_0/vpbias a_15614_6217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X860 a_30141_n921# cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_29683_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X861 a_14240_6217# cs_ring_osc_0/vpbias a_14698_6217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X862 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y freq_div_0/sky130_fd_sc_hd__inv_4_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X863 a_30933_7919# freq_div_0/sky130_fd_sc_hd__inv_4_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X864 VSS freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q a_33277_5749# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X865 a_12074_1344# cs_ring_osc_0/vpbias a_12532_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X866 VDD VDD cs_ring_osc_0/cs_ring_osc_stage_3/vin VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X867 VSS freq_div_0/sky130_fd_sc_hd__inv_4_4/A freq_div_0/sky130_fd_sc_hd__inv_4_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X868 cs_ring_osc_0/cs_ring_osc_stage_2/csinvp VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X869 VDD freq_div_0/vout a_27287_13961# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X870 a_14987_n9035# cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_14529_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X871 VSS pfd_cp_lpf_0/vRSTN a_30797_13961# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X872 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X873 a_15445_n9035# cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_14987_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=2e+06u
X874 ibiasn ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X875 freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q a_31611_5717# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X876 cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X877 a_30745_7925# a_30579_7925# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X878 a_30933_6831# freq_div_0/sky130_fd_sc_hd__inv_4_2/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X879 a_31443_7741# a_30745_7375# a_31186_7487# VSS sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=0p ps=0u w=360000u l=150000u
X880 VDD a_33884_6399# a_33811_6653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X881 a_32138_n11700# cs_ring_osc_0/vpbias a_31680_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X882 VSS a_31611_6805# a_32042_6831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X883 a_10141_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/vin a_9683_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X884 cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X885 a_34267_7209# a_33277_6837# a_34141_6831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X886 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X887 a_31018_6653# a_30745_6287# a_30933_6287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X888 a_33716_5743# a_33443_5749# a_33631_5743# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X889 a_33811_6653# a_33277_6287# a_33716_6653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X890 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X891 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y freq_div_0/sky130_fd_sc_hd__inv_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X892 a_18614_n5874# vcp VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X893 a_25750_9468# cs_ring_osc_0/cs_ring_osc_stage_5/vout a_25292_9468# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X894 a_11616_1344# cs_ring_osc_0/vpbias a_11158_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X895 a_25242_n16656# cs_ring_osc_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X896 a_32138_n11700# cs_ring_osc_0/vpbias cs_ring_osc_0/cs_ring_osc_stage_4/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X897 a_33884_6805# a_33716_6831# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X898 a_34267_6121# a_33277_5749# a_34141_5743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X899 a_31515_n921# cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_31057_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X900 VDD a_34141_7741# a_34309_7643# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X901 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X902 pfd_cp_lpf_0/vswitchh pfd_cp_lpf_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X903 VDD freq_div_0/sky130_fd_sc_hd__inv_4_0/A freq_div_0/sky130_fd_sc_hd__inv_4_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X904 cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X905 a_33716_7919# a_33277_7925# a_33631_7919# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=0p ps=0u w=360000u l=150000u
X906 a_30762_14213# a_31040_14229# a_30996_14327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X907 VSS freq_div_0/sky130_fd_sc_hd__inv_4_9/A freq_div_0/sky130_fd_sc_hd__inv_4_9/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X908 pfd_cp_lpf_0/vswitchh pfd_cp_lpf_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X909 a_16530_9468# vcp a_16072_9468# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X910 a_31222_n11700# cs_ring_osc_0/vpbias a_31680_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X911 VSS a_31611_6555# a_32042_6609# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X912 VDD a_33884_5717# a_33811_5743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X913 a_14072_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_13614_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X914 cs_ring_osc_0/cs_ring_osc_stage_1/csinvp cs_ring_osc_0/vpbias a_17138_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X915 ibiasn ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X916 a_31569_7209# a_30579_6837# a_31443_6831# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X917 a_14530_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_14072_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X918 a_33842_8297# a_33443_7925# a_33716_7919# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X919 VDD a_31611_7893# a_32042_7919# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X920 VSS a_34141_7741# a_34309_7643# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X921 a_31018_5743# a_30745_5749# a_30933_5743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X922 pfd_cp_lpf_0/vswitchh VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X923 VSS VSS ibiasn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X924 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X925 a_33811_5743# a_33277_5749# a_33716_5743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X926 a_10700_1344# cs_ring_osc_0/vpbias a_11158_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X927 a_11158_n16656# cs_ring_osc_0/vpbias a_10700_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X928 a_29071_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_28613_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X929 VDD cs_ring_osc_0/vosc2 freq_div_0/vin VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X930 VSS a_31186_7893# a_31144_8297# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X931 a_31186_6805# a_31018_6831# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X932 a_31569_6121# a_30579_5749# a_31443_5743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X933 cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X934 VDD a_31443_7741# a_31611_7643# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X935 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X936 VDD a_31611_6805# a_32042_6831# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X937 a_34225_6653# a_33443_6287# a_34141_6653# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=0p ps=0u w=420000u l=150000u
X938 a_10242_1344# cs_ring_osc_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X939 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X940 cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X941 VDD a_30391_13935# pfd_cp_lpf_0/vQA VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X942 a_30933_8463# freq_div_0/sky130_fd_sc_hd__inv_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X943 a_31018_7741# a_30579_7375# a_30933_7375# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=0p ps=0u w=360000u l=150000u
X944 cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X945 a_29765_13961# pfd_cp_lpf_0/vQB VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X946 VDD VDD a_31798_14327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X947 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X948 a_30599_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_30141_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X949 VSS freq_div_0/sky130_fd_sc_hd__inv_4_4/A freq_div_0/sky130_fd_sc_hd__inv_4_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X950 a_12074_n16656# cs_ring_osc_0/vpbias a_11616_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X951 a_11515_n921# cs_ring_osc_0/vosc a_11057_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=2e+06u
X952 a_26514_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/vin a_26056_n20414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X953 a_15306_n11700# cs_ring_osc_0/vpbias a_14848_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X954 VDD freq_div_0/vin a_30579_8463# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X955 a_14988_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_14530_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X956 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=2e+06u
X957 a_15446_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_14988_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X958 a_18613_n9035# cs_ring_osc_0/cs_ring_osc_stage_1/vin cs_ring_osc_0/cs_ring_osc_stage_1/voutcs VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X959 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_34309_6555# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X960 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X961 cs_ring_osc_0/cs_ring_osc_stage_2/csinvn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X962 a_31473_13961# pfd_cp_lpf_0/vRSTN VSS VSS sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X963 a_31144_7375# a_30745_7375# a_31018_7741# VSS sky130_fd_pr__nfet_01v8 ad=1.392e+11p pd=1.53e+06u as=0p ps=0u w=360000u l=150000u
X964 VSS a_31443_7741# a_31611_7643# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X965 freq_div_0/sky130_fd_sc_hd__inv_1_4/A a_32042_6609# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X966 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X967 a_12990_n16656# cs_ring_osc_0/vpbias a_12532_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X968 a_29987_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_29529_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X969 VDD pfd_cp_lpf_0/vpdiode pfd_cp_lpf_0/vpdiode VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X970 a_27430_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/vin a_26972_n20414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X971 a_16222_n11700# cs_ring_osc_0/vpbias a_15764_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X972 a_28368_13961# a_27287_13961# a_28021_14203# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X973 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q a_30579_7375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X974 cs_ring_osc_0/cs_ring_osc_stage_5/vout cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_32431_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X975 VSS freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_30579_7925# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X976 a_14240_6217# cs_ring_osc_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X977 VSS a_31186_7487# a_31144_7375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X978 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_33277_6837# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X979 a_10140_n21082# vcp a_9682_n21082# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X980 a_27899_13961# a_27453_13961# a_27803_13961# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X981 a_31527_6653# a_30745_6287# a_31443_6653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X982 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_34309_6555# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X983 VDD cs_ring_osc_0/vpbias a_10242_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X984 a_34225_5743# a_33443_5749# a_34141_5743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X985 freq_div_0/sky130_fd_sc_hd__inv_4_9/Y freq_div_0/sky130_fd_sc_hd__inv_4_9/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X986 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X987 freq_div_0/vout a_34309_7893# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X988 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_30579_5749# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X989 pfd_cp_lpf_0/VQBb pfd_cp_lpf_0/vQB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X990 VSS freq_div_0/sky130_fd_sc_hd__inv_4_6/A freq_div_0/sky130_fd_sc_hd__inv_4_6/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X991 cs_ring_osc_0/cs_ring_osc_stage_5/csinvn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X992 cs_ring_osc_0/vosc2 cs_ring_osc_0/vosc VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X993 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X994 VDD freq_div_0/sky130_fd_sc_hd__inv_4_0/A freq_div_0/sky130_fd_sc_hd__inv_4_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X995 a_33443_6837# a_33277_6837# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X996 a_9682_n2414# cs_ring_osc_0/vosc cs_ring_osc_0/cs_ring_osc_stage_0/csinvn VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X997 a_19529_n9035# cs_ring_osc_0/cs_ring_osc_stage_1/vin a_19071_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X998 VDD a_28021_14203# a_27911_14327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X999 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_31611_6555# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1000 a_10141_n921# cs_ring_osc_0/vosc a_9683_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1001 cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1002 a_15903_n9035# cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_15445_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1003 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_34309_6805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1004 VSS a_34309_5717# a_34740_5743# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1005 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1006 freq_div_0/sky130_fd_sc_hd__inv_1_0/A a_32042_8785# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1007 VSS freq_div_0/sky130_fd_sc_hd__inv_4_8/A freq_div_0/sky130_fd_sc_hd__inv_4_8/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1008 a_16972_n2414# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_16514_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X1009 a_31545_13961# a_31166_14327# a_31473_13961# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1010 a_17430_n2414# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_16972_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X1011 VDD pfd_cp_lpf_0/vpbias pfd_cp_lpf_0/vpbias VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1012 VDD a_31611_8731# a_32042_8785# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1013 freq_div_0/sky130_fd_sc_hd__inv_4_6/Y freq_div_0/sky130_fd_sc_hd__inv_4_6/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1014 VSS freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q a_30579_7375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1015 a_27532_1344# cs_ring_osc_0/vpbias a_27074_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1016 cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1017 cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1018 pfd_cp_lpf_0/vpdiode VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1019 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_31611_6555# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1020 a_31527_5743# a_30745_5749# a_31443_5743# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1021 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1022 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1023 cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1024 pfd_cp_lpf_0/vQB a_28543_13935# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1025 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q a_31611_7893# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1026 freq_div_0/sky130_fd_sc_hd__inv_4_4/Y freq_div_0/sky130_fd_sc_hd__inv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1027 cs_ring_osc_0/cs_ring_osc_stage_0/voutcs cs_ring_osc_0/vosc a_12431_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1028 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1029 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1030 a_29072_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_28614_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X1031 VSS freq_div_0/sky130_fd_sc_hd__inv_4_1/A freq_div_0/sky130_fd_sc_hd__inv_4_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1032 freq_div_0/sky130_fd_sc_hd__inv_4_8/Y freq_div_0/sky130_fd_sc_hd__inv_4_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1033 a_29530_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_29072_n6542# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X1034 cs_ring_osc_0/vpbias cs_ring_osc_0/vpbias a_16988_6217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1035 a_30745_6837# a_30579_6837# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1036 a_33443_6287# a_33277_6287# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1037 VDD cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_16361_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1038 a_30797_13961# a_30762_14213# a_30391_13935# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1039 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q a_31611_6805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1040 cs_ring_osc_0/cs_ring_osc_stage_1/vin cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_17430_n2414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1041 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1042 a_27532_n16656# cs_ring_osc_0/vpbias a_27990_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1043 a_14683_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1044 VSS freq_div_0/sky130_fd_sc_hd__inv_4_2/A freq_div_0/sky130_fd_sc_hd__inv_4_2/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1045 VDD VDD cs_ring_osc_0/cs_ring_osc_stage_5/voutcs VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1046 VDD pfd_cp_lpf_0/vpbias pfd_cp_lpf_0/vpbias VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1047 freq_div_0/vin cs_ring_osc_0/vosc2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1048 a_21362_n5874# vcp a_20904_n5874# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X1049 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X1050 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y freq_div_0/sky130_fd_sc_hd__inv_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1051 cs_ring_osc_0/cs_ring_osc_stage_1/csinvn vcp a_21362_n5874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1052 a_18614_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/vin cs_ring_osc_0/cs_ring_osc_stage_1/voutcs VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1053 a_29390_n11700# cs_ring_osc_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1054 a_12532_1344# cs_ring_osc_0/vpbias a_12990_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1055 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1056 VSS VSS pfd_cp_lpf_0/vpdiode VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1057 freq_div_0/sky130_fd_sc_hd__inv_4_7/A freq_div_0/sky130_fd_sc_hd__inv_1_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1058 cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1059 cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1060 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1061 a_26616_n16656# cs_ring_osc_0/vpbias a_27074_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1062 a_29988_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_29530_n6542# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1063 a_27911_14327# pfd_cp_lpf_0/vRSTN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1064 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1065 freq_div_0/sky130_fd_sc_hd__inv_4_2/Y freq_div_0/sky130_fd_sc_hd__inv_4_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1066 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1067 a_25598_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/vin a_25140_n20414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X1068 VDD VDD pfd_cp_lpf_0/vswitchh VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1069 freq_div_0/sky130_fd_sc_hd__inv_4_4/A freq_div_0/sky130_fd_sc_hd__inv_1_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1070 VDD VDD cs_ring_osc_0/cs_ring_osc_stage_1/vin VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1071 a_27431_n921# cs_ring_osc_0/cs_ring_osc_stage_5/vin a_26973_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1072 a_30745_6287# a_30579_6287# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1073 freq_div_0/sky130_fd_sc_hd__inv_4_9/Y freq_div_0/sky130_fd_sc_hd__inv_4_9/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1074 cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1075 pfd_cp_lpf_0/vswitchh pfd_cp_lpf_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1076 VSS freq_div_0/sky130_fd_sc_hd__inv_4_6/A freq_div_0/sky130_fd_sc_hd__inv_4_6/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1077 a_27708_13961# VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1078 VDD a_31235_14198# a_31166_14327# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1079 VSS VSS cs_ring_osc_0/cs_ring_osc_stage_1/csinvn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1080 VDD freq_div_0/sky130_fd_sc_hd__inv_4_10/A freq_div_0/sky130_fd_sc_hd__inv_4_10/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1081 cs_ring_osc_0/cs_ring_osc_stage_2/vin VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=2e+06u
X1082 a_25700_n16656# cs_ring_osc_0/vpbias a_25242_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1083 a_31680_n11700# cs_ring_osc_0/vpbias a_32138_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1084 a_13613_n9035# cs_ring_osc_0/cs_ring_osc_stage_1/voutcs cs_ring_osc_0/cs_ring_osc_stage_2/vin VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1085 a_33884_6399# a_33716_6653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1086 a_33884_6399# a_33716_6653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1087 a_14682_n2414# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1088 a_15904_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_15446_n6542# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1089 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1090 a_25292_9468# cs_ring_osc_0/cs_ring_osc_stage_5/vout a_24834_9468# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1091 freq_div_0/sky130_fd_sc_hd__inv_4_1/A freq_div_0/sky130_fd_sc_hd__inv_1_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1092 a_11158_1344# cs_ring_osc_0/vpbias a_10700_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1093 a_17431_n921# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_16973_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1094 a_31057_n921# cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_30599_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1095 a_26057_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/vin a_25599_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1096 a_10700_n16656# cs_ring_osc_0/vpbias a_11158_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1097 VSS freq_div_0/sky130_fd_sc_hd__inv_4_8/A freq_div_0/sky130_fd_sc_hd__inv_4_8/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1098 a_34267_7375# a_33277_7375# a_34141_7741# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X1099 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1100 freq_div_0/sky130_fd_sc_hd__inv_4_6/Y freq_div_0/sky130_fd_sc_hd__inv_4_6/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1101 VSS a_34309_7893# a_34267_8297# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1102 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1103 freq_div_0/sky130_fd_sc_hd__inv_1_7/A a_34740_7697# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1104 a_30996_14327# a_30391_13935# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1105 cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1106 a_21361_n9035# cs_ring_osc_0/cs_ring_osc_stage_1/vin a_20903_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1107 freq_div_0/sky130_fd_sc_hd__inv_4_2/A freq_div_0/sky130_fd_sc_hd__inv_1_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1108 a_16072_9468# vcp cs_ring_osc_0/vpbias VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1109 a_16072_6217# cs_ring_osc_0/vpbias a_16530_6217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1110 freq_div_0/sky130_fd_sc_hd__inv_4_4/Y freq_div_0/sky130_fd_sc_hd__inv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1111 a_26973_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/vin a_26515_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1112 cs_ring_osc_0/cs_ring_osc_stage_4/vin cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_32430_n20414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1113 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1114 VSS freq_div_0/sky130_fd_sc_hd__inv_4_1/A freq_div_0/sky130_fd_sc_hd__inv_4_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1115 freq_div_0/sky130_fd_sc_hd__inv_4_8/Y freq_div_0/sky130_fd_sc_hd__inv_4_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1116 cs_ring_osc_0/cs_ring_osc_stage_3/csinvn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1117 a_14848_n11700# cs_ring_osc_0/vpbias a_15306_n11700# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1118 freq_div_0/vin cs_ring_osc_0/vosc2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1119 VDD freq_div_0/sky130_fd_sc_hd__inv_4_5/A freq_div_0/sky130_fd_sc_hd__inv_4_5/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1120 a_28021_14203# a_27803_13961# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1121 a_31037_13961# a_30391_13935# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1122 a_11616_n16656# cs_ring_osc_0/vpbias a_11158_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1123 a_14529_n9035# cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_14071_n9035# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1124 freq_div_0/sky130_fd_sc_hd__inv_1_1/A a_32042_7919# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1125 a_31186_6399# a_31018_6653# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1126 a_15598_n2414# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_15140_n2414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1127 a_31186_6399# a_31018_6653# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1128 a_10140_n2414# cs_ring_osc_0/vosc a_9682_n2414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1129 a_27453_13961# a_27287_13961# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1130 VSS freq_div_0/sky130_fd_sc_hd__inv_4_2/A freq_div_0/sky130_fd_sc_hd__inv_4_2/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1131 freq_div_0/sky130_fd_sc_hd__inv_4_0/Y freq_div_0/sky130_fd_sc_hd__inv_4_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1132 a_11972_n2414# cs_ring_osc_0/vosc a_11514_n2414# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X1133 a_25140_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/vin a_24682_n20414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1134 pfd_cp_lpf_0/vpbias pfd_cp_lpf_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1135 a_31569_7375# a_30579_7375# a_31443_7741# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1136 a_25700_1344# cs_ring_osc_0/vpbias a_25242_1344# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1137 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1138 VSS a_31611_7893# a_31569_8297# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1139 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y freq_div_0/sky130_fd_sc_hd__inv_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1140 a_12430_n2414# cs_ring_osc_0/vosc a_11972_n2414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1141 VSS a_34309_7643# a_34267_7375# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1142 a_12532_n16656# cs_ring_osc_0/vpbias a_12074_n16656# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1143 freq_div_0/sky130_fd_sc_hd__inv_1_2/A a_32042_6831# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1144 VDD VDD cs_ring_osc_0/cs_ring_osc_stage_4/vin VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1145 VDD VDD cs_ring_osc_0/cs_ring_osc_stage_1/csinvp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1146 VSS VSS cs_ring_osc_0/vosc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1147 freq_div_0/vout a_34309_7893# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1148 a_11057_n921# cs_ring_osc_0/vosc a_10599_n921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1149 cs_ring_osc_0/cs_ring_osc_stage_2/voutcs cs_ring_osc_0/cs_ring_osc_stage_2/vin a_12431_n18921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=2e+06u
X1150 pfd_cp_lpf_0/vpbias pfd_cp_lpf_0/vpbias VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1151 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1152 ibiasn ibiasn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1153 a_15614_6217# cs_ring_osc_0/vpbias a_15156_6217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
X1154 a_36362_n5874# vcp a_35904_n5874# VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X1155 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1156 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1157 VSS freq_div_0/sky130_fd_sc_hd__inv_4_7/A freq_div_0/sky130_fd_sc_hd__inv_4_7/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1158 freq_div_0/sky130_fd_sc_hd__inv_4_2/Y freq_div_0/sky130_fd_sc_hd__inv_4_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1159 VDD a_34309_6555# a_34225_6653# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1160 a_30140_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_29682_n20414# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1161 cs_ring_osc_0/cs_ring_osc_stage_4/csinvn vcp a_36362_n5874# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
C0 VDD freq_div_0/sky130_fd_sc_hd__inv_4_10/Y 0.93fF
C1 freq_div_0/sky130_fd_sc_hd__inv_1_9/A freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.27fF
C2 VDD pfd_cp_lpf_0/vQB 0.49fF
C3 a_33277_5749# a_33884_5717# 0.37fF
C4 a_31186_8575# VDD 0.23fF
C5 VDD freq_div_0/sky130_fd_sc_hd__inv_4_4/A 0.62fF
C6 a_15599_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.03fF
C7 a_34309_7893# a_34309_7643# 0.09fF
C8 VDD a_29848_n11700# 1.55fF
C9 cs_ring_osc_0/cs_ring_osc_stage_5/vout a_27583_7037# 0.03fF
C10 a_30933_6831# a_30579_6837# 0.21fF
C11 a_31079_14103# a_31166_14327# 0.16fF
C12 a_30996_14327# a_30762_14213# 0.04fF
C13 VDD freq_div_0/sky130_fd_sc_hd__inv_4_6/Y 0.93fF
C14 pfd_cp_lpf_0/vQB a_29107_13961# 0.59fF
C15 a_31018_5743# freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 0.16fF
C16 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_31972_n2414# 0.03fF
C17 freq_div_0/sky130_fd_sc_hd__inv_1_8/A freq_div_0/sky130_fd_sc_hd__inv_4_8/Y 0.27fF
C18 a_27708_13961# a_27287_13961# 0.23fF
C19 vcp a_21362_n5874# 0.03fF
C20 pfd_cp_lpf_0/vpbias pfd_cp_lpf_0/vswitchh 0.52fF
C21 a_35903_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C22 a_34740_6609# a_34740_6831# 0.04fF
C23 a_12074_1344# a_10242_1344# 0.65fF
C24 VDD cs_ring_osc_0/cs_ring_osc_stage_4/voutcs 4.44fF
C25 freq_div_0/sky130_fd_sc_hd__inv_4_10/Y freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.08fF
C26 a_30391_13935# a_30294_13935# 0.30fF
C27 pfd_cp_lpf_0/vQA pfd_cp_lpf_0/vswitchh 0.18fF
C28 a_30762_14213# a_31166_14327# 0.13fF
C29 freq_div_0/vout freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q 0.03fF
C30 a_31443_6653# a_31443_5743# 0.07fF
C31 freq_div_0/sky130_fd_sc_hd__inv_4_10/Y a_34740_5743# 0.11fF
C32 a_30306_n11700# a_32138_n11700# 0.24fF
C33 a_31611_7893# a_31611_7643# 0.09fF
C34 a_15764_n11700# a_16680_n11700# 1.33fF
C35 a_15306_n11700# a_17138_n11700# 0.24fF
C36 VDD a_33443_7925# 0.43fF
C37 VDD freq_div_0/sky130_fd_sc_hd__inv_4_2/A 0.62fF
C38 a_29987_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs 0.03fF
C39 freq_div_0/sky130_fd_sc_hd__inv_1_0/A freq_div_0/sky130_fd_sc_hd__inv_4_0/A 0.35fF
C40 a_31018_8829# freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.16fF
C41 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q 0.38fF
C42 a_31018_6831# a_30745_6837# 0.38fF
C43 pfd_cp_lpf_0/vQAb vcp 0.08fF
C44 a_25242_n16656# cs_ring_osc_0/cs_ring_osc_stage_3/csinvp 0.08fF
C45 a_31443_7741# a_31443_6831# 0.07fF
C46 a_33277_7375# a_33716_7741# 0.63fF
C47 VDD a_10700_1344# 1.55fF
C48 a_30745_6287# a_31443_5743# 0.01fF
C49 a_33884_6399# a_33443_6287# 0.28fF
C50 a_27803_13961# a_27453_13961# 0.49fF
C51 a_33443_7375# a_33716_7741# 0.38fF
C52 cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_30904_n6542# 0.03fF
C53 VDD a_31611_8731# 0.45fF
C54 VDD freq_div_0/sky130_fd_sc_hd__inv_1_5/A 0.48fF
C55 a_16988_6217# a_16530_6217# 0.02fF
C56 cs_ring_osc_0/vpbias cs_ring_osc_0/cs_ring_osc_stage_0/csinvp 0.31fF
C57 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q a_31611_7643# 0.02fF
C58 VDD a_26616_1344# 0.69fF
C59 a_33842_8297# a_33716_7919# 0.02fF
C60 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_33277_6837# 0.51fF
C61 a_30933_6831# a_31186_6805# 0.04fF
C62 a_30579_8463# a_31018_8829# 0.63fF
C63 cs_ring_osc_0/vosc a_10598_n2414# 0.03fF
C64 VDD freq_div_0/sky130_fd_sc_hd__inv_1_9/A 0.48fF
C65 a_16222_n11700# a_14390_n11700# 0.65fF
C66 a_30579_6837# a_31018_6653# 0.02fF
C67 freq_div_0/vout a_27708_13961# 0.01fF
C68 a_32042_8785# a_31443_8829# 0.02fF
C69 a_33277_6287# a_33443_6837# 0.09fF
C70 VDD a_14240_6217# 4.03fF
C71 vcp a_25598_n3082# 0.03fF
C72 a_33716_6653# a_33884_6399# 0.59fF
C73 vcp a_25140_n21082# 0.03fF
C74 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.40fF
C75 a_31527_6653# a_31443_6653# 0.05fF
C76 a_11616_n16656# a_12990_n16656# 0.01fF
C77 cs_ring_osc_0/cs_ring_osc_stage_2/vin a_11514_n20414# 0.03fF
C78 a_31186_6399# freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.15fF
C79 a_33716_7919# a_33716_7741# 0.08fF
C80 a_15598_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.03fF
C81 a_31186_7893# a_31186_7487# 0.03fF
C82 a_30579_5749# a_30745_5749# 2.23fF
C83 cs_ring_osc_0/vpbias a_27532_1344# 0.92fF
C84 a_26209_7037# VDD 0.01fF
C85 VDD freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.91fF
C86 a_31186_6399# a_31443_6653# 0.11fF
C87 freq_div_0/vin cs_ring_osc_0/vosc2 1.01fF
C88 freq_div_0/sky130_fd_sc_hd__inv_1_5/A freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.15fF
C89 a_17138_n11700# a_16680_n11700# 0.02fF
C90 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q freq_div_0/sky130_fd_sc_hd__inv_4_8/Y 0.41fF
C91 freq_div_0/sky130_fd_sc_hd__inv_4_2/A freq_div_0/sky130_fd_sc_hd__inv_4_4/A 0.09fF
C92 VDD a_31443_6653# 0.22fF
C93 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_32431_n18921# 0.03fF
C94 a_33631_6287# freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.02fF
C95 cs_ring_osc_0/cs_ring_osc_stage_5/vout a_27125_7037# 0.03fF
C96 a_33443_7925# freq_div_0/sky130_fd_sc_hd__inv_4_6/Y 0.61fF
C97 cs_ring_osc_0/cs_ring_osc_stage_2/csinvn vcp 0.08fF
C98 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y freq_div_0/sky130_fd_sc_hd__inv_1_3/A 0.27fF
C99 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_15306_n11700# 0.22fF
C100 a_30745_6287# a_31186_6399# 0.28fF
C101 a_31443_7919# a_31527_7919# 0.05fF
C102 a_31186_8575# a_31611_8731# 0.04fF
C103 a_31611_6555# a_31186_6399# 0.04fF
C104 freq_div_0/sky130_fd_sc_hd__inv_4_0/A freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 1.64fF
C105 VDD a_30745_6287# 0.43fF
C106 a_31611_6555# VDD 0.45fF
C107 a_30745_5749# a_31186_5717# 0.28fF
C108 cs_ring_osc_0/vpbias a_32138_n11700# 0.77fF
C109 a_15156_6217# a_16072_6217# 1.98fF
C110 a_34309_5717# a_33884_5717# 0.04fF
C111 a_34141_6653# a_34309_6555# 0.67fF
C112 a_30933_7919# freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q 0.02fF
C113 a_34309_6805# a_33716_6831# 0.02fF
C114 cs_ring_osc_0/cs_ring_osc_stage_4/csinvp a_32138_n11700# 0.16fF
C115 a_30745_7375# a_30933_7375# 0.26fF
C116 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y freq_div_0/sky130_fd_sc_hd__inv_4_0/A 0.03fF
C117 vcp cs_ring_osc_0/cs_ring_osc_stage_0/csinvn 0.08fF
C118 a_30764_n11700# a_32138_n11700# 0.01fF
C119 a_33716_6831# a_33443_6837# 0.38fF
C120 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_31057_n18921# 0.03fF
C121 a_16988_6217# a_15614_6217# 0.01fF
C122 a_33884_6805# a_33277_6837# 0.37fF
C123 a_33716_6653# a_33811_6653# 0.04fF
C124 pfd_cp_lpf_0/vRSTN VDD 2.28fF
C125 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_31611_5717# 0.02fF
C126 cs_ring_osc_0/cs_ring_osc_stage_2/vin a_11057_n18921# 0.03fF
C127 a_34141_7741# a_34309_7643# 0.67fF
C128 a_31443_8829# a_31018_8829# 0.03fF
C129 pfd_cp_lpf_0/vRSTN a_28021_14203# 0.37fF
C130 a_11616_n16656# a_10700_n16656# 2.26fF
C131 VDD a_28530_14327# 0.01fF
C132 VDD freq_div_0/sky130_fd_sc_hd__inv_1_1/A 0.48fF
C133 freq_div_0/sky130_fd_sc_hd__inv_4_4/Y freq_div_0/sky130_fd_sc_hd__inv_4_4/A 1.64fF
C134 cs_ring_osc_0/cs_ring_osc_stage_1/vin a_20903_n9035# 0.03fF
C135 a_35904_n5874# vcp 0.03fF
C136 VDD pfd_cp_lpf_0/vQAb 3.39fF
C137 pfd_cp_lpf_0/vRSTN a_29107_13961# 0.10fF
C138 pfd_cp_lpf_0/vRSTN a_31079_14103# 0.86fF
C139 cs_ring_osc_0/cs_ring_osc_stage_2/vin vcp 3.55fF
C140 cs_ring_osc_0/vpbias a_14390_n11700# 0.51fF
C141 cs_ring_osc_0/vosc a_10599_n921# 0.03fF
C142 a_31611_6805# a_31611_7643# 0.09fF
C143 a_32042_5743# freq_div_0/sky130_fd_sc_hd__inv_4_5/A 0.05fF
C144 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y a_31443_7741# 0.14fF
C145 VDD a_11616_n16656# 0.69fF
C146 cs_ring_osc_0/vpbias a_27990_n16656# 0.77fF
C147 VDD a_27532_n16656# 0.09fF
C148 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_34141_6653# 0.05fF
C149 a_32042_5743# a_31611_5717# 0.31fF
C150 a_36361_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C151 VDD a_10242_1344# 0.73fF
C152 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.38fF
C153 cs_ring_osc_0/vosc a_11973_n921# 0.03fF
C154 a_27532_1344# a_25700_1344# 0.43fF
C155 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_30599_n921# 0.03fF
C156 pfd_cp_lpf_0/vndiode pfd_cp_lpf_0/vQA 0.13fF
C157 a_27803_13961# a_27708_13961# 0.13fF
C158 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q 0.04fF
C159 a_32042_7919# a_31611_7893# 0.31fF
C160 vcp a_19530_n5874# 0.03fF
C161 a_34309_6805# a_34740_6831# 0.31fF
C162 pfd_cp_lpf_0/vQA a_30294_13935# 0.59fF
C163 a_31018_6831# a_30579_6287# 0.02fF
C164 freq_div_0/vout a_27287_13961# 0.49fF
C165 pfd_cp_lpf_0/vRSTN a_30762_14213# 0.57fF
C166 cs_ring_osc_0/vosc a_11515_n921# 0.03fF
C167 a_29390_n11700# a_32138_n11700# 0.14fF
C168 cs_ring_osc_0/vpbias a_26616_n16656# 0.83fF
C169 freq_div_0/sky130_fd_sc_hd__inv_4_4/Y freq_div_0/sky130_fd_sc_hd__inv_4_2/A 0.01fF
C170 a_31018_6831# freq_div_0/sky130_fd_sc_hd__inv_4_2/Y 0.16fF
C171 a_25242_1344# a_27074_1344# 0.65fF
C172 cs_ring_osc_0/cs_ring_osc_stage_3/csinvn cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.09fF
C173 pfd_cp_lpf_0/vRSTN a_31166_14327# 0.37fF
C174 a_14683_n921# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C175 pfd_cp_lpf_0/vRSTN a_28722_13961# 0.01fF
C176 VDD a_34141_5743# 0.22fF
C177 a_30745_8463# a_31018_8829# 0.38fF
C178 cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_16056_n20414# 0.03fF
C179 pfd_cp_lpf_0/vRSTN pfd_cp_lpf_0/vQB 1.19fF
C180 a_31443_6831# a_31018_6831# 0.03fF
C181 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y a_30579_7375# 0.35fF
C182 a_30579_6837# a_30745_7375# 0.02fF
C183 vcp a_25598_n21082# 0.03fF
C184 a_12074_n16656# a_11158_n16656# 1.92fF
C185 cs_ring_osc_0/vpbias a_12074_n16656# 0.76fF
C186 a_31798_14327# a_31380_14327# 0.02fF
C187 a_32042_7919# freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 0.37fF
C188 a_30579_7925# a_31018_7919# 0.63fF
C189 a_30933_7919# a_31186_7893# 0.04fF
C190 a_30579_6837# a_30745_6837# 2.23fF
C191 VDD a_33811_7919# 0.02fF
C192 a_31144_8463# a_31018_8829# 0.02fF
C193 a_31186_7487# a_31611_7643# 0.04fF
C194 a_28368_13961# a_27453_13961# 0.29fF
C195 cs_ring_osc_0/cs_ring_osc_stage_5/vout a_26666_9468# 0.03fF
C196 a_30745_7375# a_31018_7741# 0.38fF
C197 pfd_cp_lpf_0/vQB pfd_cp_lpf_0/vQAb 0.05fF
C198 a_14698_6217# cs_ring_osc_0/vpbias 0.66fF
C199 a_33631_6287# a_33443_6287# 0.26fF
C200 VDD a_27583_7037# 0.01fF
C201 a_30933_8463# freq_div_0/vin 0.02fF
C202 a_26158_n16656# a_27990_n16656# 0.24fF
C203 a_31443_7919# a_32042_7919# 0.02fF
C204 VDD a_32042_6609# 0.37fF
C205 pfd_cp_lpf_0/vpdiode pfd_cp_lpf_0/VQBb 0.10fF
C206 freq_div_0/sky130_fd_sc_hd__inv_4_7/A freq_div_0/sky130_fd_sc_hd__inv_1_7/A 0.35fF
C207 cs_ring_osc_0/cs_ring_osc_stage_5/vout a_26208_9468# 0.03fF
C208 VDD a_32042_6831# 0.37fF
C209 vcp a_35446_n5874# 0.03fF
C210 a_34141_7741# a_33716_7741# 0.03fF
C211 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y a_33631_7375# 0.38fF
C212 freq_div_0/sky130_fd_sc_hd__inv_4_1/A freq_div_0/sky130_fd_sc_hd__inv_4_0/A 0.10fF
C213 freq_div_0/sky130_fd_sc_hd__inv_4_9/Y freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.42fF
C214 a_33716_6653# a_33631_6287# 0.11fF
C215 VDD freq_div_0/sky130_fd_sc_hd__inv_1_8/A 0.48fF
C216 a_34141_5743# a_34740_5743# 0.02fF
C217 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y a_34309_7643# 0.17fF
C218 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q freq_div_0/sky130_fd_sc_hd__inv_4_7/Y 0.42fF
C219 a_34309_7893# a_33884_7893# 0.04fF
C220 a_33614_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C221 freq_div_0/sky130_fd_sc_hd__inv_4_10/Y a_34141_5743# 0.14fF
C222 a_33716_7919# a_33884_7893# 0.59fF
C223 freq_div_0/sky130_fd_sc_hd__inv_4_9/A freq_div_0/sky130_fd_sc_hd__inv_4_8/A 0.09fF
C224 a_34309_6555# a_33277_6287# 0.11fF
C225 a_31443_6653# freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.14fF
C226 a_11158_1344# cs_ring_osc_0/vosc 0.25fF
C227 a_10140_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/vin 0.03fF
C228 a_33277_7375# a_33277_6837# 0.08fF
C229 VDD freq_div_0/sky130_fd_sc_hd__inv_1_3/A 0.48fF
C230 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_14071_n9035# 0.03fF
C231 a_14682_n2414# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C232 a_25242_1344# cs_ring_osc_0/cs_ring_osc_stage_5/csinvp 0.08fF
C233 a_34309_6805# a_33443_6837# 0.11fF
C234 a_33277_6837# a_33443_7375# 0.02fF
C235 VDD freq_div_0/vin 1.03fF
C236 a_31018_7919# a_30579_7375# 0.02fF
C237 cs_ring_osc_0/cs_ring_osc_stage_2/vin VDD 4.33fF
C238 a_15764_n11700# a_17138_n11700# 0.01fF
C239 a_30294_13935# pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N 0.14fF
C240 cs_ring_osc_0/cs_ring_osc_stage_2/vin cs_ring_osc_0/cs_ring_osc_stage_2/csinvp 0.10fF
C241 a_31235_14198# a_31040_14229# 0.49fF
C242 a_15156_6217# VDD 1.24fF
C243 cs_ring_osc_0/vpbias a_26158_1344# 0.63fF
C244 a_30579_7925# a_30745_7925# 2.23fF
C245 a_33842_7375# a_33716_7741# 0.02fF
C246 a_15306_n11700# a_16222_n11700# 1.92fF
C247 a_30745_6287# freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.61fF
C248 a_30745_6837# a_31186_6805# 0.28fF
C249 a_33631_7375# a_33631_6831# 0.02fF
C250 a_31611_6555# freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.17fF
C251 a_34141_6653# a_34267_6287# 0.04fF
C252 a_30579_5749# a_31186_5717# 0.37fF
C253 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_14530_n6542# 0.03fF
C254 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_31514_n2414# 0.03fF
C255 a_34740_6609# a_34309_6555# 0.31fF
C256 a_30745_6287# a_31443_6653# 0.44fF
C257 a_32042_6609# freq_div_0/sky130_fd_sc_hd__inv_4_4/A 0.05fF
C258 a_31611_6555# a_31443_6653# 0.67fF
C259 a_27803_13961# a_27287_13961# 0.42fF
C260 freq_div_0/sky130_fd_sc_hd__inv_4_8/Y freq_div_0/sky130_fd_sc_hd__inv_4_8/A 1.64fF
C261 a_16973_n921# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C262 a_31113_7741# a_31018_7741# 0.04fF
C263 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_34141_6831# 0.05fF
C264 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_29683_n921# 0.03fF
C265 vcp a_19988_n5874# 0.03fF
C266 VDD a_30579_7925# 0.79fF
C267 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y freq_div_0/sky130_fd_sc_hd__inv_1_7/A 0.27fF
C268 a_21362_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C269 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_33277_6287# 0.03fF
C270 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_14987_n9035# 0.03fF
C271 freq_div_0/sky130_fd_sc_hd__inv_1_4/A freq_div_0/sky130_fd_sc_hd__inv_1_2/A 0.04fF
C272 a_31611_6555# a_30745_6287# 0.11fF
C273 VDD a_33631_7375# 0.15fF
C274 freq_div_0/vout freq_div_0/sky130_fd_sc_hd__inv_1_6/A 0.07fF
C275 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y a_31443_5743# 0.14fF
C276 VDD a_31443_7741# 0.22fF
C277 cs_ring_osc_0/cs_ring_osc_stage_2/voutcs a_16973_n18921# 0.03fF
C278 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.38fF
C279 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_30579_6287# 0.03fF
C280 a_33631_5743# a_33716_5743# 0.11fF
C281 a_31113_5743# VDD 0.02fF
C282 VDD a_27125_7037# 0.01fF
C283 VDD a_34309_7643# 0.45fF
C284 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_34740_6609# 0.37fF
C285 a_33811_7741# a_33716_7741# 0.04fF
C286 a_30933_5743# a_31018_5743# 0.11fF
C287 VDD a_27074_n16656# 0.14fF
C288 cs_ring_osc_0/cs_ring_osc_stage_0/csinvp a_12074_1344# 0.10fF
C289 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q 0.38fF
C290 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y freq_div_0/sky130_fd_sc_hd__inv_4_3/Y 0.06fF
C291 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y a_33716_7741# 0.16fF
C292 a_32042_6831# freq_div_0/sky130_fd_sc_hd__inv_4_2/A 0.05fF
C293 VDD a_31113_6831# 0.02fF
C294 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.08fF
C295 a_30745_7925# a_30579_7375# 0.09fF
C296 a_27532_1344# a_27074_1344# 0.01fF
C297 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs VDD 4.44fF
C298 a_16222_n11700# a_16680_n11700# 0.01fF
C299 a_11158_1344# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.22fF
C300 a_31611_6805# freq_div_0/sky130_fd_sc_hd__inv_1_2/A 0.04fF
C301 vcp cs_ring_osc_0/cs_ring_osc_stage_3/csinvn 0.08fF
C302 a_30579_6837# a_30579_6287# 0.20fF
C303 freq_div_0/sky130_fd_sc_hd__inv_4_9/Y a_33443_6287# 0.61fF
C304 a_34141_6653# a_33884_6399# 0.11fF
C305 a_33277_6837# freq_div_0/sky130_fd_sc_hd__inv_4_2/Y 0.04fF
C306 vcp a_12430_n3082# 0.03fF
C307 cs_ring_osc_0/vpbias a_25700_n16656# 0.66fF
C308 freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.06fF
C309 a_34141_5743# a_34267_6121# 0.04fF
C310 VDD a_30579_7375# 0.79fF
C311 a_31443_7919# a_31569_8297# 0.04fF
C312 cs_ring_osc_0/vpbias a_16530_6217# 0.93fF
C313 cs_ring_osc_0/cs_ring_osc_stage_1/vin a_14390_n11700# 0.90fF
C314 VDD a_30391_13935# 0.37fF
C315 a_16988_9468# vcp 0.03fF
C316 a_30579_6837# freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.03fF
C317 a_34740_5743# freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.37fF
C318 a_30579_6837# freq_div_0/sky130_fd_sc_hd__inv_4_2/Y 0.35fF
C319 a_14682_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.03fF
C320 freq_div_0/sky130_fd_sc_hd__inv_1_10/A a_34309_5717# 0.04fF
C321 VDD a_27911_14327# 0.27fF
C322 a_34309_5717# a_34309_6555# 0.09fF
C323 a_32042_8785# freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q 0.37fF
C324 cs_ring_osc_0/cs_ring_osc_stage_5/vin a_26972_n2414# 0.03fF
C325 a_28021_14203# a_27911_14327# 0.23fF
C326 a_31798_14327# VDD 0.60fF
C327 a_15306_n11700# cs_ring_osc_0/vpbias 0.63fF
C328 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_30141_n921# 0.03fF
C329 a_30579_6837# a_31443_6831# 0.09fF
C330 pfd_cp_lpf_0/vRSTN pfd_cp_lpf_0/vQAb 0.29fF
C331 a_31079_14103# a_30391_13935# 0.12fF
C332 a_9682_n2414# cs_ring_osc_0/vosc 0.03fF
C333 freq_div_0/sky130_fd_sc_hd__inv_1_3/A freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q 0.07fF
C334 a_25242_1344# VDD 0.73fF
C335 freq_div_0/sky130_fd_sc_hd__inv_4_10/Y freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.42fF
C336 a_33716_6653# freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.16fF
C337 freq_div_0/sky130_fd_sc_hd__inv_4_7/A freq_div_0/sky130_fd_sc_hd__inv_4_8/A 0.10fF
C338 a_31798_14327# a_31079_14103# 0.23fF
C339 freq_div_0/vout a_34740_7919# 0.37fF
C340 freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q freq_div_0/sky130_fd_sc_hd__inv_4_4/A 0.02fF
C341 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_16362_n6542# 0.03fF
C342 VDD freq_div_0/sky130_fd_sc_hd__inv_1_7/A 0.48fF
C343 a_11158_1344# cs_ring_osc_0/vpbias 0.63fF
C344 freq_div_0/sky130_fd_sc_hd__inv_1_8/A freq_div_0/sky130_fd_sc_hd__inv_1_9/A 0.04fF
C345 VDD freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 0.91fF
C346 a_17431_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.03fF
C347 cs_ring_osc_0/cs_ring_osc_stage_5/vout a_24835_7037# 0.03fF
C348 freq_div_0/sky130_fd_sc_hd__inv_4_4/Y a_32042_6609# 0.11fF
C349 freq_div_0/sky130_fd_sc_hd__inv_4_8/Y a_33277_6837# 0.35fF
C350 freq_div_0/sky130_fd_sc_hd__inv_1_0/A VDD 0.48fF
C351 cs_ring_osc_0/vpbias a_12990_1344# 0.77fF
C352 a_30933_5743# a_30933_6287# 0.02fF
C353 a_31443_6653# a_32042_6609# 0.02fF
C354 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y a_31018_7919# 0.16fF
C355 a_34225_7741# a_34141_7741# 0.05fF
C356 pfd_cp_lpf_0/vpbias vcp 0.08fF
C357 a_27453_13961# a_28543_13935# 0.10fF
C358 a_31527_8829# a_31443_8829# 0.05fF
C359 a_30745_7375# freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 0.09fF
C360 cs_ring_osc_0/cs_ring_osc_stage_5/vout a_24834_9468# 0.03fF
C361 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_14988_n6542# 0.03fF
C362 a_30762_14213# a_30391_13935# 0.62fF
C363 cs_ring_osc_0/vpbias a_25242_n16656# 0.51fF
C364 a_33631_5743# a_33443_5749# 0.26fF
C365 a_30579_8463# a_31018_7919# 0.01fF
C366 a_24682_n21082# vcp 0.03fF
C367 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y a_30933_7375# 0.38fF
C368 a_31166_14327# a_30391_13935# 0.03fF
C369 VDD a_33716_7741# 0.36fF
C370 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_29682_n2414# 0.03fF
C371 a_33884_7487# a_33884_6805# 0.05fF
C372 a_31611_6555# a_32042_6609# 0.31fF
C373 cs_ring_osc_0/vpbias a_31680_n11700# 0.92fF
C374 a_30745_5749# a_31611_5717# 0.11fF
C375 a_12532_1344# a_12990_1344# 0.02fF
C376 a_18362_9468# vcp 0.03fF
C377 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.66fF
C378 a_15156_6217# a_14240_6217# 3.27fF
C379 a_30933_8463# freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.38fF
C380 a_31443_7741# freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q 0.05fF
C381 a_31144_6121# a_31018_5743# 0.02fF
C382 a_12431_n921# cs_ring_osc_0/vosc 0.03fF
C383 VDD a_33443_6287# 0.43fF
C384 cs_ring_osc_0/vpbias a_16680_n11700# 0.92fF
C385 freq_div_0/sky130_fd_sc_hd__inv_4_2/Y a_31186_6805# 0.15fF
C386 a_30764_n11700# a_31680_n11700# 1.33fF
C387 ibiasn pfd_cp_lpf_0/vswitchl 0.26fF
C388 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y freq_div_0/sky130_fd_sc_hd__inv_4_1/A 0.01fF
C389 a_31443_6831# a_31186_6805# 0.11fF
C390 a_24682_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C391 a_33884_6805# a_33716_6831# 0.59fF
C392 cs_ring_osc_0/cs_ring_osc_stage_1/csinvp a_14390_n11700# 0.08fF
C393 cs_ring_osc_0/vpbias a_15614_6217# 0.83fF
C394 a_27990_1344# cs_ring_osc_0/vpbias 0.77fF
C395 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y freq_div_0/sky130_fd_sc_hd__inv_4_4/A 0.03fF
C396 freq_div_0/sky130_fd_sc_hd__inv_1_6/A a_34740_7919# 0.25fF
C397 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_15904_n6542# 0.03fF
C398 a_34309_6805# a_34309_6555# 0.09fF
C399 a_30579_8463# a_30933_8463# 0.21fF
C400 vcp a_11056_n3082# 0.03fF
C401 a_28368_13961# a_27287_13961# 0.27fF
C402 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y freq_div_0/sky130_fd_sc_hd__inv_4_8/A 0.03fF
C403 freq_div_0/sky130_fd_sc_hd__inv_4_9/Y freq_div_0/sky130_fd_sc_hd__inv_4_8/A 0.01fF
C404 a_30306_n11700# a_31222_n11700# 1.92fF
C405 cs_ring_osc_0/cs_ring_osc_stage_3/vin a_27431_n18921# 0.03fF
C406 VDD a_33716_6653# 0.36fF
C407 pfd_cp_lpf_0/vRSTN a_29765_13961# 0.05fF
C408 a_26158_n16656# a_25242_n16656# 2.99fF
C409 a_33277_7375# freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q 0.03fF
C410 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y a_30745_7925# 0.61fF
C411 a_27430_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C412 a_33443_7375# freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q 0.03fF
C413 cs_ring_osc_0/cs_ring_osc_stage_1/vin cs_ring_osc_0/cs_ring_osc_stage_1/csinvn 0.09fF
C414 a_33631_5743# a_33277_5749# 0.21fF
C415 a_34740_7697# a_34141_7741# 0.02fF
C416 a_30579_7375# freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q 0.03fF
C417 vcp a_26514_n21082# 0.03fF
C418 VDD freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.96fF
C419 freq_div_0/sky130_fd_sc_hd__inv_1_6/A freq_div_0/sky130_fd_sc_hd__inv_4_6/A 0.35fF
C420 VDD a_31018_6831# 0.36fF
C421 a_30579_8463# a_30745_7925# 0.02fF
C422 a_33631_7919# a_33716_7919# 0.11fF
C423 freq_div_0/sky130_fd_sc_hd__inv_1_1/A freq_div_0/sky130_fd_sc_hd__inv_1_3/A 0.04fF
C424 a_34141_7919# a_33884_7893# 0.11fF
C425 freq_div_0/sky130_fd_sc_hd__inv_4_4/Y freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.04fF
C426 a_31113_8829# a_31018_8829# 0.04fF
C427 VDD cs_ring_osc_0/cs_ring_osc_stage_0/csinvp 0.48fF
C428 a_31018_6653# a_30579_5749# 0.01fF
C429 a_31018_6831# a_31144_7209# 0.02fF
C430 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y VDD 0.91fF
C431 a_33277_6287# a_33884_6399# 0.37fF
C432 vcp a_25140_n3082# 0.03fF
C433 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_34309_6805# 0.02fF
C434 a_34309_7893# freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q 0.02fF
C435 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y a_31018_7741# 0.16fF
C436 a_30579_8463# VDD 0.79fF
C437 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_33443_6837# 0.09fF
C438 a_31611_6805# a_30745_6837# 0.11fF
C439 freq_div_0/sky130_fd_sc_hd__inv_4_7/A a_34740_7697# 0.05fF
C440 pfd_cp_lpf_0/vpbias VDD 5.78fF
C441 a_31018_5743# a_30745_5749# 0.38fF
C442 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y freq_div_0/sky130_fd_sc_hd__inv_1_5/A 0.27fF
C443 VDD a_27532_1344# 0.09fF
C444 a_15764_n11700# a_16222_n11700# 0.02fF
C445 freq_div_0/sky130_fd_sc_hd__inv_1_0/A a_31611_8731# 0.04fF
C446 a_31443_8829# a_31569_8463# 0.04fF
C447 VDD pfd_cp_lpf_0/vQA 3.16fF
C448 a_33716_6653# a_33842_6287# 0.02fF
C449 a_26158_1344# a_27074_1344# 1.92fF
C450 a_32042_6831# a_32042_6609# 0.04fF
C451 VDD a_33811_6831# 0.02fF
C452 VDD freq_div_0/sky130_fd_sc_hd__inv_4_8/A 0.62fF
C453 a_19988_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C454 a_31186_8575# freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.15fF
C455 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_31515_n18921# 0.03fF
C456 a_33277_7375# a_33884_7487# 0.37fF
C457 a_34740_7919# freq_div_0/sky130_fd_sc_hd__inv_4_6/A 0.05fF
C458 a_32042_7697# a_31611_7643# 0.31fF
C459 a_33884_7487# a_33443_7375# 0.28fF
C460 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.13fF
C461 cs_ring_osc_0/vpbias a_31222_n11700# 0.76fF
C462 a_26972_n21082# vcp 0.03fF
C463 VDD a_32138_n11700# 0.06fF
C464 a_12074_n16656# a_12990_n16656# 0.79fF
C465 cs_ring_osc_0/cs_ring_osc_stage_2/vin a_11515_n18921# 0.03fF
C466 a_31222_n11700# cs_ring_osc_0/cs_ring_osc_stage_4/csinvp 0.10fF
C467 a_30745_7375# a_31186_7487# 0.28fF
C468 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_30598_n2414# 0.03fF
C469 a_11056_n21082# vcp 0.03fF
C470 a_31443_8829# a_30745_7925# 0.01fF
C471 cs_ring_osc_0/cs_ring_osc_stage_2/vin cs_ring_osc_0/cs_ring_osc_stage_2/csinvn 0.09fF
C472 a_31018_7741# a_31018_7919# 0.08fF
C473 a_31222_n11700# a_30764_n11700# 0.02fF
C474 a_31186_8575# a_30579_8463# 0.37fF
C475 a_33277_7375# a_33716_6831# 0.01fF
C476 pfd_cp_lpf_0/vQA a_30762_14213# 0.02fF
C477 pfd_cp_lpf_0/VQBb pfd_cp_lpf_0/vswitchl 0.28fF
C478 VDD a_30933_7375# 0.15fF
C479 a_27074_n16656# a_27532_n16656# 0.01fF
C480 a_34309_6805# a_33884_6805# 0.04fF
C481 a_36362_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C482 a_25242_n16656# cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.90fF
C483 a_32042_5743# a_31443_5743# 0.02fF
C484 a_12532_n16656# cs_ring_osc_0/vpbias 0.92fF
C485 a_15306_n11700# cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.25fF
C486 pfd_cp_lpf_0/vRSTN a_30391_13935# 0.70fF
C487 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y a_34740_7697# 0.11fF
C488 pfd_cp_lpf_0/vQA pfd_cp_lpf_0/vQB 0.15fF
C489 VDD a_31443_8829# 0.22fF
C490 pfd_cp_lpf_0/vRSTN a_27911_14327# 0.06fF
C491 a_33884_6805# a_33443_6837# 0.28fF
C492 VDD a_34225_7741# 0.02fF
C493 a_17138_n11700# a_16222_n11700# 0.79fF
C494 VDD a_14390_n11700# 0.73fF
C495 a_30579_5749# a_31611_5717# 0.11fF
C496 vcp cs_ring_osc_0/cs_ring_osc_stage_1/csinvn 0.08fF
C497 a_30933_8463# a_30745_8463# 0.26fF
C498 a_34141_5743# freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.05fF
C499 VDD a_27990_n16656# 0.06fF
C500 VDD a_33884_7893# 0.23fF
C501 cs_ring_osc_0/cs_ring_osc_stage_1/vin a_19529_n9035# 0.03fF
C502 cs_ring_osc_0/cs_ring_osc_stage_5/csinvp a_26158_1344# 0.09fF
C503 VDD freq_div_0/sky130_fd_sc_hd__inv_4_1/A 0.62fF
C504 a_34141_6831# a_33277_6837# 0.09fF
C505 a_33277_6837# a_33631_6831# 0.21fF
C506 a_34141_6831# a_34267_7209# 0.04fF
C507 a_32042_7697# freq_div_0/sky130_fd_sc_hd__inv_4_3/A 0.05fF
C508 a_30579_6287# a_30745_5749# 0.02fF
C509 a_31611_8731# freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.17fF
C510 a_27430_n21082# vcp 0.03fF
C511 a_12990_1344# a_11616_1344# 0.01fF
C512 a_15764_n11700# cs_ring_osc_0/vpbias 0.83fF
C513 VDD pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N 0.23fF
C514 freq_div_0/sky130_fd_sc_hd__inv_1_0/A freq_div_0/sky130_fd_sc_hd__inv_1_1/A 0.04fF
C515 a_29390_n11700# a_31222_n11700# 0.65fF
C516 a_30745_8463# a_30745_7925# 0.06fF
C517 a_14683_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.03fF
C518 a_24835_7037# VDD 0.01fF
C519 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q 0.38fF
C520 a_31611_5717# a_31186_5717# 0.04fF
C521 a_24683_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C522 a_15141_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.03fF
C523 VDD a_26616_n16656# 0.69fF
C524 a_28368_13961# a_27803_13961# 0.01fF
C525 a_33842_6121# a_33716_5743# 0.02fF
C526 a_34740_6609# freq_div_0/sky130_fd_sc_hd__inv_4_9/A 0.05fF
C527 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_15445_n9035# 0.03fF
C528 a_30579_8463# a_31611_8731# 0.11fF
C529 a_33884_6399# a_33884_5717# 0.05fF
C530 VDD a_33277_6837# 0.78fF
C531 freq_div_0/vout pfd_cp_lpf_0/VQBb 0.10fF
C532 a_33277_7375# a_33277_7925# 0.20fF
C533 a_16072_6217# a_16530_6217# 0.01fF
C534 VDD a_12074_n16656# 0.14fF
C535 VDD a_30745_8463# 0.43fF
C536 a_27287_13961# a_28543_13935# 0.12fF
C537 a_12074_n16656# cs_ring_osc_0/cs_ring_osc_stage_2/csinvp 0.10fF
C538 a_25141_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C539 a_33277_7925# a_33443_7375# 0.09fF
C540 cs_ring_osc_0/cs_ring_osc_stage_5/vin a_26973_n921# 0.03fF
C541 a_30579_6837# VDD 0.79fF
C542 a_31186_8575# a_31443_8829# 0.11fF
C543 VDD a_32042_5743# 0.37fF
C544 a_33631_5743# a_33884_5717# 0.04fF
C545 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_31515_n921# 0.03fF
C546 cs_ring_osc_0/vosc a_11057_n921# 0.03fF
C547 a_31380_14327# a_31040_14229# 0.12fF
C548 VDD a_14698_6217# 1.55fF
C549 a_27532_1344# a_26616_1344# 1.33fF
C550 cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_30445_n9035# 0.03fF
C551 freq_div_0/sky130_fd_sc_hd__inv_1_8/A freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q 0.07fF
C552 a_30745_7375# a_31611_7643# 0.11fF
C553 freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_34141_7741# 0.05fF
C554 VDD a_31018_7741# 0.36fF
C555 cs_ring_osc_0/vpbias cs_ring_osc_0/cs_ring_osc_stage_3/csinvp 0.31fF
C556 a_19987_n9035# cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C557 a_34141_6653# freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.14fF
C558 a_33277_6287# a_33631_6287# 0.21fF
C559 a_15306_n11700# cs_ring_osc_0/cs_ring_osc_stage_1/csinvp 0.09fF
C560 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.04fF
C561 VDD a_34225_5743# 0.02fF
C562 cs_ring_osc_0/cs_ring_osc_stage_5/vin cs_ring_osc_0/cs_ring_osc_stage_1/vin 1.49fF
C563 VDD pfd_cp_lpf_0/vpdiode 1.10fF
C564 vcp a_34988_n5874# 0.03fF
C565 cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_16056_n2414# 0.03fF
C566 a_11158_1344# a_12074_1344# 1.92fF
C567 VDD a_34740_7697# 0.37fF
C568 a_31611_6805# freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.39fF
C569 a_31443_7741# a_31569_7375# 0.04fF
C570 a_31611_6805# freq_div_0/sky130_fd_sc_hd__inv_4_2/Y 0.17fF
C571 freq_div_0/sky130_fd_sc_hd__inv_4_6/Y a_33884_7893# 0.15fF
C572 a_33277_7925# a_34309_7893# 0.11fF
C573 a_17430_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.03fF
C574 a_12074_1344# a_12990_1344# 0.79fF
C575 a_33277_7925# a_33716_7919# 0.63fF
C576 a_31611_6805# a_31443_6831# 0.67fF
C577 cs_ring_osc_0/vpbias a_17138_n11700# 0.77fF
C578 a_31018_5743# a_30579_5749# 0.63fF
C579 a_32042_5743# freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.45fF
C580 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 0.30fF
C581 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_34309_6555# 0.39fF
C582 a_26515_n921# cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.03fF
C583 freq_div_0/sky130_fd_sc_hd__inv_4_8/Y a_33716_6831# 0.16fF
C584 cs_ring_osc_0/cs_ring_osc_stage_4/csinvn cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.09fF
C585 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_30599_n18921# 0.03fF
C586 a_32042_7697# a_32042_7919# 0.04fF
C587 a_33443_7925# a_33884_7893# 0.28fF
C588 a_27990_1344# a_27074_1344# 0.79fF
C589 VDD a_33716_5743# 0.36fF
C590 freq_div_0/sky130_fd_sc_hd__inv_1_8/A freq_div_0/sky130_fd_sc_hd__inv_1_7/A 0.04fF
C591 a_31186_8575# a_30745_8463# 0.28fF
C592 a_34141_6653# a_34141_6831# 0.05fF
C593 a_33277_7375# a_33443_6837# 0.02fF
C594 VDD vsigin 0.12fF
C595 a_34141_5743# a_33443_6287# 0.01fF
C596 VDD a_26158_1344# 0.40fF
C597 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y freq_div_0/sky130_fd_sc_hd__inv_1_1/A 0.27fF
C598 a_33443_7375# a_33443_6837# 0.06fF
C599 a_31186_6399# a_31186_6805# 0.03fF
C600 pfd_cp_lpf_0/VQBb pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N 0.08fF
C601 a_31018_5743# a_31186_5717# 0.59fF
C602 a_31611_8731# a_31443_8829# 0.67fF
C603 cs_ring_osc_0/vpbias a_16988_6217# 0.85fF
C604 a_26158_n16656# cs_ring_osc_0/cs_ring_osc_stage_3/csinvp 0.09fF
C605 VDD a_31186_6805# 0.23fF
C606 a_31079_14103# vsigin 0.51fF
C607 VDD a_30933_5743# 0.15fF
C608 a_31611_7893# a_31018_7919# 0.02fF
C609 a_15614_6217# a_16072_6217# 0.02fF
C610 freq_div_0/vout a_34309_7893# 0.38fF
C611 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_33631_7375# 0.02fF
C612 a_17904_9468# vcp 0.03fF
C613 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_14072_n6542# 0.03fF
C614 a_33884_7487# a_34141_7741# 0.11fF
C615 cs_ring_osc_0/cs_ring_osc_stage_0/csinvp a_10242_1344# 0.08fF
C616 pfd_cp_lpf_0/vRSTN a_30797_13961# 0.01fF
C617 a_32042_8785# a_32042_7919# 0.04fF
C618 cs_ring_osc_0/cs_ring_osc_stage_5/vout cs_ring_osc_0/cs_ring_osc_stage_5/voutcs 0.38fF
C619 a_30579_7925# a_30579_7375# 0.20fF
C620 a_10242_n16656# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.82fF
C621 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_34309_7643# 0.02fF
C622 VDD a_34225_6653# 0.02fF
C623 pfd_cp_lpf_0/vRSTN pfd_cp_lpf_0/vQA 1.34fF
C624 VDD a_34141_6653# 0.22fF
C625 vcp cs_ring_osc_0/cs_ring_osc_stage_5/csinvn 0.08fF
C626 VDD a_31527_7741# 0.02fF
C627 freq_div_0/sky130_fd_sc_hd__inv_4_8/Y a_34740_6831# 0.11fF
C628 vcp cs_ring_osc_0/cs_ring_osc_stage_4/csinvn 0.08fF
C629 pfd_cp_lpf_0/vQA pfd_cp_lpf_0/vQAb 3.28fF
C630 a_31443_7741# a_30579_7375# 0.09fF
C631 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_16361_n9035# 0.03fF
C632 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q 0.29fF
C633 freq_div_0/sky130_fd_sc_hd__inv_4_10/Y a_33716_5743# 0.16fF
C634 VDD a_27453_13961# 1.24fF
C635 a_30579_6837# freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q 0.49fF
C636 a_28021_14203# a_27453_13961# 0.41fF
C637 a_27990_1344# cs_ring_osc_0/cs_ring_osc_stage_5/csinvp 0.16fF
C638 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_32431_n921# 0.03fF
C639 a_31611_8731# a_30745_8463# 0.11fF
C640 a_31443_7919# a_31018_7919# 0.03fF
C641 a_29071_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs 0.03fF
C642 a_31018_6653# a_31144_6287# 0.02fF
C643 vcp a_11972_n21082# 0.03fF
C644 a_30579_6287# a_30579_5749# 0.08fF
C645 cs_ring_osc_0/cs_ring_osc_stage_5/vin a_25140_n2414# 0.03fF
C646 cs_ring_osc_0/cs_ring_osc_stage_5/vin vcp 6.63fF
C647 cs_ring_osc_0/cs_ring_osc_stage_5/csinvp cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.10fF
C648 a_32042_5743# freq_div_0/sky130_fd_sc_hd__inv_1_5/A 0.25fF
C649 cs_ring_osc_0/cs_ring_osc_stage_3/vin a_26514_n20414# 0.03fF
C650 a_33443_5749# VDD 0.43fF
C651 a_11158_n16656# a_10242_n16656# 2.99fF
C652 cs_ring_osc_0/vpbias a_10242_n16656# 0.51fF
C653 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.42fF
C654 cs_ring_osc_0/cs_ring_osc_stage_2/vin a_9682_n20414# 0.03fF
C655 freq_div_0/sky130_fd_sc_hd__inv_1_7/A a_34309_7643# 0.04fF
C656 a_31611_7893# a_30745_7925# 0.11fF
C657 a_31527_6831# a_31443_6831# 0.05fF
C658 VDD a_25700_n16656# 1.55fF
C659 freq_div_0/sky130_fd_sc_hd__inv_1_6/A a_34309_7893# 0.04fF
C660 VDD a_16530_6217# 0.09fF
C661 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_31443_6653# 0.05fF
C662 a_30933_6831# a_30745_6837# 0.26fF
C663 a_33277_6287# freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.35fF
C664 cs_ring_osc_0/cs_ring_osc_stage_2/vin a_12431_n18921# 0.03fF
C665 a_16680_n11700# a_14848_n11700# 0.43fF
C666 vcp a_10598_n21082# 0.03fF
C667 a_15306_n11700# VDD 0.40fF
C668 a_31113_7919# a_31018_7919# 0.04fF
C669 a_33842_7209# a_33716_6831# 0.02fF
C670 a_33631_7375# a_33716_7741# 0.11fF
C671 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_30745_6287# 0.03fF
C672 VDD a_31040_14229# 1.23fF
C673 VDD a_31611_7893# 0.45fF
C674 a_27803_13961# a_28543_13935# 0.02fF
C675 a_20904_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C676 a_31611_6555# freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q 0.39fF
C677 a_11158_1344# VDD 0.40fF
C678 a_33443_5749# freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.06fF
C679 freq_div_0/sky130_fd_sc_hd__inv_1_1/A freq_div_0/sky130_fd_sc_hd__inv_4_1/A 0.35fF
C680 VDD a_33631_7919# 0.15fF
C681 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q a_30745_7925# 0.03fF
C682 freq_div_0/vin freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.05fF
C683 a_34740_6609# freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.11fF
C684 a_33716_7741# a_34309_7643# 0.02fF
C685 a_31079_14103# a_31040_14229# 1.60fF
C686 VDD a_12990_1344# 0.06fF
C687 cs_ring_osc_0/cs_ring_osc_stage_3/vin cs_ring_osc_0/cs_ring_osc_stage_3/csinvp 0.10fF
C688 a_34309_6805# freq_div_0/sky130_fd_sc_hd__inv_4_8/Y 0.17fF
C689 a_31443_5743# a_30745_5749# 0.44fF
C690 freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q a_33443_6287# 0.08fF
C691 pfd_cp_lpf_0/vRSTN pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N 0.09fF
C692 a_33884_7487# freq_div_0/sky130_fd_sc_hd__inv_4_7/Y 0.15fF
C693 freq_div_0/sky130_fd_sc_hd__inv_4_10/A freq_div_0/sky130_fd_sc_hd__inv_1_10/A 0.35fF
C694 a_33443_5749# freq_div_0/sky130_fd_sc_hd__inv_4_10/Y 0.61fF
C695 freq_div_0/sky130_fd_sc_hd__inv_4_8/Y a_33443_6837# 0.61fF
C696 a_27990_n16656# a_27532_n16656# 0.02fF
C697 VDD a_25242_n16656# 0.73fF
C698 a_31443_7919# a_30745_7925# 0.44fF
C699 a_30579_6837# a_30745_6287# 0.09fF
C700 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q 2.23fF
C701 pfd_cp_lpf_0/vQAb pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N 0.08fF
C702 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y a_31186_7487# 0.15fF
C703 a_30579_8463# freq_div_0/vin 0.41fF
C704 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 2.18fF
C705 a_34267_7375# a_34141_7741# 0.04fF
C706 VDD a_33277_5749# 0.78fF
C707 cs_ring_osc_0/vosc cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.40fF
C708 VDD a_31680_n11700# 0.09fF
C709 a_30762_14213# a_31040_14229# 0.29fF
C710 freq_div_0/sky130_fd_sc_hd__inv_1_8/A freq_div_0/sky130_fd_sc_hd__inv_4_8/A 0.35fF
C711 a_16057_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.03fF
C712 a_34740_7919# a_34309_7893# 0.31fF
C713 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_30745_7925# 0.08fF
C714 cs_ring_osc_0/cs_ring_osc_stage_5/vout a_25293_7037# 0.03fF
C715 a_16515_n921# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C716 a_31443_7919# VDD 0.22fF
C717 a_27532_n16656# a_26616_n16656# 1.33fF
C718 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y a_30579_7925# 0.35fF
C719 VDD a_16680_n11700# 0.09fF
C720 a_31166_14327# a_31040_14229# 0.41fF
C721 a_31018_6653# a_31113_6653# 0.04fF
C722 freq_div_0/sky130_fd_sc_hd__inv_4_2/Y freq_div_0/sky130_fd_sc_hd__inv_4_3/A 0.03fF
C723 a_30579_8463# a_30579_7925# 0.08fF
C724 cs_ring_osc_0/cs_ring_osc_stage_1/vin a_19530_n6542# 0.03fF
C725 VDD a_33277_6287# 0.78fF
C726 cs_ring_osc_0/cs_ring_osc_stage_2/vin a_10599_n18921# 0.03fF
C727 VDD a_15614_6217# 0.69fF
C728 a_27990_1344# VDD 0.06fF
C729 a_34309_6555# a_33884_6399# 0.04fF
C730 a_31186_7893# a_31018_7919# 0.59fF
C731 a_11616_n16656# a_12074_n16656# 0.02fF
C732 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_31057_n921# 0.03fF
C733 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q 0.38fF
C734 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_29683_n18921# 0.03fF
C735 VDD a_27708_13961# 0.60fF
C736 a_33277_5749# freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.41fF
C737 a_26972_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C738 a_31018_6831# a_31113_6831# 0.04fF
C739 a_33631_7919# freq_div_0/sky130_fd_sc_hd__inv_4_6/Y 0.38fF
C740 vcp pfd_cp_lpf_0/vswitchl 0.07fF
C741 VDD cs_ring_osc_0/cs_ring_osc_stage_5/vin 4.26fF
C742 cs_ring_osc_0/vosc cs_ring_osc_0/vpbias 2.76fF
C743 a_33443_6837# a_34141_7741# 0.01fF
C744 a_31113_7919# VDD 0.02fF
C745 a_19072_n5874# vcp 0.03fF
C746 a_34141_7919# a_33277_7925# 0.09fF
C747 a_34141_6831# a_33716_6831# 0.03fF
C748 VDD a_30745_5749# 0.43fF
C749 a_33716_6831# a_33631_6831# 0.11fF
C750 VDD a_34740_6609# 0.37fF
C751 freq_div_0/sky130_fd_sc_hd__inv_4_10/Y a_33277_5749# 0.35fF
C752 a_30933_6831# a_30933_6287# 0.02fF
C753 VDD freq_div_0/sky130_fd_sc_hd__inv_1_4/A 0.48fF
C754 a_25598_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C755 freq_div_0/sky130_fd_sc_hd__inv_4_6/Y freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q 0.30fF
C756 VDD a_33884_7487# 0.23fF
C757 a_31018_6831# a_30579_7375# 0.01fF
C758 a_31018_6653# a_31018_5743# 0.05fF
C759 a_29848_n11700# a_31680_n11700# 0.43fF
C760 cs_ring_osc_0/cs_ring_osc_stage_1/vin a_20445_n9035# 0.03fF
C761 a_33631_7919# a_33443_7925# 0.26fF
C762 a_12532_n16656# a_12990_n16656# 0.02fF
C763 VDD a_31113_8829# 0.02fF
C764 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_32042_6609# 0.37fF
C765 a_30306_n11700# cs_ring_osc_0/vpbias 0.63fF
C766 cs_ring_osc_0/vpbias a_16222_n11700# 0.76fF
C767 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_14529_n9035# 0.03fF
C768 a_16515_n18921# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.03fF
C769 a_30306_n11700# cs_ring_osc_0/cs_ring_osc_stage_4/csinvp 0.09fF
C770 a_34225_5743# a_34141_5743# 0.05fF
C771 VDD a_33716_6831# 0.36fF
C772 a_30745_5749# freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.01fF
C773 a_31611_8731# a_31611_7893# 0.09fF
C774 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y a_31611_7643# 0.17fF
C775 a_33443_7925# freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q 0.09fF
C776 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_31056_n2414# 0.03fF
C777 cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_31362_n6542# 0.03fF
C778 a_30933_6831# freq_div_0/sky130_fd_sc_hd__inv_4_2/Y 0.38fF
C779 a_31186_7893# a_30745_7925# 0.28fF
C780 VDD a_31611_6805# 0.45fF
C781 a_18820_9468# vcp 0.03fF
C782 freq_div_0/sky130_fd_sc_hd__inv_1_0/A freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.27fF
C783 cs_ring_osc_0/cs_ring_osc_stage_5/vout a_25292_9468# 0.03fF
C784 a_34740_6609# a_34740_5743# 0.04fF
C785 a_32042_5743# a_32042_6609# 0.04fF
C786 freq_div_0/vout a_34141_7919# 0.04fF
C787 a_30391_13935# a_30797_13961# 0.04fF
C788 a_34141_6831# a_34740_6831# 0.02fF
C789 cs_ring_osc_0/cs_ring_osc_stage_2/vin a_11972_n20414# 0.03fF
C790 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q 0.08fF
C791 pfd_cp_lpf_0/vQA a_30391_13935# 0.39fF
C792 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.40fF
C793 a_16072_9468# vcp 0.03fF
C794 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs VDD 4.44fF
C795 cs_ring_osc_0/cs_ring_osc_stage_1/csinvp a_17138_n11700# 0.16fF
C796 a_31186_7893# VDD 0.23fF
C797 a_33716_6653# a_33443_6287# 0.38fF
C798 a_31235_14198# a_31545_13961# 0.07fF
C799 a_11158_n16656# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.22fF
C800 freq_div_0/sky130_fd_sc_hd__inv_1_4/A freq_div_0/sky130_fd_sc_hd__inv_4_4/A 0.35fF
C801 a_33716_5743# a_34141_5743# 0.03fF
C802 cs_ring_osc_0/vosc a_11514_n2414# 0.03fF
C803 a_28368_13961# a_28543_13935# 0.62fF
C804 a_15764_n11700# a_14848_n11700# 2.26fF
C805 a_25599_n921# cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.03fF
C806 pfd_cp_lpf_0/vRSTN a_27453_13961# 0.33fF
C807 VDD a_31222_n11700# 0.14fF
C808 cs_ring_osc_0/cs_ring_osc_stage_5/vin cs_ring_osc_0/cs_ring_osc_stage_4/voutcs 0.38fF
C809 a_30745_8463# freq_div_0/vin 0.06fF
C810 a_31018_6653# a_30933_6287# 0.11fF
C811 VDD a_34309_5717# 0.45fF
C812 cs_ring_osc_0/cs_ring_osc_stage_1/vin a_19072_n6542# 0.03fF
C813 a_12532_n16656# a_10700_n16656# 0.43fF
C814 a_16988_6217# a_16072_6217# 0.79fF
C815 a_15446_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/voutcs 0.03fF
C816 a_29390_n11700# a_30306_n11700# 2.99fF
C817 VDD a_34740_6831# 0.37fF
C818 a_30579_5749# a_31443_5743# 0.09fF
C819 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y freq_div_0/sky130_fd_sc_hd__inv_4_3/A 1.64fF
C820 VDD a_31186_7487# 0.23fF
C821 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q freq_div_0/sky130_fd_sc_hd__inv_1_2/A 0.07fF
C822 freq_div_0/sky130_fd_sc_hd__inv_1_2/A freq_div_0/sky130_fd_sc_hd__inv_4_2/Y 0.27fF
C823 a_33884_6805# a_33884_6399# 0.03fF
C824 VDD a_27287_13961# 0.90fF
C825 a_27074_n16656# a_27990_n16656# 0.79fF
C826 a_28021_14203# a_27287_13961# 0.16fF
C827 a_30933_7375# a_30579_7375# 0.21fF
C828 cs_ring_osc_0/cs_ring_osc_stage_5/vout a_27582_9468# 0.03fF
C829 a_30745_7375# a_30745_6837# 0.06fF
C830 a_35445_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C831 a_25140_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C832 a_31018_6653# a_30579_6287# 0.63fF
C833 a_12532_n16656# VDD 0.09fF
C834 a_32042_8785# freq_div_0/sky130_fd_sc_hd__inv_4_0/A 0.05fF
C835 VDD a_33277_7925# 0.78fF
C836 a_27990_1344# a_26616_1344# 0.01fF
C837 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_31611_8731# 0.39fF
C838 a_30745_8463# a_30579_7925# 0.02fF
C839 a_34141_6653# a_34141_5743# 0.07fF
C840 cs_ring_osc_0/vpbias a_11158_n16656# 0.63fF
C841 a_31018_5743# a_31611_5717# 0.02fF
C842 VDD a_33884_5717# 0.23fF
C843 a_36362_n5874# vcp 0.03fF
C844 cs_ring_osc_0/vpbias cs_ring_osc_0/cs_ring_osc_stage_4/csinvp 0.31fF
C845 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q freq_div_0/sky130_fd_sc_hd__inv_4_2/Y 0.02fF
C846 pfd_cp_lpf_0/vRSTN a_31040_14229# 0.33fF
C847 a_34309_5717# a_34740_5743# 0.31fF
C848 a_31443_5743# a_31186_5717# 0.11fF
C849 a_27532_n16656# a_25700_n16656# 0.43fF
C850 a_30933_7919# a_31018_7919# 0.11fF
C851 a_27074_n16656# a_26616_n16656# 0.02fF
C852 a_30579_7925# a_31018_7741# 0.02fF
C853 a_31186_7893# a_31186_8575# 0.05fF
C854 a_34309_6805# a_34141_6831# 0.67fF
C855 freq_div_0/sky130_fd_sc_hd__inv_1_1/A a_31611_7893# 0.04fF
C856 cs_ring_osc_0/vpbias a_30764_n11700# 0.83fF
C857 pfd_cp_lpf_0/vndiode pfd_cp_lpf_0/vswitchh 0.15fF
C858 cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_31361_n9035# 0.03fF
C859 freq_div_0/sky130_fd_sc_hd__inv_1_4/A freq_div_0/sky130_fd_sc_hd__inv_1_5/A 0.04fF
C860 a_33277_6287# freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.04fF
C861 a_34309_5717# freq_div_0/sky130_fd_sc_hd__inv_4_10/Y 0.17fF
C862 a_34141_6831# a_33443_6837# 0.44fF
C863 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.13fF
C864 a_33631_6831# a_33443_6837# 0.26fF
C865 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_33277_6837# 0.03fF
C866 a_15764_n11700# VDD 0.69fF
C867 a_34740_6609# freq_div_0/sky130_fd_sc_hd__inv_1_9/A 0.25fF
C868 a_31443_7741# a_31018_7741# 0.03fF
C869 cs_ring_osc_0/cs_ring_osc_stage_5/vout a_26667_7037# 0.03fF
C870 cs_ring_osc_0/cs_ring_osc_stage_5/vout a_25750_9468# 0.03fF
C871 cs_ring_osc_0/vpbias a_12532_1344# 0.92fF
C872 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_32430_n2414# 0.03fF
C873 a_33443_5749# a_34141_5743# 0.44fF
C874 a_30579_8463# freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.35fF
C875 a_31611_6805# freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q 0.02fF
C876 pfd_cp_lpf_0/vQB pfd_cp_lpf_0/vswitchl 0.44fF
C877 a_11158_1344# a_10242_1344# 2.99fF
C878 freq_div_0/sky130_fd_sc_hd__inv_1_1/A freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 0.07fF
C879 VDD a_31527_6831# 0.02fF
C880 freq_div_0/vout VDD 0.55fF
C881 VDD a_30579_5749# 0.79fF
C882 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q freq_div_0/sky130_fd_sc_hd__inv_4_8/Y 0.30fF
C883 a_34740_7697# a_34309_7643# 0.31fF
C884 VDD a_34309_6805# 0.45fF
C885 a_12990_1344# a_10242_1344# 0.14fF
C886 a_16972_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.03fF
C887 a_31443_6653# a_30745_5749# 0.01fF
C888 a_26057_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C889 freq_div_0/sky130_fd_sc_hd__inv_1_4/A freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.27fF
C890 a_30933_7919# a_30933_8463# 0.02fF
C891 freq_div_0/sky130_fd_sc_hd__inv_4_7/A freq_div_0/sky130_fd_sc_hd__inv_4_6/A 0.09fF
C892 freq_div_0/sky130_fd_sc_hd__inv_4_10/Y a_33884_5717# 0.15fF
C893 VDD a_33443_6837# 0.43fF
C894 a_34529_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C895 a_26158_n16656# cs_ring_osc_0/vpbias 0.63fF
C896 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 0.42fF
C897 a_33277_7925# freq_div_0/sky130_fd_sc_hd__inv_4_6/Y 0.35fF
C898 a_30579_6837# a_30579_7375# 0.08fF
C899 a_27431_n921# cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.03fF
C900 a_34141_7919# a_34740_7919# 0.02fF
C901 a_29390_n11700# cs_ring_osc_0/vpbias 0.51fF
C902 VDD a_25293_7037# 0.01fF
C903 VDD cs_ring_osc_0/cs_ring_osc_stage_3/csinvp 0.48fF
C904 a_31018_7741# a_30579_7375# 0.63fF
C905 a_30745_6287# a_30745_5749# 0.06fF
C906 a_29390_n11700# cs_ring_osc_0/cs_ring_osc_stage_4/csinvp 0.08fF
C907 cs_ring_osc_0/cs_ring_osc_stage_5/vout a_25751_7037# 0.03fF
C908 a_26056_n21082# vcp 0.03fF
C909 vcp a_18614_n5874# 0.03fF
C910 VDD a_31611_7643# 0.45fF
C911 a_31186_6399# a_31186_5717# 0.05fF
C912 cs_ring_osc_0/cs_ring_osc_stage_2/vin a_10598_n20414# 0.03fF
C913 cs_ring_osc_0/cs_ring_osc_stage_5/vout cs_ring_osc_0/vosc 1.76fF
C914 a_30933_7919# a_30745_7925# 0.26fF
C915 VDD a_31186_5717# 0.23fF
C916 a_31611_6555# freq_div_0/sky130_fd_sc_hd__inv_1_4/A 0.04fF
C917 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y a_32042_5743# 0.11fF
C918 VDD a_17138_n11700# 0.06fF
C919 VDD a_33811_5743# 0.02fF
C920 cs_ring_osc_0/vpbias a_25700_1344# 0.66fF
C921 a_33277_7925# a_33443_7925# 2.23fF
C922 a_33277_5749# a_34141_5743# 0.09fF
C923 freq_div_0/sky130_fd_sc_hd__inv_1_7/A a_34740_7697# 0.25fF
C924 a_17431_n921# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C925 a_30933_7919# VDD 0.15fF
C926 freq_div_0/vout pfd_cp_lpf_0/vQB 0.12fF
C927 a_16972_n2414# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C928 a_12990_n16656# a_10242_n16656# 0.14fF
C929 a_33277_6837# a_33716_7741# 0.01fF
C930 VDD freq_div_0/sky130_fd_sc_hd__inv_1_6/A 0.48fF
C931 a_31443_8829# freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.14fF
C932 VDD a_31527_7919# 0.02fF
C933 a_31569_6287# a_31443_6653# 0.04fF
C934 a_31443_7741# a_31527_7741# 0.05fF
C935 a_32430_n20414# cs_ring_osc_0/cs_ring_osc_stage_3/voutcs 0.03fF
C936 freq_div_0/vout freq_div_0/sky130_fd_sc_hd__inv_4_6/Y 0.10fF
C937 a_33277_7375# a_33443_7375# 2.23fF
C938 a_31611_6555# a_31611_6805# 0.09fF
C939 VDD a_16988_6217# 0.06fF
C940 a_33884_6805# freq_div_0/sky130_fd_sc_hd__inv_4_8/Y 0.15fF
C941 cs_ring_osc_0/cs_ring_osc_stage_3/vin cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.38fF
C942 a_33277_6837# a_33443_6287# 0.09fF
C943 cs_ring_osc_0/vosc cs_ring_osc_0/vosc2 0.27fF
C944 VDD pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N 0.23fF
C945 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y freq_div_0/sky130_fd_sc_hd__inv_4_6/A 0.01fF
C946 vcp a_10598_n3082# 0.03fF
C947 cs_ring_osc_0/cs_ring_osc_stage_2/vin a_10141_n18921# 0.03fF
C948 freq_div_0/sky130_fd_sc_hd__inv_4_1/A freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.03fF
C949 a_31798_14327# vsigin 0.01fF
C950 a_30745_6837# a_30579_6287# 0.09fF
C951 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_31973_n921# 0.03fF
C952 VDD freq_div_0/sky130_fd_sc_hd__inv_4_3/A 0.62fF
C953 a_29107_13961# pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N 0.14fF
C954 a_30579_8463# a_31443_8829# 0.09fF
C955 a_21361_n9035# cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C956 a_25242_1344# a_26158_1344# 2.99fF
C957 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y freq_div_0/sky130_fd_sc_hd__inv_4_1/A 1.66fF
C958 a_30745_6837# freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.03fF
C959 a_30745_6837# freq_div_0/sky130_fd_sc_hd__inv_4_2/Y 0.61fF
C960 a_30745_7375# a_31443_6831# 0.01fF
C961 cs_ring_osc_0/cs_ring_osc_stage_2/vin a_11056_n20414# 0.03fF
C962 vcp a_34072_n5874# 0.03fF
C963 freq_div_0/vout a_33443_7925# 0.01fF
C964 a_33716_6653# a_33277_6837# 0.02fF
C965 a_31443_6831# a_30745_6837# 0.44fF
C966 freq_div_0/sky130_fd_sc_hd__inv_4_10/A freq_div_0/sky130_fd_sc_hd__inv_4_9/A 0.10fF
C967 a_33277_7375# a_33716_7919# 0.02fF
C968 a_33443_5749# freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.03fF
C969 VDD a_27803_13961# 0.33fF
C970 a_15598_n2414# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C971 a_32042_7697# freq_div_0/sky130_fd_sc_hd__inv_4_3/Y 0.11fF
C972 vcp a_12430_n21082# 0.03fF
C973 a_28021_14203# a_27803_13961# 0.50fF
C974 a_30933_5743# freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 0.38fF
C975 a_31380_14327# a_31235_14198# 0.21fF
C976 cs_ring_osc_0/cs_ring_osc_stage_1/vin cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.38fF
C977 a_34309_6555# freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.17fF
C978 cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_16057_n921# 0.03fF
C979 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs VDD 4.44fF
C980 a_30579_7925# a_31611_7893# 0.11fF
C981 a_30306_n11700# cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.25fF
C982 a_30745_8463# freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.61fF
C983 a_30579_6837# a_31018_6831# 0.63fF
C984 VDD a_34740_7919# 0.37fF
C985 a_30579_6287# a_31018_5743# 0.01fF
C986 cs_ring_osc_0/vosc a_9683_n921# 0.03fF
C987 a_27911_14327# a_27453_13961# 0.12fF
C988 a_34309_7893# a_33716_7919# 0.02fF
C989 pfd_cp_lpf_0/vQB pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N 0.13fF
C990 freq_div_0/sky130_fd_sc_hd__inv_1_6/A freq_div_0/sky130_fd_sc_hd__inv_4_6/Y 0.27fF
C991 a_33631_7919# a_33631_7375# 0.02fF
C992 a_31018_6831# a_31018_7741# 0.05fF
C993 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_13613_n9035# 0.03fF
C994 a_31611_7643# freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q 0.39fF
C995 cs_ring_osc_0/vosc vcp 5.08fF
C996 freq_div_0/sky130_fd_sc_hd__inv_1_4/A a_32042_6609# 0.25fF
C997 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_13614_n6542# 0.03fF
C998 pfd_cp_lpf_0/vQA pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N 0.13fF
C999 VDD a_10242_n16656# 0.73fF
C1000 cs_ring_osc_0/cs_ring_osc_stage_1/csinvp a_16222_n11700# 0.10fF
C1001 a_30579_8463# a_30745_8463# 2.23fF
C1002 pfd_cp_lpf_0/vRSTN a_27287_13961# 0.86fF
C1003 cs_ring_osc_0/cs_ring_osc_stage_2/csinvp a_10242_n16656# 0.08fF
C1004 a_30579_7925# freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 0.03fF
C1005 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q freq_div_0/vin 0.04fF
C1006 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.29fF
C1007 a_30933_6831# VDD 0.15fF
C1008 VDD freq_div_0/sky130_fd_sc_hd__inv_4_6/A 0.62fF
C1009 cs_ring_osc_0/cs_ring_osc_stage_5/vin a_26057_n921# 0.03fF
C1010 cs_ring_osc_0/vpbias a_11616_1344# 0.83fF
C1011 a_31443_7919# a_30579_7925# 0.09fF
C1012 a_33716_6653# a_33716_5743# 0.05fF
C1013 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_30598_n20414# 0.03fF
C1014 a_25242_n16656# a_27074_n16656# 0.65fF
C1015 a_33277_5749# freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.03fF
C1016 freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_34309_7643# 0.39fF
C1017 VDD a_32042_7919# 0.37fF
C1018 a_12532_n16656# a_11616_n16656# 1.33fF
C1019 a_26158_n16656# cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.25fF
C1020 a_30391_13935# a_31040_14229# 0.10fF
C1021 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_25242_n16656# 0.82fF
C1022 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q 0.08fF
C1023 a_34141_6653# a_33443_6287# 0.44fF
C1024 a_31611_6805# a_32042_6831# 0.31fF
C1025 a_31443_7919# a_31443_7741# 0.05fF
C1026 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_30579_7925# 0.49fF
C1027 freq_div_0/sky130_fd_sc_hd__inv_4_2/A freq_div_0/sky130_fd_sc_hd__inv_4_3/A 0.10fF
C1028 a_30745_6287# a_30579_5749# 0.02fF
C1029 a_34309_5717# a_34141_5743# 0.67fF
C1030 a_31798_14327# a_31040_14229# 0.22fF
C1031 VDD a_34309_6555# 0.45fF
C1032 a_12532_1344# a_11616_1344# 1.33fF
C1033 vcp pfd_cp_lpf_0/vswitchh 0.15fF
C1034 freq_div_0/sky130_fd_sc_hd__inv_1_10/A VDD 0.48fF
C1035 a_30579_6287# a_30933_6287# 0.21fF
C1036 a_31018_6831# a_31186_6805# 0.59fF
C1037 a_26973_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C1038 vcp a_9682_n21082# 0.03fF
C1039 cs_ring_osc_0/vpbias a_27074_1344# 0.76fF
C1040 vcp a_17446_9468# 0.03fF
C1041 a_33277_6287# freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.49fF
C1042 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_33631_6831# 0.02fF
C1043 a_34740_7919# freq_div_0/sky130_fd_sc_hd__inv_4_6/Y 0.11fF
C1044 a_33716_6653# a_34141_6653# 0.03fF
C1045 a_33884_6399# a_33631_6287# 0.04fF
C1046 VDD a_26667_7037# 0.01fF
C1047 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q a_30579_7375# 0.51fF
C1048 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q a_30933_6287# 0.02fF
C1049 VDD freq_div_0/sky130_fd_sc_hd__inv_1_2/A 0.48fF
C1050 a_30745_7375# freq_div_0/sky130_fd_sc_hd__inv_4_3/Y 0.61fF
C1051 a_33443_5749# a_33443_6287# 0.06fF
C1052 a_33631_5743# a_33631_6287# 0.02fF
C1053 cs_ring_osc_0/cs_ring_osc_stage_4/csinvp cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.10fF
C1054 cs_ring_osc_0/cs_ring_osc_stage_2/vin a_12430_n20414# 0.03fF
C1055 a_34141_5743# a_33884_5717# 0.11fF
C1056 a_16988_6217# a_14240_6217# 0.14fF
C1057 a_27990_n16656# a_26616_n16656# 0.01fF
C1058 cs_ring_osc_0/vpbias a_12074_1344# 0.76fF
C1059 cs_ring_osc_0/vpbias a_16072_6217# 0.77fF
C1060 cs_ring_osc_0/cs_ring_osc_stage_5/vin a_24682_n2414# 0.03fF
C1061 a_31144_8297# a_31018_7919# 0.02fF
C1062 a_31443_8829# a_30745_8463# 0.44fF
C1063 freq_div_0/sky130_fd_sc_hd__inv_1_7/A freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q 0.07fF
C1064 a_31018_6653# a_31186_6399# 0.59fF
C1065 a_30933_7375# a_31018_7741# 0.11fF
C1066 freq_div_0/sky130_fd_sc_hd__inv_4_6/A freq_div_0/sky130_fd_sc_hd__inv_4_6/Y 1.64fF
C1067 a_31018_6653# VDD 0.36fF
C1068 a_30579_6287# freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.51fF
C1069 a_33884_7487# a_33631_7375# 0.04fF
C1070 cs_ring_osc_0/cs_ring_osc_stage_1/csinvp cs_ring_osc_0/vpbias 0.31fF
C1071 a_33277_5749# freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 0.04fF
C1072 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q 2.23fF
C1073 freq_div_0/sky130_fd_sc_hd__inv_1_8/A a_34740_6831# 0.25fF
C1074 freq_div_0/sky130_fd_sc_hd__inv_1_10/A a_34740_5743# 0.25fF
C1075 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q freq_div_0/sky130_fd_sc_hd__inv_4_2/Y 0.29fF
C1076 a_33884_7487# a_34309_7643# 0.04fF
C1077 VDD a_25751_7037# 0.01fF
C1078 freq_div_0/sky130_fd_sc_hd__inv_1_10/A freq_div_0/sky130_fd_sc_hd__inv_4_10/Y 0.27fF
C1079 a_33277_7375# a_34141_7741# 0.09fF
C1080 cs_ring_osc_0/vosc VDD 8.63fF
C1081 cs_ring_osc_0/cs_ring_osc_stage_5/vin a_26514_n2414# 0.03fF
C1082 a_12074_1344# a_12532_1344# 0.01fF
C1083 a_31443_6831# freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.05fF
C1084 a_31443_6831# freq_div_0/sky130_fd_sc_hd__inv_4_2/Y 0.14fF
C1085 a_27911_14327# a_27708_13961# 0.02fF
C1086 a_33443_7375# a_34141_7741# 0.44fF
C1087 a_27990_1344# a_25242_1344# 0.14fF
C1088 VDD a_28368_13961# 0.39fF
C1089 cs_ring_osc_0/cs_ring_osc_stage_1/vin a_18613_n9035# 0.03fF
C1090 a_31443_5743# a_31611_5717# 0.67fF
C1091 a_32042_7697# VDD 0.37fF
C1092 cs_ring_osc_0/vosc a_10141_n921# 0.03fF
C1093 a_34987_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C1094 a_28368_13961# a_28021_14203# 0.13fF
C1095 cs_ring_osc_0/vpbias vcp 13.40fF
C1096 cs_ring_osc_0/vpbias cs_ring_osc_0/cs_ring_osc_stage_5/csinvp 0.31fF
C1097 a_25242_1344# cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.90fF
C1098 cs_ring_osc_0/cs_ring_osc_stage_2/vin a_11973_n18921# 0.03fF
C1099 a_33613_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C1100 a_30933_6831# freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q 0.02fF
C1101 vcp a_27430_n3082# 0.03fF
C1102 VDD a_31235_14198# 0.33fF
C1103 a_31186_7893# a_30579_7925# 0.37fF
C1104 cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_29072_n6542# 0.03fF
C1105 a_33884_6805# a_33631_6831# 0.04fF
C1106 freq_div_0/sky130_fd_sc_hd__inv_1_0/A freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q 0.07fF
C1107 a_33884_6805# a_34141_6831# 0.11fF
C1108 a_29390_n11700# cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.90fF
C1109 a_31018_7919# a_31018_8829# 0.05fF
C1110 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y a_33277_7375# 0.04fF
C1111 VDD a_30306_n11700# 0.40fF
C1112 a_31079_14103# a_31235_14198# 0.42fF
C1113 a_33277_5749# a_33443_6287# 0.02fF
C1114 VDD a_16222_n11700# 0.14fF
C1115 freq_div_0/sky130_fd_sc_hd__inv_4_9/A freq_div_0/sky130_fd_sc_hd__inv_4_8/Y 0.01fF
C1116 cs_ring_osc_0/vosc a_11972_n2414# 0.03fF
C1117 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y a_30745_5749# 0.61fF
C1118 pfd_cp_lpf_0/vRSTN pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N 0.08fF
C1119 a_16514_n2414# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C1120 a_12990_n16656# a_11158_n16656# 0.24fF
C1121 freq_div_0/sky130_fd_sc_hd__inv_4_10/A freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.03fF
C1122 cs_ring_osc_0/vpbias a_12990_n16656# 0.77fF
C1123 a_32042_8785# VDD 0.37fF
C1124 a_10140_n2414# cs_ring_osc_0/vosc 0.03fF
C1125 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_29682_n20414# 0.03fF
C1126 a_30579_6837# a_31018_7741# 0.01fF
C1127 a_25599_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C1128 a_11158_1344# cs_ring_osc_0/cs_ring_osc_stage_0/csinvp 0.09fF
C1129 VDD pfd_cp_lpf_0/vswitchh 10.21fF
C1130 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y a_31611_7893# 0.17fF
C1131 a_34309_5717# freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.39fF
C1132 a_33716_6653# a_33277_5749# 0.01fF
C1133 cs_ring_osc_0/vpbias a_14848_n11700# 0.66fF
C1134 VDD a_33884_6805# 0.23fF
C1135 freq_div_0/sky130_fd_sc_hd__inv_1_2/A freq_div_0/sky130_fd_sc_hd__inv_4_2/A 0.35fF
C1136 a_33277_6287# a_33443_6287# 2.23fF
C1137 a_34530_n5874# vcp 0.03fF
C1138 cs_ring_osc_0/cs_ring_osc_stage_0/csinvp a_12990_1344# 0.16fF
C1139 a_34309_6805# freq_div_0/sky130_fd_sc_hd__inv_1_8/A 0.04fF
C1140 a_31443_7741# a_31186_7487# 0.11fF
C1141 a_31235_14198# a_30762_14213# 0.01fF
C1142 pfd_cp_lpf_0/vRSTN a_27803_13961# 0.30fF
C1143 a_31443_5743# a_31569_6121# 0.04fF
C1144 a_28368_13961# pfd_cp_lpf_0/vQB 0.02fF
C1145 VDD freq_div_0/sky130_fd_sc_hd__inv_4_5/A 0.62fF
C1146 a_30933_8463# a_31018_8829# 0.11fF
C1147 a_34141_6831# a_34225_6831# 0.05fF
C1148 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_34740_6831# 0.37fF
C1149 a_31235_14198# a_31166_14327# 0.50fF
C1150 VDD a_31611_5717# 0.45fF
C1151 freq_div_0/sky130_fd_sc_hd__inv_1_10/A freq_div_0/sky130_fd_sc_hd__inv_1_9/A 0.04fF
C1152 a_34309_6555# freq_div_0/sky130_fd_sc_hd__inv_1_9/A 0.04fF
C1153 VDD cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 4.44fF
C1154 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q 0.02fF
C1155 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 0.29fF
C1156 a_33884_7487# a_33716_7741# 0.59fF
C1157 VDD cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 4.44fF
C1158 a_33716_6653# a_33277_6287# 0.63fF
C1159 a_33884_6399# freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.15fF
C1160 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q freq_div_0/sky130_fd_sc_hd__inv_4_2/A 0.02fF
C1161 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_30933_5743# 0.02fF
C1162 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_25242_1344# 0.82fF
C1163 a_30745_7375# a_30745_7925# 0.05fF
C1164 a_31443_7919# freq_div_0/sky130_fd_sc_hd__inv_4_1/Y 0.14fF
C1165 a_31018_5743# a_31443_5743# 0.03fF
C1166 a_33277_7375# freq_div_0/sky130_fd_sc_hd__inv_4_7/Y 0.35fF
C1167 a_34141_7919# a_34309_7893# 0.67fF
C1168 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y a_33443_7375# 0.61fF
C1169 freq_div_0/sky130_fd_sc_hd__inv_1_3/A a_31611_7643# 0.04fF
C1170 a_31186_7487# a_30579_7375# 0.37fF
C1171 a_34141_7919# a_33716_7919# 0.03fF
C1172 cs_ring_osc_0/vpbias a_10700_n16656# 0.66fF
C1173 a_33716_6831# a_33716_7741# 0.05fF
C1174 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.42fF
C1175 freq_div_0/sky130_fd_sc_hd__inv_4_5/A freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.14fF
C1176 a_30579_6837# a_31186_6805# 0.37fF
C1177 VDD a_34225_6831# 0.02fF
C1178 a_30745_7375# VDD 0.43fF
C1179 a_31611_5717# freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.38fF
C1180 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q 0.42fF
C1181 VDD a_30745_6837# 0.43fF
C1182 VDD a_31113_6653# 0.02fF
C1183 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y freq_div_0/sky130_fd_sc_hd__inv_4_2/Y 0.13fF
C1184 VDD a_31018_8829# 0.36fF
C1185 a_32042_7697# freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q 0.37fF
C1186 VDD a_11158_n16656# 0.40fF
C1187 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q freq_div_0/sky130_fd_sc_hd__inv_1_9/A 0.07fF
C1188 VDD pfd_cp_lpf_0/VQBb 0.42fF
C1189 VDD cs_ring_osc_0/vpbias 18.73fF
C1190 freq_div_0/sky130_fd_sc_hd__inv_4_10/A VDD 0.62fF
C1191 a_30306_n11700# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs 0.22fF
C1192 cs_ring_osc_0/cs_ring_osc_stage_2/csinvp a_11158_n16656# 0.09fF
C1193 cs_ring_osc_0/vpbias cs_ring_osc_0/cs_ring_osc_stage_2/csinvp 0.31fF
C1194 a_30579_8463# freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q 0.03fF
C1195 VDD cs_ring_osc_0/cs_ring_osc_stage_4/csinvp 0.48fF
C1196 freq_div_0/sky130_fd_sc_hd__inv_4_5/A freq_div_0/sky130_fd_sc_hd__inv_4_4/A 0.10fF
C1197 a_15599_n921# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C1198 a_31443_6831# a_31569_7209# 0.04fF
C1199 pfd_cp_lpf_0/VQBb a_29107_13961# 0.04fF
C1200 cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_30446_n6542# 0.03fF
C1201 VDD a_30764_n11700# 0.69fF
C1202 a_31018_6653# freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.16fF
C1203 freq_div_0/sky130_fd_sc_hd__inv_1_1/A a_32042_7919# 0.25fF
C1204 a_15306_n11700# a_14390_n11700# 2.99fF
C1205 a_27990_1344# a_27532_1344# 0.02fF
C1206 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_31514_n20414# 0.03fF
C1207 a_33716_6653# a_33716_6831# 0.08fF
C1208 a_34309_6805# a_34309_7643# 0.09fF
C1209 a_31018_6653# a_31443_6653# 0.03fF
C1210 a_31680_n11700# a_32138_n11700# 0.02fF
C1211 a_34309_6805# freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q 0.39fF
C1212 a_34141_6831# a_33443_7375# 0.01fF
C1213 VDD a_12532_1344# 0.09fF
C1214 a_33631_7919# a_33884_7893# 0.04fF
C1215 a_16514_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.03fF
C1216 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_33443_6837# 0.03fF
C1217 freq_div_0/sky130_fd_sc_hd__inv_4_7/A freq_div_0/sky130_fd_sc_hd__inv_4_8/Y 0.03fF
C1218 a_31443_7741# a_31611_7643# 0.67fF
C1219 freq_div_0/sky130_fd_sc_hd__inv_1_3/A freq_div_0/sky130_fd_sc_hd__inv_4_3/A 0.35fF
C1220 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q a_30933_7375# 0.02fF
C1221 a_25700_n16656# a_26616_n16656# 2.26fF
C1222 a_34530_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C1223 a_27074_n16656# cs_ring_osc_0/cs_ring_osc_stage_3/csinvp 0.10fF
C1224 a_31018_6653# a_30745_6287# 0.38fF
C1225 freq_div_0/sky130_fd_sc_hd__inv_4_10/A a_34740_5743# 0.05fF
C1226 VDD a_31018_5743# 0.36fF
C1227 cs_ring_osc_0/vosc a_11056_n2414# 0.03fF
C1228 VDD a_33884_6399# 0.23fF
C1229 a_32042_8785# a_31611_8731# 0.31fF
C1230 a_15156_6217# a_16988_6217# 0.24fF
C1231 a_31018_6653# a_31611_6555# 0.02fF
C1232 vcp a_10140_n3082# 0.03fF
C1233 a_31611_6805# a_31018_6831# 0.02fF
C1234 cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_28613_n9035# 0.03fF
C1235 a_30933_7919# a_30579_7925# 0.21fF
C1236 a_31037_13961# a_30762_14213# 0.04fF
C1237 a_33277_7925# a_33716_7741# 0.02fF
C1238 a_25242_n16656# a_27990_n16656# 0.14fF
C1239 vcp cs_ring_osc_0/cs_ring_osc_stage_3/vin 4.16fF
C1240 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_31973_n18921# 0.03fF
C1241 a_31186_8575# a_31018_8829# 0.59fF
C1242 VDD a_33277_7375# 0.78fF
C1243 a_26158_n16656# VDD 0.40fF
C1244 freq_div_0/sky130_fd_sc_hd__inv_4_10/A freq_div_0/sky130_fd_sc_hd__inv_4_10/Y 1.64fF
C1245 a_33631_5743# VDD 0.15fF
C1246 a_12074_1344# a_11616_1344# 0.02fF
C1247 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_15903_n9035# 0.03fF
C1248 cs_ring_osc_0/cs_ring_osc_stage_1/csinvp cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.10fF
C1249 pfd_cp_lpf_0/VQBb pfd_cp_lpf_0/vQB 1.54fF
C1250 freq_div_0/sky130_fd_sc_hd__inv_4_1/A freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q 0.02fF
C1251 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_31972_n20414# 0.03fF
C1252 a_14698_6217# a_16530_6217# 0.43fF
C1253 VDD a_33443_7375# 0.43fF
C1254 cs_ring_osc_0/vpbias a_29848_n11700# 0.66fF
C1255 a_31443_7919# a_31443_8829# 0.07fF
C1256 a_29390_n11700# VDD 0.73fF
C1257 freq_div_0/sky130_fd_sc_hd__inv_4_9/A freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 1.66fF
C1258 VDD a_31113_7741# 0.02fF
C1259 vcp a_20446_n5874# 0.03fF
C1260 VDD freq_div_0/sky130_fd_sc_hd__inv_4_0/A 0.62fF
C1261 VDD a_28543_13935# 0.37fF
C1262 a_28021_14203# a_28543_13935# 0.03fF
C1263 freq_div_0/sky130_fd_sc_hd__inv_1_5/A freq_div_0/sky130_fd_sc_hd__inv_4_5/A 0.35fF
C1264 a_30579_5749# freq_div_0/sky130_fd_sc_hd__inv_4_5/Y 0.35fF
C1265 a_29848_n11700# a_30764_n11700# 2.26fF
C1266 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs cs_ring_osc_0/cs_ring_osc_stage_2/vin 0.38fF
C1267 a_31611_7643# a_30579_7375# 0.11fF
C1268 freq_div_0/sky130_fd_sc_hd__inv_1_5/A a_31611_5717# 0.04fF
C1269 a_31186_7893# freq_div_0/sky130_fd_sc_hd__inv_4_1/Y 0.15fF
C1270 pfd_cp_lpf_0/vndiode VDD 0.32fF
C1271 a_29107_13961# a_28543_13935# 0.30fF
C1272 vcp a_11514_n3082# 0.03fF
C1273 VDD a_25700_1344# 1.55fF
C1274 VDD a_30294_13935# 0.29fF
C1275 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_31443_8829# 0.05fF
C1276 VDD a_34309_7893# 0.45fF
C1277 cs_ring_osc_0/cs_ring_osc_stage_1/vin vcp 4.28fF
C1278 VDD a_33716_7919# 0.36fF
C1279 a_33811_6831# a_33716_6831# 0.04fF
C1280 a_33631_5743# freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.02fF
C1281 pfd_cp_lpf_0/vRSTN a_28368_13961# 0.56fF
C1282 a_28368_13961# a_28530_14327# 0.04fF
C1283 a_33443_5749# a_33716_5743# 0.38fF
C1284 a_34225_6653# a_34141_6653# 0.05fF
C1285 a_30745_7375# freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q 0.03fF
C1286 a_30933_6287# a_31186_6399# 0.04fF
C1287 freq_div_0/sky130_fd_sc_hd__inv_4_8/Y freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.06fF
C1288 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y freq_div_0/sky130_fd_sc_hd__inv_4_8/Y 0.13fF
C1289 freq_div_0/sky130_fd_sc_hd__inv_4_4/Y freq_div_0/sky130_fd_sc_hd__inv_4_5/A 0.03fF
C1290 cs_ring_osc_0/cs_ring_osc_stage_2/vin a_10242_n16656# 0.90fF
C1291 cs_ring_osc_0/cs_ring_osc_stage_5/vin a_26056_n2414# 0.03fF
C1292 a_30745_6837# freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q 0.08fF
C1293 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y a_31186_5717# 0.15fF
C1294 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q freq_div_0/sky130_fd_sc_hd__inv_4_3/A 0.02fF
C1295 VDD a_30933_6287# 0.15fF
C1296 VDD a_33811_6653# 0.02fF
C1297 pfd_cp_lpf_0/vRSTN a_31235_14198# 0.30fF
C1298 a_33631_5743# freq_div_0/sky130_fd_sc_hd__inv_4_10/Y 0.38fF
C1299 cs_ring_osc_0/vosc a_10242_1344# 2.75fF
C1300 cs_ring_osc_0/vpbias a_10700_1344# 0.66fF
C1301 a_31611_8731# a_31018_8829# 0.02fF
C1302 cs_ring_osc_0/cs_ring_osc_stage_5/vin a_25598_n2414# 0.03fF
C1303 a_31443_7919# a_30745_8463# 0.01fF
C1304 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y a_33277_7925# 0.04fF
C1305 freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q a_34740_7697# 0.37fF
C1306 a_28722_13961# a_28543_13935# 0.04fF
C1307 a_33631_6287# freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.38fF
C1308 cs_ring_osc_0/vpbias a_26616_1344# 0.83fF
C1309 a_30579_6287# a_31186_6399# 0.37fF
C1310 a_33884_7487# a_33884_7893# 0.03fF
C1311 pfd_cp_lpf_0/vQB a_28543_13935# 0.39fF
C1312 a_34141_7919# a_34141_7741# 0.05fF
C1313 freq_div_0/sky130_fd_sc_hd__inv_1_2/A a_32042_6831# 0.25fF
C1314 VDD a_30579_6287# 0.79fF
C1315 a_33277_6287# a_33277_6837# 0.20fF
C1316 a_33443_6837# a_33443_6287# 0.05fF
C1317 freq_div_0/sky130_fd_sc_hd__inv_1_6/A freq_div_0/sky130_fd_sc_hd__inv_1_7/A 0.04fF
C1318 cs_ring_osc_0/cs_ring_osc_stage_5/csinvp a_27074_1344# 0.10fF
C1319 a_31040_14229# vsigin 0.04fF
C1320 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_30745_8463# 0.03fF
C1321 a_33443_5749# a_34141_6653# 0.01fF
C1322 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_30745_5749# 0.08fF
C1323 vcp a_33614_n5874# 0.03fF
C1324 a_31611_6555# a_31611_5717# 0.09fF
C1325 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q 2.18fF
C1326 VDD freq_div_0/sky130_fd_sc_hd__inv_4_2/Y 0.91fF
C1327 cs_ring_osc_0/vpbias a_14240_6217# 0.60fF
C1328 a_14698_6217# a_15614_6217# 2.26fF
C1329 vcp cs_ring_osc_0/cs_ring_osc_stage_4/vin 3.55fF
C1330 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_30140_n2414# 0.03fF
C1331 a_12532_1344# a_10700_1344# 0.43fF
C1332 a_34740_6831# freq_div_0/sky130_fd_sc_hd__inv_4_8/A 0.05fF
C1333 a_34141_6831# freq_div_0/sky130_fd_sc_hd__inv_4_8/Y 0.14fF
C1334 VDD freq_div_0/sky130_fd_sc_hd__inv_4_9/A 0.62fF
C1335 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q freq_div_0/sky130_fd_sc_hd__inv_1_4/A 0.07fF
C1336 freq_div_0/sky130_fd_sc_hd__inv_4_8/Y a_33631_6831# 0.38fF
C1337 vcp a_16530_9468# 0.03fF
C1338 pfd_cp_lpf_0/vQAb pfd_cp_lpf_0/vswitchh 1.92fF
C1339 VDD a_31443_6831# 0.22fF
C1340 a_31222_n11700# a_32138_n11700# 0.79fF
C1341 a_29390_n11700# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs 0.82fF
C1342 a_34141_7919# a_34225_7919# 0.05fF
C1343 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_30140_n20414# 0.03fF
C1344 a_33277_7375# a_33443_7925# 0.09fF
C1345 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y a_34141_7741# 0.14fF
C1346 a_34309_7893# freq_div_0/sky130_fd_sc_hd__inv_4_6/Y 0.17fF
C1347 vcp a_26056_n3082# 0.03fF
C1348 a_27911_14327# a_27803_13961# 0.21fF
C1349 freq_div_0/sky130_fd_sc_hd__inv_4_6/Y a_33716_7919# 0.16fF
C1350 freq_div_0/sky130_fd_sc_hd__inv_1_3/A freq_div_0/sky130_fd_sc_hd__inv_1_2/A 0.04fF
C1351 a_33443_7925# a_33443_7375# 0.05fF
C1352 VDD cs_ring_osc_0/cs_ring_osc_stage_3/vin 4.26fF
C1353 a_33277_5749# a_33716_5743# 0.63fF
C1354 a_33631_6287# a_33631_6831# 0.02fF
C1355 vcp a_9682_n3082# 0.03fF
C1356 a_30745_6287# a_30745_6837# 0.05fF
C1357 a_32042_7697# a_32042_6831# 0.04fF
C1358 VDD freq_div_0/sky130_fd_sc_hd__inv_4_8/Y 0.93fF
C1359 cs_ring_osc_0/vosc cs_ring_osc_0/cs_ring_osc_stage_0/csinvn 0.09fF
C1360 a_30933_7375# a_31186_7487# 0.04fF
C1361 a_34309_7893# a_33443_7925# 0.11fF
C1362 freq_div_0/sky130_fd_sc_hd__inv_4_7/A freq_div_0/sky130_fd_sc_hd__inv_4_7/Y 1.64fF
C1363 a_33716_6831# a_33277_6837# 0.63fF
C1364 a_33443_7925# a_33716_7919# 0.38fF
C1365 a_24683_n921# cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.03fF
C1366 a_33277_6287# a_33716_5743# 0.01fF
C1367 cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_10242_1344# 0.82fF
C1368 cs_ring_osc_0/cs_ring_osc_stage_5/vout VDD 9.13fF
C1369 VDD cs_ring_osc_0/cs_ring_osc_stage_1/vin 4.26fF
C1370 a_34309_6555# freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.02fF
C1371 a_34141_6831# a_34141_7741# 0.07fF
C1372 freq_div_0/sky130_fd_sc_hd__inv_4_10/Y freq_div_0/sky130_fd_sc_hd__inv_4_9/A 0.03fF
C1373 a_27990_1344# a_26158_1344# 0.24fF
C1374 freq_div_0/sky130_fd_sc_hd__inv_1_10/A freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.07fF
C1375 VDD a_33631_6287# 0.15fF
C1376 freq_div_0/sky130_fd_sc_hd__inv_4_2/Y freq_div_0/sky130_fd_sc_hd__inv_4_4/A 0.01fF
C1377 VDD a_11616_1344# 0.69fF
C1378 pfd_cp_lpf_0/vRSTN pfd_cp_lpf_0/VQBb 0.20fF
C1379 a_30579_6837# a_31611_6805# 0.11fF
C1380 a_32042_7697# freq_div_0/sky130_fd_sc_hd__inv_1_3/A 0.25fF
C1381 cs_ring_osc_0/cs_ring_osc_stage_5/vin a_26158_1344# 0.25fF
C1382 a_25700_1344# a_26616_1344# 2.26fF
C1383 a_33277_7925# a_33884_7893# 0.37fF
C1384 a_29530_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs 0.03fF
C1385 a_30933_7919# freq_div_0/sky130_fd_sc_hd__inv_4_1/Y 0.38fF
C1386 a_28368_13961# a_28477_13961# 0.04fF
C1387 cs_ring_osc_0/vpbias a_11616_n16656# 0.83fF
C1388 cs_ring_osc_0/vpbias a_27532_n16656# 0.92fF
C1389 a_34141_6653# a_33277_6287# 0.09fF
C1390 cs_ring_osc_0/cs_ring_osc_stage_5/vout freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.21fF
C1391 VDD a_34141_7741# 0.22fF
C1392 a_30933_5743# a_30745_5749# 0.26fF
C1393 cs_ring_osc_0/vpbias a_10242_1344# 0.51fF
C1394 a_35904_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C1395 a_15140_n2414# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C1396 a_31527_8829# VDD 0.02fF
C1397 a_33443_5749# a_33277_5749# 2.23fF
C1398 VDD cs_ring_osc_0/vosc2 0.58fF
C1399 VDD a_27074_1344# 0.14fF
C1400 freq_div_0/sky130_fd_sc_hd__inv_4_2/Y freq_div_0/sky130_fd_sc_hd__inv_4_2/A 1.64fF
C1401 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q 0.07fF
C1402 cs_ring_osc_0/cs_ring_osc_stage_0/voutcs a_15141_n921# 0.03fF
C1403 vcp a_26514_n3082# 0.03fF
C1404 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q 0.08fF
C1405 freq_div_0/sky130_fd_sc_hd__inv_4_2/Y freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q 0.42fF
C1406 VDD cs_ring_osc_0/cs_ring_osc_stage_4/vin 4.91fF
C1407 a_15140_n20414# cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.03fF
C1408 cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_30903_n9035# 0.03fF
C1409 a_11158_1344# a_12990_1344# 0.24fF
C1410 a_12532_n16656# a_12074_n16656# 0.01fF
C1411 a_27708_13961# a_27453_13961# 0.22fF
C1412 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y freq_div_0/sky130_fd_sc_hd__inv_4_3/A 0.01fF
C1413 a_31380_14327# VDD 0.27fF
C1414 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q 0.08fF
C1415 a_34740_6609# a_34141_6653# 0.02fF
C1416 a_11514_n21082# vcp 0.03fF
C1417 VDD a_34225_7919# 0.02fF
C1418 cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_29529_n9035# 0.03fF
C1419 a_30933_6287# freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.38fF
C1420 a_31186_7487# a_31018_7741# 0.59fF
C1421 VDD freq_div_0/sky130_fd_sc_hd__inv_4_3/Y 0.91fF
C1422 a_32042_7697# a_31443_7741# 0.02fF
C1423 VDD a_12074_1344# 0.14fF
C1424 VDD a_16072_6217# 0.52fF
C1425 a_34740_6831# a_34740_7697# 0.04fF
C1426 a_33443_5749# a_33277_6287# 0.02fF
C1427 VDD freq_div_0/sky130_fd_sc_hd__inv_4_7/A 0.62fF
C1428 a_33631_7919# freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q 0.02fF
C1429 vcp a_24682_n3082# 0.03fF
C1430 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q a_31611_7893# 0.39fF
C1431 pfd_cp_lpf_0/vpdiode pfd_cp_lpf_0/vswitchl 0.08fF
C1432 VDD cs_ring_osc_0/cs_ring_osc_stage_1/csinvp 0.48fF
C1433 a_31611_6805# a_31186_6805# 0.04fF
C1434 cs_ring_osc_0/cs_ring_osc_stage_3/vin a_26056_n20414# 0.03fF
C1435 pfd_cp_lpf_0/vRSTN a_28543_13935# 0.70fF
C1436 a_27899_13961# a_27803_13961# 0.07fF
C1437 a_31527_5743# a_31443_5743# 0.05fF
C1438 a_25141_n921# cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.03fF
C1439 freq_div_0/sky130_fd_sc_hd__inv_1_9/A freq_div_0/sky130_fd_sc_hd__inv_4_9/A 0.35fF
C1440 a_15614_6217# a_16530_6217# 1.33fF
C1441 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs a_26158_1344# 0.22fF
C1442 a_31443_7919# a_31611_7893# 0.67fF
C1443 cs_ring_osc_0/vosc a_12430_n2414# 0.03fF
C1444 a_30579_6287# freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.35fF
C1445 cs_ring_osc_0/cs_ring_osc_stage_2/vin cs_ring_osc_0/cs_ring_osc_stage_2/voutcs 0.40fF
C1446 a_30745_6287# a_30933_6287# 0.26fF
C1447 pfd_cp_lpf_0/vRSTN a_30294_13935# 0.10fF
C1448 a_30579_6287# a_31443_6653# 0.09fF
C1449 a_27990_n16656# cs_ring_osc_0/cs_ring_osc_stage_3/csinvp 0.16fF
C1450 a_34309_5717# a_33716_5743# 0.02fF
C1451 a_31380_14327# a_30762_14213# 0.01fF
C1452 a_18614_n6542# cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C1453 a_10140_n21082# vcp 0.03fF
C1454 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.30fF
C1455 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q a_30579_5749# 0.49fF
C1456 freq_div_0/sky130_fd_sc_hd__inv_4_2/Y freq_div_0/sky130_fd_sc_hd__inv_4_4/Y 0.06fF
C1457 a_30745_7925# a_31018_7919# 0.38fF
C1458 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q a_31611_7893# 0.02fF
C1459 a_30933_7919# a_30933_7375# 0.02fF
C1460 pfd_cp_lpf_0/vQAb a_30294_13935# 0.04fF
C1461 VDD vcp 5.04fF
C1462 VDD cs_ring_osc_0/cs_ring_osc_stage_5/csinvp 0.48fF
C1463 vcp a_20904_n5874# 0.03fF
C1464 VDD a_34141_7919# 0.22fF
C1465 a_17138_n11700# a_14390_n11700# 0.14fF
C1466 a_34309_6555# a_33443_6287# 0.11fF
C1467 a_31380_14327# a_31166_14327# 0.23fF
C1468 a_28368_13961# a_27911_14327# 0.01fF
C1469 a_31443_6831# a_31443_6653# 0.05fF
C1470 a_31443_7919# freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 0.05fF
C1471 a_30745_6287# a_30579_6287# 2.23fF
C1472 a_34309_6805# a_33277_6837# 0.11fF
C1473 a_30933_6831# a_31018_6831# 0.11fF
C1474 a_31611_6555# a_30579_6287# 0.11fF
C1475 cs_ring_osc_0/cs_ring_osc_stage_4/voutcs a_28614_n6542# 0.03fF
C1476 a_31235_14198# a_30391_13935# 0.02fF
C1477 a_35446_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C1478 a_10700_1344# a_11616_1344# 2.26fF
C1479 a_31186_7487# a_31186_6805# 0.05fF
C1480 a_33277_6837# a_33443_6837# 2.23fF
C1481 VDD a_31018_7919# 0.36fF
C1482 a_31144_7375# a_31018_7741# 0.02fF
C1483 a_31798_14327# a_31235_14198# 0.13fF
C1484 a_30745_6287# freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.09fF
C1485 a_31611_6555# freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q 0.02fF
C1486 cs_ring_osc_0/cs_ring_osc_stage_2/vin a_11158_n16656# 0.25fF
C1487 VDD a_33811_7741# 0.02fF
C1488 a_33716_5743# a_33884_5717# 0.59fF
C1489 a_17430_n2414# cs_ring_osc_0/cs_ring_osc_stage_0/voutcs 0.03fF
C1490 VDD a_12990_n16656# 0.06fF
C1491 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q 0.07fF
C1492 VDD freq_div_0/sky130_fd_sc_hd__inv_4_7/Y 0.93fF
C1493 a_33716_6653# a_34309_6555# 0.02fF
C1494 VDD freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.93fF
C1495 a_33277_6287# a_33277_5749# 0.08fF
C1496 cs_ring_osc_0/cs_ring_osc_stage_5/vin a_27430_n2414# 0.03fF
C1497 freq_div_0/sky130_fd_sc_hd__inv_4_7/A freq_div_0/sky130_fd_sc_hd__inv_4_6/Y 0.01fF
C1498 cs_ring_osc_0/cs_ring_osc_stage_2/csinvp a_12990_n16656# 0.16fF
C1499 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_31056_n20414# 0.03fF
C1500 a_15156_6217# cs_ring_osc_0/vpbias 0.73fF
C1501 cs_ring_osc_0/cs_ring_osc_stage_4/voutcs cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.40fF
C1502 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y a_32042_7919# 0.11fF
C1503 VDD a_31443_5743# 0.22fF
C1504 VDD a_31527_5743# 0.02fF
C1505 VDD a_14848_n11700# 1.55fF
C1506 a_26209_7037# cs_ring_osc_0/cs_ring_osc_stage_5/vout 0.03fF
C1507 a_30745_7375# a_30579_7925# 0.09fF
C1508 a_30579_7925# a_31018_8829# 0.01fF
C1509 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q a_33443_6287# 0.03fF
C1510 cs_ring_osc_0/cs_ring_osc_stage_5/vin cs_ring_osc_0/cs_ring_osc_stage_5/csinvn 0.09fF
C1511 a_34988_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C1512 a_31018_7741# a_31611_7643# 0.02fF
C1513 freq_div_0/sky130_fd_sc_hd__inv_4_1/A freq_div_0/sky130_fd_sc_hd__inv_4_3/A 0.09fF
C1514 a_33811_7919# a_33716_7919# 0.04fF
C1515 pfd_cp_lpf_0/vQB vcp 0.07fF
C1516 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y freq_div_0/sky130_fd_sc_hd__inv_4_2/A 0.03fF
C1517 a_30745_7375# a_31443_7741# 0.44fF
C1518 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs a_30141_n18921# 0.03fF
C1519 a_30933_8463# VDD 0.15fF
C1520 a_26616_1344# a_27074_1344# 0.02fF
C1521 a_29988_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/voutcs 0.03fF
C1522 a_27287_13961# a_27453_13961# 1.60fF
C1523 a_31443_7741# a_30745_6837# 0.01fF
C1524 a_32042_8785# freq_div_0/sky130_fd_sc_hd__inv_1_0/A 0.25fF
C1525 a_33443_5749# a_34309_5717# 0.11fF
C1526 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q 0.41fF
C1527 a_34141_7919# freq_div_0/sky130_fd_sc_hd__inv_4_6/Y 0.14fF
C1528 VDD a_34141_6831# 0.22fF
C1529 VDD a_33631_6831# 0.15fF
C1530 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs a_14390_n11700# 0.82fF
C1531 a_31443_5743# freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 0.04fF
C1532 a_31018_6653# a_31018_6831# 0.08fF
C1533 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y freq_div_0/sky130_fd_sc_hd__inv_4_5/A 1.64fF
C1534 freq_div_0/sky130_fd_sc_hd__inv_4_10/Y freq_div_0/sky130_fd_sc_hd__inv_4_9/Y 0.13fF
C1535 cs_ring_osc_0/cs_ring_osc_stage_5/vout a_27124_9468# 0.03fF
C1536 a_31186_7893# a_31611_7893# 0.04fF
C1537 cs_ring_osc_0/vpbias a_27074_n16656# 0.76fF
C1538 VDD a_30745_7925# 0.43fF
C1539 a_30933_5743# a_30579_5749# 0.21fF
C1540 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y a_31611_5717# 0.17fF
C1541 VDD a_31527_6653# 0.02fF
C1542 VDD a_10700_n16656# 1.55fF
C1543 a_33443_5749# a_33884_5717# 0.28fF
C1544 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y freq_div_0/sky130_fd_sc_hd__inv_4_6/Y 0.06fF
C1545 a_30933_6831# a_30933_7375# 0.02fF
C1546 a_14240_6217# a_16072_6217# 0.67fF
C1547 a_34141_7919# a_33443_7925# 0.44fF
C1548 a_30745_7375# a_30579_7375# 2.23fF
C1549 VDD a_31186_6399# 0.23fF
C1550 cs_ring_osc_0/cs_ring_osc_stage_2/vin a_9683_n18921# 0.03fF
C1551 a_34141_7919# a_34267_8297# 0.04fF
C1552 a_34071_n9035# cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C1553 a_30745_6837# a_30579_7375# 0.02fF
C1554 VDD a_28021_14203# 0.32fF
C1555 a_33716_5743# a_33811_5743# 0.04fF
C1556 cs_ring_osc_0/vosc cs_ring_osc_0/cs_ring_osc_stage_0/csinvp 1.18fF
C1557 VDD cs_ring_osc_0/cs_ring_osc_stage_2/csinvp 0.48fF
C1558 a_33277_6287# a_33716_6831# 0.02fF
C1559 VDD a_31079_14103# 0.89fF
C1560 a_30933_5743# a_31186_5717# 0.04fF
C1561 VDD a_29107_13961# 0.29fF
C1562 a_31186_8575# a_30933_8463# 0.04fF
C1563 a_31113_5743# a_31018_5743# 0.04fF
C1564 a_33277_7375# a_33631_7375# 0.21fF
C1565 freq_div_0/vout a_27453_13961# 0.04fF
C1566 a_33631_7919# a_33277_7925# 0.21fF
C1567 cs_ring_osc_0/cs_ring_osc_stage_1/vin a_20446_n6542# 0.03fF
C1568 a_26515_n18921# cs_ring_osc_0/cs_ring_osc_stage_3/vin 0.03fF
C1569 a_25242_1344# cs_ring_osc_0/vpbias 0.51fF
C1570 a_31443_7919# a_31186_7893# 0.11fF
C1571 a_33631_7375# a_33443_7375# 0.26fF
C1572 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q a_32042_6831# 0.37fF
C1573 freq_div_0/sky130_fd_sc_hd__inv_4_2/Y a_32042_6831# 0.11fF
C1574 pfd_cp_lpf_0/vpbias ibiasn 0.05fF
C1575 a_31222_n11700# a_31680_n11700# 0.01fF
C1576 a_34309_5717# a_33277_5749# 0.11fF
C1577 VDD a_30996_14327# 0.01fF
C1578 a_31443_6831# a_32042_6831# 0.02fF
C1579 a_33277_7375# a_34309_7643# 0.11fF
C1580 vcp a_26972_n3082# 0.03fF
C1581 a_26158_n16656# a_27074_n16656# 1.92fF
C1582 a_33277_7375# freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q 0.49fF
C1583 a_32042_7919# freq_div_0/sky130_fd_sc_hd__inv_4_1/A 0.05fF
C1584 a_34072_n6542# cs_ring_osc_0/cs_ring_osc_stage_4/vin 0.03fF
C1585 a_33443_7375# a_34309_7643# 0.11fF
C1586 a_32042_8785# freq_div_0/sky130_fd_sc_hd__inv_4_0/Y 0.11fF
C1587 a_26158_n16656# cs_ring_osc_0/cs_ring_osc_stage_3/voutcs 0.22fF
C1588 VDD freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q 1.02fF
C1589 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q a_33443_7375# 0.08fF
C1590 vcp a_11972_n3082# 0.03fF
C1591 VDD a_30762_14213# 0.39fF
C1592 a_33277_7925# freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q 0.51fF
C1593 VDD a_34740_5743# 0.37fF
C1594 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs cs_ring_osc_0/cs_ring_osc_stage_5/vin 0.40fF
C1595 a_12074_n16656# a_10242_n16656# 0.65fF
C1596 a_19071_n9035# cs_ring_osc_0/cs_ring_osc_stage_1/vin 0.03fF
C1597 pfd_cp_lpf_0/vRSTN a_31380_14327# 0.06fF
C1598 a_31079_14103# a_30762_14213# 0.27fF
C1599 VDD a_31166_14327# 0.32fF
C1600 a_34740_7919# a_34740_7697# 0.04fF
C1601 a_27430_n21082# VSS 0.03fF
C1602 a_26972_n21082# VSS 0.03fF
C1603 a_26514_n21082# VSS 0.03fF
C1604 a_26056_n21082# VSS 0.03fF
C1605 a_25598_n21082# VSS 0.03fF
C1606 a_25140_n21082# VSS 0.03fF
C1607 a_24682_n21082# VSS 0.03fF
C1608 a_32430_n20414# VSS 0.03fF
C1609 a_31972_n20414# VSS 0.03fF
C1610 a_31514_n20414# VSS 0.03fF
C1611 a_31056_n20414# VSS 0.03fF
C1612 a_30598_n20414# VSS 0.03fF
C1613 a_30140_n20414# VSS 0.03fF
C1614 a_29682_n20414# VSS 0.03fF
C1615 a_27430_n20414# VSS 0.03fF
C1616 a_26972_n20414# VSS 0.03fF
C1617 a_26514_n20414# VSS 0.03fF
C1618 a_26056_n20414# VSS 0.03fF
C1619 a_25598_n20414# VSS 0.03fF
C1620 a_25140_n20414# VSS 0.03fF
C1621 cs_ring_osc_0/cs_ring_osc_stage_3/csinvn VSS 0.46fF
C1622 a_12430_n21082# VSS 0.03fF
C1623 a_11972_n21082# VSS 0.03fF
C1624 a_11514_n21082# VSS 0.03fF
C1625 a_11056_n21082# VSS 0.03fF
C1626 a_10598_n21082# VSS 0.03fF
C1627 a_10140_n21082# VSS 0.03fF
C1628 a_9682_n21082# VSS 0.03fF
C1629 a_17430_n20414# VSS 0.03fF
C1630 a_16972_n20414# VSS 0.03fF
C1631 a_16514_n20414# VSS 0.03fF
C1632 a_16056_n20414# VSS 0.03fF
C1633 a_15598_n20414# VSS 0.03fF
C1634 a_15140_n20414# VSS 0.03fF
C1635 a_14682_n20414# VSS 0.03fF
C1636 a_12430_n20414# VSS 0.03fF
C1637 a_11972_n20414# VSS 0.03fF
C1638 a_11514_n20414# VSS 0.03fF
C1639 a_11056_n20414# VSS 0.03fF
C1640 a_10598_n20414# VSS 0.03fF
C1641 a_10140_n20414# VSS 0.03fF
C1642 cs_ring_osc_0/cs_ring_osc_stage_2/csinvn VSS 0.46fF
C1643 a_32431_n18921# VSS 0.03fF
C1644 a_31973_n18921# VSS 0.03fF
C1645 a_31515_n18921# VSS 0.03fF
C1646 a_31057_n18921# VSS 0.03fF
C1647 a_30599_n18921# VSS 0.03fF
C1648 a_30141_n18921# VSS 0.03fF
C1649 a_29683_n18921# VSS 0.03fF
C1650 a_27431_n18921# VSS 0.03fF
C1651 a_26973_n18921# VSS 0.03fF
C1652 a_26515_n18921# VSS 0.03fF
C1653 a_26057_n18921# VSS 0.03fF
C1654 a_25599_n18921# VSS 0.03fF
C1655 a_25141_n18921# VSS 0.03fF
C1656 a_24683_n18921# VSS 0.03fF
C1657 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs VSS 20.26fF
C1658 cs_ring_osc_0/cs_ring_osc_stage_3/csinvp VSS 2.10fF
C1659 a_27990_n16656# VSS 0.62fF
C1660 a_27532_n16656# VSS 1.00fF
C1661 a_27074_n16656# VSS 1.48fF
C1662 a_26616_n16656# VSS 1.86fF
C1663 a_26158_n16656# VSS 2.33fF
C1664 a_25700_n16656# VSS 2.71fF
C1665 a_25242_n16656# VSS 3.19fF
C1666 cs_ring_osc_0/cs_ring_osc_stage_3/vin VSS 43.02fF
C1667 a_17431_n18921# VSS 0.03fF
C1668 a_16973_n18921# VSS 0.03fF
C1669 a_16515_n18921# VSS 0.03fF
C1670 a_16057_n18921# VSS 0.03fF
C1671 a_15599_n18921# VSS 0.03fF
C1672 a_15141_n18921# VSS 0.03fF
C1673 a_14683_n18921# VSS 0.03fF
C1674 a_12431_n18921# VSS 0.03fF
C1675 a_11973_n18921# VSS 0.03fF
C1676 a_11515_n18921# VSS 0.03fF
C1677 a_11057_n18921# VSS 0.03fF
C1678 a_10599_n18921# VSS 0.03fF
C1679 a_10141_n18921# VSS 0.03fF
C1680 a_9683_n18921# VSS 0.03fF
C1681 cs_ring_osc_0/cs_ring_osc_stage_2/voutcs VSS 20.26fF
C1682 cs_ring_osc_0/cs_ring_osc_stage_2/csinvp VSS 2.10fF
C1683 a_12990_n16656# VSS 0.62fF
C1684 a_12532_n16656# VSS 1.00fF
C1685 a_12074_n16656# VSS 1.48fF
C1686 a_11616_n16656# VSS 1.86fF
C1687 a_11158_n16656# VSS 2.33fF
C1688 a_10700_n16656# VSS 2.71fF
C1689 a_10242_n16656# VSS 3.19fF
C1690 a_32138_n11700# VSS 0.62fF
C1691 a_31680_n11700# VSS 1.00fF
C1692 a_31222_n11700# VSS 1.48fF
C1693 a_30764_n11700# VSS 1.86fF
C1694 a_30306_n11700# VSS 2.33fF
C1695 a_29848_n11700# VSS 2.71fF
C1696 a_29390_n11700# VSS 3.19fF
C1697 cs_ring_osc_0/cs_ring_osc_stage_4/csinvp VSS 2.10fF
C1698 a_36361_n9035# VSS 0.03fF
C1699 a_35903_n9035# VSS 0.03fF
C1700 a_35445_n9035# VSS 0.03fF
C1701 a_34987_n9035# VSS 0.03fF
C1702 a_34529_n9035# VSS 0.03fF
C1703 a_34071_n9035# VSS 0.03fF
C1704 a_33613_n9035# VSS 0.03fF
C1705 a_31361_n9035# VSS 0.03fF
C1706 a_30903_n9035# VSS 0.03fF
C1707 a_30445_n9035# VSS 0.03fF
C1708 a_29987_n9035# VSS 0.03fF
C1709 a_29529_n9035# VSS 0.03fF
C1710 a_29071_n9035# VSS 0.03fF
C1711 a_28613_n9035# VSS 0.03fF
C1712 a_17138_n11700# VSS 0.62fF
C1713 a_16680_n11700# VSS 1.00fF
C1714 a_16222_n11700# VSS 1.48fF
C1715 a_15764_n11700# VSS 1.86fF
C1716 a_15306_n11700# VSS 2.33fF
C1717 a_14848_n11700# VSS 2.71fF
C1718 a_14390_n11700# VSS 3.19fF
C1719 cs_ring_osc_0/cs_ring_osc_stage_1/csinvp VSS 2.10fF
C1720 a_21361_n9035# VSS 0.03fF
C1721 a_20903_n9035# VSS 0.03fF
C1722 a_20445_n9035# VSS 0.03fF
C1723 a_19987_n9035# VSS 0.03fF
C1724 a_19529_n9035# VSS 0.03fF
C1725 a_19071_n9035# VSS 0.03fF
C1726 a_18613_n9035# VSS 0.03fF
C1727 a_16361_n9035# VSS 0.03fF
C1728 a_15903_n9035# VSS 0.03fF
C1729 a_15445_n9035# VSS 0.03fF
C1730 a_14987_n9035# VSS 0.03fF
C1731 a_14529_n9035# VSS 0.03fF
C1732 a_14071_n9035# VSS 0.03fF
C1733 a_13613_n9035# VSS 0.03fF
C1734 a_36362_n6542# VSS 0.03fF
C1735 a_35904_n6542# VSS 0.03fF
C1736 a_35446_n6542# VSS 0.03fF
C1737 a_34988_n6542# VSS 0.03fF
C1738 a_34530_n6542# VSS 0.03fF
C1739 a_34072_n6542# VSS 0.03fF
C1740 a_33614_n6542# VSS 0.03fF
C1741 a_31362_n6542# VSS 0.03fF
C1742 a_30904_n6542# VSS 0.03fF
C1743 a_30446_n6542# VSS 0.03fF
C1744 a_29988_n6542# VSS 0.03fF
C1745 a_29530_n6542# VSS 0.03fF
C1746 a_29072_n6542# VSS 0.03fF
C1747 a_28614_n6542# VSS 0.03fF
C1748 cs_ring_osc_0/cs_ring_osc_stage_4/vin VSS 48.60fF
C1749 cs_ring_osc_0/cs_ring_osc_stage_4/voutcs VSS 20.26fF
C1750 cs_ring_osc_0/cs_ring_osc_stage_4/csinvn VSS 0.46fF
C1751 a_36362_n5874# VSS 0.03fF
C1752 a_35904_n5874# VSS 0.03fF
C1753 a_35446_n5874# VSS 0.03fF
C1754 a_34988_n5874# VSS 0.03fF
C1755 a_34530_n5874# VSS 0.03fF
C1756 a_34072_n5874# VSS 0.03fF
C1757 a_33614_n5874# VSS 0.03fF
C1758 a_21362_n6542# VSS 0.03fF
C1759 a_20904_n6542# VSS 0.03fF
C1760 a_20446_n6542# VSS 0.03fF
C1761 a_19988_n6542# VSS 0.03fF
C1762 a_19530_n6542# VSS 0.03fF
C1763 a_19072_n6542# VSS 0.03fF
C1764 a_18614_n6542# VSS 0.03fF
C1765 a_16362_n6542# VSS 0.03fF
C1766 a_15904_n6542# VSS 0.03fF
C1767 a_15446_n6542# VSS 0.03fF
C1768 a_14988_n6542# VSS 0.03fF
C1769 a_14530_n6542# VSS 0.03fF
C1770 a_14072_n6542# VSS 0.03fF
C1771 a_13614_n6542# VSS 0.03fF
C1772 cs_ring_osc_0/cs_ring_osc_stage_2/vin VSS 1.00fF
C1773 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs VSS 20.26fF
C1774 cs_ring_osc_0/cs_ring_osc_stage_1/csinvn VSS 0.46fF
C1775 a_21362_n5874# VSS 0.03fF
C1776 a_20904_n5874# VSS 0.03fF
C1777 a_20446_n5874# VSS 0.03fF
C1778 a_19988_n5874# VSS 0.03fF
C1779 a_19530_n5874# VSS 0.03fF
C1780 a_19072_n5874# VSS 0.03fF
C1781 a_18614_n5874# VSS 0.03fF
C1782 a_27430_n3082# VSS 0.03fF
C1783 a_26972_n3082# VSS 0.03fF
C1784 a_26514_n3082# VSS 0.03fF
C1785 a_26056_n3082# VSS 0.03fF
C1786 a_25598_n3082# VSS 0.03fF
C1787 a_25140_n3082# VSS 0.03fF
C1788 a_32430_n2414# VSS 0.03fF
C1789 a_31972_n2414# VSS 0.03fF
C1790 a_31514_n2414# VSS 0.03fF
C1791 a_31056_n2414# VSS 0.03fF
C1792 a_30598_n2414# VSS 0.03fF
C1793 a_30140_n2414# VSS 0.03fF
C1794 a_29682_n2414# VSS 0.03fF
C1795 a_27430_n2414# VSS 0.03fF
C1796 a_26972_n2414# VSS 0.03fF
C1797 a_26514_n2414# VSS 0.03fF
C1798 a_26056_n2414# VSS 0.03fF
C1799 a_25598_n2414# VSS 0.03fF
C1800 a_25140_n2414# VSS 0.03fF
C1801 cs_ring_osc_0/cs_ring_osc_stage_5/csinvn VSS 0.46fF
C1802 a_12430_n3082# VSS 0.03fF
C1803 a_11972_n3082# VSS 0.03fF
C1804 a_11514_n3082# VSS 0.03fF
C1805 a_11056_n3082# VSS 0.03fF
C1806 a_10598_n3082# VSS 0.03fF
C1807 a_10140_n3082# VSS 0.03fF
C1808 a_17430_n2414# VSS 0.03fF
C1809 a_16972_n2414# VSS 0.03fF
C1810 a_16514_n2414# VSS 0.03fF
C1811 a_16056_n2414# VSS 0.03fF
C1812 a_15598_n2414# VSS 0.03fF
C1813 a_15140_n2414# VSS 0.03fF
C1814 a_14682_n2414# VSS 0.03fF
C1815 a_12430_n2414# VSS 0.03fF
C1816 a_11972_n2414# VSS 0.03fF
C1817 a_11514_n2414# VSS 0.03fF
C1818 a_11056_n2414# VSS 0.03fF
C1819 a_10598_n2414# VSS 0.03fF
C1820 a_10140_n2414# VSS 0.03fF
C1821 cs_ring_osc_0/cs_ring_osc_stage_0/csinvn VSS 0.46fF
C1822 a_32431_n921# VSS 0.03fF
C1823 a_31973_n921# VSS 0.03fF
C1824 a_31515_n921# VSS 0.03fF
C1825 a_31057_n921# VSS 0.03fF
C1826 a_30599_n921# VSS 0.03fF
C1827 a_30141_n921# VSS 0.03fF
C1828 a_29683_n921# VSS 0.03fF
C1829 a_27431_n921# VSS 0.03fF
C1830 a_26973_n921# VSS 0.03fF
C1831 a_26515_n921# VSS 0.03fF
C1832 a_26057_n921# VSS 0.03fF
C1833 a_25599_n921# VSS 0.03fF
C1834 a_25141_n921# VSS 0.03fF
C1835 a_24683_n921# VSS 0.03fF
C1836 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs VSS 20.26fF
C1837 cs_ring_osc_0/cs_ring_osc_stage_5/vin VSS 1.00fF
C1838 cs_ring_osc_0/cs_ring_osc_stage_5/csinvp VSS 2.10fF
C1839 a_27990_1344# VSS 0.62fF
C1840 a_27532_1344# VSS 1.00fF
C1841 a_27074_1344# VSS 1.48fF
C1842 a_26616_1344# VSS 1.86fF
C1843 a_26158_1344# VSS 2.33fF
C1844 a_25700_1344# VSS 2.71fF
C1845 a_25242_1344# VSS 3.19fF
C1846 cs_ring_osc_0/cs_ring_osc_stage_1/vin VSS 47.79fF
C1847 a_17431_n921# VSS 0.03fF
C1848 a_16973_n921# VSS 0.03fF
C1849 a_16515_n921# VSS 0.03fF
C1850 a_16057_n921# VSS 0.03fF
C1851 a_15599_n921# VSS 0.03fF
C1852 a_15141_n921# VSS 0.03fF
C1853 a_14683_n921# VSS 0.03fF
C1854 a_12431_n921# VSS 0.03fF
C1855 a_11973_n921# VSS 0.03fF
C1856 a_11515_n921# VSS 0.03fF
C1857 a_11057_n921# VSS 0.03fF
C1858 a_10599_n921# VSS 0.03fF
C1859 a_10141_n921# VSS 0.03fF
C1860 a_9683_n921# VSS 0.03fF
C1861 cs_ring_osc_0/cs_ring_osc_stage_0/voutcs VSS 20.26fF
C1862 cs_ring_osc_0/cs_ring_osc_stage_0/csinvp VSS 2.10fF
C1863 a_12990_1344# VSS 0.62fF
C1864 a_12532_1344# VSS 1.00fF
C1865 a_12074_1344# VSS 1.48fF
C1866 a_11616_1344# VSS 1.86fF
C1867 a_11158_1344# VSS 2.33fF
C1868 a_10700_1344# VSS 2.71fF
C1869 a_10242_1344# VSS 3.19fF
C1870 a_34267_6121# VSS 0.01fF
C1871 a_33842_6121# VSS 0.01fF
C1872 a_33631_5743# VSS 0.20fF
C1873 a_31569_6121# VSS 0.01fF
C1874 a_31144_6121# VSS 0.01fF
C1875 a_30933_5743# VSS 0.20fF
C1876 freq_div_0/sky130_fd_sc_hd__inv_4_10/A VSS 1.38fF
C1877 freq_div_0/sky130_fd_sc_hd__inv_1_10/A VSS 0.71fF
C1878 a_34740_5743# VSS 0.49fF
C1879 a_34141_5743# VSS 0.60fF
C1880 a_34309_5717# VSS 1.13fF
C1881 a_33716_5743# VSS 0.49fF
C1882 a_33884_5717# VSS 0.61fF
C1883 a_33443_5749# VSS 1.17fF
C1884 freq_div_0/sky130_fd_sc_hd__inv_4_10/Y VSS 1.31fF
C1885 a_33277_5749# VSS 1.51fF
C1886 freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q VSS 0.74fF
C1887 freq_div_0/sky130_fd_sc_hd__inv_4_5/A VSS 1.38fF
C1888 freq_div_0/sky130_fd_sc_hd__inv_1_5/A VSS 0.71fF
C1889 a_32042_5743# VSS 0.49fF
C1890 a_31443_5743# VSS 0.60fF
C1891 a_31611_5717# VSS 1.13fF
C1892 a_31018_5743# VSS 0.49fF
C1893 a_31186_5717# VSS 0.61fF
C1894 a_30745_5749# VSS 1.17fF
C1895 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y VSS 1.30fF
C1896 a_30579_5749# VSS 1.52fF
C1897 a_34267_6287# VSS 0.01fF
C1898 a_33842_6287# VSS 0.01fF
C1899 a_31569_6287# VSS 0.01fF
C1900 a_33631_6287# VSS 0.20fF
C1901 freq_div_0/sky130_fd_sc_hd__inv_4_9/A VSS 0.23fF
C1902 freq_div_0/sky130_fd_sc_hd__inv_1_9/A VSS 0.41fF
C1903 a_34740_6609# VSS 0.31fF
C1904 a_34141_6653# VSS 0.60fF
C1905 a_34309_6555# VSS 1.13fF
C1906 a_33716_6653# VSS 0.49fF
C1907 a_33884_6399# VSS 0.61fF
C1908 a_33443_6287# VSS 0.16fF
C1909 freq_div_0/sky130_fd_sc_hd__inv_4_9/Y VSS 0.25fF
C1910 a_33277_6287# VSS 0.34fF
C1911 freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q VSS 0.30fF
C1912 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q VSS 2.28fF
C1913 a_31144_6287# VSS 0.01fF
C1914 a_30933_6287# VSS 0.20fF
C1915 freq_div_0/sky130_fd_sc_hd__inv_4_4/A VSS 0.06fF
C1916 freq_div_0/sky130_fd_sc_hd__inv_1_4/A VSS 0.41fF
C1917 a_32042_6609# VSS 0.31fF
C1918 a_31443_6653# VSS 0.60fF
C1919 a_31611_6555# VSS 1.13fF
C1920 a_31018_6653# VSS 0.49fF
C1921 a_31186_6399# VSS 0.61fF
C1922 a_30745_6287# VSS 0.16fF
C1923 freq_div_0/sky130_fd_sc_hd__inv_4_4/Y VSS 0.25fF
C1924 a_30579_6287# VSS 0.34fF
C1925 a_34267_7209# VSS 0.01fF
C1926 a_33842_7209# VSS 0.01fF
C1927 a_33631_6831# VSS 0.20fF
C1928 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q VSS 0.30fF
C1929 a_31569_7209# VSS 0.01fF
C1930 a_31144_7209# VSS 0.01fF
C1931 a_30933_6831# VSS 0.20fF
C1932 freq_div_0/sky130_fd_sc_hd__inv_4_8/A VSS 0.18fF
C1933 freq_div_0/sky130_fd_sc_hd__inv_1_8/A VSS 0.34fF
C1934 a_34740_6831# VSS 0.24fF
C1935 a_34141_6831# VSS 0.60fF
C1936 a_34309_6805# VSS 1.13fF
C1937 a_33716_6831# VSS 0.49fF
C1938 a_33884_6805# VSS 0.61fF
C1939 a_33443_6837# VSS 0.11fF
C1940 freq_div_0/sky130_fd_sc_hd__inv_4_8/Y VSS 0.19fF
C1941 a_33277_6837# VSS 0.25fF
C1942 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q VSS 0.20fF
C1943 freq_div_0/sky130_fd_sc_hd__inv_4_2/A VSS 0.05fF
C1944 freq_div_0/sky130_fd_sc_hd__inv_1_2/A VSS 0.34fF
C1945 a_32042_6831# VSS 0.24fF
C1946 a_31443_6831# VSS 0.60fF
C1947 a_31611_6805# VSS 1.13fF
C1948 a_31018_6831# VSS 0.49fF
C1949 a_31186_6805# VSS 0.61fF
C1950 a_30745_6837# VSS 0.11fF
C1951 freq_div_0/sky130_fd_sc_hd__inv_4_2/Y VSS 0.19fF
C1952 a_30579_6837# VSS 0.25fF
C1953 a_34267_7375# VSS 0.01fF
C1954 a_33842_7375# VSS 0.01fF
C1955 a_31569_7375# VSS 0.01fF
C1956 a_33631_7375# VSS 0.20fF
C1957 freq_div_0/sky130_fd_sc_hd__inv_4_7/A VSS 0.23fF
C1958 freq_div_0/sky130_fd_sc_hd__inv_1_7/A VSS 0.41fF
C1959 a_34740_7697# VSS 0.31fF
C1960 a_34141_7741# VSS 0.60fF
C1961 a_34309_7643# VSS 1.13fF
C1962 a_33716_7741# VSS 0.49fF
C1963 a_33884_7487# VSS 0.61fF
C1964 a_33443_7375# VSS 0.16fF
C1965 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y VSS 0.25fF
C1966 a_33277_7375# VSS 0.34fF
C1967 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q VSS 0.30fF
C1968 freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q VSS 0.26fF
C1969 a_31144_7375# VSS 0.01fF
C1970 a_30933_7375# VSS 0.20fF
C1971 freq_div_0/sky130_fd_sc_hd__inv_4_3/A VSS 0.06fF
C1972 freq_div_0/sky130_fd_sc_hd__inv_1_3/A VSS 0.41fF
C1973 a_32042_7697# VSS 0.31fF
C1974 a_31443_7741# VSS 0.60fF
C1975 a_31611_7643# VSS 1.13fF
C1976 a_31018_7741# VSS 0.49fF
C1977 a_31186_7487# VSS 0.61fF
C1978 a_30745_7375# VSS 0.16fF
C1979 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y VSS 0.25fF
C1980 a_30579_7375# VSS 0.34fF
C1981 a_34267_8297# VSS 0.01fF
C1982 a_33842_8297# VSS 0.01fF
C1983 a_33631_7919# VSS 0.20fF
C1984 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q VSS 0.30fF
C1985 a_31569_8297# VSS 0.01fF
C1986 a_31144_8297# VSS 0.01fF
C1987 a_30933_7919# VSS 0.20fF
C1988 freq_div_0/sky130_fd_sc_hd__inv_4_6/A VSS 0.23fF
C1989 freq_div_0/sky130_fd_sc_hd__inv_1_6/A VSS 0.41fF
C1990 a_34740_7919# VSS 0.31fF
C1991 a_34141_7919# VSS 0.60fF
C1992 a_34309_7893# VSS 1.13fF
C1993 a_33716_7919# VSS 0.49fF
C1994 a_33884_7893# VSS 0.61fF
C1995 a_33443_7925# VSS 0.16fF
C1996 freq_div_0/sky130_fd_sc_hd__inv_4_6/Y VSS 0.25fF
C1997 a_33277_7925# VSS 0.34fF
C1998 freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q VSS 0.30fF
C1999 freq_div_0/sky130_fd_sc_hd__inv_4_1/A VSS 0.06fF
C2000 freq_div_0/sky130_fd_sc_hd__inv_1_1/A VSS 0.41fF
C2001 a_32042_7919# VSS 0.31fF
C2002 a_31443_7919# VSS 0.60fF
C2003 a_31611_7893# VSS 1.13fF
C2004 a_31018_7919# VSS 0.49fF
C2005 a_31186_7893# VSS 0.61fF
C2006 a_30745_7925# VSS 0.16fF
C2007 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y VSS 0.25fF
C2008 a_30579_7925# VSS 0.34fF
C2009 a_31569_8463# VSS 0.01fF
C2010 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q VSS 0.40fF
C2011 a_31144_8463# VSS 0.01fF
C2012 a_27583_7037# VSS 0.03fF
C2013 a_27125_7037# VSS 0.03fF
C2014 a_26667_7037# VSS 0.03fF
C2015 a_26209_7037# VSS 0.03fF
C2016 a_25751_7037# VSS 0.03fF
C2017 a_25293_7037# VSS 0.03fF
C2018 a_24835_7037# VSS 0.03fF
C2019 a_16988_6217# VSS 0.62fF
C2020 a_16530_6217# VSS 1.00fF
C2021 a_16072_6217# VSS 1.48fF
C2022 a_15614_6217# VSS 1.86fF
C2023 a_15156_6217# VSS 2.33fF
C2024 a_14698_6217# VSS 2.70fF
C2025 a_14240_6217# VSS 3.19fF
C2026 a_30933_8463# VSS 0.20fF
C2027 cs_ring_osc_0/vosc2 VSS 1.28fF
C2028 freq_div_0/sky130_fd_sc_hd__inv_4_0/A VSS 0.01fF
C2029 freq_div_0/sky130_fd_sc_hd__inv_1_0/A VSS 0.04fF
C2030 a_32042_8785# VSS 0.49fF
C2031 a_31443_8829# VSS 0.60fF
C2032 a_31611_8731# VSS 1.13fF
C2033 a_31018_8829# VSS 0.49fF
C2034 a_31186_8575# VSS 0.61fF
C2035 a_30745_8463# VSS 1.17fF
C2036 freq_div_0/sky130_fd_sc_hd__inv_4_0/Y VSS 0.25fF
C2037 a_30579_8463# VSS 1.52fF
C2038 freq_div_0/vin VSS 1.65fF
C2039 cs_ring_osc_0/vosc VSS 0.91fF
C2040 a_27582_9468# VSS 0.03fF
C2041 a_27124_9468# VSS 0.03fF
C2042 a_26666_9468# VSS 0.03fF
C2043 a_26208_9468# VSS 0.03fF
C2044 a_25750_9468# VSS 0.03fF
C2045 a_25292_9468# VSS 0.03fF
C2046 a_24834_9468# VSS 0.03fF
C2047 cs_ring_osc_0/cs_ring_osc_stage_5/vout VSS 48.36fF
C2048 a_18820_9468# VSS 0.03fF
C2049 a_18362_9468# VSS 0.03fF
C2050 a_17904_9468# VSS 0.03fF
C2051 a_17446_9468# VSS 0.03fF
C2052 a_16988_9468# VSS 0.03fF
C2053 a_16530_9468# VSS 0.03fF
C2054 a_16072_9468# VSS 0.03fF
C2055 cs_ring_osc_0/vpbias VSS 128.39fF
C2056 ibiasn VSS 18.07fF
C2057 a_31037_13961# VSS -0.01fF
C2058 a_30797_13961# VSS -0.01fF
C2059 vsigin VSS 0.13fF
C2060 a_31798_14327# VSS 0.23fF
C2061 a_31380_14327# VSS 0.11fF
C2062 a_28477_13961# VSS -0.01fF
C2063 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N VSS 0.07fF
C2064 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N VSS 0.07fF
C2065 pfd_cp_lpf_0/VQBb VSS 4.27fF
C2066 pfd_cp_lpf_0/vswitchl VSS 0.15fF
C2067 a_27911_14327# VSS 0.11fF
C2068 a_27708_13961# VSS 0.03fF
C2069 a_31166_14327# VSS 0.58fF
C2070 a_31235_14198# VSS 0.68fF
C2071 a_31079_14103# VSS -1.10fF
C2072 a_31040_14229# VSS 1.28fF
C2073 a_30762_14213# VSS 0.22fF
C2074 a_30391_13935# VSS 0.45fF
C2075 a_30294_13935# VSS 0.12fF
C2076 pfd_cp_lpf_0/vQB VSS 0.29fF
C2077 a_29107_13961# VSS 0.12fF
C2078 a_28368_13961# VSS -0.80fF
C2079 a_28543_13935# VSS -1.25fF
C2080 a_27803_13961# VSS 0.11fF
C2081 pfd_cp_lpf_0/vRSTN VSS -2.87fF
C2082 a_28021_14203# VSS 0.58fF
C2083 a_27453_13961# VSS 0.05fF
C2084 a_27287_13961# VSS 0.40fF
C2085 freq_div_0/vout VSS 0.13fF
C2086 pfd_cp_lpf_0/vndiode VSS 1.36fF
C2087 pfd_cp_lpf_0/vpdiode VSS 0.90fF
C2088 pfd_cp_lpf_0/vQA VSS 2.66fF
C2089 vcp VSS 110.97fF
C2090 pfd_cp_lpf_0/vQAb VSS 2.62fF
C2091 pfd_cp_lpf_0/vswitchh VSS 7.07fF
C2092 pfd_cp_lpf_0/vpbias VSS 24.46fF
C2093 VDD VSS 1995.79fF
.ends

