magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< error_p >>
rect -2101 -400 2101 400
<< nwell >>
rect -2101 -400 2101 400
<< pmoslvt >>
rect -2007 -300 -1047 300
rect -989 -300 -29 300
rect 29 -300 989 300
rect 1047 -300 2007 300
<< pdiff >>
rect -2065 288 -2007 300
rect -2065 -288 -2053 288
rect -2019 -288 -2007 288
rect -2065 -300 -2007 -288
rect -1047 288 -989 300
rect -1047 -288 -1035 288
rect -1001 -288 -989 288
rect -1047 -300 -989 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 989 288 1047 300
rect 989 -288 1001 288
rect 1035 -288 1047 288
rect 989 -300 1047 -288
rect 2007 288 2065 300
rect 2007 -288 2019 288
rect 2053 -288 2065 288
rect 2007 -300 2065 -288
<< pdiffc >>
rect -2053 -288 -2019 288
rect -1035 -288 -1001 288
rect -17 -288 17 288
rect 1001 -288 1035 288
rect 2019 -288 2053 288
<< poly >>
rect -1821 381 -1233 397
rect -1821 364 -1805 381
rect -2007 347 -1805 364
rect -1249 364 -1233 381
rect -803 381 -215 397
rect -803 364 -787 381
rect -1249 347 -1047 364
rect -2007 300 -1047 347
rect -989 347 -787 364
rect -231 364 -215 381
rect 215 381 803 397
rect 215 364 231 381
rect -231 347 -29 364
rect -989 300 -29 347
rect 29 347 231 364
rect 787 364 803 381
rect 1233 381 1821 397
rect 1233 364 1249 381
rect 787 347 989 364
rect 29 300 989 347
rect 1047 347 1249 364
rect 1805 364 1821 381
rect 1805 347 2007 364
rect 1047 300 2007 347
rect -2007 -347 -1047 -300
rect -2007 -364 -1805 -347
rect -1821 -381 -1805 -364
rect -1249 -364 -1047 -347
rect -989 -347 -29 -300
rect -989 -364 -787 -347
rect -1249 -381 -1233 -364
rect -1821 -397 -1233 -381
rect -803 -381 -787 -364
rect -231 -364 -29 -347
rect 29 -347 989 -300
rect 29 -364 231 -347
rect -231 -381 -215 -364
rect -803 -397 -215 -381
rect 215 -381 231 -364
rect 787 -364 989 -347
rect 1047 -347 2007 -300
rect 1047 -364 1249 -347
rect 787 -381 803 -364
rect 215 -397 803 -381
rect 1233 -381 1249 -364
rect 1805 -364 2007 -347
rect 1805 -381 1821 -364
rect 1233 -397 1821 -381
<< polycont >>
rect -1805 347 -1249 381
rect -787 347 -231 381
rect 231 347 787 381
rect 1249 347 1805 381
rect -1805 -381 -1249 -347
rect -787 -381 -231 -347
rect 231 -381 787 -347
rect 1249 -381 1805 -347
<< locali >>
rect -1821 347 -1805 381
rect -1249 347 -1233 381
rect -803 347 -787 381
rect -231 347 -215 381
rect 215 347 231 381
rect 787 347 803 381
rect 1233 347 1249 381
rect 1805 347 1821 381
rect -2053 288 -2019 304
rect -2053 -304 -2019 -288
rect -1035 288 -1001 304
rect -1035 -304 -1001 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 1001 288 1035 304
rect 1001 -304 1035 -288
rect 2019 288 2053 304
rect 2019 -304 2053 -288
rect -1821 -381 -1805 -347
rect -1249 -381 -1233 -347
rect -803 -381 -787 -347
rect -231 -381 -215 -347
rect 215 -381 231 -347
rect 787 -381 803 -347
rect 1233 -381 1249 -347
rect 1805 -381 1821 -347
<< viali >>
rect -1759 347 -1295 381
rect -741 347 -277 381
rect 277 347 741 381
rect 1295 347 1759 381
rect -2053 -288 -2019 288
rect -1035 -288 -1001 288
rect -17 -288 17 288
rect 1001 -288 1035 288
rect 2019 -288 2053 288
rect -1759 -381 -1295 -347
rect -741 -381 -277 -347
rect 277 -381 741 -347
rect 1295 -381 1759 -347
<< metal1 >>
rect -1771 381 -1283 387
rect -1771 347 -1759 381
rect -1295 347 -1283 381
rect -1771 341 -1283 347
rect -753 381 -265 387
rect -753 347 -741 381
rect -277 347 -265 381
rect -753 341 -265 347
rect 265 381 753 387
rect 265 347 277 381
rect 741 347 753 381
rect 265 341 753 347
rect 1283 381 1771 387
rect 1283 347 1295 381
rect 1759 347 1771 381
rect 1283 341 1771 347
rect -2059 288 -2013 300
rect -2059 -288 -2053 288
rect -2019 -288 -2013 288
rect -2059 -300 -2013 -288
rect -1041 288 -995 300
rect -1041 -288 -1035 288
rect -1001 -288 -995 288
rect -1041 -300 -995 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 995 288 1041 300
rect 995 -288 1001 288
rect 1035 -288 1041 288
rect 995 -300 1041 -288
rect 2013 288 2059 300
rect 2013 -288 2019 288
rect 2053 -288 2059 288
rect 2013 -300 2059 -288
rect -1771 -347 -1283 -341
rect -1771 -381 -1759 -347
rect -1295 -381 -1283 -347
rect -1771 -387 -1283 -381
rect -753 -347 -265 -341
rect -753 -381 -741 -347
rect -277 -381 -265 -347
rect -753 -387 -265 -381
rect 265 -347 753 -341
rect 265 -381 277 -347
rect 741 -381 753 -347
rect 265 -387 753 -381
rect 1283 -347 1771 -341
rect 1283 -381 1295 -347
rect 1759 -381 1771 -347
rect 1283 -387 1771 -381
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 3 l 4.8 m 1 nf 4 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
