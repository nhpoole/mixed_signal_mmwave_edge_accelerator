magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -3131 -1460 3131 1460
<< nwell >>
rect -1871 -200 1871 200
<< pmos >>
rect -1777 -100 -1577 100
rect -1519 -100 -1319 100
rect -1261 -100 -1061 100
rect -1003 -100 -803 100
rect -745 -100 -545 100
rect -487 -100 -287 100
rect -229 -100 -29 100
rect 29 -100 229 100
rect 287 -100 487 100
rect 545 -100 745 100
rect 803 -100 1003 100
rect 1061 -100 1261 100
rect 1319 -100 1519 100
rect 1577 -100 1777 100
<< pdiff >>
rect -1835 85 -1777 100
rect -1835 51 -1823 85
rect -1789 51 -1777 85
rect -1835 17 -1777 51
rect -1835 -17 -1823 17
rect -1789 -17 -1777 17
rect -1835 -51 -1777 -17
rect -1835 -85 -1823 -51
rect -1789 -85 -1777 -51
rect -1835 -100 -1777 -85
rect -1577 85 -1519 100
rect -1577 51 -1565 85
rect -1531 51 -1519 85
rect -1577 17 -1519 51
rect -1577 -17 -1565 17
rect -1531 -17 -1519 17
rect -1577 -51 -1519 -17
rect -1577 -85 -1565 -51
rect -1531 -85 -1519 -51
rect -1577 -100 -1519 -85
rect -1319 85 -1261 100
rect -1319 51 -1307 85
rect -1273 51 -1261 85
rect -1319 17 -1261 51
rect -1319 -17 -1307 17
rect -1273 -17 -1261 17
rect -1319 -51 -1261 -17
rect -1319 -85 -1307 -51
rect -1273 -85 -1261 -51
rect -1319 -100 -1261 -85
rect -1061 85 -1003 100
rect -1061 51 -1049 85
rect -1015 51 -1003 85
rect -1061 17 -1003 51
rect -1061 -17 -1049 17
rect -1015 -17 -1003 17
rect -1061 -51 -1003 -17
rect -1061 -85 -1049 -51
rect -1015 -85 -1003 -51
rect -1061 -100 -1003 -85
rect -803 85 -745 100
rect -803 51 -791 85
rect -757 51 -745 85
rect -803 17 -745 51
rect -803 -17 -791 17
rect -757 -17 -745 17
rect -803 -51 -745 -17
rect -803 -85 -791 -51
rect -757 -85 -745 -51
rect -803 -100 -745 -85
rect -545 85 -487 100
rect -545 51 -533 85
rect -499 51 -487 85
rect -545 17 -487 51
rect -545 -17 -533 17
rect -499 -17 -487 17
rect -545 -51 -487 -17
rect -545 -85 -533 -51
rect -499 -85 -487 -51
rect -545 -100 -487 -85
rect -287 85 -229 100
rect -287 51 -275 85
rect -241 51 -229 85
rect -287 17 -229 51
rect -287 -17 -275 17
rect -241 -17 -229 17
rect -287 -51 -229 -17
rect -287 -85 -275 -51
rect -241 -85 -229 -51
rect -287 -100 -229 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 229 85 287 100
rect 229 51 241 85
rect 275 51 287 85
rect 229 17 287 51
rect 229 -17 241 17
rect 275 -17 287 17
rect 229 -51 287 -17
rect 229 -85 241 -51
rect 275 -85 287 -51
rect 229 -100 287 -85
rect 487 85 545 100
rect 487 51 499 85
rect 533 51 545 85
rect 487 17 545 51
rect 487 -17 499 17
rect 533 -17 545 17
rect 487 -51 545 -17
rect 487 -85 499 -51
rect 533 -85 545 -51
rect 487 -100 545 -85
rect 745 85 803 100
rect 745 51 757 85
rect 791 51 803 85
rect 745 17 803 51
rect 745 -17 757 17
rect 791 -17 803 17
rect 745 -51 803 -17
rect 745 -85 757 -51
rect 791 -85 803 -51
rect 745 -100 803 -85
rect 1003 85 1061 100
rect 1003 51 1015 85
rect 1049 51 1061 85
rect 1003 17 1061 51
rect 1003 -17 1015 17
rect 1049 -17 1061 17
rect 1003 -51 1061 -17
rect 1003 -85 1015 -51
rect 1049 -85 1061 -51
rect 1003 -100 1061 -85
rect 1261 85 1319 100
rect 1261 51 1273 85
rect 1307 51 1319 85
rect 1261 17 1319 51
rect 1261 -17 1273 17
rect 1307 -17 1319 17
rect 1261 -51 1319 -17
rect 1261 -85 1273 -51
rect 1307 -85 1319 -51
rect 1261 -100 1319 -85
rect 1519 85 1577 100
rect 1519 51 1531 85
rect 1565 51 1577 85
rect 1519 17 1577 51
rect 1519 -17 1531 17
rect 1565 -17 1577 17
rect 1519 -51 1577 -17
rect 1519 -85 1531 -51
rect 1565 -85 1577 -51
rect 1519 -100 1577 -85
rect 1777 85 1835 100
rect 1777 51 1789 85
rect 1823 51 1835 85
rect 1777 17 1835 51
rect 1777 -17 1789 17
rect 1823 -17 1835 17
rect 1777 -51 1835 -17
rect 1777 -85 1789 -51
rect 1823 -85 1835 -51
rect 1777 -100 1835 -85
<< pdiffc >>
rect -1823 51 -1789 85
rect -1823 -17 -1789 17
rect -1823 -85 -1789 -51
rect -1565 51 -1531 85
rect -1565 -17 -1531 17
rect -1565 -85 -1531 -51
rect -1307 51 -1273 85
rect -1307 -17 -1273 17
rect -1307 -85 -1273 -51
rect -1049 51 -1015 85
rect -1049 -17 -1015 17
rect -1049 -85 -1015 -51
rect -791 51 -757 85
rect -791 -17 -757 17
rect -791 -85 -757 -51
rect -533 51 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -51
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
rect 499 51 533 85
rect 499 -17 533 17
rect 499 -85 533 -51
rect 757 51 791 85
rect 757 -17 791 17
rect 757 -85 791 -51
rect 1015 51 1049 85
rect 1015 -17 1049 17
rect 1015 -85 1049 -51
rect 1273 51 1307 85
rect 1273 -17 1307 17
rect 1273 -85 1307 -51
rect 1531 51 1565 85
rect 1531 -17 1565 17
rect 1531 -85 1565 -51
rect 1789 51 1823 85
rect 1789 -17 1823 17
rect 1789 -85 1823 -51
<< poly >>
rect -1743 181 -1611 197
rect -1743 164 -1694 181
rect -1777 147 -1694 164
rect -1660 164 -1611 181
rect -1485 181 -1353 197
rect -1485 164 -1436 181
rect -1660 147 -1577 164
rect -1777 100 -1577 147
rect -1519 147 -1436 164
rect -1402 164 -1353 181
rect -1227 181 -1095 197
rect -1227 164 -1178 181
rect -1402 147 -1319 164
rect -1519 100 -1319 147
rect -1261 147 -1178 164
rect -1144 164 -1095 181
rect -969 181 -837 197
rect -969 164 -920 181
rect -1144 147 -1061 164
rect -1261 100 -1061 147
rect -1003 147 -920 164
rect -886 164 -837 181
rect -711 181 -579 197
rect -711 164 -662 181
rect -886 147 -803 164
rect -1003 100 -803 147
rect -745 147 -662 164
rect -628 164 -579 181
rect -453 181 -321 197
rect -453 164 -404 181
rect -628 147 -545 164
rect -745 100 -545 147
rect -487 147 -404 164
rect -370 164 -321 181
rect -195 181 -63 197
rect -195 164 -146 181
rect -370 147 -287 164
rect -487 100 -287 147
rect -229 147 -146 164
rect -112 164 -63 181
rect 63 181 195 197
rect 63 164 112 181
rect -112 147 -29 164
rect -229 100 -29 147
rect 29 147 112 164
rect 146 164 195 181
rect 321 181 453 197
rect 321 164 370 181
rect 146 147 229 164
rect 29 100 229 147
rect 287 147 370 164
rect 404 164 453 181
rect 579 181 711 197
rect 579 164 628 181
rect 404 147 487 164
rect 287 100 487 147
rect 545 147 628 164
rect 662 164 711 181
rect 837 181 969 197
rect 837 164 886 181
rect 662 147 745 164
rect 545 100 745 147
rect 803 147 886 164
rect 920 164 969 181
rect 1095 181 1227 197
rect 1095 164 1144 181
rect 920 147 1003 164
rect 803 100 1003 147
rect 1061 147 1144 164
rect 1178 164 1227 181
rect 1353 181 1485 197
rect 1353 164 1402 181
rect 1178 147 1261 164
rect 1061 100 1261 147
rect 1319 147 1402 164
rect 1436 164 1485 181
rect 1611 181 1743 197
rect 1611 164 1660 181
rect 1436 147 1519 164
rect 1319 100 1519 147
rect 1577 147 1660 164
rect 1694 164 1743 181
rect 1694 147 1777 164
rect 1577 100 1777 147
rect -1777 -147 -1577 -100
rect -1777 -164 -1694 -147
rect -1743 -181 -1694 -164
rect -1660 -164 -1577 -147
rect -1519 -147 -1319 -100
rect -1519 -164 -1436 -147
rect -1660 -181 -1611 -164
rect -1743 -197 -1611 -181
rect -1485 -181 -1436 -164
rect -1402 -164 -1319 -147
rect -1261 -147 -1061 -100
rect -1261 -164 -1178 -147
rect -1402 -181 -1353 -164
rect -1485 -197 -1353 -181
rect -1227 -181 -1178 -164
rect -1144 -164 -1061 -147
rect -1003 -147 -803 -100
rect -1003 -164 -920 -147
rect -1144 -181 -1095 -164
rect -1227 -197 -1095 -181
rect -969 -181 -920 -164
rect -886 -164 -803 -147
rect -745 -147 -545 -100
rect -745 -164 -662 -147
rect -886 -181 -837 -164
rect -969 -197 -837 -181
rect -711 -181 -662 -164
rect -628 -164 -545 -147
rect -487 -147 -287 -100
rect -487 -164 -404 -147
rect -628 -181 -579 -164
rect -711 -197 -579 -181
rect -453 -181 -404 -164
rect -370 -164 -287 -147
rect -229 -147 -29 -100
rect -229 -164 -146 -147
rect -370 -181 -321 -164
rect -453 -197 -321 -181
rect -195 -181 -146 -164
rect -112 -164 -29 -147
rect 29 -147 229 -100
rect 29 -164 112 -147
rect -112 -181 -63 -164
rect -195 -197 -63 -181
rect 63 -181 112 -164
rect 146 -164 229 -147
rect 287 -147 487 -100
rect 287 -164 370 -147
rect 146 -181 195 -164
rect 63 -197 195 -181
rect 321 -181 370 -164
rect 404 -164 487 -147
rect 545 -147 745 -100
rect 545 -164 628 -147
rect 404 -181 453 -164
rect 321 -197 453 -181
rect 579 -181 628 -164
rect 662 -164 745 -147
rect 803 -147 1003 -100
rect 803 -164 886 -147
rect 662 -181 711 -164
rect 579 -197 711 -181
rect 837 -181 886 -164
rect 920 -164 1003 -147
rect 1061 -147 1261 -100
rect 1061 -164 1144 -147
rect 920 -181 969 -164
rect 837 -197 969 -181
rect 1095 -181 1144 -164
rect 1178 -164 1261 -147
rect 1319 -147 1519 -100
rect 1319 -164 1402 -147
rect 1178 -181 1227 -164
rect 1095 -197 1227 -181
rect 1353 -181 1402 -164
rect 1436 -164 1519 -147
rect 1577 -147 1777 -100
rect 1577 -164 1660 -147
rect 1436 -181 1485 -164
rect 1353 -197 1485 -181
rect 1611 -181 1660 -164
rect 1694 -164 1777 -147
rect 1694 -181 1743 -164
rect 1611 -197 1743 -181
<< polycont >>
rect -1694 147 -1660 181
rect -1436 147 -1402 181
rect -1178 147 -1144 181
rect -920 147 -886 181
rect -662 147 -628 181
rect -404 147 -370 181
rect -146 147 -112 181
rect 112 147 146 181
rect 370 147 404 181
rect 628 147 662 181
rect 886 147 920 181
rect 1144 147 1178 181
rect 1402 147 1436 181
rect 1660 147 1694 181
rect -1694 -181 -1660 -147
rect -1436 -181 -1402 -147
rect -1178 -181 -1144 -147
rect -920 -181 -886 -147
rect -662 -181 -628 -147
rect -404 -181 -370 -147
rect -146 -181 -112 -147
rect 112 -181 146 -147
rect 370 -181 404 -147
rect 628 -181 662 -147
rect 886 -181 920 -147
rect 1144 -181 1178 -147
rect 1402 -181 1436 -147
rect 1660 -181 1694 -147
<< locali >>
rect -1743 147 -1694 181
rect -1660 147 -1611 181
rect -1485 147 -1436 181
rect -1402 147 -1353 181
rect -1227 147 -1178 181
rect -1144 147 -1095 181
rect -969 147 -920 181
rect -886 147 -837 181
rect -711 147 -662 181
rect -628 147 -579 181
rect -453 147 -404 181
rect -370 147 -321 181
rect -195 147 -146 181
rect -112 147 -63 181
rect 63 147 112 181
rect 146 147 195 181
rect 321 147 370 181
rect 404 147 453 181
rect 579 147 628 181
rect 662 147 711 181
rect 837 147 886 181
rect 920 147 969 181
rect 1095 147 1144 181
rect 1178 147 1227 181
rect 1353 147 1402 181
rect 1436 147 1485 181
rect 1611 147 1660 181
rect 1694 147 1743 181
rect -1823 85 -1789 104
rect -1823 17 -1789 19
rect -1823 -19 -1789 -17
rect -1823 -104 -1789 -85
rect -1565 85 -1531 104
rect -1565 17 -1531 19
rect -1565 -19 -1531 -17
rect -1565 -104 -1531 -85
rect -1307 85 -1273 104
rect -1307 17 -1273 19
rect -1307 -19 -1273 -17
rect -1307 -104 -1273 -85
rect -1049 85 -1015 104
rect -1049 17 -1015 19
rect -1049 -19 -1015 -17
rect -1049 -104 -1015 -85
rect -791 85 -757 104
rect -791 17 -757 19
rect -791 -19 -757 -17
rect -791 -104 -757 -85
rect -533 85 -499 104
rect -533 17 -499 19
rect -533 -19 -499 -17
rect -533 -104 -499 -85
rect -275 85 -241 104
rect -275 17 -241 19
rect -275 -19 -241 -17
rect -275 -104 -241 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 241 85 275 104
rect 241 17 275 19
rect 241 -19 275 -17
rect 241 -104 275 -85
rect 499 85 533 104
rect 499 17 533 19
rect 499 -19 533 -17
rect 499 -104 533 -85
rect 757 85 791 104
rect 757 17 791 19
rect 757 -19 791 -17
rect 757 -104 791 -85
rect 1015 85 1049 104
rect 1015 17 1049 19
rect 1015 -19 1049 -17
rect 1015 -104 1049 -85
rect 1273 85 1307 104
rect 1273 17 1307 19
rect 1273 -19 1307 -17
rect 1273 -104 1307 -85
rect 1531 85 1565 104
rect 1531 17 1565 19
rect 1531 -19 1565 -17
rect 1531 -104 1565 -85
rect 1789 85 1823 104
rect 1789 17 1823 19
rect 1789 -19 1823 -17
rect 1789 -104 1823 -85
rect -1743 -181 -1694 -147
rect -1660 -181 -1611 -147
rect -1485 -181 -1436 -147
rect -1402 -181 -1353 -147
rect -1227 -181 -1178 -147
rect -1144 -181 -1095 -147
rect -969 -181 -920 -147
rect -886 -181 -837 -147
rect -711 -181 -662 -147
rect -628 -181 -579 -147
rect -453 -181 -404 -147
rect -370 -181 -321 -147
rect -195 -181 -146 -147
rect -112 -181 -63 -147
rect 63 -181 112 -147
rect 146 -181 195 -147
rect 321 -181 370 -147
rect 404 -181 453 -147
rect 579 -181 628 -147
rect 662 -181 711 -147
rect 837 -181 886 -147
rect 920 -181 969 -147
rect 1095 -181 1144 -147
rect 1178 -181 1227 -147
rect 1353 -181 1402 -147
rect 1436 -181 1485 -147
rect 1611 -181 1660 -147
rect 1694 -181 1743 -147
<< viali >>
rect -1694 147 -1660 181
rect -1436 147 -1402 181
rect -1178 147 -1144 181
rect -920 147 -886 181
rect -662 147 -628 181
rect -404 147 -370 181
rect -146 147 -112 181
rect 112 147 146 181
rect 370 147 404 181
rect 628 147 662 181
rect 886 147 920 181
rect 1144 147 1178 181
rect 1402 147 1436 181
rect 1660 147 1694 181
rect -1823 51 -1789 53
rect -1823 19 -1789 51
rect -1823 -51 -1789 -19
rect -1823 -53 -1789 -51
rect -1565 51 -1531 53
rect -1565 19 -1531 51
rect -1565 -51 -1531 -19
rect -1565 -53 -1531 -51
rect -1307 51 -1273 53
rect -1307 19 -1273 51
rect -1307 -51 -1273 -19
rect -1307 -53 -1273 -51
rect -1049 51 -1015 53
rect -1049 19 -1015 51
rect -1049 -51 -1015 -19
rect -1049 -53 -1015 -51
rect -791 51 -757 53
rect -791 19 -757 51
rect -791 -51 -757 -19
rect -791 -53 -757 -51
rect -533 51 -499 53
rect -533 19 -499 51
rect -533 -51 -499 -19
rect -533 -53 -499 -51
rect -275 51 -241 53
rect -275 19 -241 51
rect -275 -51 -241 -19
rect -275 -53 -241 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 241 51 275 53
rect 241 19 275 51
rect 241 -51 275 -19
rect 241 -53 275 -51
rect 499 51 533 53
rect 499 19 533 51
rect 499 -51 533 -19
rect 499 -53 533 -51
rect 757 51 791 53
rect 757 19 791 51
rect 757 -51 791 -19
rect 757 -53 791 -51
rect 1015 51 1049 53
rect 1015 19 1049 51
rect 1015 -51 1049 -19
rect 1015 -53 1049 -51
rect 1273 51 1307 53
rect 1273 19 1307 51
rect 1273 -51 1307 -19
rect 1273 -53 1307 -51
rect 1531 51 1565 53
rect 1531 19 1565 51
rect 1531 -51 1565 -19
rect 1531 -53 1565 -51
rect 1789 51 1823 53
rect 1789 19 1823 51
rect 1789 -51 1823 -19
rect 1789 -53 1823 -51
rect -1694 -181 -1660 -147
rect -1436 -181 -1402 -147
rect -1178 -181 -1144 -147
rect -920 -181 -886 -147
rect -662 -181 -628 -147
rect -404 -181 -370 -147
rect -146 -181 -112 -147
rect 112 -181 146 -147
rect 370 -181 404 -147
rect 628 -181 662 -147
rect 886 -181 920 -147
rect 1144 -181 1178 -147
rect 1402 -181 1436 -147
rect 1660 -181 1694 -147
<< metal1 >>
rect -1731 181 -1623 187
rect -1731 147 -1694 181
rect -1660 147 -1623 181
rect -1731 141 -1623 147
rect -1473 181 -1365 187
rect -1473 147 -1436 181
rect -1402 147 -1365 181
rect -1473 141 -1365 147
rect -1215 181 -1107 187
rect -1215 147 -1178 181
rect -1144 147 -1107 181
rect -1215 141 -1107 147
rect -957 181 -849 187
rect -957 147 -920 181
rect -886 147 -849 181
rect -957 141 -849 147
rect -699 181 -591 187
rect -699 147 -662 181
rect -628 147 -591 181
rect -699 141 -591 147
rect -441 181 -333 187
rect -441 147 -404 181
rect -370 147 -333 181
rect -441 141 -333 147
rect -183 181 -75 187
rect -183 147 -146 181
rect -112 147 -75 181
rect -183 141 -75 147
rect 75 181 183 187
rect 75 147 112 181
rect 146 147 183 181
rect 75 141 183 147
rect 333 181 441 187
rect 333 147 370 181
rect 404 147 441 181
rect 333 141 441 147
rect 591 181 699 187
rect 591 147 628 181
rect 662 147 699 181
rect 591 141 699 147
rect 849 181 957 187
rect 849 147 886 181
rect 920 147 957 181
rect 849 141 957 147
rect 1107 181 1215 187
rect 1107 147 1144 181
rect 1178 147 1215 181
rect 1107 141 1215 147
rect 1365 181 1473 187
rect 1365 147 1402 181
rect 1436 147 1473 181
rect 1365 141 1473 147
rect 1623 181 1731 187
rect 1623 147 1660 181
rect 1694 147 1731 181
rect 1623 141 1731 147
rect -1829 53 -1783 100
rect -1829 19 -1823 53
rect -1789 19 -1783 53
rect -1829 -19 -1783 19
rect -1829 -53 -1823 -19
rect -1789 -53 -1783 -19
rect -1829 -100 -1783 -53
rect -1571 53 -1525 100
rect -1571 19 -1565 53
rect -1531 19 -1525 53
rect -1571 -19 -1525 19
rect -1571 -53 -1565 -19
rect -1531 -53 -1525 -19
rect -1571 -100 -1525 -53
rect -1313 53 -1267 100
rect -1313 19 -1307 53
rect -1273 19 -1267 53
rect -1313 -19 -1267 19
rect -1313 -53 -1307 -19
rect -1273 -53 -1267 -19
rect -1313 -100 -1267 -53
rect -1055 53 -1009 100
rect -1055 19 -1049 53
rect -1015 19 -1009 53
rect -1055 -19 -1009 19
rect -1055 -53 -1049 -19
rect -1015 -53 -1009 -19
rect -1055 -100 -1009 -53
rect -797 53 -751 100
rect -797 19 -791 53
rect -757 19 -751 53
rect -797 -19 -751 19
rect -797 -53 -791 -19
rect -757 -53 -751 -19
rect -797 -100 -751 -53
rect -539 53 -493 100
rect -539 19 -533 53
rect -499 19 -493 53
rect -539 -19 -493 19
rect -539 -53 -533 -19
rect -499 -53 -493 -19
rect -539 -100 -493 -53
rect -281 53 -235 100
rect -281 19 -275 53
rect -241 19 -235 53
rect -281 -19 -235 19
rect -281 -53 -275 -19
rect -241 -53 -235 -19
rect -281 -100 -235 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 235 53 281 100
rect 235 19 241 53
rect 275 19 281 53
rect 235 -19 281 19
rect 235 -53 241 -19
rect 275 -53 281 -19
rect 235 -100 281 -53
rect 493 53 539 100
rect 493 19 499 53
rect 533 19 539 53
rect 493 -19 539 19
rect 493 -53 499 -19
rect 533 -53 539 -19
rect 493 -100 539 -53
rect 751 53 797 100
rect 751 19 757 53
rect 791 19 797 53
rect 751 -19 797 19
rect 751 -53 757 -19
rect 791 -53 797 -19
rect 751 -100 797 -53
rect 1009 53 1055 100
rect 1009 19 1015 53
rect 1049 19 1055 53
rect 1009 -19 1055 19
rect 1009 -53 1015 -19
rect 1049 -53 1055 -19
rect 1009 -100 1055 -53
rect 1267 53 1313 100
rect 1267 19 1273 53
rect 1307 19 1313 53
rect 1267 -19 1313 19
rect 1267 -53 1273 -19
rect 1307 -53 1313 -19
rect 1267 -100 1313 -53
rect 1525 53 1571 100
rect 1525 19 1531 53
rect 1565 19 1571 53
rect 1525 -19 1571 19
rect 1525 -53 1531 -19
rect 1565 -53 1571 -19
rect 1525 -100 1571 -53
rect 1783 53 1829 100
rect 1783 19 1789 53
rect 1823 19 1829 53
rect 1783 -19 1829 19
rect 1783 -53 1789 -19
rect 1823 -53 1829 -19
rect 1783 -100 1829 -53
rect -1731 -147 -1623 -141
rect -1731 -181 -1694 -147
rect -1660 -181 -1623 -147
rect -1731 -187 -1623 -181
rect -1473 -147 -1365 -141
rect -1473 -181 -1436 -147
rect -1402 -181 -1365 -147
rect -1473 -187 -1365 -181
rect -1215 -147 -1107 -141
rect -1215 -181 -1178 -147
rect -1144 -181 -1107 -147
rect -1215 -187 -1107 -181
rect -957 -147 -849 -141
rect -957 -181 -920 -147
rect -886 -181 -849 -147
rect -957 -187 -849 -181
rect -699 -147 -591 -141
rect -699 -181 -662 -147
rect -628 -181 -591 -147
rect -699 -187 -591 -181
rect -441 -147 -333 -141
rect -441 -181 -404 -147
rect -370 -181 -333 -147
rect -441 -187 -333 -181
rect -183 -147 -75 -141
rect -183 -181 -146 -147
rect -112 -181 -75 -147
rect -183 -187 -75 -181
rect 75 -147 183 -141
rect 75 -181 112 -147
rect 146 -181 183 -147
rect 75 -187 183 -181
rect 333 -147 441 -141
rect 333 -181 370 -147
rect 404 -181 441 -147
rect 333 -187 441 -181
rect 591 -147 699 -141
rect 591 -181 628 -147
rect 662 -181 699 -147
rect 591 -187 699 -181
rect 849 -147 957 -141
rect 849 -181 886 -147
rect 920 -181 957 -147
rect 849 -187 957 -181
rect 1107 -147 1215 -141
rect 1107 -181 1144 -147
rect 1178 -181 1215 -147
rect 1107 -187 1215 -181
rect 1365 -147 1473 -141
rect 1365 -181 1402 -147
rect 1436 -181 1473 -147
rect 1365 -187 1473 -181
rect 1623 -147 1731 -141
rect 1623 -181 1660 -147
rect 1694 -181 1731 -147
rect 1623 -187 1731 -181
<< end >>
