magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< locali >>
rect 2583 1443 3160 1477
rect 174 1372 1662 1406
rect 94 1264 1662 1298
rect 1156 1072 1662 1106
rect 1396 964 1662 998
rect 2583 893 3160 927
rect 2583 653 3160 687
rect 174 603 414 637
rect 1236 582 1662 616
rect 1316 474 1662 508
rect 1156 282 1662 316
rect 94 153 414 187
rect 1236 174 1662 208
rect 2583 103 3160 137
<< metal1 >>
rect 80 199 108 1500
rect 160 649 188 1500
rect 151 591 197 649
rect 71 141 117 199
rect 80 80 108 141
rect 160 80 188 591
rect 504 80 532 790
rect 900 80 928 790
rect 1030 644 1094 696
rect 1030 94 1094 146
rect 1142 80 1170 1500
rect 1222 80 1250 1500
rect 1302 80 1330 1500
rect 1382 80 1410 1500
rect 1788 80 1836 1610
rect 2212 80 2262 1612
rect 2602 80 2630 1580
rect 2998 80 3026 1580
<< metal2 >>
rect 1784 1168 1840 1216
rect 2209 1168 2265 1216
rect 2588 1161 2644 1209
rect 2984 1161 3040 1209
rect 1048 692 1236 720
rect 1048 670 1076 692
rect 490 371 546 419
rect 886 371 942 419
rect 1784 378 1840 426
rect 2209 378 2265 426
rect 2588 371 2644 419
rect 2984 371 3040 419
rect 1048 297 1156 325
rect 1048 120 1076 297
<< metal3 >>
rect 1763 1143 1861 1241
rect 2188 1143 2286 1241
rect 2567 1136 2665 1234
rect 2963 1136 3061 1234
rect 469 346 567 444
rect 865 346 963 444
rect 1763 353 1861 451
rect 2188 353 2286 451
rect 2567 346 2665 444
rect 2963 346 3061 444
use contact_16  contact_16_9
timestamp 1624494425
transform 1 0 61 0 1 141
box 0 0 66 58
use contact_8  contact_8_4
timestamp 1624494425
transform 1 0 486 0 1 363
box 0 0 64 64
use contact_9  contact_9_4
timestamp 1624494425
transform 1 0 485 0 1 358
box 0 0 66 74
use pinv_dec  pinv_dec_0
timestamp 1624494425
transform 1 0 320 0 -1 790
box 44 0 760 490
use pinv_dec  pinv_dec_1
timestamp 1624494425
transform 1 0 320 0 1 0
box 44 0 760 490
use contact_7  contact_7_5
timestamp 1624494425
transform 1 0 1033 0 1 87
box 0 0 58 66
use contact_8  contact_8_11
timestamp 1624494425
transform 1 0 1030 0 1 88
box 0 0 64 64
use contact_17  contact_17_1
timestamp 1624494425
transform 1 0 1124 0 1 279
box 0 0 64 64
use contact_16  contact_16_7
timestamp 1624494425
transform 1 0 1123 0 1 270
box 0 0 66 58
use contact_16  contact_16_6
timestamp 1624494425
transform 1 0 1203 0 1 162
box 0 0 66 58
use contact_16  contact_16_5
timestamp 1624494425
transform 1 0 1283 0 1 462
box 0 0 66 58
use contact_8  contact_8_9
timestamp 1624494425
transform 1 0 882 0 1 363
box 0 0 64 64
use contact_9  contact_9_9
timestamp 1624494425
transform 1 0 881 0 1 358
box 0 0 66 74
use contact_9  contact_9_2
timestamp 1624494425
transform 1 0 1779 0 1 365
box 0 0 66 74
use contact_8  contact_8_2
timestamp 1624494425
transform 1 0 1780 0 1 370
box 0 0 64 64
use contact_9  contact_9_3
timestamp 1624494425
transform 1 0 2583 0 1 358
box 0 0 66 74
use contact_8  contact_8_3
timestamp 1624494425
transform 1 0 2584 0 1 363
box 0 0 64 64
use contact_9  contact_9_7
timestamp 1624494425
transform 1 0 2979 0 1 358
box 0 0 66 74
use contact_8  contact_8_7
timestamp 1624494425
transform 1 0 2980 0 1 363
box 0 0 64 64
use contact_9  contact_9_8
timestamp 1624494425
transform 1 0 2204 0 1 365
box 0 0 66 74
use contact_8  contact_8_8
timestamp 1624494425
transform 1 0 2205 0 1 370
box 0 0 64 64
use and2_dec  and2_dec_3
timestamp 1624494425
transform 1 0 1542 0 1 0
box 70 -56 1636 490
use and2_dec  and2_dec_2
timestamp 1624494425
transform 1 0 1542 0 -1 790
box 70 -56 1636 490
use contact_16  contact_16_8
timestamp 1624494425
transform 1 0 141 0 1 591
box 0 0 66 58
use contact_7  contact_7_4
timestamp 1624494425
transform 1 0 1033 0 1 637
box 0 0 58 66
use contact_8  contact_8_10
timestamp 1624494425
transform 1 0 1030 0 1 638
box 0 0 64 64
use contact_17  contact_17_0
timestamp 1624494425
transform 1 0 1204 0 1 674
box 0 0 64 64
use contact_16  contact_16_4
timestamp 1624494425
transform 1 0 1203 0 1 570
box 0 0 66 58
use contact_16  contact_16_2
timestamp 1624494425
transform 1 0 1363 0 1 952
box 0 0 66 58
use and2_dec  and2_dec_1
timestamp 1624494425
transform 1 0 1542 0 1 790
box 70 -56 1636 490
use contact_7  contact_7_3
timestamp 1624494425
transform 1 0 65 0 1 1248
box 0 0 58 66
use contact_7  contact_7_2
timestamp 1624494425
transform 1 0 1287 0 1 1248
box 0 0 58 66
use contact_16  contact_16_3
timestamp 1624494425
transform 1 0 1123 0 1 1060
box 0 0 66 58
use contact_16  contact_16_1
timestamp 1624494425
transform 1 0 1283 0 1 1252
box 0 0 66 58
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 1780 0 1 1160
box 0 0 64 64
use contact_9  contact_9_0
timestamp 1624494425
transform 1 0 1779 0 1 1155
box 0 0 66 74
use contact_8  contact_8_6
timestamp 1624494425
transform 1 0 2205 0 1 1160
box 0 0 64 64
use contact_9  contact_9_6
timestamp 1624494425
transform 1 0 2204 0 1 1155
box 0 0 66 74
use contact_8  contact_8_1
timestamp 1624494425
transform 1 0 2584 0 1 1153
box 0 0 64 64
use contact_9  contact_9_1
timestamp 1624494425
transform 1 0 2583 0 1 1148
box 0 0 66 74
use contact_8  contact_8_5
timestamp 1624494425
transform 1 0 2980 0 1 1153
box 0 0 64 64
use contact_9  contact_9_5
timestamp 1624494425
transform 1 0 2979 0 1 1148
box 0 0 66 74
use contact_16  contact_16_0
timestamp 1624494425
transform 1 0 1363 0 1 1360
box 0 0 66 58
use contact_7  contact_7_0
timestamp 1624494425
transform 1 0 1367 0 1 1356
box 0 0 58 66
use contact_7  contact_7_1
timestamp 1624494425
transform 1 0 145 0 1 1356
box 0 0 58 66
use and2_dec  and2_dec_0
timestamp 1624494425
transform 1 0 1542 0 -1 1580
box 70 -56 1636 490
<< labels >>
rlabel metal1 s 71 141 117 199 4 in_0
rlabel metal1 s 151 591 197 649 4 in_1
rlabel locali s 2871 120 2871 120 4 out_0
rlabel locali s 2871 670 2871 670 4 out_1
rlabel locali s 2871 910 2871 910 4 out_2
rlabel locali s 2871 1460 2871 1460 4 out_3
rlabel metal3 s 2963 346 3061 444 4 vdd
rlabel metal3 s 2188 1143 2286 1241 4 vdd
rlabel metal3 s 2188 353 2286 451 4 vdd
rlabel metal3 s 2963 1136 3061 1234 4 vdd
rlabel metal3 s 865 346 963 444 4 vdd
rlabel metal3 s 2567 346 2665 444 4 gnd
rlabel metal3 s 1763 1143 1861 1241 4 gnd
rlabel metal3 s 2567 1136 2665 1234 4 gnd
rlabel metal3 s 469 346 567 444 4 gnd
rlabel metal3 s 1763 353 1861 451 4 gnd
<< properties >>
string FIXED_BBOX 0 0 3160 1580
<< end >>
