magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< nwell >>
rect 36584 12390 38738 14006
<< nsubdiff >>
rect 36718 13870 36880 13970
rect 38520 13870 38682 13970
rect 36718 13808 36818 13870
rect 36718 12526 36818 12588
rect 38582 13808 38682 13870
rect 38582 12526 38682 12588
rect 36718 12426 36880 12526
rect 38520 12426 38682 12526
<< nsubdiffcont >>
rect 36880 13870 38520 13970
rect 36718 12588 36818 13808
rect 38582 12588 38682 13808
rect 36880 12426 38520 12526
<< locali >>
rect 36718 13808 36818 13970
rect 36718 12426 36818 12588
rect 38582 13808 38682 13970
rect 38582 12426 38682 12588
<< viali >>
rect 36818 13870 36880 13970
rect 36880 13870 38520 13970
rect 38520 13870 38582 13970
rect 36718 12593 36818 13803
rect 38582 12593 38682 13803
rect 36818 12426 36880 12526
rect 36880 12426 38520 12526
rect 38520 12426 38582 12526
rect -1114 362 -914 396
rect -1188 -100 -1154 360
rect -872 -96 -836 358
rect -1116 -136 -916 -102
<< metal1 >>
rect 15638 17112 15698 17220
rect 13280 17050 13286 17110
rect 13346 17050 13352 17110
rect 15638 17046 15698 17052
rect 12484 16464 12490 16524
rect 12550 16464 13584 16524
rect 15632 16462 15638 16522
rect 15698 16462 15704 16522
rect -3432 14300 -1262 14548
rect -3432 13782 -2276 14300
rect -1748 13782 -1262 14300
rect -3432 13306 -1262 13782
rect -3432 1924 -3342 13306
rect -2908 1924 -1262 13306
rect 36712 13970 38688 13976
rect 36712 13870 36818 13970
rect 38582 13870 38688 13970
rect 36712 13864 38688 13870
rect 36712 13803 36824 13864
rect 36712 12593 36718 13803
rect 36818 12593 36824 13803
rect 37424 13564 37434 13864
rect 37966 13564 37976 13864
rect 38576 13803 38688 13864
rect 36890 13396 38514 13426
rect 36890 13300 36928 13396
rect 38480 13300 38514 13396
rect 36890 13272 38514 13300
rect 36900 13130 37084 13272
rect 36900 12658 36960 13130
rect 37024 13044 37084 13130
rect 37414 12936 37474 13272
rect 37666 13134 37672 13194
rect 37732 13134 37738 13194
rect 37028 12658 37088 12753
rect 37156 12660 37216 12876
rect 37284 12662 37344 12748
rect 37540 12662 37600 12752
rect 37672 12662 37732 13134
rect 37930 12938 37990 13272
rect 38316 13135 38502 13272
rect 38316 13044 38376 13135
rect 37802 12662 37862 12750
rect 38058 12662 38118 12752
rect 36900 12598 37088 12658
rect 37150 12600 37156 12660
rect 37216 12600 37222 12660
rect 37284 12602 38118 12662
rect 38186 12660 38246 12844
rect 38314 12660 38374 12752
rect 38442 12660 38502 13135
rect 38180 12600 38186 12660
rect 38246 12600 38252 12660
rect 38314 12600 38502 12660
rect 36712 12532 36824 12593
rect 38576 12593 38582 13803
rect 38682 12593 38688 13803
rect 38576 12532 38688 12593
rect 36712 12526 38688 12532
rect 36712 12426 36818 12526
rect 38582 12426 38688 12526
rect 36712 12420 38688 12426
rect 12492 12066 12552 12072
rect 13280 12006 13286 12066
rect 13346 12006 13352 12066
rect 12492 12000 12552 12006
rect 12492 9974 12552 9980
rect 12492 9908 12552 9914
rect 12492 8732 12552 8738
rect 12492 8666 12552 8672
rect 12492 7496 12552 7502
rect 12492 7430 12552 7436
rect 13290 6970 13350 6976
rect 12486 6910 12492 6970
rect 12552 6910 12558 6970
rect 13290 6904 13350 6910
rect 13282 5326 13288 5386
rect 13348 5326 13354 5386
rect 41288 5252 41348 5402
rect 41288 5186 41348 5192
rect 11882 4670 11888 4730
rect 11948 4670 11954 4730
rect 13280 4670 13286 4730
rect 13346 4670 13352 4730
rect -3432 1842 -1262 1924
rect 8212 1394 8424 1454
rect 47814 1394 48076 1454
rect -1266 396 -810 414
rect -1266 394 -1114 396
rect -1364 362 -1114 394
rect -914 362 -810 396
rect -1364 360 -810 362
rect -1364 -76 -1188 360
rect -1154 358 -810 360
rect -1154 344 -872 358
rect -1154 164 -1132 344
rect -1052 232 -1046 292
rect -986 232 -980 292
rect -998 166 -938 172
rect -1154 104 -1040 164
rect -1004 106 -998 166
rect -938 106 -932 166
rect -1154 -68 -1132 104
rect -998 100 -938 106
rect -1052 -18 -1046 42
rect -986 -18 -980 42
rect -894 -68 -872 344
rect -1154 -76 -872 -68
rect -836 -68 -810 358
rect -836 -76 -808 -68
rect -1364 -120 -1198 -76
rect -1266 -142 -1198 -120
rect -814 -142 -808 -76
rect -1266 -152 -808 -142
rect -1266 -154 -1140 -152
rect -894 -154 -810 -152
<< via1 >>
rect 13286 17050 13346 17110
rect 15638 17052 15698 17112
rect 12490 16464 12550 16524
rect 15638 16462 15698 16522
rect -2276 13782 -1748 14300
rect -3342 1924 -2908 13306
rect 36824 13564 37424 13864
rect 37976 13564 38576 13864
rect 36928 13300 38480 13396
rect 37672 13134 37732 13194
rect 37156 12600 37216 12660
rect 38186 12600 38246 12660
rect 12492 12006 12552 12066
rect 13286 12006 13346 12066
rect 12492 9914 12552 9974
rect 12492 8672 12552 8732
rect 12492 7436 12552 7496
rect 12492 6910 12552 6970
rect 13290 6910 13350 6970
rect 13288 5326 13348 5386
rect 41288 5192 41348 5252
rect 11888 4670 11948 4730
rect 13286 4670 13346 4730
rect -1046 232 -986 292
rect -998 106 -938 166
rect -1046 -18 -986 42
rect -1198 -100 -1188 -76
rect -1188 -100 -1154 -76
rect -1154 -96 -872 -76
rect -872 -96 -836 -76
rect -836 -96 -814 -76
rect -1154 -100 -814 -96
rect -1198 -102 -814 -100
rect -1198 -136 -1116 -102
rect -1116 -136 -916 -102
rect -916 -136 -814 -102
rect -1198 -142 -814 -136
<< metal2 >>
rect 13286 17110 13346 17116
rect 15632 17052 15638 17112
rect 15698 17052 15704 17112
rect 12490 16524 12550 16530
rect 12490 16458 12550 16464
rect 13286 16400 13346 17050
rect 15638 16522 15698 17052
rect 15638 16456 15698 16462
rect 12492 15404 12552 15426
rect 12492 15236 12552 15344
rect -3432 14300 -1262 14548
rect -3432 13782 -2276 14300
rect -1748 13782 -1262 14300
rect -3432 13306 -1262 13782
rect 36824 13864 37424 13874
rect 36824 13554 37424 13564
rect 37976 13864 38576 13874
rect 37976 13554 38576 13564
rect -3432 1924 -3342 13306
rect -2908 1924 -1262 13306
rect 36890 13396 38514 13426
rect 36890 13300 36928 13396
rect 38480 13300 38514 13396
rect 36890 13272 38514 13300
rect 37672 13194 37732 13200
rect 39132 13194 39192 13203
rect 37732 13134 39132 13194
rect 37672 13128 37732 13134
rect 39132 13125 39192 13134
rect 37136 12660 37236 12678
rect 38186 12660 38246 12666
rect 37136 12600 37156 12660
rect 37216 12600 38186 12660
rect 13286 12066 13346 12072
rect 12486 12006 12492 12066
rect 12552 12006 13286 12066
rect 13286 12000 13346 12006
rect 12486 9914 12492 9974
rect 12552 9914 13458 9974
rect 34372 9914 34708 9974
rect 34768 9914 34777 9974
rect 12486 8672 12492 8732
rect 12552 8672 13658 8732
rect 12486 7436 12492 7496
rect 12552 7436 13602 7496
rect 12492 6970 12552 6976
rect 12552 6910 13290 6970
rect 13350 6910 13356 6970
rect 12492 6904 12552 6910
rect 13288 5386 13348 5392
rect 12342 5326 13288 5386
rect 13288 5320 13348 5326
rect 33930 5192 34110 5252
rect 34170 5192 34179 5252
rect 11888 4730 11948 4736
rect 13286 4730 13346 4736
rect 11948 4670 13286 4730
rect 11888 4664 11948 4670
rect 13286 4664 13346 4670
rect 11886 2776 11946 2954
rect 11886 2716 13454 2776
rect -3432 1842 -1262 1924
rect 264 1913 273 2003
rect 363 1913 372 2003
rect -1046 292 -986 298
rect -986 232 -694 292
rect 37136 254 37236 12600
rect 38186 12594 38246 12600
rect 41279 6288 41288 6348
rect 41348 6288 41444 6348
rect 41288 5252 41348 5261
rect 41282 5192 41288 5252
rect 41348 5192 41354 5252
rect 41288 5183 41348 5192
rect 52714 2892 53274 2952
rect -1046 226 -986 232
rect -1012 168 -922 180
rect -1012 104 -1000 168
rect -934 104 -922 168
rect -1012 94 -922 104
rect -1046 42 -986 48
rect -834 42 -774 232
rect 37127 154 37136 254
rect 37236 154 37245 254
rect -986 -18 -774 42
rect -1046 -24 -986 -18
rect -1212 -76 -806 -64
rect -1212 -142 -1198 -76
rect -814 -142 -806 -76
rect -1212 -154 -806 -142
<< via2 >>
rect 12492 15344 12552 15404
rect -2276 13782 -1748 14300
rect 36824 13564 37424 13864
rect 37976 13564 38576 13864
rect -3342 1924 -2908 13306
rect 36928 13300 38480 13396
rect 39132 13134 39192 13194
rect 34708 9914 34768 9974
rect 34110 5192 34170 5252
rect 273 1913 363 2003
rect 41288 6288 41348 6348
rect 41288 5192 41348 5252
rect -1000 166 -934 168
rect -1000 106 -998 166
rect -998 106 -938 166
rect -938 106 -934 166
rect -1000 104 -934 106
rect 37136 154 37236 254
rect -1198 -142 -814 -76
<< metal3 >>
rect 12430 15424 12624 15426
rect 12430 15409 12636 15424
rect 12430 15345 12487 15409
rect 12557 15345 12636 15409
rect 12430 15344 12492 15345
rect 12552 15344 12636 15345
rect 12430 15328 12636 15344
rect 12430 15324 12624 15328
rect -3634 14544 -2794 14660
rect -16568 14398 -1528 14544
rect -16568 14388 -2374 14398
rect -16568 13698 -16416 14388
rect -15720 13700 -2374 14388
rect -1684 13700 -1528 14398
rect 52113 14346 52211 14351
rect 39110 14345 52212 14346
rect 39110 14247 52113 14345
rect 52211 14247 52212 14345
rect 39110 14246 52212 14247
rect -15720 13698 -1528 13700
rect -16568 13306 -1528 13698
rect 36814 13864 37434 13869
rect 36814 13564 36824 13864
rect 37424 13564 37434 13864
rect 36814 13559 37434 13564
rect 37966 13864 38586 13869
rect 37966 13564 37976 13864
rect 38576 13564 38586 13864
rect 37966 13559 38586 13564
rect -16568 1924 -3342 13306
rect -2908 1924 -1528 13306
rect 36890 13396 38514 13426
rect 36890 13300 36928 13396
rect 38480 13300 38514 13396
rect 36890 13272 38514 13300
rect 39110 13194 39210 14246
rect 52113 14241 52211 14246
rect 39110 13134 39132 13194
rect 39192 13134 39210 13194
rect 39110 13114 39210 13134
rect 34688 9974 41370 9992
rect 34688 9914 34708 9974
rect 34768 9914 41370 9974
rect 34688 9892 41370 9914
rect 41270 6348 41370 9892
rect 41270 6288 41288 6348
rect 41348 6288 41370 6348
rect 41270 6270 41370 6288
rect 34086 5252 41380 5270
rect 34086 5192 34110 5252
rect 34170 5192 41288 5252
rect 41348 5192 41380 5252
rect 34086 5170 41380 5192
rect -16568 360 -1528 1924
rect 268 2003 368 2008
rect 268 1913 273 2003
rect 363 1913 368 2003
rect 268 634 368 1913
rect -1016 514 -916 520
rect 268 513 370 634
rect 263 415 269 513
rect 367 415 373 513
rect 268 414 370 415
rect -16568 -458 -2656 360
rect -1016 168 -916 414
rect -1016 104 -1000 168
rect -934 104 -916 168
rect 270 254 370 414
rect 37131 254 37241 259
rect 270 154 37136 254
rect 37236 154 37241 254
rect 37131 149 37241 154
rect -1016 94 -916 104
rect -1212 -76 -806 -64
rect -1212 -142 -1198 -76
rect -814 -142 -806 -76
rect -1212 -154 -806 -142
<< via3 >>
rect 12487 15404 12557 15409
rect 12487 15345 12492 15404
rect 12492 15345 12552 15404
rect 12552 15345 12557 15404
rect -16416 13698 -15720 14388
rect -2374 14300 -1684 14398
rect -2374 13782 -2276 14300
rect -2276 13782 -1748 14300
rect -1748 13782 -1684 14300
rect -2374 13700 -1684 13782
rect 52113 14247 52211 14345
rect 36824 13564 37424 13864
rect 37976 13564 38576 13864
rect 36928 13300 38480 13396
rect -1016 414 -916 514
rect 269 415 367 513
rect -1198 -142 -814 -76
<< mimcap >>
rect -15382 14294 -9182 14344
rect -15382 13994 -9532 14294
rect -9232 13994 -9182 14294
rect -15382 13944 -9182 13994
rect -8982 14294 -2782 14344
rect -8982 13994 -3132 14294
rect -2832 13994 -2782 14294
rect -8982 13944 -2782 13994
rect -16468 13312 -15668 13362
rect -16468 7612 -16018 13312
rect -15718 7612 -15668 13312
rect -2424 13312 -1624 13362
rect -14528 12394 -9328 12444
rect -14528 7694 -9678 12394
rect -9378 7694 -9328 12394
rect -14528 7644 -9328 7694
rect -8928 12394 -3728 12444
rect -8928 7694 -4078 12394
rect -3778 7694 -3728 12394
rect -8928 7644 -3728 7694
rect -16468 7562 -15668 7612
rect -2424 7612 -1974 13312
rect -1674 7612 -1624 13312
rect -2424 7562 -1624 7612
rect -16468 6820 -15668 6870
rect -16468 1120 -16018 6820
rect -15718 1120 -15668 6820
rect -14528 6794 -9328 6844
rect -14528 2094 -9678 6794
rect -9378 2094 -9328 6794
rect -14528 2044 -9328 2094
rect -8928 6794 -3728 6844
rect -8928 2094 -4078 6794
rect -3778 2094 -3728 6794
rect -8928 2044 -3728 2094
rect -2424 6820 -1624 6870
rect -16468 1070 -15668 1120
rect -2424 1120 -1974 6820
rect -1674 1120 -1624 6820
rect -2424 1070 -1624 1120
rect -15882 394 -9682 444
rect -15882 94 -10032 394
rect -9732 94 -9682 394
rect -15882 44 -9682 94
rect -9482 394 -3282 444
rect -9482 94 -3632 394
rect -3332 94 -3282 394
rect -9482 44 -3282 94
<< mimcapcontact >>
rect -9532 13994 -9232 14294
rect -3132 13994 -2832 14294
rect -16018 7612 -15718 13312
rect -9678 7694 -9378 12394
rect -4078 7694 -3778 12394
rect -1974 7612 -1674 13312
rect -16018 1120 -15718 6820
rect -9678 2094 -9378 6794
rect -4078 2094 -3778 6794
rect -1974 1120 -1674 6820
rect -10032 94 -9732 394
rect -3632 94 -3332 394
<< metal4 >>
rect 34964 29970 35232 30770
rect 36032 29970 37598 30770
rect 12486 15409 12558 15410
rect 12486 15345 12487 15409
rect 12557 15345 12558 15409
rect 12486 15344 12558 15345
rect -4196 14544 -1528 14984
rect -16568 14398 -1528 14544
rect -16568 14388 -2374 14398
rect -16568 13698 -16416 14388
rect -15720 14294 -2374 14388
rect -15720 13994 -9532 14294
rect -9232 13994 -3132 14294
rect -2832 13994 -2374 14294
rect -15720 13700 -2374 13994
rect -1684 13700 -1528 14398
rect 52112 14345 52212 15426
rect 52112 14247 52113 14345
rect 52211 14247 52212 14345
rect 52112 14246 52212 14247
rect 35516 14048 36670 14050
rect -15720 13698 -1528 13700
rect -16568 13368 -1528 13698
rect -16568 13312 -15386 13368
rect -16568 7612 -16018 13312
rect -15718 7612 -15386 13312
rect -2828 13312 -1528 13368
rect -16568 6820 -15386 7612
rect -16568 1120 -16018 6820
rect -15718 1120 -15386 6820
rect -14628 12394 -3628 12544
rect -14628 7694 -9678 12394
rect -9378 7694 -4078 12394
rect -3778 7694 -3628 12394
rect -14628 6794 -3628 7694
rect -14628 2094 -9678 6794
rect -9378 2094 -4078 6794
rect -3778 2094 -3628 6794
rect -14628 1544 -3628 2094
rect -2828 7612 -1974 13312
rect -1674 7612 -1528 13312
rect 35232 14028 38760 14048
rect 35232 13276 35256 14028
rect 36008 13864 38760 14028
rect 36008 13564 36824 13864
rect 37424 13564 37976 13864
rect 38576 13564 38760 13864
rect 36008 13396 38760 13564
rect 36008 13300 36928 13396
rect 38480 13300 38760 13396
rect 36008 13276 38760 13300
rect 35232 13248 38760 13276
rect -2828 6820 -1528 7612
rect -2828 1760 -1974 6820
rect -3754 1496 -3628 1544
rect -3754 1396 -2814 1496
rect -16568 706 -15386 1120
rect -16568 620 -3244 706
rect -16566 394 -3244 620
rect -16566 94 -10032 394
rect -9732 94 -3632 394
rect -3332 94 -3244 394
rect -2914 340 -2814 1396
rect -2458 1120 -1974 1760
rect -1674 1120 -1528 6820
rect -2458 1002 -1528 1120
rect -2458 610 -1952 1002
rect -1017 514 -915 515
rect -1400 414 -1016 514
rect -916 513 368 514
rect -916 415 269 513
rect 367 415 368 513
rect -916 414 368 415
rect -1400 340 -1300 414
rect -1017 413 -915 414
rect -2914 240 -1300 340
rect -16566 38 -3244 94
rect -16566 -358 -16436 38
rect -16034 -32 -3244 38
rect -2652 -32 -1544 -30
rect -16034 -88 -1544 -32
rect -16034 -358 -2058 -88
rect -16566 -426 -2058 -358
rect -1690 -426 -1544 -88
rect -16566 -830 -1544 -426
rect 33872 -830 38596 -30
<< via4 >>
rect 35232 29970 36032 30770
rect -16416 13698 -15720 14388
rect -2374 13700 -1684 14398
rect 35256 13276 36008 14028
rect -16436 -358 -16034 38
rect -2058 -426 -1690 -88
<< mimcap2 >>
rect -15382 13894 -9582 14344
rect -15382 13594 -15332 13894
rect -9632 13594 -9582 13894
rect -15382 13544 -9582 13594
rect -8982 13894 -3182 14344
rect -8982 13594 -8932 13894
rect -3232 13594 -3182 13894
rect -8982 13544 -3182 13594
rect -16468 7512 -16068 13362
rect -16468 7212 -16418 7512
rect -16118 7212 -16068 7512
rect -14528 7594 -9728 12444
rect -14528 7294 -14478 7594
rect -9778 7294 -9728 7594
rect -14528 7244 -9728 7294
rect -8928 7594 -4128 12444
rect -8928 7294 -8878 7594
rect -4178 7294 -4128 7594
rect -8928 7244 -4128 7294
rect -2424 7512 -2024 13362
rect -16468 7162 -16068 7212
rect -2424 7212 -2374 7512
rect -2074 7212 -2024 7512
rect -2424 7162 -2024 7212
rect -16468 1020 -16068 6870
rect -14528 1994 -9728 6844
rect -14528 1694 -14478 1994
rect -9778 1694 -9728 1994
rect -14528 1644 -9728 1694
rect -8928 1994 -4128 6844
rect -8928 1694 -8878 1994
rect -4178 1694 -4128 1994
rect -8928 1644 -4128 1694
rect -16468 720 -16418 1020
rect -16118 720 -16068 1020
rect -16468 670 -16068 720
rect -2424 1020 -2024 6870
rect -2424 720 -2374 1020
rect -2074 720 -2024 1020
rect -2424 670 -2024 720
rect -15882 -6 -10082 444
rect -15882 -306 -15832 -6
rect -10132 -306 -10082 -6
rect -15882 -356 -10082 -306
rect -9482 -6 -3682 444
rect -9482 -306 -9432 -6
rect -3732 -306 -3682 -6
rect -9482 -356 -3682 -306
<< mimcap2contact >>
rect -15332 13594 -9632 13894
rect -8932 13594 -3232 13894
rect -16418 7212 -16118 7512
rect -14478 7294 -9778 7594
rect -8878 7294 -4178 7594
rect -2374 7212 -2074 7512
rect -14478 1694 -9778 1994
rect -8878 1694 -4178 1994
rect -16418 720 -16118 1020
rect -2374 720 -2074 1020
rect -15832 -306 -10132 -6
rect -9432 -306 -3732 -6
<< metal5 >>
rect 35208 30770 36056 30794
rect 35208 29970 35232 30770
rect 36032 29970 36056 30770
rect 35208 29946 36056 29970
rect -16568 14398 -1528 14544
rect -16568 14388 -2374 14398
rect -16568 13698 -16416 14388
rect -15720 13894 -2374 14388
rect -15720 13698 -15332 13894
rect -16568 13594 -15332 13698
rect -9632 13594 -8932 13894
rect -3232 13700 -2374 13894
rect -1684 13700 -1528 14398
rect -3232 13594 -1528 13700
rect -16568 13368 -1528 13594
rect -16568 7594 -3364 13368
rect -16568 7512 -14478 7594
rect -16568 7212 -16418 7512
rect -16118 7294 -14478 7512
rect -9778 7294 -8878 7594
rect -4178 7294 -3364 7594
rect -16118 7212 -3364 7294
rect -16568 1994 -3364 7212
rect -16568 1694 -14478 1994
rect -9778 1694 -8878 1994
rect -4178 1844 -3364 1994
rect -2828 7512 -1528 13368
rect 35232 14028 36032 29946
rect 35232 13276 35256 14028
rect 36008 13276 36032 14028
rect 35232 13252 36032 13276
rect -2828 7212 -2374 7512
rect -2074 7212 -1528 7512
rect -2828 1844 -1528 7212
rect -4178 1694 -1528 1844
rect -16568 1020 -1528 1694
rect -16568 720 -16418 1020
rect -16118 720 -2374 1020
rect -2074 720 -1528 1020
rect -16568 360 -1528 720
rect -16568 38 -1530 360
rect -16568 -358 -16436 38
rect -16034 -6 -1530 38
rect -16034 -306 -15832 -6
rect -10132 -306 -9432 -6
rect -3732 -88 -1530 -6
rect -3732 -306 -2058 -88
rect -16034 -358 -2058 -306
rect -16568 -426 -2058 -358
rect -1690 -426 -1530 -88
rect -16568 -458 -1530 -426
use sky130_fd_pr__nfet_01v8_HFLVLW  sky130_fd_pr__nfet_01v8_HFLVLW_0
timestamp 1624477805
transform 1 0 -1013 0 1 137
box -211 -279 211 275
use sky130_fd_pr__pfet_01v8_RC2RSP  sky130_fd_pr__pfet_01v8_RC2RSP_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/continuous_time_comparator
timestamp 1624477805
transform 1 0 37701 0 1 12898
box -839 -200 839 200
use se_fold_casc_wide_swing_ota  se_fold_casc_wide_swing_ota_1 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/se_fold_casc_wide_swing_ota
timestamp 1624477805
transform 1 0 51950 0 1 26370
box -15168 -27258 25000 4400
use se_fold_casc_wide_swing_ota  se_fold_casc_wide_swing_ota_0
timestamp 1624477805
transform 1 0 10950 0 1 26370
box -15168 -27258 25000 4400
<< labels >>
flabel metal2 38146 12624 38158 12636 1 FreeSans 480 0 0 0 vpeakh
flabel metal1 37310 12672 37326 12682 1 FreeSans 480 0 0 0 verr
flabel metal4 37536 14028 37548 14038 1 FreeSans 480 0 0 0 VDD
flabel metal2 -742 256 -736 264 1 FreeSans 480 0 0 0 rst
flabel metal2 53200 2918 53216 2930 1 FreeSans 480 0 0 0 vin
flabel metal2 12516 15272 12528 15284 1 FreeSans 480 0 0 0 vpeak_out
flabel metal4 36274 -344 36322 -292 1 FreeSans 480 0 0 0 VSS
flabel metal1 8324 1414 8342 1424 1 FreeSans 480 0 0 0 ibiasn2
flabel metal1 47952 1414 47972 1428 1 FreeSans 480 0 0 0 ibiasn1
flabel metal4 -1544 284 -1530 294 1 FreeSans 480 0 0 0 vpeak
<< properties >>
string FIXED_BBOX 648 33828 2512 35272
<< end >>
