magic
tech sky130A
magscale 1 2
timestamp 1620353837
<< nmoslvt >>
rect -1610 -300 -1370 300
rect -1312 -300 -1072 300
rect -1014 -300 -774 300
rect -716 -300 -476 300
rect -418 -300 -178 300
rect -120 -300 120 300
rect 178 -300 418 300
rect 476 -300 716 300
rect 774 -300 1014 300
rect 1072 -300 1312 300
rect 1370 -300 1610 300
<< ndiff >>
rect -1668 288 -1610 300
rect -1668 -288 -1656 288
rect -1622 -288 -1610 288
rect -1668 -300 -1610 -288
rect -1370 288 -1312 300
rect -1370 -288 -1358 288
rect -1324 -288 -1312 288
rect -1370 -300 -1312 -288
rect -1072 288 -1014 300
rect -1072 -288 -1060 288
rect -1026 -288 -1014 288
rect -1072 -300 -1014 -288
rect -774 288 -716 300
rect -774 -288 -762 288
rect -728 -288 -716 288
rect -774 -300 -716 -288
rect -476 288 -418 300
rect -476 -288 -464 288
rect -430 -288 -418 288
rect -476 -300 -418 -288
rect -178 288 -120 300
rect -178 -288 -166 288
rect -132 -288 -120 288
rect -178 -300 -120 -288
rect 120 288 178 300
rect 120 -288 132 288
rect 166 -288 178 288
rect 120 -300 178 -288
rect 418 288 476 300
rect 418 -288 430 288
rect 464 -288 476 288
rect 418 -300 476 -288
rect 716 288 774 300
rect 716 -288 728 288
rect 762 -288 774 288
rect 716 -300 774 -288
rect 1014 288 1072 300
rect 1014 -288 1026 288
rect 1060 -288 1072 288
rect 1014 -300 1072 -288
rect 1312 288 1370 300
rect 1312 -288 1324 288
rect 1358 -288 1370 288
rect 1312 -300 1370 -288
rect 1610 288 1668 300
rect 1610 -288 1622 288
rect 1656 -288 1668 288
rect 1610 -300 1668 -288
<< ndiffc >>
rect -1656 -288 -1622 288
rect -1358 -288 -1324 288
rect -1060 -288 -1026 288
rect -762 -288 -728 288
rect -464 -288 -430 288
rect -166 -288 -132 288
rect 132 -288 166 288
rect 430 -288 464 288
rect 728 -288 762 288
rect 1026 -288 1060 288
rect 1324 -288 1358 288
rect 1622 -288 1656 288
<< poly >>
rect -1568 372 -1412 388
rect -1568 355 -1552 372
rect -1610 338 -1552 355
rect -1428 355 -1412 372
rect -1270 372 -1114 388
rect -1270 355 -1254 372
rect -1428 338 -1370 355
rect -1610 300 -1370 338
rect -1312 338 -1254 355
rect -1130 355 -1114 372
rect -972 372 -816 388
rect -972 355 -956 372
rect -1130 338 -1072 355
rect -1312 300 -1072 338
rect -1014 338 -956 355
rect -832 355 -816 372
rect -674 372 -518 388
rect -674 355 -658 372
rect -832 338 -774 355
rect -1014 300 -774 338
rect -716 338 -658 355
rect -534 355 -518 372
rect -376 372 -220 388
rect -376 355 -360 372
rect -534 338 -476 355
rect -716 300 -476 338
rect -418 338 -360 355
rect -236 355 -220 372
rect -78 372 78 388
rect -78 355 -62 372
rect -236 338 -178 355
rect -418 300 -178 338
rect -120 338 -62 355
rect 62 355 78 372
rect 220 372 376 388
rect 220 355 236 372
rect 62 338 120 355
rect -120 300 120 338
rect 178 338 236 355
rect 360 355 376 372
rect 518 372 674 388
rect 518 355 534 372
rect 360 338 418 355
rect 178 300 418 338
rect 476 338 534 355
rect 658 355 674 372
rect 816 372 972 388
rect 816 355 832 372
rect 658 338 716 355
rect 476 300 716 338
rect 774 338 832 355
rect 956 355 972 372
rect 1114 372 1270 388
rect 1114 355 1130 372
rect 956 338 1014 355
rect 774 300 1014 338
rect 1072 338 1130 355
rect 1254 355 1270 372
rect 1412 372 1568 388
rect 1412 355 1428 372
rect 1254 338 1312 355
rect 1072 300 1312 338
rect 1370 338 1428 355
rect 1552 355 1568 372
rect 1552 338 1610 355
rect 1370 300 1610 338
rect -1610 -338 -1370 -300
rect -1610 -355 -1552 -338
rect -1568 -372 -1552 -355
rect -1428 -355 -1370 -338
rect -1312 -338 -1072 -300
rect -1312 -355 -1254 -338
rect -1428 -372 -1412 -355
rect -1568 -388 -1412 -372
rect -1270 -372 -1254 -355
rect -1130 -355 -1072 -338
rect -1014 -338 -774 -300
rect -1014 -355 -956 -338
rect -1130 -372 -1114 -355
rect -1270 -388 -1114 -372
rect -972 -372 -956 -355
rect -832 -355 -774 -338
rect -716 -338 -476 -300
rect -716 -355 -658 -338
rect -832 -372 -816 -355
rect -972 -388 -816 -372
rect -674 -372 -658 -355
rect -534 -355 -476 -338
rect -418 -338 -178 -300
rect -418 -355 -360 -338
rect -534 -372 -518 -355
rect -674 -388 -518 -372
rect -376 -372 -360 -355
rect -236 -355 -178 -338
rect -120 -338 120 -300
rect -120 -355 -62 -338
rect -236 -372 -220 -355
rect -376 -388 -220 -372
rect -78 -372 -62 -355
rect 62 -355 120 -338
rect 178 -338 418 -300
rect 178 -355 236 -338
rect 62 -372 78 -355
rect -78 -388 78 -372
rect 220 -372 236 -355
rect 360 -355 418 -338
rect 476 -338 716 -300
rect 476 -355 534 -338
rect 360 -372 376 -355
rect 220 -388 376 -372
rect 518 -372 534 -355
rect 658 -355 716 -338
rect 774 -338 1014 -300
rect 774 -355 832 -338
rect 658 -372 674 -355
rect 518 -388 674 -372
rect 816 -372 832 -355
rect 956 -355 1014 -338
rect 1072 -338 1312 -300
rect 1072 -355 1130 -338
rect 956 -372 972 -355
rect 816 -388 972 -372
rect 1114 -372 1130 -355
rect 1254 -355 1312 -338
rect 1370 -338 1610 -300
rect 1370 -355 1428 -338
rect 1254 -372 1270 -355
rect 1114 -388 1270 -372
rect 1412 -372 1428 -355
rect 1552 -355 1610 -338
rect 1552 -372 1568 -355
rect 1412 -388 1568 -372
<< polycont >>
rect -1552 338 -1428 372
rect -1254 338 -1130 372
rect -956 338 -832 372
rect -658 338 -534 372
rect -360 338 -236 372
rect -62 338 62 372
rect 236 338 360 372
rect 534 338 658 372
rect 832 338 956 372
rect 1130 338 1254 372
rect 1428 338 1552 372
rect -1552 -372 -1428 -338
rect -1254 -372 -1130 -338
rect -956 -372 -832 -338
rect -658 -372 -534 -338
rect -360 -372 -236 -338
rect -62 -372 62 -338
rect 236 -372 360 -338
rect 534 -372 658 -338
rect 832 -372 956 -338
rect 1130 -372 1254 -338
rect 1428 -372 1552 -338
<< locali >>
rect -1568 338 -1552 372
rect -1428 338 -1412 372
rect -1270 338 -1254 372
rect -1130 338 -1114 372
rect -972 338 -956 372
rect -832 338 -816 372
rect -674 338 -658 372
rect -534 338 -518 372
rect -376 338 -360 372
rect -236 338 -220 372
rect -78 338 -62 372
rect 62 338 78 372
rect 220 338 236 372
rect 360 338 376 372
rect 518 338 534 372
rect 658 338 674 372
rect 816 338 832 372
rect 956 338 972 372
rect 1114 338 1130 372
rect 1254 338 1270 372
rect 1412 338 1428 372
rect 1552 338 1568 372
rect -1656 288 -1622 304
rect -1656 -304 -1622 -288
rect -1358 288 -1324 304
rect -1358 -304 -1324 -288
rect -1060 288 -1026 304
rect -1060 -304 -1026 -288
rect -762 288 -728 304
rect -762 -304 -728 -288
rect -464 288 -430 304
rect -464 -304 -430 -288
rect -166 288 -132 304
rect -166 -304 -132 -288
rect 132 288 166 304
rect 132 -304 166 -288
rect 430 288 464 304
rect 430 -304 464 -288
rect 728 288 762 304
rect 728 -304 762 -288
rect 1026 288 1060 304
rect 1026 -304 1060 -288
rect 1324 288 1358 304
rect 1324 -304 1358 -288
rect 1622 288 1656 304
rect 1622 -304 1656 -288
rect -1568 -372 -1552 -338
rect -1428 -372 -1412 -338
rect -1270 -372 -1254 -338
rect -1130 -372 -1114 -338
rect -972 -372 -956 -338
rect -832 -372 -816 -338
rect -674 -372 -658 -338
rect -534 -372 -518 -338
rect -376 -372 -360 -338
rect -236 -372 -220 -338
rect -78 -372 -62 -338
rect 62 -372 78 -338
rect 220 -372 236 -338
rect 360 -372 376 -338
rect 518 -372 534 -338
rect 658 -372 674 -338
rect 816 -372 832 -338
rect 956 -372 972 -338
rect 1114 -372 1130 -338
rect 1254 -372 1270 -338
rect 1412 -372 1428 -338
rect 1552 -372 1568 -338
<< viali >>
rect -1532 338 -1448 372
rect -1234 338 -1150 372
rect -936 338 -852 372
rect -638 338 -554 372
rect -340 338 -256 372
rect -42 338 42 372
rect 256 338 340 372
rect 554 338 638 372
rect 852 338 936 372
rect 1150 338 1234 372
rect 1448 338 1532 372
rect -1656 -288 -1622 288
rect -1358 -288 -1324 288
rect -1060 -288 -1026 288
rect -762 -288 -728 288
rect -464 -288 -430 288
rect -166 -288 -132 288
rect 132 -288 166 288
rect 430 -288 464 288
rect 728 -288 762 288
rect 1026 -288 1060 288
rect 1324 -288 1358 288
rect 1622 -288 1656 288
rect -1532 -372 -1448 -338
rect -1234 -372 -1150 -338
rect -936 -372 -852 -338
rect -638 -372 -554 -338
rect -340 -372 -256 -338
rect -42 -372 42 -338
rect 256 -372 340 -338
rect 554 -372 638 -338
rect 852 -372 936 -338
rect 1150 -372 1234 -338
rect 1448 -372 1532 -338
<< metal1 >>
rect -1544 372 -1436 378
rect -1544 338 -1532 372
rect -1448 338 -1436 372
rect -1544 332 -1436 338
rect -1246 372 -1138 378
rect -1246 338 -1234 372
rect -1150 338 -1138 372
rect -1246 332 -1138 338
rect -948 372 -840 378
rect -948 338 -936 372
rect -852 338 -840 372
rect -948 332 -840 338
rect -650 372 -542 378
rect -650 338 -638 372
rect -554 338 -542 372
rect -650 332 -542 338
rect -352 372 -244 378
rect -352 338 -340 372
rect -256 338 -244 372
rect -352 332 -244 338
rect -54 372 54 378
rect -54 338 -42 372
rect 42 338 54 372
rect -54 332 54 338
rect 244 372 352 378
rect 244 338 256 372
rect 340 338 352 372
rect 244 332 352 338
rect 542 372 650 378
rect 542 338 554 372
rect 638 338 650 372
rect 542 332 650 338
rect 840 372 948 378
rect 840 338 852 372
rect 936 338 948 372
rect 840 332 948 338
rect 1138 372 1246 378
rect 1138 338 1150 372
rect 1234 338 1246 372
rect 1138 332 1246 338
rect 1436 372 1544 378
rect 1436 338 1448 372
rect 1532 338 1544 372
rect 1436 332 1544 338
rect -1662 288 -1616 300
rect -1662 -288 -1656 288
rect -1622 -288 -1616 288
rect -1662 -300 -1616 -288
rect -1364 288 -1318 300
rect -1364 -288 -1358 288
rect -1324 -288 -1318 288
rect -1364 -300 -1318 -288
rect -1066 288 -1020 300
rect -1066 -288 -1060 288
rect -1026 -288 -1020 288
rect -1066 -300 -1020 -288
rect -768 288 -722 300
rect -768 -288 -762 288
rect -728 -288 -722 288
rect -768 -300 -722 -288
rect -470 288 -424 300
rect -470 -288 -464 288
rect -430 -288 -424 288
rect -470 -300 -424 -288
rect -172 288 -126 300
rect -172 -288 -166 288
rect -132 -288 -126 288
rect -172 -300 -126 -288
rect 126 288 172 300
rect 126 -288 132 288
rect 166 -288 172 288
rect 126 -300 172 -288
rect 424 288 470 300
rect 424 -288 430 288
rect 464 -288 470 288
rect 424 -300 470 -288
rect 722 288 768 300
rect 722 -288 728 288
rect 762 -288 768 288
rect 722 -300 768 -288
rect 1020 288 1066 300
rect 1020 -288 1026 288
rect 1060 -288 1066 288
rect 1020 -300 1066 -288
rect 1318 288 1364 300
rect 1318 -288 1324 288
rect 1358 -288 1364 288
rect 1318 -300 1364 -288
rect 1616 288 1662 300
rect 1616 -288 1622 288
rect 1656 -288 1662 288
rect 1616 -300 1662 -288
rect -1544 -338 -1436 -332
rect -1544 -372 -1532 -338
rect -1448 -372 -1436 -338
rect -1544 -378 -1436 -372
rect -1246 -338 -1138 -332
rect -1246 -372 -1234 -338
rect -1150 -372 -1138 -338
rect -1246 -378 -1138 -372
rect -948 -338 -840 -332
rect -948 -372 -936 -338
rect -852 -372 -840 -338
rect -948 -378 -840 -372
rect -650 -338 -542 -332
rect -650 -372 -638 -338
rect -554 -372 -542 -338
rect -650 -378 -542 -372
rect -352 -338 -244 -332
rect -352 -372 -340 -338
rect -256 -372 -244 -338
rect -352 -378 -244 -372
rect -54 -338 54 -332
rect -54 -372 -42 -338
rect 42 -372 54 -338
rect -54 -378 54 -372
rect 244 -338 352 -332
rect 244 -372 256 -338
rect 340 -372 352 -338
rect 244 -378 352 -372
rect 542 -338 650 -332
rect 542 -372 554 -338
rect 638 -372 650 -338
rect 542 -378 650 -372
rect 840 -338 948 -332
rect 840 -372 852 -338
rect 936 -372 948 -338
rect 840 -378 948 -372
rect 1138 -338 1246 -332
rect 1138 -372 1150 -338
rect 1234 -372 1246 -338
rect 1138 -378 1246 -372
rect 1436 -338 1544 -332
rect 1436 -372 1448 -338
rect 1532 -372 1544 -338
rect 1436 -378 1544 -372
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string parameters w 3 l 1.2 m 1 nf 11 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 40 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
