magic
tech sky130A
timestamp 1620283077
<< nmoslvt >>
rect -805 -150 -685 150
rect -656 -150 -536 150
rect -507 -150 -387 150
rect -358 -150 -238 150
rect -209 -150 -89 150
rect -60 -150 60 150
rect 89 -150 209 150
rect 238 -150 358 150
rect 387 -150 507 150
rect 536 -150 656 150
rect 685 -150 805 150
<< ndiff >>
rect -834 144 -805 150
rect -834 -144 -828 144
rect -811 -144 -805 144
rect -834 -150 -805 -144
rect -685 144 -656 150
rect -685 -144 -679 144
rect -662 -144 -656 144
rect -685 -150 -656 -144
rect -536 144 -507 150
rect -536 -144 -530 144
rect -513 -144 -507 144
rect -536 -150 -507 -144
rect -387 144 -358 150
rect -387 -144 -381 144
rect -364 -144 -358 144
rect -387 -150 -358 -144
rect -238 144 -209 150
rect -238 -144 -232 144
rect -215 -144 -209 144
rect -238 -150 -209 -144
rect -89 144 -60 150
rect -89 -144 -83 144
rect -66 -144 -60 144
rect -89 -150 -60 -144
rect 60 144 89 150
rect 60 -144 66 144
rect 83 -144 89 144
rect 60 -150 89 -144
rect 209 144 238 150
rect 209 -144 215 144
rect 232 -144 238 144
rect 209 -150 238 -144
rect 358 144 387 150
rect 358 -144 364 144
rect 381 -144 387 144
rect 358 -150 387 -144
rect 507 144 536 150
rect 507 -144 513 144
rect 530 -144 536 144
rect 507 -150 536 -144
rect 656 144 685 150
rect 656 -144 662 144
rect 679 -144 685 144
rect 656 -150 685 -144
rect 805 144 834 150
rect 805 -144 811 144
rect 828 -144 834 144
rect 805 -150 834 -144
<< ndiffc >>
rect -828 -144 -811 144
rect -679 -144 -662 144
rect -530 -144 -513 144
rect -381 -144 -364 144
rect -232 -144 -215 144
rect -83 -144 -66 144
rect 66 -144 83 144
rect 215 -144 232 144
rect 364 -144 381 144
rect 513 -144 530 144
rect 662 -144 679 144
rect 811 -144 828 144
<< poly >>
rect -805 186 -685 194
rect -805 169 -797 186
rect -693 169 -685 186
rect -805 150 -685 169
rect -656 186 -536 194
rect -656 169 -648 186
rect -544 169 -536 186
rect -656 150 -536 169
rect -507 186 -387 194
rect -507 169 -499 186
rect -395 169 -387 186
rect -507 150 -387 169
rect -358 186 -238 194
rect -358 169 -350 186
rect -246 169 -238 186
rect -358 150 -238 169
rect -209 186 -89 194
rect -209 169 -201 186
rect -97 169 -89 186
rect -209 150 -89 169
rect -60 186 60 194
rect -60 169 -52 186
rect 52 169 60 186
rect -60 150 60 169
rect 89 186 209 194
rect 89 169 97 186
rect 201 169 209 186
rect 89 150 209 169
rect 238 186 358 194
rect 238 169 246 186
rect 350 169 358 186
rect 238 150 358 169
rect 387 186 507 194
rect 387 169 395 186
rect 499 169 507 186
rect 387 150 507 169
rect 536 186 656 194
rect 536 169 544 186
rect 648 169 656 186
rect 536 150 656 169
rect 685 186 805 194
rect 685 169 693 186
rect 797 169 805 186
rect 685 150 805 169
rect -805 -169 -685 -150
rect -805 -186 -797 -169
rect -693 -186 -685 -169
rect -805 -194 -685 -186
rect -656 -169 -536 -150
rect -656 -186 -648 -169
rect -544 -186 -536 -169
rect -656 -194 -536 -186
rect -507 -169 -387 -150
rect -507 -186 -499 -169
rect -395 -186 -387 -169
rect -507 -194 -387 -186
rect -358 -169 -238 -150
rect -358 -186 -350 -169
rect -246 -186 -238 -169
rect -358 -194 -238 -186
rect -209 -169 -89 -150
rect -209 -186 -201 -169
rect -97 -186 -89 -169
rect -209 -194 -89 -186
rect -60 -169 60 -150
rect -60 -186 -52 -169
rect 52 -186 60 -169
rect -60 -194 60 -186
rect 89 -169 209 -150
rect 89 -186 97 -169
rect 201 -186 209 -169
rect 89 -194 209 -186
rect 238 -169 358 -150
rect 238 -186 246 -169
rect 350 -186 358 -169
rect 238 -194 358 -186
rect 387 -169 507 -150
rect 387 -186 395 -169
rect 499 -186 507 -169
rect 387 -194 507 -186
rect 536 -169 656 -150
rect 536 -186 544 -169
rect 648 -186 656 -169
rect 536 -194 656 -186
rect 685 -169 805 -150
rect 685 -186 693 -169
rect 797 -186 805 -169
rect 685 -194 805 -186
<< polycont >>
rect -797 169 -693 186
rect -648 169 -544 186
rect -499 169 -395 186
rect -350 169 -246 186
rect -201 169 -97 186
rect -52 169 52 186
rect 97 169 201 186
rect 246 169 350 186
rect 395 169 499 186
rect 544 169 648 186
rect 693 169 797 186
rect -797 -186 -693 -169
rect -648 -186 -544 -169
rect -499 -186 -395 -169
rect -350 -186 -246 -169
rect -201 -186 -97 -169
rect -52 -186 52 -169
rect 97 -186 201 -169
rect 246 -186 350 -169
rect 395 -186 499 -169
rect 544 -186 648 -169
rect 693 -186 797 -169
<< locali >>
rect -805 169 -797 186
rect -693 169 -685 186
rect -656 169 -648 186
rect -544 169 -536 186
rect -507 169 -499 186
rect -395 169 -387 186
rect -358 169 -350 186
rect -246 169 -238 186
rect -209 169 -201 186
rect -97 169 -89 186
rect -60 169 -52 186
rect 52 169 60 186
rect 89 169 97 186
rect 201 169 209 186
rect 238 169 246 186
rect 350 169 358 186
rect 387 169 395 186
rect 499 169 507 186
rect 536 169 544 186
rect 648 169 656 186
rect 685 169 693 186
rect 797 169 805 186
rect -828 144 -811 152
rect -828 -152 -811 -144
rect -679 144 -662 152
rect -679 -152 -662 -144
rect -530 144 -513 152
rect -530 -152 -513 -144
rect -381 144 -364 152
rect -381 -152 -364 -144
rect -232 144 -215 152
rect -232 -152 -215 -144
rect -83 144 -66 152
rect -83 -152 -66 -144
rect 66 144 83 152
rect 66 -152 83 -144
rect 215 144 232 152
rect 215 -152 232 -144
rect 364 144 381 152
rect 364 -152 381 -144
rect 513 144 530 152
rect 513 -152 530 -144
rect 662 144 679 152
rect 662 -152 679 -144
rect 811 144 828 152
rect 811 -152 828 -144
rect -805 -186 -797 -169
rect -693 -186 -685 -169
rect -656 -186 -648 -169
rect -544 -186 -536 -169
rect -507 -186 -499 -169
rect -395 -186 -387 -169
rect -358 -186 -350 -169
rect -246 -186 -238 -169
rect -209 -186 -201 -169
rect -97 -186 -89 -169
rect -60 -186 -52 -169
rect 52 -186 60 -169
rect 89 -186 97 -169
rect 201 -186 209 -169
rect 238 -186 246 -169
rect 350 -186 358 -169
rect 387 -186 395 -169
rect 499 -186 507 -169
rect 536 -186 544 -169
rect 648 -186 656 -169
rect 685 -186 693 -169
rect 797 -186 805 -169
<< viali >>
rect -771 169 -719 186
rect -622 169 -570 186
rect -473 169 -421 186
rect -324 169 -272 186
rect -175 169 -123 186
rect -26 169 26 186
rect 123 169 175 186
rect 272 169 324 186
rect 421 169 473 186
rect 570 169 622 186
rect 719 169 771 186
rect -828 -144 -811 144
rect -679 -144 -662 144
rect -530 -144 -513 144
rect -381 -144 -364 144
rect -232 -144 -215 144
rect -83 -144 -66 144
rect 66 -144 83 144
rect 215 -144 232 144
rect 364 -144 381 144
rect 513 -144 530 144
rect 662 -144 679 144
rect 811 -144 828 144
rect -771 -186 -719 -169
rect -622 -186 -570 -169
rect -473 -186 -421 -169
rect -324 -186 -272 -169
rect -175 -186 -123 -169
rect -26 -186 26 -169
rect 123 -186 175 -169
rect 272 -186 324 -169
rect 421 -186 473 -169
rect 570 -186 622 -169
rect 719 -186 771 -169
<< metal1 >>
rect -777 186 -713 189
rect -777 169 -771 186
rect -719 169 -713 186
rect -777 166 -713 169
rect -628 186 -564 189
rect -628 169 -622 186
rect -570 169 -564 186
rect -628 166 -564 169
rect -479 186 -415 189
rect -479 169 -473 186
rect -421 169 -415 186
rect -479 166 -415 169
rect -330 186 -266 189
rect -330 169 -324 186
rect -272 169 -266 186
rect -330 166 -266 169
rect -181 186 -117 189
rect -181 169 -175 186
rect -123 169 -117 186
rect -181 166 -117 169
rect -32 186 32 189
rect -32 169 -26 186
rect 26 169 32 186
rect -32 166 32 169
rect 117 186 181 189
rect 117 169 123 186
rect 175 169 181 186
rect 117 166 181 169
rect 266 186 330 189
rect 266 169 272 186
rect 324 169 330 186
rect 266 166 330 169
rect 415 186 479 189
rect 415 169 421 186
rect 473 169 479 186
rect 415 166 479 169
rect 564 186 628 189
rect 564 169 570 186
rect 622 169 628 186
rect 564 166 628 169
rect 713 186 777 189
rect 713 169 719 186
rect 771 169 777 186
rect 713 166 777 169
rect -831 144 -808 150
rect -831 -144 -828 144
rect -811 -144 -808 144
rect -831 -150 -808 -144
rect -682 144 -659 150
rect -682 -144 -679 144
rect -662 -144 -659 144
rect -682 -150 -659 -144
rect -533 144 -510 150
rect -533 -144 -530 144
rect -513 -144 -510 144
rect -533 -150 -510 -144
rect -384 144 -361 150
rect -384 -144 -381 144
rect -364 -144 -361 144
rect -384 -150 -361 -144
rect -235 144 -212 150
rect -235 -144 -232 144
rect -215 -144 -212 144
rect -235 -150 -212 -144
rect -86 144 -63 150
rect -86 -144 -83 144
rect -66 -144 -63 144
rect -86 -150 -63 -144
rect 63 144 86 150
rect 63 -144 66 144
rect 83 -144 86 144
rect 63 -150 86 -144
rect 212 144 235 150
rect 212 -144 215 144
rect 232 -144 235 144
rect 212 -150 235 -144
rect 361 144 384 150
rect 361 -144 364 144
rect 381 -144 384 144
rect 361 -150 384 -144
rect 510 144 533 150
rect 510 -144 513 144
rect 530 -144 533 144
rect 510 -150 533 -144
rect 659 144 682 150
rect 659 -144 662 144
rect 679 -144 682 144
rect 659 -150 682 -144
rect 808 144 831 150
rect 808 -144 811 144
rect 828 -144 831 144
rect 808 -150 831 -144
rect -777 -169 -713 -166
rect -777 -186 -771 -169
rect -719 -186 -713 -169
rect -777 -189 -713 -186
rect -628 -169 -564 -166
rect -628 -186 -622 -169
rect -570 -186 -564 -169
rect -628 -189 -564 -186
rect -479 -169 -415 -166
rect -479 -186 -473 -169
rect -421 -186 -415 -169
rect -479 -189 -415 -186
rect -330 -169 -266 -166
rect -330 -186 -324 -169
rect -272 -186 -266 -169
rect -330 -189 -266 -186
rect -181 -169 -117 -166
rect -181 -186 -175 -169
rect -123 -186 -117 -169
rect -181 -189 -117 -186
rect -32 -169 32 -166
rect -32 -186 -26 -169
rect 26 -186 32 -169
rect -32 -189 32 -186
rect 117 -169 181 -166
rect 117 -186 123 -169
rect 175 -186 181 -169
rect 117 -189 181 -186
rect 266 -169 330 -166
rect 266 -186 272 -169
rect 324 -186 330 -169
rect 266 -189 330 -186
rect 415 -169 479 -166
rect 415 -186 421 -169
rect 473 -186 479 -169
rect 415 -189 479 -186
rect 564 -169 628 -166
rect 564 -186 570 -169
rect 622 -186 628 -169
rect 564 -189 628 -186
rect 713 -169 777 -166
rect 713 -186 719 -169
rect 771 -186 777 -169
rect 713 -189 777 -186
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string parameters w 3 l 1.2 m 1 nf 11 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
