magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< error_p >>
rect -5119 -300 -5061 300
rect -4101 -300 -4043 300
rect -3083 -300 -3025 300
rect -2065 -300 -2007 300
rect -1047 -300 -989 300
rect -29 -300 29 300
rect 989 -300 1047 300
rect 2007 -300 2065 300
rect 3025 -300 3083 300
rect 4043 -300 4101 300
rect 5061 -300 5119 300
<< nmos >>
rect -5061 -300 -4101 300
rect -4043 -300 -3083 300
rect -3025 -300 -2065 300
rect -2007 -300 -1047 300
rect -989 -300 -29 300
rect 29 -300 989 300
rect 1047 -300 2007 300
rect 2065 -300 3025 300
rect 3083 -300 4043 300
rect 4101 -300 5061 300
<< ndiff >>
rect -5119 288 -5061 300
rect -5119 -288 -5107 288
rect -5073 -288 -5061 288
rect -5119 -300 -5061 -288
rect -4101 288 -4043 300
rect -4101 -288 -4089 288
rect -4055 -288 -4043 288
rect -4101 -300 -4043 -288
rect -3083 288 -3025 300
rect -3083 -288 -3071 288
rect -3037 -288 -3025 288
rect -3083 -300 -3025 -288
rect -2065 288 -2007 300
rect -2065 -288 -2053 288
rect -2019 -288 -2007 288
rect -2065 -300 -2007 -288
rect -1047 288 -989 300
rect -1047 -288 -1035 288
rect -1001 -288 -989 288
rect -1047 -300 -989 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 989 288 1047 300
rect 989 -288 1001 288
rect 1035 -288 1047 288
rect 989 -300 1047 -288
rect 2007 288 2065 300
rect 2007 -288 2019 288
rect 2053 -288 2065 288
rect 2007 -300 2065 -288
rect 3025 288 3083 300
rect 3025 -288 3037 288
rect 3071 -288 3083 288
rect 3025 -300 3083 -288
rect 4043 288 4101 300
rect 4043 -288 4055 288
rect 4089 -288 4101 288
rect 4043 -300 4101 -288
rect 5061 288 5119 300
rect 5061 -288 5073 288
rect 5107 -288 5119 288
rect 5061 -300 5119 -288
<< ndiffc >>
rect -5107 -288 -5073 288
rect -4089 -288 -4055 288
rect -3071 -288 -3037 288
rect -2053 -288 -2019 288
rect -1035 -288 -1001 288
rect -17 -288 17 288
rect 1001 -288 1035 288
rect 2019 -288 2053 288
rect 3037 -288 3071 288
rect 4055 -288 4089 288
rect 5073 -288 5107 288
<< poly >>
rect -4875 372 -4287 388
rect -4875 355 -4859 372
rect -5061 338 -4859 355
rect -4303 355 -4287 372
rect -3857 372 -3269 388
rect -3857 355 -3841 372
rect -4303 338 -4101 355
rect -5061 300 -4101 338
rect -4043 338 -3841 355
rect -3285 355 -3269 372
rect -2839 372 -2251 388
rect -2839 355 -2823 372
rect -3285 338 -3083 355
rect -4043 300 -3083 338
rect -3025 338 -2823 355
rect -2267 355 -2251 372
rect -1821 372 -1233 388
rect -1821 355 -1805 372
rect -2267 338 -2065 355
rect -3025 300 -2065 338
rect -2007 338 -1805 355
rect -1249 355 -1233 372
rect -803 372 -215 388
rect -803 355 -787 372
rect -1249 338 -1047 355
rect -2007 300 -1047 338
rect -989 338 -787 355
rect -231 355 -215 372
rect 215 372 803 388
rect 215 355 231 372
rect -231 338 -29 355
rect -989 300 -29 338
rect 29 338 231 355
rect 787 355 803 372
rect 1233 372 1821 388
rect 1233 355 1249 372
rect 787 338 989 355
rect 29 300 989 338
rect 1047 338 1249 355
rect 1805 355 1821 372
rect 2251 372 2839 388
rect 2251 355 2267 372
rect 1805 338 2007 355
rect 1047 300 2007 338
rect 2065 338 2267 355
rect 2823 355 2839 372
rect 3269 372 3857 388
rect 3269 355 3285 372
rect 2823 338 3025 355
rect 2065 300 3025 338
rect 3083 338 3285 355
rect 3841 355 3857 372
rect 4287 372 4875 388
rect 4287 355 4303 372
rect 3841 338 4043 355
rect 3083 300 4043 338
rect 4101 338 4303 355
rect 4859 355 4875 372
rect 4859 338 5061 355
rect 4101 300 5061 338
rect -5061 -338 -4101 -300
rect -5061 -355 -4859 -338
rect -4875 -372 -4859 -355
rect -4303 -355 -4101 -338
rect -4043 -338 -3083 -300
rect -4043 -355 -3841 -338
rect -4303 -372 -4287 -355
rect -4875 -388 -4287 -372
rect -3857 -372 -3841 -355
rect -3285 -355 -3083 -338
rect -3025 -338 -2065 -300
rect -3025 -355 -2823 -338
rect -3285 -372 -3269 -355
rect -3857 -388 -3269 -372
rect -2839 -372 -2823 -355
rect -2267 -355 -2065 -338
rect -2007 -338 -1047 -300
rect -2007 -355 -1805 -338
rect -2267 -372 -2251 -355
rect -2839 -388 -2251 -372
rect -1821 -372 -1805 -355
rect -1249 -355 -1047 -338
rect -989 -338 -29 -300
rect -989 -355 -787 -338
rect -1249 -372 -1233 -355
rect -1821 -388 -1233 -372
rect -803 -372 -787 -355
rect -231 -355 -29 -338
rect 29 -338 989 -300
rect 29 -355 231 -338
rect -231 -372 -215 -355
rect -803 -388 -215 -372
rect 215 -372 231 -355
rect 787 -355 989 -338
rect 1047 -338 2007 -300
rect 1047 -355 1249 -338
rect 787 -372 803 -355
rect 215 -388 803 -372
rect 1233 -372 1249 -355
rect 1805 -355 2007 -338
rect 2065 -338 3025 -300
rect 2065 -355 2267 -338
rect 1805 -372 1821 -355
rect 1233 -388 1821 -372
rect 2251 -372 2267 -355
rect 2823 -355 3025 -338
rect 3083 -338 4043 -300
rect 3083 -355 3285 -338
rect 2823 -372 2839 -355
rect 2251 -388 2839 -372
rect 3269 -372 3285 -355
rect 3841 -355 4043 -338
rect 4101 -338 5061 -300
rect 4101 -355 4303 -338
rect 3841 -372 3857 -355
rect 3269 -388 3857 -372
rect 4287 -372 4303 -355
rect 4859 -355 5061 -338
rect 4859 -372 4875 -355
rect 4287 -388 4875 -372
<< polycont >>
rect -4859 338 -4303 372
rect -3841 338 -3285 372
rect -2823 338 -2267 372
rect -1805 338 -1249 372
rect -787 338 -231 372
rect 231 338 787 372
rect 1249 338 1805 372
rect 2267 338 2823 372
rect 3285 338 3841 372
rect 4303 338 4859 372
rect -4859 -372 -4303 -338
rect -3841 -372 -3285 -338
rect -2823 -372 -2267 -338
rect -1805 -372 -1249 -338
rect -787 -372 -231 -338
rect 231 -372 787 -338
rect 1249 -372 1805 -338
rect 2267 -372 2823 -338
rect 3285 -372 3841 -338
rect 4303 -372 4859 -338
<< locali >>
rect -4875 338 -4859 372
rect -4303 338 -4287 372
rect -3857 338 -3841 372
rect -3285 338 -3269 372
rect -2839 338 -2823 372
rect -2267 338 -2251 372
rect -1821 338 -1805 372
rect -1249 338 -1233 372
rect -803 338 -787 372
rect -231 338 -215 372
rect 215 338 231 372
rect 787 338 803 372
rect 1233 338 1249 372
rect 1805 338 1821 372
rect 2251 338 2267 372
rect 2823 338 2839 372
rect 3269 338 3285 372
rect 3841 338 3857 372
rect 4287 338 4303 372
rect 4859 338 4875 372
rect -5107 288 -5073 304
rect -5107 -304 -5073 -288
rect -4089 288 -4055 304
rect -4089 -304 -4055 -288
rect -3071 288 -3037 304
rect -3071 -304 -3037 -288
rect -2053 288 -2019 304
rect -2053 -304 -2019 -288
rect -1035 288 -1001 304
rect -1035 -304 -1001 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 1001 288 1035 304
rect 1001 -304 1035 -288
rect 2019 288 2053 304
rect 2019 -304 2053 -288
rect 3037 288 3071 304
rect 3037 -304 3071 -288
rect 4055 288 4089 304
rect 4055 -304 4089 -288
rect 5073 288 5107 304
rect 5073 -304 5107 -288
rect -4875 -372 -4859 -338
rect -4303 -372 -4287 -338
rect -3857 -372 -3841 -338
rect -3285 -372 -3269 -338
rect -2839 -372 -2823 -338
rect -2267 -372 -2251 -338
rect -1821 -372 -1805 -338
rect -1249 -372 -1233 -338
rect -803 -372 -787 -338
rect -231 -372 -215 -338
rect 215 -372 231 -338
rect 787 -372 803 -338
rect 1233 -372 1249 -338
rect 1805 -372 1821 -338
rect 2251 -372 2267 -338
rect 2823 -372 2839 -338
rect 3269 -372 3285 -338
rect 3841 -372 3857 -338
rect 4287 -372 4303 -338
rect 4859 -372 4875 -338
<< viali >>
rect -4813 338 -4349 372
rect -3795 338 -3331 372
rect -2777 338 -2313 372
rect -1759 338 -1295 372
rect -741 338 -277 372
rect 277 338 741 372
rect 1295 338 1759 372
rect 2313 338 2777 372
rect 3331 338 3795 372
rect 4349 338 4813 372
rect -5107 -288 -5073 288
rect -4089 -288 -4055 288
rect -3071 -288 -3037 288
rect -2053 -288 -2019 288
rect -1035 -288 -1001 288
rect -17 -288 17 288
rect 1001 -288 1035 288
rect 2019 -288 2053 288
rect 3037 -288 3071 288
rect 4055 -288 4089 288
rect 5073 -288 5107 288
rect -4813 -372 -4349 -338
rect -3795 -372 -3331 -338
rect -2777 -372 -2313 -338
rect -1759 -372 -1295 -338
rect -741 -372 -277 -338
rect 277 -372 741 -338
rect 1295 -372 1759 -338
rect 2313 -372 2777 -338
rect 3331 -372 3795 -338
rect 4349 -372 4813 -338
<< metal1 >>
rect -4825 372 -4337 378
rect -4825 338 -4813 372
rect -4349 338 -4337 372
rect -4825 332 -4337 338
rect -3807 372 -3319 378
rect -3807 338 -3795 372
rect -3331 338 -3319 372
rect -3807 332 -3319 338
rect -2789 372 -2301 378
rect -2789 338 -2777 372
rect -2313 338 -2301 372
rect -2789 332 -2301 338
rect -1771 372 -1283 378
rect -1771 338 -1759 372
rect -1295 338 -1283 372
rect -1771 332 -1283 338
rect -753 372 -265 378
rect -753 338 -741 372
rect -277 338 -265 372
rect -753 332 -265 338
rect 265 372 753 378
rect 265 338 277 372
rect 741 338 753 372
rect 265 332 753 338
rect 1283 372 1771 378
rect 1283 338 1295 372
rect 1759 338 1771 372
rect 1283 332 1771 338
rect 2301 372 2789 378
rect 2301 338 2313 372
rect 2777 338 2789 372
rect 2301 332 2789 338
rect 3319 372 3807 378
rect 3319 338 3331 372
rect 3795 338 3807 372
rect 3319 332 3807 338
rect 4337 372 4825 378
rect 4337 338 4349 372
rect 4813 338 4825 372
rect 4337 332 4825 338
rect -5113 288 -5067 300
rect -5113 -288 -5107 288
rect -5073 -288 -5067 288
rect -5113 -300 -5067 -288
rect -4095 288 -4049 300
rect -4095 -288 -4089 288
rect -4055 -288 -4049 288
rect -4095 -300 -4049 -288
rect -3077 288 -3031 300
rect -3077 -288 -3071 288
rect -3037 -288 -3031 288
rect -3077 -300 -3031 -288
rect -2059 288 -2013 300
rect -2059 -288 -2053 288
rect -2019 -288 -2013 288
rect -2059 -300 -2013 -288
rect -1041 288 -995 300
rect -1041 -288 -1035 288
rect -1001 -288 -995 288
rect -1041 -300 -995 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 995 288 1041 300
rect 995 -288 1001 288
rect 1035 -288 1041 288
rect 995 -300 1041 -288
rect 2013 288 2059 300
rect 2013 -288 2019 288
rect 2053 -288 2059 288
rect 2013 -300 2059 -288
rect 3031 288 3077 300
rect 3031 -288 3037 288
rect 3071 -288 3077 288
rect 3031 -300 3077 -288
rect 4049 288 4095 300
rect 4049 -288 4055 288
rect 4089 -288 4095 288
rect 4049 -300 4095 -288
rect 5067 288 5113 300
rect 5067 -288 5073 288
rect 5107 -288 5113 288
rect 5067 -300 5113 -288
rect -4825 -338 -4337 -332
rect -4825 -372 -4813 -338
rect -4349 -372 -4337 -338
rect -4825 -378 -4337 -372
rect -3807 -338 -3319 -332
rect -3807 -372 -3795 -338
rect -3331 -372 -3319 -338
rect -3807 -378 -3319 -372
rect -2789 -338 -2301 -332
rect -2789 -372 -2777 -338
rect -2313 -372 -2301 -338
rect -2789 -378 -2301 -372
rect -1771 -338 -1283 -332
rect -1771 -372 -1759 -338
rect -1295 -372 -1283 -338
rect -1771 -378 -1283 -372
rect -753 -338 -265 -332
rect -753 -372 -741 -338
rect -277 -372 -265 -338
rect -753 -378 -265 -372
rect 265 -338 753 -332
rect 265 -372 277 -338
rect 741 -372 753 -338
rect 265 -378 753 -372
rect 1283 -338 1771 -332
rect 1283 -372 1295 -338
rect 1759 -372 1771 -338
rect 1283 -378 1771 -372
rect 2301 -338 2789 -332
rect 2301 -372 2313 -338
rect 2777 -372 2789 -338
rect 2301 -378 2789 -372
rect 3319 -338 3807 -332
rect 3319 -372 3331 -338
rect 3795 -372 3807 -338
rect 3319 -378 3807 -372
rect 4337 -338 4825 -332
rect 4337 -372 4349 -338
rect 4813 -372 4825 -338
rect 4337 -378 4825 -372
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 3 l 4.8 m 1 nf 10 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
