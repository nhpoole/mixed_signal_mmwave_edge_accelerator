magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1320 -1617 1320 1617
<< metal1 >>
rect -60 300 60 357
rect -60 -357 60 -300
<< rmetal1 >>
rect -60 -300 60 300
<< end >>
