* NGSPICE file created from peak_detector_flat.ext - technology: sky130A

.subckt peak_detector_flat vin ibiasn1 vpeak_out VDD VSS vpeakh rst ibiasn2
X0 se_fold_casc_wide_swing_ota_0/M7d se_fold_casc_wide_swing_ota_0/M7d se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X2 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X4 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X5 se_fold_casc_wide_swing_ota_0/M9d se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X6 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X7 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X8 se_fold_casc_wide_swing_ota_0/vcascpm vpeakh se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X9 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X10 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X11 se_fold_casc_wide_swing_ota_1/vcascpm se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X12 VDD se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X13 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X14 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X15 se_fold_casc_wide_swing_ota_0/vcascpm se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X16 se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X17 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X18 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X19 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X20 VSS vpeakh sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X21 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X22 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X23 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X24 VSS se_fold_casc_wide_swing_ota_1/vbias4 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X25 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X26 se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vbias3 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X27 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X28 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X29 VDD se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X30 se_fold_casc_wide_swing_ota_0/M9d se_fold_casc_wide_swing_ota_0/M9d se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X31 VDD VDD verr VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X32 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X33 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X34 se_fold_casc_wide_swing_ota_1/vtail_cascn vin se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X35 VDD se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X36 se_fold_casc_wide_swing_ota_1/M7d se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X37 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X38 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X39 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X40 se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X41 se_fold_casc_wide_swing_ota_0/vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X42 se_fold_casc_wide_swing_ota_1/vcascnp vin se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X43 VSS se_fold_casc_wide_swing_ota_0/vbias4 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X44 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X45 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X46 VDD VDD se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X47 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X48 VDD se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X49 vpeakh VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X50 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X51 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X52 VDD VDD se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X53 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X54 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X55 se_fold_casc_wide_swing_ota_0/vtail_cascp vpeakh se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X56 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X57 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X58 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X59 se_fold_casc_wide_swing_ota_1/vcascpm vpeak_out se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X60 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X61 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias3 verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X62 se_fold_casc_wide_swing_ota_1/vcascnm vpeak_out se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X63 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X64 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X65 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X66 se_fold_casc_wide_swing_ota_0/vtail_cascp se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X67 se_fold_casc_wide_swing_ota_0/vcascpm se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X68 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X69 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X70 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X71 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X72 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X73 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X74 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X75 se_fold_casc_wide_swing_ota_0/vcascpm se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X76 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X77 VSS ibiasn2 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X78 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X79 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X80 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X81 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X82 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X83 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X84 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X85 se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X86 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X87 se_fold_casc_wide_swing_ota_1/vtail_cascn vin se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X88 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X89 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X90 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X91 VDD se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X92 VDD VDD se_fold_casc_wide_swing_ota_1/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X93 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X94 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X95 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X96 se_fold_casc_wide_swing_ota_1/vcascpp vin se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X97 se_fold_casc_wide_swing_ota_1/vcascpm vpeak_out se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X98 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X99 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X100 se_fold_casc_wide_swing_ota_0/M13d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X101 se_fold_casc_wide_swing_ota_1/vcascpp se_fold_casc_wide_swing_ota_1/vbias2 verr VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X102 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X103 vpeak_out VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X104 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X105 se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X106 VDD VDD se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X107 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X108 VSS ibiasn1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X109 VDD se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X110 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X111 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X112 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X113 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X114 se_fold_casc_wide_swing_ota_1/vtail_cascn vin se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X115 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X116 se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vbias3 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X117 VDD se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X118 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X119 se_fold_casc_wide_swing_ota_1/vcascpp vin se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X120 se_fold_casc_wide_swing_ota_0/M7d se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X121 VDD se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X122 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X123 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X124 se_fold_casc_wide_swing_ota_1/vcascpp vin se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X125 VDD se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X126 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X127 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X128 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X129 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X130 se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X131 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X132 ibiasn2 ibiasn2 ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X133 se_fold_casc_wide_swing_ota_0/vtail_cascp se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X134 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X135 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X136 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X137 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X138 vpeak_out vpeak_out vpeak_out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X139 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X140 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X141 se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X142 se_fold_casc_wide_swing_ota_0/vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X143 se_fold_casc_wide_swing_ota_0/vcascpp se_fold_casc_wide_swing_ota_0/vcascpp se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X144 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X145 se_fold_casc_wide_swing_ota_1/M13d se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X146 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X147 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X148 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X149 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeakh se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X150 VDD se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X151 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X152 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X153 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias3 vpeak_out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X154 se_fold_casc_wide_swing_ota_1/vcascpp vin se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X155 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X156 verr se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X157 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X158 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X159 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X160 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X161 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias3 vpeak_out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X162 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X163 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X164 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X165 se_fold_casc_wide_swing_ota_1/M7d se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X166 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X167 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X168 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X169 se_fold_casc_wide_swing_ota_0/vcascpm vpeakh se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X170 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X171 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X172 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X173 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X174 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X175 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X176 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X177 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X178 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X179 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X180 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X181 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X182 verr se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X183 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias3 vpeak_out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X184 VSS se_fold_casc_wide_swing_ota_0/vbias4 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X185 se_fold_casc_wide_swing_ota_0/M13d se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X186 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X187 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X188 se_fold_casc_wide_swing_ota_0/vcascpm se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X189 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X190 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X191 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X192 se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vbias3 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X193 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X194 se_fold_casc_wide_swing_ota_1/vcascpm se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X195 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X196 se_fold_casc_wide_swing_ota_0/vbias2 ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X197 vpeak_out se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X198 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X199 se_fold_casc_wide_swing_ota_0/vcascpm vpeakh se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X200 verr verr VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X201 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X202 se_fold_casc_wide_swing_ota_1/vtail_cascn vin se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X203 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X204 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X205 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X206 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X207 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X208 se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X209 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X210 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X211 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X212 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X213 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X214 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X215 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X216 se_fold_casc_wide_swing_ota_0/vtail_cascp se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X217 VDD se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X218 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X219 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X220 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X221 se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X222 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X223 verr se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X224 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X225 VSS se_fold_casc_wide_swing_ota_0/vbias4 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X226 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X227 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X228 se_fold_casc_wide_swing_ota_1/vbias2 ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X229 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X230 VDD se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X231 se_fold_casc_wide_swing_ota_0/vcascpp se_fold_casc_wide_swing_ota_0/vcascpp se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X232 se_fold_casc_wide_swing_ota_1/M8d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X233 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X234 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X235 se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X236 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X237 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X238 se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X239 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X240 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X241 se_fold_casc_wide_swing_ota_1/M16d se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X242 vpeakh VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X243 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X244 se_fold_casc_wide_swing_ota_1/M16d se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X245 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X246 se_fold_casc_wide_swing_ota_0/vcascpm se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X247 se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X248 VDD verr vpeakh VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X249 se_fold_casc_wide_swing_ota_1/vtail_cascn vin se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X250 verr se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X251 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X252 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias3 vpeak_out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X253 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X254 VSS vpeakh sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X255 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X256 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X257 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X258 VDD VDD vpeak_out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X259 VDD se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X260 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X261 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X262 se_fold_casc_wide_swing_ota_0/M7d se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X263 se_fold_casc_wide_swing_ota_0/vcascnp vpeak_out se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X264 se_fold_casc_wide_swing_ota_1/vcascpp se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X265 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X266 se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X267 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X268 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X269 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X270 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X271 VDD se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X272 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X273 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X274 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X275 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X276 VDD se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X277 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X278 se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X279 se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X280 VSS vpeak_out sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X281 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X282 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X283 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X284 se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X285 se_fold_casc_wide_swing_ota_0/vcascnm vpeakh se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X286 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X287 se_fold_casc_wide_swing_ota_1/vtail_cascn vin se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X288 VDD se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X289 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X290 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X291 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X292 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X293 VDD se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X294 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X295 se_fold_casc_wide_swing_ota_1/vcascnp vin se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X296 se_fold_casc_wide_swing_ota_1/vtail_cascp se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X297 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X298 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X299 se_fold_casc_wide_swing_ota_1/vcascpm se_fold_casc_wide_swing_ota_1/vcascpm se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X300 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X301 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X302 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X303 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X304 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X305 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X306 se_fold_casc_wide_swing_ota_0/vcascpp se_fold_casc_wide_swing_ota_0/vcascpp se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X307 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X308 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X309 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X310 se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X311 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X312 se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X313 VDD VDD se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X314 se_fold_casc_wide_swing_ota_1/M13d se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X315 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X316 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X317 se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X318 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X319 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X320 se_fold_casc_wide_swing_ota_1/vcascpp se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X321 VSS ibiasn2 ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X322 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X323 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X324 verr verr verr VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X325 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X326 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X327 se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X328 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X329 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X330 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X331 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X332 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X333 se_fold_casc_wide_swing_ota_1/M7d se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X334 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X335 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X336 se_fold_casc_wide_swing_ota_1/M13d se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X337 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X338 se_fold_casc_wide_swing_ota_0/vcascpm se_fold_casc_wide_swing_ota_0/vcascpm se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X339 se_fold_casc_wide_swing_ota_0/vcascpm vpeakh se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X340 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X341 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X342 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X343 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X344 VDD se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X345 se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X346 verr verr verr VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X347 se_fold_casc_wide_swing_ota_1/vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X348 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X349 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X350 VSS ibiasn1 ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X351 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias3 verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X352 se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X353 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X354 se_fold_casc_wide_swing_ota_1/vcascpp vin se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X355 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X356 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X357 vpeak_out se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X358 ibiasn1 ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X359 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X360 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X361 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X362 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X363 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X364 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X365 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X366 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X367 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X368 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X369 se_fold_casc_wide_swing_ota_0/M13d se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X370 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X371 se_fold_casc_wide_swing_ota_0/vcascpp vpeak_out se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X372 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X373 se_fold_casc_wide_swing_ota_0/vcascpm se_fold_casc_wide_swing_ota_0/vcascpm se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X374 se_fold_casc_wide_swing_ota_0/vcascpm vpeakh se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X375 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X376 verr VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X377 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X378 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X379 se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vbias3 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X380 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias3 verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X381 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X382 vpeak_out se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X383 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X384 se_fold_casc_wide_swing_ota_1/vtail_cascp vin se_fold_casc_wide_swing_ota_1/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X385 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X386 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X387 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X388 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X389 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X390 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X391 vpeak_out VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X392 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X393 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X394 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X395 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X396 se_fold_casc_wide_swing_ota_0/M7d se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X397 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias3 verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X398 se_fold_casc_wide_swing_ota_1/M9d se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X399 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X400 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X401 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X402 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X403 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X404 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X405 se_fold_casc_wide_swing_ota_0/vcascpp vpeak_out se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X406 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X407 se_fold_casc_wide_swing_ota_0/vcascpp vpeak_out se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X408 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X409 se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X410 se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X411 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X412 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X413 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X414 se_fold_casc_wide_swing_ota_1/M13d se_fold_casc_wide_swing_ota_1/M13d se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X415 se_fold_casc_wide_swing_ota_1/M9d se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X416 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X417 se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vbias3 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X418 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X419 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X420 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X421 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X422 verr se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X423 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X424 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X425 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X426 VDD se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X427 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X428 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X429 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X430 se_fold_casc_wide_swing_ota_1/M7d se_fold_casc_wide_swing_ota_1/M7d se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X431 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X432 se_fold_casc_wide_swing_ota_0/vcascpp vpeak_out se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X433 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X434 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X435 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X436 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X437 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X438 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X439 se_fold_casc_wide_swing_ota_1/vcascpm se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X440 ibiasn2 ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X441 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X442 se_fold_casc_wide_swing_ota_1/M13d se_fold_casc_wide_swing_ota_1/M13d se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X443 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X444 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X445 se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X446 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X447 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X448 vpeak_out se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X449 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X450 VDD se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X451 se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X452 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X453 se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X454 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X455 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X456 vpeak_out se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X457 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X458 se_fold_casc_wide_swing_ota_0/M8d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X459 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X460 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X461 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X462 se_fold_casc_wide_swing_ota_1/vtail_cascp se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X463 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X464 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X465 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X466 se_fold_casc_wide_swing_ota_0/M16d se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X467 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X468 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X469 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X470 se_fold_casc_wide_swing_ota_0/M16d se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X471 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X472 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X473 VSS vpeak_out sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X474 ibiasn1 ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X475 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X476 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X477 se_fold_casc_wide_swing_ota_1/M16d se_fold_casc_wide_swing_ota_1/M16d VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X478 verr VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X479 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X480 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X481 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X482 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X483 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X484 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X485 VDD se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X486 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X487 se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X488 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X489 VDD se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X490 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X491 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X492 se_fold_casc_wide_swing_ota_0/vcascpp se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X493 se_fold_casc_wide_swing_ota_1/M9d se_fold_casc_wide_swing_ota_1/M9d se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X494 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X495 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X496 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X497 VSS se_fold_casc_wide_swing_ota_1/vbias4 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X498 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X499 se_fold_casc_wide_swing_ota_1/vcascpp se_fold_casc_wide_swing_ota_1/vcascpp se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X500 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X501 VDD se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X502 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X503 VDD se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X504 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X505 ibiasn2 ibiasn2 ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X506 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X507 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X508 vpeak_out se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X509 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X510 VSS se_fold_casc_wide_swing_ota_1/vbias4 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X511 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X512 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X513 se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X514 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X515 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X516 se_fold_casc_wide_swing_ota_1/M7d se_fold_casc_wide_swing_ota_1/M7d se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X517 VSS ibiasn2 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X518 se_fold_casc_wide_swing_ota_1/vcascpp vin se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X519 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X520 se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X521 VDD se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X522 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X523 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X524 se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X525 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X526 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X527 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X528 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X529 se_fold_casc_wide_swing_ota_0/vcascnp vpeak_out se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X530 VDD verr verr VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X531 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X532 VDD se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X533 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X534 se_fold_casc_wide_swing_ota_0/vcascpm se_fold_casc_wide_swing_ota_0/vcascpm se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X535 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X536 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X537 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X538 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X539 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X540 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X541 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X542 VDD se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X543 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X544 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X545 se_fold_casc_wide_swing_ota_0/M13d se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X546 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X547 se_fold_casc_wide_swing_ota_1/M9d se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X548 se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X549 se_fold_casc_wide_swing_ota_0/vcascpp se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X550 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X551 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X552 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias3 vpeak_out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X553 VSS ibiasn1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X554 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X555 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X556 se_fold_casc_wide_swing_ota_1/vcascpp se_fold_casc_wide_swing_ota_1/vcascpp se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X557 vpeak_out vpeak_out vpeak_out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X558 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X559 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X560 se_fold_casc_wide_swing_ota_1/vcascpm vpeak_out se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X561 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X562 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X563 se_fold_casc_wide_swing_ota_1/M9d se_fold_casc_wide_swing_ota_1/M9d se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X564 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X565 ibiasn1 ibiasn1 ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X566 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X567 se_fold_casc_wide_swing_ota_1/vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X568 se_fold_casc_wide_swing_ota_0/M7d se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X569 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X570 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeakh se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X571 verr VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X572 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X573 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias3 verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X574 verr se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X575 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X576 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X577 se_fold_casc_wide_swing_ota_0/M13d se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X578 VSS se_fold_casc_wide_swing_ota_1/vbias4 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X579 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X580 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias3 vpeak_out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X581 vpeak_out vpeak_out vpeak_out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X582 vpeak_out VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X583 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X584 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X585 se_fold_casc_wide_swing_ota_0/vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X586 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X587 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X588 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X589 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X590 se_fold_casc_wide_swing_ota_1/vcascpm vpeak_out se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X591 se_fold_casc_wide_swing_ota_1/vcascpp se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X592 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X593 vpeakh VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X594 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X595 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X596 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias3 vpeak_out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X597 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X598 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X599 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X600 VDD se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X601 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X602 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X603 se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vbias3 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X604 se_fold_casc_wide_swing_ota_1/vcascpp vin se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X605 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X606 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeakh se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X607 se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X608 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeakh se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X609 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X610 se_fold_casc_wide_swing_ota_0/vtail_cascp se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X611 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X612 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X613 se_fold_casc_wide_swing_ota_0/vtail_cascp vpeak_out se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X614 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X615 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X616 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X617 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X618 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X619 se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vbias3 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X620 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X621 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X622 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X623 verr verr verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X624 se_fold_casc_wide_swing_ota_0/M7d se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X625 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X626 se_fold_casc_wide_swing_ota_0/M9d se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X627 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X628 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X629 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X630 se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vbias3 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X631 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X632 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X633 se_fold_casc_wide_swing_ota_1/vcascpp se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X634 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X635 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeakh se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X636 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X637 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X638 se_fold_casc_wide_swing_ota_0/vcascpp vpeak_out se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X639 se_fold_casc_wide_swing_ota_0/vbias2 ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X640 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X641 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X642 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X643 se_fold_casc_wide_swing_ota_1/vcascpp se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X644 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeakh se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X645 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X646 se_fold_casc_wide_swing_ota_0/M13d se_fold_casc_wide_swing_ota_0/M13d se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X647 se_fold_casc_wide_swing_ota_0/M9d se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X648 se_fold_casc_wide_swing_ota_1/M9d se_fold_casc_wide_swing_ota_1/M9d se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X649 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X650 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X651 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X652 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X653 se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X654 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X655 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X656 VDD se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X657 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X658 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X659 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X660 verr se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X661 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X662 se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vbias3 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X663 se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vbias3 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X664 se_fold_casc_wide_swing_ota_0/M7d se_fold_casc_wide_swing_ota_0/M7d se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X665 se_fold_casc_wide_swing_ota_1/vtail_cascp vpeak_out se_fold_casc_wide_swing_ota_1/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X666 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X667 se_fold_casc_wide_swing_ota_1/vbias2 ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X668 se_fold_casc_wide_swing_ota_1/vcascpp se_fold_casc_wide_swing_ota_1/vbias2 verr VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X669 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X670 se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X671 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X672 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X673 verr VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X674 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X675 se_fold_casc_wide_swing_ota_0/M13d se_fold_casc_wide_swing_ota_0/M13d se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X676 se_fold_casc_wide_swing_ota_0/vcascpm se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X677 se_fold_casc_wide_swing_ota_0/M16d se_fold_casc_wide_swing_ota_0/M16d VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X678 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeakh se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X679 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X680 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X681 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X682 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X683 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X684 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X685 se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X686 se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X687 VDD se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X688 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X689 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X690 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X691 VDD se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X692 se_fold_casc_wide_swing_ota_1/vtail_cascp vin se_fold_casc_wide_swing_ota_1/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X693 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X694 se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X695 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X696 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X697 se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X698 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X699 vpeakh rst VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X700 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X701 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X702 se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vbias3 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X703 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X704 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X705 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X706 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X707 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X708 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X709 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X710 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X711 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X712 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X713 se_fold_casc_wide_swing_ota_1/M13d se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X714 se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X715 VSS se_fold_casc_wide_swing_ota_0/vbias4 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X716 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X717 VDD se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X718 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X719 se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X720 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X721 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X722 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X723 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X724 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X725 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X726 se_fold_casc_wide_swing_ota_0/M9d se_fold_casc_wide_swing_ota_0/M9d se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X727 VSS vpeakh sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X728 se_fold_casc_wide_swing_ota_1/vcascpp se_fold_casc_wide_swing_ota_1/vcascpp se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X729 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X730 se_fold_casc_wide_swing_ota_0/vcascpp se_fold_casc_wide_swing_ota_0/vcascpp se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X731 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X732 VDD se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X733 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X734 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X735 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X736 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X737 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X738 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X739 vpeak_out se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X740 VSS verr sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X741 se_fold_casc_wide_swing_ota_1/vcascpp se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X742 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X743 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X744 se_fold_casc_wide_swing_ota_0/M7d se_fold_casc_wide_swing_ota_0/M7d se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X745 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X746 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X747 se_fold_casc_wide_swing_ota_1/vtail_cascn vin se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X748 se_fold_casc_wide_swing_ota_1/vcascpm se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X749 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X750 verr se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X751 se_fold_casc_wide_swing_ota_1/vcascpm se_fold_casc_wide_swing_ota_1/vcascpm se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X752 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X753 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X754 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X755 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X756 VSS ibiasn2 ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X757 VSS vpeak_out sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X758 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X759 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X760 vpeakh verr VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X761 verr se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X762 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias3 vpeak_out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X763 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X764 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X765 VDD VDD se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X766 se_fold_casc_wide_swing_ota_1/vcascpm se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X767 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X768 se_fold_casc_wide_swing_ota_1/vcascpp vin se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X769 VDD se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X770 se_fold_casc_wide_swing_ota_1/M7d se_fold_casc_wide_swing_ota_1/M7d se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X771 VSS se_fold_casc_wide_swing_ota_1/vbias4 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X772 se_fold_casc_wide_swing_ota_0/M9d se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X773 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X774 se_fold_casc_wide_swing_ota_1/M7d se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X775 se_fold_casc_wide_swing_ota_1/M9d se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X776 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X777 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X778 se_fold_casc_wide_swing_ota_0/vtail_cascp se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X779 se_fold_casc_wide_swing_ota_1/vtail_cascn vin se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X780 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X781 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X782 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X783 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X784 VSS ibiasn1 ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X785 se_fold_casc_wide_swing_ota_1/vcascpm se_fold_casc_wide_swing_ota_1/vcascpm se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X786 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X787 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X788 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X789 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X790 se_fold_casc_wide_swing_ota_0/vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X791 se_fold_casc_wide_swing_ota_0/M9d se_fold_casc_wide_swing_ota_0/M9d se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X792 se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X793 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X794 VDD se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X795 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X796 se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vbias3 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X797 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X798 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X799 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X800 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X801 vpeak_out se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X802 se_fold_casc_wide_swing_ota_1/vcascpm vpeak_out se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X803 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X804 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X805 se_fold_casc_wide_swing_ota_1/M13d se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X806 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X807 se_fold_casc_wide_swing_ota_1/vcascpm se_fold_casc_wide_swing_ota_1/vcascpm se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X808 se_fold_casc_wide_swing_ota_0/vcascpp vpeak_out se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X809 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X810 VDD VDD se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X811 VSS se_fold_casc_wide_swing_ota_1/vbias4 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X812 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X813 se_fold_casc_wide_swing_ota_1/M16d se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X814 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X815 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X816 se_fold_casc_wide_swing_ota_0/vcascpp se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X817 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X818 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X819 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X820 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X821 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X822 vpeak_out vpeak_out vpeak_out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X823 VSS se_fold_casc_wide_swing_ota_0/vbias4 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X824 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X825 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X826 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X827 se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vbias3 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X828 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X829 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X830 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X831 se_fold_casc_wide_swing_ota_1/vcascpm vpeak_out se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X832 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X833 VDD se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X834 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeakh se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X835 verr se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X836 VDD se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X837 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X838 se_fold_casc_wide_swing_ota_0/M9d se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X839 se_fold_casc_wide_swing_ota_0/vcascpm vpeakh se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X840 VDD se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X841 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias3 verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X842 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X843 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X844 se_fold_casc_wide_swing_ota_1/vtail_cascp se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X845 se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X846 VDD se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X847 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X848 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X849 VSS verr sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X850 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X851 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X852 se_fold_casc_wide_swing_ota_1/vcascnm vpeak_out se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X853 se_fold_casc_wide_swing_ota_1/vcascpp se_fold_casc_wide_swing_ota_1/vbias2 verr VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X854 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X855 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X856 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X857 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X858 verr se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X859 se_fold_casc_wide_swing_ota_0/vcascpp se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X860 se_fold_casc_wide_swing_ota_1/vtail_cascp se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X861 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X862 se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vbias3 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X863 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X864 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X865 se_fold_casc_wide_swing_ota_1/M16d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X866 se_fold_casc_wide_swing_ota_1/M7d se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X867 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X868 verr se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X869 VDD VDD se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X870 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X871 se_fold_casc_wide_swing_ota_0/vcascpm vpeakh se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X872 se_fold_casc_wide_swing_ota_0/vcascpp se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X873 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X874 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X875 se_fold_casc_wide_swing_ota_0/M9d se_fold_casc_wide_swing_ota_0/M9d se_fold_casc_wide_swing_ota_0/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X876 se_fold_casc_wide_swing_ota_1/M7d se_fold_casc_wide_swing_ota_1/M7d se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X877 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X878 se_fold_casc_wide_swing_ota_0/vcascpp vpeak_out se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X879 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X880 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X881 se_fold_casc_wide_swing_ota_1/M9d se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X882 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X883 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X884 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X885 vpeak_out se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X886 VDD se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X887 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X888 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X889 se_fold_casc_wide_swing_ota_1/vcascpm se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X890 se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X891 VSS se_fold_casc_wide_swing_ota_1/vbias4 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X892 se_fold_casc_wide_swing_ota_0/vtail_cascp vpeakh se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X893 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X894 VSS se_fold_casc_wide_swing_ota_0/vbias4 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X895 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X896 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X897 se_fold_casc_wide_swing_ota_0/vcascpp se_fold_casc_wide_swing_ota_0/vbias2 vpeak_out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X898 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X899 se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X900 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X901 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X902 VDD se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X903 se_fold_casc_wide_swing_ota_1/M9d se_fold_casc_wide_swing_ota_1/M9d se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X904 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X905 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X906 VDD se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X907 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X908 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X909 se_fold_casc_wide_swing_ota_1/vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X910 se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X911 ibiasn1 ibiasn1 ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X912 VDD VDD se_fold_casc_wide_swing_ota_1/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X913 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X914 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X915 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X916 VDD se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X917 se_fold_casc_wide_swing_ota_0/vtail_cascp vpeak_out se_fold_casc_wide_swing_ota_0/vcascnp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X918 VDD se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/M13d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X919 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X920 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X921 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X922 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X923 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X924 VDD VDD se_fold_casc_wide_swing_ota_1/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X925 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X926 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X927 se_fold_casc_wide_swing_ota_1/vtail_cascp vpeak_out se_fold_casc_wide_swing_ota_1/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X928 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X929 se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vbias3 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X930 se_fold_casc_wide_swing_ota_1/vcascpm se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X931 VSS verr sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X932 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X933 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X934 VSS se_fold_casc_wide_swing_ota_1/vbias4 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X935 se_fold_casc_wide_swing_ota_0/M13d se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/M16d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X936 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vmirror VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X937 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X938 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X939 vpeakh VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X940 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X941 se_fold_casc_wide_swing_ota_1/vcascpm se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X942 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X943 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X944 VSS vpeak_out sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X945 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X946 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X947 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X948 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X949 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X950 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X951 se_fold_casc_wide_swing_ota_0/vcascpp se_fold_casc_wide_swing_ota_0/vbias2 vpeak_out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X952 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X953 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X954 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X955 VDD se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X956 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X957 VSS vpeakh sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X958 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X959 se_fold_casc_wide_swing_ota_1/vcascnm se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X960 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X961 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X962 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X963 VDD VDD vpeakh VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X964 se_fold_casc_wide_swing_ota_1/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_1/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X965 se_fold_casc_wide_swing_ota_1/M13d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X966 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X967 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X968 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X969 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=3.1e+07u
X970 VSS se_fold_casc_wide_swing_ota_0/vbias4 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X971 VDD VDD se_fold_casc_wide_swing_ota_1/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X972 se_fold_casc_wide_swing_ota_0/vcascpp se_fold_casc_wide_swing_ota_0/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X973 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X974 VDD se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/M9d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X975 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X976 se_fold_casc_wide_swing_ota_0/vcascpm se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X977 se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vbias3 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X978 vpeakh VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X979 se_fold_casc_wide_swing_ota_1/vcascpm vpeak_out se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X980 a_56554_4138# se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X981 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X982 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X983 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X984 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X985 VDD se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X986 se_fold_casc_wide_swing_ota_1/M7d se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X987 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X988 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X989 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X990 VDD se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X991 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X992 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X993 se_fold_casc_wide_swing_ota_1/vtail_cascn vin se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X994 VDD VDD se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X995 se_fold_casc_wide_swing_ota_0/vcascpm se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X996 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X997 se_fold_casc_wide_swing_ota_0/M7d se_fold_casc_wide_swing_ota_0/M7d se_fold_casc_wide_swing_ota_0/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X998 se_fold_casc_wide_swing_ota_1/vtail_cascp se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X999 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeakh se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1000 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1001 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1002 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1003 se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1004 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1005 se_fold_casc_wide_swing_ota_0/M7d se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1006 se_fold_casc_wide_swing_ota_0/M9d se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1007 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1008 VSS se_fold_casc_wide_swing_ota_0/vbias4 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1009 se_fold_casc_wide_swing_ota_1/vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1010 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1011 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1012 vpeak_out VSS sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.6e+07u
X1013 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1014 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1015 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1016 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1017 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1018 VDD se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1019 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1020 se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vbias3 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1021 se_fold_casc_wide_swing_ota_1/vcascpm vpeak_out se_fold_casc_wide_swing_ota_1/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1022 VDD se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1023 se_fold_casc_wide_swing_ota_1/vtail_cascp se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1024 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1025 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1026 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vbias4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1027 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1028 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1029 se_fold_casc_wide_swing_ota_1/vtail_cascn vin se_fold_casc_wide_swing_ota_1/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1030 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1031 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1032 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1033 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1034 vpeak_out se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1035 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1036 se_fold_casc_wide_swing_ota_0/M13d se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1037 se_fold_casc_wide_swing_ota_0/vcascpm se_fold_casc_wide_swing_ota_0/vcascpm se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1038 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1039 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1040 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X1041 se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1042 verr verr verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1043 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1044 VDD VDD se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1045 se_fold_casc_wide_swing_ota_0/vcascnp se_fold_casc_wide_swing_ota_0/vbias3 vpeak_out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1046 VSS verr sky130_fd_pr__cap_mim_m3_2 l=2.6e+07u w=2.4e+07u
X1047 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1048 se_fold_casc_wide_swing_ota_0/M16d se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/M13d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1049 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1050 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X1051 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1052 se_fold_casc_wide_swing_ota_0/vcascpp vpeak_out se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1053 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1054 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1055 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias3 verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1056 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1057 ibiasn2 ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1058 se_fold_casc_wide_swing_ota_0/vcascpm se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vmirror VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1059 vpeak_out se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1060 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1061 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vcascnm VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1062 se_fold_casc_wide_swing_ota_1/M13d se_fold_casc_wide_swing_ota_1/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1063 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1064 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/vbias3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1065 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1066 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias3 verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1067 VSS se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1068 se_fold_casc_wide_swing_ota_1/vcascpm se_fold_casc_wide_swing_ota_1/vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1069 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeak_out se_fold_casc_wide_swing_ota_0/vcascpp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1070 vpeak_out se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1071 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1072 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1073 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1074 VDD se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1075 se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/M8d se_fold_casc_wide_swing_ota_0/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1076 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1077 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1078 VDD se_fold_casc_wide_swing_ota_1/vmirror se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1079 se_fold_casc_wide_swing_ota_0/vtail_cascn vpeakh se_fold_casc_wide_swing_ota_0/vcascpm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1080 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1081 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=2e+06u
X1082 VDD se_fold_casc_wide_swing_ota_0/vmirror se_fold_casc_wide_swing_ota_0/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1083 se_fold_casc_wide_swing_ota_1/M9d se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/M8d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1084 se_fold_casc_wide_swing_ota_0/vbias2 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1085 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X1086 se_fold_casc_wide_swing_ota_1/vtail_cascn se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1087 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1088 se_fold_casc_wide_swing_ota_0/vcascpm vpeakh se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1089 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1090 se_fold_casc_wide_swing_ota_0/vcascnm vpeakh se_fold_casc_wide_swing_ota_0/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1091 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1092 se_fold_casc_wide_swing_ota_0/vcascpp se_fold_casc_wide_swing_ota_0/vbias2 vpeak_out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1093 vpeak_out se_fold_casc_wide_swing_ota_0/vbias3 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1094 se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vtail_cascn se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1095 se_fold_casc_wide_swing_ota_0/vcascnm se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1096 VSS se_fold_casc_wide_swing_ota_1/vbias4 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1097 se_fold_casc_wide_swing_ota_1/vcascnp se_fold_casc_wide_swing_ota_1/vbias3 verr VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1098 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1099 a_15554_4138# se_fold_casc_wide_swing_ota_0/vbias4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1100 se_fold_casc_wide_swing_ota_0/vtail_cascp se_fold_casc_wide_swing_ota_0/vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1101 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 se_fold_casc_wide_swing_ota_1/M7d VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1102 VSS se_fold_casc_wide_swing_ota_0/vbias4 a_15554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1103 VSS VSS sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=2.9e+07u
X1104 se_fold_casc_wide_swing_ota_0/M16d VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1105 VSS se_fold_casc_wide_swing_ota_0/vbias4 se_fold_casc_wide_swing_ota_0/vtail_cascn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1106 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=2.9e+07u w=4e+06u
X1107 se_fold_casc_wide_swing_ota_1/vbias4 se_fold_casc_wide_swing_ota_1/vbias3 a_56554_4138# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1108 VDD VDD se_fold_casc_wide_swing_ota_0/vcascpm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1109 se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/M8d se_fold_casc_wide_swing_ota_1/M8d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1110 se_fold_casc_wide_swing_ota_1/vcascpp se_fold_casc_wide_swing_ota_1/vcascpp se_fold_casc_wide_swing_ota_1/vcascpp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1111 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias1 se_fold_casc_wide_swing_ota_0/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1112 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vbias2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1113 VDD se_fold_casc_wide_swing_ota_1/vbias1 se_fold_casc_wide_swing_ota_1/vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
X1114 verr se_fold_casc_wide_swing_ota_1/vbias3 se_fold_casc_wide_swing_ota_1/vcascnp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=4.8e+06u
.ends

