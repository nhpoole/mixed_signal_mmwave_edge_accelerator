magic
tech sky130A
timestamp 1626065694
<< checkpaint >>
rect -798 -798 798 798
<< metal4 >>
rect -168 139 168 168
rect -168 -139 -139 139
rect 139 -139 168 139
rect -168 -168 168 -139
<< via4 >>
rect -139 -139 139 139
<< metal5 >>
rect -168 139 168 168
rect -168 -139 -139 139
rect 139 -139 168 139
rect -168 -168 168 -139
<< end >>
