magic
tech sky130A
magscale 1 2
timestamp 1622780374
<< nwell >>
rect 94 333 4678 654
rect 370 -510 4126 -189
<< pwell >>
rect 135 110 221 267
rect 266 93 452 275
rect 1204 229 1386 273
rect 1694 229 2247 275
rect 2952 229 3134 273
rect 3442 229 3995 275
rect 501 93 2247 229
rect 2249 93 3995 229
rect 3997 93 4267 275
rect 4314 93 4500 275
rect 4551 110 4637 267
rect 266 89 287 93
rect 253 55 287 89
rect 529 51 563 93
rect 2277 51 2311 93
rect 4210 55 4244 93
rect 4314 89 4335 93
rect 4301 55 4335 89
rect 411 -123 497 34
rect 501 -85 2247 51
rect 2249 -85 3995 51
rect 1204 -129 1386 -85
rect 1694 -131 2247 -85
rect 2952 -129 3134 -85
rect 3442 -131 3995 -85
rect 3999 -123 4085 34
<< scnmos >>
rect 344 119 374 249
rect 579 119 609 203
rect 663 119 693 203
rect 851 119 881 203
rect 963 119 993 191
rect 1062 119 1092 191
rect 1161 119 1191 203
rect 1280 119 1310 247
rect 1381 119 1411 191
rect 1487 119 1517 191
rect 1582 119 1612 203
rect 1772 119 1802 249
rect 1856 119 1886 249
rect 2044 119 2074 203
rect 2139 119 2169 249
rect 2327 119 2357 203
rect 2411 119 2441 203
rect 2599 119 2629 203
rect 2711 119 2741 191
rect 2810 119 2840 191
rect 2909 119 2939 203
rect 3028 119 3058 247
rect 3129 119 3159 191
rect 3235 119 3265 191
rect 3330 119 3360 203
rect 3520 119 3550 249
rect 3604 119 3634 249
rect 3792 119 3822 203
rect 3887 119 3917 249
rect 4075 119 4105 249
rect 4159 119 4189 249
rect 4392 119 4422 249
rect 579 -59 609 25
rect 663 -59 693 25
rect 851 -59 881 25
rect 963 -47 993 25
rect 1062 -47 1092 25
rect 1161 -59 1191 25
rect 1280 -103 1310 25
rect 1381 -47 1411 25
rect 1487 -47 1517 25
rect 1582 -59 1612 25
rect 1772 -105 1802 25
rect 1856 -105 1886 25
rect 2044 -59 2074 25
rect 2139 -105 2169 25
rect 2327 -59 2357 25
rect 2411 -59 2441 25
rect 2599 -59 2629 25
rect 2711 -47 2741 25
rect 2810 -47 2840 25
rect 2909 -59 2939 25
rect 3028 -103 3058 25
rect 3129 -47 3159 25
rect 3235 -47 3265 25
rect 3330 -59 3360 25
rect 3520 -105 3550 25
rect 3604 -105 3634 25
rect 3792 -59 3822 25
rect 3887 -105 3917 25
<< scpmoshvt >>
rect 344 369 374 569
rect 579 435 609 563
rect 663 435 693 563
rect 851 485 881 569
rect 936 485 966 569
rect 1031 485 1061 569
rect 1134 485 1164 569
rect 1266 419 1296 569
rect 1361 485 1391 569
rect 1445 485 1475 569
rect 1559 485 1589 569
rect 1770 369 1800 569
rect 1854 369 1884 569
rect 2042 441 2072 569
rect 2139 369 2169 569
rect 2327 435 2357 563
rect 2411 435 2441 563
rect 2599 485 2629 569
rect 2684 485 2714 569
rect 2779 485 2809 569
rect 2882 485 2912 569
rect 3014 419 3044 569
rect 3109 485 3139 569
rect 3193 485 3223 569
rect 3307 485 3337 569
rect 3518 369 3548 569
rect 3602 369 3632 569
rect 3790 441 3820 569
rect 3887 369 3917 569
rect 4075 369 4105 569
rect 4159 369 4189 569
rect 4392 369 4422 569
rect 579 -419 609 -291
rect 663 -419 693 -291
rect 851 -425 881 -341
rect 936 -425 966 -341
rect 1031 -425 1061 -341
rect 1134 -425 1164 -341
rect 1266 -425 1296 -275
rect 1361 -425 1391 -341
rect 1445 -425 1475 -341
rect 1559 -425 1589 -341
rect 1770 -425 1800 -225
rect 1854 -425 1884 -225
rect 2042 -425 2072 -297
rect 2139 -425 2169 -225
rect 2327 -419 2357 -291
rect 2411 -419 2441 -291
rect 2599 -425 2629 -341
rect 2684 -425 2714 -341
rect 2779 -425 2809 -341
rect 2882 -425 2912 -341
rect 3014 -425 3044 -275
rect 3109 -425 3139 -341
rect 3193 -425 3223 -341
rect 3307 -425 3337 -341
rect 3518 -425 3548 -225
rect 3602 -425 3632 -225
rect 3790 -425 3820 -297
rect 3887 -425 3917 -225
<< ndiff >>
rect 292 237 344 249
rect 292 203 300 237
rect 334 203 344 237
rect 292 169 344 203
rect 292 135 300 169
rect 334 135 344 169
rect 292 119 344 135
rect 374 237 426 249
rect 374 203 384 237
rect 418 203 426 237
rect 374 169 426 203
rect 374 135 384 169
rect 418 135 426 169
rect 374 119 426 135
rect 527 191 579 203
rect 527 157 535 191
rect 569 157 579 191
rect 527 119 579 157
rect 609 165 663 203
rect 609 131 619 165
rect 653 131 663 165
rect 609 119 663 131
rect 693 191 745 203
rect 693 157 703 191
rect 737 157 745 191
rect 693 119 745 157
rect 799 165 851 203
rect 799 131 807 165
rect 841 131 851 165
rect 799 119 851 131
rect 881 191 931 203
rect 1230 203 1280 247
rect 1111 191 1161 203
rect 881 179 963 191
rect 881 145 892 179
rect 926 145 963 179
rect 881 119 963 145
rect 993 179 1062 191
rect 993 145 1003 179
rect 1037 145 1062 179
rect 993 119 1062 145
rect 1092 119 1161 191
rect 1191 173 1280 203
rect 1191 139 1202 173
rect 1236 139 1280 173
rect 1191 119 1280 139
rect 1310 191 1360 247
rect 1720 234 1772 249
rect 1532 191 1582 203
rect 1310 179 1381 191
rect 1310 145 1321 179
rect 1355 145 1381 179
rect 1310 119 1381 145
rect 1411 179 1487 191
rect 1411 145 1424 179
rect 1458 145 1487 179
rect 1411 119 1487 145
rect 1517 119 1582 191
rect 1612 179 1664 203
rect 1612 145 1622 179
rect 1656 145 1664 179
rect 1612 119 1664 145
rect 1720 200 1728 234
rect 1762 200 1772 234
rect 1720 166 1772 200
rect 1720 132 1728 166
rect 1762 132 1772 166
rect 1720 119 1772 132
rect 1802 195 1856 249
rect 1802 161 1812 195
rect 1846 161 1856 195
rect 1802 119 1856 161
rect 1886 236 1938 249
rect 1886 202 1896 236
rect 1930 202 1938 236
rect 2089 203 2139 249
rect 1886 168 1938 202
rect 1886 134 1896 168
rect 1930 134 1938 168
rect 1886 119 1938 134
rect 1992 191 2044 203
rect 1992 157 2000 191
rect 2034 157 2044 191
rect 1992 119 2044 157
rect 2074 165 2139 203
rect 2074 131 2095 165
rect 2129 131 2139 165
rect 2074 119 2139 131
rect 2169 203 2221 249
rect 2169 169 2179 203
rect 2213 169 2221 203
rect 2169 119 2221 169
rect 2275 191 2327 203
rect 2275 157 2283 191
rect 2317 157 2327 191
rect 2275 119 2327 157
rect 2357 165 2411 203
rect 2357 131 2367 165
rect 2401 131 2411 165
rect 2357 119 2411 131
rect 2441 191 2493 203
rect 2441 157 2451 191
rect 2485 157 2493 191
rect 2441 119 2493 157
rect 2547 165 2599 203
rect 2547 131 2555 165
rect 2589 131 2599 165
rect 2547 119 2599 131
rect 2629 191 2679 203
rect 2978 203 3028 247
rect 2859 191 2909 203
rect 2629 179 2711 191
rect 2629 145 2640 179
rect 2674 145 2711 179
rect 2629 119 2711 145
rect 2741 179 2810 191
rect 2741 145 2751 179
rect 2785 145 2810 179
rect 2741 119 2810 145
rect 2840 119 2909 191
rect 2939 173 3028 203
rect 2939 139 2950 173
rect 2984 139 3028 173
rect 2939 119 3028 139
rect 3058 191 3108 247
rect 3468 234 3520 249
rect 3280 191 3330 203
rect 3058 179 3129 191
rect 3058 145 3069 179
rect 3103 145 3129 179
rect 3058 119 3129 145
rect 3159 179 3235 191
rect 3159 145 3172 179
rect 3206 145 3235 179
rect 3159 119 3235 145
rect 3265 119 3330 191
rect 3360 179 3412 203
rect 3360 145 3370 179
rect 3404 145 3412 179
rect 3360 119 3412 145
rect 3468 200 3476 234
rect 3510 200 3520 234
rect 3468 166 3520 200
rect 3468 132 3476 166
rect 3510 132 3520 166
rect 3468 119 3520 132
rect 3550 195 3604 249
rect 3550 161 3560 195
rect 3594 161 3604 195
rect 3550 119 3604 161
rect 3634 236 3686 249
rect 3634 202 3644 236
rect 3678 202 3686 236
rect 3837 203 3887 249
rect 3634 168 3686 202
rect 3634 134 3644 168
rect 3678 134 3686 168
rect 3634 119 3686 134
rect 3740 191 3792 203
rect 3740 157 3748 191
rect 3782 157 3792 191
rect 3740 119 3792 157
rect 3822 165 3887 203
rect 3822 131 3843 165
rect 3877 131 3887 165
rect 3822 119 3887 131
rect 3917 203 3969 249
rect 3917 169 3927 203
rect 3961 169 3969 203
rect 3917 119 3969 169
rect 4023 233 4075 249
rect 4023 199 4031 233
rect 4065 199 4075 233
rect 4023 165 4075 199
rect 4023 131 4031 165
rect 4065 131 4075 165
rect 4023 119 4075 131
rect 4105 119 4159 249
rect 4189 233 4241 249
rect 4189 199 4199 233
rect 4233 199 4241 233
rect 4189 165 4241 199
rect 4189 131 4199 165
rect 4233 131 4241 165
rect 4189 119 4241 131
rect 4340 237 4392 249
rect 4340 203 4348 237
rect 4382 203 4392 237
rect 4340 169 4392 203
rect 4340 135 4348 169
rect 4382 135 4392 169
rect 4340 119 4392 135
rect 4422 237 4474 249
rect 4422 203 4432 237
rect 4466 203 4474 237
rect 4422 169 4474 203
rect 4422 135 4432 169
rect 4466 135 4474 169
rect 4422 119 4474 135
rect 527 -13 579 25
rect 527 -47 535 -13
rect 569 -47 579 -13
rect 527 -59 579 -47
rect 609 13 663 25
rect 609 -21 619 13
rect 653 -21 663 13
rect 609 -59 663 -21
rect 693 -13 745 25
rect 693 -47 703 -13
rect 737 -47 745 -13
rect 693 -59 745 -47
rect 799 13 851 25
rect 799 -21 807 13
rect 841 -21 851 13
rect 799 -59 851 -21
rect 881 -1 963 25
rect 881 -35 892 -1
rect 926 -35 963 -1
rect 881 -47 963 -35
rect 993 -1 1062 25
rect 993 -35 1003 -1
rect 1037 -35 1062 -1
rect 993 -47 1062 -35
rect 1092 -47 1161 25
rect 881 -59 931 -47
rect 1111 -59 1161 -47
rect 1191 5 1280 25
rect 1191 -29 1202 5
rect 1236 -29 1280 5
rect 1191 -59 1280 -29
rect 1230 -103 1280 -59
rect 1310 -1 1381 25
rect 1310 -35 1321 -1
rect 1355 -35 1381 -1
rect 1310 -47 1381 -35
rect 1411 -1 1487 25
rect 1411 -35 1424 -1
rect 1458 -35 1487 -1
rect 1411 -47 1487 -35
rect 1517 -47 1582 25
rect 1310 -103 1360 -47
rect 1532 -59 1582 -47
rect 1612 -1 1664 25
rect 1612 -35 1622 -1
rect 1656 -35 1664 -1
rect 1612 -59 1664 -35
rect 1720 12 1772 25
rect 1720 -22 1728 12
rect 1762 -22 1772 12
rect 1720 -56 1772 -22
rect 1720 -90 1728 -56
rect 1762 -90 1772 -56
rect 1720 -105 1772 -90
rect 1802 -17 1856 25
rect 1802 -51 1812 -17
rect 1846 -51 1856 -17
rect 1802 -105 1856 -51
rect 1886 10 1938 25
rect 1886 -24 1896 10
rect 1930 -24 1938 10
rect 1886 -58 1938 -24
rect 1886 -92 1896 -58
rect 1930 -92 1938 -58
rect 1992 -13 2044 25
rect 1992 -47 2000 -13
rect 2034 -47 2044 -13
rect 1992 -59 2044 -47
rect 2074 13 2139 25
rect 2074 -21 2095 13
rect 2129 -21 2139 13
rect 2074 -59 2139 -21
rect 1886 -105 1938 -92
rect 2089 -105 2139 -59
rect 2169 -25 2221 25
rect 2169 -59 2179 -25
rect 2213 -59 2221 -25
rect 2275 -13 2327 25
rect 2275 -47 2283 -13
rect 2317 -47 2327 -13
rect 2275 -59 2327 -47
rect 2357 13 2411 25
rect 2357 -21 2367 13
rect 2401 -21 2411 13
rect 2357 -59 2411 -21
rect 2441 -13 2493 25
rect 2441 -47 2451 -13
rect 2485 -47 2493 -13
rect 2441 -59 2493 -47
rect 2547 13 2599 25
rect 2547 -21 2555 13
rect 2589 -21 2599 13
rect 2547 -59 2599 -21
rect 2629 -1 2711 25
rect 2629 -35 2640 -1
rect 2674 -35 2711 -1
rect 2629 -47 2711 -35
rect 2741 -1 2810 25
rect 2741 -35 2751 -1
rect 2785 -35 2810 -1
rect 2741 -47 2810 -35
rect 2840 -47 2909 25
rect 2629 -59 2679 -47
rect 2169 -105 2221 -59
rect 2859 -59 2909 -47
rect 2939 5 3028 25
rect 2939 -29 2950 5
rect 2984 -29 3028 5
rect 2939 -59 3028 -29
rect 2978 -103 3028 -59
rect 3058 -1 3129 25
rect 3058 -35 3069 -1
rect 3103 -35 3129 -1
rect 3058 -47 3129 -35
rect 3159 -1 3235 25
rect 3159 -35 3172 -1
rect 3206 -35 3235 -1
rect 3159 -47 3235 -35
rect 3265 -47 3330 25
rect 3058 -103 3108 -47
rect 3280 -59 3330 -47
rect 3360 -1 3412 25
rect 3360 -35 3370 -1
rect 3404 -35 3412 -1
rect 3360 -59 3412 -35
rect 3468 12 3520 25
rect 3468 -22 3476 12
rect 3510 -22 3520 12
rect 3468 -56 3520 -22
rect 3468 -90 3476 -56
rect 3510 -90 3520 -56
rect 3468 -105 3520 -90
rect 3550 -17 3604 25
rect 3550 -51 3560 -17
rect 3594 -51 3604 -17
rect 3550 -105 3604 -51
rect 3634 10 3686 25
rect 3634 -24 3644 10
rect 3678 -24 3686 10
rect 3634 -58 3686 -24
rect 3634 -92 3644 -58
rect 3678 -92 3686 -58
rect 3740 -13 3792 25
rect 3740 -47 3748 -13
rect 3782 -47 3792 -13
rect 3740 -59 3792 -47
rect 3822 13 3887 25
rect 3822 -21 3843 13
rect 3877 -21 3887 13
rect 3822 -59 3887 -21
rect 3634 -105 3686 -92
rect 3837 -105 3887 -59
rect 3917 -25 3969 25
rect 3917 -59 3927 -25
rect 3961 -59 3969 -25
rect 3917 -105 3969 -59
<< pdiff >>
rect 292 557 344 569
rect 292 523 300 557
rect 334 523 344 557
rect 292 489 344 523
rect 292 455 300 489
rect 334 455 344 489
rect 292 421 344 455
rect 292 387 300 421
rect 334 387 344 421
rect 292 369 344 387
rect 374 557 426 569
rect 374 523 384 557
rect 418 523 426 557
rect 374 489 426 523
rect 374 455 384 489
rect 418 455 426 489
rect 374 421 426 455
rect 527 549 579 563
rect 527 515 535 549
rect 569 515 579 549
rect 527 481 579 515
rect 527 447 535 481
rect 569 447 579 481
rect 527 435 579 447
rect 609 533 663 563
rect 609 499 619 533
rect 653 499 663 533
rect 609 435 663 499
rect 693 549 745 563
rect 693 515 703 549
rect 737 515 745 549
rect 693 481 745 515
rect 799 557 851 569
rect 799 523 807 557
rect 841 523 851 557
rect 799 485 851 523
rect 881 549 936 569
rect 881 515 891 549
rect 925 515 936 549
rect 881 485 936 515
rect 966 544 1031 569
rect 966 510 983 544
rect 1017 510 1031 544
rect 966 485 1031 510
rect 1061 485 1134 569
rect 1164 557 1266 569
rect 1164 523 1222 557
rect 1256 523 1266 557
rect 1164 489 1266 523
rect 1164 485 1222 489
rect 693 447 703 481
rect 737 447 745 481
rect 693 435 745 447
rect 374 387 384 421
rect 418 387 426 421
rect 374 369 426 387
rect 1179 455 1222 485
rect 1256 455 1266 489
rect 1179 419 1266 455
rect 1296 549 1361 569
rect 1296 515 1306 549
rect 1340 515 1361 549
rect 1296 485 1361 515
rect 1391 539 1445 569
rect 1391 505 1401 539
rect 1435 505 1445 539
rect 1391 485 1445 505
rect 1475 485 1559 569
rect 1589 549 1642 569
rect 1589 515 1600 549
rect 1634 515 1642 549
rect 1589 485 1642 515
rect 1716 557 1770 569
rect 1716 523 1724 557
rect 1758 523 1770 557
rect 1716 486 1770 523
rect 1296 419 1346 485
rect 1716 452 1724 486
rect 1758 452 1770 486
rect 1716 415 1770 452
rect 1716 381 1724 415
rect 1758 381 1770 415
rect 1716 369 1770 381
rect 1800 527 1854 569
rect 1800 493 1810 527
rect 1844 493 1854 527
rect 1800 447 1854 493
rect 1800 413 1810 447
rect 1844 413 1854 447
rect 1800 369 1854 413
rect 1884 551 1936 569
rect 1884 517 1894 551
rect 1928 517 1936 551
rect 1884 483 1936 517
rect 1884 449 1894 483
rect 1928 449 1936 483
rect 1884 415 1936 449
rect 1990 557 2042 569
rect 1990 523 1998 557
rect 2032 523 2042 557
rect 1990 489 2042 523
rect 1990 455 1998 489
rect 2032 455 2042 489
rect 1990 441 2042 455
rect 2072 557 2139 569
rect 2072 523 2095 557
rect 2129 523 2139 557
rect 2072 489 2139 523
rect 2072 455 2095 489
rect 2129 455 2139 489
rect 2072 441 2139 455
rect 1884 381 1894 415
rect 1928 381 1936 415
rect 1884 369 1936 381
rect 2087 421 2139 441
rect 2087 387 2095 421
rect 2129 387 2139 421
rect 2087 369 2139 387
rect 2169 557 2221 569
rect 2169 523 2179 557
rect 2213 523 2221 557
rect 2169 486 2221 523
rect 2169 452 2179 486
rect 2213 452 2221 486
rect 2169 415 2221 452
rect 2275 549 2327 563
rect 2275 515 2283 549
rect 2317 515 2327 549
rect 2275 481 2327 515
rect 2275 447 2283 481
rect 2317 447 2327 481
rect 2275 435 2327 447
rect 2357 533 2411 563
rect 2357 499 2367 533
rect 2401 499 2411 533
rect 2357 435 2411 499
rect 2441 549 2493 563
rect 2441 515 2451 549
rect 2485 515 2493 549
rect 2441 481 2493 515
rect 2547 557 2599 569
rect 2547 523 2555 557
rect 2589 523 2599 557
rect 2547 485 2599 523
rect 2629 549 2684 569
rect 2629 515 2639 549
rect 2673 515 2684 549
rect 2629 485 2684 515
rect 2714 544 2779 569
rect 2714 510 2731 544
rect 2765 510 2779 544
rect 2714 485 2779 510
rect 2809 485 2882 569
rect 2912 557 3014 569
rect 2912 523 2970 557
rect 3004 523 3014 557
rect 2912 489 3014 523
rect 2912 485 2970 489
rect 2441 447 2451 481
rect 2485 447 2493 481
rect 2441 435 2493 447
rect 2169 381 2179 415
rect 2213 381 2221 415
rect 2169 369 2221 381
rect 2927 455 2970 485
rect 3004 455 3014 489
rect 2927 419 3014 455
rect 3044 549 3109 569
rect 3044 515 3054 549
rect 3088 515 3109 549
rect 3044 485 3109 515
rect 3139 539 3193 569
rect 3139 505 3149 539
rect 3183 505 3193 539
rect 3139 485 3193 505
rect 3223 485 3307 569
rect 3337 549 3390 569
rect 3337 515 3348 549
rect 3382 515 3390 549
rect 3337 485 3390 515
rect 3464 557 3518 569
rect 3464 523 3472 557
rect 3506 523 3518 557
rect 3464 486 3518 523
rect 3044 419 3094 485
rect 3464 452 3472 486
rect 3506 452 3518 486
rect 3464 415 3518 452
rect 3464 381 3472 415
rect 3506 381 3518 415
rect 3464 369 3518 381
rect 3548 527 3602 569
rect 3548 493 3558 527
rect 3592 493 3602 527
rect 3548 447 3602 493
rect 3548 413 3558 447
rect 3592 413 3602 447
rect 3548 369 3602 413
rect 3632 551 3684 569
rect 3632 517 3642 551
rect 3676 517 3684 551
rect 3632 483 3684 517
rect 3632 449 3642 483
rect 3676 449 3684 483
rect 3632 415 3684 449
rect 3738 557 3790 569
rect 3738 523 3746 557
rect 3780 523 3790 557
rect 3738 489 3790 523
rect 3738 455 3746 489
rect 3780 455 3790 489
rect 3738 441 3790 455
rect 3820 557 3887 569
rect 3820 523 3843 557
rect 3877 523 3887 557
rect 3820 489 3887 523
rect 3820 455 3843 489
rect 3877 455 3887 489
rect 3820 441 3887 455
rect 3632 381 3642 415
rect 3676 381 3684 415
rect 3632 369 3684 381
rect 3835 421 3887 441
rect 3835 387 3843 421
rect 3877 387 3887 421
rect 3835 369 3887 387
rect 3917 557 3969 569
rect 3917 523 3927 557
rect 3961 523 3969 557
rect 3917 486 3969 523
rect 3917 452 3927 486
rect 3961 452 3969 486
rect 3917 415 3969 452
rect 3917 381 3927 415
rect 3961 381 3969 415
rect 3917 369 3969 381
rect 4023 557 4075 569
rect 4023 523 4031 557
rect 4065 523 4075 557
rect 4023 489 4075 523
rect 4023 455 4031 489
rect 4065 455 4075 489
rect 4023 421 4075 455
rect 4023 387 4031 421
rect 4065 387 4075 421
rect 4023 369 4075 387
rect 4105 557 4159 569
rect 4105 523 4115 557
rect 4149 523 4159 557
rect 4105 489 4159 523
rect 4105 455 4115 489
rect 4149 455 4159 489
rect 4105 421 4159 455
rect 4105 387 4115 421
rect 4149 387 4159 421
rect 4105 369 4159 387
rect 4189 557 4241 569
rect 4189 523 4199 557
rect 4233 523 4241 557
rect 4189 489 4241 523
rect 4189 455 4199 489
rect 4233 455 4241 489
rect 4189 421 4241 455
rect 4189 387 4199 421
rect 4233 387 4241 421
rect 4189 369 4241 387
rect 4340 557 4392 569
rect 4340 523 4348 557
rect 4382 523 4392 557
rect 4340 489 4392 523
rect 4340 455 4348 489
rect 4382 455 4392 489
rect 4340 421 4392 455
rect 4340 387 4348 421
rect 4382 387 4392 421
rect 4340 369 4392 387
rect 4422 557 4474 569
rect 4422 523 4432 557
rect 4466 523 4474 557
rect 4422 489 4474 523
rect 4422 455 4432 489
rect 4466 455 4474 489
rect 4422 421 4474 455
rect 4422 387 4432 421
rect 4466 387 4474 421
rect 4422 369 4474 387
rect 527 -303 579 -291
rect 527 -337 535 -303
rect 569 -337 579 -303
rect 527 -371 579 -337
rect 527 -405 535 -371
rect 569 -405 579 -371
rect 527 -419 579 -405
rect 609 -355 663 -291
rect 609 -389 619 -355
rect 653 -389 663 -355
rect 609 -419 663 -389
rect 693 -303 745 -291
rect 693 -337 703 -303
rect 737 -337 745 -303
rect 693 -371 745 -337
rect 1716 -237 1770 -225
rect 1179 -311 1266 -275
rect 1179 -341 1222 -311
rect 693 -405 703 -371
rect 737 -405 745 -371
rect 693 -419 745 -405
rect 799 -379 851 -341
rect 799 -413 807 -379
rect 841 -413 851 -379
rect 799 -425 851 -413
rect 881 -371 936 -341
rect 881 -405 891 -371
rect 925 -405 936 -371
rect 881 -425 936 -405
rect 966 -366 1031 -341
rect 966 -400 983 -366
rect 1017 -400 1031 -366
rect 966 -425 1031 -400
rect 1061 -425 1134 -341
rect 1164 -345 1222 -341
rect 1256 -345 1266 -311
rect 1164 -379 1266 -345
rect 1164 -413 1222 -379
rect 1256 -413 1266 -379
rect 1164 -425 1266 -413
rect 1296 -341 1346 -275
rect 1716 -271 1724 -237
rect 1758 -271 1770 -237
rect 1716 -308 1770 -271
rect 1296 -371 1361 -341
rect 1296 -405 1306 -371
rect 1340 -405 1361 -371
rect 1296 -425 1361 -405
rect 1391 -361 1445 -341
rect 1391 -395 1401 -361
rect 1435 -395 1445 -361
rect 1391 -425 1445 -395
rect 1475 -425 1559 -341
rect 1589 -371 1642 -341
rect 1589 -405 1600 -371
rect 1634 -405 1642 -371
rect 1589 -425 1642 -405
rect 1716 -342 1724 -308
rect 1758 -342 1770 -308
rect 1716 -379 1770 -342
rect 1716 -413 1724 -379
rect 1758 -413 1770 -379
rect 1716 -425 1770 -413
rect 1800 -269 1854 -225
rect 1800 -303 1810 -269
rect 1844 -303 1854 -269
rect 1800 -349 1854 -303
rect 1800 -383 1810 -349
rect 1844 -383 1854 -349
rect 1800 -425 1854 -383
rect 1884 -237 1936 -225
rect 1884 -271 1894 -237
rect 1928 -271 1936 -237
rect 1884 -305 1936 -271
rect 2087 -243 2139 -225
rect 2087 -277 2095 -243
rect 2129 -277 2139 -243
rect 2087 -297 2139 -277
rect 1884 -339 1894 -305
rect 1928 -339 1936 -305
rect 1884 -373 1936 -339
rect 1884 -407 1894 -373
rect 1928 -407 1936 -373
rect 1884 -425 1936 -407
rect 1990 -311 2042 -297
rect 1990 -345 1998 -311
rect 2032 -345 2042 -311
rect 1990 -379 2042 -345
rect 1990 -413 1998 -379
rect 2032 -413 2042 -379
rect 1990 -425 2042 -413
rect 2072 -311 2139 -297
rect 2072 -345 2095 -311
rect 2129 -345 2139 -311
rect 2072 -379 2139 -345
rect 2072 -413 2095 -379
rect 2129 -413 2139 -379
rect 2072 -425 2139 -413
rect 2169 -237 2221 -225
rect 2169 -271 2179 -237
rect 2213 -271 2221 -237
rect 2169 -308 2221 -271
rect 2169 -342 2179 -308
rect 2213 -342 2221 -308
rect 2169 -379 2221 -342
rect 2169 -413 2179 -379
rect 2213 -413 2221 -379
rect 2169 -425 2221 -413
rect 2275 -303 2327 -291
rect 2275 -337 2283 -303
rect 2317 -337 2327 -303
rect 2275 -371 2327 -337
rect 2275 -405 2283 -371
rect 2317 -405 2327 -371
rect 2275 -419 2327 -405
rect 2357 -355 2411 -291
rect 2357 -389 2367 -355
rect 2401 -389 2411 -355
rect 2357 -419 2411 -389
rect 2441 -303 2493 -291
rect 2441 -337 2451 -303
rect 2485 -337 2493 -303
rect 2441 -371 2493 -337
rect 3464 -237 3518 -225
rect 2927 -311 3014 -275
rect 2927 -341 2970 -311
rect 2441 -405 2451 -371
rect 2485 -405 2493 -371
rect 2441 -419 2493 -405
rect 2547 -379 2599 -341
rect 2547 -413 2555 -379
rect 2589 -413 2599 -379
rect 2547 -425 2599 -413
rect 2629 -371 2684 -341
rect 2629 -405 2639 -371
rect 2673 -405 2684 -371
rect 2629 -425 2684 -405
rect 2714 -366 2779 -341
rect 2714 -400 2731 -366
rect 2765 -400 2779 -366
rect 2714 -425 2779 -400
rect 2809 -425 2882 -341
rect 2912 -345 2970 -341
rect 3004 -345 3014 -311
rect 2912 -379 3014 -345
rect 2912 -413 2970 -379
rect 3004 -413 3014 -379
rect 2912 -425 3014 -413
rect 3044 -341 3094 -275
rect 3464 -271 3472 -237
rect 3506 -271 3518 -237
rect 3464 -308 3518 -271
rect 3044 -371 3109 -341
rect 3044 -405 3054 -371
rect 3088 -405 3109 -371
rect 3044 -425 3109 -405
rect 3139 -361 3193 -341
rect 3139 -395 3149 -361
rect 3183 -395 3193 -361
rect 3139 -425 3193 -395
rect 3223 -425 3307 -341
rect 3337 -371 3390 -341
rect 3337 -405 3348 -371
rect 3382 -405 3390 -371
rect 3337 -425 3390 -405
rect 3464 -342 3472 -308
rect 3506 -342 3518 -308
rect 3464 -379 3518 -342
rect 3464 -413 3472 -379
rect 3506 -413 3518 -379
rect 3464 -425 3518 -413
rect 3548 -269 3602 -225
rect 3548 -303 3558 -269
rect 3592 -303 3602 -269
rect 3548 -349 3602 -303
rect 3548 -383 3558 -349
rect 3592 -383 3602 -349
rect 3548 -425 3602 -383
rect 3632 -237 3684 -225
rect 3632 -271 3642 -237
rect 3676 -271 3684 -237
rect 3632 -305 3684 -271
rect 3835 -243 3887 -225
rect 3835 -277 3843 -243
rect 3877 -277 3887 -243
rect 3835 -297 3887 -277
rect 3632 -339 3642 -305
rect 3676 -339 3684 -305
rect 3632 -373 3684 -339
rect 3632 -407 3642 -373
rect 3676 -407 3684 -373
rect 3632 -425 3684 -407
rect 3738 -311 3790 -297
rect 3738 -345 3746 -311
rect 3780 -345 3790 -311
rect 3738 -379 3790 -345
rect 3738 -413 3746 -379
rect 3780 -413 3790 -379
rect 3738 -425 3790 -413
rect 3820 -311 3887 -297
rect 3820 -345 3843 -311
rect 3877 -345 3887 -311
rect 3820 -379 3887 -345
rect 3820 -413 3843 -379
rect 3877 -413 3887 -379
rect 3820 -425 3887 -413
rect 3917 -237 3969 -225
rect 3917 -271 3927 -237
rect 3961 -271 3969 -237
rect 3917 -308 3969 -271
rect 3917 -342 3927 -308
rect 3961 -342 3969 -308
rect 3917 -379 3969 -342
rect 3917 -413 3927 -379
rect 3961 -413 3969 -379
rect 3917 -425 3969 -413
<< ndiffc >>
rect 300 203 334 237
rect 300 135 334 169
rect 384 203 418 237
rect 384 135 418 169
rect 535 157 569 191
rect 619 131 653 165
rect 703 157 737 191
rect 807 131 841 165
rect 892 145 926 179
rect 1003 145 1037 179
rect 1202 139 1236 173
rect 1321 145 1355 179
rect 1424 145 1458 179
rect 1622 145 1656 179
rect 1728 200 1762 234
rect 1728 132 1762 166
rect 1812 161 1846 195
rect 1896 202 1930 236
rect 1896 134 1930 168
rect 2000 157 2034 191
rect 2095 131 2129 165
rect 2179 169 2213 203
rect 2283 157 2317 191
rect 2367 131 2401 165
rect 2451 157 2485 191
rect 2555 131 2589 165
rect 2640 145 2674 179
rect 2751 145 2785 179
rect 2950 139 2984 173
rect 3069 145 3103 179
rect 3172 145 3206 179
rect 3370 145 3404 179
rect 3476 200 3510 234
rect 3476 132 3510 166
rect 3560 161 3594 195
rect 3644 202 3678 236
rect 3644 134 3678 168
rect 3748 157 3782 191
rect 3843 131 3877 165
rect 3927 169 3961 203
rect 4031 199 4065 233
rect 4031 131 4065 165
rect 4199 199 4233 233
rect 4199 131 4233 165
rect 4348 203 4382 237
rect 4348 135 4382 169
rect 4432 203 4466 237
rect 4432 135 4466 169
rect 535 -47 569 -13
rect 619 -21 653 13
rect 703 -47 737 -13
rect 807 -21 841 13
rect 892 -35 926 -1
rect 1003 -35 1037 -1
rect 1202 -29 1236 5
rect 1321 -35 1355 -1
rect 1424 -35 1458 -1
rect 1622 -35 1656 -1
rect 1728 -22 1762 12
rect 1728 -90 1762 -56
rect 1812 -51 1846 -17
rect 1896 -24 1930 10
rect 1896 -92 1930 -58
rect 2000 -47 2034 -13
rect 2095 -21 2129 13
rect 2179 -59 2213 -25
rect 2283 -47 2317 -13
rect 2367 -21 2401 13
rect 2451 -47 2485 -13
rect 2555 -21 2589 13
rect 2640 -35 2674 -1
rect 2751 -35 2785 -1
rect 2950 -29 2984 5
rect 3069 -35 3103 -1
rect 3172 -35 3206 -1
rect 3370 -35 3404 -1
rect 3476 -22 3510 12
rect 3476 -90 3510 -56
rect 3560 -51 3594 -17
rect 3644 -24 3678 10
rect 3644 -92 3678 -58
rect 3748 -47 3782 -13
rect 3843 -21 3877 13
rect 3927 -59 3961 -25
<< pdiffc >>
rect 300 523 334 557
rect 300 455 334 489
rect 300 387 334 421
rect 384 523 418 557
rect 384 455 418 489
rect 535 515 569 549
rect 535 447 569 481
rect 619 499 653 533
rect 703 515 737 549
rect 807 523 841 557
rect 891 515 925 549
rect 983 510 1017 544
rect 1222 523 1256 557
rect 703 447 737 481
rect 384 387 418 421
rect 1222 455 1256 489
rect 1306 515 1340 549
rect 1401 505 1435 539
rect 1600 515 1634 549
rect 1724 523 1758 557
rect 1724 452 1758 486
rect 1724 381 1758 415
rect 1810 493 1844 527
rect 1810 413 1844 447
rect 1894 517 1928 551
rect 1894 449 1928 483
rect 1998 523 2032 557
rect 1998 455 2032 489
rect 2095 523 2129 557
rect 2095 455 2129 489
rect 1894 381 1928 415
rect 2095 387 2129 421
rect 2179 523 2213 557
rect 2179 452 2213 486
rect 2283 515 2317 549
rect 2283 447 2317 481
rect 2367 499 2401 533
rect 2451 515 2485 549
rect 2555 523 2589 557
rect 2639 515 2673 549
rect 2731 510 2765 544
rect 2970 523 3004 557
rect 2451 447 2485 481
rect 2179 381 2213 415
rect 2970 455 3004 489
rect 3054 515 3088 549
rect 3149 505 3183 539
rect 3348 515 3382 549
rect 3472 523 3506 557
rect 3472 452 3506 486
rect 3472 381 3506 415
rect 3558 493 3592 527
rect 3558 413 3592 447
rect 3642 517 3676 551
rect 3642 449 3676 483
rect 3746 523 3780 557
rect 3746 455 3780 489
rect 3843 523 3877 557
rect 3843 455 3877 489
rect 3642 381 3676 415
rect 3843 387 3877 421
rect 3927 523 3961 557
rect 3927 452 3961 486
rect 3927 381 3961 415
rect 4031 523 4065 557
rect 4031 455 4065 489
rect 4031 387 4065 421
rect 4115 523 4149 557
rect 4115 455 4149 489
rect 4115 387 4149 421
rect 4199 523 4233 557
rect 4199 455 4233 489
rect 4199 387 4233 421
rect 4348 523 4382 557
rect 4348 455 4382 489
rect 4348 387 4382 421
rect 4432 523 4466 557
rect 4432 455 4466 489
rect 4432 387 4466 421
rect 535 -337 569 -303
rect 535 -405 569 -371
rect 619 -389 653 -355
rect 703 -337 737 -303
rect 703 -405 737 -371
rect 807 -413 841 -379
rect 891 -405 925 -371
rect 983 -400 1017 -366
rect 1222 -345 1256 -311
rect 1222 -413 1256 -379
rect 1724 -271 1758 -237
rect 1306 -405 1340 -371
rect 1401 -395 1435 -361
rect 1600 -405 1634 -371
rect 1724 -342 1758 -308
rect 1724 -413 1758 -379
rect 1810 -303 1844 -269
rect 1810 -383 1844 -349
rect 1894 -271 1928 -237
rect 2095 -277 2129 -243
rect 1894 -339 1928 -305
rect 1894 -407 1928 -373
rect 1998 -345 2032 -311
rect 1998 -413 2032 -379
rect 2095 -345 2129 -311
rect 2095 -413 2129 -379
rect 2179 -271 2213 -237
rect 2179 -342 2213 -308
rect 2179 -413 2213 -379
rect 2283 -337 2317 -303
rect 2283 -405 2317 -371
rect 2367 -389 2401 -355
rect 2451 -337 2485 -303
rect 2451 -405 2485 -371
rect 2555 -413 2589 -379
rect 2639 -405 2673 -371
rect 2731 -400 2765 -366
rect 2970 -345 3004 -311
rect 2970 -413 3004 -379
rect 3472 -271 3506 -237
rect 3054 -405 3088 -371
rect 3149 -395 3183 -361
rect 3348 -405 3382 -371
rect 3472 -342 3506 -308
rect 3472 -413 3506 -379
rect 3558 -303 3592 -269
rect 3558 -383 3592 -349
rect 3642 -271 3676 -237
rect 3843 -277 3877 -243
rect 3642 -339 3676 -305
rect 3642 -407 3676 -373
rect 3746 -345 3780 -311
rect 3746 -413 3780 -379
rect 3843 -345 3877 -311
rect 3843 -413 3877 -379
rect 3927 -271 3961 -237
rect 3927 -342 3961 -308
rect 3927 -413 3961 -379
<< psubdiff >>
rect 161 217 195 241
rect 161 136 195 183
rect 4577 217 4611 241
rect 4577 136 4611 183
rect 437 -39 471 8
rect 437 -97 471 -73
rect 4025 -39 4059 8
rect 4025 -97 4059 -73
<< nsubdiff >>
rect 161 528 195 552
rect 161 435 195 494
rect 161 377 195 401
rect 4577 528 4611 552
rect 4577 435 4611 494
rect 4577 377 4611 401
rect 437 -257 471 -233
rect 437 -350 471 -291
rect 437 -408 471 -384
rect 4025 -257 4059 -233
rect 4025 -350 4059 -291
rect 4025 -408 4059 -384
<< psubdiffcont >>
rect 161 183 195 217
rect 4577 183 4611 217
rect 437 -73 471 -39
rect 4025 -73 4059 -39
<< nsubdiffcont >>
rect 161 494 195 528
rect 161 401 195 435
rect 4577 494 4611 528
rect 4577 401 4611 435
rect 437 -291 471 -257
rect 437 -384 471 -350
rect 4025 -291 4059 -257
rect 4025 -384 4059 -350
<< poly >>
rect 344 569 374 595
rect 579 563 609 589
rect 663 563 693 589
rect 851 569 881 595
rect 936 569 966 595
rect 1031 569 1061 595
rect 1134 569 1164 595
rect 1266 569 1296 595
rect 1361 569 1391 595
rect 1445 569 1475 595
rect 1559 569 1589 595
rect 1770 569 1800 595
rect 1854 569 1884 595
rect 2042 569 2072 595
rect 2139 569 2169 595
rect 579 420 609 435
rect 546 390 609 420
rect 344 337 374 369
rect 546 337 576 390
rect 663 346 693 435
rect 851 405 881 485
rect 288 321 374 337
rect 288 287 304 321
rect 338 287 374 321
rect 288 271 374 287
rect 522 321 576 337
rect 522 287 532 321
rect 566 287 576 321
rect 618 336 693 346
rect 786 389 881 405
rect 786 355 796 389
rect 830 355 881 389
rect 936 369 966 485
rect 1031 453 1061 485
rect 1031 437 1092 453
rect 1031 403 1048 437
rect 1082 403 1092 437
rect 1031 387 1092 403
rect 786 339 881 355
rect 618 302 634 336
rect 668 302 693 336
rect 618 292 693 302
rect 522 271 576 287
rect 344 249 374 271
rect 546 248 576 271
rect 546 218 609 248
rect 579 203 609 218
rect 663 203 693 292
rect 851 203 881 339
rect 923 359 989 369
rect 923 325 939 359
rect 973 345 989 359
rect 973 325 1092 345
rect 923 315 1092 325
rect 943 263 1009 273
rect 943 229 959 263
rect 993 229 1009 263
rect 943 219 1009 229
rect 963 191 993 219
rect 1062 191 1092 315
rect 1134 285 1164 485
rect 1266 381 1296 419
rect 1361 387 1391 485
rect 1445 447 1475 485
rect 1559 453 1589 485
rect 1444 437 1510 447
rect 1444 403 1460 437
rect 1494 403 1510 437
rect 1444 393 1510 403
rect 1559 437 1640 453
rect 1559 403 1596 437
rect 1630 403 1640 437
rect 1559 387 1640 403
rect 1206 371 1296 381
rect 1206 337 1222 371
rect 1256 337 1296 371
rect 1206 327 1296 337
rect 1266 292 1296 327
rect 1348 371 1402 387
rect 1348 337 1358 371
rect 1392 351 1402 371
rect 1392 337 1517 351
rect 1348 321 1517 337
rect 1134 275 1208 285
rect 1134 241 1158 275
rect 1192 241 1208 275
rect 1266 262 1310 292
rect 1280 247 1310 262
rect 1381 263 1445 279
rect 1134 231 1208 241
rect 1161 203 1191 231
rect 1381 229 1401 263
rect 1435 229 1445 263
rect 1381 213 1445 229
rect 1381 191 1411 213
rect 1487 191 1517 321
rect 1582 203 1612 387
rect 2042 405 2072 441
rect 2033 375 2072 405
rect 1770 337 1800 369
rect 1854 337 1884 369
rect 2033 337 2063 375
rect 2327 563 2357 589
rect 2411 563 2441 589
rect 2599 569 2629 595
rect 2684 569 2714 595
rect 2779 569 2809 595
rect 2882 569 2912 595
rect 3014 569 3044 595
rect 3109 569 3139 595
rect 3193 569 3223 595
rect 3307 569 3337 595
rect 3518 569 3548 595
rect 3602 569 3632 595
rect 3790 569 3820 595
rect 3887 569 3917 595
rect 4075 569 4105 595
rect 4159 569 4189 595
rect 4392 569 4422 595
rect 2327 420 2357 435
rect 2294 390 2357 420
rect 2139 337 2169 369
rect 2294 337 2324 390
rect 2411 346 2441 435
rect 2599 405 2629 485
rect 1660 321 1802 337
rect 1660 287 1670 321
rect 1704 287 1802 321
rect 1660 271 1802 287
rect 1844 321 2063 337
rect 1844 287 1854 321
rect 1888 287 2063 321
rect 1844 271 2063 287
rect 2105 321 2169 337
rect 2105 287 2115 321
rect 2149 287 2169 321
rect 2105 271 2169 287
rect 2270 321 2324 337
rect 2270 287 2280 321
rect 2314 287 2324 321
rect 2366 336 2441 346
rect 2534 389 2629 405
rect 2534 355 2544 389
rect 2578 355 2629 389
rect 2684 369 2714 485
rect 2779 453 2809 485
rect 2779 437 2840 453
rect 2779 403 2796 437
rect 2830 403 2840 437
rect 2779 387 2840 403
rect 2534 339 2629 355
rect 2366 302 2382 336
rect 2416 302 2441 336
rect 2366 292 2441 302
rect 2270 271 2324 287
rect 1772 249 1802 271
rect 1856 249 1886 271
rect 2033 242 2063 271
rect 2139 249 2169 271
rect 2033 218 2074 242
rect 2044 203 2074 218
rect 2294 248 2324 271
rect 2294 218 2357 248
rect 2327 203 2357 218
rect 2411 203 2441 292
rect 2599 203 2629 339
rect 2671 359 2737 369
rect 2671 325 2687 359
rect 2721 345 2737 359
rect 2721 325 2840 345
rect 2671 315 2840 325
rect 2691 263 2757 273
rect 2691 229 2707 263
rect 2741 229 2757 263
rect 2691 219 2757 229
rect 2711 191 2741 219
rect 2810 191 2840 315
rect 2882 285 2912 485
rect 3014 381 3044 419
rect 3109 387 3139 485
rect 3193 447 3223 485
rect 3307 453 3337 485
rect 3192 437 3258 447
rect 3192 403 3208 437
rect 3242 403 3258 437
rect 3192 393 3258 403
rect 3307 437 3388 453
rect 3307 403 3344 437
rect 3378 403 3388 437
rect 3307 387 3388 403
rect 2954 371 3044 381
rect 2954 337 2970 371
rect 3004 337 3044 371
rect 2954 327 3044 337
rect 3014 292 3044 327
rect 3096 371 3150 387
rect 3096 337 3106 371
rect 3140 351 3150 371
rect 3140 337 3265 351
rect 3096 321 3265 337
rect 2882 275 2956 285
rect 2882 241 2906 275
rect 2940 241 2956 275
rect 3014 262 3058 292
rect 3028 247 3058 262
rect 3129 263 3193 279
rect 2882 231 2956 241
rect 2909 203 2939 231
rect 3129 229 3149 263
rect 3183 229 3193 263
rect 3129 213 3193 229
rect 3129 191 3159 213
rect 3235 191 3265 321
rect 3330 203 3360 387
rect 3790 405 3820 441
rect 3781 375 3820 405
rect 3518 337 3548 369
rect 3602 337 3632 369
rect 3781 337 3811 375
rect 3887 337 3917 369
rect 4075 337 4105 369
rect 3408 321 3550 337
rect 3408 287 3418 321
rect 3452 287 3550 321
rect 3408 271 3550 287
rect 3592 321 3811 337
rect 3592 287 3602 321
rect 3636 287 3811 321
rect 3592 271 3811 287
rect 3853 321 3917 337
rect 3853 287 3863 321
rect 3897 287 3917 321
rect 3853 271 3917 287
rect 4017 321 4105 337
rect 4017 287 4034 321
rect 4068 287 4105 321
rect 4017 271 4105 287
rect 3520 249 3550 271
rect 3604 249 3634 271
rect 3781 242 3811 271
rect 3887 249 3917 271
rect 4075 249 4105 271
rect 4159 337 4189 369
rect 4392 337 4422 369
rect 4159 321 4251 337
rect 4159 287 4202 321
rect 4236 287 4251 321
rect 4159 271 4251 287
rect 4336 321 4422 337
rect 4336 287 4352 321
rect 4386 287 4422 321
rect 4336 271 4422 287
rect 4159 249 4189 271
rect 4392 249 4422 271
rect 3781 218 3822 242
rect 3792 203 3822 218
rect 344 93 374 119
rect 579 93 609 119
rect 663 93 693 119
rect 851 93 881 119
rect 963 93 993 119
rect 1062 93 1092 119
rect 1161 93 1191 119
rect 1280 93 1310 119
rect 1381 93 1411 119
rect 1487 93 1517 119
rect 1582 93 1612 119
rect 1772 93 1802 119
rect 1856 93 1886 119
rect 2044 93 2074 119
rect 2139 93 2169 119
rect 2327 93 2357 119
rect 2411 93 2441 119
rect 2599 93 2629 119
rect 2711 93 2741 119
rect 2810 93 2840 119
rect 2909 93 2939 119
rect 3028 93 3058 119
rect 3129 93 3159 119
rect 3235 93 3265 119
rect 3330 93 3360 119
rect 3520 93 3550 119
rect 3604 93 3634 119
rect 3792 93 3822 119
rect 3887 93 3917 119
rect 4075 93 4105 119
rect 4159 93 4189 119
rect 4392 93 4422 119
rect 579 25 609 51
rect 663 25 693 51
rect 851 25 881 51
rect 963 25 993 51
rect 1062 25 1092 51
rect 1161 25 1191 51
rect 1280 25 1310 51
rect 1381 25 1411 51
rect 1487 25 1517 51
rect 1582 25 1612 51
rect 1772 25 1802 51
rect 1856 25 1886 51
rect 2044 25 2074 51
rect 2139 25 2169 51
rect 2327 25 2357 51
rect 2411 25 2441 51
rect 2599 25 2629 51
rect 2711 25 2741 51
rect 2810 25 2840 51
rect 2909 25 2939 51
rect 3028 25 3058 51
rect 3129 25 3159 51
rect 3235 25 3265 51
rect 3330 25 3360 51
rect 3520 25 3550 51
rect 3604 25 3634 51
rect 3792 25 3822 51
rect 3887 25 3917 51
rect 579 -74 609 -59
rect 546 -104 609 -74
rect 546 -127 576 -104
rect 522 -143 576 -127
rect 522 -177 532 -143
rect 566 -177 576 -143
rect 663 -148 693 -59
rect 522 -193 576 -177
rect 546 -246 576 -193
rect 618 -158 693 -148
rect 618 -192 634 -158
rect 668 -192 693 -158
rect 618 -202 693 -192
rect 851 -195 881 -59
rect 963 -75 993 -47
rect 943 -85 1009 -75
rect 943 -119 959 -85
rect 993 -119 1009 -85
rect 943 -129 1009 -119
rect 1062 -171 1092 -47
rect 1161 -87 1191 -59
rect 546 -276 609 -246
rect 579 -291 609 -276
rect 663 -291 693 -202
rect 786 -211 881 -195
rect 786 -245 796 -211
rect 830 -245 881 -211
rect 923 -181 1092 -171
rect 923 -215 939 -181
rect 973 -201 1092 -181
rect 1134 -97 1208 -87
rect 1134 -131 1158 -97
rect 1192 -131 1208 -97
rect 1381 -69 1411 -47
rect 1381 -85 1445 -69
rect 1280 -118 1310 -103
rect 1134 -141 1208 -131
rect 973 -215 989 -201
rect 923 -225 989 -215
rect 786 -261 881 -245
rect 851 -341 881 -261
rect 936 -341 966 -225
rect 1031 -259 1092 -243
rect 1031 -293 1048 -259
rect 1082 -293 1092 -259
rect 1031 -309 1092 -293
rect 1031 -341 1061 -309
rect 1134 -341 1164 -141
rect 1266 -148 1310 -118
rect 1381 -119 1401 -85
rect 1435 -119 1445 -85
rect 1381 -135 1445 -119
rect 1266 -183 1296 -148
rect 1487 -177 1517 -47
rect 1206 -193 1296 -183
rect 1206 -227 1222 -193
rect 1256 -227 1296 -193
rect 1206 -237 1296 -227
rect 1266 -275 1296 -237
rect 1348 -193 1517 -177
rect 1348 -227 1358 -193
rect 1392 -207 1517 -193
rect 1392 -227 1402 -207
rect 1348 -243 1402 -227
rect 1582 -243 1612 -59
rect 2044 -74 2074 -59
rect 2033 -98 2074 -74
rect 1772 -127 1802 -105
rect 1856 -127 1886 -105
rect 2033 -127 2063 -98
rect 2327 -74 2357 -59
rect 2294 -104 2357 -74
rect 2139 -127 2169 -105
rect 2294 -127 2324 -104
rect 1660 -143 1802 -127
rect 1660 -177 1670 -143
rect 1704 -177 1802 -143
rect 1660 -193 1802 -177
rect 1844 -143 2063 -127
rect 1844 -177 1854 -143
rect 1888 -177 2063 -143
rect 1844 -193 2063 -177
rect 2105 -143 2169 -127
rect 2105 -177 2115 -143
rect 2149 -177 2169 -143
rect 2105 -193 2169 -177
rect 2270 -143 2324 -127
rect 2270 -177 2280 -143
rect 2314 -177 2324 -143
rect 2411 -148 2441 -59
rect 2270 -193 2324 -177
rect 1770 -225 1800 -193
rect 1854 -225 1884 -193
rect 579 -445 609 -419
rect 663 -445 693 -419
rect 1361 -341 1391 -243
rect 1444 -259 1510 -249
rect 1444 -293 1460 -259
rect 1494 -293 1510 -259
rect 1444 -303 1510 -293
rect 1559 -259 1640 -243
rect 1559 -293 1596 -259
rect 1630 -293 1640 -259
rect 1445 -341 1475 -303
rect 1559 -309 1640 -293
rect 1559 -341 1589 -309
rect 2033 -231 2063 -193
rect 2139 -225 2169 -193
rect 2033 -261 2072 -231
rect 2042 -297 2072 -261
rect 2294 -246 2324 -193
rect 2366 -158 2441 -148
rect 2366 -192 2382 -158
rect 2416 -192 2441 -158
rect 2366 -202 2441 -192
rect 2599 -195 2629 -59
rect 2711 -75 2741 -47
rect 2691 -85 2757 -75
rect 2691 -119 2707 -85
rect 2741 -119 2757 -85
rect 2691 -129 2757 -119
rect 2810 -171 2840 -47
rect 2909 -87 2939 -59
rect 2294 -276 2357 -246
rect 2327 -291 2357 -276
rect 2411 -291 2441 -202
rect 2534 -211 2629 -195
rect 2534 -245 2544 -211
rect 2578 -245 2629 -211
rect 2671 -181 2840 -171
rect 2671 -215 2687 -181
rect 2721 -201 2840 -181
rect 2882 -97 2956 -87
rect 2882 -131 2906 -97
rect 2940 -131 2956 -97
rect 3129 -69 3159 -47
rect 3129 -85 3193 -69
rect 3028 -118 3058 -103
rect 2882 -141 2956 -131
rect 2721 -215 2737 -201
rect 2671 -225 2737 -215
rect 2534 -261 2629 -245
rect 2599 -341 2629 -261
rect 2684 -341 2714 -225
rect 2779 -259 2840 -243
rect 2779 -293 2796 -259
rect 2830 -293 2840 -259
rect 2779 -309 2840 -293
rect 2779 -341 2809 -309
rect 2882 -341 2912 -141
rect 3014 -148 3058 -118
rect 3129 -119 3149 -85
rect 3183 -119 3193 -85
rect 3129 -135 3193 -119
rect 3014 -183 3044 -148
rect 3235 -177 3265 -47
rect 2954 -193 3044 -183
rect 2954 -227 2970 -193
rect 3004 -227 3044 -193
rect 2954 -237 3044 -227
rect 3014 -275 3044 -237
rect 3096 -193 3265 -177
rect 3096 -227 3106 -193
rect 3140 -207 3265 -193
rect 3140 -227 3150 -207
rect 3096 -243 3150 -227
rect 3330 -243 3360 -59
rect 3792 -74 3822 -59
rect 3781 -98 3822 -74
rect 3520 -127 3550 -105
rect 3604 -127 3634 -105
rect 3781 -127 3811 -98
rect 3887 -127 3917 -105
rect 3408 -143 3550 -127
rect 3408 -177 3418 -143
rect 3452 -177 3550 -143
rect 3408 -193 3550 -177
rect 3592 -143 3811 -127
rect 3592 -177 3602 -143
rect 3636 -177 3811 -143
rect 3592 -193 3811 -177
rect 3853 -143 3917 -127
rect 3853 -177 3863 -143
rect 3897 -177 3917 -143
rect 3853 -193 3917 -177
rect 3518 -225 3548 -193
rect 3602 -225 3632 -193
rect 851 -451 881 -425
rect 936 -451 966 -425
rect 1031 -451 1061 -425
rect 1134 -451 1164 -425
rect 1266 -451 1296 -425
rect 1361 -451 1391 -425
rect 1445 -451 1475 -425
rect 1559 -451 1589 -425
rect 1770 -451 1800 -425
rect 1854 -451 1884 -425
rect 2042 -451 2072 -425
rect 2139 -451 2169 -425
rect 2327 -445 2357 -419
rect 2411 -445 2441 -419
rect 3109 -341 3139 -243
rect 3192 -259 3258 -249
rect 3192 -293 3208 -259
rect 3242 -293 3258 -259
rect 3192 -303 3258 -293
rect 3307 -259 3388 -243
rect 3307 -293 3344 -259
rect 3378 -293 3388 -259
rect 3193 -341 3223 -303
rect 3307 -309 3388 -293
rect 3307 -341 3337 -309
rect 3781 -231 3811 -193
rect 3887 -225 3917 -193
rect 3781 -261 3820 -231
rect 3790 -297 3820 -261
rect 2599 -451 2629 -425
rect 2684 -451 2714 -425
rect 2779 -451 2809 -425
rect 2882 -451 2912 -425
rect 3014 -451 3044 -425
rect 3109 -451 3139 -425
rect 3193 -451 3223 -425
rect 3307 -451 3337 -425
rect 3518 -451 3548 -425
rect 3602 -451 3632 -425
rect 3790 -451 3820 -425
rect 3887 -451 3917 -425
<< polycont >>
rect 304 287 338 321
rect 532 287 566 321
rect 796 355 830 389
rect 1048 403 1082 437
rect 634 302 668 336
rect 939 325 973 359
rect 959 229 993 263
rect 1460 403 1494 437
rect 1596 403 1630 437
rect 1222 337 1256 371
rect 1358 337 1392 371
rect 1158 241 1192 275
rect 1401 229 1435 263
rect 1670 287 1704 321
rect 1854 287 1888 321
rect 2115 287 2149 321
rect 2280 287 2314 321
rect 2544 355 2578 389
rect 2796 403 2830 437
rect 2382 302 2416 336
rect 2687 325 2721 359
rect 2707 229 2741 263
rect 3208 403 3242 437
rect 3344 403 3378 437
rect 2970 337 3004 371
rect 3106 337 3140 371
rect 2906 241 2940 275
rect 3149 229 3183 263
rect 3418 287 3452 321
rect 3602 287 3636 321
rect 3863 287 3897 321
rect 4034 287 4068 321
rect 4202 287 4236 321
rect 4352 287 4386 321
rect 532 -177 566 -143
rect 634 -192 668 -158
rect 959 -119 993 -85
rect 796 -245 830 -211
rect 939 -215 973 -181
rect 1158 -131 1192 -97
rect 1048 -293 1082 -259
rect 1401 -119 1435 -85
rect 1222 -227 1256 -193
rect 1358 -227 1392 -193
rect 1670 -177 1704 -143
rect 1854 -177 1888 -143
rect 2115 -177 2149 -143
rect 2280 -177 2314 -143
rect 1460 -293 1494 -259
rect 1596 -293 1630 -259
rect 2382 -192 2416 -158
rect 2707 -119 2741 -85
rect 2544 -245 2578 -211
rect 2687 -215 2721 -181
rect 2906 -131 2940 -97
rect 2796 -293 2830 -259
rect 3149 -119 3183 -85
rect 2970 -227 3004 -193
rect 3106 -227 3140 -193
rect 3418 -177 3452 -143
rect 3602 -177 3636 -143
rect 3863 -177 3897 -143
rect 3208 -293 3242 -259
rect 3344 -293 3378 -259
<< locali >>
rect 132 599 161 633
rect 195 599 253 633
rect 287 599 345 633
rect 379 599 437 633
rect 471 599 529 633
rect 563 599 621 633
rect 655 599 713 633
rect 747 599 805 633
rect 839 599 897 633
rect 931 599 989 633
rect 1023 599 1081 633
rect 1115 599 1173 633
rect 1207 599 1265 633
rect 1299 599 1357 633
rect 1391 599 1449 633
rect 1483 599 1541 633
rect 1575 599 1633 633
rect 1667 599 1725 633
rect 1759 599 1817 633
rect 1851 599 1909 633
rect 1943 599 2001 633
rect 2035 599 2093 633
rect 2127 599 2185 633
rect 2219 599 2277 633
rect 2311 599 2369 633
rect 2403 599 2461 633
rect 2495 599 2553 633
rect 2587 599 2645 633
rect 2679 599 2737 633
rect 2771 599 2829 633
rect 2863 599 2921 633
rect 2955 599 3013 633
rect 3047 599 3105 633
rect 3139 599 3197 633
rect 3231 599 3289 633
rect 3323 599 3381 633
rect 3415 599 3473 633
rect 3507 599 3565 633
rect 3599 599 3657 633
rect 3691 599 3749 633
rect 3783 599 3841 633
rect 3875 599 3933 633
rect 3967 599 4025 633
rect 4059 599 4117 633
rect 4151 599 4209 633
rect 4243 599 4301 633
rect 4335 599 4393 633
rect 4427 599 4485 633
rect 4519 599 4577 633
rect 4611 599 4640 633
rect 149 528 207 599
rect 149 494 161 528
rect 195 494 207 528
rect 149 435 207 494
rect 149 401 161 435
rect 195 401 207 435
rect 149 366 207 401
rect 292 557 334 599
rect 292 523 300 557
rect 292 489 334 523
rect 292 455 300 489
rect 292 421 334 455
rect 292 387 300 421
rect 292 371 334 387
rect 368 557 434 565
rect 368 523 384 557
rect 418 523 434 557
rect 368 489 434 523
rect 368 455 384 489
rect 418 455 434 489
rect 368 421 434 455
rect 535 549 569 565
rect 535 481 569 515
rect 603 533 669 599
rect 603 499 619 533
rect 653 499 669 533
rect 703 549 740 565
rect 737 515 740 549
rect 703 481 740 515
rect 788 557 841 599
rect 788 523 807 557
rect 788 507 841 523
rect 875 549 925 565
rect 875 515 891 549
rect 1222 557 1256 599
rect 569 463 668 465
rect 569 447 626 463
rect 535 431 626 447
rect 368 387 384 421
rect 418 387 434 421
rect 622 429 626 431
rect 660 429 668 463
rect 368 369 434 387
rect 336 321 354 335
rect 288 287 304 288
rect 338 287 354 321
rect 288 237 334 253
rect 388 249 434 369
rect 518 376 588 397
rect 518 328 520 376
rect 568 328 588 376
rect 518 321 588 328
rect 518 287 532 321
rect 566 287 588 321
rect 518 267 588 287
rect 622 336 668 429
rect 622 302 634 336
rect 149 217 207 234
rect 149 183 161 217
rect 195 183 207 217
rect 149 89 207 183
rect 288 203 300 237
rect 288 169 334 203
rect 288 135 300 169
rect 288 89 334 135
rect 368 242 434 249
rect 368 194 384 242
rect 432 194 434 242
rect 622 233 668 302
rect 368 169 434 194
rect 368 135 384 169
rect 418 135 434 169
rect 535 199 668 233
rect 737 447 740 481
rect 875 480 925 515
rect 967 510 983 544
rect 1017 510 1188 544
rect 703 395 740 447
rect 864 454 925 480
rect 1014 463 1120 476
rect 703 361 705 395
rect 739 361 740 395
rect 535 191 569 199
rect 703 191 740 361
rect 774 389 830 405
rect 774 355 796 389
rect 774 292 830 355
rect 774 244 780 292
rect 828 244 830 292
rect 774 215 830 244
rect 864 233 898 454
rect 1014 429 1046 463
rect 1080 437 1120 463
rect 932 395 980 416
rect 932 361 943 395
rect 977 361 980 395
rect 932 359 980 361
rect 932 325 939 359
rect 973 325 980 359
rect 932 297 980 325
rect 1014 263 1048 429
rect 1082 403 1120 437
rect 1154 387 1188 510
rect 1222 489 1256 523
rect 1222 439 1256 455
rect 1290 549 1340 565
rect 1290 515 1306 549
rect 1598 549 1661 599
rect 1290 499 1340 515
rect 1385 505 1401 539
rect 1435 505 1562 539
rect 1154 371 1256 387
rect 1154 369 1222 371
rect 864 207 909 233
rect 943 229 959 263
rect 993 229 1048 263
rect 943 219 1048 229
rect 1082 337 1222 369
rect 1082 335 1256 337
rect 535 141 569 157
rect 368 123 434 135
rect 603 131 619 165
rect 653 131 669 165
rect 737 157 740 191
rect 703 141 740 157
rect 791 165 841 181
rect 603 89 669 131
rect 791 131 807 165
rect 875 179 909 207
rect 1082 179 1116 335
rect 1222 321 1256 335
rect 1158 285 1198 291
rect 1290 285 1324 499
rect 1358 463 1396 465
rect 1358 429 1360 463
rect 1394 429 1396 463
rect 1358 371 1396 429
rect 1392 337 1396 371
rect 1358 321 1396 337
rect 1430 437 1494 471
rect 1430 403 1460 437
rect 1430 395 1494 403
rect 1430 361 1447 395
rect 1481 361 1494 395
rect 1158 275 1324 285
rect 1430 279 1494 361
rect 1192 241 1324 275
rect 1158 225 1324 241
rect 875 145 892 179
rect 926 145 942 179
rect 981 145 1003 179
rect 1037 145 1116 179
rect 1180 173 1254 189
rect 791 89 841 131
rect 1180 139 1202 173
rect 1236 139 1254 173
rect 1290 179 1324 225
rect 1401 263 1494 279
rect 1435 229 1494 263
rect 1401 213 1494 229
rect 1528 337 1562 505
rect 1598 515 1600 549
rect 1634 515 1661 549
rect 1598 499 1661 515
rect 1708 557 1776 565
rect 1708 523 1724 557
rect 1758 523 1776 557
rect 1708 486 1776 523
rect 1708 453 1724 486
rect 1596 452 1724 453
rect 1758 452 1776 486
rect 1596 437 1776 452
rect 1630 415 1776 437
rect 1630 403 1724 415
rect 1596 381 1724 403
rect 1758 381 1776 415
rect 1810 527 1844 599
rect 1982 557 2048 561
rect 1810 447 1844 493
rect 1810 397 1844 413
rect 1878 551 1944 556
rect 1878 517 1894 551
rect 1928 517 1944 551
rect 1878 483 1944 517
rect 1878 449 1894 483
rect 1928 449 1944 483
rect 1878 415 1944 449
rect 1982 523 1998 557
rect 2032 523 2048 557
rect 1982 489 2048 523
rect 1982 455 1998 489
rect 2032 455 2048 489
rect 1982 415 2048 455
rect 1596 378 1776 381
rect 1738 337 1776 378
rect 1878 381 1894 415
rect 1928 387 1944 415
rect 1928 381 1960 387
rect 1878 371 1960 381
rect 1913 361 1960 371
rect 1528 321 1704 337
rect 1528 287 1670 321
rect 1528 271 1704 287
rect 1738 321 1888 337
rect 1738 287 1854 321
rect 1738 271 1888 287
rect 1528 179 1562 271
rect 1738 237 1778 271
rect 1922 245 1960 361
rect 1911 237 1960 245
rect 1712 234 1778 237
rect 1712 200 1728 234
rect 1762 200 1778 234
rect 1880 236 1960 237
rect 1880 230 1896 236
rect 1930 230 1960 236
rect 1290 145 1321 179
rect 1355 145 1371 179
rect 1405 145 1424 179
rect 1458 145 1562 179
rect 1617 179 1659 195
rect 1617 145 1622 179
rect 1656 145 1659 179
rect 1180 89 1254 139
rect 1617 89 1659 145
rect 1712 166 1778 200
rect 1712 132 1728 166
rect 1762 132 1778 166
rect 1812 195 1846 211
rect 1812 89 1846 161
rect 1880 182 1886 230
rect 1934 220 1960 230
rect 1994 337 2048 415
rect 2086 557 2129 599
rect 2086 523 2095 557
rect 2086 489 2129 523
rect 2086 455 2095 489
rect 2086 421 2129 455
rect 2086 387 2095 421
rect 2086 371 2129 387
rect 2163 557 2230 565
rect 2163 523 2179 557
rect 2213 523 2230 557
rect 2163 486 2230 523
rect 2163 452 2179 486
rect 2213 452 2230 486
rect 2163 415 2230 452
rect 2283 549 2317 565
rect 2283 481 2317 515
rect 2351 533 2417 599
rect 2351 499 2367 533
rect 2401 499 2417 533
rect 2451 549 2488 565
rect 2485 515 2488 549
rect 2451 481 2488 515
rect 2536 557 2589 599
rect 2536 523 2555 557
rect 2536 507 2589 523
rect 2623 549 2673 565
rect 2623 515 2639 549
rect 2970 557 3004 599
rect 2317 463 2416 465
rect 2317 447 2374 463
rect 2283 431 2374 447
rect 2163 381 2179 415
rect 2213 381 2230 415
rect 2370 429 2374 431
rect 2408 429 2416 463
rect 2163 368 2230 381
rect 1994 321 2149 337
rect 1994 287 2115 321
rect 1994 271 2149 287
rect 1934 182 1946 220
rect 1994 195 2034 271
rect 2183 254 2230 368
rect 2266 384 2336 397
rect 2266 336 2274 384
rect 2322 336 2336 384
rect 2266 321 2336 336
rect 2266 287 2280 321
rect 2314 287 2336 321
rect 2266 267 2336 287
rect 2370 336 2416 429
rect 2370 302 2382 336
rect 1880 168 1946 182
rect 1880 134 1896 168
rect 1930 134 1946 168
rect 1984 191 2034 195
rect 1984 157 2000 191
rect 2179 203 2230 254
rect 2370 233 2416 302
rect 1984 141 2034 157
rect 2081 165 2145 181
rect 1880 133 1946 134
rect 2081 131 2095 165
rect 2129 131 2145 165
rect 2081 89 2145 131
rect 2213 169 2230 203
rect 2179 123 2230 169
rect 2283 199 2416 233
rect 2485 447 2488 481
rect 2623 480 2673 515
rect 2715 510 2731 544
rect 2765 510 2936 544
rect 2451 395 2488 447
rect 2612 454 2673 480
rect 2762 463 2868 476
rect 2451 361 2453 395
rect 2487 361 2488 395
rect 2283 191 2317 199
rect 2451 191 2488 361
rect 2522 389 2578 405
rect 2522 355 2544 389
rect 2522 280 2578 355
rect 2522 232 2526 280
rect 2574 232 2578 280
rect 2522 215 2578 232
rect 2612 233 2646 454
rect 2762 429 2794 463
rect 2828 437 2868 463
rect 2680 395 2728 416
rect 2680 361 2691 395
rect 2725 361 2728 395
rect 2680 359 2728 361
rect 2680 325 2687 359
rect 2721 325 2728 359
rect 2680 297 2728 325
rect 2762 263 2796 429
rect 2830 403 2868 437
rect 2902 387 2936 510
rect 2970 489 3004 523
rect 2970 439 3004 455
rect 3038 549 3088 565
rect 3038 515 3054 549
rect 3346 549 3409 599
rect 3038 499 3088 515
rect 3133 505 3149 539
rect 3183 505 3310 539
rect 2902 371 3004 387
rect 2902 369 2970 371
rect 2612 207 2657 233
rect 2691 229 2707 263
rect 2741 229 2796 263
rect 2691 219 2796 229
rect 2830 337 2970 369
rect 2830 335 3004 337
rect 2283 141 2317 157
rect 2351 131 2367 165
rect 2401 131 2417 165
rect 2485 157 2488 191
rect 2451 141 2488 157
rect 2539 165 2589 181
rect 2351 89 2417 131
rect 2539 131 2555 165
rect 2623 179 2657 207
rect 2830 179 2864 335
rect 2970 321 3004 335
rect 2906 285 2946 291
rect 3038 285 3072 499
rect 3106 463 3144 465
rect 3106 429 3108 463
rect 3142 429 3144 463
rect 3106 371 3144 429
rect 3140 337 3144 371
rect 3106 321 3144 337
rect 3178 437 3242 471
rect 3178 403 3208 437
rect 3178 395 3242 403
rect 3178 361 3195 395
rect 3229 361 3242 395
rect 2906 275 3072 285
rect 3178 279 3242 361
rect 2940 241 3072 275
rect 2906 225 3072 241
rect 2623 145 2640 179
rect 2674 145 2690 179
rect 2729 145 2751 179
rect 2785 145 2864 179
rect 2928 173 3002 189
rect 2539 89 2589 131
rect 2928 139 2950 173
rect 2984 139 3002 173
rect 3038 179 3072 225
rect 3149 263 3242 279
rect 3183 229 3242 263
rect 3149 213 3242 229
rect 3276 337 3310 505
rect 3346 515 3348 549
rect 3382 515 3409 549
rect 3346 499 3409 515
rect 3456 557 3524 565
rect 3456 523 3472 557
rect 3506 523 3524 557
rect 3456 486 3524 523
rect 3456 453 3472 486
rect 3344 452 3472 453
rect 3506 452 3524 486
rect 3344 437 3524 452
rect 3378 415 3524 437
rect 3378 403 3472 415
rect 3344 381 3472 403
rect 3506 381 3524 415
rect 3558 527 3592 599
rect 3730 557 3796 561
rect 3558 447 3592 493
rect 3558 397 3592 413
rect 3626 551 3692 556
rect 3626 517 3642 551
rect 3676 517 3692 551
rect 3626 483 3692 517
rect 3626 449 3642 483
rect 3676 449 3692 483
rect 3626 415 3692 449
rect 3730 523 3746 557
rect 3780 523 3796 557
rect 3730 489 3796 523
rect 3730 455 3746 489
rect 3780 455 3796 489
rect 3730 415 3796 455
rect 3344 378 3524 381
rect 3486 337 3524 378
rect 3626 381 3642 415
rect 3676 387 3692 415
rect 3676 381 3708 387
rect 3626 371 3708 381
rect 3661 361 3708 371
rect 3276 321 3452 337
rect 3276 287 3418 321
rect 3276 271 3452 287
rect 3486 321 3636 337
rect 3486 287 3602 321
rect 3486 271 3636 287
rect 3276 179 3310 271
rect 3486 237 3526 271
rect 3670 245 3708 361
rect 3659 237 3708 245
rect 3460 234 3526 237
rect 3460 200 3476 234
rect 3510 200 3526 234
rect 3628 236 3708 237
rect 3628 230 3644 236
rect 3678 230 3708 236
rect 3038 145 3069 179
rect 3103 145 3119 179
rect 3153 145 3172 179
rect 3206 145 3310 179
rect 3365 179 3407 195
rect 3365 145 3370 179
rect 3404 145 3407 179
rect 2928 89 3002 139
rect 3365 89 3407 145
rect 3460 166 3526 200
rect 3460 132 3476 166
rect 3510 132 3526 166
rect 3560 195 3594 211
rect 3560 89 3594 161
rect 3628 182 3634 230
rect 3682 220 3708 230
rect 3742 337 3796 415
rect 3834 557 3877 599
rect 3834 523 3843 557
rect 3834 489 3877 523
rect 3834 455 3843 489
rect 3834 421 3877 455
rect 3834 387 3843 421
rect 3834 371 3877 387
rect 3911 557 3978 565
rect 3911 523 3927 557
rect 3961 523 3978 557
rect 3911 486 3978 523
rect 3911 452 3927 486
rect 3961 452 3978 486
rect 3911 415 3978 452
rect 3911 381 3927 415
rect 3961 381 3978 415
rect 3911 368 3978 381
rect 4013 557 4065 599
rect 4013 523 4031 557
rect 4013 489 4065 523
rect 4013 455 4031 489
rect 4013 421 4065 455
rect 4013 387 4031 421
rect 4013 371 4065 387
rect 4099 557 4165 565
rect 4099 523 4115 557
rect 4149 523 4165 557
rect 4099 489 4165 523
rect 4099 460 4115 489
rect 4149 460 4165 489
rect 4099 412 4104 460
rect 4152 412 4165 460
rect 4099 387 4115 412
rect 4149 387 4165 412
rect 4099 369 4165 387
rect 4199 557 4255 599
rect 4233 523 4255 557
rect 4199 489 4255 523
rect 4233 455 4255 489
rect 4199 421 4255 455
rect 4233 387 4255 421
rect 4199 371 4255 387
rect 4340 557 4382 599
rect 4340 523 4348 557
rect 4340 489 4382 523
rect 4340 455 4348 489
rect 4340 421 4382 455
rect 4340 387 4348 421
rect 4340 371 4382 387
rect 4416 557 4482 565
rect 4416 523 4432 557
rect 4466 523 4482 557
rect 4416 489 4482 523
rect 4416 455 4432 489
rect 4466 455 4482 489
rect 4416 421 4482 455
rect 4416 387 4432 421
rect 4466 387 4482 421
rect 4416 369 4482 387
rect 3742 321 3897 337
rect 3742 287 3863 321
rect 3742 271 3897 287
rect 3682 182 3694 220
rect 3742 195 3782 271
rect 3931 254 3978 368
rect 4017 332 4084 337
rect 4017 287 4026 332
rect 4074 287 4084 332
rect 3628 168 3694 182
rect 3628 134 3644 168
rect 3678 134 3694 168
rect 3732 191 3782 195
rect 3732 157 3748 191
rect 3927 203 3978 254
rect 4118 249 4152 369
rect 4186 332 4253 337
rect 4186 284 4198 332
rect 4246 284 4253 332
rect 4336 288 4340 335
rect 4388 288 4402 335
rect 4336 287 4352 288
rect 4386 287 4402 288
rect 4436 332 4482 369
rect 4565 528 4623 599
rect 4565 494 4577 528
rect 4611 494 4623 528
rect 4565 435 4623 494
rect 4565 401 4577 435
rect 4611 401 4623 435
rect 4565 366 4623 401
rect 4186 283 4253 284
rect 4436 284 4442 332
rect 3732 141 3782 157
rect 3829 165 3893 181
rect 3628 133 3694 134
rect 3829 131 3843 165
rect 3877 131 3893 165
rect 3829 89 3893 131
rect 3961 169 3978 203
rect 3927 123 3978 169
rect 4013 233 4152 249
rect 4013 199 4031 233
rect 4065 199 4152 233
rect 4013 165 4152 199
rect 4013 131 4031 165
rect 4065 131 4152 165
rect 4013 123 4152 131
rect 4193 233 4255 249
rect 4193 199 4199 233
rect 4233 199 4255 233
rect 4193 165 4255 199
rect 4193 131 4199 165
rect 4233 131 4255 165
rect 4193 89 4255 131
rect 4336 237 4382 253
rect 4436 249 4482 284
rect 4336 203 4348 237
rect 4336 169 4382 203
rect 4336 135 4348 169
rect 4336 89 4382 135
rect 4416 237 4482 249
rect 4416 203 4432 237
rect 4466 203 4482 237
rect 4416 169 4482 203
rect 4416 135 4432 169
rect 4466 135 4482 169
rect 4416 123 4482 135
rect 4565 217 4623 234
rect 4565 183 4577 217
rect 4611 183 4623 217
rect 4565 89 4623 183
rect 132 55 161 89
rect 195 55 253 89
rect 287 55 345 89
rect 379 55 437 89
rect 471 55 529 89
rect 563 55 621 89
rect 655 55 713 89
rect 747 55 805 89
rect 839 55 897 89
rect 931 55 989 89
rect 1023 55 1081 89
rect 1115 55 1173 89
rect 1207 55 1265 89
rect 1299 55 1357 89
rect 1391 55 1449 89
rect 1483 55 1541 89
rect 1575 55 1633 89
rect 1667 55 1725 89
rect 1759 55 1817 89
rect 1851 55 1909 89
rect 1943 55 2001 89
rect 2035 55 2093 89
rect 2127 55 2185 89
rect 2219 55 2277 89
rect 2311 55 2369 89
rect 2403 55 2461 89
rect 2495 55 2553 89
rect 2587 55 2645 89
rect 2679 55 2737 89
rect 2771 55 2829 89
rect 2863 55 2921 89
rect 2955 55 3013 89
rect 3047 55 3105 89
rect 3139 55 3197 89
rect 3231 55 3289 89
rect 3323 55 3381 89
rect 3415 55 3473 89
rect 3507 55 3565 89
rect 3599 55 3657 89
rect 3691 55 3749 89
rect 3783 55 3841 89
rect 3875 55 3933 89
rect 3967 55 4025 89
rect 4059 55 4117 89
rect 4151 55 4209 89
rect 4243 55 4301 89
rect 4335 55 4393 89
rect 4427 55 4485 89
rect 4519 55 4577 89
rect 4611 55 4640 89
rect 425 -39 483 55
rect 603 13 669 55
rect 425 -73 437 -39
rect 471 -73 483 -39
rect 425 -90 483 -73
rect 535 -13 569 3
rect 603 -21 619 13
rect 653 -21 669 13
rect 791 13 841 55
rect 703 -13 740 3
rect 535 -55 569 -47
rect 737 -47 740 -13
rect 791 -21 807 13
rect 1180 5 1254 55
rect 791 -37 841 -21
rect 875 -35 892 -1
rect 926 -35 942 -1
rect 981 -35 1003 -1
rect 1037 -35 1116 -1
rect 535 -89 668 -55
rect 518 -138 588 -123
rect 518 -186 520 -138
rect 568 -186 588 -138
rect 425 -257 483 -222
rect 518 -253 588 -186
rect 622 -158 668 -89
rect 622 -192 634 -158
rect 425 -291 437 -257
rect 471 -291 483 -257
rect 622 -285 668 -192
rect 622 -287 626 -285
rect 425 -350 483 -291
rect 425 -384 437 -350
rect 471 -384 483 -350
rect 425 -455 483 -384
rect 535 -303 626 -287
rect 569 -319 626 -303
rect 660 -319 668 -285
rect 569 -321 668 -319
rect 703 -217 740 -47
rect 875 -63 909 -35
rect 703 -251 705 -217
rect 739 -251 740 -217
rect 703 -303 740 -251
rect 774 -78 830 -71
rect 774 -126 780 -78
rect 828 -126 830 -78
rect 774 -211 830 -126
rect 774 -245 796 -211
rect 774 -261 830 -245
rect 864 -89 909 -63
rect 943 -85 1048 -75
rect 535 -371 569 -337
rect 737 -337 740 -303
rect 864 -310 898 -89
rect 943 -119 959 -85
rect 993 -119 1048 -85
rect 932 -181 980 -153
rect 932 -215 939 -181
rect 973 -215 980 -181
rect 932 -217 980 -215
rect 932 -251 943 -217
rect 977 -251 980 -217
rect 932 -272 980 -251
rect 1014 -285 1048 -119
rect 1082 -191 1116 -35
rect 1180 -29 1202 5
rect 1236 -29 1254 5
rect 1617 -1 1659 55
rect 1180 -45 1254 -29
rect 1290 -35 1321 -1
rect 1355 -35 1371 -1
rect 1405 -35 1424 -1
rect 1458 -35 1562 -1
rect 1290 -81 1324 -35
rect 1158 -97 1324 -81
rect 1192 -131 1324 -97
rect 1158 -141 1324 -131
rect 1401 -85 1494 -69
rect 1435 -119 1494 -85
rect 1401 -135 1494 -119
rect 1158 -147 1198 -141
rect 1222 -191 1256 -177
rect 1082 -193 1256 -191
rect 1082 -225 1222 -193
rect 1154 -227 1222 -225
rect 1154 -243 1256 -227
rect 864 -336 925 -310
rect 1014 -319 1046 -285
rect 1082 -293 1120 -259
rect 1080 -319 1120 -293
rect 1014 -332 1120 -319
rect 535 -421 569 -405
rect 603 -389 619 -355
rect 653 -389 669 -355
rect 603 -455 669 -389
rect 703 -371 740 -337
rect 737 -405 740 -371
rect 703 -421 740 -405
rect 788 -379 841 -363
rect 788 -413 807 -379
rect 788 -455 841 -413
rect 875 -371 925 -336
rect 1154 -366 1188 -243
rect 875 -405 891 -371
rect 967 -400 983 -366
rect 1017 -400 1188 -366
rect 1222 -311 1256 -295
rect 1222 -379 1256 -345
rect 875 -421 925 -405
rect 1222 -455 1256 -413
rect 1290 -355 1324 -141
rect 1358 -193 1396 -177
rect 1392 -227 1396 -193
rect 1358 -285 1396 -227
rect 1358 -319 1360 -285
rect 1394 -319 1396 -285
rect 1358 -321 1396 -319
rect 1430 -217 1494 -135
rect 1430 -251 1447 -217
rect 1481 -251 1494 -217
rect 1430 -259 1494 -251
rect 1430 -293 1460 -259
rect 1430 -327 1494 -293
rect 1528 -127 1562 -35
rect 1617 -35 1622 -1
rect 1656 -35 1659 -1
rect 1617 -51 1659 -35
rect 1712 -22 1728 12
rect 1762 -22 1778 12
rect 1712 -56 1778 -22
rect 1712 -90 1728 -56
rect 1762 -90 1778 -56
rect 1812 -17 1846 55
rect 2081 13 2145 55
rect 1812 -67 1846 -51
rect 1880 10 1946 11
rect 1880 -24 1896 10
rect 1930 -24 1946 10
rect 1880 -58 1946 -24
rect 1984 -13 2034 3
rect 1984 -47 2000 -13
rect 2081 -21 2095 13
rect 2129 -21 2145 13
rect 2081 -37 2145 -21
rect 2179 -25 2230 21
rect 2351 13 2417 55
rect 2213 -30 2230 -25
rect 2283 -13 2317 3
rect 1984 -51 2034 -47
rect 1712 -93 1778 -90
rect 1880 -92 1896 -58
rect 1930 -76 1946 -58
rect 1930 -92 1960 -76
rect 1880 -93 1960 -92
rect 1738 -127 1778 -93
rect 1911 -101 1960 -93
rect 1528 -143 1704 -127
rect 1528 -177 1670 -143
rect 1528 -193 1704 -177
rect 1738 -143 1888 -127
rect 1738 -177 1854 -143
rect 1738 -193 1888 -177
rect 1290 -371 1340 -355
rect 1528 -361 1562 -193
rect 1738 -234 1776 -193
rect 1922 -217 1960 -101
rect 1913 -227 1960 -217
rect 1596 -237 1776 -234
rect 1596 -259 1724 -237
rect 1630 -271 1724 -259
rect 1758 -271 1776 -237
rect 1878 -237 1960 -227
rect 1630 -293 1776 -271
rect 1596 -308 1776 -293
rect 1596 -309 1724 -308
rect 1708 -342 1724 -309
rect 1758 -342 1776 -308
rect 1290 -405 1306 -371
rect 1385 -395 1401 -361
rect 1435 -395 1562 -361
rect 1598 -371 1661 -355
rect 1290 -421 1340 -405
rect 1598 -405 1600 -371
rect 1634 -405 1661 -371
rect 1598 -455 1661 -405
rect 1708 -379 1776 -342
rect 1708 -413 1724 -379
rect 1758 -413 1776 -379
rect 1708 -421 1776 -413
rect 1810 -269 1844 -253
rect 1810 -349 1844 -303
rect 1810 -455 1844 -383
rect 1878 -271 1894 -237
rect 1928 -243 1960 -237
rect 1994 -127 2034 -51
rect 2179 -78 2186 -59
rect 2351 -21 2367 13
rect 2401 -21 2417 13
rect 2539 13 2589 55
rect 2451 -13 2488 3
rect 2283 -55 2317 -47
rect 2485 -47 2488 -13
rect 2539 -21 2555 13
rect 2928 5 3002 55
rect 2539 -37 2589 -21
rect 2623 -35 2640 -1
rect 2674 -35 2690 -1
rect 2729 -35 2751 -1
rect 2785 -35 2864 -1
rect 2179 -110 2230 -78
rect 2283 -89 2416 -55
rect 1994 -143 2149 -127
rect 1994 -177 2115 -143
rect 1994 -193 2149 -177
rect 1928 -271 1944 -243
rect 1994 -271 2048 -193
rect 2183 -224 2230 -110
rect 1878 -305 1944 -271
rect 1878 -339 1894 -305
rect 1928 -339 1944 -305
rect 1878 -373 1944 -339
rect 1878 -407 1894 -373
rect 1928 -407 1944 -373
rect 1878 -412 1944 -407
rect 1982 -311 2048 -271
rect 1982 -345 1998 -311
rect 2032 -345 2048 -311
rect 1982 -379 2048 -345
rect 1982 -413 1998 -379
rect 2032 -413 2048 -379
rect 1982 -417 2048 -413
rect 2086 -243 2129 -227
rect 2086 -277 2095 -243
rect 2086 -311 2129 -277
rect 2086 -345 2095 -311
rect 2086 -379 2129 -345
rect 2086 -413 2095 -379
rect 2086 -455 2129 -413
rect 2163 -237 2230 -224
rect 2163 -271 2179 -237
rect 2213 -271 2230 -237
rect 2266 -142 2336 -123
rect 2266 -190 2280 -142
rect 2328 -190 2336 -142
rect 2266 -253 2336 -190
rect 2370 -158 2416 -89
rect 2370 -192 2382 -158
rect 2163 -308 2230 -271
rect 2370 -285 2416 -192
rect 2370 -287 2374 -285
rect 2163 -342 2179 -308
rect 2213 -342 2230 -308
rect 2163 -379 2230 -342
rect 2163 -413 2179 -379
rect 2213 -413 2230 -379
rect 2163 -421 2230 -413
rect 2283 -303 2374 -287
rect 2317 -319 2374 -303
rect 2408 -319 2416 -285
rect 2317 -321 2416 -319
rect 2451 -217 2488 -47
rect 2623 -63 2657 -35
rect 2451 -251 2453 -217
rect 2487 -251 2488 -217
rect 2451 -303 2488 -251
rect 2522 -84 2578 -71
rect 2522 -132 2526 -84
rect 2574 -132 2578 -84
rect 2522 -211 2578 -132
rect 2522 -245 2544 -211
rect 2522 -261 2578 -245
rect 2612 -89 2657 -63
rect 2691 -85 2796 -75
rect 2283 -371 2317 -337
rect 2485 -337 2488 -303
rect 2612 -310 2646 -89
rect 2691 -119 2707 -85
rect 2741 -119 2796 -85
rect 2680 -181 2728 -153
rect 2680 -215 2687 -181
rect 2721 -215 2728 -181
rect 2680 -217 2728 -215
rect 2680 -251 2691 -217
rect 2725 -251 2728 -217
rect 2680 -272 2728 -251
rect 2762 -285 2796 -119
rect 2830 -191 2864 -35
rect 2928 -29 2950 5
rect 2984 -29 3002 5
rect 3365 -1 3407 55
rect 2928 -45 3002 -29
rect 3038 -35 3069 -1
rect 3103 -35 3119 -1
rect 3153 -35 3172 -1
rect 3206 -35 3310 -1
rect 3038 -81 3072 -35
rect 2906 -97 3072 -81
rect 2940 -131 3072 -97
rect 2906 -141 3072 -131
rect 3149 -85 3242 -69
rect 3183 -119 3242 -85
rect 3149 -135 3242 -119
rect 2906 -147 2946 -141
rect 2970 -191 3004 -177
rect 2830 -193 3004 -191
rect 2830 -225 2970 -193
rect 2902 -227 2970 -225
rect 2902 -243 3004 -227
rect 2612 -336 2673 -310
rect 2762 -319 2794 -285
rect 2830 -293 2868 -259
rect 2828 -319 2868 -293
rect 2762 -332 2868 -319
rect 2283 -421 2317 -405
rect 2351 -389 2367 -355
rect 2401 -389 2417 -355
rect 2351 -455 2417 -389
rect 2451 -371 2488 -337
rect 2485 -405 2488 -371
rect 2451 -421 2488 -405
rect 2536 -379 2589 -363
rect 2536 -413 2555 -379
rect 2536 -455 2589 -413
rect 2623 -371 2673 -336
rect 2902 -366 2936 -243
rect 2623 -405 2639 -371
rect 2715 -400 2731 -366
rect 2765 -400 2936 -366
rect 2970 -311 3004 -295
rect 2970 -379 3004 -345
rect 2623 -421 2673 -405
rect 2970 -455 3004 -413
rect 3038 -355 3072 -141
rect 3106 -193 3144 -177
rect 3140 -227 3144 -193
rect 3106 -285 3144 -227
rect 3106 -319 3108 -285
rect 3142 -319 3144 -285
rect 3106 -321 3144 -319
rect 3178 -217 3242 -135
rect 3178 -251 3195 -217
rect 3229 -251 3242 -217
rect 3178 -259 3242 -251
rect 3178 -293 3208 -259
rect 3178 -327 3242 -293
rect 3276 -127 3310 -35
rect 3365 -35 3370 -1
rect 3404 -35 3407 -1
rect 3365 -51 3407 -35
rect 3460 -22 3476 12
rect 3510 -22 3526 12
rect 3460 -56 3526 -22
rect 3460 -90 3476 -56
rect 3510 -90 3526 -56
rect 3560 -17 3594 55
rect 3829 13 3893 55
rect 3560 -67 3594 -51
rect 3628 10 3694 11
rect 3628 -24 3644 10
rect 3678 -24 3694 10
rect 3628 -34 3694 -24
rect 3460 -93 3526 -90
rect 3628 -82 3636 -34
rect 3684 -76 3694 -34
rect 3732 -13 3782 3
rect 3732 -47 3748 -13
rect 3829 -21 3843 13
rect 3877 -21 3893 13
rect 3829 -37 3893 -21
rect 3927 -25 3978 21
rect 3732 -51 3782 -47
rect 3684 -82 3708 -76
rect 3628 -92 3644 -82
rect 3678 -92 3708 -82
rect 3628 -93 3708 -92
rect 3486 -127 3526 -93
rect 3659 -101 3708 -93
rect 3276 -143 3452 -127
rect 3276 -177 3418 -143
rect 3276 -193 3452 -177
rect 3486 -143 3636 -127
rect 3486 -177 3602 -143
rect 3486 -193 3636 -177
rect 3038 -371 3088 -355
rect 3276 -361 3310 -193
rect 3486 -234 3524 -193
rect 3670 -217 3708 -101
rect 3661 -227 3708 -217
rect 3344 -237 3524 -234
rect 3344 -259 3472 -237
rect 3378 -271 3472 -259
rect 3506 -271 3524 -237
rect 3626 -237 3708 -227
rect 3378 -293 3524 -271
rect 3344 -308 3524 -293
rect 3344 -309 3472 -308
rect 3456 -342 3472 -309
rect 3506 -342 3524 -308
rect 3038 -405 3054 -371
rect 3133 -395 3149 -361
rect 3183 -395 3310 -361
rect 3346 -371 3409 -355
rect 3038 -421 3088 -405
rect 3346 -405 3348 -371
rect 3382 -405 3409 -371
rect 3346 -455 3409 -405
rect 3456 -379 3524 -342
rect 3456 -413 3472 -379
rect 3506 -413 3524 -379
rect 3456 -421 3524 -413
rect 3558 -269 3592 -253
rect 3558 -349 3592 -303
rect 3558 -455 3592 -383
rect 3626 -271 3642 -237
rect 3676 -243 3708 -237
rect 3742 -127 3782 -51
rect 3961 -59 3978 -25
rect 3927 -110 3978 -59
rect 4013 -39 4071 55
rect 4013 -73 4025 -39
rect 4059 -73 4071 -39
rect 4013 -90 4071 -73
rect 3742 -143 3897 -127
rect 3742 -177 3863 -143
rect 3742 -193 3897 -177
rect 3676 -271 3692 -243
rect 3742 -271 3796 -193
rect 3931 -224 3978 -110
rect 3626 -305 3692 -271
rect 3626 -339 3642 -305
rect 3676 -339 3692 -305
rect 3626 -373 3692 -339
rect 3626 -407 3642 -373
rect 3676 -407 3692 -373
rect 3626 -412 3692 -407
rect 3730 -311 3796 -271
rect 3730 -345 3746 -311
rect 3780 -345 3796 -311
rect 3730 -379 3796 -345
rect 3730 -413 3746 -379
rect 3780 -413 3796 -379
rect 3730 -417 3796 -413
rect 3834 -243 3877 -227
rect 3834 -277 3843 -243
rect 3834 -311 3877 -277
rect 3834 -345 3843 -311
rect 3834 -379 3877 -345
rect 3834 -413 3843 -379
rect 3834 -455 3877 -413
rect 3911 -237 3978 -224
rect 3911 -271 3927 -237
rect 3961 -271 3978 -237
rect 3911 -308 3978 -271
rect 3911 -342 3927 -308
rect 3961 -342 3978 -308
rect 3911 -379 3978 -342
rect 3911 -413 3927 -379
rect 3961 -413 3978 -379
rect 3911 -421 3978 -413
rect 4013 -257 4071 -222
rect 4013 -291 4025 -257
rect 4059 -291 4071 -257
rect 4013 -350 4071 -291
rect 4013 -384 4025 -350
rect 4059 -384 4071 -350
rect 4013 -455 4071 -384
rect 408 -489 437 -455
rect 471 -489 529 -455
rect 563 -489 621 -455
rect 655 -489 713 -455
rect 747 -489 805 -455
rect 839 -489 897 -455
rect 931 -489 989 -455
rect 1023 -489 1081 -455
rect 1115 -489 1173 -455
rect 1207 -489 1265 -455
rect 1299 -489 1357 -455
rect 1391 -489 1449 -455
rect 1483 -489 1541 -455
rect 1575 -489 1633 -455
rect 1667 -489 1725 -455
rect 1759 -489 1817 -455
rect 1851 -489 1909 -455
rect 1943 -489 2001 -455
rect 2035 -489 2093 -455
rect 2127 -489 2185 -455
rect 2219 -489 2277 -455
rect 2311 -489 2369 -455
rect 2403 -489 2461 -455
rect 2495 -489 2553 -455
rect 2587 -489 2645 -455
rect 2679 -489 2737 -455
rect 2771 -489 2829 -455
rect 2863 -489 2921 -455
rect 2955 -489 3013 -455
rect 3047 -489 3105 -455
rect 3139 -489 3197 -455
rect 3231 -489 3289 -455
rect 3323 -489 3381 -455
rect 3415 -489 3473 -455
rect 3507 -489 3565 -455
rect 3599 -489 3657 -455
rect 3691 -489 3749 -455
rect 3783 -489 3841 -455
rect 3875 -489 3933 -455
rect 3967 -489 4025 -455
rect 4059 -489 4088 -455
<< viali >>
rect 161 599 195 633
rect 253 599 287 633
rect 345 599 379 633
rect 437 599 471 633
rect 529 599 563 633
rect 621 599 655 633
rect 713 599 747 633
rect 805 599 839 633
rect 897 599 931 633
rect 989 599 1023 633
rect 1081 599 1115 633
rect 1173 599 1207 633
rect 1265 599 1299 633
rect 1357 599 1391 633
rect 1449 599 1483 633
rect 1541 599 1575 633
rect 1633 599 1667 633
rect 1725 599 1759 633
rect 1817 599 1851 633
rect 1909 599 1943 633
rect 2001 599 2035 633
rect 2093 599 2127 633
rect 2185 599 2219 633
rect 2277 599 2311 633
rect 2369 599 2403 633
rect 2461 599 2495 633
rect 2553 599 2587 633
rect 2645 599 2679 633
rect 2737 599 2771 633
rect 2829 599 2863 633
rect 2921 599 2955 633
rect 3013 599 3047 633
rect 3105 599 3139 633
rect 3197 599 3231 633
rect 3289 599 3323 633
rect 3381 599 3415 633
rect 3473 599 3507 633
rect 3565 599 3599 633
rect 3657 599 3691 633
rect 3749 599 3783 633
rect 3841 599 3875 633
rect 3933 599 3967 633
rect 4025 599 4059 633
rect 4117 599 4151 633
rect 4209 599 4243 633
rect 4301 599 4335 633
rect 4393 599 4427 633
rect 4485 599 4519 633
rect 4577 599 4611 633
rect 626 429 660 463
rect 288 321 336 336
rect 288 288 304 321
rect 304 288 336 321
rect 520 328 568 376
rect 384 237 432 242
rect 384 203 418 237
rect 418 203 432 237
rect 384 194 432 203
rect 705 361 739 395
rect 780 244 828 292
rect 1046 437 1080 463
rect 1046 429 1048 437
rect 1048 429 1080 437
rect 943 361 977 395
rect 1360 429 1394 463
rect 1447 361 1481 395
rect 1886 202 1896 230
rect 1896 202 1930 230
rect 1930 202 1934 230
rect 2374 429 2408 463
rect 1886 182 1934 202
rect 2274 336 2322 384
rect 2453 361 2487 395
rect 2526 232 2574 280
rect 2794 437 2828 463
rect 2794 429 2796 437
rect 2796 429 2828 437
rect 2691 361 2725 395
rect 3108 429 3142 463
rect 3195 361 3229 395
rect 3634 202 3644 230
rect 3644 202 3678 230
rect 3678 202 3682 230
rect 4104 455 4115 460
rect 4115 455 4149 460
rect 4149 455 4152 460
rect 4104 421 4152 455
rect 4104 412 4115 421
rect 4115 412 4149 421
rect 4149 412 4152 421
rect 3634 182 3682 202
rect 4026 321 4074 332
rect 4026 287 4034 321
rect 4034 287 4068 321
rect 4068 287 4074 321
rect 4026 284 4074 287
rect 4198 321 4246 332
rect 4198 287 4202 321
rect 4202 287 4236 321
rect 4236 287 4246 321
rect 4198 284 4246 287
rect 4340 321 4388 336
rect 4340 288 4352 321
rect 4352 288 4386 321
rect 4386 288 4388 321
rect 4442 284 4490 332
rect 161 55 195 89
rect 253 55 287 89
rect 345 55 379 89
rect 437 55 471 89
rect 529 55 563 89
rect 621 55 655 89
rect 713 55 747 89
rect 805 55 839 89
rect 897 55 931 89
rect 989 55 1023 89
rect 1081 55 1115 89
rect 1173 55 1207 89
rect 1265 55 1299 89
rect 1357 55 1391 89
rect 1449 55 1483 89
rect 1541 55 1575 89
rect 1633 55 1667 89
rect 1725 55 1759 89
rect 1817 55 1851 89
rect 1909 55 1943 89
rect 2001 55 2035 89
rect 2093 55 2127 89
rect 2185 55 2219 89
rect 2277 55 2311 89
rect 2369 55 2403 89
rect 2461 55 2495 89
rect 2553 55 2587 89
rect 2645 55 2679 89
rect 2737 55 2771 89
rect 2829 55 2863 89
rect 2921 55 2955 89
rect 3013 55 3047 89
rect 3105 55 3139 89
rect 3197 55 3231 89
rect 3289 55 3323 89
rect 3381 55 3415 89
rect 3473 55 3507 89
rect 3565 55 3599 89
rect 3657 55 3691 89
rect 3749 55 3783 89
rect 3841 55 3875 89
rect 3933 55 3967 89
rect 4025 55 4059 89
rect 4117 55 4151 89
rect 4209 55 4243 89
rect 4301 55 4335 89
rect 4393 55 4427 89
rect 4485 55 4519 89
rect 4577 55 4611 89
rect 520 -143 568 -138
rect 520 -177 532 -143
rect 532 -177 566 -143
rect 566 -177 568 -143
rect 520 -186 568 -177
rect 626 -319 660 -285
rect 705 -251 739 -217
rect 780 -126 828 -78
rect 943 -251 977 -217
rect 1046 -293 1048 -285
rect 1048 -293 1080 -285
rect 1046 -319 1080 -293
rect 1360 -319 1394 -285
rect 1447 -251 1481 -217
rect 2186 -59 2213 -30
rect 2213 -59 2234 -30
rect 2186 -78 2234 -59
rect 2280 -143 2328 -142
rect 2280 -177 2314 -143
rect 2314 -177 2328 -143
rect 2280 -190 2328 -177
rect 2374 -319 2408 -285
rect 2453 -251 2487 -217
rect 2526 -132 2574 -84
rect 2691 -251 2725 -217
rect 2794 -293 2796 -285
rect 2796 -293 2828 -285
rect 2794 -319 2828 -293
rect 3108 -319 3142 -285
rect 3195 -251 3229 -217
rect 3636 -58 3684 -34
rect 3636 -82 3644 -58
rect 3644 -82 3678 -58
rect 3678 -82 3684 -58
rect 437 -489 471 -455
rect 529 -489 563 -455
rect 621 -489 655 -455
rect 713 -489 747 -455
rect 805 -489 839 -455
rect 897 -489 931 -455
rect 989 -489 1023 -455
rect 1081 -489 1115 -455
rect 1173 -489 1207 -455
rect 1265 -489 1299 -455
rect 1357 -489 1391 -455
rect 1449 -489 1483 -455
rect 1541 -489 1575 -455
rect 1633 -489 1667 -455
rect 1725 -489 1759 -455
rect 1817 -489 1851 -455
rect 1909 -489 1943 -455
rect 2001 -489 2035 -455
rect 2093 -489 2127 -455
rect 2185 -489 2219 -455
rect 2277 -489 2311 -455
rect 2369 -489 2403 -455
rect 2461 -489 2495 -455
rect 2553 -489 2587 -455
rect 2645 -489 2679 -455
rect 2737 -489 2771 -455
rect 2829 -489 2863 -455
rect 2921 -489 2955 -455
rect 3013 -489 3047 -455
rect 3105 -489 3139 -455
rect 3197 -489 3231 -455
rect 3289 -489 3323 -455
rect 3381 -489 3415 -455
rect 3473 -489 3507 -455
rect 3565 -489 3599 -455
rect 3657 -489 3691 -455
rect 3749 -489 3783 -455
rect 3841 -489 3875 -455
rect 3933 -489 3967 -455
rect 4025 -489 4059 -455
<< metal1 >>
rect -10 664 86 670
rect 86 633 4640 664
rect 86 599 161 633
rect 195 599 253 633
rect 287 599 345 633
rect 379 599 437 633
rect 471 599 529 633
rect 563 599 621 633
rect 655 599 713 633
rect 747 599 805 633
rect 839 599 897 633
rect 931 599 989 633
rect 1023 599 1081 633
rect 1115 599 1173 633
rect 1207 599 1265 633
rect 1299 599 1357 633
rect 1391 599 1449 633
rect 1483 599 1541 633
rect 1575 599 1633 633
rect 1667 599 1725 633
rect 1759 599 1817 633
rect 1851 599 1909 633
rect 1943 599 2001 633
rect 2035 599 2093 633
rect 2127 599 2185 633
rect 2219 599 2277 633
rect 2311 599 2369 633
rect 2403 599 2461 633
rect 2495 599 2553 633
rect 2587 599 2645 633
rect 2679 599 2737 633
rect 2771 599 2829 633
rect 2863 599 2921 633
rect 2955 599 3013 633
rect 3047 599 3105 633
rect 3139 599 3197 633
rect 3231 599 3289 633
rect 3323 599 3381 633
rect 3415 599 3473 633
rect 3507 599 3565 633
rect 3599 599 3657 633
rect 3691 599 3749 633
rect 3783 599 3841 633
rect 3875 599 3933 633
rect 3967 599 4025 633
rect 4059 599 4117 633
rect 4151 599 4209 633
rect 4243 599 4301 633
rect 4335 599 4393 633
rect 4427 599 4485 633
rect 4519 599 4577 633
rect 4611 599 4640 633
rect 86 568 4640 599
rect -10 562 86 568
rect -72 406 514 466
rect 574 406 580 466
rect 614 463 672 469
rect 614 429 626 463
rect 660 460 672 463
rect 1034 463 1092 469
rect 1034 460 1046 463
rect 660 432 1046 460
rect 660 429 672 432
rect 614 423 672 429
rect 1034 429 1046 432
rect 1080 460 1092 463
rect 1348 463 1406 469
rect 1348 460 1360 463
rect 1080 432 1360 460
rect 1080 429 1092 432
rect 1034 423 1092 429
rect 1348 429 1360 432
rect 1394 429 1406 463
rect 1348 423 1406 429
rect 2362 463 2420 469
rect 2362 429 2374 463
rect 2408 460 2420 463
rect 2782 463 2840 469
rect 2782 460 2794 463
rect 2408 432 2794 460
rect 2408 429 2420 432
rect 2362 423 2420 429
rect 2782 429 2794 432
rect 2828 460 2840 463
rect 3096 463 3154 469
rect 3096 460 3108 463
rect 2828 432 3108 460
rect 2828 429 2840 432
rect 2782 423 2840 429
rect 3096 429 3108 432
rect 3142 429 3154 463
rect 3096 423 3154 429
rect 4092 460 4394 466
rect 4092 412 4104 460
rect 4152 412 4394 460
rect 4092 406 4394 412
rect 514 376 574 406
rect -72 336 348 342
rect -72 288 288 336
rect 336 288 348 336
rect 514 328 520 376
rect 568 328 574 376
rect 693 395 751 401
rect 693 361 705 395
rect 739 392 751 395
rect 931 395 989 401
rect 931 392 943 395
rect 739 364 943 392
rect 739 361 751 364
rect 693 355 751 361
rect 931 361 943 364
rect 977 392 989 395
rect 1435 395 1493 401
rect 1435 392 1447 395
rect 977 364 1447 392
rect 977 361 989 364
rect 931 355 989 361
rect 1435 361 1447 364
rect 1481 361 1493 395
rect 2268 390 2328 396
rect 2441 395 2499 401
rect 1435 355 1493 361
rect 2262 330 2268 390
rect 2328 330 2334 390
rect 2441 361 2453 395
rect 2487 392 2499 395
rect 2679 395 2737 401
rect 2679 392 2691 395
rect 2487 364 2691 392
rect 2487 361 2499 364
rect 2441 355 2499 361
rect 2679 361 2691 364
rect 2725 392 2737 395
rect 3183 395 3241 401
rect 3183 392 3195 395
rect 2725 364 3195 392
rect 2725 361 2737 364
rect 2679 355 2737 361
rect 3183 361 3195 364
rect 3229 361 3241 395
rect 3183 355 3241 361
rect 4192 338 4252 344
rect 3934 332 4086 338
rect 514 316 574 328
rect 2268 324 2328 330
rect -72 282 348 288
rect 774 292 834 304
rect 774 248 780 292
rect 372 244 780 248
rect 828 244 834 292
rect 372 242 834 244
rect 372 194 384 242
rect 432 194 834 242
rect 2520 280 2580 292
rect 2520 236 2526 280
rect 372 188 834 194
rect 1874 232 2526 236
rect 2574 232 2580 280
rect 3934 284 4026 332
rect 4074 284 4086 332
rect 3934 278 4086 284
rect 4186 278 4192 338
rect 4252 278 4258 338
rect 4334 336 4394 406
rect 4334 288 4340 336
rect 4388 288 4394 336
rect 3624 236 3684 242
rect 3934 236 3994 278
rect 4192 272 4252 278
rect 4334 276 4394 288
rect 4430 332 4688 338
rect 4430 284 4442 332
rect 4490 284 4688 332
rect 4430 278 4688 284
rect 1874 230 2580 232
rect 1874 182 1886 230
rect 1934 182 2580 230
rect 1874 176 2580 182
rect 3622 176 3624 236
rect 3684 176 3994 236
rect 3624 170 3684 176
rect -10 89 4640 120
rect -10 55 161 89
rect 195 55 253 89
rect 287 55 345 89
rect 379 55 437 89
rect 471 55 529 89
rect 563 55 621 89
rect 655 55 713 89
rect 747 55 805 89
rect 839 55 897 89
rect 931 55 989 89
rect 1023 55 1081 89
rect 1115 55 1173 89
rect 1207 55 1265 89
rect 1299 55 1357 89
rect 1391 55 1449 89
rect 1483 55 1541 89
rect 1575 55 1633 89
rect 1667 55 1725 89
rect 1759 55 1817 89
rect 1851 55 1909 89
rect 1943 55 2001 89
rect 2035 55 2093 89
rect 2127 55 2185 89
rect 2219 55 2277 89
rect 2311 55 2369 89
rect 2403 55 2461 89
rect 2495 55 2553 89
rect 2587 55 2645 89
rect 2679 55 2737 89
rect 2771 55 2829 89
rect 2863 55 2921 89
rect 2955 55 3013 89
rect 3047 55 3105 89
rect 3139 55 3197 89
rect 3231 55 3289 89
rect 3323 55 3381 89
rect 3415 55 3473 89
rect 3507 55 3565 89
rect 3599 55 3657 89
rect 3691 55 3749 89
rect 3783 55 3841 89
rect 3875 55 3933 89
rect 3967 55 4025 89
rect 4059 55 4117 89
rect 4151 55 4209 89
rect 4243 55 4301 89
rect 4335 55 4393 89
rect 4427 55 4485 89
rect 4519 55 4577 89
rect 4611 55 4640 89
rect -10 24 4640 55
rect 2174 -30 2580 -24
rect 3934 -28 3994 -22
rect 774 -72 834 -66
rect 514 -132 574 -126
rect 768 -132 774 -72
rect 834 -132 840 -72
rect 2174 -78 2186 -30
rect 2234 -78 2580 -30
rect 2174 -84 2580 -78
rect 508 -192 514 -132
rect 574 -192 580 -132
rect 774 -138 834 -132
rect 2274 -136 2334 -130
rect 2520 -132 2526 -84
rect 2574 -132 2580 -84
rect 3624 -34 3934 -28
rect 3624 -82 3636 -34
rect 3684 -82 3934 -34
rect 3624 -88 3934 -82
rect 3934 -94 3994 -88
rect 514 -198 574 -192
rect 2268 -196 2274 -136
rect 2334 -196 2340 -136
rect 2520 -144 2580 -132
rect 2274 -202 2334 -196
rect 693 -217 751 -211
rect 693 -251 705 -217
rect 739 -220 751 -217
rect 931 -217 989 -211
rect 931 -220 943 -217
rect 739 -248 943 -220
rect 739 -251 751 -248
rect 693 -257 751 -251
rect 931 -251 943 -248
rect 977 -220 989 -217
rect 1435 -217 1493 -211
rect 1435 -220 1447 -217
rect 977 -248 1447 -220
rect 977 -251 989 -248
rect 931 -257 989 -251
rect 1435 -251 1447 -248
rect 1481 -251 1493 -217
rect 1435 -257 1493 -251
rect 2441 -217 2499 -211
rect 2441 -251 2453 -217
rect 2487 -220 2499 -217
rect 2679 -217 2737 -211
rect 2679 -220 2691 -217
rect 2487 -248 2691 -220
rect 2487 -251 2499 -248
rect 2441 -257 2499 -251
rect 2679 -251 2691 -248
rect 2725 -220 2737 -217
rect 3183 -217 3241 -211
rect 3183 -220 3195 -217
rect 2725 -248 3195 -220
rect 2725 -251 2737 -248
rect 2679 -257 2737 -251
rect 3183 -251 3195 -248
rect 3229 -251 3241 -217
rect 3183 -257 3241 -251
rect 614 -285 672 -279
rect 614 -319 626 -285
rect 660 -288 672 -285
rect 1034 -285 1092 -279
rect 1034 -288 1046 -285
rect 660 -316 1046 -288
rect 660 -319 672 -316
rect 614 -325 672 -319
rect 1034 -319 1046 -316
rect 1080 -288 1092 -285
rect 1348 -285 1406 -279
rect 1348 -288 1360 -285
rect 1080 -316 1360 -288
rect 1080 -319 1092 -316
rect 1034 -325 1092 -319
rect 1348 -319 1360 -316
rect 1394 -319 1406 -285
rect 1348 -325 1406 -319
rect 2362 -285 2420 -279
rect 2362 -319 2374 -285
rect 2408 -288 2420 -285
rect 2782 -285 2840 -279
rect 2782 -288 2794 -285
rect 2408 -316 2794 -288
rect 2408 -319 2420 -316
rect 2362 -325 2420 -319
rect 2782 -319 2794 -316
rect 2828 -288 2840 -285
rect 3096 -285 3154 -279
rect 3096 -288 3108 -285
rect 2828 -316 3108 -288
rect 2828 -319 2840 -316
rect 2782 -325 2840 -319
rect 3096 -319 3108 -316
rect 3142 -319 3154 -285
rect 3096 -325 3154 -319
rect -10 -424 86 -418
rect 86 -455 4088 -424
rect 86 -489 437 -455
rect 471 -489 529 -455
rect 563 -489 621 -455
rect 655 -489 713 -455
rect 747 -489 805 -455
rect 839 -489 897 -455
rect 931 -489 989 -455
rect 1023 -489 1081 -455
rect 1115 -489 1173 -455
rect 1207 -489 1265 -455
rect 1299 -489 1357 -455
rect 1391 -489 1449 -455
rect 1483 -489 1541 -455
rect 1575 -489 1633 -455
rect 1667 -489 1725 -455
rect 1759 -489 1817 -455
rect 1851 -489 1909 -455
rect 1943 -489 2001 -455
rect 2035 -489 2093 -455
rect 2127 -489 2185 -455
rect 2219 -489 2277 -455
rect 2311 -489 2369 -455
rect 2403 -489 2461 -455
rect 2495 -489 2553 -455
rect 2587 -489 2645 -455
rect 2679 -489 2737 -455
rect 2771 -489 2829 -455
rect 2863 -489 2921 -455
rect 2955 -489 3013 -455
rect 3047 -489 3105 -455
rect 3139 -489 3197 -455
rect 3231 -489 3289 -455
rect 3323 -489 3381 -455
rect 3415 -489 3473 -455
rect 3507 -489 3565 -455
rect 3599 -489 3657 -455
rect 3691 -489 3749 -455
rect 3783 -489 3841 -455
rect 3875 -489 3933 -455
rect 3967 -489 4025 -455
rect 4059 -489 4088 -455
rect 86 -520 4088 -489
rect -10 -526 86 -520
<< via1 >>
rect -10 568 86 664
rect 514 406 574 466
rect 2268 384 2328 390
rect 2268 336 2274 384
rect 2274 336 2322 384
rect 2322 336 2328 384
rect 2268 330 2328 336
rect 4192 332 4252 338
rect 4192 284 4198 332
rect 4198 284 4246 332
rect 4246 284 4252 332
rect 4192 278 4252 284
rect 3624 230 3684 236
rect 3624 182 3634 230
rect 3634 182 3682 230
rect 3682 182 3684 230
rect 3624 176 3684 182
rect 774 -78 834 -72
rect 774 -126 780 -78
rect 780 -126 828 -78
rect 828 -126 834 -78
rect 774 -132 834 -126
rect 514 -138 574 -132
rect 514 -186 520 -138
rect 520 -186 568 -138
rect 568 -186 574 -138
rect 514 -192 574 -186
rect 3934 -88 3994 -28
rect 2274 -142 2334 -136
rect 2274 -190 2280 -142
rect 2280 -190 2328 -142
rect 2328 -190 2334 -142
rect 2274 -196 2334 -190
rect -10 -520 86 -424
<< metal2 >>
rect -16 568 -10 664
rect 86 568 92 664
rect -10 -424 86 568
rect 514 466 574 472
rect 510 406 514 466
rect 574 406 2332 466
rect 514 -132 574 406
rect 2268 390 2328 406
rect 2268 324 2328 330
rect 3934 278 4192 338
rect 4252 278 4258 338
rect 3618 176 3624 236
rect 3684 176 3690 236
rect 3624 102 3684 176
rect 774 42 3684 102
rect 774 -72 834 42
rect 3934 -28 3994 278
rect 3928 -88 3934 -28
rect 3994 -88 4000 -28
rect 774 -138 834 -132
rect 2274 -136 2334 -130
rect 514 -214 574 -192
rect 2274 -214 2334 -196
rect 514 -274 2334 -214
rect -16 -520 -10 -424
rect 86 -520 92 -424
<< labels >>
flabel metal2 20 502 26 506 1 FreeSans 480 0 0 0 VDD
port 2 n power bidirectional
flabel metal1 94 100 96 104 1 FreeSans 480 0 0 0 VSS
port 3 n ground bidirectional
flabel metal1 -52 310 -44 318 1 FreeSans 480 0 0 0 trigb
port 1 n
flabel metal1 -52 434 -42 442 1 FreeSans 480 0 0 0 clk
port 4 n
flabel metal1 4644 304 4650 308 1 FreeSans 480 0 0 0 pulse
port 5 n
flabel metal1 4570 596 4623 625 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_3/VPWR
flabel metal1 4569 54 4620 92 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_3/VGND
rlabel comment 4548 72 4548 72 4 sky130_fd_sc_hd__tapvpwrvgnd_1_3/tapvpwrvgnd_1
flabel metal1 4018 -481 4071 -452 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VPWR
flabel metal1 4017 52 4068 90 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VGND
rlabel comment 3996 72 3996 72 2 sky130_fd_sc_hd__tapvpwrvgnd_1_0/tapvpwrvgnd_1
flabel locali 4118 157 4152 191 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/Y
flabel locali 4118 225 4152 259 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/Y
flabel locali 4118 293 4152 327 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/Y
flabel locali 4210 293 4244 327 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/B
flabel locali 4026 293 4060 327 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/A
flabel nwell 4210 599 4244 633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VPB
flabel pwell 4210 55 4244 89 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VNB
flabel metal1 4210 55 4244 89 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VGND
flabel metal1 4210 599 4244 633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VPWR
rlabel comment 4272 72 4272 72 6 sky130_fd_sc_hd__nand2_1_0/nand2_1
flabel locali 4436 361 4470 395 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/Y
flabel locali 4436 293 4470 327 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/Y
flabel locali 4344 293 4378 327 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/A
flabel nwell 4301 599 4335 633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VPB
flabel pwell 4301 55 4335 89 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VNB
flabel metal1 4301 55 4335 89 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VGND
flabel metal1 4301 599 4335 633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VPWR
rlabel comment 4272 72 4272 72 4 sky130_fd_sc_hd__inv_1_1/inv_1
flabel metal1 2277 55 2311 89 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/VGND
flabel metal1 2277 -489 2311 -455 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/VPWR
flabel locali 3933 -266 3967 -232 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/Q_N
flabel locali 2537 -183 2571 -149 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/D
flabel locali 2277 -183 2311 -149 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/CLK
flabel locali 3638 -47 3672 -13 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/Q
flabel pwell 2277 55 2311 89 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/VNB
flabel pwell 2294 72 2294 72 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/VNB
flabel nwell 2277 -489 2311 -455 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/VPB
flabel nwell 2294 -472 2294 -472 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/VPB
rlabel comment 2248 72 2248 72 2 sky130_fd_sc_hd__dfxbp_1_3/dfxbp_1
flabel metal1 2277 55 2311 89 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VGND
flabel metal1 2277 599 2311 633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VPWR
flabel locali 3933 376 3967 410 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/Q_N
flabel locali 2537 293 2571 327 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/D
flabel locali 2277 293 2311 327 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/CLK
flabel locali 3638 157 3672 191 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/Q
flabel pwell 2277 55 2311 89 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VNB
flabel pwell 2294 72 2294 72 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VNB
flabel nwell 2277 599 2311 633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VPB
flabel nwell 2294 616 2294 616 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VPB
rlabel comment 2248 72 2248 72 4 sky130_fd_sc_hd__dfxbp_1_1/dfxbp_1
flabel metal1 154 596 207 625 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_2/VPWR
flabel metal1 153 54 204 92 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_2/VGND
rlabel comment 132 72 132 72 4 sky130_fd_sc_hd__tapvpwrvgnd_1_2/tapvpwrvgnd_1
flabel metal1 430 -481 483 -452 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VPWR
flabel metal1 429 52 480 90 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VGND
rlabel comment 408 72 408 72 2 sky130_fd_sc_hd__tapvpwrvgnd_1_1/tapvpwrvgnd_1
flabel metal1 529 55 563 89 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/VGND
flabel metal1 529 -489 563 -455 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/VPWR
flabel locali 2185 -266 2219 -232 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/Q_N
flabel locali 789 -183 823 -149 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/D
flabel locali 529 -183 563 -149 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/CLK
flabel locali 1890 -47 1924 -13 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/Q
flabel pwell 529 55 563 89 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/VNB
flabel pwell 546 72 546 72 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/VNB
flabel nwell 529 -489 563 -455 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/VPB
flabel nwell 546 -472 546 -472 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/VPB
rlabel comment 500 72 500 72 2 sky130_fd_sc_hd__dfxbp_1_2/dfxbp_1
flabel metal1 529 55 563 89 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VGND
flabel metal1 529 599 563 633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VPWR
flabel locali 2185 376 2219 410 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/Q_N
flabel locali 789 293 823 327 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/D
flabel locali 529 293 563 327 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/CLK
flabel locali 1890 157 1924 191 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/Q
flabel pwell 529 55 563 89 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VNB
flabel pwell 546 72 546 72 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VNB
flabel nwell 529 599 563 633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VPB
flabel nwell 546 616 546 616 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VPB
rlabel comment 500 72 500 72 4 sky130_fd_sc_hd__dfxbp_1_0/dfxbp_1
flabel locali 388 361 422 395 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 388 293 422 327 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 296 293 330 327 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/A
flabel nwell 253 599 287 633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 253 55 287 89 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 253 55 287 89 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 253 599 287 633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 224 72 224 72 4 sky130_fd_sc_hd__inv_1_0/inv_1
<< end >>
