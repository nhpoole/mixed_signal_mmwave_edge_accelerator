magic
tech sky130A
magscale 1 2
timestamp 1622435379
<< nwell >>
rect -358 582 11058 2438
<< pwell >>
rect -358 -3058 11058 418
<< nmos >>
rect 782 -578 982 -178
rect 1040 -578 1240 -178
rect 1298 -578 1498 -178
rect 1556 -578 1756 -178
rect 1814 -578 2014 -178
rect 2072 -578 2272 -178
rect 2330 -578 2530 -178
rect 2588 -578 2788 -178
rect 2846 -578 3046 -178
rect 3104 -578 3304 -178
rect 7374 -578 7574 -178
rect 7632 -578 7832 -178
rect 7890 -578 8090 -178
rect 8148 -578 8348 -178
rect 8406 -578 8606 -178
rect 8664 -578 8864 -178
rect 8922 -578 9122 -178
rect 9180 -578 9380 -178
rect 9438 -578 9638 -178
rect 9696 -578 9896 -178
rect 234 -1486 1034 -1286
rect 1092 -1486 1892 -1286
rect 1950 -1486 2750 -1286
rect 2808 -1486 3608 -1286
rect 3666 -1486 4466 -1286
rect 4524 -1486 5324 -1286
rect 5382 -1486 6182 -1286
rect 6240 -1486 7040 -1286
rect 7098 -1486 7898 -1286
rect 7956 -1486 8756 -1286
rect 8814 -1486 9614 -1286
rect 9672 -1486 10472 -1286
rect 234 -2026 1034 -1826
rect 1092 -2026 1892 -1826
rect 1950 -2026 2750 -1826
rect 2808 -2026 3608 -1826
rect 3666 -2026 4466 -1826
rect 4524 -2026 5324 -1826
rect 5382 -2026 6182 -1826
rect 6240 -2026 7040 -1826
rect 7098 -2026 7898 -1826
rect 7956 -2026 8756 -1826
rect 8814 -2026 9614 -1826
rect 9672 -2026 10472 -1826
<< pmos >>
rect 3566 1090 3766 1290
rect 3824 1090 4024 1290
rect 4082 1090 4282 1290
rect 4340 1090 4540 1290
rect 4598 1090 4798 1290
rect 4856 1090 5056 1290
rect 5114 1090 5314 1290
rect 5372 1090 5572 1290
rect 5630 1090 5830 1290
rect 5888 1090 6088 1290
rect 6146 1090 6346 1290
rect 6404 1090 6604 1290
rect 6662 1090 6862 1290
rect 6920 1090 7120 1290
<< nmoslvt >>
rect 4078 -578 4278 -178
rect 4336 -578 4536 -178
rect 4594 -578 4794 -178
rect 4852 -578 5052 -178
rect 5110 -578 5310 -178
rect 5368 -578 5568 -178
rect 5626 -578 5826 -178
rect 5884 -578 6084 -178
rect 6142 -578 6342 -178
rect 6400 -578 6600 -178
<< ndiff >>
rect 724 -190 782 -178
rect 724 -566 736 -190
rect 770 -566 782 -190
rect 724 -578 782 -566
rect 982 -190 1040 -178
rect 982 -566 994 -190
rect 1028 -566 1040 -190
rect 982 -578 1040 -566
rect 1240 -190 1298 -178
rect 1240 -566 1252 -190
rect 1286 -566 1298 -190
rect 1240 -578 1298 -566
rect 1498 -190 1556 -178
rect 1498 -566 1510 -190
rect 1544 -566 1556 -190
rect 1498 -578 1556 -566
rect 1756 -190 1814 -178
rect 1756 -566 1768 -190
rect 1802 -566 1814 -190
rect 1756 -578 1814 -566
rect 2014 -190 2072 -178
rect 2014 -566 2026 -190
rect 2060 -566 2072 -190
rect 2014 -578 2072 -566
rect 2272 -190 2330 -178
rect 2272 -566 2284 -190
rect 2318 -566 2330 -190
rect 2272 -578 2330 -566
rect 2530 -190 2588 -178
rect 2530 -566 2542 -190
rect 2576 -566 2588 -190
rect 2530 -578 2588 -566
rect 2788 -190 2846 -178
rect 2788 -566 2800 -190
rect 2834 -566 2846 -190
rect 2788 -578 2846 -566
rect 3046 -190 3104 -178
rect 3046 -566 3058 -190
rect 3092 -566 3104 -190
rect 3046 -578 3104 -566
rect 3304 -190 3362 -178
rect 3304 -566 3316 -190
rect 3350 -566 3362 -190
rect 3304 -578 3362 -566
rect 4020 -190 4078 -178
rect 4020 -566 4032 -190
rect 4066 -566 4078 -190
rect 4020 -578 4078 -566
rect 4278 -190 4336 -178
rect 4278 -566 4290 -190
rect 4324 -566 4336 -190
rect 4278 -578 4336 -566
rect 4536 -190 4594 -178
rect 4536 -566 4548 -190
rect 4582 -566 4594 -190
rect 4536 -578 4594 -566
rect 4794 -190 4852 -178
rect 4794 -566 4806 -190
rect 4840 -566 4852 -190
rect 4794 -578 4852 -566
rect 5052 -190 5110 -178
rect 5052 -566 5064 -190
rect 5098 -566 5110 -190
rect 5052 -578 5110 -566
rect 5310 -190 5368 -178
rect 5310 -566 5322 -190
rect 5356 -566 5368 -190
rect 5310 -578 5368 -566
rect 5568 -190 5626 -178
rect 5568 -566 5580 -190
rect 5614 -566 5626 -190
rect 5568 -578 5626 -566
rect 5826 -190 5884 -178
rect 5826 -566 5838 -190
rect 5872 -566 5884 -190
rect 5826 -578 5884 -566
rect 6084 -190 6142 -178
rect 6084 -566 6096 -190
rect 6130 -566 6142 -190
rect 6084 -578 6142 -566
rect 6342 -190 6400 -178
rect 6342 -566 6354 -190
rect 6388 -566 6400 -190
rect 6342 -578 6400 -566
rect 6600 -190 6658 -178
rect 6600 -566 6612 -190
rect 6646 -566 6658 -190
rect 6600 -578 6658 -566
rect 7316 -190 7374 -178
rect 7316 -566 7328 -190
rect 7362 -566 7374 -190
rect 7316 -578 7374 -566
rect 7574 -190 7632 -178
rect 7574 -566 7586 -190
rect 7620 -566 7632 -190
rect 7574 -578 7632 -566
rect 7832 -190 7890 -178
rect 7832 -566 7844 -190
rect 7878 -566 7890 -190
rect 7832 -578 7890 -566
rect 8090 -190 8148 -178
rect 8090 -566 8102 -190
rect 8136 -566 8148 -190
rect 8090 -578 8148 -566
rect 8348 -190 8406 -178
rect 8348 -566 8360 -190
rect 8394 -566 8406 -190
rect 8348 -578 8406 -566
rect 8606 -190 8664 -178
rect 8606 -566 8618 -190
rect 8652 -566 8664 -190
rect 8606 -578 8664 -566
rect 8864 -190 8922 -178
rect 8864 -566 8876 -190
rect 8910 -566 8922 -190
rect 8864 -578 8922 -566
rect 9122 -190 9180 -178
rect 9122 -566 9134 -190
rect 9168 -566 9180 -190
rect 9122 -578 9180 -566
rect 9380 -190 9438 -178
rect 9380 -566 9392 -190
rect 9426 -566 9438 -190
rect 9380 -578 9438 -566
rect 9638 -190 9696 -178
rect 9638 -566 9650 -190
rect 9684 -566 9696 -190
rect 9638 -578 9696 -566
rect 9896 -190 9954 -178
rect 9896 -566 9908 -190
rect 9942 -566 9954 -190
rect 9896 -578 9954 -566
rect 176 -1298 234 -1286
rect 176 -1474 188 -1298
rect 222 -1474 234 -1298
rect 176 -1486 234 -1474
rect 1034 -1298 1092 -1286
rect 1034 -1474 1046 -1298
rect 1080 -1474 1092 -1298
rect 1034 -1486 1092 -1474
rect 1892 -1298 1950 -1286
rect 1892 -1474 1904 -1298
rect 1938 -1474 1950 -1298
rect 1892 -1486 1950 -1474
rect 2750 -1298 2808 -1286
rect 2750 -1474 2762 -1298
rect 2796 -1474 2808 -1298
rect 2750 -1486 2808 -1474
rect 3608 -1298 3666 -1286
rect 3608 -1474 3620 -1298
rect 3654 -1474 3666 -1298
rect 3608 -1486 3666 -1474
rect 4466 -1298 4524 -1286
rect 4466 -1474 4478 -1298
rect 4512 -1474 4524 -1298
rect 4466 -1486 4524 -1474
rect 5324 -1298 5382 -1286
rect 5324 -1474 5336 -1298
rect 5370 -1474 5382 -1298
rect 5324 -1486 5382 -1474
rect 6182 -1298 6240 -1286
rect 6182 -1474 6194 -1298
rect 6228 -1474 6240 -1298
rect 6182 -1486 6240 -1474
rect 7040 -1298 7098 -1286
rect 7040 -1474 7052 -1298
rect 7086 -1474 7098 -1298
rect 7040 -1486 7098 -1474
rect 7898 -1298 7956 -1286
rect 7898 -1474 7910 -1298
rect 7944 -1474 7956 -1298
rect 7898 -1486 7956 -1474
rect 8756 -1298 8814 -1286
rect 8756 -1474 8768 -1298
rect 8802 -1474 8814 -1298
rect 8756 -1486 8814 -1474
rect 9614 -1298 9672 -1286
rect 9614 -1474 9626 -1298
rect 9660 -1474 9672 -1298
rect 9614 -1486 9672 -1474
rect 10472 -1298 10530 -1286
rect 10472 -1474 10484 -1298
rect 10518 -1474 10530 -1298
rect 10472 -1486 10530 -1474
rect 176 -1838 234 -1826
rect 176 -2014 188 -1838
rect 222 -2014 234 -1838
rect 176 -2026 234 -2014
rect 1034 -1838 1092 -1826
rect 1034 -2014 1046 -1838
rect 1080 -2014 1092 -1838
rect 1034 -2026 1092 -2014
rect 1892 -1838 1950 -1826
rect 1892 -2014 1904 -1838
rect 1938 -2014 1950 -1838
rect 1892 -2026 1950 -2014
rect 2750 -1838 2808 -1826
rect 2750 -2014 2762 -1838
rect 2796 -2014 2808 -1838
rect 2750 -2026 2808 -2014
rect 3608 -1838 3666 -1826
rect 3608 -2014 3620 -1838
rect 3654 -2014 3666 -1838
rect 3608 -2026 3666 -2014
rect 4466 -1838 4524 -1826
rect 4466 -2014 4478 -1838
rect 4512 -2014 4524 -1838
rect 4466 -2026 4524 -2014
rect 5324 -1838 5382 -1826
rect 5324 -2014 5336 -1838
rect 5370 -2014 5382 -1838
rect 5324 -2026 5382 -2014
rect 6182 -1838 6240 -1826
rect 6182 -2014 6194 -1838
rect 6228 -2014 6240 -1838
rect 6182 -2026 6240 -2014
rect 7040 -1838 7098 -1826
rect 7040 -2014 7052 -1838
rect 7086 -2014 7098 -1838
rect 7040 -2026 7098 -2014
rect 7898 -1838 7956 -1826
rect 7898 -2014 7910 -1838
rect 7944 -2014 7956 -1838
rect 7898 -2026 7956 -2014
rect 8756 -1838 8814 -1826
rect 8756 -2014 8768 -1838
rect 8802 -2014 8814 -1838
rect 8756 -2026 8814 -2014
rect 9614 -1838 9672 -1826
rect 9614 -2014 9626 -1838
rect 9660 -2014 9672 -1838
rect 9614 -2026 9672 -2014
rect 10472 -1838 10530 -1826
rect 10472 -2014 10484 -1838
rect 10518 -2014 10530 -1838
rect 10472 -2026 10530 -2014
<< pdiff >>
rect 3508 1278 3566 1290
rect 3508 1102 3520 1278
rect 3554 1102 3566 1278
rect 3508 1090 3566 1102
rect 3766 1278 3824 1290
rect 3766 1102 3778 1278
rect 3812 1102 3824 1278
rect 3766 1090 3824 1102
rect 4024 1278 4082 1290
rect 4024 1102 4036 1278
rect 4070 1102 4082 1278
rect 4024 1090 4082 1102
rect 4282 1278 4340 1290
rect 4282 1102 4294 1278
rect 4328 1102 4340 1278
rect 4282 1090 4340 1102
rect 4540 1278 4598 1290
rect 4540 1102 4552 1278
rect 4586 1102 4598 1278
rect 4540 1090 4598 1102
rect 4798 1278 4856 1290
rect 4798 1102 4810 1278
rect 4844 1102 4856 1278
rect 4798 1090 4856 1102
rect 5056 1278 5114 1290
rect 5056 1102 5068 1278
rect 5102 1102 5114 1278
rect 5056 1090 5114 1102
rect 5314 1278 5372 1290
rect 5314 1102 5326 1278
rect 5360 1102 5372 1278
rect 5314 1090 5372 1102
rect 5572 1278 5630 1290
rect 5572 1102 5584 1278
rect 5618 1102 5630 1278
rect 5572 1090 5630 1102
rect 5830 1278 5888 1290
rect 5830 1102 5842 1278
rect 5876 1102 5888 1278
rect 5830 1090 5888 1102
rect 6088 1278 6146 1290
rect 6088 1102 6100 1278
rect 6134 1102 6146 1278
rect 6088 1090 6146 1102
rect 6346 1278 6404 1290
rect 6346 1102 6358 1278
rect 6392 1102 6404 1278
rect 6346 1090 6404 1102
rect 6604 1278 6662 1290
rect 6604 1102 6616 1278
rect 6650 1102 6662 1278
rect 6604 1090 6662 1102
rect 6862 1278 6920 1290
rect 6862 1102 6874 1278
rect 6908 1102 6920 1278
rect 6862 1090 6920 1102
rect 7120 1278 7178 1290
rect 7120 1102 7132 1278
rect 7166 1102 7178 1278
rect 7120 1090 7178 1102
<< ndiffc >>
rect 736 -566 770 -190
rect 994 -566 1028 -190
rect 1252 -566 1286 -190
rect 1510 -566 1544 -190
rect 1768 -566 1802 -190
rect 2026 -566 2060 -190
rect 2284 -566 2318 -190
rect 2542 -566 2576 -190
rect 2800 -566 2834 -190
rect 3058 -566 3092 -190
rect 3316 -566 3350 -190
rect 4032 -566 4066 -190
rect 4290 -566 4324 -190
rect 4548 -566 4582 -190
rect 4806 -566 4840 -190
rect 5064 -566 5098 -190
rect 5322 -566 5356 -190
rect 5580 -566 5614 -190
rect 5838 -566 5872 -190
rect 6096 -566 6130 -190
rect 6354 -566 6388 -190
rect 6612 -566 6646 -190
rect 7328 -566 7362 -190
rect 7586 -566 7620 -190
rect 7844 -566 7878 -190
rect 8102 -566 8136 -190
rect 8360 -566 8394 -190
rect 8618 -566 8652 -190
rect 8876 -566 8910 -190
rect 9134 -566 9168 -190
rect 9392 -566 9426 -190
rect 9650 -566 9684 -190
rect 9908 -566 9942 -190
rect 188 -1474 222 -1298
rect 1046 -1474 1080 -1298
rect 1904 -1474 1938 -1298
rect 2762 -1474 2796 -1298
rect 3620 -1474 3654 -1298
rect 4478 -1474 4512 -1298
rect 5336 -1474 5370 -1298
rect 6194 -1474 6228 -1298
rect 7052 -1474 7086 -1298
rect 7910 -1474 7944 -1298
rect 8768 -1474 8802 -1298
rect 9626 -1474 9660 -1298
rect 10484 -1474 10518 -1298
rect 188 -2014 222 -1838
rect 1046 -2014 1080 -1838
rect 1904 -2014 1938 -1838
rect 2762 -2014 2796 -1838
rect 3620 -2014 3654 -1838
rect 4478 -2014 4512 -1838
rect 5336 -2014 5370 -1838
rect 6194 -2014 6228 -1838
rect 7052 -2014 7086 -1838
rect 7910 -2014 7944 -1838
rect 8768 -2014 8802 -1838
rect 9626 -2014 9660 -1838
rect 10484 -2014 10518 -1838
<< pdiffc >>
rect 3520 1102 3554 1278
rect 3778 1102 3812 1278
rect 4036 1102 4070 1278
rect 4294 1102 4328 1278
rect 4552 1102 4586 1278
rect 4810 1102 4844 1278
rect 5068 1102 5102 1278
rect 5326 1102 5360 1278
rect 5584 1102 5618 1278
rect 5842 1102 5876 1278
rect 6100 1102 6134 1278
rect 6358 1102 6392 1278
rect 6616 1102 6650 1278
rect 6874 1102 6908 1278
rect 7132 1102 7166 1278
<< psubdiff >>
rect -322 282 -160 382
rect 10860 282 11022 382
rect -322 220 -222 282
rect 10922 220 11022 282
rect -322 -2922 -222 -2860
rect 10922 -2922 11022 -2860
rect -322 -3022 -160 -2922
rect 10860 -3022 11022 -2922
<< nsubdiff >>
rect -322 2302 -160 2402
rect 10860 2302 11022 2402
rect -322 2240 -222 2302
rect 10922 2240 11022 2302
rect -322 718 -222 780
rect 10922 718 11022 780
rect -322 618 -160 718
rect 10860 618 11022 718
<< psubdiffcont >>
rect -160 282 10860 382
rect -322 -2860 -222 220
rect 10922 -2860 11022 220
rect -160 -3022 10860 -2922
<< nsubdiffcont >>
rect -160 2302 10860 2402
rect -322 780 -222 2240
rect 10922 780 11022 2240
rect -160 618 10860 718
<< poly >>
rect 3600 1371 3732 1387
rect 3600 1354 3616 1371
rect 3566 1337 3616 1354
rect 3716 1354 3732 1371
rect 3858 1371 3990 1387
rect 3858 1354 3874 1371
rect 3716 1337 3766 1354
rect 3566 1290 3766 1337
rect 3824 1337 3874 1354
rect 3974 1354 3990 1371
rect 4116 1371 4248 1387
rect 4116 1354 4132 1371
rect 3974 1337 4024 1354
rect 3824 1290 4024 1337
rect 4082 1337 4132 1354
rect 4232 1354 4248 1371
rect 4374 1371 4506 1387
rect 4374 1354 4390 1371
rect 4232 1337 4282 1354
rect 4082 1290 4282 1337
rect 4340 1337 4390 1354
rect 4490 1354 4506 1371
rect 4632 1371 4764 1387
rect 4632 1354 4648 1371
rect 4490 1337 4540 1354
rect 4340 1290 4540 1337
rect 4598 1337 4648 1354
rect 4748 1354 4764 1371
rect 4890 1371 5022 1387
rect 4890 1354 4906 1371
rect 4748 1337 4798 1354
rect 4598 1290 4798 1337
rect 4856 1337 4906 1354
rect 5006 1354 5022 1371
rect 5148 1371 5280 1387
rect 5148 1354 5164 1371
rect 5006 1337 5056 1354
rect 4856 1290 5056 1337
rect 5114 1337 5164 1354
rect 5264 1354 5280 1371
rect 5406 1371 5538 1387
rect 5406 1354 5422 1371
rect 5264 1337 5314 1354
rect 5114 1290 5314 1337
rect 5372 1337 5422 1354
rect 5522 1354 5538 1371
rect 5664 1371 5796 1387
rect 5664 1354 5680 1371
rect 5522 1337 5572 1354
rect 5372 1290 5572 1337
rect 5630 1337 5680 1354
rect 5780 1354 5796 1371
rect 5922 1371 6054 1387
rect 5922 1354 5938 1371
rect 5780 1337 5830 1354
rect 5630 1290 5830 1337
rect 5888 1337 5938 1354
rect 6038 1354 6054 1371
rect 6180 1371 6312 1387
rect 6180 1354 6196 1371
rect 6038 1337 6088 1354
rect 5888 1290 6088 1337
rect 6146 1337 6196 1354
rect 6296 1354 6312 1371
rect 6438 1371 6570 1387
rect 6438 1354 6454 1371
rect 6296 1337 6346 1354
rect 6146 1290 6346 1337
rect 6404 1337 6454 1354
rect 6554 1354 6570 1371
rect 6696 1371 6828 1387
rect 6696 1354 6712 1371
rect 6554 1337 6604 1354
rect 6404 1290 6604 1337
rect 6662 1337 6712 1354
rect 6812 1354 6828 1371
rect 6954 1371 7086 1387
rect 6954 1354 6970 1371
rect 6812 1337 6862 1354
rect 6662 1290 6862 1337
rect 6920 1337 6970 1354
rect 7070 1354 7086 1371
rect 7070 1337 7120 1354
rect 6920 1290 7120 1337
rect 3566 1043 3766 1090
rect 3566 1026 3616 1043
rect 3600 1009 3616 1026
rect 3716 1026 3766 1043
rect 3824 1043 4024 1090
rect 3824 1026 3874 1043
rect 3716 1009 3732 1026
rect 3600 993 3732 1009
rect 3858 1009 3874 1026
rect 3974 1026 4024 1043
rect 4082 1043 4282 1090
rect 4082 1026 4132 1043
rect 3974 1009 3990 1026
rect 3858 993 3990 1009
rect 4116 1009 4132 1026
rect 4232 1026 4282 1043
rect 4340 1043 4540 1090
rect 4340 1026 4390 1043
rect 4232 1009 4248 1026
rect 4116 993 4248 1009
rect 4374 1009 4390 1026
rect 4490 1026 4540 1043
rect 4598 1043 4798 1090
rect 4598 1026 4648 1043
rect 4490 1009 4506 1026
rect 4374 993 4506 1009
rect 4632 1009 4648 1026
rect 4748 1026 4798 1043
rect 4856 1043 5056 1090
rect 4856 1026 4906 1043
rect 4748 1009 4764 1026
rect 4632 993 4764 1009
rect 4890 1009 4906 1026
rect 5006 1026 5056 1043
rect 5114 1043 5314 1090
rect 5114 1026 5164 1043
rect 5006 1009 5022 1026
rect 4890 993 5022 1009
rect 5148 1009 5164 1026
rect 5264 1026 5314 1043
rect 5372 1043 5572 1090
rect 5372 1026 5422 1043
rect 5264 1009 5280 1026
rect 5148 993 5280 1009
rect 5406 1009 5422 1026
rect 5522 1026 5572 1043
rect 5630 1043 5830 1090
rect 5630 1026 5680 1043
rect 5522 1009 5538 1026
rect 5406 993 5538 1009
rect 5664 1009 5680 1026
rect 5780 1026 5830 1043
rect 5888 1043 6088 1090
rect 5888 1026 5938 1043
rect 5780 1009 5796 1026
rect 5664 993 5796 1009
rect 5922 1009 5938 1026
rect 6038 1026 6088 1043
rect 6146 1043 6346 1090
rect 6146 1026 6196 1043
rect 6038 1009 6054 1026
rect 5922 993 6054 1009
rect 6180 1009 6196 1026
rect 6296 1026 6346 1043
rect 6404 1043 6604 1090
rect 6404 1026 6454 1043
rect 6296 1009 6312 1026
rect 6180 993 6312 1009
rect 6438 1009 6454 1026
rect 6554 1026 6604 1043
rect 6662 1043 6862 1090
rect 6662 1026 6712 1043
rect 6554 1009 6570 1026
rect 6438 993 6570 1009
rect 6696 1009 6712 1026
rect 6812 1026 6862 1043
rect 6920 1043 7120 1090
rect 6920 1026 6970 1043
rect 6812 1009 6828 1026
rect 6696 993 6828 1009
rect 6954 1009 6970 1026
rect 7070 1026 7120 1043
rect 7070 1009 7086 1026
rect 6954 993 7086 1009
rect 816 -106 948 -90
rect 816 -123 832 -106
rect 782 -140 832 -123
rect 932 -123 948 -106
rect 1074 -106 1206 -90
rect 1074 -123 1090 -106
rect 932 -140 982 -123
rect 782 -178 982 -140
rect 1040 -140 1090 -123
rect 1190 -123 1206 -106
rect 1332 -106 1464 -90
rect 1332 -123 1348 -106
rect 1190 -140 1240 -123
rect 1040 -178 1240 -140
rect 1298 -140 1348 -123
rect 1448 -123 1464 -106
rect 1590 -106 1722 -90
rect 1590 -123 1606 -106
rect 1448 -140 1498 -123
rect 1298 -178 1498 -140
rect 1556 -140 1606 -123
rect 1706 -123 1722 -106
rect 1848 -106 1980 -90
rect 1848 -123 1864 -106
rect 1706 -140 1756 -123
rect 1556 -178 1756 -140
rect 1814 -140 1864 -123
rect 1964 -123 1980 -106
rect 2106 -106 2238 -90
rect 2106 -123 2122 -106
rect 1964 -140 2014 -123
rect 1814 -178 2014 -140
rect 2072 -140 2122 -123
rect 2222 -123 2238 -106
rect 2364 -106 2496 -90
rect 2364 -123 2380 -106
rect 2222 -140 2272 -123
rect 2072 -178 2272 -140
rect 2330 -140 2380 -123
rect 2480 -123 2496 -106
rect 2622 -106 2754 -90
rect 2622 -123 2638 -106
rect 2480 -140 2530 -123
rect 2330 -178 2530 -140
rect 2588 -140 2638 -123
rect 2738 -123 2754 -106
rect 2880 -106 3012 -90
rect 2880 -123 2896 -106
rect 2738 -140 2788 -123
rect 2588 -178 2788 -140
rect 2846 -140 2896 -123
rect 2996 -123 3012 -106
rect 3138 -106 3270 -90
rect 3138 -123 3154 -106
rect 2996 -140 3046 -123
rect 2846 -178 3046 -140
rect 3104 -140 3154 -123
rect 3254 -123 3270 -106
rect 4112 -106 4244 -90
rect 4112 -123 4128 -106
rect 3254 -140 3304 -123
rect 3104 -178 3304 -140
rect 4078 -140 4128 -123
rect 4228 -123 4244 -106
rect 4370 -106 4502 -90
rect 4370 -123 4386 -106
rect 4228 -140 4278 -123
rect 4078 -178 4278 -140
rect 4336 -140 4386 -123
rect 4486 -123 4502 -106
rect 4628 -106 4760 -90
rect 4628 -123 4644 -106
rect 4486 -140 4536 -123
rect 4336 -178 4536 -140
rect 4594 -140 4644 -123
rect 4744 -123 4760 -106
rect 4886 -106 5018 -90
rect 4886 -123 4902 -106
rect 4744 -140 4794 -123
rect 4594 -178 4794 -140
rect 4852 -140 4902 -123
rect 5002 -123 5018 -106
rect 5144 -106 5276 -90
rect 5144 -123 5160 -106
rect 5002 -140 5052 -123
rect 4852 -178 5052 -140
rect 5110 -140 5160 -123
rect 5260 -123 5276 -106
rect 5402 -106 5534 -90
rect 5402 -123 5418 -106
rect 5260 -140 5310 -123
rect 5110 -178 5310 -140
rect 5368 -140 5418 -123
rect 5518 -123 5534 -106
rect 5660 -106 5792 -90
rect 5660 -123 5676 -106
rect 5518 -140 5568 -123
rect 5368 -178 5568 -140
rect 5626 -140 5676 -123
rect 5776 -123 5792 -106
rect 5918 -106 6050 -90
rect 5918 -123 5934 -106
rect 5776 -140 5826 -123
rect 5626 -178 5826 -140
rect 5884 -140 5934 -123
rect 6034 -123 6050 -106
rect 6176 -106 6308 -90
rect 6176 -123 6192 -106
rect 6034 -140 6084 -123
rect 5884 -178 6084 -140
rect 6142 -140 6192 -123
rect 6292 -123 6308 -106
rect 6434 -106 6566 -90
rect 6434 -123 6450 -106
rect 6292 -140 6342 -123
rect 6142 -178 6342 -140
rect 6400 -140 6450 -123
rect 6550 -123 6566 -106
rect 7408 -106 7540 -90
rect 7408 -123 7424 -106
rect 6550 -140 6600 -123
rect 6400 -178 6600 -140
rect 7374 -140 7424 -123
rect 7524 -123 7540 -106
rect 7666 -106 7798 -90
rect 7666 -123 7682 -106
rect 7524 -140 7574 -123
rect 7374 -178 7574 -140
rect 7632 -140 7682 -123
rect 7782 -123 7798 -106
rect 7924 -106 8056 -90
rect 7924 -123 7940 -106
rect 7782 -140 7832 -123
rect 7632 -178 7832 -140
rect 7890 -140 7940 -123
rect 8040 -123 8056 -106
rect 8182 -106 8314 -90
rect 8182 -123 8198 -106
rect 8040 -140 8090 -123
rect 7890 -178 8090 -140
rect 8148 -140 8198 -123
rect 8298 -123 8314 -106
rect 8440 -106 8572 -90
rect 8440 -123 8456 -106
rect 8298 -140 8348 -123
rect 8148 -178 8348 -140
rect 8406 -140 8456 -123
rect 8556 -123 8572 -106
rect 8698 -106 8830 -90
rect 8698 -123 8714 -106
rect 8556 -140 8606 -123
rect 8406 -178 8606 -140
rect 8664 -140 8714 -123
rect 8814 -123 8830 -106
rect 8956 -106 9088 -90
rect 8956 -123 8972 -106
rect 8814 -140 8864 -123
rect 8664 -178 8864 -140
rect 8922 -140 8972 -123
rect 9072 -123 9088 -106
rect 9214 -106 9346 -90
rect 9214 -123 9230 -106
rect 9072 -140 9122 -123
rect 8922 -178 9122 -140
rect 9180 -140 9230 -123
rect 9330 -123 9346 -106
rect 9472 -106 9604 -90
rect 9472 -123 9488 -106
rect 9330 -140 9380 -123
rect 9180 -178 9380 -140
rect 9438 -140 9488 -123
rect 9588 -123 9604 -106
rect 9730 -106 9862 -90
rect 9730 -123 9746 -106
rect 9588 -140 9638 -123
rect 9438 -178 9638 -140
rect 9696 -140 9746 -123
rect 9846 -123 9862 -106
rect 9846 -140 9896 -123
rect 9696 -178 9896 -140
rect 782 -616 982 -578
rect 782 -633 832 -616
rect 816 -650 832 -633
rect 932 -633 982 -616
rect 1040 -616 1240 -578
rect 1040 -633 1090 -616
rect 932 -650 948 -633
rect 816 -666 948 -650
rect 1074 -650 1090 -633
rect 1190 -633 1240 -616
rect 1298 -616 1498 -578
rect 1298 -633 1348 -616
rect 1190 -650 1206 -633
rect 1074 -666 1206 -650
rect 1332 -650 1348 -633
rect 1448 -633 1498 -616
rect 1556 -616 1756 -578
rect 1556 -633 1606 -616
rect 1448 -650 1464 -633
rect 1332 -666 1464 -650
rect 1590 -650 1606 -633
rect 1706 -633 1756 -616
rect 1814 -616 2014 -578
rect 1814 -633 1864 -616
rect 1706 -650 1722 -633
rect 1590 -666 1722 -650
rect 1848 -650 1864 -633
rect 1964 -633 2014 -616
rect 2072 -616 2272 -578
rect 2072 -633 2122 -616
rect 1964 -650 1980 -633
rect 1848 -666 1980 -650
rect 2106 -650 2122 -633
rect 2222 -633 2272 -616
rect 2330 -616 2530 -578
rect 2330 -633 2380 -616
rect 2222 -650 2238 -633
rect 2106 -666 2238 -650
rect 2364 -650 2380 -633
rect 2480 -633 2530 -616
rect 2588 -616 2788 -578
rect 2588 -633 2638 -616
rect 2480 -650 2496 -633
rect 2364 -666 2496 -650
rect 2622 -650 2638 -633
rect 2738 -633 2788 -616
rect 2846 -616 3046 -578
rect 2846 -633 2896 -616
rect 2738 -650 2754 -633
rect 2622 -666 2754 -650
rect 2880 -650 2896 -633
rect 2996 -633 3046 -616
rect 3104 -616 3304 -578
rect 3104 -633 3154 -616
rect 2996 -650 3012 -633
rect 2880 -666 3012 -650
rect 3138 -650 3154 -633
rect 3254 -633 3304 -616
rect 4078 -616 4278 -578
rect 4078 -633 4128 -616
rect 3254 -650 3270 -633
rect 3138 -666 3270 -650
rect 4112 -650 4128 -633
rect 4228 -633 4278 -616
rect 4336 -616 4536 -578
rect 4336 -633 4386 -616
rect 4228 -650 4244 -633
rect 4112 -666 4244 -650
rect 4370 -650 4386 -633
rect 4486 -633 4536 -616
rect 4594 -616 4794 -578
rect 4594 -633 4644 -616
rect 4486 -650 4502 -633
rect 4370 -666 4502 -650
rect 4628 -650 4644 -633
rect 4744 -633 4794 -616
rect 4852 -616 5052 -578
rect 4852 -633 4902 -616
rect 4744 -650 4760 -633
rect 4628 -666 4760 -650
rect 4886 -650 4902 -633
rect 5002 -633 5052 -616
rect 5110 -616 5310 -578
rect 5110 -633 5160 -616
rect 5002 -650 5018 -633
rect 4886 -666 5018 -650
rect 5144 -650 5160 -633
rect 5260 -633 5310 -616
rect 5368 -616 5568 -578
rect 5368 -633 5418 -616
rect 5260 -650 5276 -633
rect 5144 -666 5276 -650
rect 5402 -650 5418 -633
rect 5518 -633 5568 -616
rect 5626 -616 5826 -578
rect 5626 -633 5676 -616
rect 5518 -650 5534 -633
rect 5402 -666 5534 -650
rect 5660 -650 5676 -633
rect 5776 -633 5826 -616
rect 5884 -616 6084 -578
rect 5884 -633 5934 -616
rect 5776 -650 5792 -633
rect 5660 -666 5792 -650
rect 5918 -650 5934 -633
rect 6034 -633 6084 -616
rect 6142 -616 6342 -578
rect 6142 -633 6192 -616
rect 6034 -650 6050 -633
rect 5918 -666 6050 -650
rect 6176 -650 6192 -633
rect 6292 -633 6342 -616
rect 6400 -616 6600 -578
rect 6400 -633 6450 -616
rect 6292 -650 6308 -633
rect 6176 -666 6308 -650
rect 6434 -650 6450 -633
rect 6550 -633 6600 -616
rect 7374 -616 7574 -578
rect 7374 -633 7424 -616
rect 6550 -650 6566 -633
rect 6434 -666 6566 -650
rect 7408 -650 7424 -633
rect 7524 -633 7574 -616
rect 7632 -616 7832 -578
rect 7632 -633 7682 -616
rect 7524 -650 7540 -633
rect 7408 -666 7540 -650
rect 7666 -650 7682 -633
rect 7782 -633 7832 -616
rect 7890 -616 8090 -578
rect 7890 -633 7940 -616
rect 7782 -650 7798 -633
rect 7666 -666 7798 -650
rect 7924 -650 7940 -633
rect 8040 -633 8090 -616
rect 8148 -616 8348 -578
rect 8148 -633 8198 -616
rect 8040 -650 8056 -633
rect 7924 -666 8056 -650
rect 8182 -650 8198 -633
rect 8298 -633 8348 -616
rect 8406 -616 8606 -578
rect 8406 -633 8456 -616
rect 8298 -650 8314 -633
rect 8182 -666 8314 -650
rect 8440 -650 8456 -633
rect 8556 -633 8606 -616
rect 8664 -616 8864 -578
rect 8664 -633 8714 -616
rect 8556 -650 8572 -633
rect 8440 -666 8572 -650
rect 8698 -650 8714 -633
rect 8814 -633 8864 -616
rect 8922 -616 9122 -578
rect 8922 -633 8972 -616
rect 8814 -650 8830 -633
rect 8698 -666 8830 -650
rect 8956 -650 8972 -633
rect 9072 -633 9122 -616
rect 9180 -616 9380 -578
rect 9180 -633 9230 -616
rect 9072 -650 9088 -633
rect 8956 -666 9088 -650
rect 9214 -650 9230 -633
rect 9330 -633 9380 -616
rect 9438 -616 9638 -578
rect 9438 -633 9488 -616
rect 9330 -650 9346 -633
rect 9214 -666 9346 -650
rect 9472 -650 9488 -633
rect 9588 -633 9638 -616
rect 9696 -616 9896 -578
rect 9696 -633 9746 -616
rect 9588 -650 9604 -633
rect 9472 -666 9604 -650
rect 9730 -650 9746 -633
rect 9846 -633 9896 -616
rect 9846 -650 9862 -633
rect 9730 -666 9862 -650
rect 388 -1214 880 -1198
rect 388 -1231 404 -1214
rect 234 -1248 404 -1231
rect 864 -1231 880 -1214
rect 1246 -1214 1738 -1198
rect 1246 -1231 1262 -1214
rect 864 -1248 1034 -1231
rect 234 -1286 1034 -1248
rect 1092 -1248 1262 -1231
rect 1722 -1231 1738 -1214
rect 2104 -1214 2596 -1198
rect 2104 -1231 2120 -1214
rect 1722 -1248 1892 -1231
rect 1092 -1286 1892 -1248
rect 1950 -1248 2120 -1231
rect 2580 -1231 2596 -1214
rect 2962 -1214 3454 -1198
rect 2962 -1231 2978 -1214
rect 2580 -1248 2750 -1231
rect 1950 -1286 2750 -1248
rect 2808 -1248 2978 -1231
rect 3438 -1231 3454 -1214
rect 3820 -1214 4312 -1198
rect 3820 -1231 3836 -1214
rect 3438 -1248 3608 -1231
rect 2808 -1286 3608 -1248
rect 3666 -1248 3836 -1231
rect 4296 -1231 4312 -1214
rect 4678 -1214 5170 -1198
rect 4678 -1231 4694 -1214
rect 4296 -1248 4466 -1231
rect 3666 -1286 4466 -1248
rect 4524 -1248 4694 -1231
rect 5154 -1231 5170 -1214
rect 5536 -1214 6028 -1198
rect 5536 -1231 5552 -1214
rect 5154 -1248 5324 -1231
rect 4524 -1286 5324 -1248
rect 5382 -1248 5552 -1231
rect 6012 -1231 6028 -1214
rect 6394 -1214 6886 -1198
rect 6394 -1231 6410 -1214
rect 6012 -1248 6182 -1231
rect 5382 -1286 6182 -1248
rect 6240 -1248 6410 -1231
rect 6870 -1231 6886 -1214
rect 7252 -1214 7744 -1198
rect 7252 -1231 7268 -1214
rect 6870 -1248 7040 -1231
rect 6240 -1286 7040 -1248
rect 7098 -1248 7268 -1231
rect 7728 -1231 7744 -1214
rect 8110 -1214 8602 -1198
rect 8110 -1231 8126 -1214
rect 7728 -1248 7898 -1231
rect 7098 -1286 7898 -1248
rect 7956 -1248 8126 -1231
rect 8586 -1231 8602 -1214
rect 8968 -1214 9460 -1198
rect 8968 -1231 8984 -1214
rect 8586 -1248 8756 -1231
rect 7956 -1286 8756 -1248
rect 8814 -1248 8984 -1231
rect 9444 -1231 9460 -1214
rect 9826 -1214 10318 -1198
rect 9826 -1231 9842 -1214
rect 9444 -1248 9614 -1231
rect 8814 -1286 9614 -1248
rect 9672 -1248 9842 -1231
rect 10302 -1231 10318 -1214
rect 10302 -1248 10472 -1231
rect 9672 -1286 10472 -1248
rect 234 -1524 1034 -1486
rect 234 -1541 404 -1524
rect 388 -1558 404 -1541
rect 864 -1541 1034 -1524
rect 1092 -1524 1892 -1486
rect 1092 -1541 1262 -1524
rect 864 -1558 880 -1541
rect 388 -1574 880 -1558
rect 1246 -1558 1262 -1541
rect 1722 -1541 1892 -1524
rect 1950 -1524 2750 -1486
rect 1950 -1541 2120 -1524
rect 1722 -1558 1738 -1541
rect 1246 -1574 1738 -1558
rect 2104 -1558 2120 -1541
rect 2580 -1541 2750 -1524
rect 2808 -1524 3608 -1486
rect 2808 -1541 2978 -1524
rect 2580 -1558 2596 -1541
rect 2104 -1574 2596 -1558
rect 2962 -1558 2978 -1541
rect 3438 -1541 3608 -1524
rect 3666 -1524 4466 -1486
rect 3666 -1541 3836 -1524
rect 3438 -1558 3454 -1541
rect 2962 -1574 3454 -1558
rect 3820 -1558 3836 -1541
rect 4296 -1541 4466 -1524
rect 4524 -1524 5324 -1486
rect 4524 -1541 4694 -1524
rect 4296 -1558 4312 -1541
rect 3820 -1574 4312 -1558
rect 4678 -1558 4694 -1541
rect 5154 -1541 5324 -1524
rect 5382 -1524 6182 -1486
rect 5382 -1541 5552 -1524
rect 5154 -1558 5170 -1541
rect 4678 -1574 5170 -1558
rect 5536 -1558 5552 -1541
rect 6012 -1541 6182 -1524
rect 6240 -1524 7040 -1486
rect 6240 -1541 6410 -1524
rect 6012 -1558 6028 -1541
rect 5536 -1574 6028 -1558
rect 6394 -1558 6410 -1541
rect 6870 -1541 7040 -1524
rect 7098 -1524 7898 -1486
rect 7098 -1541 7268 -1524
rect 6870 -1558 6886 -1541
rect 6394 -1574 6886 -1558
rect 7252 -1558 7268 -1541
rect 7728 -1541 7898 -1524
rect 7956 -1524 8756 -1486
rect 7956 -1541 8126 -1524
rect 7728 -1558 7744 -1541
rect 7252 -1574 7744 -1558
rect 8110 -1558 8126 -1541
rect 8586 -1541 8756 -1524
rect 8814 -1524 9614 -1486
rect 8814 -1541 8984 -1524
rect 8586 -1558 8602 -1541
rect 8110 -1574 8602 -1558
rect 8968 -1558 8984 -1541
rect 9444 -1541 9614 -1524
rect 9672 -1524 10472 -1486
rect 9672 -1541 9842 -1524
rect 9444 -1558 9460 -1541
rect 8968 -1574 9460 -1558
rect 9826 -1558 9842 -1541
rect 10302 -1541 10472 -1524
rect 10302 -1558 10318 -1541
rect 9826 -1574 10318 -1558
rect 388 -1754 880 -1738
rect 388 -1771 404 -1754
rect 234 -1788 404 -1771
rect 864 -1771 880 -1754
rect 1246 -1754 1738 -1738
rect 1246 -1771 1262 -1754
rect 864 -1788 1034 -1771
rect 234 -1826 1034 -1788
rect 1092 -1788 1262 -1771
rect 1722 -1771 1738 -1754
rect 2104 -1754 2596 -1738
rect 2104 -1771 2120 -1754
rect 1722 -1788 1892 -1771
rect 1092 -1826 1892 -1788
rect 1950 -1788 2120 -1771
rect 2580 -1771 2596 -1754
rect 2962 -1754 3454 -1738
rect 2962 -1771 2978 -1754
rect 2580 -1788 2750 -1771
rect 1950 -1826 2750 -1788
rect 2808 -1788 2978 -1771
rect 3438 -1771 3454 -1754
rect 3820 -1754 4312 -1738
rect 3820 -1771 3836 -1754
rect 3438 -1788 3608 -1771
rect 2808 -1826 3608 -1788
rect 3666 -1788 3836 -1771
rect 4296 -1771 4312 -1754
rect 4678 -1754 5170 -1738
rect 4678 -1771 4694 -1754
rect 4296 -1788 4466 -1771
rect 3666 -1826 4466 -1788
rect 4524 -1788 4694 -1771
rect 5154 -1771 5170 -1754
rect 5536 -1754 6028 -1738
rect 5536 -1771 5552 -1754
rect 5154 -1788 5324 -1771
rect 4524 -1826 5324 -1788
rect 5382 -1788 5552 -1771
rect 6012 -1771 6028 -1754
rect 6394 -1754 6886 -1738
rect 6394 -1771 6410 -1754
rect 6012 -1788 6182 -1771
rect 5382 -1826 6182 -1788
rect 6240 -1788 6410 -1771
rect 6870 -1771 6886 -1754
rect 7252 -1754 7744 -1738
rect 7252 -1771 7268 -1754
rect 6870 -1788 7040 -1771
rect 6240 -1826 7040 -1788
rect 7098 -1788 7268 -1771
rect 7728 -1771 7744 -1754
rect 8110 -1754 8602 -1738
rect 8110 -1771 8126 -1754
rect 7728 -1788 7898 -1771
rect 7098 -1826 7898 -1788
rect 7956 -1788 8126 -1771
rect 8586 -1771 8602 -1754
rect 8968 -1754 9460 -1738
rect 8968 -1771 8984 -1754
rect 8586 -1788 8756 -1771
rect 7956 -1826 8756 -1788
rect 8814 -1788 8984 -1771
rect 9444 -1771 9460 -1754
rect 9826 -1754 10318 -1738
rect 9826 -1771 9842 -1754
rect 9444 -1788 9614 -1771
rect 8814 -1826 9614 -1788
rect 9672 -1788 9842 -1771
rect 10302 -1771 10318 -1754
rect 10302 -1788 10472 -1771
rect 9672 -1826 10472 -1788
rect 234 -2064 1034 -2026
rect 234 -2081 404 -2064
rect 388 -2098 404 -2081
rect 864 -2081 1034 -2064
rect 1092 -2064 1892 -2026
rect 1092 -2081 1262 -2064
rect 864 -2098 880 -2081
rect 388 -2114 880 -2098
rect 1246 -2098 1262 -2081
rect 1722 -2081 1892 -2064
rect 1950 -2064 2750 -2026
rect 1950 -2081 2120 -2064
rect 1722 -2098 1738 -2081
rect 1246 -2114 1738 -2098
rect 2104 -2098 2120 -2081
rect 2580 -2081 2750 -2064
rect 2808 -2064 3608 -2026
rect 2808 -2081 2978 -2064
rect 2580 -2098 2596 -2081
rect 2104 -2114 2596 -2098
rect 2962 -2098 2978 -2081
rect 3438 -2081 3608 -2064
rect 3666 -2064 4466 -2026
rect 3666 -2081 3836 -2064
rect 3438 -2098 3454 -2081
rect 2962 -2114 3454 -2098
rect 3820 -2098 3836 -2081
rect 4296 -2081 4466 -2064
rect 4524 -2064 5324 -2026
rect 4524 -2081 4694 -2064
rect 4296 -2098 4312 -2081
rect 3820 -2114 4312 -2098
rect 4678 -2098 4694 -2081
rect 5154 -2081 5324 -2064
rect 5382 -2064 6182 -2026
rect 5382 -2081 5552 -2064
rect 5154 -2098 5170 -2081
rect 4678 -2114 5170 -2098
rect 5536 -2098 5552 -2081
rect 6012 -2081 6182 -2064
rect 6240 -2064 7040 -2026
rect 6240 -2081 6410 -2064
rect 6012 -2098 6028 -2081
rect 5536 -2114 6028 -2098
rect 6394 -2098 6410 -2081
rect 6870 -2081 7040 -2064
rect 7098 -2064 7898 -2026
rect 7098 -2081 7268 -2064
rect 6870 -2098 6886 -2081
rect 6394 -2114 6886 -2098
rect 7252 -2098 7268 -2081
rect 7728 -2081 7898 -2064
rect 7956 -2064 8756 -2026
rect 7956 -2081 8126 -2064
rect 7728 -2098 7744 -2081
rect 7252 -2114 7744 -2098
rect 8110 -2098 8126 -2081
rect 8586 -2081 8756 -2064
rect 8814 -2064 9614 -2026
rect 8814 -2081 8984 -2064
rect 8586 -2098 8602 -2081
rect 8110 -2114 8602 -2098
rect 8968 -2098 8984 -2081
rect 9444 -2081 9614 -2064
rect 9672 -2064 10472 -2026
rect 9672 -2081 9842 -2064
rect 9444 -2098 9460 -2081
rect 8968 -2114 9460 -2098
rect 9826 -2098 9842 -2081
rect 10302 -2081 10472 -2064
rect 10302 -2098 10318 -2081
rect 9826 -2114 10318 -2098
<< polycont >>
rect 3616 1337 3716 1371
rect 3874 1337 3974 1371
rect 4132 1337 4232 1371
rect 4390 1337 4490 1371
rect 4648 1337 4748 1371
rect 4906 1337 5006 1371
rect 5164 1337 5264 1371
rect 5422 1337 5522 1371
rect 5680 1337 5780 1371
rect 5938 1337 6038 1371
rect 6196 1337 6296 1371
rect 6454 1337 6554 1371
rect 6712 1337 6812 1371
rect 6970 1337 7070 1371
rect 3616 1009 3716 1043
rect 3874 1009 3974 1043
rect 4132 1009 4232 1043
rect 4390 1009 4490 1043
rect 4648 1009 4748 1043
rect 4906 1009 5006 1043
rect 5164 1009 5264 1043
rect 5422 1009 5522 1043
rect 5680 1009 5780 1043
rect 5938 1009 6038 1043
rect 6196 1009 6296 1043
rect 6454 1009 6554 1043
rect 6712 1009 6812 1043
rect 6970 1009 7070 1043
rect 832 -140 932 -106
rect 1090 -140 1190 -106
rect 1348 -140 1448 -106
rect 1606 -140 1706 -106
rect 1864 -140 1964 -106
rect 2122 -140 2222 -106
rect 2380 -140 2480 -106
rect 2638 -140 2738 -106
rect 2896 -140 2996 -106
rect 3154 -140 3254 -106
rect 4128 -140 4228 -106
rect 4386 -140 4486 -106
rect 4644 -140 4744 -106
rect 4902 -140 5002 -106
rect 5160 -140 5260 -106
rect 5418 -140 5518 -106
rect 5676 -140 5776 -106
rect 5934 -140 6034 -106
rect 6192 -140 6292 -106
rect 6450 -140 6550 -106
rect 7424 -140 7524 -106
rect 7682 -140 7782 -106
rect 7940 -140 8040 -106
rect 8198 -140 8298 -106
rect 8456 -140 8556 -106
rect 8714 -140 8814 -106
rect 8972 -140 9072 -106
rect 9230 -140 9330 -106
rect 9488 -140 9588 -106
rect 9746 -140 9846 -106
rect 832 -650 932 -616
rect 1090 -650 1190 -616
rect 1348 -650 1448 -616
rect 1606 -650 1706 -616
rect 1864 -650 1964 -616
rect 2122 -650 2222 -616
rect 2380 -650 2480 -616
rect 2638 -650 2738 -616
rect 2896 -650 2996 -616
rect 3154 -650 3254 -616
rect 4128 -650 4228 -616
rect 4386 -650 4486 -616
rect 4644 -650 4744 -616
rect 4902 -650 5002 -616
rect 5160 -650 5260 -616
rect 5418 -650 5518 -616
rect 5676 -650 5776 -616
rect 5934 -650 6034 -616
rect 6192 -650 6292 -616
rect 6450 -650 6550 -616
rect 7424 -650 7524 -616
rect 7682 -650 7782 -616
rect 7940 -650 8040 -616
rect 8198 -650 8298 -616
rect 8456 -650 8556 -616
rect 8714 -650 8814 -616
rect 8972 -650 9072 -616
rect 9230 -650 9330 -616
rect 9488 -650 9588 -616
rect 9746 -650 9846 -616
rect 404 -1248 864 -1214
rect 1262 -1248 1722 -1214
rect 2120 -1248 2580 -1214
rect 2978 -1248 3438 -1214
rect 3836 -1248 4296 -1214
rect 4694 -1248 5154 -1214
rect 5552 -1248 6012 -1214
rect 6410 -1248 6870 -1214
rect 7268 -1248 7728 -1214
rect 8126 -1248 8586 -1214
rect 8984 -1248 9444 -1214
rect 9842 -1248 10302 -1214
rect 404 -1558 864 -1524
rect 1262 -1558 1722 -1524
rect 2120 -1558 2580 -1524
rect 2978 -1558 3438 -1524
rect 3836 -1558 4296 -1524
rect 4694 -1558 5154 -1524
rect 5552 -1558 6012 -1524
rect 6410 -1558 6870 -1524
rect 7268 -1558 7728 -1524
rect 8126 -1558 8586 -1524
rect 8984 -1558 9444 -1524
rect 9842 -1558 10302 -1524
rect 404 -1788 864 -1754
rect 1262 -1788 1722 -1754
rect 2120 -1788 2580 -1754
rect 2978 -1788 3438 -1754
rect 3836 -1788 4296 -1754
rect 4694 -1788 5154 -1754
rect 5552 -1788 6012 -1754
rect 6410 -1788 6870 -1754
rect 7268 -1788 7728 -1754
rect 8126 -1788 8586 -1754
rect 8984 -1788 9444 -1754
rect 9842 -1788 10302 -1754
rect 404 -2098 864 -2064
rect 1262 -2098 1722 -2064
rect 2120 -2098 2580 -2064
rect 2978 -2098 3438 -2064
rect 3836 -2098 4296 -2064
rect 4694 -2098 5154 -2064
rect 5552 -2098 6012 -2064
rect 6410 -2098 6870 -2064
rect 7268 -2098 7728 -2064
rect 8126 -2098 8586 -2064
rect 8984 -2098 9444 -2064
rect 9842 -2098 10302 -2064
<< locali >>
rect -322 2242 -222 2402
rect 10922 2242 11022 2402
rect 3600 1337 3616 1371
rect 3716 1337 3732 1371
rect 3858 1337 3874 1371
rect 3974 1337 3990 1371
rect 4116 1337 4132 1371
rect 4232 1337 4248 1371
rect 4374 1337 4390 1371
rect 4490 1337 4506 1371
rect 4632 1337 4648 1371
rect 4748 1337 4764 1371
rect 4890 1337 4906 1371
rect 5006 1337 5022 1371
rect 5148 1337 5164 1371
rect 5264 1337 5280 1371
rect 5406 1337 5422 1371
rect 5522 1337 5538 1371
rect 5664 1337 5680 1371
rect 5780 1337 5796 1371
rect 5922 1337 5938 1371
rect 6038 1337 6054 1371
rect 6180 1337 6196 1371
rect 6296 1337 6312 1371
rect 6438 1337 6454 1371
rect 6554 1337 6570 1371
rect 6696 1337 6712 1371
rect 6812 1337 6828 1371
rect 6954 1337 6970 1371
rect 7070 1337 7086 1371
rect 3520 1278 3554 1294
rect 3520 1086 3554 1102
rect 3778 1278 3812 1294
rect 3778 1086 3812 1102
rect 4036 1278 4070 1294
rect 4036 1086 4070 1102
rect 4294 1278 4328 1294
rect 4294 1086 4328 1102
rect 4552 1278 4586 1294
rect 4552 1086 4586 1102
rect 4810 1278 4844 1294
rect 4810 1086 4844 1102
rect 5068 1278 5102 1294
rect 5068 1086 5102 1102
rect 5326 1278 5360 1294
rect 5326 1086 5360 1102
rect 5584 1278 5618 1294
rect 5584 1086 5618 1102
rect 5842 1278 5876 1294
rect 5842 1086 5876 1102
rect 6100 1278 6134 1294
rect 6100 1086 6134 1102
rect 6358 1278 6392 1294
rect 6358 1086 6392 1102
rect 6616 1278 6650 1294
rect 6616 1086 6650 1102
rect 6874 1278 6908 1294
rect 6874 1086 6908 1102
rect 7132 1278 7166 1294
rect 7132 1086 7166 1102
rect 3600 1009 3616 1043
rect 3716 1009 3732 1043
rect 3858 1009 3874 1043
rect 3974 1009 3990 1043
rect 4116 1009 4132 1043
rect 4232 1009 4248 1043
rect 4374 1009 4390 1043
rect 4490 1009 4506 1043
rect 4632 1009 4648 1043
rect 4748 1009 4764 1043
rect 4890 1009 4906 1043
rect 5006 1009 5022 1043
rect 5148 1009 5164 1043
rect 5264 1009 5280 1043
rect 5406 1009 5422 1043
rect 5522 1009 5538 1043
rect 5664 1009 5680 1043
rect 5780 1009 5796 1043
rect 5922 1009 5938 1043
rect 6038 1009 6054 1043
rect 6180 1009 6196 1043
rect 6296 1009 6312 1043
rect 6438 1009 6454 1043
rect 6554 1009 6570 1043
rect 6696 1009 6712 1043
rect 6812 1009 6828 1043
rect 6954 1009 6970 1043
rect 7070 1009 7086 1043
rect -322 618 -222 778
rect 10922 618 11022 778
rect -322 220 -222 382
rect 10922 220 11022 382
rect 816 -140 832 -106
rect 932 -140 948 -106
rect 1074 -140 1090 -106
rect 1190 -140 1206 -106
rect 1332 -140 1348 -106
rect 1448 -140 1464 -106
rect 1590 -140 1606 -106
rect 1706 -140 1722 -106
rect 1848 -140 1864 -106
rect 1964 -140 1980 -106
rect 2106 -140 2122 -106
rect 2222 -140 2238 -106
rect 2364 -140 2380 -106
rect 2480 -140 2496 -106
rect 2622 -140 2638 -106
rect 2738 -140 2754 -106
rect 2880 -140 2896 -106
rect 2996 -140 3012 -106
rect 3138 -140 3154 -106
rect 3254 -140 3270 -106
rect 4112 -140 4128 -106
rect 4228 -140 4244 -106
rect 4370 -140 4386 -106
rect 4486 -140 4502 -106
rect 4628 -140 4644 -106
rect 4744 -140 4760 -106
rect 4886 -140 4902 -106
rect 5002 -140 5018 -106
rect 5144 -140 5160 -106
rect 5260 -140 5276 -106
rect 5402 -140 5418 -106
rect 5518 -140 5534 -106
rect 5660 -140 5676 -106
rect 5776 -140 5792 -106
rect 5918 -140 5934 -106
rect 6034 -140 6050 -106
rect 6176 -140 6192 -106
rect 6292 -140 6308 -106
rect 6434 -140 6450 -106
rect 6550 -140 6566 -106
rect 7408 -140 7424 -106
rect 7524 -140 7540 -106
rect 7666 -140 7682 -106
rect 7782 -140 7798 -106
rect 7924 -140 7940 -106
rect 8040 -140 8056 -106
rect 8182 -140 8198 -106
rect 8298 -140 8314 -106
rect 8440 -140 8456 -106
rect 8556 -140 8572 -106
rect 8698 -140 8714 -106
rect 8814 -140 8830 -106
rect 8956 -140 8972 -106
rect 9072 -140 9088 -106
rect 9214 -140 9230 -106
rect 9330 -140 9346 -106
rect 9472 -140 9488 -106
rect 9588 -140 9604 -106
rect 9730 -140 9746 -106
rect 9846 -140 9862 -106
rect 736 -190 770 -174
rect 736 -582 770 -566
rect 994 -190 1028 -174
rect 994 -582 1028 -566
rect 1252 -190 1286 -174
rect 1252 -582 1286 -566
rect 1510 -190 1544 -174
rect 1510 -582 1544 -566
rect 1768 -190 1802 -174
rect 1768 -582 1802 -566
rect 2026 -190 2060 -174
rect 2026 -582 2060 -566
rect 2284 -190 2318 -174
rect 2284 -582 2318 -566
rect 2542 -190 2576 -174
rect 2542 -582 2576 -566
rect 2800 -190 2834 -174
rect 2800 -582 2834 -566
rect 3058 -190 3092 -174
rect 3058 -582 3092 -566
rect 3316 -190 3350 -174
rect 3316 -582 3350 -566
rect 4032 -190 4066 -174
rect 4032 -582 4066 -566
rect 4290 -190 4324 -174
rect 4290 -582 4324 -566
rect 4548 -190 4582 -174
rect 4548 -582 4582 -566
rect 4806 -190 4840 -174
rect 4806 -582 4840 -566
rect 5064 -190 5098 -174
rect 5064 -582 5098 -566
rect 5322 -190 5356 -174
rect 5322 -582 5356 -566
rect 5580 -190 5614 -174
rect 5580 -582 5614 -566
rect 5838 -190 5872 -174
rect 5838 -582 5872 -566
rect 6096 -190 6130 -174
rect 6096 -582 6130 -566
rect 6354 -190 6388 -174
rect 6354 -582 6388 -566
rect 6612 -190 6646 -174
rect 6612 -582 6646 -566
rect 7328 -190 7362 -174
rect 7328 -582 7362 -566
rect 7586 -190 7620 -174
rect 7586 -582 7620 -566
rect 7844 -190 7878 -174
rect 7844 -582 7878 -566
rect 8102 -190 8136 -174
rect 8102 -582 8136 -566
rect 8360 -190 8394 -174
rect 8360 -582 8394 -566
rect 8618 -190 8652 -174
rect 8618 -582 8652 -566
rect 8876 -190 8910 -174
rect 8876 -582 8910 -566
rect 9134 -190 9168 -174
rect 9134 -582 9168 -566
rect 9392 -190 9426 -174
rect 9392 -582 9426 -566
rect 9650 -190 9684 -174
rect 9650 -582 9684 -566
rect 9908 -190 9942 -174
rect 9908 -582 9942 -566
rect 816 -650 832 -616
rect 932 -650 948 -616
rect 1074 -650 1090 -616
rect 1190 -650 1206 -616
rect 1332 -650 1348 -616
rect 1448 -650 1464 -616
rect 1590 -650 1606 -616
rect 1706 -650 1722 -616
rect 1848 -650 1864 -616
rect 1964 -650 1980 -616
rect 2106 -650 2122 -616
rect 2222 -650 2238 -616
rect 2364 -650 2380 -616
rect 2480 -650 2496 -616
rect 2622 -650 2638 -616
rect 2738 -650 2754 -616
rect 2880 -650 2896 -616
rect 2996 -650 3012 -616
rect 3138 -650 3154 -616
rect 3254 -650 3270 -616
rect 4112 -650 4128 -616
rect 4228 -650 4244 -616
rect 4370 -650 4386 -616
rect 4486 -650 4502 -616
rect 4628 -650 4644 -616
rect 4744 -650 4760 -616
rect 4886 -650 4902 -616
rect 5002 -650 5018 -616
rect 5144 -650 5160 -616
rect 5260 -650 5276 -616
rect 5402 -650 5418 -616
rect 5518 -650 5534 -616
rect 5660 -650 5676 -616
rect 5776 -650 5792 -616
rect 5918 -650 5934 -616
rect 6034 -650 6050 -616
rect 6176 -650 6192 -616
rect 6292 -650 6308 -616
rect 6434 -650 6450 -616
rect 6550 -650 6566 -616
rect 7408 -650 7424 -616
rect 7524 -650 7540 -616
rect 7666 -650 7682 -616
rect 7782 -650 7798 -616
rect 7924 -650 7940 -616
rect 8040 -650 8056 -616
rect 8182 -650 8198 -616
rect 8298 -650 8314 -616
rect 8440 -650 8456 -616
rect 8556 -650 8572 -616
rect 8698 -650 8714 -616
rect 8814 -650 8830 -616
rect 8956 -650 8972 -616
rect 9072 -650 9088 -616
rect 9214 -650 9230 -616
rect 9330 -650 9346 -616
rect 9472 -650 9488 -616
rect 9588 -650 9604 -616
rect 9730 -650 9746 -616
rect 9846 -650 9862 -616
rect 388 -1248 404 -1214
rect 864 -1248 880 -1214
rect 1246 -1248 1262 -1214
rect 1722 -1248 1738 -1214
rect 2104 -1248 2120 -1214
rect 2580 -1248 2596 -1214
rect 2962 -1248 2978 -1214
rect 3438 -1248 3454 -1214
rect 3820 -1248 3836 -1214
rect 4296 -1248 4312 -1214
rect 4678 -1248 4694 -1214
rect 5154 -1248 5170 -1214
rect 5536 -1248 5552 -1214
rect 6012 -1248 6028 -1214
rect 6394 -1248 6410 -1214
rect 6870 -1248 6886 -1214
rect 7252 -1248 7268 -1214
rect 7728 -1248 7744 -1214
rect 8110 -1248 8126 -1214
rect 8586 -1248 8602 -1214
rect 8968 -1248 8984 -1214
rect 9444 -1248 9460 -1214
rect 9826 -1248 9842 -1214
rect 10302 -1248 10318 -1214
rect 188 -1298 222 -1282
rect 188 -1490 222 -1474
rect 1046 -1298 1080 -1282
rect 1046 -1490 1080 -1474
rect 1904 -1298 1938 -1282
rect 1904 -1490 1938 -1474
rect 2762 -1298 2796 -1282
rect 2762 -1490 2796 -1474
rect 3620 -1298 3654 -1282
rect 3620 -1490 3654 -1474
rect 4478 -1298 4512 -1282
rect 4478 -1490 4512 -1474
rect 5336 -1298 5370 -1282
rect 5336 -1490 5370 -1474
rect 6194 -1298 6228 -1282
rect 6194 -1490 6228 -1474
rect 7052 -1298 7086 -1282
rect 7052 -1490 7086 -1474
rect 7910 -1298 7944 -1282
rect 7910 -1490 7944 -1474
rect 8768 -1298 8802 -1282
rect 8768 -1490 8802 -1474
rect 9626 -1298 9660 -1282
rect 9626 -1490 9660 -1474
rect 10484 -1298 10518 -1282
rect 10484 -1490 10518 -1474
rect 388 -1558 404 -1524
rect 864 -1558 880 -1524
rect 1246 -1558 1262 -1524
rect 1722 -1558 1738 -1524
rect 2104 -1558 2120 -1524
rect 2580 -1558 2596 -1524
rect 2962 -1558 2978 -1524
rect 3438 -1558 3454 -1524
rect 3820 -1558 3836 -1524
rect 4296 -1558 4312 -1524
rect 4678 -1558 4694 -1524
rect 5154 -1558 5170 -1524
rect 5536 -1558 5552 -1524
rect 6012 -1558 6028 -1524
rect 6394 -1558 6410 -1524
rect 6870 -1558 6886 -1524
rect 7252 -1558 7268 -1524
rect 7728 -1558 7744 -1524
rect 8110 -1558 8126 -1524
rect 8586 -1558 8602 -1524
rect 8968 -1558 8984 -1524
rect 9444 -1558 9460 -1524
rect 9826 -1558 9842 -1524
rect 10302 -1558 10318 -1524
rect 388 -1788 404 -1754
rect 864 -1788 880 -1754
rect 1246 -1788 1262 -1754
rect 1722 -1788 1738 -1754
rect 2104 -1788 2120 -1754
rect 2580 -1788 2596 -1754
rect 2962 -1788 2978 -1754
rect 3438 -1788 3454 -1754
rect 3820 -1788 3836 -1754
rect 4296 -1788 4312 -1754
rect 4678 -1788 4694 -1754
rect 5154 -1788 5170 -1754
rect 5536 -1788 5552 -1754
rect 6012 -1788 6028 -1754
rect 6394 -1788 6410 -1754
rect 6870 -1788 6886 -1754
rect 7252 -1788 7268 -1754
rect 7728 -1788 7744 -1754
rect 8110 -1788 8126 -1754
rect 8586 -1788 8602 -1754
rect 8968 -1788 8984 -1754
rect 9444 -1788 9460 -1754
rect 9826 -1788 9842 -1754
rect 10302 -1788 10318 -1754
rect 188 -1838 222 -1822
rect 188 -2030 222 -2014
rect 1046 -1838 1080 -1822
rect 1046 -2030 1080 -2014
rect 1904 -1838 1938 -1822
rect 1904 -2030 1938 -2014
rect 2762 -1838 2796 -1822
rect 2762 -2030 2796 -2014
rect 3620 -1838 3654 -1822
rect 3620 -2030 3654 -2014
rect 4478 -1838 4512 -1822
rect 4478 -2030 4512 -2014
rect 5336 -1838 5370 -1822
rect 5336 -2030 5370 -2014
rect 6194 -1838 6228 -1822
rect 6194 -2030 6228 -2014
rect 7052 -1838 7086 -1822
rect 7052 -2030 7086 -2014
rect 7910 -1838 7944 -1822
rect 7910 -2030 7944 -2014
rect 8768 -1838 8802 -1822
rect 8768 -2030 8802 -2014
rect 9626 -1838 9660 -1822
rect 9626 -2030 9660 -2014
rect 10484 -1838 10518 -1822
rect 10484 -2030 10518 -2014
rect 388 -2098 404 -2064
rect 864 -2098 880 -2064
rect 1246 -2098 1262 -2064
rect 1722 -2098 1738 -2064
rect 2104 -2098 2120 -2064
rect 2580 -2098 2596 -2064
rect 2962 -2098 2978 -2064
rect 3438 -2098 3454 -2064
rect 3820 -2098 3836 -2064
rect 4296 -2098 4312 -2064
rect 4678 -2098 4694 -2064
rect 5154 -2098 5170 -2064
rect 5536 -2098 5552 -2064
rect 6012 -2098 6028 -2064
rect 6394 -2098 6410 -2064
rect 6870 -2098 6886 -2064
rect 7252 -2098 7268 -2064
rect 7728 -2098 7744 -2064
rect 8110 -2098 8126 -2064
rect 8586 -2098 8602 -2064
rect 8968 -2098 8984 -2064
rect 9444 -2098 9460 -2064
rect 9826 -2098 9842 -2064
rect 10302 -2098 10318 -2064
rect -322 -3022 -222 -2860
rect 10922 -3022 11022 -2860
<< viali >>
rect -222 2302 -160 2402
rect -160 2302 10860 2402
rect 10860 2302 10922 2402
rect -322 2240 -222 2242
rect -322 780 -222 2240
rect 10922 2240 11022 2242
rect 3624 1337 3708 1371
rect 3882 1337 3966 1371
rect 4140 1337 4224 1371
rect 4398 1337 4482 1371
rect 4656 1337 4740 1371
rect 4914 1337 4998 1371
rect 5172 1337 5256 1371
rect 5430 1337 5514 1371
rect 5688 1337 5772 1371
rect 5946 1337 6030 1371
rect 6204 1337 6288 1371
rect 6462 1337 6546 1371
rect 6720 1337 6804 1371
rect 6978 1337 7062 1371
rect 3520 1102 3554 1278
rect 3778 1102 3812 1278
rect 4036 1102 4070 1278
rect 4294 1102 4328 1278
rect 4552 1102 4586 1278
rect 4810 1102 4844 1278
rect 5068 1102 5102 1278
rect 5326 1102 5360 1278
rect 5584 1102 5618 1278
rect 5842 1102 5876 1278
rect 6100 1102 6134 1278
rect 6358 1102 6392 1278
rect 6616 1102 6650 1278
rect 6874 1102 6908 1278
rect 7132 1102 7166 1278
rect 3624 1009 3708 1043
rect 3882 1009 3966 1043
rect 4140 1009 4224 1043
rect 4398 1009 4482 1043
rect 4656 1009 4740 1043
rect 4914 1009 4998 1043
rect 5172 1009 5256 1043
rect 5430 1009 5514 1043
rect 5688 1009 5772 1043
rect 5946 1009 6030 1043
rect 6204 1009 6288 1043
rect 6462 1009 6546 1043
rect 6720 1009 6804 1043
rect 6978 1009 7062 1043
rect -322 778 -222 780
rect 10922 780 11022 2240
rect 10922 778 11022 780
rect -222 618 -160 718
rect -160 618 10860 718
rect 10860 618 10922 718
rect -222 282 -160 382
rect -160 282 10860 382
rect 10860 282 10922 382
rect -322 -2762 -222 122
rect 840 -140 924 -106
rect 1098 -140 1182 -106
rect 1356 -140 1440 -106
rect 1614 -140 1698 -106
rect 1872 -140 1956 -106
rect 2130 -140 2214 -106
rect 2388 -140 2472 -106
rect 2646 -140 2730 -106
rect 2904 -140 2988 -106
rect 3162 -140 3246 -106
rect 4136 -140 4220 -106
rect 4394 -140 4478 -106
rect 4652 -140 4736 -106
rect 4910 -140 4994 -106
rect 5168 -140 5252 -106
rect 5426 -140 5510 -106
rect 5684 -140 5768 -106
rect 5942 -140 6026 -106
rect 6200 -140 6284 -106
rect 6458 -140 6542 -106
rect 7432 -140 7516 -106
rect 7690 -140 7774 -106
rect 7948 -140 8032 -106
rect 8206 -140 8290 -106
rect 8464 -140 8548 -106
rect 8722 -140 8806 -106
rect 8980 -140 9064 -106
rect 9238 -140 9322 -106
rect 9496 -140 9580 -106
rect 9754 -140 9838 -106
rect 736 -566 770 -190
rect 994 -566 1028 -190
rect 1252 -566 1286 -190
rect 1510 -566 1544 -190
rect 1768 -566 1802 -190
rect 2026 -566 2060 -190
rect 2284 -566 2318 -190
rect 2542 -566 2576 -190
rect 2800 -566 2834 -190
rect 3058 -566 3092 -190
rect 3316 -566 3350 -190
rect 4032 -566 4066 -190
rect 4290 -566 4324 -190
rect 4548 -566 4582 -190
rect 4806 -566 4840 -190
rect 5064 -566 5098 -190
rect 5322 -566 5356 -190
rect 5580 -566 5614 -190
rect 5838 -566 5872 -190
rect 6096 -566 6130 -190
rect 6354 -566 6388 -190
rect 6612 -566 6646 -190
rect 7328 -566 7362 -190
rect 7586 -566 7620 -190
rect 7844 -566 7878 -190
rect 8102 -566 8136 -190
rect 8360 -566 8394 -190
rect 8618 -566 8652 -190
rect 8876 -566 8910 -190
rect 9134 -566 9168 -190
rect 9392 -566 9426 -190
rect 9650 -566 9684 -190
rect 9908 -566 9942 -190
rect 840 -650 924 -616
rect 1098 -650 1182 -616
rect 1356 -650 1440 -616
rect 1614 -650 1698 -616
rect 1872 -650 1956 -616
rect 2130 -650 2214 -616
rect 2388 -650 2472 -616
rect 2646 -650 2730 -616
rect 2904 -650 2988 -616
rect 3162 -650 3246 -616
rect 4136 -650 4220 -616
rect 4394 -650 4478 -616
rect 4652 -650 4736 -616
rect 4910 -650 4994 -616
rect 5168 -650 5252 -616
rect 5426 -650 5510 -616
rect 5684 -650 5768 -616
rect 5942 -650 6026 -616
rect 6200 -650 6284 -616
rect 6458 -650 6542 -616
rect 7432 -650 7516 -616
rect 7690 -650 7774 -616
rect 7948 -650 8032 -616
rect 8206 -650 8290 -616
rect 8464 -650 8548 -616
rect 8722 -650 8806 -616
rect 8980 -650 9064 -616
rect 9238 -650 9322 -616
rect 9496 -650 9580 -616
rect 9754 -650 9838 -616
rect 442 -1248 826 -1214
rect 1300 -1248 1684 -1214
rect 2158 -1248 2542 -1214
rect 3016 -1248 3400 -1214
rect 3874 -1248 4258 -1214
rect 4732 -1248 5116 -1214
rect 5590 -1248 5974 -1214
rect 6448 -1248 6832 -1214
rect 7306 -1248 7690 -1214
rect 8164 -1248 8548 -1214
rect 9022 -1248 9406 -1214
rect 9880 -1248 10264 -1214
rect 188 -1474 222 -1298
rect 1046 -1474 1080 -1298
rect 1904 -1474 1938 -1298
rect 2762 -1474 2796 -1298
rect 3620 -1474 3654 -1298
rect 4478 -1474 4512 -1298
rect 5336 -1474 5370 -1298
rect 6194 -1474 6228 -1298
rect 7052 -1474 7086 -1298
rect 7910 -1474 7944 -1298
rect 8768 -1474 8802 -1298
rect 9626 -1474 9660 -1298
rect 10484 -1474 10518 -1298
rect 442 -1558 826 -1524
rect 1300 -1558 1684 -1524
rect 2158 -1558 2542 -1524
rect 3016 -1558 3400 -1524
rect 3874 -1558 4258 -1524
rect 4732 -1558 5116 -1524
rect 5590 -1558 5974 -1524
rect 6448 -1558 6832 -1524
rect 7306 -1558 7690 -1524
rect 8164 -1558 8548 -1524
rect 9022 -1558 9406 -1524
rect 9880 -1558 10264 -1524
rect 442 -1788 826 -1754
rect 1300 -1788 1684 -1754
rect 2158 -1788 2542 -1754
rect 3016 -1788 3400 -1754
rect 3874 -1788 4258 -1754
rect 4732 -1788 5116 -1754
rect 5590 -1788 5974 -1754
rect 6448 -1788 6832 -1754
rect 7306 -1788 7690 -1754
rect 8164 -1788 8548 -1754
rect 9022 -1788 9406 -1754
rect 9880 -1788 10264 -1754
rect 188 -2014 222 -1838
rect 1046 -2014 1080 -1838
rect 1904 -2014 1938 -1838
rect 2762 -2014 2796 -1838
rect 3620 -2014 3654 -1838
rect 4478 -2014 4512 -1838
rect 5336 -2014 5370 -1838
rect 6194 -2014 6228 -1838
rect 7052 -2014 7086 -1838
rect 7910 -2014 7944 -1838
rect 8768 -2014 8802 -1838
rect 9626 -2014 9660 -1838
rect 10484 -2014 10518 -1838
rect 442 -2098 826 -2064
rect 1300 -2098 1684 -2064
rect 2158 -2098 2542 -2064
rect 3016 -2098 3400 -2064
rect 3874 -2098 4258 -2064
rect 4732 -2098 5116 -2064
rect 5590 -2098 5974 -2064
rect 6448 -2098 6832 -2064
rect 7306 -2098 7690 -2064
rect 8164 -2098 8548 -2064
rect 9022 -2098 9406 -2064
rect 9880 -2098 10264 -2064
rect 10922 -2762 11022 122
rect -222 -3022 -160 -2922
rect -160 -3022 10860 -2922
rect 10860 -3022 10922 -2922
<< metal1 >>
rect -328 2402 11028 2408
rect -328 2302 -222 2402
rect 10922 2302 11028 2402
rect -328 2296 11028 2302
rect -328 2242 -216 2296
rect -328 778 -322 2242
rect -222 778 -216 2242
rect 384 1996 394 2296
rect 10306 1996 10316 2296
rect 10916 2242 11028 2296
rect 3466 1910 7322 1950
rect 3466 1758 3514 1910
rect 7278 1758 7322 1910
rect 3466 1720 7322 1758
rect -328 724 -216 778
rect 3504 1503 3564 1720
rect 3640 1503 3700 1720
rect 3504 1443 3700 1503
rect 3504 1278 3564 1443
rect 3640 1377 3700 1443
rect 3612 1371 3720 1377
rect 3612 1337 3624 1371
rect 3708 1337 3720 1371
rect 3612 1331 3720 1337
rect 3870 1371 3978 1377
rect 3870 1337 3882 1371
rect 3966 1337 3978 1371
rect 3870 1331 3978 1337
rect 3504 1102 3520 1278
rect 3554 1102 3564 1278
rect 3772 1278 3818 1290
rect 3772 1142 3778 1278
rect 3504 956 3564 1102
rect 3764 1102 3778 1142
rect 3812 1142 3818 1278
rect 4022 1278 4082 1720
rect 4412 1498 4472 1720
rect 4538 1498 4598 1720
rect 4412 1438 4598 1498
rect 4412 1377 4472 1438
rect 4128 1371 4236 1377
rect 4128 1337 4140 1371
rect 4224 1337 4236 1371
rect 4128 1331 4236 1337
rect 4386 1371 4494 1377
rect 4386 1337 4398 1371
rect 4482 1337 4494 1371
rect 4386 1331 4494 1337
rect 4022 1248 4036 1278
rect 3812 1102 3824 1142
rect 3612 1043 3720 1049
rect 3612 1009 3624 1043
rect 3708 1009 3720 1043
rect 3612 1003 3720 1009
rect 3636 956 3696 1003
rect 3504 896 3696 956
rect 3504 724 3564 896
rect 3636 724 3696 896
rect 3764 952 3824 1102
rect 4030 1102 4036 1248
rect 4070 1248 4082 1278
rect 4288 1278 4334 1290
rect 4070 1102 4076 1248
rect 4288 1125 4294 1278
rect 4030 1090 4076 1102
rect 4280 1102 4294 1125
rect 4328 1125 4334 1278
rect 4538 1278 4598 1438
rect 4926 1503 4986 1720
rect 5054 1503 5114 1720
rect 5178 1503 5238 1720
rect 5302 1556 5308 1616
rect 5368 1556 5374 1616
rect 4926 1443 5238 1503
rect 4926 1377 4986 1443
rect 4644 1371 4752 1377
rect 4644 1337 4656 1371
rect 4740 1337 4752 1371
rect 4644 1331 4752 1337
rect 4902 1371 5010 1377
rect 4902 1337 4914 1371
rect 4998 1337 5010 1371
rect 4902 1331 5010 1337
rect 4328 1102 4340 1125
rect 3870 1043 3978 1049
rect 3870 1009 3882 1043
rect 3966 1009 3978 1043
rect 3870 1003 3978 1009
rect 4128 1043 4236 1049
rect 4128 1009 4140 1043
rect 4224 1009 4236 1043
rect 4128 1003 4236 1009
rect 3896 952 3956 1003
rect 4152 952 4212 1003
rect 3764 892 4152 952
rect 4212 892 4218 952
rect 4280 842 4340 1102
rect 4538 1102 4552 1278
rect 4586 1102 4598 1278
rect 4804 1278 4850 1290
rect 4804 1157 4810 1278
rect 4386 1043 4494 1049
rect 4386 1009 4398 1043
rect 4482 1009 4494 1043
rect 4386 1003 4494 1009
rect 4280 776 4340 782
rect 4538 724 4598 1102
rect 4794 1102 4810 1157
rect 4844 1157 4850 1278
rect 5054 1278 5114 1443
rect 5178 1377 5238 1443
rect 5160 1371 5268 1377
rect 5160 1337 5172 1371
rect 5256 1337 5268 1371
rect 5160 1331 5268 1337
rect 4844 1102 4854 1157
rect 4644 1043 4752 1049
rect 4644 1009 4656 1043
rect 4740 1009 4752 1043
rect 4644 1003 4752 1009
rect 4668 952 4728 1003
rect 4662 892 4668 952
rect 4728 892 4734 952
rect 4794 840 4854 1102
rect 5054 1102 5068 1278
rect 5102 1102 5114 1278
rect 5308 1278 5368 1556
rect 5418 1371 5526 1377
rect 5418 1337 5430 1371
rect 5514 1337 5526 1371
rect 5418 1331 5526 1337
rect 5308 1238 5326 1278
rect 4902 1043 5010 1049
rect 4902 1009 4914 1043
rect 4998 1009 5010 1043
rect 4902 1003 5010 1009
rect 4794 774 4854 780
rect 4926 956 4986 1003
rect 5054 956 5114 1102
rect 5320 1102 5326 1238
rect 5360 1238 5368 1278
rect 5568 1278 5628 1720
rect 5958 1497 6018 1720
rect 6086 1497 6146 1720
rect 6218 1497 6278 1720
rect 5958 1437 6278 1497
rect 5958 1377 6018 1437
rect 5676 1371 5784 1377
rect 5676 1337 5688 1371
rect 5772 1337 5784 1371
rect 5676 1331 5784 1337
rect 5934 1371 6042 1377
rect 5934 1337 5946 1371
rect 6030 1337 6042 1371
rect 5934 1331 6042 1337
rect 5568 1248 5584 1278
rect 5360 1102 5366 1238
rect 5320 1090 5366 1102
rect 5578 1102 5584 1248
rect 5618 1248 5628 1278
rect 5836 1278 5882 1290
rect 5618 1102 5624 1248
rect 5836 1140 5842 1278
rect 5578 1090 5624 1102
rect 5826 1102 5842 1140
rect 5876 1140 5882 1278
rect 6086 1278 6146 1437
rect 6218 1377 6278 1437
rect 6340 1434 6346 1494
rect 6406 1434 6412 1494
rect 6192 1371 6300 1377
rect 6192 1337 6204 1371
rect 6288 1337 6300 1371
rect 6192 1331 6300 1337
rect 5876 1102 5886 1140
rect 5160 1043 5268 1049
rect 5160 1009 5172 1043
rect 5256 1009 5268 1043
rect 5160 1003 5268 1009
rect 5418 1043 5526 1049
rect 5418 1009 5430 1043
rect 5514 1009 5526 1043
rect 5418 1003 5526 1009
rect 5676 1043 5784 1049
rect 5676 1009 5688 1043
rect 5772 1009 5784 1043
rect 5676 1003 5784 1009
rect 5182 956 5242 1003
rect 4926 896 5242 956
rect 4926 724 4986 896
rect 5054 724 5114 896
rect 5182 724 5242 896
rect 5440 950 5500 1003
rect 5700 950 5760 1003
rect 5826 950 5886 1102
rect 6086 1102 6100 1278
rect 6134 1102 6146 1278
rect 5934 1043 6042 1049
rect 5934 1009 5946 1043
rect 6030 1009 6042 1043
rect 5934 1003 6042 1009
rect 5440 890 5886 950
rect 5956 950 6016 1003
rect 6086 950 6146 1102
rect 6346 1278 6406 1434
rect 6450 1371 6558 1377
rect 6450 1337 6462 1371
rect 6546 1337 6558 1371
rect 6450 1331 6558 1337
rect 6346 1102 6358 1278
rect 6392 1102 6406 1278
rect 6192 1043 6300 1049
rect 6192 1009 6204 1043
rect 6288 1009 6300 1043
rect 6192 1003 6300 1009
rect 6210 950 6270 1003
rect 5956 890 6270 950
rect 5700 838 5760 890
rect 5700 772 5760 778
rect 5956 724 6016 890
rect 6086 724 6146 890
rect 6210 724 6270 890
rect 6346 948 6406 1102
rect 6602 1278 6662 1720
rect 6988 1496 7048 1720
rect 7118 1496 7178 1720
rect 6988 1436 7178 1496
rect 6988 1377 7048 1436
rect 6708 1371 6816 1377
rect 6708 1337 6720 1371
rect 6804 1337 6816 1371
rect 6708 1331 6816 1337
rect 6966 1371 7074 1377
rect 6966 1337 6978 1371
rect 7062 1337 7074 1371
rect 6966 1331 7074 1337
rect 6602 1102 6616 1278
rect 6650 1102 6662 1278
rect 6868 1278 6914 1290
rect 6868 1148 6874 1278
rect 6450 1043 6558 1049
rect 6450 1009 6462 1043
rect 6546 1009 6558 1043
rect 6450 1003 6558 1009
rect 6472 948 6532 1003
rect 6346 888 6532 948
rect 6602 724 6662 1102
rect 6864 1102 6874 1148
rect 6908 1148 6914 1278
rect 7118 1278 7178 1436
rect 6908 1102 6924 1148
rect 6708 1043 6816 1049
rect 6708 1009 6720 1043
rect 6804 1009 6816 1043
rect 6708 1003 6816 1009
rect 6736 948 6796 1003
rect 6864 948 6924 1102
rect 7118 1102 7132 1278
rect 7166 1102 7178 1278
rect 6966 1043 7074 1049
rect 6966 1009 6978 1043
rect 7062 1009 7074 1043
rect 6966 1003 7074 1009
rect 6736 888 6924 948
rect 6864 836 6924 888
rect 6988 952 7048 1003
rect 7118 952 7178 1102
rect 6988 892 7178 952
rect 6858 776 6864 836
rect 6924 776 6930 836
rect 6988 724 7048 892
rect 7118 724 7178 892
rect 10916 778 10922 2242
rect 11022 778 11028 2242
rect 10916 724 11028 778
rect -328 718 11028 724
rect -328 618 -222 718
rect 10922 618 11028 718
rect -328 612 11028 618
rect 3052 524 3112 530
rect 5700 524 5760 530
rect 8088 524 8148 530
rect 3112 464 5700 524
rect 5760 464 8088 524
rect 3052 458 3112 464
rect 5700 458 5760 464
rect 8088 458 8148 464
rect -328 382 11028 388
rect -328 282 -222 382
rect 10922 282 11028 382
rect -328 276 11028 282
rect -328 122 -216 276
rect -328 -2762 -322 122
rect -222 4 -216 122
rect 726 4 786 276
rect 852 4 912 276
rect 1488 170 1494 230
rect 1554 170 1560 230
rect 2524 170 2530 230
rect 2590 170 2596 230
rect 974 54 980 114
rect 1040 54 1046 114
rect -222 -56 912 4
rect -222 -728 -216 -56
rect 726 -190 786 -56
rect 852 -100 912 -56
rect 828 -106 936 -100
rect 828 -140 840 -106
rect 924 -140 936 -106
rect 828 -146 936 -140
rect 726 -566 736 -190
rect 770 -566 786 -190
rect 980 -190 1040 54
rect 1364 -56 1370 4
rect 1430 -56 1436 4
rect 1370 -100 1430 -56
rect 1086 -106 1194 -100
rect 1086 -140 1098 -106
rect 1182 -140 1194 -106
rect 1086 -146 1194 -140
rect 1344 -106 1452 -100
rect 1344 -140 1356 -106
rect 1440 -140 1452 -106
rect 1344 -146 1452 -140
rect 980 -240 994 -190
rect 726 -728 786 -566
rect 988 -566 994 -240
rect 1028 -240 1040 -190
rect 1246 -190 1292 -178
rect 1028 -566 1034 -240
rect 1246 -546 1252 -190
rect 988 -578 1034 -566
rect 1240 -566 1252 -546
rect 1286 -546 1292 -190
rect 1494 -190 1554 170
rect 2006 54 2012 114
rect 2072 54 2078 114
rect 1618 -56 1624 4
rect 1684 -56 1690 4
rect 1624 -100 1684 -56
rect 1602 -106 1710 -100
rect 1602 -140 1614 -106
rect 1698 -140 1710 -106
rect 1602 -146 1710 -140
rect 1860 -106 1968 -100
rect 1860 -140 1872 -106
rect 1956 -140 1968 -106
rect 1860 -146 1968 -140
rect 1494 -236 1510 -190
rect 1286 -566 1300 -546
rect 828 -616 936 -610
rect 828 -650 840 -616
rect 924 -650 936 -616
rect 828 -656 936 -650
rect 1086 -616 1194 -610
rect 1086 -650 1098 -616
rect 1182 -650 1194 -616
rect 1086 -656 1194 -650
rect 852 -728 912 -656
rect 1110 -726 1170 -656
rect -222 -788 912 -728
rect 1104 -786 1110 -726
rect 1170 -786 1176 -726
rect -222 -2762 -216 -788
rect 26 -896 32 -836
rect 92 -896 98 -836
rect 32 -2170 92 -896
rect 172 -1082 232 -788
rect 1240 -836 1300 -566
rect 1504 -566 1510 -236
rect 1544 -236 1554 -190
rect 1762 -190 1808 -178
rect 1544 -566 1550 -236
rect 1762 -546 1768 -190
rect 1504 -578 1550 -566
rect 1752 -566 1768 -546
rect 1802 -546 1808 -190
rect 2012 -190 2072 54
rect 2390 -56 2396 4
rect 2456 -56 2462 4
rect 2396 -100 2456 -56
rect 2118 -106 2226 -100
rect 2118 -140 2130 -106
rect 2214 -140 2226 -106
rect 2118 -146 2226 -140
rect 2376 -106 2484 -100
rect 2376 -140 2388 -106
rect 2472 -140 2484 -106
rect 2376 -146 2484 -140
rect 2396 -150 2456 -146
rect 2012 -250 2026 -190
rect 1802 -566 1812 -546
rect 1344 -616 1452 -610
rect 1344 -650 1356 -616
rect 1440 -650 1452 -616
rect 1344 -656 1452 -650
rect 1602 -616 1710 -610
rect 1602 -650 1614 -616
rect 1698 -650 1710 -616
rect 1602 -656 1710 -650
rect 1752 -836 1812 -566
rect 2020 -566 2026 -250
rect 2060 -250 2072 -190
rect 2278 -190 2324 -178
rect 2060 -566 2066 -250
rect 2278 -542 2284 -190
rect 2020 -578 2066 -566
rect 2272 -566 2284 -542
rect 2318 -542 2324 -190
rect 2530 -190 2590 170
rect 3042 54 3048 114
rect 3108 54 3114 114
rect 2652 -56 2658 4
rect 2718 -56 2724 4
rect 2658 -100 2718 -56
rect 2634 -106 2742 -100
rect 2634 -140 2646 -106
rect 2730 -140 2742 -106
rect 2634 -146 2742 -140
rect 2892 -106 3000 -100
rect 2892 -140 2904 -106
rect 2988 -140 3000 -106
rect 2892 -146 3000 -140
rect 2530 -240 2542 -190
rect 2318 -566 2332 -542
rect 1860 -616 1968 -610
rect 1860 -650 1872 -616
rect 1956 -650 1968 -616
rect 1860 -656 1968 -650
rect 2118 -616 2226 -610
rect 2118 -650 2130 -616
rect 2214 -650 2226 -616
rect 2118 -656 2226 -650
rect 1886 -726 1946 -656
rect 2140 -726 2200 -656
rect 1880 -786 1886 -726
rect 1946 -786 1952 -726
rect 2134 -786 2140 -726
rect 2200 -786 2206 -726
rect 2272 -836 2332 -566
rect 2536 -566 2542 -240
rect 2576 -240 2590 -190
rect 2794 -190 2840 -178
rect 2576 -566 2582 -240
rect 2794 -542 2800 -190
rect 2536 -578 2582 -566
rect 2788 -566 2800 -542
rect 2834 -542 2840 -190
rect 3048 -190 3108 54
rect 3172 4 3232 276
rect 3306 4 3366 276
rect 4022 4 4082 276
rect 4146 4 4206 276
rect 4784 176 4790 236
rect 4850 176 4856 236
rect 5820 176 5826 236
rect 5886 176 5892 236
rect 4270 60 4276 120
rect 4336 60 4342 120
rect 3172 -56 4206 4
rect 3172 -100 3232 -56
rect 3150 -106 3258 -100
rect 3150 -140 3162 -106
rect 3246 -140 3258 -106
rect 3150 -146 3258 -140
rect 3048 -246 3058 -190
rect 2834 -566 2848 -542
rect 2376 -616 2484 -610
rect 2376 -650 2388 -616
rect 2472 -650 2484 -616
rect 2376 -656 2484 -650
rect 2634 -616 2742 -610
rect 2634 -650 2646 -616
rect 2730 -650 2742 -616
rect 2634 -656 2742 -650
rect 2788 -836 2848 -566
rect 3052 -566 3058 -246
rect 3092 -246 3108 -190
rect 3306 -190 3366 -56
rect 3092 -566 3098 -246
rect 3052 -578 3098 -566
rect 3306 -566 3316 -190
rect 3350 -566 3366 -190
rect 2892 -616 3000 -610
rect 2892 -650 2904 -616
rect 2988 -650 3000 -616
rect 2892 -656 3000 -650
rect 3150 -616 3258 -610
rect 3150 -650 3162 -616
rect 3246 -650 3258 -616
rect 3150 -656 3258 -650
rect 2918 -726 2978 -656
rect 2912 -786 2918 -726
rect 2978 -786 2984 -726
rect 3172 -728 3232 -656
rect 3306 -728 3366 -566
rect 4022 -190 4082 -56
rect 4146 -100 4206 -56
rect 4124 -106 4232 -100
rect 4124 -140 4136 -106
rect 4220 -140 4232 -106
rect 4124 -146 4232 -140
rect 4022 -566 4032 -190
rect 4066 -566 4082 -190
rect 4276 -190 4336 60
rect 4660 -50 4666 10
rect 4726 -50 4732 10
rect 4666 -100 4726 -50
rect 4382 -106 4490 -100
rect 4382 -140 4394 -106
rect 4478 -140 4490 -106
rect 4382 -146 4490 -140
rect 4640 -106 4748 -100
rect 4640 -140 4652 -106
rect 4736 -140 4748 -106
rect 4640 -146 4748 -140
rect 4276 -234 4290 -190
rect 4022 -728 4082 -566
rect 4284 -566 4290 -234
rect 4324 -234 4336 -190
rect 4542 -190 4588 -178
rect 4324 -566 4330 -234
rect 4542 -540 4548 -190
rect 4284 -578 4330 -566
rect 4536 -566 4548 -540
rect 4582 -540 4588 -190
rect 4790 -190 4850 176
rect 5302 60 5308 120
rect 5368 60 5374 120
rect 4914 -50 4920 10
rect 4980 -50 4986 10
rect 4920 -100 4980 -50
rect 4898 -106 5006 -100
rect 4898 -140 4910 -106
rect 4994 -140 5006 -106
rect 4898 -146 5006 -140
rect 5156 -106 5264 -100
rect 5156 -140 5168 -106
rect 5252 -140 5264 -106
rect 5156 -146 5264 -140
rect 4790 -230 4806 -190
rect 4800 -478 4806 -230
rect 4582 -566 4596 -540
rect 4124 -616 4232 -610
rect 4124 -650 4136 -616
rect 4220 -650 4232 -616
rect 4124 -656 4232 -650
rect 4382 -616 4490 -610
rect 4382 -650 4394 -616
rect 4478 -650 4490 -616
rect 4382 -656 4490 -650
rect 4148 -728 4208 -656
rect 4406 -720 4466 -656
rect 1746 -896 1752 -836
rect 1812 -896 1818 -836
rect 2266 -896 2272 -836
rect 2332 -896 2338 -836
rect 2782 -896 2788 -836
rect 2848 -896 2854 -836
rect 1240 -902 1300 -896
rect 2918 -958 2978 -786
rect 3172 -788 4208 -728
rect 4400 -780 4406 -720
rect 4466 -780 4472 -720
rect 2912 -1018 2918 -958
rect 2978 -1018 2984 -958
rect 172 -1142 654 -1082
rect 1024 -1142 1030 -1082
rect 1090 -1142 1096 -1082
rect 172 -1298 232 -1142
rect 594 -1208 654 -1142
rect 430 -1214 838 -1208
rect 430 -1248 442 -1214
rect 826 -1248 838 -1214
rect 430 -1254 838 -1248
rect 172 -1474 188 -1298
rect 222 -1474 232 -1298
rect 1030 -1298 1090 -1142
rect 1288 -1214 1696 -1208
rect 1288 -1248 1300 -1214
rect 1684 -1248 1696 -1214
rect 1288 -1254 1696 -1248
rect 2146 -1214 2554 -1208
rect 2146 -1248 2158 -1214
rect 2542 -1248 2554 -1214
rect 2146 -1254 2554 -1248
rect 3004 -1214 3412 -1208
rect 3004 -1248 3016 -1214
rect 3400 -1248 3412 -1214
rect 3004 -1254 3412 -1248
rect 1030 -1336 1046 -1298
rect 172 -1632 232 -1474
rect 1040 -1474 1046 -1336
rect 1080 -1336 1090 -1298
rect 1898 -1298 1944 -1286
rect 1080 -1474 1086 -1336
rect 1898 -1394 1904 -1298
rect 1040 -1486 1086 -1474
rect 1890 -1474 1904 -1394
rect 1938 -1394 1944 -1298
rect 2756 -1298 2802 -1286
rect 1938 -1474 1950 -1394
rect 2756 -1424 2762 -1298
rect 430 -1524 838 -1518
rect 430 -1558 442 -1524
rect 826 -1558 838 -1524
rect 430 -1564 838 -1558
rect 1288 -1524 1696 -1518
rect 1288 -1558 1300 -1524
rect 1684 -1558 1696 -1524
rect 1288 -1564 1696 -1558
rect 596 -1632 656 -1564
rect 1456 -1626 1516 -1564
rect 172 -1692 656 -1632
rect 1026 -1686 1032 -1626
rect 1092 -1686 1516 -1626
rect 172 -1838 232 -1692
rect 596 -1748 656 -1692
rect 430 -1754 838 -1748
rect 430 -1788 442 -1754
rect 826 -1788 838 -1754
rect 430 -1794 838 -1788
rect 172 -2014 188 -1838
rect 222 -2014 232 -1838
rect 1032 -1838 1092 -1686
rect 1456 -1748 1516 -1686
rect 1288 -1754 1696 -1748
rect 1288 -1788 1300 -1754
rect 1684 -1788 1696 -1754
rect 1288 -1794 1696 -1788
rect 1032 -1890 1046 -1838
rect 172 -2162 232 -2014
rect 1040 -2014 1046 -1890
rect 1080 -1890 1092 -1838
rect 1890 -1838 1950 -1474
rect 2748 -1474 2762 -1424
rect 2796 -1424 2802 -1298
rect 3606 -1298 3666 -788
rect 4536 -830 4596 -566
rect 4798 -566 4806 -478
rect 4840 -230 4850 -190
rect 5058 -190 5104 -178
rect 4840 -478 4846 -230
rect 4840 -566 4858 -478
rect 5058 -540 5064 -190
rect 4640 -616 4748 -610
rect 4640 -650 4652 -616
rect 4736 -650 4748 -616
rect 4640 -656 4748 -650
rect 4536 -1082 4596 -890
rect 4798 -958 4858 -566
rect 5048 -566 5064 -540
rect 5098 -540 5104 -190
rect 5308 -190 5368 60
rect 5686 -50 5692 10
rect 5752 -50 5758 10
rect 5692 -100 5752 -50
rect 5414 -106 5522 -100
rect 5414 -140 5426 -106
rect 5510 -140 5522 -106
rect 5414 -146 5522 -140
rect 5672 -106 5780 -100
rect 5672 -140 5684 -106
rect 5768 -140 5780 -106
rect 5672 -146 5780 -140
rect 5308 -244 5322 -190
rect 5098 -566 5108 -540
rect 4898 -616 5006 -610
rect 4898 -650 4910 -616
rect 4994 -650 5006 -616
rect 4898 -656 5006 -650
rect 5048 -830 5108 -566
rect 5316 -566 5322 -244
rect 5356 -244 5368 -190
rect 5574 -190 5620 -178
rect 5356 -566 5362 -244
rect 5574 -536 5580 -190
rect 5316 -578 5362 -566
rect 5568 -566 5580 -536
rect 5614 -536 5620 -190
rect 5826 -190 5886 176
rect 6338 60 6344 120
rect 6404 60 6410 120
rect 5948 -50 5954 10
rect 6014 -50 6020 10
rect 5954 -100 6014 -50
rect 5930 -106 6038 -100
rect 5930 -140 5942 -106
rect 6026 -140 6038 -106
rect 5930 -146 6038 -140
rect 6188 -106 6296 -100
rect 6188 -140 6200 -106
rect 6284 -140 6296 -106
rect 6188 -146 6296 -140
rect 5826 -234 5838 -190
rect 5614 -566 5628 -536
rect 5156 -616 5264 -610
rect 5156 -650 5168 -616
rect 5252 -650 5264 -616
rect 5156 -656 5264 -650
rect 5414 -616 5522 -610
rect 5414 -650 5426 -616
rect 5510 -650 5522 -616
rect 5414 -656 5522 -650
rect 5182 -720 5242 -656
rect 5436 -720 5496 -656
rect 5176 -780 5182 -720
rect 5242 -780 5248 -720
rect 5430 -780 5436 -720
rect 5496 -780 5502 -720
rect 5568 -830 5628 -566
rect 5832 -566 5838 -234
rect 5872 -234 5886 -190
rect 6090 -190 6136 -178
rect 5872 -566 5878 -234
rect 6090 -536 6096 -190
rect 5832 -578 5878 -566
rect 6084 -566 6096 -536
rect 6130 -536 6136 -190
rect 6344 -190 6404 60
rect 6470 10 6530 276
rect 6602 10 6662 276
rect 7318 10 7378 276
rect 7442 10 7502 276
rect 8080 170 8086 230
rect 8146 170 8152 230
rect 9116 170 9122 230
rect 9182 170 9188 230
rect 7566 54 7572 114
rect 7632 54 7638 114
rect 6470 -50 7502 10
rect 6470 -100 6530 -50
rect 6446 -106 6554 -100
rect 6446 -140 6458 -106
rect 6542 -140 6554 -106
rect 6446 -146 6554 -140
rect 6344 -240 6354 -190
rect 6130 -566 6144 -536
rect 5672 -616 5780 -610
rect 5672 -650 5684 -616
rect 5768 -650 5780 -616
rect 5672 -656 5780 -650
rect 5930 -616 6038 -610
rect 5930 -650 5942 -616
rect 6026 -650 6038 -616
rect 5930 -656 6038 -650
rect 6084 -830 6144 -566
rect 6348 -566 6354 -240
rect 6388 -240 6404 -190
rect 6602 -190 6662 -50
rect 6388 -566 6394 -240
rect 6348 -578 6394 -566
rect 6602 -566 6612 -190
rect 6646 -566 6662 -190
rect 6188 -616 6296 -610
rect 6188 -650 6200 -616
rect 6284 -650 6296 -616
rect 6188 -656 6296 -650
rect 6446 -616 6554 -610
rect 6446 -650 6458 -616
rect 6542 -650 6554 -616
rect 6446 -656 6554 -650
rect 6214 -720 6274 -656
rect 6208 -780 6214 -720
rect 6274 -780 6280 -720
rect 6468 -722 6528 -656
rect 6602 -722 6662 -566
rect 7318 -190 7378 -50
rect 7442 -100 7502 -50
rect 7420 -106 7528 -100
rect 7420 -140 7432 -106
rect 7516 -140 7528 -106
rect 7420 -146 7528 -140
rect 7318 -566 7328 -190
rect 7362 -566 7378 -190
rect 7572 -190 7632 54
rect 7956 -56 7962 4
rect 8022 -56 8028 4
rect 7962 -100 8022 -56
rect 7678 -106 7786 -100
rect 7678 -140 7690 -106
rect 7774 -140 7786 -106
rect 7678 -146 7786 -140
rect 7936 -106 8044 -100
rect 7936 -140 7948 -106
rect 8032 -140 8044 -106
rect 7936 -146 8044 -140
rect 7572 -240 7586 -190
rect 7318 -722 7378 -566
rect 7580 -566 7586 -240
rect 7620 -240 7632 -190
rect 7838 -190 7884 -178
rect 7620 -566 7626 -240
rect 7838 -546 7844 -190
rect 7580 -578 7626 -566
rect 7832 -566 7844 -546
rect 7878 -546 7884 -190
rect 8086 -190 8146 170
rect 8598 54 8604 114
rect 8664 54 8670 114
rect 8210 -56 8216 4
rect 8276 -56 8282 4
rect 8216 -100 8276 -56
rect 8194 -106 8302 -100
rect 8194 -140 8206 -106
rect 8290 -140 8302 -106
rect 8194 -146 8302 -140
rect 8452 -106 8560 -100
rect 8452 -140 8464 -106
rect 8548 -140 8560 -106
rect 8452 -146 8560 -140
rect 8086 -236 8102 -190
rect 7878 -566 7892 -546
rect 7420 -616 7528 -610
rect 7420 -650 7432 -616
rect 7516 -650 7528 -616
rect 7420 -656 7528 -650
rect 7678 -616 7786 -610
rect 7678 -650 7690 -616
rect 7774 -650 7786 -616
rect 7678 -656 7786 -650
rect 7444 -722 7504 -656
rect 6468 -782 7504 -722
rect 7702 -726 7762 -656
rect 5042 -890 5048 -830
rect 5108 -890 5114 -830
rect 5562 -890 5568 -830
rect 5628 -890 5634 -830
rect 6078 -890 6084 -830
rect 6144 -890 6150 -830
rect 4792 -1018 4798 -958
rect 4858 -1018 4864 -958
rect 4458 -1142 4464 -1082
rect 4524 -1142 4596 -1082
rect 4894 -1140 5818 -1080
rect 3862 -1214 4270 -1208
rect 3862 -1248 3874 -1214
rect 4258 -1248 4270 -1214
rect 3862 -1254 4270 -1248
rect 2796 -1474 2808 -1424
rect 2146 -1524 2554 -1518
rect 2146 -1558 2158 -1524
rect 2542 -1558 2554 -1524
rect 2146 -1564 2554 -1558
rect 2314 -1626 2374 -1564
rect 2748 -1626 2808 -1474
rect 3606 -1474 3620 -1298
rect 3654 -1474 3666 -1298
rect 4464 -1298 4524 -1142
rect 4894 -1208 4954 -1140
rect 4720 -1214 5128 -1208
rect 4720 -1248 4732 -1214
rect 5116 -1248 5128 -1214
rect 4720 -1254 5128 -1248
rect 4464 -1340 4478 -1298
rect 3004 -1524 3412 -1518
rect 3004 -1558 3016 -1524
rect 3400 -1558 3412 -1524
rect 3004 -1564 3412 -1558
rect 3178 -1626 3238 -1564
rect 2308 -1682 2314 -1626
rect 2374 -1682 2380 -1626
rect 2308 -1686 2380 -1682
rect 2742 -1686 2748 -1626
rect 2808 -1686 2814 -1626
rect 2314 -1748 2374 -1686
rect 2146 -1754 2554 -1748
rect 2146 -1788 2158 -1754
rect 2542 -1788 2554 -1754
rect 2146 -1794 2554 -1788
rect 1080 -2014 1086 -1890
rect 1040 -2026 1086 -2014
rect 1890 -2014 1904 -1838
rect 1938 -2014 1950 -1838
rect 2748 -1838 2808 -1686
rect 3178 -1748 3238 -1682
rect 3004 -1754 3412 -1748
rect 3004 -1788 3016 -1754
rect 3400 -1788 3412 -1754
rect 3004 -1794 3412 -1788
rect 2748 -1866 2762 -1838
rect 430 -2064 838 -2058
rect 430 -2098 442 -2064
rect 826 -2098 838 -2064
rect 430 -2104 838 -2098
rect 1288 -2064 1696 -2058
rect 1288 -2098 1300 -2064
rect 1684 -2098 1696 -2064
rect 1288 -2104 1696 -2098
rect 592 -2162 652 -2104
rect 26 -2230 32 -2170
rect 92 -2230 98 -2170
rect 172 -2222 652 -2162
rect 172 -2336 232 -2222
rect 592 -2336 652 -2222
rect 1890 -2336 1950 -2014
rect 2756 -2014 2762 -1866
rect 2796 -1866 2808 -1838
rect 3606 -1838 3666 -1474
rect 4472 -1474 4478 -1340
rect 4512 -1340 4524 -1298
rect 5320 -1298 5380 -1140
rect 5758 -1208 5818 -1140
rect 5578 -1214 5986 -1208
rect 5578 -1248 5590 -1214
rect 5974 -1248 5986 -1214
rect 5578 -1254 5986 -1248
rect 6436 -1214 6844 -1208
rect 6436 -1248 6448 -1214
rect 6832 -1248 6844 -1214
rect 6436 -1254 6844 -1248
rect 4512 -1474 4518 -1340
rect 4472 -1486 4518 -1474
rect 5320 -1474 5336 -1298
rect 5370 -1474 5380 -1298
rect 6188 -1298 6234 -1286
rect 6188 -1426 6194 -1298
rect 3862 -1524 4270 -1518
rect 3862 -1558 3874 -1524
rect 4258 -1558 4270 -1524
rect 3862 -1564 4270 -1558
rect 4720 -1524 5128 -1518
rect 4720 -1558 4732 -1524
rect 5116 -1558 5128 -1524
rect 4720 -1564 5128 -1558
rect 4038 -1626 4098 -1564
rect 4896 -1624 4956 -1564
rect 5320 -1624 5380 -1474
rect 6184 -1474 6194 -1426
rect 6228 -1426 6234 -1298
rect 7038 -1298 7098 -782
rect 7696 -786 7702 -726
rect 7762 -786 7768 -726
rect 7832 -836 7892 -566
rect 8096 -566 8102 -236
rect 8136 -236 8146 -190
rect 8354 -190 8400 -178
rect 8136 -566 8142 -236
rect 8354 -546 8360 -190
rect 8096 -578 8142 -566
rect 8344 -566 8360 -546
rect 8394 -546 8400 -190
rect 8604 -190 8664 54
rect 8982 -56 8988 4
rect 9048 -56 9054 4
rect 8988 -100 9048 -56
rect 8710 -106 8818 -100
rect 8710 -140 8722 -106
rect 8806 -140 8818 -106
rect 8710 -146 8818 -140
rect 8968 -106 9076 -100
rect 8968 -140 8980 -106
rect 9064 -140 9076 -106
rect 8968 -146 9076 -140
rect 8988 -150 9048 -146
rect 8604 -250 8618 -190
rect 8394 -566 8404 -546
rect 7936 -616 8044 -610
rect 7936 -650 7948 -616
rect 8032 -650 8044 -616
rect 7936 -656 8044 -650
rect 8194 -616 8302 -610
rect 8194 -650 8206 -616
rect 8290 -650 8302 -616
rect 8194 -656 8302 -650
rect 8344 -836 8404 -566
rect 8612 -566 8618 -250
rect 8652 -250 8664 -190
rect 8870 -190 8916 -178
rect 8652 -566 8658 -250
rect 8870 -542 8876 -190
rect 8612 -578 8658 -566
rect 8864 -566 8876 -542
rect 8910 -542 8916 -190
rect 9122 -190 9182 170
rect 9634 54 9640 114
rect 9700 54 9706 114
rect 9244 -56 9250 4
rect 9310 -56 9316 4
rect 9250 -100 9310 -56
rect 9226 -106 9334 -100
rect 9226 -140 9238 -106
rect 9322 -140 9334 -106
rect 9226 -146 9334 -140
rect 9484 -106 9592 -100
rect 9484 -140 9496 -106
rect 9580 -140 9592 -106
rect 9484 -146 9592 -140
rect 9122 -240 9134 -190
rect 8910 -566 8924 -542
rect 8452 -616 8560 -610
rect 8452 -650 8464 -616
rect 8548 -650 8560 -616
rect 8452 -656 8560 -650
rect 8710 -616 8818 -610
rect 8710 -650 8722 -616
rect 8806 -650 8818 -616
rect 8710 -656 8818 -650
rect 8478 -726 8538 -656
rect 8732 -726 8792 -656
rect 8472 -786 8478 -726
rect 8538 -786 8544 -726
rect 8726 -786 8732 -726
rect 8792 -786 8798 -726
rect 8864 -836 8924 -566
rect 9128 -566 9134 -240
rect 9168 -240 9182 -190
rect 9386 -190 9432 -178
rect 9168 -566 9174 -240
rect 9386 -542 9392 -190
rect 9128 -578 9174 -566
rect 9380 -566 9392 -542
rect 9426 -542 9432 -190
rect 9640 -190 9700 54
rect 9766 2 9826 276
rect 9898 2 9958 276
rect 10916 122 11028 276
rect 10916 2 10922 122
rect 9766 -58 10922 2
rect 9766 -100 9826 -58
rect 9742 -106 9850 -100
rect 9742 -140 9754 -106
rect 9838 -140 9850 -106
rect 9742 -146 9850 -140
rect 9640 -246 9650 -190
rect 9426 -566 9440 -542
rect 8968 -616 9076 -610
rect 8968 -650 8980 -616
rect 9064 -650 9076 -616
rect 8968 -656 9076 -650
rect 9226 -616 9334 -610
rect 9226 -650 9238 -616
rect 9322 -650 9334 -616
rect 9226 -656 9334 -650
rect 9380 -836 9440 -566
rect 9644 -566 9650 -246
rect 9684 -246 9700 -190
rect 9898 -190 9958 -58
rect 9684 -566 9690 -246
rect 9644 -578 9690 -566
rect 9898 -566 9908 -190
rect 9942 -566 9958 -190
rect 9484 -616 9592 -610
rect 9484 -650 9496 -616
rect 9580 -650 9592 -616
rect 9484 -656 9592 -650
rect 9742 -616 9850 -610
rect 9742 -650 9754 -616
rect 9838 -650 9850 -616
rect 9742 -656 9850 -650
rect 9510 -726 9570 -656
rect 9504 -786 9510 -726
rect 9570 -786 9576 -726
rect 9764 -728 9824 -656
rect 9898 -728 9958 -566
rect 10916 -728 10922 -58
rect 9764 -788 10922 -728
rect 7826 -896 7832 -836
rect 7892 -896 7898 -836
rect 8338 -896 8344 -836
rect 8404 -896 8410 -836
rect 8858 -896 8864 -836
rect 8924 -896 8930 -836
rect 9374 -896 9380 -836
rect 9440 -896 9446 -836
rect 9608 -1026 9614 -966
rect 9674 -1026 9680 -966
rect 7294 -1214 7702 -1208
rect 7294 -1248 7306 -1214
rect 7690 -1248 7702 -1214
rect 7294 -1254 7702 -1248
rect 8152 -1214 8560 -1208
rect 8152 -1248 8164 -1214
rect 8548 -1248 8560 -1214
rect 8152 -1254 8560 -1248
rect 9010 -1214 9418 -1208
rect 9010 -1248 9022 -1214
rect 9406 -1248 9418 -1214
rect 9010 -1254 9418 -1248
rect 6228 -1474 6244 -1426
rect 5578 -1524 5986 -1518
rect 5578 -1558 5590 -1524
rect 5974 -1558 5986 -1524
rect 5578 -1564 5986 -1558
rect 5756 -1624 5816 -1564
rect 4038 -1748 4098 -1682
rect 4462 -1686 4468 -1626
rect 4528 -1686 4534 -1626
rect 4896 -1684 5816 -1624
rect 6184 -1626 6244 -1474
rect 7038 -1474 7052 -1298
rect 7086 -1474 7098 -1298
rect 7904 -1298 7950 -1286
rect 7904 -1410 7910 -1298
rect 6436 -1524 6844 -1518
rect 6436 -1558 6448 -1524
rect 6832 -1558 6844 -1524
rect 6436 -1564 6844 -1558
rect 6610 -1626 6670 -1564
rect 3862 -1754 4270 -1748
rect 3862 -1788 3874 -1754
rect 4258 -1788 4270 -1754
rect 3862 -1794 4270 -1788
rect 2796 -2014 2802 -1866
rect 2756 -2026 2802 -2014
rect 3606 -2014 3620 -1838
rect 3654 -2014 3666 -1838
rect 4468 -1838 4528 -1686
rect 4896 -1748 4956 -1684
rect 4720 -1754 5128 -1748
rect 4720 -1788 4732 -1754
rect 5116 -1788 5128 -1754
rect 4720 -1794 5128 -1788
rect 4468 -1890 4478 -1838
rect 2146 -2064 2554 -2058
rect 2146 -2098 2158 -2064
rect 2542 -2098 2554 -2064
rect 2146 -2104 2554 -2098
rect 3004 -2064 3412 -2058
rect 3004 -2098 3016 -2064
rect 3400 -2098 3412 -2064
rect 3004 -2104 3412 -2098
rect 3606 -2336 3666 -2014
rect 4472 -2014 4478 -1890
rect 4512 -1890 4528 -1838
rect 5320 -1838 5380 -1684
rect 5756 -1748 5816 -1684
rect 6178 -1686 6184 -1626
rect 6244 -1686 6250 -1626
rect 6604 -1682 6610 -1626
rect 6670 -1682 6676 -1626
rect 6604 -1686 6676 -1682
rect 6610 -1748 6670 -1686
rect 5578 -1754 5986 -1748
rect 5578 -1788 5590 -1754
rect 5974 -1788 5986 -1754
rect 5578 -1794 5986 -1788
rect 6436 -1754 6844 -1748
rect 6436 -1788 6448 -1754
rect 6832 -1788 6844 -1754
rect 6436 -1794 6844 -1788
rect 4512 -2014 4518 -1890
rect 4472 -2026 4518 -2014
rect 5320 -2014 5336 -1838
rect 5370 -2014 5380 -1838
rect 6188 -1838 6234 -1826
rect 6188 -1984 6194 -1838
rect 3862 -2064 4270 -2058
rect 3862 -2098 3874 -2064
rect 4258 -2098 4270 -2064
rect 3862 -2104 4270 -2098
rect 4720 -2064 5128 -2058
rect 4720 -2098 4732 -2064
rect 5116 -2098 5128 -2064
rect 4720 -2104 5128 -2098
rect 4894 -2168 4954 -2104
rect 5320 -2168 5380 -2014
rect 6180 -2014 6194 -1984
rect 6228 -1984 6234 -1838
rect 7038 -1838 7098 -1474
rect 7896 -1474 7910 -1410
rect 7944 -1410 7950 -1298
rect 8762 -1298 8808 -1286
rect 7944 -1474 7956 -1410
rect 8762 -1418 8768 -1298
rect 7294 -1524 7702 -1518
rect 7294 -1558 7306 -1524
rect 7690 -1558 7702 -1524
rect 7294 -1564 7702 -1558
rect 7468 -1626 7528 -1564
rect 7896 -1626 7956 -1474
rect 8756 -1474 8768 -1418
rect 8802 -1418 8808 -1298
rect 9614 -1298 9674 -1026
rect 10044 -1096 10104 -788
rect 10468 -1096 10528 -788
rect 10594 -896 10600 -836
rect 10660 -896 10666 -836
rect 10044 -1156 10528 -1096
rect 10044 -1208 10104 -1156
rect 9868 -1214 10276 -1208
rect 9868 -1248 9880 -1214
rect 10264 -1248 10276 -1214
rect 9868 -1254 10276 -1248
rect 9614 -1332 9626 -1298
rect 8802 -1474 8816 -1418
rect 8152 -1524 8560 -1518
rect 8152 -1558 8164 -1524
rect 8548 -1558 8560 -1524
rect 8152 -1564 8560 -1558
rect 8322 -1626 8382 -1564
rect 7468 -1748 7528 -1682
rect 7890 -1686 7896 -1626
rect 7956 -1686 7962 -1626
rect 7294 -1754 7702 -1748
rect 7294 -1788 7306 -1754
rect 7690 -1788 7702 -1754
rect 7294 -1794 7702 -1788
rect 6228 -2014 6240 -1984
rect 5578 -2064 5986 -2058
rect 5578 -2098 5590 -2064
rect 5974 -2098 5986 -2064
rect 5578 -2104 5986 -2098
rect 5756 -2168 5816 -2104
rect 4894 -2228 5816 -2168
rect 6180 -2170 6240 -2014
rect 7038 -2014 7052 -1838
rect 7086 -2014 7098 -1838
rect 7896 -1838 7956 -1686
rect 8322 -1748 8382 -1682
rect 8152 -1754 8560 -1748
rect 8152 -1788 8164 -1754
rect 8548 -1788 8560 -1754
rect 8152 -1794 8560 -1788
rect 7896 -1880 7910 -1838
rect 6436 -2064 6844 -2058
rect 6436 -2098 6448 -2064
rect 6832 -2098 6844 -2064
rect 6436 -2104 6844 -2098
rect 4894 -2336 4954 -2228
rect 5320 -2336 5380 -2228
rect 5756 -2336 5816 -2228
rect 6174 -2230 6180 -2170
rect 6240 -2230 6246 -2170
rect 7038 -2336 7098 -2014
rect 7904 -2014 7910 -1880
rect 7944 -1880 7956 -1838
rect 8756 -1838 8816 -1474
rect 9620 -1474 9626 -1332
rect 9660 -1332 9674 -1298
rect 10468 -1298 10528 -1156
rect 9660 -1474 9666 -1332
rect 9620 -1486 9666 -1474
rect 10468 -1474 10484 -1298
rect 10518 -1474 10528 -1298
rect 9010 -1524 9418 -1518
rect 9010 -1558 9022 -1524
rect 9406 -1558 9418 -1524
rect 9010 -1564 9418 -1558
rect 9868 -1524 10276 -1518
rect 9868 -1558 9880 -1524
rect 10264 -1558 10276 -1524
rect 9868 -1564 10276 -1558
rect 9186 -1620 9246 -1564
rect 9186 -1626 9248 -1620
rect 9186 -1686 9188 -1626
rect 9186 -1692 9248 -1686
rect 10042 -1630 10102 -1564
rect 10468 -1630 10528 -1474
rect 10042 -1690 10528 -1630
rect 9186 -1748 9246 -1692
rect 10042 -1748 10102 -1690
rect 9010 -1754 9418 -1748
rect 9010 -1788 9022 -1754
rect 9406 -1788 9418 -1754
rect 9010 -1794 9418 -1788
rect 9868 -1754 10276 -1748
rect 9868 -1788 9880 -1754
rect 10264 -1788 10276 -1754
rect 9868 -1794 10276 -1788
rect 7944 -2014 7950 -1880
rect 7904 -2026 7950 -2014
rect 8756 -2014 8768 -1838
rect 8802 -2014 8816 -1838
rect 9620 -1838 9666 -1826
rect 9620 -1982 9626 -1838
rect 7294 -2064 7702 -2058
rect 7294 -2098 7306 -2064
rect 7690 -2098 7702 -2064
rect 7294 -2104 7702 -2098
rect 8152 -2064 8560 -2058
rect 8152 -2098 8164 -2064
rect 8548 -2098 8560 -2064
rect 8152 -2104 8560 -2098
rect 8756 -2336 8816 -2014
rect 9612 -2014 9626 -1982
rect 9660 -1982 9666 -1838
rect 10468 -1838 10528 -1690
rect 9660 -2014 9672 -1982
rect 9010 -2064 9418 -2058
rect 9010 -2098 9022 -2064
rect 9406 -2098 9418 -2064
rect 9010 -2104 9418 -2098
rect 9612 -2164 9672 -2014
rect 10468 -2014 10484 -1838
rect 10518 -2014 10528 -1838
rect 9868 -2064 10276 -2058
rect 9868 -2098 9880 -2064
rect 10264 -2098 10276 -2064
rect 9868 -2104 10276 -2098
rect 10044 -2164 10104 -2104
rect 10468 -2164 10528 -2014
rect 10600 -2164 10660 -896
rect 9606 -2224 9612 -2164
rect 9672 -2224 9678 -2164
rect 10044 -2224 10528 -2164
rect 10594 -2224 10600 -2164
rect 10660 -2224 10666 -2164
rect 10044 -2336 10104 -2224
rect 10468 -2336 10528 -2224
rect -66 -2384 10708 -2336
rect -66 -2494 -4 -2384
rect 10652 -2494 10708 -2384
rect -66 -2550 10708 -2494
rect -328 -2916 -216 -2762
rect 384 -2916 394 -2616
rect 10306 -2916 10316 -2616
rect 10916 -2762 10922 -788
rect 11022 -2762 11028 122
rect 10916 -2916 11028 -2762
rect -328 -2922 11028 -2916
rect -328 -3022 -222 -2922
rect 10922 -3022 11028 -2922
rect -328 -3028 11028 -3022
<< via1 >>
rect -216 1996 384 2296
rect 10316 1996 10916 2296
rect 3514 1758 7278 1910
rect 5308 1556 5368 1616
rect 4152 892 4212 952
rect 4280 782 4340 842
rect 4668 892 4728 952
rect 4794 780 4854 840
rect 6346 1434 6406 1494
rect 5700 778 5760 838
rect 6864 776 6924 836
rect 3052 464 3112 524
rect 5700 464 5760 524
rect 8088 464 8148 524
rect 1494 170 1554 230
rect 2530 170 2590 230
rect 980 54 1040 114
rect 1370 -56 1430 4
rect 2012 54 2072 114
rect 1624 -56 1684 4
rect 1110 -786 1170 -726
rect 32 -896 92 -836
rect 2396 -56 2456 4
rect 3048 54 3108 114
rect 2658 -56 2718 4
rect 1886 -786 1946 -726
rect 2140 -786 2200 -726
rect 4790 176 4850 236
rect 5826 176 5886 236
rect 4276 60 4336 120
rect 2918 -786 2978 -726
rect 4666 -50 4726 10
rect 5308 60 5368 120
rect 4920 -50 4980 10
rect 1240 -896 1300 -836
rect 1752 -896 1812 -836
rect 2272 -896 2332 -836
rect 2788 -896 2848 -836
rect 4406 -780 4466 -720
rect 2918 -1018 2978 -958
rect 1030 -1142 1090 -1082
rect 1032 -1686 1092 -1626
rect 4536 -890 4596 -830
rect 5692 -50 5752 10
rect 6344 60 6404 120
rect 5954 -50 6014 10
rect 5182 -780 5242 -720
rect 5436 -780 5496 -720
rect 8086 170 8146 230
rect 9122 170 9182 230
rect 7572 54 7632 114
rect 6214 -780 6274 -720
rect 7962 -56 8022 4
rect 8604 54 8664 114
rect 8216 -56 8276 4
rect 5048 -890 5108 -830
rect 5568 -890 5628 -830
rect 6084 -890 6144 -830
rect 4798 -1018 4858 -958
rect 4464 -1142 4524 -1082
rect 2314 -1682 2374 -1626
rect 2748 -1686 2808 -1626
rect 3178 -1682 3238 -1626
rect 32 -2230 92 -2170
rect 7702 -786 7762 -726
rect 8988 -56 9048 4
rect 9640 54 9700 114
rect 9250 -56 9310 4
rect 8478 -786 8538 -726
rect 8732 -786 8792 -726
rect 9510 -786 9570 -726
rect 7832 -896 7892 -836
rect 8344 -896 8404 -836
rect 8864 -896 8924 -836
rect 9380 -896 9440 -836
rect 9614 -1026 9674 -966
rect 4038 -1682 4098 -1626
rect 4468 -1686 4528 -1626
rect 6184 -1686 6244 -1626
rect 6610 -1682 6670 -1626
rect 10600 -896 10660 -836
rect 7468 -1682 7528 -1626
rect 7896 -1686 7956 -1626
rect 8322 -1682 8382 -1626
rect 6180 -2230 6240 -2170
rect 9188 -1686 9248 -1626
rect 9612 -2224 9672 -2164
rect 10600 -2224 10660 -2164
rect -4 -2494 10652 -2384
rect -216 -2916 384 -2616
rect 10316 -2916 10916 -2616
<< metal2 >>
rect -216 2296 384 2306
rect -216 1986 384 1996
rect 10316 2296 10916 2306
rect 10316 1986 10916 1996
rect 3466 1910 7322 1950
rect 3466 1758 3514 1910
rect 7278 1758 7322 1910
rect 3466 1720 7322 1758
rect 5308 1616 5368 1622
rect 602 1556 5308 1616
rect 602 168 662 1556
rect 5308 1550 5368 1556
rect 6346 1494 6406 1500
rect 2532 1434 6346 1494
rect 2532 236 2592 1434
rect 6346 1428 6406 1434
rect 4152 952 4212 958
rect 4668 952 4728 958
rect 4212 892 4668 952
rect 4728 892 10792 952
rect 4152 886 4212 892
rect 4668 886 4728 892
rect 4274 782 4280 842
rect 4340 782 4346 842
rect 3046 464 3052 524
rect 3112 464 3118 524
rect -84 108 662 168
rect 1494 230 1554 236
rect 2530 230 2592 236
rect 1554 170 2530 230
rect 2590 170 2592 230
rect 1494 164 1554 170
rect 2530 164 2590 170
rect 3052 120 3112 464
rect 4280 126 4340 782
rect 4788 780 4794 840
rect 4854 780 4860 840
rect 4794 242 4854 780
rect 5694 778 5700 838
rect 5760 778 5766 838
rect 6864 836 6924 842
rect 5700 524 5760 778
rect 6924 776 7632 836
rect 6864 770 6924 776
rect 5694 464 5700 524
rect 5760 464 5766 524
rect 4790 236 4854 242
rect 5826 236 5886 242
rect 4850 176 5826 236
rect 4790 170 4850 176
rect 5826 170 5886 176
rect 980 114 1040 120
rect 2012 114 2072 120
rect 3048 114 3112 120
rect -84 -1626 -24 108
rect 1040 54 2012 114
rect 2072 54 3048 114
rect 3108 54 3112 114
rect 4276 120 4340 126
rect 5308 120 5368 126
rect 6344 120 6404 126
rect 4336 60 5308 120
rect 5368 60 6344 120
rect 6404 60 7262 120
rect 4276 54 4336 60
rect 5308 54 5368 60
rect 6344 54 6404 60
rect 980 48 1040 54
rect 2012 48 2072 54
rect 3048 48 3108 54
rect 4666 10 4726 16
rect 4920 10 4980 16
rect 5692 10 5752 16
rect 5954 10 6014 16
rect 1370 4 1430 10
rect 1624 4 1684 10
rect 2396 4 2456 10
rect 2658 4 2718 10
rect 1430 -56 1624 4
rect 1684 -56 2396 4
rect 2456 -56 2658 4
rect 2718 -56 3716 4
rect 4726 -50 4920 10
rect 4980 -50 5692 10
rect 5752 -50 5954 10
rect 4666 -56 4726 -50
rect 4920 -56 4980 -50
rect 5692 -56 5752 -50
rect 5954 -56 6014 -50
rect 7202 4 7262 60
rect 7572 114 7632 776
rect 8082 464 8088 524
rect 8148 464 8154 524
rect 8088 236 8148 464
rect 8086 230 8148 236
rect 9122 230 9182 236
rect 8146 170 9122 230
rect 8086 164 8146 170
rect 9122 164 9182 170
rect 8604 114 8664 120
rect 9640 114 9700 120
rect 7632 54 8604 114
rect 8664 54 9640 114
rect 7572 48 7632 54
rect 8604 48 8664 54
rect 9640 48 9700 54
rect 7962 4 8022 10
rect 8216 4 8276 10
rect 8988 4 9048 10
rect 9250 4 9310 10
rect 7202 -56 7962 4
rect 8022 -56 8216 4
rect 8276 -56 8988 4
rect 9048 -56 9250 4
rect 1370 -62 1430 -56
rect 1624 -62 1684 -56
rect 2396 -62 2456 -56
rect 2658 -62 2718 -56
rect 1110 -726 1170 -720
rect 1886 -726 1946 -720
rect 2140 -726 2200 -720
rect 2918 -726 2978 -720
rect 1170 -786 1886 -726
rect 1946 -786 2140 -726
rect 2200 -786 2918 -726
rect 1110 -792 1170 -786
rect 1886 -792 1946 -786
rect 2140 -792 2200 -786
rect 2918 -792 2978 -786
rect 32 -836 92 -830
rect 1752 -836 1812 -830
rect 2272 -836 2332 -830
rect 2788 -836 2848 -830
rect 92 -896 1240 -836
rect 1300 -896 1752 -836
rect 1812 -896 2272 -836
rect 2332 -896 2788 -836
rect 3656 -838 3716 -56
rect 7962 -62 8022 -56
rect 8216 -62 8276 -56
rect 8988 -62 9048 -56
rect 9250 -62 9310 -56
rect 4406 -720 4466 -714
rect 5182 -720 5242 -714
rect 5436 -720 5496 -714
rect 6214 -720 6274 -714
rect 4466 -780 5182 -720
rect 5242 -780 5436 -720
rect 5496 -780 6214 -720
rect 4406 -786 4466 -780
rect 5182 -786 5242 -780
rect 5436 -786 5496 -780
rect 6214 -786 6274 -780
rect 7702 -726 7762 -720
rect 8478 -726 8538 -720
rect 8732 -726 8792 -720
rect 9510 -726 9570 -720
rect 7762 -786 8478 -726
rect 8538 -786 8732 -726
rect 8792 -786 9510 -726
rect 7702 -792 7764 -786
rect 8478 -792 8538 -786
rect 8732 -792 8792 -786
rect 9510 -792 9570 -786
rect 5048 -830 5108 -824
rect 5568 -830 5628 -824
rect 6084 -830 6144 -824
rect 32 -902 92 -896
rect 1752 -902 1812 -896
rect 2272 -902 2332 -896
rect 2788 -902 2848 -896
rect 3647 -898 3656 -838
rect 3716 -898 3725 -838
rect 4530 -890 4536 -830
rect 4596 -890 5048 -830
rect 5108 -890 5568 -830
rect 5628 -890 6084 -830
rect 7704 -840 7764 -792
rect 7832 -836 7892 -830
rect 8344 -836 8404 -830
rect 8864 -836 8924 -830
rect 9380 -836 9440 -830
rect 10600 -836 10660 -830
rect 5048 -896 5108 -890
rect 5568 -896 5628 -890
rect 6084 -896 6144 -890
rect 7697 -896 7706 -840
rect 7762 -896 7771 -840
rect 7892 -896 8344 -836
rect 8404 -896 8864 -836
rect 8924 -896 9380 -836
rect 9440 -896 10600 -836
rect 7704 -898 7764 -896
rect 7832 -902 7892 -896
rect 8344 -902 8404 -896
rect 8864 -902 8924 -896
rect 9380 -902 9440 -896
rect 10600 -902 10660 -896
rect 2918 -958 2978 -952
rect 4798 -958 4858 -952
rect 2978 -1018 4798 -958
rect 2918 -1024 2978 -1018
rect 4798 -1024 4858 -1018
rect 9614 -966 9674 -960
rect 10732 -966 10792 892
rect 9674 -1026 10792 -966
rect 9614 -1032 9674 -1026
rect 1030 -1082 1090 -1076
rect 4464 -1082 4524 -1076
rect 1090 -1142 4464 -1082
rect 1030 -1148 1090 -1142
rect 4464 -1148 4524 -1142
rect 1032 -1626 1092 -1620
rect -84 -1686 1032 -1626
rect 1032 -1692 1092 -1686
rect 2314 -1626 2374 -1620
rect 2748 -1626 2808 -1620
rect 4468 -1626 4528 -1620
rect 6184 -1626 6244 -1620
rect 6610 -1626 6670 -1620
rect 7896 -1626 7956 -1620
rect 2374 -1682 2748 -1626
rect 2314 -1686 2748 -1682
rect 2808 -1682 3178 -1626
rect 3238 -1682 4038 -1626
rect 4098 -1682 4468 -1626
rect 2808 -1686 4468 -1682
rect 4528 -1686 6184 -1626
rect 6244 -1682 6610 -1626
rect 6670 -1682 7468 -1626
rect 7528 -1682 7896 -1626
rect 6244 -1686 7896 -1682
rect 7956 -1682 8322 -1626
rect 8382 -1682 9188 -1626
rect 7956 -1686 9188 -1682
rect 9248 -1686 9254 -1626
rect 2314 -1692 2374 -1686
rect 2748 -1692 2808 -1686
rect 4468 -1692 4528 -1686
rect 6184 -1692 6244 -1686
rect 6610 -1692 6670 -1686
rect 7896 -1692 7956 -1686
rect 9612 -2164 9672 -2158
rect 10600 -2164 10660 -2158
rect 32 -2170 92 -2164
rect 6180 -2170 6240 -2164
rect 92 -2230 6180 -2170
rect 9672 -2224 10600 -2164
rect 9612 -2230 9672 -2224
rect 10600 -2230 10660 -2224
rect 32 -2236 92 -2230
rect 6180 -2236 6240 -2230
rect -66 -2384 10708 -2336
rect -66 -2494 -4 -2384
rect 10652 -2494 10708 -2384
rect -66 -2550 10708 -2494
rect -216 -2616 384 -2606
rect -216 -2926 384 -2916
rect 10316 -2616 10916 -2606
rect 10316 -2926 10916 -2916
<< via2 >>
rect -216 1996 384 2296
rect 10316 1996 10916 2296
rect 3514 1758 7278 1910
rect 3656 -898 3716 -838
rect 7706 -896 7762 -840
rect -4 -2494 10652 -2384
rect -216 -2916 384 -2616
rect 10316 -2916 10916 -2616
<< metal3 >>
rect -226 2296 394 2301
rect -226 1996 -216 2296
rect 384 1996 394 2296
rect -226 1991 394 1996
rect 10306 2296 10926 2301
rect 10306 1996 10316 2296
rect 10916 1996 10926 2296
rect 10306 1991 10926 1996
rect 3466 1910 7322 1950
rect 3466 1758 3514 1910
rect 7278 1758 7322 1910
rect 3466 1720 7322 1758
rect 3628 -838 7786 -820
rect 3628 -898 3656 -838
rect 3716 -840 7786 -838
rect 3716 -896 7706 -840
rect 7762 -896 7786 -840
rect 3716 -898 7786 -896
rect 3628 -920 7786 -898
rect -66 -2384 10708 -2336
rect -66 -2494 -4 -2384
rect 10652 -2494 10708 -2384
rect -66 -2550 10708 -2494
rect -226 -2616 394 -2611
rect -226 -2916 -216 -2616
rect 384 -2916 394 -2616
rect -226 -2921 394 -2916
rect 10306 -2616 10926 -2611
rect 10306 -2916 10316 -2616
rect 10916 -2916 10926 -2616
rect 10306 -2921 10926 -2916
<< via3 >>
rect -216 1996 384 2296
rect 10316 1996 10916 2296
rect 3514 1758 7278 1910
rect -4 -2494 10652 -2384
rect -216 -2916 384 -2616
rect 10316 -2916 10916 -2616
<< metal4 >>
rect -400 2296 11100 2480
rect -400 1996 -216 2296
rect 384 1996 10316 2296
rect 10916 1996 11100 2296
rect -400 1910 11100 1996
rect -400 1758 3514 1910
rect 7278 1758 11100 1910
rect -400 1680 11100 1758
rect -400 -2384 11100 -2300
rect -400 -2494 -4 -2384
rect 10652 -2494 11100 -2384
rect -400 -2616 11100 -2494
rect -400 -2916 -216 -2616
rect 384 -2916 10316 -2616
rect 10916 -2916 11100 -2616
rect -400 -3100 11100 -2916
<< labels >>
flabel metal1 1044 -1164 1062 -1152 1 FreeSans 480 0 0 0 vtail_diff
flabel metal1 9634 -1132 9650 -1116 1 FreeSans 480 0 0 0 vbiasp
flabel metal1 9628 -2132 9644 -2122 1 FreeSans 480 0 0 0 vcmn_tail2
flabel metal1 6202 -2146 6214 -2134 1 FreeSans 480 0 0 0 vcmn_tail1
flabel metal1 1262 -1662 1270 -1654 1 FreeSans 480 0 0 0 vcmc
flabel metal2 6878 -1662 6892 -1652 1 FreeSans 480 0 0 0 ibiasn
port 6 n
flabel metal2 8640 -872 8650 -858 1 FreeSans 480 0 0 0 vcmn_tail2
flabel metal2 8428 -30 8440 -14 1 FreeSans 480 0 0 0 vom
port 5 n
flabel metal2 8082 -768 8104 -750 1 FreeSans 480 0 0 0 vocm
port 3 n
flabel metal2 7816 84 7828 94 1 FreeSans 480 0 0 0 vcmcn2
flabel metal2 8638 196 8648 208 1 FreeSans 480 0 0 0 vcmcn
flabel metal2 4368 918 4374 930 1 FreeSans 480 0 0 0 vbiasp
flabel metal2 5334 -876 5352 -860 1 FreeSans 480 0 0 0 vtail_diff
flabel metal2 5154 -28 5172 -12 1 FreeSans 480 0 0 0 vim
port 2 n
flabel metal2 4486 84 4506 96 1 FreeSans 480 0 0 0 vom
flabel metal2 5310 198 5330 214 1 FreeSans 480 0 0 0 vop
port 4 n
flabel metal2 2032 190 2050 210 1 FreeSans 480 0 0 0 vcmcn1
flabel metal2 1136 72 1156 86 1 FreeSans 480 0 0 0 vcmcn
flabel metal2 1856 -42 1878 -30 1 FreeSans 480 0 0 0 vocm
flabel metal2 1492 -760 1510 -748 1 FreeSans 480 0 0 0 vop
flabel metal2 2030 -874 2050 -858 1 FreeSans 480 0 0 0 vcmn_tail1
flabel metal2 4684 -754 4692 -748 1 FreeSans 480 0 0 0 vip
port 1 n
flabel metal1 5328 1322 5346 1338 1 FreeSans 480 0 0 0 vcmc
flabel metal2 4306 554 4312 558 1 FreeSans 480 0 0 0 vom
flabel metal2 4818 552 4824 558 1 FreeSans 480 0 0 0 vop
flabel metal4 -66 2456 -54 2470 1 FreeSans 480 0 0 0 VDD
port 7 n power bidirectional
flabel metal4 172 -3088 186 -3074 1 FreeSans 480 0 0 0 VSS
port 8 n ground bidirectional
<< end >>
