magic
tech sky130A
magscale 1 2
timestamp 1623661481
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 28 -17 62 17
<< locali >>
rect 17 299 94 491
rect 17 165 52 299
rect 297 265 362 425
rect 201 215 251 265
rect 201 199 235 215
rect 293 199 362 265
rect 396 199 451 332
rect 488 199 559 332
rect 664 199 719 265
rect 17 51 119 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 137 367 195 527
rect 229 459 502 493
rect 229 333 263 459
rect 128 299 263 333
rect 128 265 162 299
rect 436 417 502 459
rect 436 367 627 417
rect 89 215 162 265
rect 89 199 127 215
rect 593 165 627 367
rect 661 299 719 527
rect 228 131 508 165
rect 153 17 187 129
rect 228 51 294 131
rect 329 17 395 97
rect 442 93 508 131
rect 542 127 627 165
rect 661 93 719 147
rect 442 51 719 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 201 215 251 265 6 A1
port 1 nsew signal input
rlabel locali s 201 199 235 215 6 A1
port 1 nsew signal input
rlabel locali s 297 265 362 425 6 A2
port 2 nsew signal input
rlabel locali s 293 199 362 265 6 A2
port 2 nsew signal input
rlabel locali s 396 199 451 332 6 A3
port 3 nsew signal input
rlabel locali s 664 199 719 265 6 B1
port 4 nsew signal input
rlabel locali s 488 199 559 332 6 B2
port 5 nsew signal input
rlabel locali s 17 299 94 491 6 X
port 6 nsew signal output
rlabel locali s 17 165 52 299 6 X
port 6 nsew signal output
rlabel locali s 17 51 119 165 6 X
port 6 nsew signal output
rlabel metal1 s 0 -48 736 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel pwell s 28 -17 62 17 8 VNB
port 8 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 10 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
