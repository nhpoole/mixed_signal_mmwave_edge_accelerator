../../0-lvs_setup/outputs/user_analog_project_wrapper.spice