magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -2415 -1560 2415 1560
<< nwell >>
rect -1155 -300 1155 300
<< pmos >>
rect -1061 -200 -901 200
rect -843 -200 -683 200
rect -625 -200 -465 200
rect -407 -200 -247 200
rect -189 -200 -29 200
rect 29 -200 189 200
rect 247 -200 407 200
rect 465 -200 625 200
rect 683 -200 843 200
rect 901 -200 1061 200
<< pdiff >>
rect -1119 187 -1061 200
rect -1119 153 -1107 187
rect -1073 153 -1061 187
rect -1119 119 -1061 153
rect -1119 85 -1107 119
rect -1073 85 -1061 119
rect -1119 51 -1061 85
rect -1119 17 -1107 51
rect -1073 17 -1061 51
rect -1119 -17 -1061 17
rect -1119 -51 -1107 -17
rect -1073 -51 -1061 -17
rect -1119 -85 -1061 -51
rect -1119 -119 -1107 -85
rect -1073 -119 -1061 -85
rect -1119 -153 -1061 -119
rect -1119 -187 -1107 -153
rect -1073 -187 -1061 -153
rect -1119 -200 -1061 -187
rect -901 187 -843 200
rect -901 153 -889 187
rect -855 153 -843 187
rect -901 119 -843 153
rect -901 85 -889 119
rect -855 85 -843 119
rect -901 51 -843 85
rect -901 17 -889 51
rect -855 17 -843 51
rect -901 -17 -843 17
rect -901 -51 -889 -17
rect -855 -51 -843 -17
rect -901 -85 -843 -51
rect -901 -119 -889 -85
rect -855 -119 -843 -85
rect -901 -153 -843 -119
rect -901 -187 -889 -153
rect -855 -187 -843 -153
rect -901 -200 -843 -187
rect -683 187 -625 200
rect -683 153 -671 187
rect -637 153 -625 187
rect -683 119 -625 153
rect -683 85 -671 119
rect -637 85 -625 119
rect -683 51 -625 85
rect -683 17 -671 51
rect -637 17 -625 51
rect -683 -17 -625 17
rect -683 -51 -671 -17
rect -637 -51 -625 -17
rect -683 -85 -625 -51
rect -683 -119 -671 -85
rect -637 -119 -625 -85
rect -683 -153 -625 -119
rect -683 -187 -671 -153
rect -637 -187 -625 -153
rect -683 -200 -625 -187
rect -465 187 -407 200
rect -465 153 -453 187
rect -419 153 -407 187
rect -465 119 -407 153
rect -465 85 -453 119
rect -419 85 -407 119
rect -465 51 -407 85
rect -465 17 -453 51
rect -419 17 -407 51
rect -465 -17 -407 17
rect -465 -51 -453 -17
rect -419 -51 -407 -17
rect -465 -85 -407 -51
rect -465 -119 -453 -85
rect -419 -119 -407 -85
rect -465 -153 -407 -119
rect -465 -187 -453 -153
rect -419 -187 -407 -153
rect -465 -200 -407 -187
rect -247 187 -189 200
rect -247 153 -235 187
rect -201 153 -189 187
rect -247 119 -189 153
rect -247 85 -235 119
rect -201 85 -189 119
rect -247 51 -189 85
rect -247 17 -235 51
rect -201 17 -189 51
rect -247 -17 -189 17
rect -247 -51 -235 -17
rect -201 -51 -189 -17
rect -247 -85 -189 -51
rect -247 -119 -235 -85
rect -201 -119 -189 -85
rect -247 -153 -189 -119
rect -247 -187 -235 -153
rect -201 -187 -189 -153
rect -247 -200 -189 -187
rect -29 187 29 200
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -200 29 -187
rect 189 187 247 200
rect 189 153 201 187
rect 235 153 247 187
rect 189 119 247 153
rect 189 85 201 119
rect 235 85 247 119
rect 189 51 247 85
rect 189 17 201 51
rect 235 17 247 51
rect 189 -17 247 17
rect 189 -51 201 -17
rect 235 -51 247 -17
rect 189 -85 247 -51
rect 189 -119 201 -85
rect 235 -119 247 -85
rect 189 -153 247 -119
rect 189 -187 201 -153
rect 235 -187 247 -153
rect 189 -200 247 -187
rect 407 187 465 200
rect 407 153 419 187
rect 453 153 465 187
rect 407 119 465 153
rect 407 85 419 119
rect 453 85 465 119
rect 407 51 465 85
rect 407 17 419 51
rect 453 17 465 51
rect 407 -17 465 17
rect 407 -51 419 -17
rect 453 -51 465 -17
rect 407 -85 465 -51
rect 407 -119 419 -85
rect 453 -119 465 -85
rect 407 -153 465 -119
rect 407 -187 419 -153
rect 453 -187 465 -153
rect 407 -200 465 -187
rect 625 187 683 200
rect 625 153 637 187
rect 671 153 683 187
rect 625 119 683 153
rect 625 85 637 119
rect 671 85 683 119
rect 625 51 683 85
rect 625 17 637 51
rect 671 17 683 51
rect 625 -17 683 17
rect 625 -51 637 -17
rect 671 -51 683 -17
rect 625 -85 683 -51
rect 625 -119 637 -85
rect 671 -119 683 -85
rect 625 -153 683 -119
rect 625 -187 637 -153
rect 671 -187 683 -153
rect 625 -200 683 -187
rect 843 187 901 200
rect 843 153 855 187
rect 889 153 901 187
rect 843 119 901 153
rect 843 85 855 119
rect 889 85 901 119
rect 843 51 901 85
rect 843 17 855 51
rect 889 17 901 51
rect 843 -17 901 17
rect 843 -51 855 -17
rect 889 -51 901 -17
rect 843 -85 901 -51
rect 843 -119 855 -85
rect 889 -119 901 -85
rect 843 -153 901 -119
rect 843 -187 855 -153
rect 889 -187 901 -153
rect 843 -200 901 -187
rect 1061 187 1119 200
rect 1061 153 1073 187
rect 1107 153 1119 187
rect 1061 119 1119 153
rect 1061 85 1073 119
rect 1107 85 1119 119
rect 1061 51 1119 85
rect 1061 17 1073 51
rect 1107 17 1119 51
rect 1061 -17 1119 17
rect 1061 -51 1073 -17
rect 1107 -51 1119 -17
rect 1061 -85 1119 -51
rect 1061 -119 1073 -85
rect 1107 -119 1119 -85
rect 1061 -153 1119 -119
rect 1061 -187 1073 -153
rect 1107 -187 1119 -153
rect 1061 -200 1119 -187
<< pdiffc >>
rect -1107 153 -1073 187
rect -1107 85 -1073 119
rect -1107 17 -1073 51
rect -1107 -51 -1073 -17
rect -1107 -119 -1073 -85
rect -1107 -187 -1073 -153
rect -889 153 -855 187
rect -889 85 -855 119
rect -889 17 -855 51
rect -889 -51 -855 -17
rect -889 -119 -855 -85
rect -889 -187 -855 -153
rect -671 153 -637 187
rect -671 85 -637 119
rect -671 17 -637 51
rect -671 -51 -637 -17
rect -671 -119 -637 -85
rect -671 -187 -637 -153
rect -453 153 -419 187
rect -453 85 -419 119
rect -453 17 -419 51
rect -453 -51 -419 -17
rect -453 -119 -419 -85
rect -453 -187 -419 -153
rect -235 153 -201 187
rect -235 85 -201 119
rect -235 17 -201 51
rect -235 -51 -201 -17
rect -235 -119 -201 -85
rect -235 -187 -201 -153
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect 201 153 235 187
rect 201 85 235 119
rect 201 17 235 51
rect 201 -51 235 -17
rect 201 -119 235 -85
rect 201 -187 235 -153
rect 419 153 453 187
rect 419 85 453 119
rect 419 17 453 51
rect 419 -51 453 -17
rect 419 -119 453 -85
rect 419 -187 453 -153
rect 637 153 671 187
rect 637 85 671 119
rect 637 17 671 51
rect 637 -51 671 -17
rect 637 -119 671 -85
rect 637 -187 671 -153
rect 855 153 889 187
rect 855 85 889 119
rect 855 17 889 51
rect 855 -51 889 -17
rect 855 -119 889 -85
rect 855 -187 889 -153
rect 1073 153 1107 187
rect 1073 85 1107 119
rect 1073 17 1107 51
rect 1073 -51 1107 -17
rect 1073 -119 1107 -85
rect 1073 -187 1107 -153
<< poly >>
rect -1035 281 -927 297
rect -1035 264 -998 281
rect -1061 247 -998 264
rect -964 264 -927 281
rect -817 281 -709 297
rect -817 264 -780 281
rect -964 247 -901 264
rect -1061 200 -901 247
rect -843 247 -780 264
rect -746 264 -709 281
rect -599 281 -491 297
rect -599 264 -562 281
rect -746 247 -683 264
rect -843 200 -683 247
rect -625 247 -562 264
rect -528 264 -491 281
rect -381 281 -273 297
rect -381 264 -344 281
rect -528 247 -465 264
rect -625 200 -465 247
rect -407 247 -344 264
rect -310 264 -273 281
rect -163 281 -55 297
rect -163 264 -126 281
rect -310 247 -247 264
rect -407 200 -247 247
rect -189 247 -126 264
rect -92 264 -55 281
rect 55 281 163 297
rect 55 264 92 281
rect -92 247 -29 264
rect -189 200 -29 247
rect 29 247 92 264
rect 126 264 163 281
rect 273 281 381 297
rect 273 264 310 281
rect 126 247 189 264
rect 29 200 189 247
rect 247 247 310 264
rect 344 264 381 281
rect 491 281 599 297
rect 491 264 528 281
rect 344 247 407 264
rect 247 200 407 247
rect 465 247 528 264
rect 562 264 599 281
rect 709 281 817 297
rect 709 264 746 281
rect 562 247 625 264
rect 465 200 625 247
rect 683 247 746 264
rect 780 264 817 281
rect 927 281 1035 297
rect 927 264 964 281
rect 780 247 843 264
rect 683 200 843 247
rect 901 247 964 264
rect 998 264 1035 281
rect 998 247 1061 264
rect 901 200 1061 247
rect -1061 -247 -901 -200
rect -1061 -264 -998 -247
rect -1035 -281 -998 -264
rect -964 -264 -901 -247
rect -843 -247 -683 -200
rect -843 -264 -780 -247
rect -964 -281 -927 -264
rect -1035 -297 -927 -281
rect -817 -281 -780 -264
rect -746 -264 -683 -247
rect -625 -247 -465 -200
rect -625 -264 -562 -247
rect -746 -281 -709 -264
rect -817 -297 -709 -281
rect -599 -281 -562 -264
rect -528 -264 -465 -247
rect -407 -247 -247 -200
rect -407 -264 -344 -247
rect -528 -281 -491 -264
rect -599 -297 -491 -281
rect -381 -281 -344 -264
rect -310 -264 -247 -247
rect -189 -247 -29 -200
rect -189 -264 -126 -247
rect -310 -281 -273 -264
rect -381 -297 -273 -281
rect -163 -281 -126 -264
rect -92 -264 -29 -247
rect 29 -247 189 -200
rect 29 -264 92 -247
rect -92 -281 -55 -264
rect -163 -297 -55 -281
rect 55 -281 92 -264
rect 126 -264 189 -247
rect 247 -247 407 -200
rect 247 -264 310 -247
rect 126 -281 163 -264
rect 55 -297 163 -281
rect 273 -281 310 -264
rect 344 -264 407 -247
rect 465 -247 625 -200
rect 465 -264 528 -247
rect 344 -281 381 -264
rect 273 -297 381 -281
rect 491 -281 528 -264
rect 562 -264 625 -247
rect 683 -247 843 -200
rect 683 -264 746 -247
rect 562 -281 599 -264
rect 491 -297 599 -281
rect 709 -281 746 -264
rect 780 -264 843 -247
rect 901 -247 1061 -200
rect 901 -264 964 -247
rect 780 -281 817 -264
rect 709 -297 817 -281
rect 927 -281 964 -264
rect 998 -264 1061 -247
rect 998 -281 1035 -264
rect 927 -297 1035 -281
<< polycont >>
rect -998 247 -964 281
rect -780 247 -746 281
rect -562 247 -528 281
rect -344 247 -310 281
rect -126 247 -92 281
rect 92 247 126 281
rect 310 247 344 281
rect 528 247 562 281
rect 746 247 780 281
rect 964 247 998 281
rect -998 -281 -964 -247
rect -780 -281 -746 -247
rect -562 -281 -528 -247
rect -344 -281 -310 -247
rect -126 -281 -92 -247
rect 92 -281 126 -247
rect 310 -281 344 -247
rect 528 -281 562 -247
rect 746 -281 780 -247
rect 964 -281 998 -247
<< locali >>
rect -1035 247 -998 281
rect -964 247 -927 281
rect -817 247 -780 281
rect -746 247 -709 281
rect -599 247 -562 281
rect -528 247 -491 281
rect -381 247 -344 281
rect -310 247 -273 281
rect -163 247 -126 281
rect -92 247 -55 281
rect 55 247 92 281
rect 126 247 163 281
rect 273 247 310 281
rect 344 247 381 281
rect 491 247 528 281
rect 562 247 599 281
rect 709 247 746 281
rect 780 247 817 281
rect 927 247 964 281
rect 998 247 1035 281
rect -1107 187 -1073 204
rect -1107 119 -1073 127
rect -1107 51 -1073 55
rect -1107 -55 -1073 -51
rect -1107 -127 -1073 -119
rect -1107 -204 -1073 -187
rect -889 187 -855 204
rect -889 119 -855 127
rect -889 51 -855 55
rect -889 -55 -855 -51
rect -889 -127 -855 -119
rect -889 -204 -855 -187
rect -671 187 -637 204
rect -671 119 -637 127
rect -671 51 -637 55
rect -671 -55 -637 -51
rect -671 -127 -637 -119
rect -671 -204 -637 -187
rect -453 187 -419 204
rect -453 119 -419 127
rect -453 51 -419 55
rect -453 -55 -419 -51
rect -453 -127 -419 -119
rect -453 -204 -419 -187
rect -235 187 -201 204
rect -235 119 -201 127
rect -235 51 -201 55
rect -235 -55 -201 -51
rect -235 -127 -201 -119
rect -235 -204 -201 -187
rect -17 187 17 204
rect -17 119 17 127
rect -17 51 17 55
rect -17 -55 17 -51
rect -17 -127 17 -119
rect -17 -204 17 -187
rect 201 187 235 204
rect 201 119 235 127
rect 201 51 235 55
rect 201 -55 235 -51
rect 201 -127 235 -119
rect 201 -204 235 -187
rect 419 187 453 204
rect 419 119 453 127
rect 419 51 453 55
rect 419 -55 453 -51
rect 419 -127 453 -119
rect 419 -204 453 -187
rect 637 187 671 204
rect 637 119 671 127
rect 637 51 671 55
rect 637 -55 671 -51
rect 637 -127 671 -119
rect 637 -204 671 -187
rect 855 187 889 204
rect 855 119 889 127
rect 855 51 889 55
rect 855 -55 889 -51
rect 855 -127 889 -119
rect 855 -204 889 -187
rect 1073 187 1107 204
rect 1073 119 1107 127
rect 1073 51 1107 55
rect 1073 -55 1107 -51
rect 1073 -127 1107 -119
rect 1073 -204 1107 -187
rect -1035 -281 -998 -247
rect -964 -281 -927 -247
rect -817 -281 -780 -247
rect -746 -281 -709 -247
rect -599 -281 -562 -247
rect -528 -281 -491 -247
rect -381 -281 -344 -247
rect -310 -281 -273 -247
rect -163 -281 -126 -247
rect -92 -281 -55 -247
rect 55 -281 92 -247
rect 126 -281 163 -247
rect 273 -281 310 -247
rect 344 -281 381 -247
rect 491 -281 528 -247
rect 562 -281 599 -247
rect 709 -281 746 -247
rect 780 -281 817 -247
rect 927 -281 964 -247
rect 998 -281 1035 -247
<< viali >>
rect -998 247 -964 281
rect -780 247 -746 281
rect -562 247 -528 281
rect -344 247 -310 281
rect -126 247 -92 281
rect 92 247 126 281
rect 310 247 344 281
rect 528 247 562 281
rect 746 247 780 281
rect 964 247 998 281
rect -1107 153 -1073 161
rect -1107 127 -1073 153
rect -1107 85 -1073 89
rect -1107 55 -1073 85
rect -1107 -17 -1073 17
rect -1107 -85 -1073 -55
rect -1107 -89 -1073 -85
rect -1107 -153 -1073 -127
rect -1107 -161 -1073 -153
rect -889 153 -855 161
rect -889 127 -855 153
rect -889 85 -855 89
rect -889 55 -855 85
rect -889 -17 -855 17
rect -889 -85 -855 -55
rect -889 -89 -855 -85
rect -889 -153 -855 -127
rect -889 -161 -855 -153
rect -671 153 -637 161
rect -671 127 -637 153
rect -671 85 -637 89
rect -671 55 -637 85
rect -671 -17 -637 17
rect -671 -85 -637 -55
rect -671 -89 -637 -85
rect -671 -153 -637 -127
rect -671 -161 -637 -153
rect -453 153 -419 161
rect -453 127 -419 153
rect -453 85 -419 89
rect -453 55 -419 85
rect -453 -17 -419 17
rect -453 -85 -419 -55
rect -453 -89 -419 -85
rect -453 -153 -419 -127
rect -453 -161 -419 -153
rect -235 153 -201 161
rect -235 127 -201 153
rect -235 85 -201 89
rect -235 55 -201 85
rect -235 -17 -201 17
rect -235 -85 -201 -55
rect -235 -89 -201 -85
rect -235 -153 -201 -127
rect -235 -161 -201 -153
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect 201 153 235 161
rect 201 127 235 153
rect 201 85 235 89
rect 201 55 235 85
rect 201 -17 235 17
rect 201 -85 235 -55
rect 201 -89 235 -85
rect 201 -153 235 -127
rect 201 -161 235 -153
rect 419 153 453 161
rect 419 127 453 153
rect 419 85 453 89
rect 419 55 453 85
rect 419 -17 453 17
rect 419 -85 453 -55
rect 419 -89 453 -85
rect 419 -153 453 -127
rect 419 -161 453 -153
rect 637 153 671 161
rect 637 127 671 153
rect 637 85 671 89
rect 637 55 671 85
rect 637 -17 671 17
rect 637 -85 671 -55
rect 637 -89 671 -85
rect 637 -153 671 -127
rect 637 -161 671 -153
rect 855 153 889 161
rect 855 127 889 153
rect 855 85 889 89
rect 855 55 889 85
rect 855 -17 889 17
rect 855 -85 889 -55
rect 855 -89 889 -85
rect 855 -153 889 -127
rect 855 -161 889 -153
rect 1073 153 1107 161
rect 1073 127 1107 153
rect 1073 85 1107 89
rect 1073 55 1107 85
rect 1073 -17 1107 17
rect 1073 -85 1107 -55
rect 1073 -89 1107 -85
rect 1073 -153 1107 -127
rect 1073 -161 1107 -153
rect -998 -281 -964 -247
rect -780 -281 -746 -247
rect -562 -281 -528 -247
rect -344 -281 -310 -247
rect -126 -281 -92 -247
rect 92 -281 126 -247
rect 310 -281 344 -247
rect 528 -281 562 -247
rect 746 -281 780 -247
rect 964 -281 998 -247
<< metal1 >>
rect -1025 281 -937 287
rect -1025 247 -998 281
rect -964 247 -937 281
rect -1025 241 -937 247
rect -807 281 -719 287
rect -807 247 -780 281
rect -746 247 -719 281
rect -807 241 -719 247
rect -589 281 -501 287
rect -589 247 -562 281
rect -528 247 -501 281
rect -589 241 -501 247
rect -371 281 -283 287
rect -371 247 -344 281
rect -310 247 -283 281
rect -371 241 -283 247
rect -153 281 -65 287
rect -153 247 -126 281
rect -92 247 -65 281
rect -153 241 -65 247
rect 65 281 153 287
rect 65 247 92 281
rect 126 247 153 281
rect 65 241 153 247
rect 283 281 371 287
rect 283 247 310 281
rect 344 247 371 281
rect 283 241 371 247
rect 501 281 589 287
rect 501 247 528 281
rect 562 247 589 281
rect 501 241 589 247
rect 719 281 807 287
rect 719 247 746 281
rect 780 247 807 281
rect 719 241 807 247
rect 937 281 1025 287
rect 937 247 964 281
rect 998 247 1025 281
rect 937 241 1025 247
rect -1113 161 -1067 200
rect -1113 127 -1107 161
rect -1073 127 -1067 161
rect -1113 89 -1067 127
rect -1113 55 -1107 89
rect -1073 55 -1067 89
rect -1113 17 -1067 55
rect -1113 -17 -1107 17
rect -1073 -17 -1067 17
rect -1113 -55 -1067 -17
rect -1113 -89 -1107 -55
rect -1073 -89 -1067 -55
rect -1113 -127 -1067 -89
rect -1113 -161 -1107 -127
rect -1073 -161 -1067 -127
rect -1113 -200 -1067 -161
rect -895 161 -849 200
rect -895 127 -889 161
rect -855 127 -849 161
rect -895 89 -849 127
rect -895 55 -889 89
rect -855 55 -849 89
rect -895 17 -849 55
rect -895 -17 -889 17
rect -855 -17 -849 17
rect -895 -55 -849 -17
rect -895 -89 -889 -55
rect -855 -89 -849 -55
rect -895 -127 -849 -89
rect -895 -161 -889 -127
rect -855 -161 -849 -127
rect -895 -200 -849 -161
rect -677 161 -631 200
rect -677 127 -671 161
rect -637 127 -631 161
rect -677 89 -631 127
rect -677 55 -671 89
rect -637 55 -631 89
rect -677 17 -631 55
rect -677 -17 -671 17
rect -637 -17 -631 17
rect -677 -55 -631 -17
rect -677 -89 -671 -55
rect -637 -89 -631 -55
rect -677 -127 -631 -89
rect -677 -161 -671 -127
rect -637 -161 -631 -127
rect -677 -200 -631 -161
rect -459 161 -413 200
rect -459 127 -453 161
rect -419 127 -413 161
rect -459 89 -413 127
rect -459 55 -453 89
rect -419 55 -413 89
rect -459 17 -413 55
rect -459 -17 -453 17
rect -419 -17 -413 17
rect -459 -55 -413 -17
rect -459 -89 -453 -55
rect -419 -89 -413 -55
rect -459 -127 -413 -89
rect -459 -161 -453 -127
rect -419 -161 -413 -127
rect -459 -200 -413 -161
rect -241 161 -195 200
rect -241 127 -235 161
rect -201 127 -195 161
rect -241 89 -195 127
rect -241 55 -235 89
rect -201 55 -195 89
rect -241 17 -195 55
rect -241 -17 -235 17
rect -201 -17 -195 17
rect -241 -55 -195 -17
rect -241 -89 -235 -55
rect -201 -89 -195 -55
rect -241 -127 -195 -89
rect -241 -161 -235 -127
rect -201 -161 -195 -127
rect -241 -200 -195 -161
rect -23 161 23 200
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -200 23 -161
rect 195 161 241 200
rect 195 127 201 161
rect 235 127 241 161
rect 195 89 241 127
rect 195 55 201 89
rect 235 55 241 89
rect 195 17 241 55
rect 195 -17 201 17
rect 235 -17 241 17
rect 195 -55 241 -17
rect 195 -89 201 -55
rect 235 -89 241 -55
rect 195 -127 241 -89
rect 195 -161 201 -127
rect 235 -161 241 -127
rect 195 -200 241 -161
rect 413 161 459 200
rect 413 127 419 161
rect 453 127 459 161
rect 413 89 459 127
rect 413 55 419 89
rect 453 55 459 89
rect 413 17 459 55
rect 413 -17 419 17
rect 453 -17 459 17
rect 413 -55 459 -17
rect 413 -89 419 -55
rect 453 -89 459 -55
rect 413 -127 459 -89
rect 413 -161 419 -127
rect 453 -161 459 -127
rect 413 -200 459 -161
rect 631 161 677 200
rect 631 127 637 161
rect 671 127 677 161
rect 631 89 677 127
rect 631 55 637 89
rect 671 55 677 89
rect 631 17 677 55
rect 631 -17 637 17
rect 671 -17 677 17
rect 631 -55 677 -17
rect 631 -89 637 -55
rect 671 -89 677 -55
rect 631 -127 677 -89
rect 631 -161 637 -127
rect 671 -161 677 -127
rect 631 -200 677 -161
rect 849 161 895 200
rect 849 127 855 161
rect 889 127 895 161
rect 849 89 895 127
rect 849 55 855 89
rect 889 55 895 89
rect 849 17 895 55
rect 849 -17 855 17
rect 889 -17 895 17
rect 849 -55 895 -17
rect 849 -89 855 -55
rect 889 -89 895 -55
rect 849 -127 895 -89
rect 849 -161 855 -127
rect 889 -161 895 -127
rect 849 -200 895 -161
rect 1067 161 1113 200
rect 1067 127 1073 161
rect 1107 127 1113 161
rect 1067 89 1113 127
rect 1067 55 1073 89
rect 1107 55 1113 89
rect 1067 17 1113 55
rect 1067 -17 1073 17
rect 1107 -17 1113 17
rect 1067 -55 1113 -17
rect 1067 -89 1073 -55
rect 1107 -89 1113 -55
rect 1067 -127 1113 -89
rect 1067 -161 1073 -127
rect 1107 -161 1113 -127
rect 1067 -200 1113 -161
rect -1025 -247 -937 -241
rect -1025 -281 -998 -247
rect -964 -281 -937 -247
rect -1025 -287 -937 -281
rect -807 -247 -719 -241
rect -807 -281 -780 -247
rect -746 -281 -719 -247
rect -807 -287 -719 -281
rect -589 -247 -501 -241
rect -589 -281 -562 -247
rect -528 -281 -501 -247
rect -589 -287 -501 -281
rect -371 -247 -283 -241
rect -371 -281 -344 -247
rect -310 -281 -283 -247
rect -371 -287 -283 -281
rect -153 -247 -65 -241
rect -153 -281 -126 -247
rect -92 -281 -65 -247
rect -153 -287 -65 -281
rect 65 -247 153 -241
rect 65 -281 92 -247
rect 126 -281 153 -247
rect 65 -287 153 -281
rect 283 -247 371 -241
rect 283 -281 310 -247
rect 344 -281 371 -247
rect 283 -287 371 -281
rect 501 -247 589 -241
rect 501 -281 528 -247
rect 562 -281 589 -247
rect 501 -287 589 -281
rect 719 -247 807 -241
rect 719 -281 746 -247
rect 780 -281 807 -247
rect 719 -287 807 -281
rect 937 -247 1025 -241
rect 937 -281 964 -247
rect 998 -281 1025 -247
rect 937 -287 1025 -281
<< end >>
