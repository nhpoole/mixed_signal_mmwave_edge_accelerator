magic
tech sky130A
timestamp 1626065694
<< checkpaint >>
rect -732 -654 732 654
<< metal2 >>
rect -102 14 102 24
rect -102 -14 -94 14
rect -66 -14 -54 14
rect -26 -14 -14 14
rect 14 -14 26 14
rect 54 -14 66 14
rect 94 -14 102 14
rect -102 -24 102 -14
<< via2 >>
rect -94 -14 -66 14
rect -54 -14 -26 14
rect -14 -14 14 14
rect 26 -14 54 14
rect 66 -14 94 14
<< metal3 >>
rect -102 14 102 24
rect -102 -14 -94 14
rect -66 -14 -54 14
rect -26 -14 -14 14
rect 14 -14 26 14
rect 54 -14 66 14
rect 94 -14 102 14
rect -102 -24 102 -14
<< end >>
