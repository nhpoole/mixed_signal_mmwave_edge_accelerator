magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -30495 -77163 59785 1272
<< nwell >>
rect 10260 -57542 12494 -56702
<< locali >>
rect 10342 -56772 10363 -56738
rect 10397 -56772 10435 -56738
rect 10469 -56772 10507 -56738
rect 10541 -56772 10562 -56738
rect 11834 -56772 11846 -56738
rect 11880 -56772 11918 -56738
rect 11952 -56772 11990 -56738
rect 12024 -56772 12036 -56738
rect 10294 -56853 10332 -56836
rect 10294 -56887 10296 -56853
rect 10330 -56887 10332 -56853
rect 10294 -56925 10332 -56887
rect 10294 -56959 10296 -56925
rect 10330 -56959 10332 -56925
rect 10294 -56997 10332 -56959
rect 10294 -57031 10296 -56997
rect 10330 -57031 10332 -56997
rect 10294 -57069 10332 -57031
rect 10294 -57103 10296 -57069
rect 10330 -57103 10332 -57069
rect 10294 -57141 10332 -57103
rect 10294 -57175 10296 -57141
rect 10330 -57175 10332 -57141
rect 10294 -57213 10332 -57175
rect 10294 -57247 10296 -57213
rect 10330 -57247 10332 -57213
rect 10294 -57285 10332 -57247
rect 10294 -57319 10296 -57285
rect 10330 -57319 10332 -57285
rect 10294 -57357 10332 -57319
rect 10294 -57391 10296 -57357
rect 10330 -57391 10332 -57357
rect 10294 -57408 10332 -57391
rect 12070 -56853 12106 -56834
rect 12070 -56887 12071 -56853
rect 12105 -56887 12106 -56853
rect 12070 -56925 12106 -56887
rect 12070 -56959 12071 -56925
rect 12105 -56959 12106 -56925
rect 12070 -56997 12106 -56959
rect 12070 -57031 12071 -56997
rect 12105 -57031 12106 -56997
rect 12070 -57069 12106 -57031
rect 12070 -57103 12071 -57069
rect 12105 -57103 12106 -57069
rect 12070 -57141 12106 -57103
rect 12070 -57175 12071 -57141
rect 12105 -57175 12106 -57141
rect 12070 -57213 12106 -57175
rect 12070 -57247 12071 -57213
rect 12105 -57247 12106 -57213
rect 12070 -57285 12106 -57247
rect 12070 -57319 12071 -57285
rect 12105 -57319 12106 -57285
rect 12070 -57357 12106 -57319
rect 12070 -57391 12071 -57357
rect 12105 -57391 12106 -57357
rect 12070 -57410 12106 -57391
rect 10342 -57506 10363 -57472
rect 10397 -57506 10435 -57472
rect 10469 -57506 10507 -57472
rect 10541 -57506 10562 -57472
rect 11834 -57504 11846 -57470
rect 11880 -57504 11918 -57470
rect 11952 -57504 11990 -57470
rect 12024 -57504 12036 -57470
rect 12238 -57545 12286 -57538
rect 12238 -57579 12245 -57545
rect 12279 -57579 12286 -57545
rect 12238 -57586 12286 -57579
rect 12342 -57545 12390 -57538
rect 12342 -57579 12349 -57545
rect 12383 -57579 12390 -57545
rect 12342 -57586 12390 -57579
rect 11838 -57670 12036 -57668
rect 10366 -57672 10574 -57670
rect 10366 -57706 10381 -57672
rect 10415 -57706 10453 -57672
rect 10487 -57706 10525 -57672
rect 10559 -57706 10574 -57672
rect 11838 -57704 11848 -57670
rect 11882 -57704 11920 -57670
rect 11954 -57704 11992 -57670
rect 12026 -57704 12036 -57670
rect 11838 -57706 12036 -57704
rect 10366 -57708 10574 -57706
rect 10294 -57785 10330 -57768
rect 10294 -57819 10295 -57785
rect 10329 -57819 10330 -57785
rect 10294 -57857 10330 -57819
rect 10294 -57891 10295 -57857
rect 10329 -57891 10330 -57857
rect 10294 -57929 10330 -57891
rect 10294 -57963 10295 -57929
rect 10329 -57963 10330 -57929
rect 10294 -58001 10330 -57963
rect 10294 -58035 10295 -58001
rect 10329 -58035 10330 -58001
rect 10294 -58073 10330 -58035
rect 10294 -58107 10295 -58073
rect 10329 -58107 10330 -58073
rect 10294 -58124 10330 -58107
rect 12070 -57785 12108 -57768
rect 12070 -57819 12072 -57785
rect 12106 -57819 12108 -57785
rect 12070 -57857 12108 -57819
rect 12070 -57891 12072 -57857
rect 12106 -57891 12108 -57857
rect 12070 -57929 12108 -57891
rect 12070 -57963 12072 -57929
rect 12106 -57963 12108 -57929
rect 12070 -58001 12108 -57963
rect 12070 -58035 12072 -58001
rect 12106 -58035 12108 -58001
rect 12070 -58073 12108 -58035
rect 12070 -58107 12072 -58073
rect 12106 -58107 12108 -58073
rect 12070 -58124 12108 -58107
rect 10364 -58185 10572 -58184
rect 10364 -58219 10379 -58185
rect 10413 -58219 10451 -58185
rect 10485 -58219 10523 -58185
rect 10557 -58219 10572 -58185
rect 10364 -58220 10572 -58219
rect 11836 -58187 12038 -58186
rect 11836 -58221 11848 -58187
rect 11882 -58221 11920 -58187
rect 11954 -58221 11992 -58187
rect 12026 -58221 12038 -58187
rect 11836 -58222 12038 -58221
<< viali >>
rect 10363 -56772 10397 -56738
rect 10435 -56772 10469 -56738
rect 10507 -56772 10541 -56738
rect 11846 -56772 11880 -56738
rect 11918 -56772 11952 -56738
rect 11990 -56772 12024 -56738
rect 10296 -56887 10330 -56853
rect 10296 -56959 10330 -56925
rect 10296 -57031 10330 -56997
rect 10296 -57103 10330 -57069
rect 10296 -57175 10330 -57141
rect 10296 -57247 10330 -57213
rect 10296 -57319 10330 -57285
rect 10296 -57391 10330 -57357
rect 12071 -56887 12105 -56853
rect 12071 -56959 12105 -56925
rect 12071 -57031 12105 -56997
rect 12071 -57103 12105 -57069
rect 12071 -57175 12105 -57141
rect 12071 -57247 12105 -57213
rect 12071 -57319 12105 -57285
rect 12071 -57391 12105 -57357
rect 10363 -57506 10397 -57472
rect 10435 -57506 10469 -57472
rect 10507 -57506 10541 -57472
rect 11846 -57504 11880 -57470
rect 11918 -57504 11952 -57470
rect 11990 -57504 12024 -57470
rect 12245 -57579 12279 -57545
rect 12349 -57579 12383 -57545
rect 10381 -57706 10415 -57672
rect 10453 -57706 10487 -57672
rect 10525 -57706 10559 -57672
rect 11848 -57704 11882 -57670
rect 11920 -57704 11954 -57670
rect 11992 -57704 12026 -57670
rect 10295 -57819 10329 -57785
rect 10295 -57891 10329 -57857
rect 10295 -57963 10329 -57929
rect 10295 -58035 10329 -58001
rect 10295 -58107 10329 -58073
rect 12072 -57819 12106 -57785
rect 12072 -57891 12106 -57857
rect 12072 -57963 12106 -57929
rect 12072 -58035 12106 -58001
rect 12072 -58107 12106 -58073
rect 10379 -58219 10413 -58185
rect 10451 -58219 10485 -58185
rect 10523 -58219 10557 -58185
rect 11848 -58221 11882 -58187
rect 11920 -58221 11954 -58187
rect 11992 -58221 12026 -58187
<< metal1 >>
rect -74 -48 106 12
rect 53108 -40021 53424 -40017
rect 53108 -40073 53118 -40021
rect 53170 -40073 53424 -40021
rect 53108 -40077 53424 -40073
rect 30132 -41244 30192 -41148
rect 30132 -41296 30136 -41244
rect 30188 -41296 30192 -41244
rect 30132 -41306 30192 -41296
rect 30132 -41826 30192 -41816
rect 30132 -41878 30136 -41826
rect 30188 -41878 30192 -41826
rect 30132 -41888 30192 -41878
rect 57134 -41984 57194 -41978
rect 57034 -41988 57194 -41984
rect 57034 -42040 57138 -41988
rect 57190 -42040 57194 -41988
rect 57034 -42044 57194 -42040
rect 57134 -42050 57194 -42044
rect 26980 -45108 27052 -45104
rect 26980 -45160 26990 -45108
rect 27042 -45160 27052 -45108
rect 26980 -45164 27052 -45160
rect 27774 -45108 27846 -45104
rect 27774 -45160 27784 -45108
rect 27836 -45160 27846 -45108
rect 27774 -45164 27846 -45160
rect 26980 -46864 27052 -46860
rect 26980 -46916 26990 -46864
rect 27042 -46916 27052 -46864
rect 26980 -46920 27052 -46916
rect 27774 -46864 27846 -46860
rect 27774 -46916 27784 -46864
rect 27836 -46916 27846 -46864
rect 27774 -46920 27846 -46916
rect 26980 -48378 27052 -48374
rect 26980 -48430 26990 -48378
rect 27042 -48430 27052 -48378
rect 26980 -48434 27052 -48430
rect 26976 -49620 27048 -49616
rect 26976 -49672 26986 -49620
rect 27038 -49672 27048 -49620
rect 26976 -49676 27048 -49672
rect 26980 -50856 27052 -50852
rect 26980 -50908 26990 -50856
rect 27042 -50908 27052 -50856
rect 26980 -50912 27052 -50908
rect 14762 -52972 14862 -52942
rect 14762 -53024 14786 -52972
rect 14838 -53024 14862 -52972
rect 27776 -52966 27848 -52962
rect 27776 -53018 27786 -52966
rect 27838 -53018 27848 -52966
rect 27776 -53022 27848 -53018
rect 14762 -53054 14862 -53024
rect 26374 -53568 26446 -53564
rect 26374 -53620 26384 -53568
rect 26436 -53620 26446 -53568
rect 26374 -53624 26446 -53620
rect 27774 -53568 27846 -53564
rect 27774 -53620 27784 -53568
rect 27836 -53620 27846 -53568
rect 27774 -53624 27846 -53620
rect 26380 -53734 26440 -53624
rect 14764 -53966 14864 -53936
rect 14764 -54018 14788 -53966
rect 14840 -54018 14864 -53966
rect 14764 -54048 14864 -54018
rect 14764 -54972 14864 -54942
rect 14764 -55024 14788 -54972
rect 14840 -55024 14864 -54972
rect 14764 -55054 14864 -55024
rect 27774 -55400 27846 -55396
rect 27774 -55452 27784 -55400
rect 27836 -55452 27846 -55400
rect 27774 -55456 27846 -55452
rect 10528 -56672 11876 -56612
rect 9350 -56724 9452 -56700
rect 9350 -56726 10454 -56724
rect 10528 -56726 10588 -56672
rect 9350 -56738 10588 -56726
rect 9350 -56743 10363 -56738
rect 9350 -56795 9378 -56743
rect 9430 -56772 10363 -56743
rect 10397 -56772 10435 -56738
rect 10469 -56772 10507 -56738
rect 10541 -56772 10588 -56738
rect 9430 -56784 10588 -56772
rect 9430 -56795 9452 -56784
rect 9350 -56807 9452 -56795
rect 9350 -56859 9378 -56807
rect 9430 -56859 9452 -56807
rect 9350 -56871 9452 -56859
rect 9350 -56923 9378 -56871
rect 9430 -56923 9452 -56871
rect 9350 -56935 9452 -56923
rect 9350 -56987 9378 -56935
rect 9430 -56987 9452 -56935
rect 9350 -56999 9452 -56987
rect 9350 -57051 9378 -56999
rect 9430 -57051 9452 -56999
rect 9350 -57063 9452 -57051
rect 9350 -57115 9378 -57063
rect 9430 -57094 9452 -57063
rect 10284 -56786 10588 -56784
rect 10284 -56853 10344 -56786
rect 10284 -56887 10296 -56853
rect 10330 -56887 10344 -56853
rect 10284 -56925 10344 -56887
rect 10284 -56959 10296 -56925
rect 10330 -56959 10344 -56925
rect 10284 -56997 10344 -56959
rect 10284 -57031 10296 -56997
rect 10330 -57031 10344 -56997
rect 10284 -57069 10344 -57031
rect 10284 -57094 10296 -57069
rect 9430 -57103 10296 -57094
rect 10330 -57094 10344 -57069
rect 10394 -57094 10454 -56786
rect 10528 -56877 10588 -56786
rect 10784 -56720 10844 -56719
rect 11560 -56720 11620 -56714
rect 10784 -56724 11620 -56720
rect 10784 -56776 11564 -56724
rect 11616 -56776 11620 -56724
rect 10784 -56780 11620 -56776
rect 10784 -56875 10844 -56780
rect 11042 -56877 11102 -56780
rect 11300 -56875 11360 -56780
rect 11560 -56875 11620 -56780
rect 11816 -56722 11876 -56672
rect 11816 -56738 12118 -56722
rect 11816 -56772 11846 -56738
rect 11880 -56772 11918 -56738
rect 11952 -56772 11990 -56738
rect 12024 -56772 12118 -56738
rect 11816 -56786 12118 -56772
rect 11816 -56877 11876 -56786
rect 10330 -57103 10454 -57094
rect 9430 -57115 10454 -57103
rect 9350 -57127 10454 -57115
rect 9350 -57179 9378 -57127
rect 9430 -57141 10454 -57127
rect 9430 -57154 10296 -57141
rect 9430 -57179 9452 -57154
rect 9350 -57191 9452 -57179
rect 9350 -57243 9378 -57191
rect 9430 -57243 9452 -57191
rect 9350 -57255 9452 -57243
rect 9350 -57307 9378 -57255
rect 9430 -57307 9452 -57255
rect 9350 -57319 9452 -57307
rect 9350 -57371 9378 -57319
rect 9430 -57371 9452 -57319
rect 9350 -57383 9452 -57371
rect 9350 -57435 9378 -57383
rect 9430 -57435 9452 -57383
rect 9350 -57447 9452 -57435
rect 9350 -57499 9378 -57447
rect 9430 -57458 9452 -57447
rect 10284 -57175 10296 -57154
rect 10330 -57154 10454 -57141
rect 11944 -57092 12004 -56786
rect 12058 -56853 12118 -56786
rect 12058 -56887 12071 -56853
rect 12105 -56887 12118 -56853
rect 12058 -56925 12118 -56887
rect 12058 -56959 12071 -56925
rect 12105 -56959 12118 -56925
rect 15194 -56954 15562 -56894
rect 17356 -56954 17566 -56894
rect 12058 -56997 12118 -56959
rect 12058 -57031 12071 -56997
rect 12105 -57031 12118 -56997
rect 12058 -57069 12118 -57031
rect 12058 -57092 12071 -57069
rect 11944 -57103 12071 -57092
rect 12105 -57103 12118 -57069
rect 11944 -57141 12118 -57103
rect 11944 -57152 12071 -57141
rect 10330 -57175 10344 -57154
rect 10284 -57213 10344 -57175
rect 10284 -57247 10296 -57213
rect 10330 -57247 10344 -57213
rect 10284 -57285 10344 -57247
rect 12058 -57175 12071 -57152
rect 12105 -57175 12118 -57141
rect 12058 -57210 12118 -57175
rect 12058 -57213 12184 -57210
rect 12058 -57247 12071 -57213
rect 12105 -57247 12184 -57213
rect 10284 -57319 10296 -57285
rect 10330 -57319 10344 -57285
rect 10284 -57357 10344 -57319
rect 10284 -57391 10296 -57357
rect 10330 -57391 10344 -57357
rect 10284 -57458 10344 -57391
rect 10396 -57458 10456 -57276
rect 10524 -57458 10584 -57370
rect 9430 -57472 10584 -57458
rect 9430 -57499 10363 -57472
rect 9350 -57506 10363 -57499
rect 10397 -57506 10435 -57472
rect 10469 -57506 10507 -57472
rect 10541 -57506 10584 -57472
rect 9350 -57518 10584 -57506
rect 9350 -57536 9452 -57518
rect 10654 -57635 10714 -57265
rect 10912 -57486 10972 -57290
rect 10906 -57490 10978 -57486
rect 10906 -57542 10916 -57490
rect 10968 -57542 10978 -57490
rect 10906 -57546 10978 -57542
rect 10648 -57639 10720 -57635
rect 10282 -57672 10586 -57660
rect 10282 -57706 10381 -57672
rect 10415 -57706 10453 -57672
rect 10487 -57706 10525 -57672
rect 10559 -57706 10586 -57672
rect 10648 -57691 10658 -57639
rect 10710 -57691 10720 -57639
rect 10648 -57695 10720 -57691
rect 10282 -57720 10586 -57706
rect 10282 -57785 10342 -57720
rect 10282 -57819 10295 -57785
rect 10329 -57819 10342 -57785
rect 10282 -57857 10342 -57819
rect 10282 -57891 10295 -57857
rect 10329 -57891 10342 -57857
rect 10282 -57929 10342 -57891
rect 10396 -57908 10456 -57720
rect 10526 -57808 10586 -57720
rect 10654 -57895 10714 -57695
rect 10912 -57828 10972 -57546
rect 11170 -57635 11230 -57267
rect 11430 -57486 11490 -57272
rect 11424 -57490 11496 -57486
rect 11424 -57542 11434 -57490
rect 11486 -57542 11496 -57490
rect 11424 -57546 11496 -57542
rect 11164 -57639 11236 -57635
rect 11164 -57691 11174 -57639
rect 11226 -57691 11236 -57639
rect 11164 -57695 11236 -57691
rect 10912 -57894 10974 -57828
rect 10282 -57963 10295 -57929
rect 10329 -57963 10342 -57929
rect 10282 -58001 10342 -57963
rect 10282 -58035 10295 -58001
rect 10329 -58035 10342 -58001
rect 10282 -58073 10342 -58035
rect 10282 -58107 10295 -58073
rect 10329 -58107 10342 -58073
rect 10282 -58173 10342 -58107
rect 10398 -58173 10458 -57995
rect 10914 -58074 10974 -57894
rect 11170 -58014 11230 -57695
rect 11430 -58074 11490 -57546
rect 11688 -57639 11748 -57267
rect 11812 -57458 11872 -57370
rect 11946 -57458 12006 -57280
rect 12058 -57285 12184 -57247
rect 12058 -57319 12071 -57285
rect 12105 -57306 12184 -57285
rect 12105 -57319 12118 -57306
rect 12058 -57357 12118 -57319
rect 12058 -57391 12071 -57357
rect 12105 -57391 12118 -57357
rect 12058 -57458 12118 -57391
rect 11812 -57470 12118 -57458
rect 11812 -57504 11846 -57470
rect 11880 -57504 11918 -57470
rect 11952 -57504 11990 -57470
rect 12024 -57504 12118 -57470
rect 11812 -57518 12118 -57504
rect 12176 -57532 12236 -57526
rect 12524 -57532 12584 -57526
rect 12176 -57536 12298 -57532
rect 12176 -57588 12180 -57536
rect 12232 -57545 12298 -57536
rect 12232 -57579 12245 -57545
rect 12279 -57579 12298 -57545
rect 12232 -57588 12298 -57579
rect 12176 -57592 12298 -57588
rect 12330 -57536 12584 -57532
rect 12330 -57545 12528 -57536
rect 12330 -57579 12349 -57545
rect 12383 -57579 12528 -57545
rect 12330 -57588 12528 -57579
rect 12580 -57588 12584 -57536
rect 12330 -57592 12584 -57588
rect 12176 -57598 12236 -57592
rect 12524 -57598 12584 -57592
rect 11688 -57691 11692 -57639
rect 11744 -57691 11748 -57639
rect 11688 -57897 11748 -57691
rect 11818 -57670 12120 -57658
rect 11818 -57704 11848 -57670
rect 11882 -57704 11920 -57670
rect 11954 -57704 11992 -57670
rect 12026 -57704 12120 -57670
rect 11818 -57718 12120 -57704
rect 11818 -57806 11878 -57718
rect 11946 -57904 12006 -57718
rect 12060 -57754 12120 -57718
rect 12060 -57785 12190 -57754
rect 12060 -57819 12072 -57785
rect 12106 -57819 12190 -57785
rect 12060 -57850 12190 -57819
rect 12436 -57850 13132 -57754
rect 12060 -57857 12120 -57850
rect 12060 -57891 12072 -57857
rect 12106 -57891 12120 -57857
rect 12060 -57929 12120 -57891
rect 12060 -57963 12072 -57929
rect 12106 -57963 12120 -57929
rect 12060 -58001 12120 -57963
rect 10908 -58078 10980 -58074
rect 10526 -58173 10586 -58084
rect 10282 -58185 10586 -58173
rect 10282 -58219 10379 -58185
rect 10413 -58219 10451 -58185
rect 10485 -58219 10523 -58185
rect 10557 -58219 10586 -58185
rect 10282 -58233 10586 -58219
rect 10282 -58390 10342 -58233
rect 10398 -58390 10458 -58233
rect 10526 -58390 10586 -58233
rect 10784 -58183 10844 -58083
rect 10908 -58130 10918 -58078
rect 10970 -58130 10980 -58078
rect 11424 -58078 11496 -58074
rect 10908 -58134 10980 -58130
rect 11044 -58183 11104 -58083
rect 11302 -58183 11362 -58085
rect 11424 -58130 11434 -58078
rect 11486 -58130 11496 -58078
rect 11424 -58134 11496 -58130
rect 11558 -58183 11618 -58085
rect 11816 -58173 11876 -58082
rect 11944 -58173 12004 -58001
rect 12060 -58035 12072 -58001
rect 12106 -58035 12120 -58001
rect 12060 -58073 12120 -58035
rect 12060 -58107 12072 -58073
rect 12106 -58107 12120 -58073
rect 12060 -58173 12120 -58107
rect 10784 -58187 11624 -58183
rect 10784 -58239 11562 -58187
rect 11614 -58239 11624 -58187
rect 10784 -58243 11624 -58239
rect 11816 -58187 12120 -58173
rect 11816 -58221 11848 -58187
rect 11882 -58221 11920 -58187
rect 11954 -58221 11992 -58187
rect 12026 -58221 12120 -58187
rect 11816 -58233 12120 -58221
rect 11816 -58390 11876 -58233
rect 11944 -58390 12004 -58233
rect 12060 -58390 12120 -58233
rect 10276 -58435 12130 -58390
rect 10276 -58487 10312 -58435
rect 10364 -58487 10376 -58435
rect 10428 -58487 10440 -58435
rect 10492 -58487 10504 -58435
rect 10556 -58487 10568 -58435
rect 10620 -58487 10632 -58435
rect 10684 -58487 10696 -58435
rect 10748 -58487 10760 -58435
rect 10812 -58487 10824 -58435
rect 10876 -58487 10888 -58435
rect 10940 -58487 10952 -58435
rect 11004 -58487 11016 -58435
rect 11068 -58487 11080 -58435
rect 11132 -58487 11144 -58435
rect 11196 -58487 11208 -58435
rect 11260 -58487 11272 -58435
rect 11324 -58487 11336 -58435
rect 11388 -58487 11400 -58435
rect 11452 -58487 11464 -58435
rect 11516 -58487 11528 -58435
rect 11580 -58487 11592 -58435
rect 11644 -58487 11656 -58435
rect 11708 -58487 11720 -58435
rect 11772 -58487 11784 -58435
rect 11836 -58487 11848 -58435
rect 11900 -58487 11912 -58435
rect 11964 -58487 11976 -58435
rect 12028 -58487 12040 -58435
rect 12092 -58487 12130 -58435
rect 10276 -58528 12130 -58487
rect -3252 -72336 -3180 -72332
rect -3252 -72388 -3242 -72336
rect -3190 -72388 -3180 -72336
rect -3252 -72392 -3180 -72388
rect -2708 -72404 -2648 -71934
rect -2452 -72384 -2392 -71934
rect -28374 -72640 -28084 -72580
rect -24360 -72640 -24032 -72580
rect -20376 -72640 -20040 -72580
rect -16390 -72640 -16040 -72580
rect -12428 -72640 -12040 -72580
rect -8402 -72640 -8076 -72580
rect -392 -72640 -52 -72580
rect 3606 -72640 3958 -72580
rect -27092 -74870 -27032 -74054
rect -23092 -74868 -23032 -74034
rect -19092 -74868 -19032 -74042
rect -15092 -74868 -15032 -74048
rect -27098 -74874 -27026 -74870
rect -27098 -74926 -27088 -74874
rect -27036 -74926 -27026 -74874
rect -27098 -74930 -27026 -74926
rect -23098 -74872 -23026 -74868
rect -23098 -74924 -23088 -74872
rect -23036 -74924 -23026 -74872
rect -23098 -74928 -23026 -74924
rect -19098 -74872 -19026 -74868
rect -19098 -74924 -19088 -74872
rect -19036 -74924 -19026 -74872
rect -19098 -74928 -19026 -74924
rect -15098 -74872 -15026 -74868
rect -11092 -74870 -11032 -74034
rect -7092 -74870 -7032 -74036
rect -3092 -74868 -3032 -74034
rect 908 -74868 968 -74028
rect 4908 -74866 4968 -74040
rect -15098 -74924 -15088 -74872
rect -15036 -74924 -15026 -74872
rect -15098 -74928 -15026 -74924
rect -11098 -74874 -11026 -74870
rect -11098 -74926 -11088 -74874
rect -11036 -74926 -11026 -74874
rect -11098 -74930 -11026 -74926
rect -7098 -74874 -7026 -74870
rect -7098 -74926 -7088 -74874
rect -7036 -74926 -7026 -74874
rect -7098 -74930 -7026 -74926
rect -3098 -74872 -3026 -74868
rect -3098 -74924 -3088 -74872
rect -3036 -74924 -3026 -74872
rect -3098 -74928 -3026 -74924
rect 902 -74872 974 -74868
rect 902 -74924 912 -74872
rect 964 -74924 974 -74872
rect 902 -74928 974 -74924
rect 4902 -74870 4974 -74866
rect 4902 -74922 4912 -74870
rect 4964 -74922 4974 -74870
rect 4902 -74926 4974 -74922
<< via1 >>
rect 53118 -40073 53170 -40021
rect 30136 -41296 30188 -41244
rect 30136 -41878 30188 -41826
rect 57138 -42040 57190 -41988
rect 26990 -45160 27042 -45108
rect 27784 -45160 27836 -45108
rect 26990 -46916 27042 -46864
rect 27784 -46916 27836 -46864
rect 26990 -48430 27042 -48378
rect 26986 -49672 27038 -49620
rect 26990 -50908 27042 -50856
rect 14786 -53024 14838 -52972
rect 27786 -53018 27838 -52966
rect 26384 -53620 26436 -53568
rect 27784 -53620 27836 -53568
rect 14788 -54018 14840 -53966
rect 14788 -55024 14840 -54972
rect 27784 -55452 27836 -55400
rect 9378 -56795 9430 -56743
rect 9378 -56859 9430 -56807
rect 9378 -56923 9430 -56871
rect 9378 -56987 9430 -56935
rect 9378 -57051 9430 -56999
rect 9378 -57115 9430 -57063
rect 11564 -56776 11616 -56724
rect 9378 -57179 9430 -57127
rect 9378 -57243 9430 -57191
rect 9378 -57307 9430 -57255
rect 9378 -57371 9430 -57319
rect 9378 -57435 9430 -57383
rect 9378 -57499 9430 -57447
rect 10916 -57542 10968 -57490
rect 10658 -57691 10710 -57639
rect 11434 -57542 11486 -57490
rect 11174 -57691 11226 -57639
rect 12180 -57588 12232 -57536
rect 12528 -57588 12580 -57536
rect 11692 -57691 11744 -57639
rect 10918 -58130 10970 -58078
rect 11434 -58130 11486 -58078
rect 11562 -58239 11614 -58187
rect 10312 -58487 10364 -58435
rect 10376 -58487 10428 -58435
rect 10440 -58487 10492 -58435
rect 10504 -58487 10556 -58435
rect 10568 -58487 10620 -58435
rect 10632 -58487 10684 -58435
rect 10696 -58487 10748 -58435
rect 10760 -58487 10812 -58435
rect 10824 -58487 10876 -58435
rect 10888 -58487 10940 -58435
rect 10952 -58487 11004 -58435
rect 11016 -58487 11068 -58435
rect 11080 -58487 11132 -58435
rect 11144 -58487 11196 -58435
rect 11208 -58487 11260 -58435
rect 11272 -58487 11324 -58435
rect 11336 -58487 11388 -58435
rect 11400 -58487 11452 -58435
rect 11464 -58487 11516 -58435
rect 11528 -58487 11580 -58435
rect 11592 -58487 11644 -58435
rect 11656 -58487 11708 -58435
rect 11720 -58487 11772 -58435
rect 11784 -58487 11836 -58435
rect 11848 -58487 11900 -58435
rect 11912 -58487 11964 -58435
rect 11976 -58487 12028 -58435
rect 12040 -58487 12092 -58435
rect -3242 -72388 -3190 -72336
rect -27088 -74926 -27036 -74874
rect -23088 -74924 -23036 -74872
rect -19088 -74924 -19036 -74872
rect -15088 -74924 -15036 -74872
rect -11088 -74926 -11036 -74874
rect -7088 -74926 -7036 -74874
rect -3088 -74924 -3036 -74872
rect 912 -74924 964 -74872
rect 4912 -74922 4964 -74870
<< metal2 >>
rect 53114 -40017 53174 -40011
rect 52006 -40021 53174 -40017
rect 52006 -40073 53118 -40021
rect 53170 -40073 53174 -40021
rect 52006 -40077 53174 -40073
rect 53114 -40083 53174 -40077
rect -14318 -40796 -14218 -40765
rect -14318 -40852 -14296 -40796
rect -14240 -40852 -14218 -40796
rect -7399 -40852 -7309 -40848
rect -15855 -41124 -15765 -41120
rect -14318 -41124 -14218 -40852
rect -7404 -40874 -5210 -40852
rect -7404 -40930 -7382 -40874
rect -7326 -40930 -5210 -40874
rect -7404 -40952 -5210 -40930
rect -7399 -40956 -7309 -40952
rect -7973 -41094 -7883 -41090
rect -15860 -41146 -14218 -41124
rect -15860 -41202 -15838 -41146
rect -15782 -41202 -14218 -41146
rect -13177 -41116 -7878 -41094
rect -13177 -41172 -13146 -41116
rect -13090 -41172 -7956 -41116
rect -7900 -41172 -7878 -41116
rect -13177 -41194 -7878 -41172
rect -5310 -41168 -5210 -40952
rect -7973 -41198 -7883 -41194
rect -15860 -41224 -14218 -41202
rect -5310 -41224 -5288 -41168
rect -5232 -41224 -5210 -41168
rect 49182 -41108 49290 -41091
rect 49182 -41164 49208 -41108
rect 49264 -41164 49290 -41108
rect 49182 -41181 49290 -41164
rect 51909 -41108 53320 -41106
rect 51909 -41164 51920 -41108
rect 51976 -41164 53320 -41108
rect 51909 -41166 53320 -41164
rect -15855 -41228 -15765 -41224
rect -5310 -41255 -5210 -41224
rect 30126 -41244 30198 -41240
rect 30126 -41296 30136 -41244
rect 30188 -41296 30198 -41244
rect 30126 -41300 30198 -41296
rect 30132 -41822 30192 -41300
rect 30126 -41826 30198 -41822
rect 30126 -41878 30136 -41826
rect 30188 -41878 30198 -41826
rect 30126 -41882 30198 -41878
rect 52380 -41962 52440 -41953
rect 52380 -41964 52500 -41962
rect 52380 -42020 52382 -41964
rect 52438 -42020 52500 -41964
rect 52380 -42022 52500 -42020
rect 57128 -41988 57200 -41984
rect 52380 -42031 52440 -42022
rect 57128 -42040 57138 -41988
rect 57190 -42040 57200 -41988
rect 58200 -41992 58452 -41932
rect 57128 -42044 57200 -42040
rect 57134 -42132 57194 -42044
rect 57134 -42192 58450 -42132
rect -14632 -42469 -14532 -42464
rect -14636 -42486 -14528 -42469
rect -14636 -42542 -14610 -42486
rect -14554 -42542 -14528 -42486
rect 51994 -42484 53383 -42482
rect -6432 -42537 -6332 -42532
rect -14636 -42559 -14528 -42542
rect -6436 -42554 -6328 -42537
rect 51994 -42540 53316 -42484
rect 53372 -42540 53383 -42484
rect 51994 -42542 53383 -42540
rect -14632 -47446 -14532 -42559
rect -6436 -42610 -6410 -42554
rect -6354 -42610 -6328 -42554
rect -6436 -42627 -6328 -42610
rect -11643 -42836 -11553 -42832
rect -9531 -42836 -9441 -42832
rect -13746 -42858 -11548 -42836
rect -13746 -42914 -11626 -42858
rect -11570 -42914 -11548 -42858
rect -13746 -42936 -11548 -42914
rect -9536 -42858 -7342 -42836
rect -9536 -42914 -9514 -42858
rect -9458 -42914 -7342 -42858
rect -9536 -42936 -7342 -42914
rect -13746 -43142 -13646 -42936
rect -11643 -42940 -11553 -42936
rect -9531 -42940 -9441 -42936
rect -13746 -43198 -13724 -43142
rect -13668 -43198 -13646 -43142
rect -13746 -43229 -13646 -43198
rect -7442 -43134 -7342 -42936
rect -7442 -43190 -7420 -43134
rect -7364 -43190 -7342 -43134
rect -7442 -43221 -7342 -43190
rect -10917 -44832 -10827 -44828
rect -10922 -44854 -10064 -44832
rect -10922 -44910 -10900 -44854
rect -10844 -44910 -10064 -44854
rect -10922 -44932 -10064 -44910
rect -10917 -44936 -10827 -44932
rect -10164 -45146 -10064 -44932
rect -10164 -45202 -10142 -45146
rect -10086 -45202 -10064 -45146
rect -10164 -45233 -10064 -45202
rect -7444 -46780 -7344 -46749
rect -13741 -46836 -13651 -46832
rect -7444 -46836 -7422 -46780
rect -7366 -46836 -7344 -46780
rect -13746 -46858 -11544 -46836
rect -13746 -46914 -13724 -46858
rect -13668 -46914 -11544 -46858
rect -13746 -46936 -11544 -46914
rect -13741 -46940 -13651 -46936
rect -11644 -47156 -11544 -46936
rect -9537 -47104 -9447 -47100
rect -7444 -47104 -7344 -46836
rect -11644 -47212 -11622 -47156
rect -11566 -47212 -11544 -47156
rect -9542 -47126 -7344 -47104
rect -9542 -47182 -9520 -47126
rect -9464 -47182 -7344 -47126
rect -9542 -47204 -7344 -47182
rect -9537 -47208 -9447 -47204
rect -11644 -47243 -11544 -47212
rect -14632 -47502 -14610 -47446
rect -14554 -47502 -14532 -47446
rect -14632 -47533 -14532 -47502
rect -6432 -47552 -6332 -42627
rect 26986 -42944 27046 -42933
rect 26986 -43000 26988 -42944
rect 27044 -43000 27046 -42944
rect 26986 -43098 27046 -43000
rect 26986 -45104 27046 -45098
rect 27780 -45104 27840 -45098
rect 26986 -45108 27840 -45104
rect 26986 -45160 26990 -45108
rect 27042 -45160 27784 -45108
rect 27836 -45160 27840 -45108
rect 26986 -45164 27840 -45160
rect 26986 -45170 27046 -45164
rect 27780 -45170 27840 -45164
rect 26986 -46860 27046 -46854
rect 27780 -46860 27840 -46854
rect 26986 -46864 27840 -46860
rect 26986 -46916 26990 -46864
rect 27042 -46916 27784 -46864
rect 27836 -46916 27840 -46864
rect 26986 -46920 27840 -46916
rect 26986 -46926 27046 -46920
rect 27780 -46926 27840 -46920
rect -6432 -47608 -6410 -47552
rect -6354 -47608 -6332 -47552
rect -6432 -47639 -6332 -47608
rect 26986 -48374 27046 -48368
rect 26986 -48378 27900 -48374
rect 26986 -48430 26990 -48378
rect 27042 -48430 27900 -48378
rect 26986 -48434 27900 -48430
rect 26986 -48440 27046 -48434
rect -5312 -48800 -5212 -48769
rect -15855 -48852 -15765 -48848
rect -12999 -48850 -12909 -48846
rect -8060 -48850 -7960 -48841
rect -15860 -48874 -13656 -48852
rect -15860 -48930 -15838 -48874
rect -15782 -48930 -13656 -48874
rect -15860 -48952 -13656 -48930
rect -13004 -48872 -7960 -48850
rect -13004 -48928 -12982 -48872
rect -12926 -48928 -8038 -48872
rect -7982 -48928 -7960 -48872
rect -13004 -48950 -7960 -48928
rect -15855 -48956 -15765 -48952
rect -13756 -49170 -13656 -48952
rect -12999 -48954 -12909 -48950
rect -8060 -48959 -7960 -48950
rect -5312 -48856 -5290 -48800
rect -5234 -48856 -5212 -48800
rect -7431 -49046 -7341 -49042
rect -5312 -49046 -5212 -48856
rect -7436 -49068 -5212 -49046
rect -7436 -49124 -7414 -49068
rect -7358 -49124 -5212 -49068
rect -7436 -49146 -5212 -49124
rect -7431 -49150 -7341 -49146
rect -13756 -49226 -13734 -49170
rect -13678 -49226 -13656 -49170
rect -13756 -49257 -13656 -49226
rect 26982 -49616 27042 -49610
rect 26982 -49620 28044 -49616
rect 26982 -49672 26986 -49620
rect 27038 -49672 28044 -49620
rect 26982 -49676 28044 -49672
rect 26982 -49682 27042 -49676
rect 26986 -50852 27046 -50846
rect 26986 -50856 28070 -50852
rect 26986 -50908 26990 -50856
rect 27042 -50908 28070 -50856
rect 26986 -50912 28070 -50908
rect 26986 -50918 27046 -50912
rect 14775 -52004 14865 -51978
rect 14775 -52060 14792 -52004
rect 14848 -52060 14865 -52004
rect 14775 -52086 14865 -52060
rect 14767 -52948 14857 -52944
rect 14756 -52970 14868 -52948
rect 27782 -52962 27842 -52956
rect 14756 -53026 14784 -52970
rect 14840 -53026 14868 -52970
rect 26732 -52966 27842 -52962
rect 26732 -53018 27786 -52966
rect 27838 -53018 27842 -52966
rect 26732 -53022 27842 -53018
rect 14756 -53048 14868 -53026
rect 27782 -53028 27842 -53022
rect 14767 -53052 14857 -53048
rect 26380 -53564 26440 -53558
rect 27780 -53564 27840 -53558
rect 26380 -53568 27840 -53564
rect 26380 -53620 26384 -53568
rect 26436 -53620 27784 -53568
rect 27836 -53620 27840 -53568
rect 26380 -53624 27840 -53620
rect 26380 -53630 26440 -53624
rect 27780 -53630 27840 -53624
rect 14769 -53942 14859 -53938
rect 14758 -53964 14870 -53942
rect 14758 -54020 14786 -53964
rect 14842 -54020 14870 -53964
rect 14758 -54042 14870 -54020
rect 14769 -54046 14859 -54042
rect 14769 -54948 14859 -54944
rect 14758 -54970 14870 -54948
rect 14758 -55026 14786 -54970
rect 14842 -55026 14870 -54970
rect 14758 -55048 14870 -55026
rect 14769 -55052 14859 -55048
rect 27780 -55396 27840 -55390
rect 26320 -55400 27840 -55396
rect 26320 -55452 27784 -55400
rect 27836 -55452 27840 -55400
rect 26320 -55456 27840 -55452
rect 27780 -55462 27840 -55456
rect 14779 -56356 14869 -56330
rect 14779 -56412 14796 -56356
rect 14852 -56412 14869 -56356
rect 14779 -56438 14869 -56412
rect 9350 -56733 9452 -56700
rect 9350 -56789 9376 -56733
rect 9432 -56789 9452 -56733
rect 11554 -56724 12236 -56720
rect 11554 -56776 11564 -56724
rect 11616 -56776 12236 -56724
rect 11554 -56780 12236 -56776
rect 9350 -56795 9378 -56789
rect 9430 -56795 9452 -56789
rect 9350 -56807 9452 -56795
rect 9350 -56813 9378 -56807
rect 9430 -56813 9452 -56807
rect 9350 -56869 9376 -56813
rect 9432 -56869 9452 -56813
rect 9350 -56871 9452 -56869
rect 9350 -56893 9378 -56871
rect 9430 -56893 9452 -56871
rect 9350 -56949 9376 -56893
rect 9432 -56949 9452 -56893
rect 9350 -56973 9378 -56949
rect 9430 -56973 9452 -56949
rect 9350 -57029 9376 -56973
rect 9432 -57029 9452 -56973
rect 9350 -57051 9378 -57029
rect 9430 -57051 9452 -57029
rect 9350 -57053 9452 -57051
rect 9350 -57109 9376 -57053
rect 9432 -57109 9452 -57053
rect 9350 -57115 9378 -57109
rect 9430 -57115 9452 -57109
rect 9350 -57127 9452 -57115
rect 9350 -57133 9378 -57127
rect 9430 -57133 9452 -57127
rect 9350 -57189 9376 -57133
rect 9432 -57189 9452 -57133
rect 9350 -57191 9452 -57189
rect 9350 -57213 9378 -57191
rect 9430 -57213 9452 -57191
rect 9350 -57269 9376 -57213
rect 9432 -57269 9452 -57213
rect 9350 -57293 9378 -57269
rect 9430 -57293 9452 -57269
rect 9350 -57349 9376 -57293
rect 9432 -57349 9452 -57293
rect 9350 -57371 9378 -57349
rect 9430 -57371 9452 -57349
rect 9350 -57373 9452 -57371
rect 9350 -57429 9376 -57373
rect 9432 -57429 9452 -57373
rect 9350 -57435 9378 -57429
rect 9430 -57435 9452 -57429
rect 9350 -57447 9452 -57435
rect 9350 -57453 9378 -57447
rect 9430 -57453 9452 -57447
rect 9350 -57509 9376 -57453
rect 9432 -57509 9452 -57453
rect 9350 -57536 9452 -57509
rect 10912 -57486 10972 -57480
rect 11430 -57486 11490 -57480
rect 10912 -57490 11490 -57486
rect 10912 -57542 10916 -57490
rect 10968 -57542 11434 -57490
rect 11486 -57542 11490 -57490
rect 12176 -57532 12236 -56780
rect 12524 -57532 12584 -57523
rect 10912 -57546 11490 -57542
rect 10912 -57552 10972 -57546
rect 11430 -57552 11490 -57546
rect 12170 -57536 12242 -57532
rect 12170 -57588 12180 -57536
rect 12232 -57588 12242 -57536
rect 12170 -57592 12242 -57588
rect 12518 -57534 12590 -57532
rect 12518 -57590 12526 -57534
rect 12582 -57590 12590 -57534
rect 12518 -57592 12590 -57590
rect 12524 -57601 12584 -57592
rect 10654 -57635 10714 -57629
rect 11170 -57635 11230 -57629
rect 10643 -57637 11754 -57635
rect 10643 -57693 10654 -57637
rect 10710 -57639 11754 -57637
rect 10710 -57691 11174 -57639
rect 11226 -57691 11692 -57639
rect 11744 -57691 11754 -57639
rect 10710 -57693 11754 -57691
rect 10643 -57695 11754 -57693
rect 10654 -57701 10714 -57695
rect 11170 -57701 11230 -57695
rect 10914 -58078 10974 -58068
rect 10914 -58130 10918 -58078
rect 10970 -58130 10974 -58078
rect 10914 -58286 10974 -58130
rect 11430 -58078 11490 -58068
rect 11430 -58130 11434 -58078
rect 11486 -58130 11490 -58078
rect 11430 -58286 11490 -58130
rect 11558 -58183 11618 -58177
rect 11558 -58185 12595 -58183
rect 11558 -58187 12528 -58185
rect 11558 -58239 11562 -58187
rect 11614 -58239 12528 -58187
rect 11558 -58241 12528 -58239
rect 12584 -58241 12595 -58185
rect 11558 -58243 12595 -58241
rect 11558 -58249 11618 -58243
rect 10914 -58346 13076 -58286
rect 10276 -58433 12130 -58390
rect 10276 -58489 10294 -58433
rect 10350 -58435 10374 -58433
rect 10430 -58435 10454 -58433
rect 10510 -58435 10534 -58433
rect 10590 -58435 10614 -58433
rect 10670 -58435 10694 -58433
rect 10750 -58435 10774 -58433
rect 10830 -58435 10854 -58433
rect 10910 -58435 10934 -58433
rect 10990 -58435 11014 -58433
rect 11070 -58435 11094 -58433
rect 11150 -58435 11174 -58433
rect 11230 -58435 11254 -58433
rect 11310 -58435 11334 -58433
rect 11390 -58435 11414 -58433
rect 11470 -58435 11494 -58433
rect 11550 -58435 11574 -58433
rect 11630 -58435 11654 -58433
rect 11710 -58435 11734 -58433
rect 11790 -58435 11814 -58433
rect 11870 -58435 11894 -58433
rect 11950 -58435 11974 -58433
rect 12030 -58435 12054 -58433
rect 10364 -58487 10374 -58435
rect 10430 -58487 10440 -58435
rect 10684 -58487 10694 -58435
rect 10750 -58487 10760 -58435
rect 11004 -58487 11014 -58435
rect 11070 -58487 11080 -58435
rect 11324 -58487 11334 -58435
rect 11390 -58487 11400 -58435
rect 11644 -58487 11654 -58435
rect 11710 -58487 11720 -58435
rect 11964 -58487 11974 -58435
rect 12030 -58487 12040 -58435
rect 10350 -58489 10374 -58487
rect 10430 -58489 10454 -58487
rect 10510 -58489 10534 -58487
rect 10590 -58489 10614 -58487
rect 10670 -58489 10694 -58487
rect 10750 -58489 10774 -58487
rect 10830 -58489 10854 -58487
rect 10910 -58489 10934 -58487
rect 10990 -58489 11014 -58487
rect 11070 -58489 11094 -58487
rect 11150 -58489 11174 -58487
rect 11230 -58489 11254 -58487
rect 11310 -58489 11334 -58487
rect 11390 -58489 11414 -58487
rect 11470 -58489 11494 -58487
rect 11550 -58489 11574 -58487
rect 11630 -58489 11654 -58487
rect 11710 -58489 11734 -58487
rect 11790 -58489 11814 -58487
rect 11870 -58489 11894 -58487
rect 11950 -58489 11974 -58487
rect 12030 -58489 12054 -58487
rect 12110 -58489 12130 -58433
rect 10276 -58528 12130 -58489
rect 13016 -59714 13076 -58346
rect 13007 -59716 13085 -59714
rect 13007 -59772 13018 -59716
rect 13074 -59772 13085 -59716
rect 13007 -59774 13085 -59772
rect -9207 -64028 -9129 -64026
rect -9207 -64084 -9196 -64028
rect -9140 -64084 -9129 -64028
rect -9207 -64086 -9129 -64084
rect -25195 -65212 -25105 -65186
rect -25195 -65214 -25178 -65212
rect -26400 -65268 -25178 -65214
rect -25122 -65268 -25105 -65212
rect -21031 -65214 -20941 -65188
rect -17109 -65214 -17019 -65188
rect -26400 -65274 -25105 -65268
rect -22446 -65270 -21014 -65214
rect -20958 -65270 -20941 -65214
rect -22446 -65274 -20941 -65270
rect -18454 -65270 -17092 -65214
rect -17036 -65270 -17019 -65214
rect -18454 -65274 -17019 -65270
rect -25195 -65294 -25105 -65274
rect -21031 -65296 -20941 -65274
rect -17109 -65296 -17019 -65274
rect -16087 -65214 -15997 -65188
rect -9198 -65214 -9138 -64086
rect -4097 -65214 -4007 -65188
rect -39 -65214 51 -65192
rect 4015 -65214 4105 -65190
rect -16087 -65270 -16070 -65214
rect -16014 -65270 -14694 -65214
rect -16087 -65274 -14694 -65270
rect -10484 -65274 -9138 -65214
rect -7965 -65216 -6710 -65214
rect -7965 -65272 -7954 -65216
rect -7898 -65272 -6710 -65216
rect -7965 -65274 -6710 -65272
rect -4097 -65270 -4080 -65214
rect -4024 -65270 -2662 -65214
rect -4097 -65274 -2662 -65270
rect -39 -65218 1320 -65214
rect -39 -65274 -22 -65218
rect 34 -65274 1320 -65218
rect 4015 -65216 5342 -65214
rect 4015 -65272 4032 -65216
rect 4088 -65272 5342 -65216
rect 4015 -65274 5342 -65272
rect -16087 -65296 -15997 -65274
rect -4097 -65296 -4007 -65274
rect -39 -65300 51 -65274
rect 4015 -65298 4105 -65274
rect -26630 -65448 -26379 -65446
rect -26630 -65504 -26446 -65448
rect -26390 -65504 -26379 -65448
rect -26630 -65506 -26379 -65504
rect -22516 -65448 -22379 -65446
rect -22516 -65504 -22446 -65448
rect -22390 -65504 -22379 -65448
rect -22516 -65506 -22379 -65504
rect -18518 -65448 -18381 -65446
rect -18518 -65504 -18448 -65448
rect -18392 -65504 -18381 -65448
rect -18518 -65506 -18381 -65504
rect -14522 -65448 -14381 -65446
rect -14522 -65504 -14448 -65448
rect -14392 -65504 -14381 -65448
rect -14522 -65506 -14381 -65504
rect -10518 -65448 -10381 -65446
rect -10518 -65504 -10448 -65448
rect -10392 -65504 -10381 -65448
rect -10518 -65506 -10381 -65504
rect -6522 -65448 -6379 -65446
rect -6522 -65504 -6446 -65448
rect -6390 -65504 -6379 -65448
rect -6522 -65506 -6379 -65504
rect -2518 -65448 -2383 -65446
rect -2518 -65504 -2450 -65448
rect -2394 -65504 -2383 -65448
rect -2518 -65506 -2383 -65504
rect 1476 -65448 1621 -65446
rect 1476 -65504 1554 -65448
rect 1610 -65504 1621 -65448
rect 1476 -65506 1621 -65504
rect 5490 -65448 5623 -65446
rect 5490 -65504 5556 -65448
rect 5612 -65504 5623 -65448
rect 5490 -65506 5623 -65504
rect -26578 -67920 -26518 -67858
rect -22578 -67920 -22518 -67856
rect -18578 -67920 -18518 -67858
rect -14578 -67920 -14518 -67854
rect -10578 -67920 -10518 -67854
rect -6578 -67920 -6518 -67854
rect -2578 -67920 -2518 -67858
rect 1422 -67920 1482 -67854
rect -26587 -67922 -26509 -67920
rect -26587 -67978 -26576 -67922
rect -26520 -67978 -26509 -67922
rect -26587 -67980 -26509 -67978
rect -22587 -67922 -22509 -67920
rect -22587 -67978 -22576 -67922
rect -22520 -67978 -22509 -67922
rect -22587 -67980 -22509 -67978
rect -18587 -67922 -18509 -67920
rect -18587 -67978 -18576 -67922
rect -18520 -67978 -18509 -67922
rect -18587 -67980 -18509 -67978
rect -14587 -67922 -14509 -67920
rect -14587 -67978 -14576 -67922
rect -14520 -67978 -14509 -67922
rect -14587 -67980 -14509 -67978
rect -10587 -67922 -10509 -67920
rect -10587 -67978 -10576 -67922
rect -10520 -67978 -10509 -67922
rect -10587 -67980 -10509 -67978
rect -6587 -67922 -6509 -67920
rect -6587 -67978 -6576 -67922
rect -6520 -67978 -6509 -67922
rect -6587 -67980 -6509 -67978
rect -2587 -67922 -2509 -67920
rect -2587 -67978 -2576 -67922
rect -2520 -67978 -2509 -67922
rect -2587 -67980 -2509 -67978
rect 1413 -67922 1491 -67920
rect 5422 -67922 5482 -67860
rect 1413 -67978 1424 -67922
rect 1480 -67978 1491 -67922
rect 1413 -67980 1491 -67978
rect 5413 -67924 5491 -67922
rect 5413 -67980 5424 -67924
rect 5480 -67980 5491 -67924
rect 5413 -67982 5491 -67980
rect -26324 -68954 -25163 -68952
rect -26324 -69010 -25230 -68954
rect -25174 -69010 -25163 -68954
rect -26324 -69012 -25163 -69010
rect -22300 -68954 -21163 -68952
rect -22300 -69010 -21230 -68954
rect -21174 -69010 -21163 -68954
rect -22300 -69012 -21163 -69010
rect -18274 -68954 -17163 -68952
rect -18274 -69010 -17230 -68954
rect -17174 -69010 -17163 -68954
rect -18274 -69012 -17163 -69010
rect -14234 -68954 -13163 -68952
rect -14234 -69010 -13230 -68954
rect -13174 -69010 -13163 -68954
rect -14234 -69012 -13163 -69010
rect -10196 -68954 -9163 -68952
rect -10196 -69010 -9230 -68954
rect -9174 -69010 -9163 -68954
rect -10196 -69012 -9163 -69010
rect -6386 -68954 -5163 -68952
rect -6386 -69010 -5230 -68954
rect -5174 -69010 -5163 -68954
rect -6386 -69012 -5163 -69010
rect -2252 -68954 -1163 -68952
rect -2252 -69010 -1230 -68954
rect -1174 -69010 -1163 -68954
rect -2252 -69012 -1163 -69010
rect 1768 -68954 2837 -68952
rect 1768 -69010 2770 -68954
rect 2826 -69010 2837 -68954
rect 1768 -69012 2837 -69010
rect 5834 -68954 6837 -68952
rect 5834 -69010 6770 -68954
rect 6826 -69010 6837 -68954
rect 5834 -69012 6837 -69010
rect -25238 -72106 -25178 -72097
rect -21238 -72106 -21178 -72097
rect -17238 -72106 -17178 -72097
rect -13238 -72106 -13178 -72097
rect -9238 -72106 -9178 -72097
rect -5238 -72106 -5178 -72097
rect -1238 -72106 -1178 -72097
rect 2762 -72106 2822 -72097
rect 6762 -72106 6822 -72097
rect -26424 -72108 -25178 -72106
rect -26424 -72164 -25236 -72108
rect -25180 -72164 -25178 -72108
rect -26424 -72166 -25178 -72164
rect -22452 -72108 -21178 -72106
rect -22452 -72164 -21236 -72108
rect -21180 -72164 -21178 -72108
rect -22452 -72166 -21178 -72164
rect -18416 -72108 -17178 -72106
rect -18416 -72164 -17236 -72108
rect -17180 -72164 -17178 -72108
rect -18416 -72166 -17178 -72164
rect -14438 -72108 -13178 -72106
rect -14438 -72164 -13236 -72108
rect -13180 -72164 -13178 -72108
rect -14438 -72166 -13178 -72164
rect -10442 -72108 -9178 -72106
rect -10442 -72164 -9236 -72108
rect -9180 -72164 -9178 -72108
rect -10442 -72166 -9178 -72164
rect -6444 -72108 -5178 -72106
rect -6444 -72164 -5236 -72108
rect -5180 -72164 -5178 -72108
rect -6444 -72166 -5178 -72164
rect -2442 -72108 -1178 -72106
rect -2442 -72164 -1236 -72108
rect -1180 -72164 -1178 -72108
rect -2442 -72166 -1178 -72164
rect 1550 -72108 2822 -72106
rect 1550 -72164 2764 -72108
rect 2820 -72164 2822 -72108
rect 1550 -72166 2822 -72164
rect 5566 -72108 6822 -72106
rect 5566 -72164 6764 -72108
rect 6820 -72164 6822 -72108
rect 5566 -72166 6822 -72164
rect -25238 -72175 -25178 -72166
rect -21238 -72175 -21178 -72166
rect -17238 -72175 -17178 -72166
rect -13238 -72175 -13178 -72166
rect -9238 -72175 -9178 -72166
rect -5238 -72175 -5178 -72166
rect -1238 -72175 -1178 -72166
rect 2762 -72175 2822 -72166
rect 6762 -72175 6822 -72166
rect -3246 -72336 -3186 -72326
rect -3246 -72388 -3242 -72336
rect -3190 -72388 -3186 -72336
rect -3246 -72552 -3186 -72388
rect -27094 -72882 -27034 -72800
rect -23094 -72882 -23034 -72808
rect -19094 -72882 -19034 -72780
rect -15094 -72882 -15034 -72776
rect -11094 -72880 -11034 -72786
rect -11103 -72882 -11025 -72880
rect -7094 -72882 -7034 -72796
rect -3094 -72882 -3034 -72788
rect 906 -72882 966 -72786
rect -27103 -72884 -27025 -72882
rect -27103 -72940 -27092 -72884
rect -27036 -72940 -27025 -72884
rect -27103 -72942 -27025 -72940
rect -23103 -72884 -23025 -72882
rect -23103 -72940 -23092 -72884
rect -23036 -72940 -23025 -72884
rect -23103 -72942 -23025 -72940
rect -19103 -72884 -19025 -72882
rect -19103 -72940 -19092 -72884
rect -19036 -72940 -19025 -72884
rect -19103 -72942 -19025 -72940
rect -15103 -72884 -15025 -72882
rect -15103 -72940 -15092 -72884
rect -15036 -72940 -15025 -72884
rect -11103 -72938 -11092 -72882
rect -11036 -72938 -11025 -72882
rect -11103 -72940 -11025 -72938
rect -7103 -72884 -7025 -72882
rect -7103 -72940 -7092 -72884
rect -7036 -72940 -7025 -72884
rect -15103 -72942 -15025 -72940
rect -7103 -72942 -7025 -72940
rect -3103 -72884 -3025 -72882
rect -3103 -72940 -3092 -72884
rect -3036 -72940 -3025 -72884
rect -3103 -72942 -3025 -72940
rect 897 -72884 975 -72882
rect 897 -72940 908 -72884
rect 964 -72940 975 -72884
rect 897 -72942 975 -72940
rect 4897 -72884 4975 -72882
rect 4897 -72940 4908 -72884
rect 4964 -72940 4975 -72884
rect 4897 -72942 4975 -72940
rect -27092 -74870 -27032 -74864
rect -23092 -74868 -23032 -74862
rect -19092 -74868 -19032 -74862
rect -15092 -74868 -15032 -74862
rect -23101 -74870 -23023 -74868
rect -27101 -74872 -27023 -74870
rect -27101 -74928 -27090 -74872
rect -27034 -74928 -27023 -74872
rect -23101 -74926 -23090 -74870
rect -23034 -74926 -23023 -74870
rect -23101 -74928 -23023 -74926
rect -19101 -74870 -19023 -74868
rect -19101 -74926 -19090 -74870
rect -19034 -74926 -19023 -74870
rect -19101 -74928 -19023 -74926
rect -15101 -74870 -15023 -74868
rect -11092 -74870 -11032 -74864
rect -7092 -74870 -7032 -74864
rect -3092 -74868 -3032 -74862
rect 908 -74868 968 -74862
rect 4908 -74866 4968 -74860
rect 4899 -74868 4977 -74866
rect -3101 -74870 -3023 -74868
rect -15101 -74926 -15090 -74870
rect -15034 -74926 -15023 -74870
rect -15101 -74928 -15023 -74926
rect -11101 -74872 -11023 -74870
rect -11101 -74928 -11090 -74872
rect -11034 -74928 -11023 -74872
rect -27101 -74930 -27023 -74928
rect -27092 -74936 -27032 -74930
rect -23092 -74934 -23032 -74928
rect -19092 -74934 -19032 -74928
rect -15092 -74934 -15032 -74928
rect -11101 -74930 -11023 -74928
rect -7101 -74872 -7023 -74870
rect -7101 -74928 -7090 -74872
rect -7034 -74928 -7023 -74872
rect -3101 -74926 -3090 -74870
rect -3034 -74926 -3023 -74870
rect -3101 -74928 -3023 -74926
rect 899 -74870 977 -74868
rect 899 -74926 910 -74870
rect 966 -74926 977 -74870
rect 4899 -74924 4910 -74868
rect 4966 -74924 4977 -74868
rect 4899 -74926 4977 -74924
rect 899 -74928 977 -74926
rect -7101 -74930 -7023 -74928
rect -11092 -74936 -11032 -74930
rect -7092 -74936 -7032 -74930
rect -3092 -74934 -3032 -74928
rect 908 -74934 968 -74928
rect 4908 -74932 4968 -74926
<< via2 >>
rect -14296 -40852 -14240 -40796
rect -7382 -40930 -7326 -40874
rect -15838 -41202 -15782 -41146
rect -13146 -41172 -13090 -41116
rect -7956 -41172 -7900 -41116
rect -5288 -41224 -5232 -41168
rect 49208 -41164 49264 -41108
rect 51920 -41164 51976 -41108
rect 52382 -42020 52438 -41964
rect -14610 -42542 -14554 -42486
rect 53316 -42540 53372 -42484
rect -6410 -42610 -6354 -42554
rect -11626 -42914 -11570 -42858
rect -9514 -42914 -9458 -42858
rect -13724 -43198 -13668 -43142
rect -7420 -43190 -7364 -43134
rect -10900 -44910 -10844 -44854
rect -10142 -45202 -10086 -45146
rect -7422 -46836 -7366 -46780
rect -13724 -46914 -13668 -46858
rect -11622 -47212 -11566 -47156
rect -9520 -47182 -9464 -47126
rect -14610 -47502 -14554 -47446
rect 26988 -43000 27044 -42944
rect -6410 -47608 -6354 -47552
rect -15838 -48930 -15782 -48874
rect -12982 -48928 -12926 -48872
rect -8038 -48928 -7982 -48872
rect -5290 -48856 -5234 -48800
rect -7414 -49124 -7358 -49068
rect -13734 -49226 -13678 -49170
rect 14792 -52060 14848 -52004
rect 14784 -52972 14840 -52970
rect 14784 -53024 14786 -52972
rect 14786 -53024 14838 -52972
rect 14838 -53024 14840 -52972
rect 14784 -53026 14840 -53024
rect 14786 -53966 14842 -53964
rect 14786 -54018 14788 -53966
rect 14788 -54018 14840 -53966
rect 14840 -54018 14842 -53966
rect 14786 -54020 14842 -54018
rect 14786 -54972 14842 -54970
rect 14786 -55024 14788 -54972
rect 14788 -55024 14840 -54972
rect 14840 -55024 14842 -54972
rect 14786 -55026 14842 -55024
rect 14796 -56412 14852 -56356
rect 9376 -56743 9432 -56733
rect 9376 -56789 9378 -56743
rect 9378 -56789 9430 -56743
rect 9430 -56789 9432 -56743
rect 9376 -56859 9378 -56813
rect 9378 -56859 9430 -56813
rect 9430 -56859 9432 -56813
rect 9376 -56869 9432 -56859
rect 9376 -56923 9378 -56893
rect 9378 -56923 9430 -56893
rect 9430 -56923 9432 -56893
rect 9376 -56935 9432 -56923
rect 9376 -56949 9378 -56935
rect 9378 -56949 9430 -56935
rect 9430 -56949 9432 -56935
rect 9376 -56987 9378 -56973
rect 9378 -56987 9430 -56973
rect 9430 -56987 9432 -56973
rect 9376 -56999 9432 -56987
rect 9376 -57029 9378 -56999
rect 9378 -57029 9430 -56999
rect 9430 -57029 9432 -56999
rect 9376 -57063 9432 -57053
rect 9376 -57109 9378 -57063
rect 9378 -57109 9430 -57063
rect 9430 -57109 9432 -57063
rect 9376 -57179 9378 -57133
rect 9378 -57179 9430 -57133
rect 9430 -57179 9432 -57133
rect 9376 -57189 9432 -57179
rect 9376 -57243 9378 -57213
rect 9378 -57243 9430 -57213
rect 9430 -57243 9432 -57213
rect 9376 -57255 9432 -57243
rect 9376 -57269 9378 -57255
rect 9378 -57269 9430 -57255
rect 9430 -57269 9432 -57255
rect 9376 -57307 9378 -57293
rect 9378 -57307 9430 -57293
rect 9430 -57307 9432 -57293
rect 9376 -57319 9432 -57307
rect 9376 -57349 9378 -57319
rect 9378 -57349 9430 -57319
rect 9430 -57349 9432 -57319
rect 9376 -57383 9432 -57373
rect 9376 -57429 9378 -57383
rect 9378 -57429 9430 -57383
rect 9430 -57429 9432 -57383
rect 9376 -57499 9378 -57453
rect 9378 -57499 9430 -57453
rect 9430 -57499 9432 -57453
rect 9376 -57509 9432 -57499
rect 12526 -57536 12582 -57534
rect 12526 -57588 12528 -57536
rect 12528 -57588 12580 -57536
rect 12580 -57588 12582 -57536
rect 12526 -57590 12582 -57588
rect 10654 -57639 10710 -57637
rect 10654 -57691 10658 -57639
rect 10658 -57691 10710 -57639
rect 10654 -57693 10710 -57691
rect 12528 -58241 12584 -58185
rect 10294 -58435 10350 -58433
rect 10374 -58435 10430 -58433
rect 10454 -58435 10510 -58433
rect 10534 -58435 10590 -58433
rect 10614 -58435 10670 -58433
rect 10694 -58435 10750 -58433
rect 10774 -58435 10830 -58433
rect 10854 -58435 10910 -58433
rect 10934 -58435 10990 -58433
rect 11014 -58435 11070 -58433
rect 11094 -58435 11150 -58433
rect 11174 -58435 11230 -58433
rect 11254 -58435 11310 -58433
rect 11334 -58435 11390 -58433
rect 11414 -58435 11470 -58433
rect 11494 -58435 11550 -58433
rect 11574 -58435 11630 -58433
rect 11654 -58435 11710 -58433
rect 11734 -58435 11790 -58433
rect 11814 -58435 11870 -58433
rect 11894 -58435 11950 -58433
rect 11974 -58435 12030 -58433
rect 12054 -58435 12110 -58433
rect 10294 -58487 10312 -58435
rect 10312 -58487 10350 -58435
rect 10374 -58487 10376 -58435
rect 10376 -58487 10428 -58435
rect 10428 -58487 10430 -58435
rect 10454 -58487 10492 -58435
rect 10492 -58487 10504 -58435
rect 10504 -58487 10510 -58435
rect 10534 -58487 10556 -58435
rect 10556 -58487 10568 -58435
rect 10568 -58487 10590 -58435
rect 10614 -58487 10620 -58435
rect 10620 -58487 10632 -58435
rect 10632 -58487 10670 -58435
rect 10694 -58487 10696 -58435
rect 10696 -58487 10748 -58435
rect 10748 -58487 10750 -58435
rect 10774 -58487 10812 -58435
rect 10812 -58487 10824 -58435
rect 10824 -58487 10830 -58435
rect 10854 -58487 10876 -58435
rect 10876 -58487 10888 -58435
rect 10888 -58487 10910 -58435
rect 10934 -58487 10940 -58435
rect 10940 -58487 10952 -58435
rect 10952 -58487 10990 -58435
rect 11014 -58487 11016 -58435
rect 11016 -58487 11068 -58435
rect 11068 -58487 11070 -58435
rect 11094 -58487 11132 -58435
rect 11132 -58487 11144 -58435
rect 11144 -58487 11150 -58435
rect 11174 -58487 11196 -58435
rect 11196 -58487 11208 -58435
rect 11208 -58487 11230 -58435
rect 11254 -58487 11260 -58435
rect 11260 -58487 11272 -58435
rect 11272 -58487 11310 -58435
rect 11334 -58487 11336 -58435
rect 11336 -58487 11388 -58435
rect 11388 -58487 11390 -58435
rect 11414 -58487 11452 -58435
rect 11452 -58487 11464 -58435
rect 11464 -58487 11470 -58435
rect 11494 -58487 11516 -58435
rect 11516 -58487 11528 -58435
rect 11528 -58487 11550 -58435
rect 11574 -58487 11580 -58435
rect 11580 -58487 11592 -58435
rect 11592 -58487 11630 -58435
rect 11654 -58487 11656 -58435
rect 11656 -58487 11708 -58435
rect 11708 -58487 11710 -58435
rect 11734 -58487 11772 -58435
rect 11772 -58487 11784 -58435
rect 11784 -58487 11790 -58435
rect 11814 -58487 11836 -58435
rect 11836 -58487 11848 -58435
rect 11848 -58487 11870 -58435
rect 11894 -58487 11900 -58435
rect 11900 -58487 11912 -58435
rect 11912 -58487 11950 -58435
rect 11974 -58487 11976 -58435
rect 11976 -58487 12028 -58435
rect 12028 -58487 12030 -58435
rect 12054 -58487 12092 -58435
rect 12092 -58487 12110 -58435
rect 10294 -58489 10350 -58487
rect 10374 -58489 10430 -58487
rect 10454 -58489 10510 -58487
rect 10534 -58489 10590 -58487
rect 10614 -58489 10670 -58487
rect 10694 -58489 10750 -58487
rect 10774 -58489 10830 -58487
rect 10854 -58489 10910 -58487
rect 10934 -58489 10990 -58487
rect 11014 -58489 11070 -58487
rect 11094 -58489 11150 -58487
rect 11174 -58489 11230 -58487
rect 11254 -58489 11310 -58487
rect 11334 -58489 11390 -58487
rect 11414 -58489 11470 -58487
rect 11494 -58489 11550 -58487
rect 11574 -58489 11630 -58487
rect 11654 -58489 11710 -58487
rect 11734 -58489 11790 -58487
rect 11814 -58489 11870 -58487
rect 11894 -58489 11950 -58487
rect 11974 -58489 12030 -58487
rect 12054 -58489 12110 -58487
rect 13018 -59772 13074 -59716
rect -9196 -64084 -9140 -64028
rect -25178 -65268 -25122 -65212
rect -21014 -65270 -20958 -65214
rect -17092 -65270 -17036 -65214
rect -16070 -65270 -16014 -65214
rect -7954 -65272 -7898 -65216
rect -4080 -65270 -4024 -65214
rect -22 -65274 34 -65218
rect 4032 -65272 4088 -65216
rect -26446 -65504 -26390 -65448
rect -22446 -65504 -22390 -65448
rect -18448 -65504 -18392 -65448
rect -14448 -65504 -14392 -65448
rect -10448 -65504 -10392 -65448
rect -6446 -65504 -6390 -65448
rect -2450 -65504 -2394 -65448
rect 1554 -65504 1610 -65448
rect 5556 -65504 5612 -65448
rect -26576 -67978 -26520 -67922
rect -22576 -67978 -22520 -67922
rect -18576 -67978 -18520 -67922
rect -14576 -67978 -14520 -67922
rect -10576 -67978 -10520 -67922
rect -6576 -67978 -6520 -67922
rect -2576 -67978 -2520 -67922
rect 1424 -67978 1480 -67922
rect 5424 -67980 5480 -67924
rect -25230 -69010 -25174 -68954
rect -21230 -69010 -21174 -68954
rect -17230 -69010 -17174 -68954
rect -13230 -69010 -13174 -68954
rect -9230 -69010 -9174 -68954
rect -5230 -69010 -5174 -68954
rect -1230 -69010 -1174 -68954
rect 2770 -69010 2826 -68954
rect 6770 -69010 6826 -68954
rect -25236 -72164 -25180 -72108
rect -21236 -72164 -21180 -72108
rect -17236 -72164 -17180 -72108
rect -13236 -72164 -13180 -72108
rect -9236 -72164 -9180 -72108
rect -5236 -72164 -5180 -72108
rect -1236 -72164 -1180 -72108
rect 2764 -72164 2820 -72108
rect 6764 -72164 6820 -72108
rect -27092 -72940 -27036 -72884
rect -23092 -72940 -23036 -72884
rect -19092 -72940 -19036 -72884
rect -15092 -72940 -15036 -72884
rect -11092 -72938 -11036 -72882
rect -7092 -72940 -7036 -72884
rect -3092 -72940 -3036 -72884
rect 908 -72940 964 -72884
rect 4908 -72940 4964 -72884
rect -27090 -74874 -27034 -74872
rect -27090 -74926 -27088 -74874
rect -27088 -74926 -27036 -74874
rect -27036 -74926 -27034 -74874
rect -27090 -74928 -27034 -74926
rect -23090 -74872 -23034 -74870
rect -23090 -74924 -23088 -74872
rect -23088 -74924 -23036 -74872
rect -23036 -74924 -23034 -74872
rect -23090 -74926 -23034 -74924
rect -19090 -74872 -19034 -74870
rect -19090 -74924 -19088 -74872
rect -19088 -74924 -19036 -74872
rect -19036 -74924 -19034 -74872
rect -19090 -74926 -19034 -74924
rect -15090 -74872 -15034 -74870
rect -15090 -74924 -15088 -74872
rect -15088 -74924 -15036 -74872
rect -15036 -74924 -15034 -74872
rect -15090 -74926 -15034 -74924
rect -11090 -74874 -11034 -74872
rect -11090 -74926 -11088 -74874
rect -11088 -74926 -11036 -74874
rect -11036 -74926 -11034 -74874
rect -11090 -74928 -11034 -74926
rect -7090 -74874 -7034 -74872
rect -7090 -74926 -7088 -74874
rect -7088 -74926 -7036 -74874
rect -7036 -74926 -7034 -74874
rect -7090 -74928 -7034 -74926
rect -3090 -74872 -3034 -74870
rect -3090 -74924 -3088 -74872
rect -3088 -74924 -3036 -74872
rect -3036 -74924 -3034 -74872
rect -3090 -74926 -3034 -74924
rect 910 -74872 966 -74870
rect 910 -74924 912 -74872
rect 912 -74924 964 -74872
rect 964 -74924 966 -74872
rect 910 -74926 966 -74924
rect 4910 -74870 4966 -74868
rect 4910 -74922 4912 -74870
rect 4912 -74922 4964 -74870
rect 4964 -74922 4966 -74870
rect 4910 -74924 4966 -74922
<< metal3 >>
rect -24278 -29944 -24178 -29206
rect -22172 -29944 -22072 -29206
rect -20066 -29944 -19966 -29206
rect -17960 -29944 -17860 -29206
rect -15854 -29944 -15754 -29206
rect -13748 -29944 -13648 -29206
rect -11642 -29944 -11542 -29206
rect -9536 -29944 -9436 -29206
rect -7430 -29944 -7330 -29206
rect -5324 -29944 -5224 -29206
rect -3218 -29944 -3118 -29206
rect -1112 -29944 -1012 -29206
rect 3060 -29944 3160 -29942
rect -26452 -30044 5328 -29944
rect -26392 -31934 -26292 -30782
rect -24286 -31934 -24178 -30044
rect -22172 -31934 -22072 -30044
rect -20066 -31934 -19966 -30044
rect -17960 -31934 -17860 -30044
rect -15854 -31934 -15754 -30044
rect -13748 -31934 -13648 -30044
rect -11642 -31934 -11542 -30044
rect -9536 -31934 -9436 -30044
rect -7430 -31934 -7330 -30044
rect -5324 -31934 -5224 -30044
rect -3218 -31934 -3118 -30044
rect -1112 -31934 -1012 -30044
rect 994 -31900 1094 -30044
rect 964 -31934 1094 -31900
rect 3060 -31934 3160 -30044
rect -26450 -31950 3160 -31934
rect 5228 -31950 5328 -30044
rect -26450 -32034 6076 -31950
rect -26392 -33956 -26292 -32034
rect -24286 -32806 -24178 -32034
rect -22172 -32408 -22072 -32034
rect -22172 -32806 -22034 -32408
rect -20066 -32806 -19936 -32034
rect -17960 -32806 -17792 -32034
rect -15854 -32806 -15754 -32034
rect -13748 -32806 -13648 -32034
rect -11642 -32806 -11542 -32034
rect -9536 -32806 -9436 -32034
rect -7430 -32806 -7330 -32034
rect -5324 -32806 -5224 -32034
rect -3218 -32806 -3118 -32034
rect -1112 -32362 -1012 -32034
rect -1134 -32806 -1012 -32362
rect 964 -32078 1094 -32034
rect 2355 -32050 6076 -32034
rect -24286 -33956 -24186 -32806
rect -22134 -33956 -22034 -32806
rect -20036 -33956 -19936 -32806
rect -17892 -33956 -17792 -32806
rect -26392 -34056 -17792 -33956
rect -26392 -35916 -26292 -34056
rect -24286 -35916 -24186 -34056
rect -22180 -35916 -22080 -34056
rect -26392 -36016 -22080 -35916
rect -20078 -35958 -19978 -35928
rect -15854 -35958 -15754 -33872
rect -13748 -33920 -13648 -33206
rect -11642 -33920 -11542 -33206
rect -9536 -33920 -9436 -33206
rect -7430 -33920 -7330 -33206
rect -5324 -33920 -5224 -33206
rect -15046 -34020 -3164 -33920
rect -13748 -35958 -13648 -34020
rect -11642 -35958 -11542 -34020
rect -9536 -35958 -9436 -34020
rect -7430 -35958 -7330 -34020
rect -5324 -35958 -5224 -34020
rect -3264 -35958 -3164 -34020
rect -1134 -33950 -1034 -32806
rect 964 -33950 1064 -32078
rect 3060 -33950 3160 -32050
rect 5228 -33950 5328 -32050
rect -1134 -34050 6076 -33950
rect 964 -35934 1064 -34050
rect 964 -35950 2978 -35934
rect 3060 -35950 3160 -34050
rect 5228 -35950 5328 -34050
rect -26392 -37942 -26292 -36016
rect -24286 -37942 -24186 -36016
rect -20134 -36058 -994 -35958
rect 964 -36034 6076 -35950
rect -26392 -38042 -24186 -37942
rect -22154 -37980 -22054 -37968
rect -20078 -37980 -19978 -36058
rect -13748 -36806 -13648 -36058
rect -11642 -36806 -11542 -36058
rect -9536 -36806 -9436 -36058
rect -7430 -36806 -7330 -36058
rect -5324 -36806 -5224 -36058
rect -26392 -39962 -26292 -38042
rect -24286 -39962 -24186 -38042
rect -22214 -38080 -19978 -37980
rect -26392 -40062 -24186 -39962
rect -22154 -39980 -22054 -38080
rect -20078 -39980 -19978 -38080
rect -17986 -38036 -3080 -37936
rect -17986 -39928 -17886 -38036
rect -15882 -39928 -15782 -38036
rect -26392 -41954 -26292 -40062
rect -24286 -41954 -24186 -40062
rect -22917 -40080 -19196 -39980
rect -17986 -40028 -15782 -39928
rect -12934 -40006 -7304 -39906
rect -26392 -42054 -24186 -41954
rect -22154 -41980 -22054 -40080
rect -20078 -41980 -19978 -40080
rect -26392 -43954 -26292 -42054
rect -24286 -43954 -24186 -42054
rect -22917 -42080 -19196 -41980
rect -27129 -44054 -23408 -43954
rect -22154 -43980 -22054 -42080
rect -20078 -43980 -19978 -42080
rect -26392 -45954 -26292 -44054
rect -24286 -45954 -24186 -44054
rect -22917 -44080 -19196 -43980
rect -27129 -46054 -23408 -45954
rect -22154 -45980 -22054 -44080
rect -20078 -45980 -19978 -44080
rect -26392 -47954 -26292 -46054
rect -24286 -47954 -24186 -46054
rect -22917 -46080 -19196 -45980
rect -27129 -48054 -23408 -47954
rect -22154 -47980 -22054 -46080
rect -20078 -47980 -19978 -46080
rect -26392 -49954 -26292 -48054
rect -24286 -49954 -24186 -48054
rect -22917 -48080 -19196 -47980
rect -27129 -50054 -23408 -49954
rect -22154 -49980 -22054 -48080
rect -20078 -49980 -19978 -48080
rect -17986 -49922 -17886 -40028
rect -14318 -40769 -14218 -40574
rect -13736 -40648 -13636 -40574
rect -14323 -40796 -14213 -40769
rect -14323 -40852 -14296 -40796
rect -14240 -40852 -14213 -40796
rect -14323 -40879 -14213 -40852
rect -7404 -40874 -7304 -40006
rect -5340 -39968 -5240 -38036
rect -3180 -39968 -3080 -38036
rect -5340 -40068 -3080 -39968
rect -7404 -40930 -7382 -40874
rect -7326 -40930 -7304 -40874
rect -7404 -40952 -7304 -40930
rect -13180 -41116 -13048 -41088
rect -15860 -41146 -15760 -41124
rect -15860 -41202 -15838 -41146
rect -15782 -41202 -15760 -41146
rect -15860 -48874 -15760 -41202
rect -13180 -41172 -13146 -41116
rect -13090 -41172 -13048 -41116
rect -13180 -41472 -13048 -41172
rect -7978 -41116 -7878 -41094
rect -7978 -41172 -7956 -41116
rect -7900 -41172 -7878 -41116
rect -7978 -41466 -7878 -41172
rect -5315 -41168 -5205 -41141
rect -5315 -41224 -5288 -41168
rect -5232 -41224 -5205 -41168
rect -5315 -41251 -5205 -41224
rect -5310 -41484 -5210 -41251
rect -5310 -41570 -5206 -41484
rect -10842 -42024 -9436 -41924
rect -14632 -42486 -14060 -42464
rect -14632 -42542 -14610 -42486
rect -14554 -42542 -14060 -42486
rect -14632 -42564 -14060 -42542
rect -11648 -42858 -11548 -42180
rect -11648 -42914 -11626 -42858
rect -11570 -42914 -11548 -42858
rect -11648 -42936 -11548 -42914
rect -9536 -42858 -9436 -42024
rect -6634 -42554 -6332 -42532
rect -6634 -42610 -6410 -42554
rect -6354 -42610 -6332 -42554
rect -6634 -42632 -6332 -42610
rect -9536 -42914 -9514 -42858
rect -9458 -42914 -9436 -42858
rect -9536 -42936 -9436 -42914
rect -13751 -43142 -13641 -43115
rect -13751 -43198 -13724 -43142
rect -13668 -43198 -13641 -43142
rect -13751 -43225 -13641 -43198
rect -7447 -43134 -7337 -43107
rect -7447 -43190 -7420 -43134
rect -7364 -43190 -7337 -43134
rect -7447 -43217 -7337 -43190
rect -13746 -46858 -13646 -43225
rect -7442 -43426 -7342 -43217
rect -7444 -43498 -7342 -43426
rect -10922 -44854 -10822 -44592
rect -10922 -44910 -10900 -44854
rect -10844 -44910 -10822 -44854
rect -10922 -44932 -10822 -44910
rect -10169 -45146 -10059 -45119
rect -10169 -45202 -10142 -45146
rect -10086 -45202 -10059 -45146
rect -10169 -45229 -10059 -45202
rect -10164 -45450 -10064 -45229
rect -7444 -46753 -7344 -43498
rect -13746 -46914 -13724 -46858
rect -13668 -46914 -13646 -46858
rect -7449 -46780 -7339 -46753
rect -7449 -46836 -7422 -46780
rect -7366 -46836 -7339 -46780
rect -7449 -46863 -7339 -46836
rect -13746 -46936 -13646 -46914
rect -9542 -47126 -9442 -47104
rect -11649 -47156 -11539 -47129
rect -11649 -47212 -11622 -47156
rect -11566 -47212 -11539 -47156
rect -11649 -47239 -11539 -47212
rect -9542 -47182 -9520 -47126
rect -9464 -47182 -9442 -47126
rect -14654 -47428 -14296 -47406
rect -14654 -47446 -14274 -47428
rect -14654 -47502 -14610 -47446
rect -14554 -47502 -14274 -47446
rect -14654 -47528 -14274 -47502
rect -14654 -47554 -14296 -47528
rect -11644 -47550 -11544 -47239
rect -11648 -47554 -11544 -47550
rect -11648 -47914 -11548 -47554
rect -9542 -47914 -9442 -47182
rect -6652 -47524 -6320 -47516
rect -6982 -47552 -6320 -47524
rect -6982 -47608 -6410 -47552
rect -6354 -47608 -6320 -47552
rect -6982 -47624 -6320 -47608
rect -6652 -47648 -6320 -47624
rect -11648 -48014 -9442 -47914
rect -15860 -48930 -15838 -48874
rect -15782 -48930 -15760 -48874
rect -15860 -48952 -15760 -48930
rect -13004 -48872 -12904 -48584
rect -9542 -48662 -9442 -48014
rect -5306 -48498 -5206 -41570
rect -8052 -48658 -7952 -48568
rect -13004 -48928 -12982 -48872
rect -12926 -48928 -12904 -48872
rect -13004 -48950 -12904 -48928
rect -8074 -48872 -7938 -48658
rect -5312 -48773 -5212 -48580
rect -8074 -48928 -8038 -48872
rect -7982 -48928 -7938 -48872
rect -5317 -48800 -5207 -48773
rect -5317 -48856 -5290 -48800
rect -5234 -48856 -5207 -48800
rect -5317 -48883 -5207 -48856
rect -8074 -48966 -7938 -48928
rect -7436 -49068 -7336 -49046
rect -7436 -49124 -7414 -49068
rect -7358 -49124 -7336 -49068
rect -13761 -49170 -13651 -49143
rect -13761 -49226 -13734 -49170
rect -13678 -49226 -13651 -49170
rect -13761 -49253 -13651 -49226
rect -13756 -49572 -13656 -49253
rect -7436 -49906 -7336 -49124
rect -26392 -51954 -26292 -50054
rect -24286 -51954 -24186 -50054
rect -22917 -50080 -19196 -49980
rect -17986 -50022 -15768 -49922
rect -14493 -50006 -6560 -49906
rect -3180 -49940 -3080 -40068
rect -1110 -39950 -1010 -36058
rect 964 -37918 1064 -36034
rect 2355 -36050 6076 -36034
rect 3060 -37918 3160 -36050
rect 964 -37950 3162 -37918
rect 5228 -37950 5328 -36050
rect 964 -38018 6076 -37950
rect 2355 -38050 6076 -38018
rect 3060 -39950 3160 -38050
rect 5228 -39950 5328 -38050
rect -1110 -40050 1110 -39950
rect 2355 -40050 6076 -39950
rect -1110 -41946 -1010 -40050
rect 1010 -41946 1110 -40050
rect -1154 -42046 1110 -41946
rect 3060 -41950 3160 -40050
rect 5228 -41950 5328 -40050
rect 49186 -41108 52004 -41086
rect 49186 -41164 49208 -41108
rect 49264 -41164 51920 -41108
rect 51976 -41164 52004 -41108
rect 49186 -41186 52004 -41164
rect -1110 -43916 -1010 -42046
rect 1010 -43916 1110 -42046
rect 2355 -42050 6076 -41950
rect 52310 -41964 52510 -41908
rect 52310 -42020 52382 -41964
rect 52438 -42020 52510 -41964
rect -1110 -44016 1110 -43916
rect 3060 -43950 3160 -42050
rect 5228 -43950 5328 -42050
rect 26958 -42937 27090 -42924
rect 26958 -43001 26984 -42937
rect 27048 -43001 27090 -42937
rect 26958 -43018 27090 -43001
rect -1110 -45948 -1010 -44016
rect 1010 -45948 1110 -44016
rect 2355 -44050 6076 -43950
rect -1154 -46048 1110 -45948
rect 3060 -45950 3160 -44050
rect 5228 -45950 5328 -44050
rect -1110 -47944 -1010 -46048
rect 1010 -47944 1110 -46048
rect 2355 -46050 6076 -45950
rect -1130 -48044 1110 -47944
rect 3060 -47950 3160 -46050
rect 5228 -47950 5328 -46050
rect -27129 -51956 -23408 -51954
rect -27129 -52054 -22126 -51956
rect -26392 -53954 -26292 -52054
rect -24286 -52056 -22126 -52054
rect -24286 -53954 -24186 -52056
rect -22226 -53954 -22126 -52056
rect -27129 -54054 -22080 -53954
rect -26392 -55954 -26292 -54054
rect -24286 -55954 -24186 -54054
rect -22180 -55954 -22080 -54054
rect -20078 -53970 -19978 -50080
rect -17986 -51980 -17886 -50022
rect -15868 -51980 -15768 -50022
rect -5324 -50040 -3080 -49940
rect -5324 -51980 -5224 -50040
rect -17986 -52080 -3918 -51980
rect -3180 -52114 -3080 -50040
rect -1110 -49926 -1010 -48044
rect 1010 -49926 1110 -48044
rect 2355 -48050 6076 -47950
rect -1110 -50026 1110 -49926
rect 3060 -49950 3160 -48050
rect 5228 -49950 5328 -48050
rect -1110 -51970 -1010 -50026
rect 1010 -51970 1110 -50026
rect 2355 -50050 6076 -49950
rect 3060 -51950 3160 -50050
rect 5228 -51950 5328 -50050
rect -1110 -52070 1110 -51970
rect 2355 -52050 6076 -51950
rect 7906 -52004 14870 -51982
rect -17970 -53970 -17870 -53966
rect -15864 -53970 -15764 -53206
rect -13758 -53970 -13658 -53206
rect -11652 -53970 -11552 -53206
rect -9546 -53970 -9446 -53206
rect -7440 -53970 -7340 -53206
rect -1110 -53970 -1010 -52070
rect 3060 -53950 3160 -52050
rect 5228 -53950 5328 -52050
rect 7906 -52060 14792 -52004
rect 14848 -52060 14870 -52004
rect 7906 -52082 14870 -52060
rect 8165 -52948 8263 -52943
rect 8164 -52966 14862 -52948
rect 8164 -53030 8182 -52966
rect 8246 -52970 14862 -52966
rect 8246 -53026 14784 -52970
rect 14840 -53026 14862 -52970
rect 8246 -53030 14862 -53026
rect 8164 -53048 14862 -53030
rect 8165 -53053 8263 -53048
rect -20078 -54070 -1010 -53970
rect 1010 -54050 6076 -53950
rect 8138 -53964 14864 -53942
rect 8138 -54020 14786 -53964
rect 14842 -54020 14864 -53964
rect 8138 -54042 14864 -54020
rect -27129 -56054 -19912 -55954
rect -26392 -57954 -26292 -56054
rect -24286 -57930 -24186 -56054
rect -22156 -57930 -22056 -56054
rect -20012 -57206 -19912 -56054
rect -17970 -55976 -17870 -54070
rect -15864 -55976 -15764 -54070
rect -13758 -55976 -13658 -54070
rect -11652 -55976 -11552 -54070
rect -9546 -55976 -9446 -54070
rect -7440 -55976 -7340 -54070
rect -5340 -55976 -5240 -54070
rect 1010 -55950 1110 -54050
rect 3060 -55950 3160 -54050
rect 5228 -55950 5328 -54050
rect 8163 -54948 8261 -54943
rect 8162 -54966 14864 -54948
rect 8162 -55030 8180 -54966
rect 8244 -54970 14864 -54966
rect 8244 -55026 14786 -54970
rect 14842 -55026 14864 -54970
rect 8244 -55030 14864 -55026
rect 8162 -55048 14864 -55030
rect 8163 -55053 8261 -55048
rect -17970 -56076 -5240 -55976
rect -3278 -56050 5328 -55950
rect -15864 -56806 -15764 -56076
rect -13758 -56806 -13658 -56076
rect -11652 -56806 -11552 -56076
rect -9546 -56806 -9446 -56076
rect -7440 -56806 -7340 -56076
rect -3278 -57206 -3178 -56050
rect -1156 -57206 -1056 -56050
rect 1010 -57206 1110 -56050
rect -20060 -57930 -19912 -57206
rect -17954 -57930 -17854 -57206
rect -15848 -57930 -15748 -57206
rect -13742 -57930 -13642 -57206
rect -11636 -57930 -11536 -57206
rect -9530 -57930 -9430 -57206
rect -7424 -57930 -7324 -57206
rect -5318 -57930 -5218 -57206
rect -3278 -57930 -3112 -57206
rect -1156 -57930 -1006 -57206
rect 1000 -57930 1110 -57206
rect 3060 -57206 3160 -56050
rect 3060 -57930 3206 -57206
rect 5228 -57930 5328 -56050
rect 8100 -56356 14874 -56334
rect 8100 -56412 14796 -56356
rect 14852 -56412 14874 -56356
rect 8100 -56434 14874 -56412
rect 9350 -56729 9452 -56700
rect 9350 -56793 9372 -56729
rect 9436 -56793 9452 -56729
rect 9350 -56809 9452 -56793
rect 9350 -56873 9372 -56809
rect 9436 -56873 9452 -56809
rect 9350 -56889 9452 -56873
rect 9350 -56953 9372 -56889
rect 9436 -56953 9452 -56889
rect 9350 -56969 9452 -56953
rect 9350 -57033 9372 -56969
rect 9436 -57033 9452 -56969
rect 9350 -57049 9452 -57033
rect 9350 -57113 9372 -57049
rect 9436 -57113 9452 -57049
rect 9350 -57129 9452 -57113
rect 9350 -57193 9372 -57129
rect 9436 -57193 9452 -57129
rect 9350 -57209 9452 -57193
rect 9350 -57273 9372 -57209
rect 9436 -57273 9452 -57209
rect 9350 -57289 9452 -57273
rect 9350 -57353 9372 -57289
rect 9436 -57353 9452 -57289
rect 9350 -57369 9452 -57353
rect 9350 -57433 9372 -57369
rect 9436 -57433 9452 -57369
rect 9350 -57449 9452 -57433
rect 9350 -57513 9372 -57449
rect 9436 -57513 9452 -57449
rect 9350 -57536 9452 -57513
rect 12504 -57534 12604 -57512
rect 12504 -57590 12526 -57534
rect 12582 -57590 12604 -57534
rect 8086 -57637 10734 -57614
rect 8086 -57693 10654 -57637
rect 10710 -57693 10734 -57637
rect 8086 -57712 10734 -57693
rect 8086 -57714 10652 -57712
rect -24286 -57954 5328 -57930
rect -27129 -58030 5328 -57954
rect -27129 -58054 -23408 -58030
rect -26392 -59206 -26292 -58054
rect -26392 -60076 -26344 -59206
rect -24286 -59946 -24186 -58054
rect -22166 -58072 -22056 -58030
rect -20060 -58072 -19912 -58030
rect -22166 -59946 -22066 -58072
rect -20060 -59946 -19960 -58072
rect -17954 -59946 -17854 -58030
rect -15848 -59946 -15748 -58030
rect -13742 -59946 -13642 -58030
rect -11636 -59946 -11536 -58030
rect -9530 -59946 -9430 -58030
rect -7424 -59946 -7324 -58030
rect -5318 -59946 -5218 -58030
rect -3278 -58050 -3112 -58030
rect -3212 -59946 -3112 -58050
rect -1156 -58118 -1006 -58030
rect -1106 -59946 -1006 -58118
rect 1000 -58142 1110 -58030
rect 1000 -59946 1100 -58142
rect 3106 -59946 3206 -58030
rect 5228 -59946 5328 -58030
rect 12504 -58185 12604 -57590
rect 12504 -58241 12528 -58185
rect 12584 -58241 12604 -58185
rect 10276 -58429 12130 -58390
rect 10276 -58433 10330 -58429
rect 10394 -58433 10410 -58429
rect 10474 -58433 10490 -58429
rect 10554 -58433 10570 -58429
rect 10634 -58433 10650 -58429
rect 10714 -58433 10730 -58429
rect 10794 -58433 10810 -58429
rect 10874 -58433 10890 -58429
rect 10954 -58433 10970 -58429
rect 11034 -58433 11050 -58429
rect 11114 -58433 11130 -58429
rect 11194 -58433 11210 -58429
rect 11274 -58433 11290 -58429
rect 11354 -58433 11370 -58429
rect 11434 -58433 11450 -58429
rect 11514 -58433 11530 -58429
rect 11594 -58433 11610 -58429
rect 11674 -58433 11690 -58429
rect 11754 -58433 11770 -58429
rect 11834 -58433 11850 -58429
rect 11914 -58433 11930 -58429
rect 11994 -58433 12010 -58429
rect 12074 -58433 12130 -58429
rect 10276 -58489 10294 -58433
rect 12110 -58489 12130 -58433
rect 10276 -58493 10330 -58489
rect 10394 -58493 10410 -58489
rect 10474 -58493 10490 -58489
rect 10554 -58493 10570 -58489
rect 10634 -58493 10650 -58489
rect 10714 -58493 10730 -58489
rect 10794 -58493 10810 -58489
rect 10874 -58493 10890 -58489
rect 10954 -58493 10970 -58489
rect 11034 -58493 11050 -58489
rect 11114 -58493 11130 -58489
rect 11194 -58493 11210 -58489
rect 11274 -58493 11290 -58489
rect 11354 -58493 11370 -58489
rect 11434 -58493 11450 -58489
rect 11514 -58493 11530 -58489
rect 11594 -58493 11610 -58489
rect 11674 -58493 11690 -58489
rect 11754 -58493 11770 -58489
rect 11834 -58493 11850 -58489
rect 11914 -58493 11930 -58489
rect 11994 -58493 12010 -58489
rect 12074 -58493 12130 -58489
rect 10276 -58528 12130 -58493
rect -26244 -60046 5328 -59946
rect -24286 -60066 -24186 -60046
rect -22166 -60114 -22066 -60046
rect -20060 -60806 -19960 -60046
rect -17954 -60806 -17854 -60046
rect -15848 -60806 -15748 -60046
rect -13742 -60806 -13642 -60046
rect -11636 -60806 -11536 -60046
rect -9530 -60806 -9430 -60046
rect -7424 -60806 -7324 -60046
rect -5318 -60806 -5218 -60046
rect -3212 -60806 -3112 -60046
rect -1106 -60806 -1006 -60046
rect 1000 -60806 1100 -60046
rect 3106 -60806 3206 -60046
rect -25590 -62040 -24772 -61936
rect -9938 -63001 -9838 -63000
rect -14752 -63009 -14652 -63008
rect -16848 -63011 -16748 -63010
rect -18964 -63015 -18864 -63014
rect -18969 -63032 -18859 -63015
rect -18969 -63096 -18946 -63032
rect -18882 -63096 -18859 -63032
rect -18969 -63113 -18859 -63096
rect -16853 -63028 -16743 -63011
rect -16853 -63092 -16830 -63028
rect -16766 -63092 -16743 -63028
rect -16853 -63109 -16743 -63092
rect -14757 -63026 -14647 -63009
rect -10592 -63011 -10492 -63010
rect -12628 -63019 -12528 -63018
rect -14757 -63090 -14734 -63026
rect -14670 -63090 -14647 -63026
rect -14757 -63107 -14647 -63090
rect -12633 -63036 -12523 -63019
rect -12633 -63100 -12610 -63036
rect -12546 -63100 -12523 -63036
rect -25200 -63296 -25100 -63272
rect -25200 -63360 -25182 -63296
rect -25118 -63360 -25100 -63296
rect -18964 -63326 -18864 -63113
rect -16848 -63310 -16748 -63109
rect -25200 -65212 -25100 -63360
rect -25200 -65268 -25178 -65212
rect -25122 -65268 -25100 -65212
rect -25200 -65290 -25100 -65268
rect -21036 -63426 -18864 -63326
rect -17114 -63410 -16748 -63310
rect -21036 -65214 -20936 -63426
rect -21036 -65270 -21014 -65214
rect -20958 -65270 -20936 -65214
rect -21036 -65292 -20936 -65270
rect -17114 -65214 -17014 -63410
rect -14752 -63634 -14652 -63107
rect -12633 -63117 -12523 -63100
rect -10597 -63028 -10487 -63011
rect -10597 -63092 -10574 -63028
rect -10510 -63092 -10487 -63028
rect -10597 -63109 -10487 -63092
rect -9943 -63018 -9833 -63001
rect -9943 -63082 -9920 -63018
rect -9856 -63082 -9833 -63018
rect -8496 -63019 -8396 -63018
rect -9943 -63099 -9833 -63082
rect -8501 -63036 -8391 -63019
rect -7927 -63022 -7829 -63017
rect -17114 -65270 -17092 -65214
rect -17036 -65270 -17014 -65214
rect -17114 -65292 -17014 -65270
rect -16092 -63734 -14652 -63634
rect -16092 -65214 -15992 -63734
rect -12628 -64188 -12528 -63117
rect -10592 -64004 -10492 -63109
rect -9938 -63640 -9838 -63099
rect -8501 -63100 -8478 -63036
rect -8414 -63100 -8391 -63036
rect -8501 -63117 -8391 -63100
rect -7928 -63040 4110 -63022
rect -7928 -63104 -7910 -63040
rect -7846 -63104 4110 -63040
rect -8496 -63322 -8396 -63117
rect -7928 -63122 4110 -63104
rect -7927 -63127 -7829 -63122
rect -8496 -63422 56 -63322
rect -9938 -63740 -4002 -63640
rect -10592 -64028 -9114 -64004
rect -10592 -64084 -9196 -64028
rect -9140 -64084 -9114 -64028
rect -10592 -64104 -9114 -64084
rect -12628 -64288 -7874 -64188
rect -16092 -65270 -16070 -65214
rect -16014 -65270 -15992 -65214
rect -16092 -65292 -15992 -65270
rect -7974 -65216 -7874 -64288
rect -7974 -65272 -7954 -65216
rect -7898 -65272 -7874 -65216
rect -7974 -65298 -7874 -65272
rect -4102 -65214 -4002 -63740
rect -4102 -65270 -4080 -65214
rect -4024 -65270 -4002 -65214
rect -4102 -65292 -4002 -65270
rect -44 -65218 56 -63422
rect -44 -65274 -22 -65218
rect 34 -65274 56 -65218
rect -44 -65296 56 -65274
rect 4010 -65216 4110 -63122
rect 4010 -65272 4032 -65216
rect 4088 -65272 4110 -65216
rect 4010 -65294 4110 -65272
rect 12504 -65426 12604 -58241
rect 52310 -59666 52510 -42020
rect 53309 -42484 53379 -42477
rect 53309 -42540 53316 -42484
rect 53372 -42540 53379 -42484
rect 53309 -42547 53379 -42540
rect -26472 -65448 12604 -65426
rect -26472 -65504 -26446 -65448
rect -26390 -65504 -22446 -65448
rect -22390 -65504 -18448 -65448
rect -18392 -65504 -14448 -65448
rect -14392 -65504 -10448 -65448
rect -10392 -65504 -6446 -65448
rect -6390 -65504 -2450 -65448
rect -2394 -65504 1554 -65448
rect 1610 -65504 5556 -65448
rect 5612 -65504 12604 -65448
rect -26472 -65526 12604 -65504
rect 12962 -59716 52510 -59666
rect 12962 -59772 13018 -59716
rect 13074 -59772 52510 -59716
rect 12962 -59866 52510 -59772
rect -28296 -67922 5506 -67902
rect -28296 -67978 -26576 -67922
rect -26520 -67978 -22576 -67922
rect -22520 -67978 -18576 -67922
rect -18520 -67978 -14576 -67922
rect -14520 -67978 -10576 -67922
rect -10520 -67978 -6576 -67922
rect -6520 -67978 -2576 -67922
rect -2520 -67978 1424 -67922
rect 1480 -67924 5506 -67922
rect 1480 -67978 5424 -67924
rect -28296 -67980 5424 -67978
rect 5480 -67980 5506 -67924
rect -28296 -68002 5506 -67980
rect -25254 -68954 -25154 -68924
rect -25254 -69010 -25230 -68954
rect -25174 -69010 -25154 -68954
rect -25254 -72108 -25154 -69010
rect -25254 -72164 -25236 -72108
rect -25180 -72164 -25154 -72108
rect -25254 -72192 -25154 -72164
rect -21254 -68954 -21154 -68924
rect -21254 -69010 -21230 -68954
rect -21174 -69010 -21154 -68954
rect -21254 -72108 -21154 -69010
rect -21254 -72164 -21236 -72108
rect -21180 -72164 -21154 -72108
rect -21254 -72192 -21154 -72164
rect -17254 -68954 -17154 -68924
rect -17254 -69010 -17230 -68954
rect -17174 -69010 -17154 -68954
rect -17254 -72108 -17154 -69010
rect -17254 -72164 -17236 -72108
rect -17180 -72164 -17154 -72108
rect -17254 -72192 -17154 -72164
rect -13254 -68954 -13154 -68924
rect -13254 -69010 -13230 -68954
rect -13174 -69010 -13154 -68954
rect -13254 -72108 -13154 -69010
rect -13254 -72164 -13236 -72108
rect -13180 -72164 -13154 -72108
rect -13254 -72192 -13154 -72164
rect -9254 -68954 -9154 -68924
rect -9254 -69010 -9230 -68954
rect -9174 -69010 -9154 -68954
rect -9254 -72108 -9154 -69010
rect -9254 -72164 -9236 -72108
rect -9180 -72164 -9154 -72108
rect -9254 -72192 -9154 -72164
rect -5254 -68954 -5154 -68924
rect -5254 -69010 -5230 -68954
rect -5174 -69010 -5154 -68954
rect -5254 -72108 -5154 -69010
rect -5254 -72164 -5236 -72108
rect -5180 -72164 -5154 -72108
rect -5254 -72192 -5154 -72164
rect -1254 -68954 -1154 -68924
rect -1254 -69010 -1230 -68954
rect -1174 -69010 -1154 -68954
rect -1254 -72108 -1154 -69010
rect -1254 -72164 -1236 -72108
rect -1180 -72164 -1154 -72108
rect -1254 -72192 -1154 -72164
rect 2746 -68954 2846 -68924
rect 2746 -69010 2770 -68954
rect 2826 -69010 2846 -68954
rect 2746 -72108 2846 -69010
rect 2746 -72164 2764 -72108
rect 2820 -72164 2846 -72108
rect 2746 -72192 2846 -72164
rect 6746 -68954 6846 -68924
rect 6746 -69010 6770 -68954
rect 6826 -69010 6846 -68954
rect 6746 -72108 6846 -69010
rect 6746 -72164 6764 -72108
rect 6820 -72164 6846 -72108
rect 6746 -72192 6846 -72164
rect 12962 -72808 13162 -59866
rect 4844 -72864 13162 -72808
rect -28500 -72882 13162 -72864
rect -28500 -72884 -11092 -72882
rect -28500 -72940 -27092 -72884
rect -27036 -72940 -23092 -72884
rect -23036 -72940 -19092 -72884
rect -19036 -72940 -15092 -72884
rect -15036 -72938 -11092 -72884
rect -11036 -72884 13162 -72882
rect -11036 -72938 -7092 -72884
rect -15036 -72940 -7092 -72938
rect -7036 -72940 -3092 -72884
rect -3036 -72940 908 -72884
rect 964 -72940 4908 -72884
rect 4964 -72940 13162 -72884
rect -28500 -72964 13162 -72940
rect 4844 -73008 13162 -72964
rect -28238 -74868 4986 -74848
rect -28238 -74870 4910 -74868
rect -28238 -74872 -23090 -74870
rect -28238 -74928 -27090 -74872
rect -27034 -74926 -23090 -74872
rect -23034 -74926 -19090 -74870
rect -19034 -74926 -15090 -74870
rect -15034 -74872 -3090 -74870
rect -15034 -74926 -11090 -74872
rect -27034 -74928 -11090 -74926
rect -11034 -74928 -7090 -74872
rect -7034 -74926 -3090 -74872
rect -3034 -74926 910 -74870
rect 966 -74924 4910 -74870
rect 4966 -74924 4986 -74868
rect 966 -74926 4986 -74924
rect -7034 -74928 4986 -74926
rect -28238 -74948 4986 -74928
<< via3 >>
rect 26984 -42944 27048 -42937
rect 26984 -43000 26988 -42944
rect 26988 -43000 27044 -42944
rect 27044 -43000 27048 -42944
rect 26984 -43001 27048 -43000
rect 8182 -53030 8246 -52966
rect 8180 -55030 8244 -54966
rect 9372 -56733 9436 -56729
rect 9372 -56789 9376 -56733
rect 9376 -56789 9432 -56733
rect 9432 -56789 9436 -56733
rect 9372 -56793 9436 -56789
rect 9372 -56813 9436 -56809
rect 9372 -56869 9376 -56813
rect 9376 -56869 9432 -56813
rect 9432 -56869 9436 -56813
rect 9372 -56873 9436 -56869
rect 9372 -56893 9436 -56889
rect 9372 -56949 9376 -56893
rect 9376 -56949 9432 -56893
rect 9432 -56949 9436 -56893
rect 9372 -56953 9436 -56949
rect 9372 -56973 9436 -56969
rect 9372 -57029 9376 -56973
rect 9376 -57029 9432 -56973
rect 9432 -57029 9436 -56973
rect 9372 -57033 9436 -57029
rect 9372 -57053 9436 -57049
rect 9372 -57109 9376 -57053
rect 9376 -57109 9432 -57053
rect 9432 -57109 9436 -57053
rect 9372 -57113 9436 -57109
rect 9372 -57133 9436 -57129
rect 9372 -57189 9376 -57133
rect 9376 -57189 9432 -57133
rect 9432 -57189 9436 -57133
rect 9372 -57193 9436 -57189
rect 9372 -57213 9436 -57209
rect 9372 -57269 9376 -57213
rect 9376 -57269 9432 -57213
rect 9432 -57269 9436 -57213
rect 9372 -57273 9436 -57269
rect 9372 -57293 9436 -57289
rect 9372 -57349 9376 -57293
rect 9376 -57349 9432 -57293
rect 9432 -57349 9436 -57293
rect 9372 -57353 9436 -57349
rect 9372 -57373 9436 -57369
rect 9372 -57429 9376 -57373
rect 9376 -57429 9432 -57373
rect 9432 -57429 9436 -57373
rect 9372 -57433 9436 -57429
rect 9372 -57453 9436 -57449
rect 9372 -57509 9376 -57453
rect 9376 -57509 9432 -57453
rect 9432 -57509 9436 -57453
rect 9372 -57513 9436 -57509
rect 10330 -58433 10394 -58429
rect 10410 -58433 10474 -58429
rect 10490 -58433 10554 -58429
rect 10570 -58433 10634 -58429
rect 10650 -58433 10714 -58429
rect 10730 -58433 10794 -58429
rect 10810 -58433 10874 -58429
rect 10890 -58433 10954 -58429
rect 10970 -58433 11034 -58429
rect 11050 -58433 11114 -58429
rect 11130 -58433 11194 -58429
rect 11210 -58433 11274 -58429
rect 11290 -58433 11354 -58429
rect 11370 -58433 11434 -58429
rect 11450 -58433 11514 -58429
rect 11530 -58433 11594 -58429
rect 11610 -58433 11674 -58429
rect 11690 -58433 11754 -58429
rect 11770 -58433 11834 -58429
rect 11850 -58433 11914 -58429
rect 11930 -58433 11994 -58429
rect 12010 -58433 12074 -58429
rect 10330 -58489 10350 -58433
rect 10350 -58489 10374 -58433
rect 10374 -58489 10394 -58433
rect 10410 -58489 10430 -58433
rect 10430 -58489 10454 -58433
rect 10454 -58489 10474 -58433
rect 10490 -58489 10510 -58433
rect 10510 -58489 10534 -58433
rect 10534 -58489 10554 -58433
rect 10570 -58489 10590 -58433
rect 10590 -58489 10614 -58433
rect 10614 -58489 10634 -58433
rect 10650 -58489 10670 -58433
rect 10670 -58489 10694 -58433
rect 10694 -58489 10714 -58433
rect 10730 -58489 10750 -58433
rect 10750 -58489 10774 -58433
rect 10774 -58489 10794 -58433
rect 10810 -58489 10830 -58433
rect 10830 -58489 10854 -58433
rect 10854 -58489 10874 -58433
rect 10890 -58489 10910 -58433
rect 10910 -58489 10934 -58433
rect 10934 -58489 10954 -58433
rect 10970 -58489 10990 -58433
rect 10990 -58489 11014 -58433
rect 11014 -58489 11034 -58433
rect 11050 -58489 11070 -58433
rect 11070 -58489 11094 -58433
rect 11094 -58489 11114 -58433
rect 11130 -58489 11150 -58433
rect 11150 -58489 11174 -58433
rect 11174 -58489 11194 -58433
rect 11210 -58489 11230 -58433
rect 11230 -58489 11254 -58433
rect 11254 -58489 11274 -58433
rect 11290 -58489 11310 -58433
rect 11310 -58489 11334 -58433
rect 11334 -58489 11354 -58433
rect 11370 -58489 11390 -58433
rect 11390 -58489 11414 -58433
rect 11414 -58489 11434 -58433
rect 11450 -58489 11470 -58433
rect 11470 -58489 11494 -58433
rect 11494 -58489 11514 -58433
rect 11530 -58489 11550 -58433
rect 11550 -58489 11574 -58433
rect 11574 -58489 11594 -58433
rect 11610 -58489 11630 -58433
rect 11630 -58489 11654 -58433
rect 11654 -58489 11674 -58433
rect 11690 -58489 11710 -58433
rect 11710 -58489 11734 -58433
rect 11734 -58489 11754 -58433
rect 11770 -58489 11790 -58433
rect 11790 -58489 11814 -58433
rect 11814 -58489 11834 -58433
rect 11850 -58489 11870 -58433
rect 11870 -58489 11894 -58433
rect 11894 -58489 11914 -58433
rect 11930 -58489 11950 -58433
rect 11950 -58489 11974 -58433
rect 11974 -58489 11994 -58433
rect 12010 -58489 12030 -58433
rect 12030 -58489 12054 -58433
rect 12054 -58489 12074 -58433
rect 10330 -58493 10394 -58489
rect 10410 -58493 10474 -58489
rect 10490 -58493 10554 -58489
rect 10570 -58493 10634 -58489
rect 10650 -58493 10714 -58489
rect 10730 -58493 10794 -58489
rect 10810 -58493 10874 -58489
rect 10890 -58493 10954 -58489
rect 10970 -58493 11034 -58489
rect 11050 -58493 11114 -58489
rect 11130 -58493 11194 -58489
rect 11210 -58493 11274 -58489
rect 11290 -58493 11354 -58489
rect 11370 -58493 11434 -58489
rect 11450 -58493 11514 -58489
rect 11530 -58493 11594 -58489
rect 11610 -58493 11674 -58489
rect 11690 -58493 11754 -58489
rect 11770 -58493 11834 -58489
rect 11850 -58493 11914 -58489
rect 11930 -58493 11994 -58489
rect 12010 -58493 12074 -58489
rect -18946 -63096 -18882 -63032
rect -16830 -63092 -16766 -63028
rect -14734 -63090 -14670 -63026
rect -12610 -63100 -12546 -63036
rect -25182 -63360 -25118 -63296
rect -10574 -63092 -10510 -63028
rect -9920 -63082 -9856 -63018
rect -8478 -63100 -8414 -63036
rect -7910 -63104 -7846 -63040
<< metal4 >>
rect 8788 -27700 11212 -27578
rect 7330 -27958 8260 -27942
rect -28478 -28058 8276 -27958
rect -28470 -28948 -28370 -28058
rect -27640 -28948 -27540 -28058
rect -26348 -28948 -26248 -28058
rect -24242 -28948 -24142 -28058
rect -22136 -28948 -22036 -28058
rect -20030 -28948 -19930 -28058
rect -17924 -28948 -17824 -28058
rect -15818 -28948 -15718 -28058
rect -13712 -28948 -13612 -28058
rect -11606 -28948 -11506 -28058
rect -9500 -28948 -9400 -28058
rect -7394 -28948 -7294 -28058
rect -5288 -28948 -5188 -28058
rect -3182 -28948 -3082 -28058
rect -1076 -28948 -976 -28058
rect 1030 -28948 1130 -28058
rect 3136 -28948 3236 -28058
rect 5242 -28948 5342 -28058
rect 7368 -28948 7468 -28058
rect 8160 -28948 8260 -28058
rect 8788 -28256 8910 -27700
rect 9466 -28256 11212 -27700
rect 8788 -28378 11212 -28256
rect 48760 -27700 51352 -27578
rect 48760 -28256 50674 -27700
rect 51230 -28256 51352 -27700
rect 48760 -28378 51352 -28256
rect -28470 -29048 8260 -28948
rect -28470 -29938 -28370 -29048
rect -27640 -29938 -27540 -29048
rect -28470 -30038 -27540 -29938
rect -28470 -30948 -28370 -30038
rect -27640 -30948 -27540 -30038
rect -26348 -30948 -26248 -29048
rect -24242 -30948 -24142 -29048
rect -22136 -30948 -22036 -29048
rect -20030 -30948 -19930 -29048
rect -17924 -30948 -17824 -29048
rect -15818 -30948 -15718 -29048
rect -13712 -30948 -13612 -29048
rect -11606 -30948 -11506 -29048
rect -9500 -30948 -9400 -29048
rect -7394 -30948 -7294 -29048
rect -5288 -30948 -5188 -29048
rect -3182 -30948 -3082 -29048
rect -1076 -30948 -976 -29048
rect 1030 -30948 1130 -29048
rect 3136 -30948 3236 -29048
rect 5242 -30948 5342 -29048
rect 7368 -29942 7468 -29048
rect 8160 -29942 8260 -29048
rect 7330 -30042 8260 -29942
rect 7368 -30948 7468 -30042
rect 8160 -30948 8260 -30042
rect -28470 -31048 8260 -30948
rect -28470 -31938 -28370 -31048
rect -27640 -31938 -27540 -31048
rect -28470 -32038 -27540 -31938
rect -28470 -32948 -28370 -32038
rect -27640 -32948 -27540 -32038
rect -26348 -32948 -26248 -31048
rect -24242 -32948 -24142 -31048
rect -22136 -32948 -22036 -31048
rect -20030 -32948 -19930 -31048
rect -17924 -32948 -17824 -31048
rect -15818 -32948 -15718 -31048
rect -13712 -32948 -13612 -31048
rect -11606 -32948 -11506 -31048
rect -9500 -32948 -9400 -31048
rect -7394 -32948 -7294 -31048
rect -5288 -32948 -5188 -31048
rect -3182 -32948 -3082 -31048
rect -1076 -32948 -976 -31048
rect 1030 -32948 1130 -31048
rect 3136 -32948 3236 -31048
rect 5242 -32948 5342 -31048
rect 7368 -31942 7468 -31048
rect 8160 -31942 8260 -31048
rect 7330 -32042 8260 -31942
rect 7368 -32948 7468 -32042
rect 8160 -32948 8260 -32042
rect -28470 -33048 8260 -32948
rect -28470 -33938 -28370 -33048
rect -27640 -33938 -27540 -33048
rect -28470 -34038 -27540 -33938
rect -28470 -34948 -28370 -34038
rect -27640 -34948 -27540 -34038
rect -26348 -34948 -26248 -33048
rect -24242 -34948 -24142 -33048
rect -22136 -34948 -22036 -33048
rect -20030 -34948 -19930 -33048
rect -17924 -34948 -17824 -33048
rect -15818 -34948 -15718 -33048
rect -13712 -34948 -13612 -33048
rect -11606 -34948 -11506 -33048
rect -9500 -34948 -9400 -33048
rect -7394 -34948 -7294 -33048
rect -5288 -34948 -5188 -33048
rect -3182 -34948 -3082 -33048
rect -1076 -34948 -976 -33048
rect 1030 -34948 1130 -33048
rect 3136 -34948 3236 -33048
rect 5242 -34948 5342 -33048
rect 7368 -33942 7468 -33048
rect 8160 -33942 8260 -33048
rect 7330 -34042 8260 -33942
rect 7368 -34948 7468 -34042
rect 8160 -34948 8260 -34042
rect -28470 -35048 8260 -34948
rect -28470 -35938 -28370 -35048
rect -27640 -35938 -27540 -35048
rect -28470 -36038 -27540 -35938
rect -28470 -36948 -28370 -36038
rect -27640 -36948 -27540 -36038
rect -26348 -36948 -26248 -35048
rect -24242 -36948 -24142 -35048
rect -22136 -36948 -22036 -35048
rect -20030 -36948 -19930 -35048
rect -17924 -36948 -17824 -35048
rect -15818 -36948 -15718 -35048
rect -13712 -36948 -13612 -35048
rect -11606 -36948 -11506 -35048
rect -9500 -36948 -9400 -35048
rect -7394 -36948 -7294 -35048
rect -5288 -36948 -5188 -35048
rect -3182 -36948 -3082 -35048
rect -1076 -36948 -976 -35048
rect 1030 -36948 1130 -35048
rect 3136 -36948 3236 -35048
rect 5242 -36948 5342 -35048
rect 7368 -35942 7468 -35048
rect 8160 -35942 8260 -35048
rect 7330 -36042 8260 -35942
rect 7368 -36948 7468 -36042
rect 8160 -36948 8260 -36042
rect -28470 -37048 8260 -36948
rect -28470 -37938 -28370 -37048
rect -27640 -37938 -27540 -37048
rect -28470 -38038 -27540 -37938
rect -28470 -38948 -28370 -38038
rect -27640 -38948 -27540 -38038
rect -26348 -38948 -26248 -37048
rect -24242 -38948 -24142 -37048
rect -22136 -38948 -22036 -37048
rect -20030 -38948 -19930 -37048
rect -17924 -38948 -17824 -37048
rect -15818 -38948 -15718 -37048
rect -13712 -38948 -13612 -37048
rect -11606 -38948 -11506 -37048
rect -9500 -38948 -9400 -37048
rect -7394 -38948 -7294 -37048
rect -5288 -38948 -5188 -37048
rect -3182 -38948 -3082 -37048
rect -1076 -38948 -976 -37048
rect 1030 -38948 1130 -37048
rect 3136 -38948 3236 -37048
rect 5242 -38948 5342 -37048
rect 7368 -37942 7468 -37048
rect 8160 -37942 8260 -37048
rect 7330 -38042 8260 -37942
rect 7368 -38948 7468 -38042
rect 8160 -38948 8260 -38042
rect -28470 -39048 8260 -38948
rect -28470 -39938 -28370 -39048
rect -27640 -39938 -27540 -39048
rect -28470 -40038 -27540 -39938
rect -28470 -40948 -28370 -40038
rect -27640 -40948 -27540 -40038
rect -26348 -40948 -26248 -39048
rect -24242 -40948 -24142 -39048
rect -22136 -40948 -22036 -39048
rect -20030 -40948 -19930 -39048
rect -17924 -40948 -17824 -39048
rect -15818 -40948 -15718 -39048
rect -13712 -40948 -13612 -39048
rect -11606 -40948 -11506 -39048
rect -9500 -40948 -9400 -39048
rect -7394 -40948 -7294 -39048
rect -5288 -40948 -5188 -39048
rect -3182 -40948 -3082 -39048
rect -1076 -40948 -976 -39048
rect 1030 -40948 1130 -39048
rect 3136 -40948 3236 -39048
rect 5242 -40948 5342 -39048
rect 7368 -39942 7468 -39048
rect 8160 -39942 8260 -39048
rect 50552 -38802 52664 -38680
rect 50552 -39358 50674 -38802
rect 51230 -39358 52664 -38802
rect 50552 -39480 52664 -39358
rect 7330 -40042 8260 -39942
rect 7368 -40948 7468 -40042
rect 8160 -40948 8260 -40042
rect -28470 -41048 8260 -40948
rect -28470 -41938 -28370 -41048
rect -27640 -41938 -27540 -41048
rect -28470 -42038 -27540 -41938
rect -28470 -42948 -28370 -42038
rect -27640 -42948 -27540 -42038
rect -26348 -42948 -26248 -41048
rect -24242 -42948 -24142 -41048
rect -22136 -42948 -22036 -41048
rect -20030 -42948 -19930 -41048
rect -17924 -42948 -17824 -41048
rect -15818 -42948 -15718 -41048
rect -13712 -42948 -13612 -41048
rect -11606 -42948 -11506 -41048
rect -9500 -42948 -9400 -41048
rect -7394 -42948 -7294 -41048
rect -5288 -42948 -5188 -41048
rect -3182 -42948 -3082 -41048
rect -1076 -42948 -976 -41048
rect 1030 -42948 1130 -41048
rect 3136 -42948 3236 -41048
rect 5242 -42948 5342 -41048
rect 7368 -41942 7468 -41048
rect 8160 -41942 8260 -41048
rect 7330 -42042 8260 -41942
rect 7368 -42948 7468 -42042
rect 8160 -42948 8260 -42042
rect -28470 -43048 8260 -42948
rect 26980 -42937 27052 -42936
rect 26980 -43001 26984 -42937
rect 27048 -43001 27052 -42937
rect 26980 -43002 27052 -43001
rect -28470 -43938 -28370 -43048
rect -27640 -43938 -27540 -43048
rect -28470 -44038 -27540 -43938
rect -28470 -44942 -28370 -44038
rect -27640 -44942 -27540 -44038
rect -26348 -44942 -26248 -43048
rect -24242 -44942 -24142 -43048
rect -22136 -44942 -22036 -43048
rect -20030 -44942 -19930 -43048
rect -17924 -44942 -17824 -43048
rect -15818 -44942 -15718 -43048
rect -13712 -44942 -13612 -43410
rect -11606 -44942 -11506 -43048
rect -9500 -44942 -9400 -43048
rect -28470 -45042 -9400 -44942
rect -8684 -44864 -8584 -44560
rect -8684 -44964 -8182 -44864
rect -7394 -44948 -7294 -43426
rect -5288 -44948 -5188 -43048
rect -3182 -44948 -3082 -43048
rect -1076 -44948 -976 -43048
rect 1030 -44948 1130 -43048
rect 3136 -44948 3236 -43048
rect 5242 -44948 5342 -43048
rect 7368 -43942 7468 -43048
rect 8160 -43942 8260 -43048
rect 7330 -44042 8260 -43942
rect 50544 -43306 53126 -43184
rect 50544 -43862 50666 -43306
rect 51222 -43862 53126 -43306
rect 50544 -43984 53126 -43862
rect 7368 -44948 7468 -44042
rect 8160 -44948 8260 -44042
rect -28470 -45938 -28370 -45042
rect -27640 -45938 -27540 -45042
rect -28470 -46038 -27540 -45938
rect -28470 -46950 -28370 -46038
rect -27640 -46950 -27540 -46038
rect -26348 -46950 -26248 -45042
rect -24242 -46950 -24142 -45042
rect -22136 -46950 -22036 -45042
rect -20030 -46950 -19930 -45042
rect -17924 -46950 -17824 -45042
rect -15818 -46950 -15718 -45042
rect -13712 -46950 -13612 -45042
rect -11606 -46950 -11506 -45042
rect -28470 -47050 -11506 -46950
rect -10794 -46922 -10694 -46420
rect -10794 -47022 -10292 -46922
rect -28470 -47938 -28370 -47050
rect -27640 -47938 -27540 -47050
rect -28470 -48038 -27540 -47938
rect -28470 -48952 -28370 -48038
rect -27640 -48952 -27540 -48038
rect -26348 -48952 -26248 -47050
rect -24242 -48952 -24142 -47050
rect -22136 -48952 -22036 -47050
rect -20030 -48952 -19930 -47050
rect -17924 -48952 -17824 -47050
rect -15818 -48952 -15718 -47050
rect -28470 -49052 -15718 -48952
rect -15000 -48900 -14900 -48486
rect -15000 -49000 -14652 -48900
rect -28470 -49938 -28370 -49052
rect -27640 -49938 -27540 -49052
rect -28470 -50038 -27540 -49938
rect -28470 -50966 -28370 -50038
rect -27640 -50966 -27540 -50038
rect -26348 -50966 -26248 -49052
rect -24242 -50966 -24142 -49052
rect -22136 -50966 -22036 -49052
rect -20030 -50966 -19930 -49052
rect -17924 -50966 -17824 -49052
rect -15818 -50966 -15718 -49052
rect -28470 -51066 -15718 -50966
rect -28470 -51938 -28370 -51066
rect -27640 -51938 -27540 -51066
rect -28470 -52038 -27540 -51938
rect -28470 -52962 -28370 -52038
rect -27640 -52962 -27540 -52038
rect -26348 -52962 -26248 -51066
rect -24242 -52962 -24142 -51066
rect -22136 -52962 -22036 -51066
rect -20030 -52962 -19930 -51066
rect -17924 -52962 -17824 -51066
rect -28470 -53062 -17824 -52962
rect -28470 -53938 -28370 -53062
rect -27640 -53938 -27540 -53062
rect -28470 -54038 -27540 -53938
rect -28470 -54956 -28370 -54038
rect -27640 -54956 -27540 -54038
rect -26348 -54956 -26248 -53062
rect -24242 -54956 -24142 -53062
rect -22136 -54956 -22036 -53062
rect -20030 -54956 -19930 -53062
rect -28470 -55056 -19930 -54956
rect -19212 -54926 -19112 -54450
rect -19212 -55026 -18864 -54926
rect -28470 -55938 -28370 -55056
rect -27640 -55938 -27540 -55056
rect -28470 -56038 -27540 -55938
rect -28470 -56966 -28370 -56038
rect -27640 -56966 -27540 -56038
rect -26348 -56966 -26248 -55056
rect -24242 -56966 -24142 -55056
rect -22136 -56966 -22036 -55056
rect -20030 -56966 -19930 -55056
rect -28470 -57066 -19930 -56966
rect -28470 -57938 -28370 -57066
rect -27640 -57938 -27540 -57066
rect -28470 -58038 -27540 -57938
rect -28470 -58934 -28370 -58038
rect -27640 -58934 -27540 -58038
rect -26348 -58934 -26248 -57066
rect -24242 -58934 -24142 -57066
rect -22136 -58934 -22036 -57066
rect -20030 -58934 -19930 -57066
rect -28470 -59034 -19930 -58934
rect -28470 -59938 -28370 -59034
rect -27640 -59938 -27540 -59034
rect -28470 -60038 -27540 -59938
rect -28470 -60942 -28370 -60038
rect -27640 -60942 -27540 -60038
rect -26348 -60942 -26248 -59034
rect -28470 -61042 -26248 -60942
rect -25530 -60938 -25434 -60554
rect -25530 -61034 -25104 -60938
rect -28470 -61936 -28370 -61042
rect -27640 -61936 -27540 -61042
rect -26348 -61936 -26248 -61042
rect -28470 -62036 -25436 -61936
rect -25200 -63050 -25104 -61034
rect -24242 -60942 -24142 -59034
rect -22136 -60942 -22036 -59034
rect -20030 -60942 -19930 -59034
rect -24242 -61042 -19930 -60942
rect -24242 -61930 -24142 -61042
rect -22136 -61908 -22036 -61042
rect -20030 -61908 -19930 -61042
rect -24242 -61936 -23350 -61930
rect -22136 -61936 -21244 -61930
rect -20030 -61936 -19138 -61930
rect -24884 -62030 -19138 -61936
rect -24884 -62036 -19570 -62030
rect -18964 -63032 -18864 -55026
rect -17924 -61908 -17824 -53062
rect -17114 -52968 -17014 -52416
rect -17114 -53068 -16748 -52968
rect -17924 -62030 -17032 -61930
rect -25200 -63277 -25100 -63050
rect -18964 -63096 -18946 -63032
rect -18882 -63096 -18864 -63032
rect -18964 -63114 -18864 -63096
rect -16848 -63028 -16748 -53068
rect -15818 -61908 -15718 -51066
rect -15818 -62030 -14926 -61930
rect -16848 -63092 -16830 -63028
rect -16766 -63092 -16748 -63028
rect -16848 -63110 -16748 -63092
rect -14752 -63026 -14652 -49000
rect -13712 -61908 -13612 -47050
rect -12906 -48898 -12806 -48394
rect -12906 -48998 -12528 -48898
rect -13712 -62030 -12820 -61930
rect -14752 -63090 -14734 -63026
rect -14670 -63090 -14652 -63026
rect -14752 -63108 -14652 -63090
rect -12628 -63036 -12528 -48998
rect -11606 -61908 -11506 -47050
rect -10794 -48956 -10694 -48326
rect -10794 -49056 -10492 -48956
rect -11606 -62030 -10714 -61930
rect -12628 -63100 -12610 -63036
rect -12546 -63100 -12528 -63036
rect -12628 -63118 -12528 -63100
rect -10592 -63028 -10492 -49056
rect -10592 -63092 -10574 -63028
rect -10510 -63092 -10492 -63028
rect -10592 -63110 -10492 -63092
rect -10392 -63000 -10292 -47022
rect -9500 -61908 -9400 -45042
rect -8688 -47012 -8588 -46382
rect -8688 -47112 -8396 -47012
rect -9500 -62030 -8608 -61930
rect -10392 -63018 -9838 -63000
rect -10392 -63082 -9920 -63018
rect -9856 -63082 -9838 -63018
rect -10392 -63100 -9838 -63082
rect -8496 -63036 -8396 -47112
rect -8496 -63100 -8478 -63036
rect -8414 -63100 -8396 -63036
rect -8496 -63118 -8396 -63100
rect -8282 -63022 -8182 -44964
rect -7408 -45048 8260 -44948
rect -7394 -46948 -7294 -45048
rect -5288 -46948 -5188 -45048
rect -3182 -46948 -3082 -45048
rect -1076 -46948 -976 -45048
rect 1030 -46948 1130 -45048
rect 3136 -46948 3236 -45048
rect 5242 -46948 5342 -45048
rect 7368 -45942 7468 -45048
rect 8160 -45942 8260 -45048
rect 7330 -46042 8260 -45942
rect 7368 -46948 7468 -46042
rect 8160 -46948 8260 -46042
rect -7394 -47048 8260 -46948
rect -7394 -48948 -7294 -47048
rect -5288 -48948 -5188 -47048
rect -3182 -48948 -3082 -47048
rect -1076 -48948 -976 -47048
rect 1030 -48948 1130 -47048
rect 3136 -48948 3236 -47048
rect 5242 -48948 5342 -47048
rect 7368 -47942 7468 -47048
rect 8160 -47942 8260 -47048
rect 7330 -48042 8260 -47942
rect 7368 -48948 7468 -48042
rect 8160 -48948 8260 -48042
rect -7394 -49048 8260 -48948
rect -7394 -61908 -7294 -49048
rect -5288 -50948 -5188 -49048
rect -3182 -50948 -3082 -49048
rect -1076 -50948 -976 -49048
rect 1030 -50948 1130 -49048
rect 3136 -50948 3236 -49048
rect 5242 -50948 5342 -49048
rect 7368 -49942 7468 -49048
rect 8160 -49942 8260 -49048
rect 7330 -50042 8260 -49942
rect 7368 -50948 7468 -50042
rect 8160 -50948 8260 -50042
rect -5288 -51048 8260 -50948
rect -5288 -52948 -5188 -51048
rect -3182 -52948 -3082 -51048
rect -1076 -52948 -976 -51048
rect 1030 -52948 1130 -51048
rect 3136 -52948 3236 -51048
rect 5242 -52948 5342 -51048
rect 7368 -51942 7468 -51048
rect 8160 -51942 8260 -51048
rect 7330 -52042 8260 -51942
rect 7368 -52948 7468 -52042
rect 8160 -52948 8260 -52042
rect -5288 -52966 8264 -52948
rect -5288 -53030 8182 -52966
rect 8246 -53030 8264 -52966
rect -5288 -53048 8264 -53030
rect -5288 -54948 -5188 -53048
rect -3182 -54948 -3082 -53048
rect -1076 -54948 -976 -53048
rect 1030 -54948 1130 -53048
rect 3136 -54948 3236 -53048
rect 5242 -54948 5342 -53048
rect 7368 -53942 7468 -53048
rect 8160 -53942 8260 -53048
rect 7330 -54042 8260 -53942
rect 7368 -54948 7468 -54042
rect 8160 -54948 8260 -54042
rect -5288 -54966 8262 -54948
rect -5288 -55030 8180 -54966
rect 8244 -55030 8262 -54966
rect -5288 -55048 8262 -55030
rect -5288 -56948 -5188 -55048
rect -3182 -56948 -3082 -55048
rect -1076 -56948 -976 -55048
rect 1030 -56948 1130 -55048
rect 3136 -56948 3236 -55048
rect 5242 -56948 5342 -55048
rect 7368 -55942 7468 -55048
rect 8160 -55942 8260 -55048
rect 7330 -56042 8260 -55942
rect 7368 -56948 7468 -56042
rect 8160 -56948 8260 -56042
rect -5288 -57048 8260 -56948
rect -5288 -58948 -5188 -57048
rect -3182 -58948 -3082 -57048
rect -1076 -58948 -976 -57048
rect 1030 -58948 1130 -57048
rect 3136 -58948 3236 -57048
rect 5242 -58948 5342 -57048
rect 7368 -57942 7468 -57048
rect 8160 -57942 8260 -57048
rect 9250 -56658 9554 -56598
rect 9250 -56894 9284 -56658
rect 9520 -56894 9554 -56658
rect 9250 -56953 9372 -56894
rect 9436 -56953 9554 -56894
rect 9250 -56969 9554 -56953
rect 9250 -56978 9372 -56969
rect 9436 -56978 9554 -56969
rect 9250 -57214 9284 -56978
rect 9520 -57214 9554 -56978
rect 9250 -57273 9372 -57214
rect 9436 -57273 9554 -57214
rect 9250 -57289 9554 -57273
rect 9250 -57298 9372 -57289
rect 9436 -57298 9554 -57289
rect 9250 -57534 9284 -57298
rect 9520 -57534 9554 -57298
rect 9250 -57594 9554 -57534
rect 7330 -58042 8260 -57942
rect 7368 -58948 7468 -58042
rect 8160 -58948 8260 -58042
rect -5288 -59048 8260 -58948
rect -5288 -60968 -5188 -59048
rect -3182 -60968 -3082 -59048
rect -1076 -60968 -976 -59048
rect 1030 -60968 1130 -59048
rect 3136 -60968 3236 -59048
rect 5242 -60968 5342 -59048
rect 7368 -59942 7468 -59048
rect 8160 -59942 8260 -59048
rect 10276 -58408 11076 -58378
rect 10276 -58429 12110 -58408
rect 10276 -58493 10330 -58429
rect 10394 -58493 10410 -58429
rect 10474 -58493 10490 -58429
rect 10554 -58493 10570 -58429
rect 10634 -58493 10650 -58429
rect 10714 -58493 10730 -58429
rect 10794 -58493 10810 -58429
rect 10874 -58493 10890 -58429
rect 10954 -58493 10970 -58429
rect 11034 -58493 11050 -58429
rect 11114 -58493 11130 -58429
rect 11194 -58493 11210 -58429
rect 11274 -58493 11290 -58429
rect 11354 -58493 11370 -58429
rect 11434 -58493 11450 -58429
rect 11514 -58493 11530 -58429
rect 11594 -58493 11610 -58429
rect 11674 -58493 11690 -58429
rect 11754 -58493 11770 -58429
rect 11834 -58493 11850 -58429
rect 11914 -58493 11930 -58429
rect 11994 -58493 12010 -58429
rect 12074 -58493 12110 -58429
rect 10276 -58500 12110 -58493
rect 10276 -59056 10398 -58500
rect 10954 -58514 12110 -58500
rect 49716 -58502 51344 -58380
rect 10954 -59056 11076 -58514
rect 10276 -59178 11076 -59056
rect 49716 -59058 50666 -58502
rect 51222 -59058 51344 -58502
rect 49716 -59180 51344 -59058
rect 7330 -60042 8260 -59942
rect 7368 -60968 7468 -60042
rect 8160 -60968 8260 -60042
rect -5288 -61068 8260 -60968
rect -5288 -61908 -5188 -61068
rect -3182 -61908 -3082 -61068
rect -1076 -61908 -976 -61068
rect 1030 -61908 1130 -61068
rect 3136 -61908 3236 -61068
rect 5242 -61930 5342 -61068
rect 7368 -61930 7468 -61068
rect -7394 -62030 -6502 -61930
rect -5288 -61936 7476 -61930
rect 8160 -61936 8260 -61068
rect -5288 -62030 8260 -61936
rect 5202 -62036 8260 -62030
rect 8160 -62122 8260 -62036
rect -8282 -63040 -7828 -63022
rect -8282 -63104 -7910 -63040
rect -7846 -63104 -7828 -63040
rect -8282 -63122 -7828 -63104
rect -25201 -63296 -25099 -63277
rect -25201 -63360 -25182 -63296
rect -25118 -63360 -25099 -63296
rect -25201 -63379 -25099 -63360
rect -27764 -64414 9542 -64348
rect -27764 -64970 7106 -64414
rect 7662 -64970 8920 -64414
rect 9476 -64970 9542 -64414
rect -27764 -65036 9542 -64970
rect -26889 -69716 -26223 -69222
rect -22859 -69716 -22193 -69222
rect -18837 -69716 -18171 -69222
rect -14853 -69716 -14187 -69222
rect -10909 -69716 -10243 -69222
rect -6853 -69716 -6187 -69222
rect -2875 -69716 -2209 -69222
rect 1153 -69716 1819 -69222
rect 5131 -69716 5797 -69222
rect 9356 -69716 11076 -69714
rect -27762 -69836 11076 -69716
rect -27762 -70392 10398 -69836
rect 10954 -70392 11076 -69836
rect -27762 -70514 11076 -70392
rect -27762 -70516 10276 -70514
rect -26889 -70941 -26223 -70516
rect -22859 -70875 -22193 -70516
rect -18837 -70901 -18171 -70516
rect -14853 -70913 -14187 -70516
rect -10909 -70853 -10243 -70516
rect -6853 -70859 -6187 -70516
rect -2875 -70877 -2209 -70516
rect 1153 -70889 1819 -70516
rect 5131 -70871 5797 -70516
rect -27760 -75220 7728 -75160
rect -27760 -75776 7106 -75220
rect 7662 -75776 7728 -75220
rect -27760 -75848 7728 -75776
<< via4 >>
rect 8910 -28256 9466 -27700
rect 50674 -28256 51230 -27700
rect 50674 -39358 51230 -38802
rect 50666 -43862 51222 -43306
rect 9284 -56729 9520 -56658
rect 9284 -56793 9372 -56729
rect 9372 -56793 9436 -56729
rect 9436 -56793 9520 -56729
rect 9284 -56809 9520 -56793
rect 9284 -56873 9372 -56809
rect 9372 -56873 9436 -56809
rect 9436 -56873 9520 -56809
rect 9284 -56889 9520 -56873
rect 9284 -56894 9372 -56889
rect 9372 -56894 9436 -56889
rect 9436 -56894 9520 -56889
rect 9284 -57033 9372 -56978
rect 9372 -57033 9436 -56978
rect 9436 -57033 9520 -56978
rect 9284 -57049 9520 -57033
rect 9284 -57113 9372 -57049
rect 9372 -57113 9436 -57049
rect 9436 -57113 9520 -57049
rect 9284 -57129 9520 -57113
rect 9284 -57193 9372 -57129
rect 9372 -57193 9436 -57129
rect 9436 -57193 9520 -57129
rect 9284 -57209 9520 -57193
rect 9284 -57214 9372 -57209
rect 9372 -57214 9436 -57209
rect 9436 -57214 9520 -57209
rect 9284 -57353 9372 -57298
rect 9372 -57353 9436 -57298
rect 9436 -57353 9520 -57298
rect 9284 -57369 9520 -57353
rect 9284 -57433 9372 -57369
rect 9372 -57433 9436 -57369
rect 9436 -57433 9520 -57369
rect 9284 -57449 9520 -57433
rect 9284 -57513 9372 -57449
rect 9372 -57513 9436 -57449
rect 9436 -57513 9520 -57449
rect 9284 -57534 9520 -57513
rect 10398 -59056 10954 -58500
rect 50666 -59058 51222 -58502
rect 7106 -64970 7662 -64414
rect 8920 -64970 9476 -64414
rect 10398 -70392 10954 -69836
rect 7106 -75776 7662 -75220
<< metal5 >>
rect 8764 -27700 9612 -27554
rect 8764 -28256 8910 -27700
rect 9466 -28256 9612 -27700
rect 8764 -28402 9612 -28256
rect 50528 -27700 51376 -27554
rect 50528 -28256 50674 -27700
rect 51230 -28256 51376 -27700
rect 50528 -28402 51376 -28256
rect 8788 -56658 9588 -28402
rect 50552 -38802 51352 -28402
rect 50552 -39358 50674 -38802
rect 51230 -39358 51352 -38802
rect 50552 -39480 51352 -39358
rect 50520 -43306 51368 -43160
rect 50520 -43862 50666 -43306
rect 51222 -43862 51368 -43306
rect 50520 -44008 51368 -43862
rect 8788 -56894 9284 -56658
rect 9520 -56894 9588 -56658
rect 8788 -56978 9588 -56894
rect 8788 -57214 9284 -56978
rect 9520 -57214 9588 -56978
rect 8788 -57298 9588 -57214
rect 8788 -57534 9284 -57298
rect 9520 -57534 9588 -57298
rect 7016 -64414 7752 -64324
rect 7016 -64970 7106 -64414
rect 7662 -64970 7752 -64414
rect 7016 -65060 7752 -64970
rect 8788 -64414 9588 -57534
rect 10252 -58500 11100 -58354
rect 10252 -59056 10398 -58500
rect 10954 -59056 11100 -58500
rect 10252 -59202 11100 -59056
rect 50544 -58502 51344 -44008
rect 50544 -59058 50666 -58502
rect 51222 -59058 51344 -58502
rect 50544 -59180 51344 -59058
rect 8788 -64970 8920 -64414
rect 9476 -64970 9588 -64414
rect 7040 -75220 7728 -65060
rect 8788 -65088 9588 -64970
rect 10276 -69836 11076 -59202
rect 10276 -70392 10398 -69836
rect 10954 -70392 11076 -69836
rect 10276 -70514 11076 -70392
rect 7040 -75776 7106 -75220
rect 7662 -75776 7728 -75220
rect 7040 -75842 7728 -75776
use amux_2to1  amux_2to1_17
timestamp 1626065694
transform 1 0 -28122 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_16
timestamp 1626065694
transform 1 0 -24122 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_15
timestamp 1626065694
transform 1 0 -20122 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_14
timestamp 1626065694
transform 1 0 -16122 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_13
timestamp 1626065694
transform 1 0 -12122 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_12
timestamp 1626065694
transform 1 0 -8122 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_11
timestamp 1626065694
transform 1 0 -4122 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_10
timestamp 1626065694
transform 1 0 -122 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_9
timestamp 1626065694
transform 1 0 3878 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_8
timestamp 1626065694
transform 1 0 -28122 0 1 -68088
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_7
timestamp 1626065694
transform 1 0 -24122 0 1 -68088
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_6
timestamp 1626065694
transform 1 0 -20122 0 1 -68088
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_5
timestamp 1626065694
transform 1 0 -16122 0 1 -68088
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_4
timestamp 1626065694
transform 1 0 -12122 0 1 -68088
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_3
timestamp 1626065694
transform 1 0 -8122 0 1 -68088
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_2
timestamp 1626065694
transform 1 0 -4122 0 1 -68088
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_1
timestamp 1626065694
transform 1 0 -122 0 1 -68088
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_0
timestamp 1626065694
transform 1 0 3878 0 1 -68088
box -114 -1800 2840 3740
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_320
timestamp 1626065694
transform 1 0 -26279 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_321
timestamp 1626065694
transform 1 0 -26279 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_322
timestamp 1626065694
transform 1 0 -28385 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_323
timestamp 1626065694
transform 1 0 -28385 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_318
timestamp 1626065694
transform 1 0 -24173 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_319
timestamp 1626065694
transform 1 0 -24173 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_314
timestamp 1626065694
transform 1 0 -19961 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_315
timestamp 1626065694
transform 1 0 -19961 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_316
timestamp 1626065694
transform 1 0 -22067 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_317
timestamp 1626065694
transform 1 0 -22067 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_312
timestamp 1626065694
transform 1 0 -17855 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_313
timestamp 1626065694
transform 1 0 -17855 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_308
timestamp 1626065694
transform 1 0 -13643 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_309
timestamp 1626065694
transform 1 0 -13643 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_310
timestamp 1626065694
transform 1 0 -15749 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_311
timestamp 1626065694
transform 1 0 -15749 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_306
timestamp 1626065694
transform 1 0 -11537 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_307
timestamp 1626065694
transform 1 0 -11537 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_304
timestamp 1626065694
transform 1 0 -9431 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_305
timestamp 1626065694
transform 1 0 -9431 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_300
timestamp 1626065694
transform 1 0 -5219 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_301
timestamp 1626065694
transform 1 0 -5219 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_302
timestamp 1626065694
transform 1 0 -7325 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_303
timestamp 1626065694
transform 1 0 -7325 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_298
timestamp 1626065694
transform 1 0 -3113 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_299
timestamp 1626065694
transform 1 0 -3113 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_294
timestamp 1626065694
transform 1 0 1099 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_295
timestamp 1626065694
transform 1 0 1099 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_296
timestamp 1626065694
transform 1 0 -1007 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_297
timestamp 1626065694
transform 1 0 -1007 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_292
timestamp 1626065694
transform 1 0 3205 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_293
timestamp 1626065694
transform 1 0 3205 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_290
timestamp 1626065694
transform 1 0 5311 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_291
timestamp 1626065694
transform 1 0 5311 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_288
timestamp 1626065694
transform 1 0 7417 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_289
timestamp 1626065694
transform 1 0 7417 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_282
timestamp 1626065694
transform 1 0 -26279 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_283
timestamp 1626065694
transform 1 0 -28385 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_284
timestamp 1626065694
transform 1 0 -26279 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_285
timestamp 1626065694
transform 1 0 -28385 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_286
timestamp 1626065694
transform 1 0 -26279 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_287
timestamp 1626065694
transform 1 0 -28385 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_279
timestamp 1626065694
transform 1 0 -24173 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_280
timestamp 1626065694
transform 1 0 -24173 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_281
timestamp 1626065694
transform 1 0 -24173 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_273
timestamp 1626065694
transform 1 0 -19961 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_274
timestamp 1626065694
transform 1 0 -19961 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_275
timestamp 1626065694
transform 1 0 -19961 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_276
timestamp 1626065694
transform 1 0 -22067 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_277
timestamp 1626065694
transform 1 0 -22067 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_278
timestamp 1626065694
transform 1 0 -22067 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_270
timestamp 1626065694
transform 1 0 -17855 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_271
timestamp 1626065694
transform 1 0 -17855 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_272
timestamp 1626065694
transform 1 0 -17855 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_264
timestamp 1626065694
transform 1 0 -13643 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_265
timestamp 1626065694
transform 1 0 -15749 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_266
timestamp 1626065694
transform 1 0 -13643 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_267
timestamp 1626065694
transform 1 0 -15749 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_268
timestamp 1626065694
transform 1 0 -13643 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_269
timestamp 1626065694
transform 1 0 -15749 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_261
timestamp 1626065694
transform 1 0 -11537 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_262
timestamp 1626065694
transform 1 0 -11537 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_263
timestamp 1626065694
transform 1 0 -11537 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_258
timestamp 1626065694
transform 1 0 -9431 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_259
timestamp 1626065694
transform 1 0 -9431 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_260
timestamp 1626065694
transform 1 0 -9431 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_252
timestamp 1626065694
transform 1 0 -5219 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_253
timestamp 1626065694
transform 1 0 -5219 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_254
timestamp 1626065694
transform 1 0 -5219 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_255
timestamp 1626065694
transform 1 0 -7325 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_256
timestamp 1626065694
transform 1 0 -7325 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_257
timestamp 1626065694
transform 1 0 -7325 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_249
timestamp 1626065694
transform 1 0 -3113 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_250
timestamp 1626065694
transform 1 0 -3113 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_251
timestamp 1626065694
transform 1 0 -3113 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_243
timestamp 1626065694
transform 1 0 1099 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_244
timestamp 1626065694
transform 1 0 -1007 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_245
timestamp 1626065694
transform 1 0 1099 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_246
timestamp 1626065694
transform 1 0 -1007 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_247
timestamp 1626065694
transform 1 0 1099 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_248
timestamp 1626065694
transform 1 0 -1007 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_240
timestamp 1626065694
transform 1 0 3205 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_241
timestamp 1626065694
transform 1 0 3205 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_242
timestamp 1626065694
transform 1 0 3205 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_237
timestamp 1626065694
transform 1 0 5311 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_238
timestamp 1626065694
transform 1 0 5311 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_239
timestamp 1626065694
transform 1 0 5311 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_234
timestamp 1626065694
transform 1 0 7417 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_235
timestamp 1626065694
transform 1 0 7417 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_236
timestamp 1626065694
transform 1 0 7417 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__nfet_01v8_N6QVV6  sky130_fd_pr__nfet_01v8_N6QVV6_0
timestamp 1626065694
transform 1 0 11201 0 1 -57946
box -931 -300 931 300
use sky130_fd_pr__pfet_01v8_hvt_SCHXZ7  sky130_fd_pr__pfet_01v8_hvt_SCHXZ7_0
timestamp 1626065694
transform 1 0 11201 0 1 -57122
box -941 -419 941 419
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_232
timestamp 1626065694
transform 1 0 -26279 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_233
timestamp 1626065694
transform 1 0 -28385 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_231
timestamp 1626065694
transform 1 0 -24173 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_229
timestamp 1626065694
transform 1 0 -19961 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_230
timestamp 1626065694
transform 1 0 -22067 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_228
timestamp 1626065694
transform 1 0 -17855 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_226
timestamp 1626065694
transform 1 0 -13643 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_227
timestamp 1626065694
transform 1 0 -15749 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_225
timestamp 1626065694
transform 1 0 -11537 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_224
timestamp 1626065694
transform 1 0 -9431 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_222
timestamp 1626065694
transform 1 0 -5219 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_223
timestamp 1626065694
transform 1 0 -7325 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_221
timestamp 1626065694
transform 1 0 -3113 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_219
timestamp 1626065694
transform 1 0 1099 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_220
timestamp 1626065694
transform 1 0 -1007 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_218
timestamp 1626065694
transform 1 0 3205 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_217
timestamp 1626065694
transform 1 0 5311 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_216
timestamp 1626065694
transform 1 0 7417 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_214
timestamp 1626065694
transform 1 0 -26279 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_215
timestamp 1626065694
transform 1 0 -28385 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_213
timestamp 1626065694
transform 1 0 -24173 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_212
timestamp 1626065694
transform 1 0 -22067 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_211
timestamp 1626065694
transform 1 0 -19961 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_210
timestamp 1626065694
transform 1 0 -17855 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_209
timestamp 1626065694
transform 1 0 -15749 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_208
timestamp 1626065694
transform 1 0 -13643 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_207
timestamp 1626065694
transform 1 0 -11537 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_206
timestamp 1626065694
transform 1 0 -9431 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_205
timestamp 1626065694
transform 1 0 -7325 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_204
timestamp 1626065694
transform 1 0 -5219 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_203
timestamp 1626065694
transform 1 0 -3113 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_202
timestamp 1626065694
transform 1 0 -1007 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_201
timestamp 1626065694
transform 1 0 1099 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_200
timestamp 1626065694
transform 1 0 3205 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_199
timestamp 1626065694
transform 1 0 5311 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_198
timestamp 1626065694
transform 1 0 7417 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_196
timestamp 1626065694
transform 1 0 -26279 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_197
timestamp 1626065694
transform 1 0 -28385 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_195
timestamp 1626065694
transform 1 0 -24173 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_194
timestamp 1626065694
transform 1 0 -22067 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_193
timestamp 1626065694
transform 1 0 -19961 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_192
timestamp 1626065694
transform 1 0 -17855 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_191
timestamp 1626065694
transform 1 0 -15749 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_190
timestamp 1626065694
transform 1 0 -13643 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_189
timestamp 1626065694
transform 1 0 -11537 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_188
timestamp 1626065694
transform 1 0 -9431 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_187
timestamp 1626065694
transform 1 0 -7325 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_186
timestamp 1626065694
transform 1 0 -5219 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_185
timestamp 1626065694
transform 1 0 -3113 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_184
timestamp 1626065694
transform 1 0 -1007 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_183
timestamp 1626065694
transform 1 0 1099 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_182
timestamp 1626065694
transform 1 0 3205 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_181
timestamp 1626065694
transform 1 0 5311 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_180
timestamp 1626065694
transform 1 0 7417 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_178
timestamp 1626065694
transform 1 0 -26279 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_179
timestamp 1626065694
transform 1 0 -28385 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_177
timestamp 1626065694
transform 1 0 -24173 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_176
timestamp 1626065694
transform 1 0 -22067 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_175
timestamp 1626065694
transform 1 0 -19961 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_174
timestamp 1626065694
transform 1 0 -17855 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_173
timestamp 1626065694
transform 1 0 -15749 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_172
timestamp 1626065694
transform 1 0 -13643 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_171
timestamp 1626065694
transform 1 0 -11537 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_170
timestamp 1626065694
transform 1 0 -9431 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_169
timestamp 1626065694
transform 1 0 -7325 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_168
timestamp 1626065694
transform 1 0 -5219 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_167
timestamp 1626065694
transform 1 0 -3113 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_166
timestamp 1626065694
transform 1 0 -1007 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_165
timestamp 1626065694
transform 1 0 1099 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_164
timestamp 1626065694
transform 1 0 3205 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_163
timestamp 1626065694
transform 1 0 5311 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_162
timestamp 1626065694
transform 1 0 7417 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_160
timestamp 1626065694
transform 1 0 -26279 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_161
timestamp 1626065694
transform 1 0 -28385 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_159
timestamp 1626065694
transform 1 0 -24173 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_158
timestamp 1626065694
transform 1 0 -22067 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_157
timestamp 1626065694
transform 1 0 -19961 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_156
timestamp 1626065694
transform 1 0 -17855 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_155
timestamp 1626065694
transform 1 0 -15749 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_154
timestamp 1626065694
transform 1 0 -13643 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_153
timestamp 1626065694
transform 1 0 -11537 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_152
timestamp 1626065694
transform 1 0 -9431 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_151
timestamp 1626065694
transform 1 0 -7325 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_150
timestamp 1626065694
transform 1 0 -5219 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_149
timestamp 1626065694
transform 1 0 -3113 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_148
timestamp 1626065694
transform 1 0 -1007 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_147
timestamp 1626065694
transform 1 0 1099 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_146
timestamp 1626065694
transform 1 0 3205 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_145
timestamp 1626065694
transform 1 0 5311 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_144
timestamp 1626065694
transform 1 0 7417 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_142
timestamp 1626065694
transform 1 0 -26279 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_143
timestamp 1626065694
transform 1 0 -28385 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_141
timestamp 1626065694
transform 1 0 -24173 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_140
timestamp 1626065694
transform 1 0 -22067 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_139
timestamp 1626065694
transform 1 0 -19961 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_138
timestamp 1626065694
transform 1 0 -17855 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_137
timestamp 1626065694
transform 1 0 -15749 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_136
timestamp 1626065694
transform 1 0 -13643 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_135
timestamp 1626065694
transform 1 0 -11537 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_134
timestamp 1626065694
transform 1 0 -9431 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_133
timestamp 1626065694
transform 1 0 -7325 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_132
timestamp 1626065694
transform 1 0 -5219 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_131
timestamp 1626065694
transform 1 0 -3113 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_130
timestamp 1626065694
transform 1 0 -1007 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_129
timestamp 1626065694
transform 1 0 1099 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_128
timestamp 1626065694
transform 1 0 3205 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_127
timestamp 1626065694
transform 1 0 5311 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_126
timestamp 1626065694
transform 1 0 7417 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_122
timestamp 1626065694
transform 1 0 -26279 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_123
timestamp 1626065694
transform 1 0 -28385 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_124
timestamp 1626065694
transform 1 0 -26279 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_125
timestamp 1626065694
transform 1 0 -28385 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_120
timestamp 1626065694
transform 1 0 -24173 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_121
timestamp 1626065694
transform 1 0 -24173 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_118
timestamp 1626065694
transform 1 0 -22067 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_119
timestamp 1626065694
transform 1 0 -22067 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_116
timestamp 1626065694
transform 1 0 -19961 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_117
timestamp 1626065694
transform 1 0 -19961 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_114
timestamp 1626065694
transform 1 0 -17855 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_115
timestamp 1626065694
transform 1 0 -17855 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_112
timestamp 1626065694
transform 1 0 -15749 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_113
timestamp 1626065694
transform 1 0 -15749 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_110
timestamp 1626065694
transform 1 0 -13643 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_111
timestamp 1626065694
transform 1 0 -13643 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_108
timestamp 1626065694
transform 1 0 -11537 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_109
timestamp 1626065694
transform 1 0 -11537 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_106
timestamp 1626065694
transform 1 0 -9431 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_107
timestamp 1626065694
transform 1 0 -9431 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_104
timestamp 1626065694
transform 1 0 -7325 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_105
timestamp 1626065694
transform 1 0 -7325 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_102
timestamp 1626065694
transform 1 0 -5219 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_103
timestamp 1626065694
transform 1 0 -5219 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_100
timestamp 1626065694
transform 1 0 -3113 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_101
timestamp 1626065694
transform 1 0 -3113 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_98
timestamp 1626065694
transform 1 0 -1007 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_99
timestamp 1626065694
transform 1 0 -1007 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_96
timestamp 1626065694
transform 1 0 1099 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_97
timestamp 1626065694
transform 1 0 1099 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_94
timestamp 1626065694
transform 1 0 3205 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_95
timestamp 1626065694
transform 1 0 3205 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_92
timestamp 1626065694
transform 1 0 5311 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_93
timestamp 1626065694
transform 1 0 5311 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_90
timestamp 1626065694
transform 1 0 7417 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_91
timestamp 1626065694
transform 1 0 7417 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_88
timestamp 1626065694
transform 1 0 -26279 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_89
timestamp 1626065694
transform 1 0 -28385 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_87
timestamp 1626065694
transform 1 0 -24173 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_86
timestamp 1626065694
transform 1 0 -22067 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_85
timestamp 1626065694
transform 1 0 -19961 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_84
timestamp 1626065694
transform 1 0 -17855 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_83
timestamp 1626065694
transform 1 0 -15749 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_82
timestamp 1626065694
transform 1 0 -13643 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_81
timestamp 1626065694
transform 1 0 -11537 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_80
timestamp 1626065694
transform 1 0 -9431 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_79
timestamp 1626065694
transform 1 0 -7325 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_78
timestamp 1626065694
transform 1 0 -5219 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_77
timestamp 1626065694
transform 1 0 -3113 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_76
timestamp 1626065694
transform 1 0 -1007 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_75
timestamp 1626065694
transform 1 0 1099 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_74
timestamp 1626065694
transform 1 0 3205 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_73
timestamp 1626065694
transform 1 0 5311 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_72
timestamp 1626065694
transform 1 0 7417 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_70
timestamp 1626065694
transform 1 0 -26279 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_71
timestamp 1626065694
transform 1 0 -28385 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_69
timestamp 1626065694
transform 1 0 -24173 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_68
timestamp 1626065694
transform 1 0 -22067 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_67
timestamp 1626065694
transform 1 0 -19961 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_66
timestamp 1626065694
transform 1 0 -17855 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_65
timestamp 1626065694
transform 1 0 -15749 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_64
timestamp 1626065694
transform 1 0 -13643 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_63
timestamp 1626065694
transform 1 0 -11537 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_62
timestamp 1626065694
transform 1 0 -9431 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_61
timestamp 1626065694
transform 1 0 -7325 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_60
timestamp 1626065694
transform 1 0 -5219 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_59
timestamp 1626065694
transform 1 0 -3113 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_58
timestamp 1626065694
transform 1 0 -1007 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_57
timestamp 1626065694
transform 1 0 1099 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_56
timestamp 1626065694
transform 1 0 3205 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_55
timestamp 1626065694
transform 1 0 5311 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_54
timestamp 1626065694
transform 1 0 7417 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_52
timestamp 1626065694
transform 1 0 -26279 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_53
timestamp 1626065694
transform 1 0 -28385 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_51
timestamp 1626065694
transform 1 0 -24173 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_50
timestamp 1626065694
transform 1 0 -22067 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_49
timestamp 1626065694
transform 1 0 -19961 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_48
timestamp 1626065694
transform 1 0 -17855 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_47
timestamp 1626065694
transform 1 0 -15749 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_46
timestamp 1626065694
transform 1 0 -13643 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_45
timestamp 1626065694
transform 1 0 -11537 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_44
timestamp 1626065694
transform 1 0 -9431 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_43
timestamp 1626065694
transform 1 0 -7325 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_42
timestamp 1626065694
transform 1 0 -5219 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_41
timestamp 1626065694
transform 1 0 -3113 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_40
timestamp 1626065694
transform 1 0 -1007 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_39
timestamp 1626065694
transform 1 0 1099 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_38
timestamp 1626065694
transform 1 0 3205 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_37
timestamp 1626065694
transform 1 0 5311 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_36
timestamp 1626065694
transform 1 0 7417 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_34
timestamp 1626065694
transform 1 0 -26279 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_35
timestamp 1626065694
transform 1 0 -28385 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_33
timestamp 1626065694
transform 1 0 -24173 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_32
timestamp 1626065694
transform 1 0 -22067 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_31
timestamp 1626065694
transform 1 0 -19961 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_30
timestamp 1626065694
transform 1 0 -17855 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_29
timestamp 1626065694
transform 1 0 -15749 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_28
timestamp 1626065694
transform 1 0 -13643 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_27
timestamp 1626065694
transform 1 0 -11537 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_26
timestamp 1626065694
transform 1 0 -9431 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_25
timestamp 1626065694
transform 1 0 -7325 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_24
timestamp 1626065694
transform 1 0 -5219 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_23
timestamp 1626065694
transform 1 0 -3113 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_22
timestamp 1626065694
transform 1 0 -1007 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_21
timestamp 1626065694
transform 1 0 1099 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_20
timestamp 1626065694
transform 1 0 3205 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_19
timestamp 1626065694
transform 1 0 5311 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_18
timestamp 1626065694
transform 1 0 7417 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_16
timestamp 1626065694
transform 1 0 -26279 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_17
timestamp 1626065694
transform 1 0 -28385 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_15
timestamp 1626065694
transform 1 0 -24173 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_14
timestamp 1626065694
transform 1 0 -22067 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_13
timestamp 1626065694
transform 1 0 -19961 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_12
timestamp 1626065694
transform 1 0 -17855 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_11
timestamp 1626065694
transform 1 0 -15749 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_10
timestamp 1626065694
transform 1 0 -13643 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_9
timestamp 1626065694
transform 1 0 -11537 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_8
timestamp 1626065694
transform 1 0 -9431 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_7
timestamp 1626065694
transform 1 0 -7325 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_6
timestamp 1626065694
transform 1 0 -5219 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_5
timestamp 1626065694
transform 1 0 -3113 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_4
timestamp 1626065694
transform 1 0 -1007 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_3
timestamp 1626065694
transform 1 0 1099 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_2
timestamp 1626065694
transform 1 0 3205 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_1
timestamp 1626065694
transform 1 0 5311 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_0
timestamp 1626065694
transform 1 0 7417 0 1 -28006
box -850 -800 849 800
use se_fold_casc_wide_swing_ota  se_fold_casc_wide_swing_ota_0
timestamp 1626065694
transform 1 0 25444 0 1 -31978
box -15168 -27248 25000 4400
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1626065694
transform -1 0 12456 0 1 -57802
box -38 -48 314 592
use latched_comparator_folded  latched_comparator_folded_0
timestamp 1626065694
transform 1 0 55478 0 1 -40970
box -3400 -3014 3047 2278
<< labels >>
flabel metal3 s -18928 -63224 -18910 -63206 1 FreeSans 600 0 0 0 c6m
flabel metal3 s -16804 -63244 -16796 -63228 1 FreeSans 600 0 0 0 c5m
flabel metal3 s -14718 -63246 -14704 -63230 1 FreeSans 600 0 0 0 c4m
flabel metal3 s -8458 -63254 -8442 -63236 1 FreeSans 600 0 0 0 c1m
flabel metal3 s -9900 -63276 -9878 -63242 1 FreeSans 600 0 0 0 cdumm
flabel metal3 s -7508 -63088 -7478 -63062 1 FreeSans 600 0 0 0 c0m
flabel metal4 s -27544 -70138 -27514 -70094 1 FreeSans 600 0 0 0 VSS
flabel metal4 s -27740 -64374 -27728 -64364 1 FreeSans 600 0 0 0 VDD
flabel metal3 s -28160 -74900 -28146 -74892 1 FreeSans 600 0 0 0 vref
flabel metal3 s -28452 -72922 -28438 -72906 1 FreeSans 600 0 0 0 vlow
flabel metal3 s -28232 -67966 -28214 -67946 1 FreeSans 600 0 0 0 vin
flabel metal3 s 12544 -58056 12562 -58044 1 FreeSans 600 0 0 0 sample
flabel metal2 s 12200 -57048 12212 -57040 1 FreeSans 600 0 0 0 adc_run
flabel metal1 s -28342 -72610 -28336 -72600 1 FreeSans 600 0 0 0 q7
flabel metal1 s -24328 -72616 -24316 -72604 1 FreeSans 600 0 0 0 q6
flabel metal1 s -20346 -72616 -20340 -72608 1 FreeSans 600 0 0 0 q5
flabel metal1 s -16352 -72620 -16346 -72608 1 FreeSans 600 0 0 0 q4
flabel metal1 s -12382 -72614 -12370 -72604 1 FreeSans 600 0 0 0 q3
flabel metal1 s -8362 -72620 -8352 -72608 1 FreeSans 600 0 0 0 q2
flabel metal1 s -356 -72608 -350 -72602 1 FreeSans 600 0 0 0 q1
flabel metal1 s 3634 -72616 3644 -72606 1 FreeSans 600 0 0 0 q0
flabel metal1 s 15262 -56936 15270 -56922 1 FreeSans 600 0 0 0 ibiasn
flabel metal3 s 10682 -52044 10722 -52028 1 FreeSans 600 0 0 0 vcom
flabel metal2 s 27012 -43058 27020 -43048 1 FreeSans 600 0 0 0 vcom_buf
flabel metal2 s 52036 -40050 52042 -40042 1 FreeSans 600 0 0 0 ibiasp
flabel metal2 s 52026 -42516 52034 -42508 1 FreeSans 600 0 0 0 adc_clk
flabel metal2 s 58410 -41968 58422 -41960 1 FreeSans 600 0 0 0 comp_out
flabel metal2 s 58400 -42168 58406 -42162 1 FreeSans 600 0 0 0 comp_outm
flabel metal3 s -25158 -63656 -25132 -63634 1 FreeSans 600 0 0 0 c7m
flabel metal3 s -12584 -63246 -12564 -63222 1 FreeSans 600 0 0 0 c2m
flabel metal3 s -10558 -63254 -10540 -63232 1 FreeSans 600 0 0 0 c3m
<< end >>
