.subckt user_analog_project_wrapper vdda1 vdda2 vssa1 vssa2 vccd1 vccd2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_stb_i wbs_cyc_i wbs_we_i wbs_sel_i[3],wbs_sel_i[2],wbs_sel_i[1],wbs_sel_i[0]
+ wbs_dat_i[31],wbs_dat_i[30],wbs_dat_i[29],wbs_dat_i[28],wbs_dat_i[27],wbs_dat_i[26],wbs_dat_i[25],wbs_dat_i[24],wbs_dat_i[23],wbs_dat_i[22],wbs_dat_i[21],wbs_dat_i[20],wbs_dat_i[19],wbs_dat_i[18],wbs_dat_i[17],wbs_dat_i[16],wbs_dat_i[15],wbs_dat_i[14],wbs_dat_i[13],wbs_dat_i[12],wbs_dat_i[11],wbs_dat_i[10],wbs_dat_i[9],wbs_dat_i[8],wbs_dat_i[7],wbs_dat_i[6],wbs_dat_i[5],wbs_dat_i[4],wbs_dat_i[3],wbs_dat_i[2],wbs_dat_i[1],wbs_dat_i[0]
+ wbs_adr_i[31],wbs_adr_i[30],wbs_adr_i[29],wbs_adr_i[28],wbs_adr_i[27],wbs_adr_i[26],wbs_adr_i[25],wbs_adr_i[24],wbs_adr_i[23],wbs_adr_i[22],wbs_adr_i[21],wbs_adr_i[20],wbs_adr_i[19],wbs_adr_i[18],wbs_adr_i[17],wbs_adr_i[16],wbs_adr_i[15],wbs_adr_i[14],wbs_adr_i[13],wbs_adr_i[12],wbs_adr_i[11],wbs_adr_i[10],wbs_adr_i[9],wbs_adr_i[8],wbs_adr_i[7],wbs_adr_i[6],wbs_adr_i[5],wbs_adr_i[4],wbs_adr_i[3],wbs_adr_i[2],wbs_adr_i[1],wbs_adr_i[0] wbs_ack_o
+ wbs_dat_o[31],wbs_dat_o[30],wbs_dat_o[29],wbs_dat_o[28],wbs_dat_o[27],wbs_dat_o[26],wbs_dat_o[25],wbs_dat_o[24],wbs_dat_o[23],wbs_dat_o[22],wbs_dat_o[21],wbs_dat_o[20],wbs_dat_o[19],wbs_dat_o[18],wbs_dat_o[17],wbs_dat_o[16],wbs_dat_o[15],wbs_dat_o[14],wbs_dat_o[13],wbs_dat_o[12],wbs_dat_o[11],wbs_dat_o[10],wbs_dat_o[9],wbs_dat_o[8],wbs_dat_o[7],wbs_dat_o[6],wbs_dat_o[5],wbs_dat_o[4],wbs_dat_o[3],wbs_dat_o[2],wbs_dat_o[1],wbs_dat_o[0]
+ la_data_in[127],la_data_in[126],la_data_in[125],la_data_in[124],la_data_in[123],la_data_in[122],la_data_in[121],la_data_in[120],la_data_in[119],la_data_in[118],la_data_in[117],la_data_in[116],la_data_in[115],la_data_in[114],la_data_in[113],la_data_in[112],la_data_in[111],la_data_in[110],la_data_in[109],la_data_in[108],la_data_in[107],la_data_in[106],la_data_in[105],la_data_in[104],la_data_in[103],la_data_in[102],la_data_in[101],la_data_in[100],la_data_in[99],la_data_in[98],la_data_in[97],la_data_in[96],la_data_in[95],la_data_in[94],la_data_in[93],la_data_in[92],la_data_in[91],la_data_in[90],la_data_in[89],la_data_in[88],la_data_in[87],la_data_in[86],la_data_in[85],la_data_in[84],la_data_in[83],la_data_in[82],la_data_in[81],la_data_in[80],la_data_in[79],la_data_in[78],la_data_in[77],la_data_in[76],la_data_in[75],la_data_in[74],la_data_in[73],la_data_in[72],la_data_in[71],la_data_in[70],la_data_in[69],la_data_in[68],la_data_in[67],la_data_in[66],la_data_in[65],la_data_in[64],la_data_in[63],la_data_in[62],la_data_in[61],la_data_in[60],la_data_in[59],la_data_in[58],la_data_in[57],la_data_in[56],la_data_in[55],la_data_in[54],la_data_in[53],la_data_in[52],la_data_in[51],la_data_in[50],la_data_in[49],la_data_in[48],la_data_in[47],la_data_in[46],la_data_in[45],la_data_in[44],la_data_in[43],la_data_in[42],la_data_in[41],la_data_in[40],la_data_in[39],la_data_in[38],la_data_in[37],la_data_in[36],la_data_in[35],la_data_in[34],la_data_in[33],la_data_in[32],la_data_in[31],la_data_in[30],la_data_in[29],la_data_in[28],la_data_in[27],la_data_in[26],la_data_in[25],la_data_in[24],la_data_in[23],la_data_in[22],la_data_in[21],la_data_in[20],la_data_in[19],la_data_in[18],la_data_in[17],la_data_in[16],la_data_in[15],la_data_in[14],la_data_in[13],la_data_in[12],la_data_in[11],la_data_in[10],la_data_in[9],la_data_in[8],la_data_in[7],la_data_in[6],la_data_in[5],la_data_in[4],la_data_in[3],la_data_in[2],la_data_in[1],la_data_in[0]
+ la_data_out[127],la_data_out[126],la_data_out[125],la_data_out[124],la_data_out[123],la_data_out[122],la_data_out[121],la_data_out[120],la_data_out[119],la_data_out[118],la_data_out[117],la_data_out[116],la_data_out[115],la_data_out[114],la_data_out[113],la_data_out[112],la_data_out[111],la_data_out[110],la_data_out[109],la_data_out[108],la_data_out[107],la_data_out[106],la_data_out[105],la_data_out[104],la_data_out[103],la_data_out[102],la_data_out[101],la_data_out[100],la_data_out[99],la_data_out[98],la_data_out[97],la_data_out[96],la_data_out[95],la_data_out[94],la_data_out[93],la_data_out[92],la_data_out[91],la_data_out[90],la_data_out[89],la_data_out[88],la_data_out[87],la_data_out[86],la_data_out[85],la_data_out[84],la_data_out[83],la_data_out[82],la_data_out[81],la_data_out[80],la_data_out[79],la_data_out[78],la_data_out[77],la_data_out[76],la_data_out[75],la_data_out[74],la_data_out[73],la_data_out[72],la_data_out[71],la_data_out[70],la_data_out[69],la_data_out[68],la_data_out[67],la_data_out[66],la_data_out[65],la_data_out[64],la_data_out[63],la_data_out[62],la_data_out[61],la_data_out[60],la_data_out[59],la_data_out[58],la_data_out[57],la_data_out[56],la_data_out[55],la_data_out[54],la_data_out[53],la_data_out[52],la_data_out[51],la_data_out[50],la_data_out[49],la_data_out[48],la_data_out[47],la_data_out[46],la_data_out[45],la_data_out[44],la_data_out[43],la_data_out[42],la_data_out[41],la_data_out[40],la_data_out[39],la_data_out[38],la_data_out[37],la_data_out[36],la_data_out[35],la_data_out[34],la_data_out[33],la_data_out[32],la_data_out[31],la_data_out[30],la_data_out[29],la_data_out[28],la_data_out[27],la_data_out[26],la_data_out[25],la_data_out[24],la_data_out[23],la_data_out[22],la_data_out[21],la_data_out[20],la_data_out[19],la_data_out[18],la_data_out[17],la_data_out[16],la_data_out[15],la_data_out[14],la_data_out[13],la_data_out[12],la_data_out[11],la_data_out[10],la_data_out[9],la_data_out[8],la_data_out[7],la_data_out[6],la_data_out[5],la_data_out[4],la_data_out[3],la_data_out[2],la_data_out[1],la_data_out[0]
+ io_in[26],io_in[25],io_in[24],io_in[23],io_in[22],io_in[21],io_in[20],io_in[19],io_in[18],io_in[17],io_in[16],io_in[15],io_in[14],io_in[13],io_in[12],io_in[11],io_in[10],io_in[9],io_in[8],io_in[7],io_in[6],io_in[5],io_in[4],io_in[3],io_in[2],io_in[1],io_in[0]
+ io_in_3v3[26],io_in_3v3[25],io_in_3v3[24],io_in_3v3[23],io_in_3v3[22],io_in_3v3[21],io_in_3v3[20],io_in_3v3[19],io_in_3v3[18],io_in_3v3[17],io_in_3v3[16],io_in_3v3[15],io_in_3v3[14],io_in_3v3[13],io_in_3v3[12],io_in_3v3[11],io_in_3v3[10],io_in_3v3[9],io_in_3v3[8],io_in_3v3[7],io_in_3v3[6],io_in_3v3[5],io_in_3v3[4],io_in_3v3[3],io_in_3v3[2],io_in_3v3[1],io_in_3v3[0] user_clock2
+ io_out[26],io_out[25],io_out[24],io_out[23],io_out[22],io_out[21],io_out[20],io_out[19],io_out[18],io_out[17],io_out[16],io_out[15],io_out[14],io_out[13],io_out[12],io_out[11],io_out[10],io_out[9],io_out[8],io_out[7],io_out[6],io_out[5],io_out[4],io_out[3],io_out[2],io_out[1],io_out[0]
+ io_oeb[26],io_oeb[25],io_oeb[24],io_oeb[23],io_oeb[22],io_oeb[21],io_oeb[20],io_oeb[19],io_oeb[18],io_oeb[17],io_oeb[16],io_oeb[15],io_oeb[14],io_oeb[13],io_oeb[12],io_oeb[11],io_oeb[10],io_oeb[9],io_oeb[8],io_oeb[7],io_oeb[6],io_oeb[5],io_oeb[4],io_oeb[3],io_oeb[2],io_oeb[1],io_oeb[0]
+ gpio_analog[17],gpio_analog[16],gpio_analog[15],gpio_analog[14],gpio_analog[13],gpio_analog[12],gpio_analog[11],gpio_analog[10],gpio_analog[9],gpio_analog[8],gpio_analog[7],gpio_analog[6],gpio_analog[5],gpio_analog[4],gpio_analog[3],gpio_analog[2],gpio_analog[1],gpio_analog[0]
+ gpio_noesd[17],gpio_noesd[16],gpio_noesd[15],gpio_noesd[14],gpio_noesd[13],gpio_noesd[12],gpio_noesd[11],gpio_noesd[10],gpio_noesd[9],gpio_noesd[8],gpio_noesd[7],gpio_noesd[6],gpio_noesd[5],gpio_noesd[4],gpio_noesd[3],gpio_noesd[2],gpio_noesd[1],gpio_noesd[0]
+ io_analog[10],io_analog[9],io_analog[8],io_analog[7],io_analog[6],io_analog[5],io_analog[4],io_analog[3],io_analog[2],io_analog[1],io_analog[0] io_clamp_high[2],io_clamp_high[1],io_clamp_high[0] io_clamp_low[2],io_clamp_low[1],io_clamp_low[0]
+ user_irq[2],user_irq[1],user_irq[0]
+ la_oenb[127],la_oenb[126],la_oenb[125],la_oenb[124],la_oenb[123],la_oenb[122],la_oenb[121],la_oenb[120],la_oenb[119],la_oenb[118],la_oenb[117],la_oenb[116],la_oenb[115],la_oenb[114],la_oenb[113],la_oenb[112],la_oenb[111],la_oenb[110],la_oenb[109],la_oenb[108],la_oenb[107],la_oenb[106],la_oenb[105],la_oenb[104],la_oenb[103],la_oenb[102],la_oenb[101],la_oenb[100],la_oenb[99],la_oenb[98],la_oenb[97],la_oenb[96],la_oenb[95],la_oenb[94],la_oenb[93],la_oenb[92],la_oenb[91],la_oenb[90],la_oenb[89],la_oenb[88],la_oenb[87],la_oenb[86],la_oenb[85],la_oenb[84],la_oenb[83],la_oenb[82],la_oenb[81],la_oenb[80],la_oenb[79],la_oenb[78],la_oenb[77],la_oenb[76],la_oenb[75],la_oenb[74],la_oenb[73],la_oenb[72],la_oenb[71],la_oenb[70],la_oenb[69],la_oenb[68],la_oenb[67],la_oenb[66],la_oenb[65],la_oenb[64],la_oenb[63],la_oenb[62],la_oenb[61],la_oenb[60],la_oenb[59],la_oenb[58],la_oenb[57],la_oenb[56],la_oenb[55],la_oenb[54],la_oenb[53],la_oenb[52],la_oenb[51],la_oenb[50],la_oenb[49],la_oenb[48],la_oenb[47],la_oenb[46],la_oenb[45],la_oenb[44],la_oenb[43],la_oenb[42],la_oenb[41],la_oenb[40],la_oenb[39],la_oenb[38],la_oenb[37],la_oenb[36],la_oenb[35],la_oenb[34],la_oenb[33],la_oenb[32],la_oenb[31],la_oenb[30],la_oenb[29],la_oenb[28],la_oenb[27],la_oenb[26],la_oenb[25],la_oenb[24],la_oenb[23],la_oenb[22],la_oenb[21],la_oenb[20],la_oenb[19],la_oenb[18],la_oenb[17],la_oenb[16],la_oenb[15],la_oenb[14],la_oenb[13],la_oenb[12],la_oenb[11],la_oenb[10],la_oenb[9],la_oenb[8],la_oenb[7],la_oenb[6],la_oenb[5],la_oenb[4],la_oenb[3],la_oenb[2],la_oenb[1],la_oenb[0]
*.iopin vdda1
*.iopin vdda2
*.iopin vssa1
*.iopin vssa2
*.iopin vccd1
*.iopin vccd2
*.iopin vssd1
*.iopin vssd2
*.ipin wb_clk_i
*.ipin wb_rst_i
*.ipin wbs_stb_i
*.ipin wbs_cyc_i
*.ipin wbs_we_i
*.ipin wbs_sel_i[3],wbs_sel_i[2],wbs_sel_i[1],wbs_sel_i[0]
*.ipin
*+ wbs_dat_i[31],wbs_dat_i[30],wbs_dat_i[29],wbs_dat_i[28],wbs_dat_i[27],wbs_dat_i[26],wbs_dat_i[25],wbs_dat_i[24],wbs_dat_i[23],wbs_dat_i[22],wbs_dat_i[21],wbs_dat_i[20],wbs_dat_i[19],wbs_dat_i[18],wbs_dat_i[17],wbs_dat_i[16],wbs_dat_i[15],wbs_dat_i[14],wbs_dat_i[13],wbs_dat_i[12],wbs_dat_i[11],wbs_dat_i[10],wbs_dat_i[9],wbs_dat_i[8],wbs_dat_i[7],wbs_dat_i[6],wbs_dat_i[5],wbs_dat_i[4],wbs_dat_i[3],wbs_dat_i[2],wbs_dat_i[1],wbs_dat_i[0]
*.ipin
*+ wbs_adr_i[31],wbs_adr_i[30],wbs_adr_i[29],wbs_adr_i[28],wbs_adr_i[27],wbs_adr_i[26],wbs_adr_i[25],wbs_adr_i[24],wbs_adr_i[23],wbs_adr_i[22],wbs_adr_i[21],wbs_adr_i[20],wbs_adr_i[19],wbs_adr_i[18],wbs_adr_i[17],wbs_adr_i[16],wbs_adr_i[15],wbs_adr_i[14],wbs_adr_i[13],wbs_adr_i[12],wbs_adr_i[11],wbs_adr_i[10],wbs_adr_i[9],wbs_adr_i[8],wbs_adr_i[7],wbs_adr_i[6],wbs_adr_i[5],wbs_adr_i[4],wbs_adr_i[3],wbs_adr_i[2],wbs_adr_i[1],wbs_adr_i[0]
*.opin wbs_ack_o
*.opin
*+ wbs_dat_o[31],wbs_dat_o[30],wbs_dat_o[29],wbs_dat_o[28],wbs_dat_o[27],wbs_dat_o[26],wbs_dat_o[25],wbs_dat_o[24],wbs_dat_o[23],wbs_dat_o[22],wbs_dat_o[21],wbs_dat_o[20],wbs_dat_o[19],wbs_dat_o[18],wbs_dat_o[17],wbs_dat_o[16],wbs_dat_o[15],wbs_dat_o[14],wbs_dat_o[13],wbs_dat_o[12],wbs_dat_o[11],wbs_dat_o[10],wbs_dat_o[9],wbs_dat_o[8],wbs_dat_o[7],wbs_dat_o[6],wbs_dat_o[5],wbs_dat_o[4],wbs_dat_o[3],wbs_dat_o[2],wbs_dat_o[1],wbs_dat_o[0]
*.ipin
*+ la_data_in[127],la_data_in[126],la_data_in[125],la_data_in[124],la_data_in[123],la_data_in[122],la_data_in[121],la_data_in[120],la_data_in[119],la_data_in[118],la_data_in[117],la_data_in[116],la_data_in[115],la_data_in[114],la_data_in[113],la_data_in[112],la_data_in[111],la_data_in[110],la_data_in[109],la_data_in[108],la_data_in[107],la_data_in[106],la_data_in[105],la_data_in[104],la_data_in[103],la_data_in[102],la_data_in[101],la_data_in[100],la_data_in[99],la_data_in[98],la_data_in[97],la_data_in[96],la_data_in[95],la_data_in[94],la_data_in[93],la_data_in[92],la_data_in[91],la_data_in[90],la_data_in[89],la_data_in[88],la_data_in[87],la_data_in[86],la_data_in[85],la_data_in[84],la_data_in[83],la_data_in[82],la_data_in[81],la_data_in[80],la_data_in[79],la_data_in[78],la_data_in[77],la_data_in[76],la_data_in[75],la_data_in[74],la_data_in[73],la_data_in[72],la_data_in[71],la_data_in[70],la_data_in[69],la_data_in[68],la_data_in[67],la_data_in[66],la_data_in[65],la_data_in[64],la_data_in[63],la_data_in[62],la_data_in[61],la_data_in[60],la_data_in[59],la_data_in[58],la_data_in[57],la_data_in[56],la_data_in[55],la_data_in[54],la_data_in[53],la_data_in[52],la_data_in[51],la_data_in[50],la_data_in[49],la_data_in[48],la_data_in[47],la_data_in[46],la_data_in[45],la_data_in[44],la_data_in[43],la_data_in[42],la_data_in[41],la_data_in[40],la_data_in[39],la_data_in[38],la_data_in[37],la_data_in[36],la_data_in[35],la_data_in[34],la_data_in[33],la_data_in[32],la_data_in[31],la_data_in[30],la_data_in[29],la_data_in[28],la_data_in[27],la_data_in[26],la_data_in[25],la_data_in[24],la_data_in[23],la_data_in[22],la_data_in[21],la_data_in[20],la_data_in[19],la_data_in[18],la_data_in[17],la_data_in[16],la_data_in[15],la_data_in[14],la_data_in[13],la_data_in[12],la_data_in[11],la_data_in[10],la_data_in[9],la_data_in[8],la_data_in[7],la_data_in[6],la_data_in[5],la_data_in[4],la_data_in[3],la_data_in[2],la_data_in[1],la_data_in[0]
*.opin
*+ la_data_out[127],la_data_out[126],la_data_out[125],la_data_out[124],la_data_out[123],la_data_out[122],la_data_out[121],la_data_out[120],la_data_out[119],la_data_out[118],la_data_out[117],la_data_out[116],la_data_out[115],la_data_out[114],la_data_out[113],la_data_out[112],la_data_out[111],la_data_out[110],la_data_out[109],la_data_out[108],la_data_out[107],la_data_out[106],la_data_out[105],la_data_out[104],la_data_out[103],la_data_out[102],la_data_out[101],la_data_out[100],la_data_out[99],la_data_out[98],la_data_out[97],la_data_out[96],la_data_out[95],la_data_out[94],la_data_out[93],la_data_out[92],la_data_out[91],la_data_out[90],la_data_out[89],la_data_out[88],la_data_out[87],la_data_out[86],la_data_out[85],la_data_out[84],la_data_out[83],la_data_out[82],la_data_out[81],la_data_out[80],la_data_out[79],la_data_out[78],la_data_out[77],la_data_out[76],la_data_out[75],la_data_out[74],la_data_out[73],la_data_out[72],la_data_out[71],la_data_out[70],la_data_out[69],la_data_out[68],la_data_out[67],la_data_out[66],la_data_out[65],la_data_out[64],la_data_out[63],la_data_out[62],la_data_out[61],la_data_out[60],la_data_out[59],la_data_out[58],la_data_out[57],la_data_out[56],la_data_out[55],la_data_out[54],la_data_out[53],la_data_out[52],la_data_out[51],la_data_out[50],la_data_out[49],la_data_out[48],la_data_out[47],la_data_out[46],la_data_out[45],la_data_out[44],la_data_out[43],la_data_out[42],la_data_out[41],la_data_out[40],la_data_out[39],la_data_out[38],la_data_out[37],la_data_out[36],la_data_out[35],la_data_out[34],la_data_out[33],la_data_out[32],la_data_out[31],la_data_out[30],la_data_out[29],la_data_out[28],la_data_out[27],la_data_out[26],la_data_out[25],la_data_out[24],la_data_out[23],la_data_out[22],la_data_out[21],la_data_out[20],la_data_out[19],la_data_out[18],la_data_out[17],la_data_out[16],la_data_out[15],la_data_out[14],la_data_out[13],la_data_out[12],la_data_out[11],la_data_out[10],la_data_out[9],la_data_out[8],la_data_out[7],la_data_out[6],la_data_out[5],la_data_out[4],la_data_out[3],la_data_out[2],la_data_out[1],la_data_out[0]
*.ipin
*+ io_in[26],io_in[25],io_in[24],io_in[23],io_in[22],io_in[21],io_in[20],io_in[19],io_in[18],io_in[17],io_in[16],io_in[15],io_in[14],io_in[13],io_in[12],io_in[11],io_in[10],io_in[9],io_in[8],io_in[7],io_in[6],io_in[5],io_in[4],io_in[3],io_in[2],io_in[1],io_in[0]
*.ipin
*+ io_in_3v3[26],io_in_3v3[25],io_in_3v3[24],io_in_3v3[23],io_in_3v3[22],io_in_3v3[21],io_in_3v3[20],io_in_3v3[19],io_in_3v3[18],io_in_3v3[17],io_in_3v3[16],io_in_3v3[15],io_in_3v3[14],io_in_3v3[13],io_in_3v3[12],io_in_3v3[11],io_in_3v3[10],io_in_3v3[9],io_in_3v3[8],io_in_3v3[7],io_in_3v3[6],io_in_3v3[5],io_in_3v3[4],io_in_3v3[3],io_in_3v3[2],io_in_3v3[1],io_in_3v3[0]
*.ipin user_clock2
*.opin
*+ io_out[26],io_out[25],io_out[24],io_out[23],io_out[22],io_out[21],io_out[20],io_out[19],io_out[18],io_out[17],io_out[16],io_out[15],io_out[14],io_out[13],io_out[12],io_out[11],io_out[10],io_out[9],io_out[8],io_out[7],io_out[6],io_out[5],io_out[4],io_out[3],io_out[2],io_out[1],io_out[0]
*.opin
*+ io_oeb[26],io_oeb[25],io_oeb[24],io_oeb[23],io_oeb[22],io_oeb[21],io_oeb[20],io_oeb[19],io_oeb[18],io_oeb[17],io_oeb[16],io_oeb[15],io_oeb[14],io_oeb[13],io_oeb[12],io_oeb[11],io_oeb[10],io_oeb[9],io_oeb[8],io_oeb[7],io_oeb[6],io_oeb[5],io_oeb[4],io_oeb[3],io_oeb[2],io_oeb[1],io_oeb[0]
*.iopin
*+ gpio_analog[17],gpio_analog[16],gpio_analog[15],gpio_analog[14],gpio_analog[13],gpio_analog[12],gpio_analog[11],gpio_analog[10],gpio_analog[9],gpio_analog[8],gpio_analog[7],gpio_analog[6],gpio_analog[5],gpio_analog[4],gpio_analog[3],gpio_analog[2],gpio_analog[1],gpio_analog[0]
*.iopin
*+ gpio_noesd[17],gpio_noesd[16],gpio_noesd[15],gpio_noesd[14],gpio_noesd[13],gpio_noesd[12],gpio_noesd[11],gpio_noesd[10],gpio_noesd[9],gpio_noesd[8],gpio_noesd[7],gpio_noesd[6],gpio_noesd[5],gpio_noesd[4],gpio_noesd[3],gpio_noesd[2],gpio_noesd[1],gpio_noesd[0]
*.iopin
*+ io_analog[10],io_analog[9],io_analog[8],io_analog[7],io_analog[6],io_analog[5],io_analog[4],io_analog[3],io_analog[2],io_analog[1],io_analog[0]
*.iopin io_clamp_high[2],io_clamp_high[1],io_clamp_high[0]
*.iopin io_clamp_low[2],io_clamp_low[1],io_clamp_low[0]
*.opin user_irq[2],user_irq[1],user_irq[0]
*.ipin
*+ la_oenb[127],la_oenb[126],la_oenb[125],la_oenb[124],la_oenb[123],la_oenb[122],la_oenb[121],la_oenb[120],la_oenb[119],la_oenb[118],la_oenb[117],la_oenb[116],la_oenb[115],la_oenb[114],la_oenb[113],la_oenb[112],la_oenb[111],la_oenb[110],la_oenb[109],la_oenb[108],la_oenb[107],la_oenb[106],la_oenb[105],la_oenb[104],la_oenb[103],la_oenb[102],la_oenb[101],la_oenb[100],la_oenb[99],la_oenb[98],la_oenb[97],la_oenb[96],la_oenb[95],la_oenb[94],la_oenb[93],la_oenb[92],la_oenb[91],la_oenb[90],la_oenb[89],la_oenb[88],la_oenb[87],la_oenb[86],la_oenb[85],la_oenb[84],la_oenb[83],la_oenb[82],la_oenb[81],la_oenb[80],la_oenb[79],la_oenb[78],la_oenb[77],la_oenb[76],la_oenb[75],la_oenb[74],la_oenb[73],la_oenb[72],la_oenb[71],la_oenb[70],la_oenb[69],la_oenb[68],la_oenb[67],la_oenb[66],la_oenb[65],la_oenb[64],la_oenb[63],la_oenb[62],la_oenb[61],la_oenb[60],la_oenb[59],la_oenb[58],la_oenb[57],la_oenb[56],la_oenb[55],la_oenb[54],la_oenb[53],la_oenb[52],la_oenb[51],la_oenb[50],la_oenb[49],la_oenb[48],la_oenb[47],la_oenb[46],la_oenb[45],la_oenb[44],la_oenb[43],la_oenb[42],la_oenb[41],la_oenb[40],la_oenb[39],la_oenb[38],la_oenb[37],la_oenb[36],la_oenb[35],la_oenb[34],la_oenb[33],la_oenb[32],la_oenb[31],la_oenb[30],la_oenb[29],la_oenb[28],la_oenb[27],la_oenb[26],la_oenb[25],la_oenb[24],la_oenb[23],la_oenb[22],la_oenb[21],la_oenb[20],la_oenb[19],la_oenb[18],la_oenb[17],la_oenb[16],la_oenb[15],la_oenb[14],la_oenb[13],la_oenb[12],la_oenb[11],la_oenb[10],la_oenb[9],la_oenb[8],la_oenb[7],la_oenb[6],la_oenb[5],la_oenb[4],la_oenb[3],la_oenb[2],la_oenb[1],la_oenb[0]
x1 io_in[25] io_in[20] gpio_analog[9] io_in[14] io_in[24] io_out[0] gpio_analog[8] io_in[5] io_in[6]
+ io_in[23] io_in[21] io_in[26] io_out[2] io_out[1] io_in[4] io_in[3] gpio_analog[2] gpio_analog[3]
+ io_analog[7] io_analog[6] vccd1 vccd2 io_analog[1] io_analog[4] io_analog[5] io_analog[0] gpio_analog[6]
+ gpio_analog[10] gpio_analog[11] gpio_analog[5] gpio_analog[4] gpio_analog[15] io_analog[9] gpio_analog[0]
+ gpio_analog[1] io_analog[2] io_analog[3] io_analog[10] io_analog[8] gpio_analog[12] vssa1 vssd1 chip_top_level
R7 vssa1 io_clamp_low[2] sky130_fd_pr__res_generic_m1 W=0.6 L=3 mult=1 m=1
x2 vccd2 vssa1 io_analog[0] esd_cell
x3 vccd2 vssa1 io_analog[1] esd_cell
x4 vccd2 vssa1 io_analog[2] esd_cell
x5 vccd2 vssa1 io_analog[3] esd_cell
x6 vccd2 vssa1 io_analog[4] esd_cell
x7 vccd2 vssa1 io_analog[5] esd_cell
x8 vccd2 vssa1 io_analog[6] esd_cell
x9 vccd2 vssa1 io_analog[7] esd_cell
x10 vccd2 vssa1 io_analog[8] esd_cell
x11 vccd2 vssa1 io_analog[9] esd_cell
x12 vccd2 vssa1 io_analog[10] esd_cell
R1 vssd1 io_oeb[2] sky130_fd_pr__res_generic_m1 W=0.6 L=3 mult=1 m=1
R2 vssd1 io_oeb[1] sky130_fd_pr__res_generic_m1 W=0.6 L=3 mult=1 m=1
R3 vssd1 io_oeb[0] sky130_fd_pr__res_generic_m1 W=0.6 L=3 mult=1 m=1
R4 vssa1 io_clamp_high[2] sky130_fd_pr__res_generic_m1 W=0.6 L=3 mult=1 m=1
R5 vssa1 io_clamp_high[1] sky130_fd_pr__res_generic_m1 W=0.6 L=3 mult=1 m=1
R6 vssa1 io_clamp_high[0] sky130_fd_pr__res_generic_m1 W=0.6 L=3 mult=1 m=1
R8 vssa1 io_clamp_low[1] sky130_fd_pr__res_generic_m1 W=0.6 L=3 mult=1 m=1
R9 vssa1 io_clamp_low[0] sky130_fd_pr__res_generic_m1 W=0.6 L=3 mult=1 m=1
.ends

* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/chip_top_level.sym # of pins=42
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/chip_top_level.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/chip_top_level.sch
.subckt chip_top_level  adc_bypass_en adc_start amplitude_comparator_val clk debug_en freq_eval_done
+ frequency_comparator_val gain_ctrl_0 gain_ctrl_1 load_en rst_n serial_in serial_out serial_out_valid sram_select_0
+ sram_select_1 vampm vampp vbiasn vbiasp vccd1 vccd2 vcomp vcp vcp_sampled vfiltm vfiltp vhpf vincm vintm vintp
+ vlow_amplitude vlow_frequency vocm vocm_filt vpeak vpeak_sampled vref_amplitude vref_frequency vse vssa1 vssd1
*.ipin vssd1
*.ipin vssa1
*.opin vse
*.ipin vref_frequency
*.ipin vref_amplitude
*.opin vpeak_sampled
*.opin vpeak
*.ipin vocm_filt
*.ipin vocm
*.ipin vlow_frequency
*.ipin vlow_amplitude
*.opin vintp
*.opin vintm
*.ipin vincm
*.ipin vhpf
*.opin vfiltp
*.opin vfiltm
*.opin vcp_sampled
*.opin vcp
*.opin vcomp
*.ipin vccd2
*.ipin vccd1
*.ipin vbiasp
*.ipin vbiasn
*.opin vampp
*.opin vampm
*.ipin sram_select_1
*.opin serial_out_valid
*.opin serial_out
*.ipin serial_in
*.ipin rst_n
*.ipin load_en
*.ipin gain_ctrl_1
*.ipin gain_ctrl_0
*.opin frequency_comparator_val
*.opin freq_eval_done
*.ipin debug_en
*.ipin clk
*.opin amplitude_comparator_val
*.ipin adc_start
*.ipin adc_bypass_en
*.ipin sram_select_0
x1 vintp vfiltp vfiltm vintm vampm vampp vocm_filt vse vincm vccd2 vhpf vssa1 gain_ctrl_0
+ gain_ctrl_1 vocm sample clk net3 rst_n frequency_comparator_val vbiasp vbiasn sig_frequency_0 sig_frequency_1
+ sig_frequency_2 vcp sig_frequency_3 sig_frequency_4 sig_frequency_5 sig_frequency_6 vcp_sampled sig_frequency_7
+ vref_frequency vlow_frequency vcomp net4 amplitude_comparator_val vpeak_sampled net5 vpeak sig_amplitude_0
+ sig_amplitude_1 sig_amplitude_2 sig_amplitude_3 sig_amplitude_4 sig_amplitude_5 sig_amplitude_6 sig_amplitude_7
+ vref_amplitude vlow_amplitude analog_top_level_lvs

x2 clk rst_n adc_start frequency_comparator_val sample 
+ sig_frequency_7 sig_frequency_6 sig_frequency_5 sig_frequency_4 sig_frequency_3 sig_frequency_2
+ sig_frequency_1 sig_frequency_0 frequency_adc_done vssd1 vccd1 sar_adc_controller
*x2 sample vccd1 vssd1 sig_frequency_0 sig_frequency_1 clk sig_frequency_2 rst_n adc_start
*+ sig_frequency_3 sig_frequency_4 frequency_comparator_val sig_frequency_5 sig_frequency_6 sig_frequency_7 net2
*+ sar_adc_controller

x3 clk rst_n adc_start amplitude_comparator_val amplitude_run_adc_n 
+ sig_amplitude_7 sig_amplitude_6 sig_amplitude_5 sig_amplitude_4 sig_amplitude_3 sig_amplitude_2
+ sig_amplitude_1 sig_amplitude_0 amplitude_adc_done vssd1 vccd1 sar_adc_controller
*x3 net6 vccd1 vssd1 sig_amplitude_0 sig_amplitude_1 clk sig_amplitude_2 rst_n adc_start
*+ sig_amplitude_3 sig_amplitude_4 amplitude_comparator_val sig_amplitude_5 sig_amplitude_6 sig_amplitude_7 net1
*+ sar_adc_controller

x4 clk rst_n load_en debug_en serial_in 
+ sram_select_1 sram_select_0 frequency_adc_done amplitude_adc_done 
+ sig_frequency_7 sig_frequency_6 sig_frequency_5 sig_frequency_4 
+ sig_frequency_3 sig_frequency_2 sig_frequency_1 sig_frequency_0 
+ sig_amplitude_7 sig_amplitude_6 sig_amplitude_5 sig_amplitude_4 
+ sig_amplitude_3 sig_amplitude_2 sig_amplitude_1 sig_amplitude_0 
+ adc_bypass_en serial_out serial_out_valid freq_eval_done vssd1 vccd1 deconv_kernel_estimator_top_level
*x4 serial_out vccd1 serial_out_valid vssd1 clk freq_eval_done rst_n load_en debug_en serial_in
*+ sram_select_0 sram_select_1 net2 net1 sig_frequency_0 sig_frequency_1 sig_frequency_2 sig_frequency_3
*+ sig_frequency_4 sig_frequency_5 sig_frequency_6 sig_frequency_7 sig_amplitude_0 sig_amplitude_1 sig_amplitude_2
*+ sig_amplitude_3 sig_amplitude_4 sig_amplitude_5 sig_amplitude_6 sig_amplitude_7 adc_bypass_en
*+ deconv_kernel_estimator_top_level
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/esd_cell.sym # of pins=3
* sym_path: /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/esd_cell.sym
* sch_path: /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/esd_cell.sch
.subckt esd_cell  VDD VSS clamp
*.iopin clamp
*.ipin VDD
*.ipin VSS
XM1 clamp VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=20 m=20 
XM2 clamp VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=20 m=20 
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/analog_top_level_lvs.sym # of pins=50
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/analog_top_level_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/analog_top_level_lvs.sch
.subckt analog_top_level_lvs  vintp vfiltp vfiltm vintm vampm vampp vocm_filt vse vincm VDD vhpf VSS
+ gain_ctrl_0 gain_ctrl_1 vocm sample adc_clk adc_vcaparrayA rst_n adc_compA vbiasp vbiasn q0A q1A q2A vcp q3A
+ q4A q5A q6A vcp_sampled q7A vrefA vlowA vcomp adc_vcaparrayB adc_compB vpeak_sampled peak_detector_rst
+ vpeak q0B q1B q2B q3B q4B q5B q6B q7B vrefB vlowB
*.opin vintp
*.opin vintm
*.opin vfiltp
*.opin vfiltm
*.ipin vlowA
*.ipin vrefA
*.ipin q7A
*.ipin q6A
*.ipin q5A
*.ipin q4A
*.ipin q3A
*.ipin q2A
*.ipin q1A
*.ipin q0A
*.ipin adc_clk
*.ipin sample
*.ipin vlowB
*.ipin vrefB
*.ipin q7B
*.ipin q6B
*.ipin q5B
*.ipin q4B
*.ipin q3B
*.ipin q2B
*.ipin q1B
*.ipin q0B
*.opin adc_compA
*.opin adc_compB
*.opin vcp
*.opin vcp_sampled
*.opin vpeak_sampled
*.opin vpeak
*.opin vse
*.opin vcomp
*.ipin vhpf
*.ipin VDD
*.ipin VSS
*.ipin vincm
*.ipin vocm
*.ipin vocm_filt
*.ipin gain_ctrl_0
*.ipin gain_ctrl_1
*.ipin vbiasp
*.ipin vbiasn
*.opin peak_detector_rst
*.opin vampm
*.opin vampp
*.opin adc_vcaparrayB
*.opin adc_vcaparrayA
*.ipin rst_n
x1 VDD VSS vincm vhpf gain_ctrl_0 gain_ctrl_1 vocm net1 net2 rst_n vampm vampp input_amplifier_lvs
x2 VDD VSS vampp vampm net6 net5 net4 net3 vocm_filt vfiltp vfiltm vintp vintm
+ biquad_gm_c_filter_lvs
x3 vocm_filt VDD VSS vfiltp vse net7 vfiltm rst_n diff_to_se_converter_lvs
x5 VDD VSS net16 net15 vbiasp vbiasn net9 net17 net7 net13 net14 net8 net6 net5 net11 net12 net3
+ net4 net10 net2 net1 bias_current_distribution_lvs
x6 vfiltp vfiltm vcomp net8 VDD VSS comparator_lvs
x4 VDD VSS vse net9 net18 vpeak net10 peak_detector_rst peak_detector_lvs
x7 VDD sample VSS net19 vcp vcp_sampled net12 sample_and_hold_lvs
x8 VDD sample VSS net20 vpeak vpeak_sampled net13 sample_and_hold_lvs
x9 vcp VDD VSS vcomp net11 low_freq_pll_block_lvs
x10 adc_vcaparrayA VDD sample net14 net21 VSS adc_compA adc_clk net15 vcp_sampled q0A q1A q2A q7A
+ q3A q4A q5A q6A vrefA vlowA dac_8bit_lvs
x11 adc_vcaparrayB VDD sample net17 net22 VSS adc_compB adc_clk net16 vpeak_sampled q0B q1B q2B q7B
+ q3B q4B q5B q6B vrefB vlowB dac_8bit_lvs
x12 VDD VSS sample peak_detector_rst adc_clk pulse_generator_lvs
.ends


** expanding   symbol:
**+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/sar_adc_controller.sym # of pins=16
** sym_path:
**+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/sar_adc_controller.sym
** sch_path:
**+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/sar_adc_controller.sch
*.subckt sar_adc_controller  run_adc_n VDD VSS adc_val[0] adc_val[1] clk adc_val[2] rst_n adc_start
*+ adc_val[3] adc_val[4] comparator_val adc_val[5] adc_val[6] adc_val[7] out_valid
**.ipin VDD
**.ipin VSS
**.ipin clk
**.ipin rst_n
**.ipin adc_start
**.ipin comparator_val
**.opin run_adc_n
**.opin adc_val[0]
**.opin out_valid
**.opin adc_val[1]
**.opin adc_val[2]
**.opin adc_val[3]
**.opin adc_val[4]
**.opin adc_val[5]
**.opin adc_val[6]
**.opin adc_val[7]
*.ends
*
*
** expanding   symbol:
**+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/deconv_kernel_estimator_top_level.sym # of pins=31
** sym_path:
**+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/deconv_kernel_estimator_top_level.sym
** sch_path:
**+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/deconv_kernel_estimator_top_level.sch
*.subckt deconv_kernel_estimator_top_level  serial_out VDD serial_out_valid VSS clk freq_eval_done
*+ rst_n load_en debug_en serial_in sram_select[0] sram_select[1] frequency_adc_done amplitude_adc_done
*+ sig_frequency[0] sig_frequency[1] sig_frequency[2] sig_frequency[3] sig_frequency[4] sig_frequency[5]
*+ sig_frequency[6] sig_frequency[7] sig_amplitude[0] sig_amplitude[1] sig_amplitude[2] sig_amplitude[3]
*+ sig_amplitude[4] sig_amplitude[5] sig_amplitude[6] sig_amplitude[7] adc_bypass_en
**.ipin VDD
**.ipin VSS
**.ipin clk
**.ipin rst_n
**.ipin load_en
**.ipin debug_en
**.opin serial_out
**.opin serial_out_valid
**.opin freq_eval_done
**.ipin serial_in
**.ipin sram_select[0]
**.ipin sram_select[1]
**.ipin frequency_adc_done
**.ipin amplitude_adc_done
**.ipin sig_frequency[0]
**.ipin sig_frequency[1]
**.ipin sig_frequency[2]
**.ipin sig_frequency[3]
**.ipin sig_frequency[4]
**.ipin sig_frequency[5]
**.ipin sig_frequency[6]
**.ipin sig_frequency[7]
**.ipin sig_amplitude[0]
**.ipin sig_amplitude[1]
**.ipin sig_amplitude[2]
**.ipin sig_amplitude[3]
**.ipin sig_amplitude[4]
**.ipin sig_amplitude[5]
**.ipin sig_amplitude[6]
**.ipin sig_amplitude[7]
**.ipin adc_bypass_en
*.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/input_amplifier_lvs.sym # of pins=12
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/input_amplifier_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/input_amplifier_lvs.sch
.subckt input_amplifier_lvs  VDD VSS vincm vhpf gain_ctrl_0 gain_ctrl_1 vocm ibiasn1 ibiasn2 rst_n
+ vom vop
*.ipin VDD
*.ipin VSS
*.ipin vincm
*.ipin vhpf
*.ipin gain_ctrl_0
*.ipin gain_ctrl_1
*.ipin vocm
*.ipin ibiasn1
*.opin vom
*.opin vop
*.ipin ibiasn2
*.ipin rst_n
x5 VDD gain_ctrl_1 VSS vom venm2 txgate_lvs
x6 VDD gain_ctrl_1 VSS vop venp2 txgate_lvs
x7 VDD gain_ctrl_0 VSS vip2 venm1 txgate_lvs
x8 VDD gain_ctrl_0 VSS vim2 venp1 txgate_lvs
XC1 vom vip2 sky130_fd_pr__cap_mim_m3_1 W=8 L=8 MF=2 m=2
XC2 vop vim2 sky130_fd_pr__cap_mim_m3_1 W=8 L=8 MF=2 m=2
XC4 venm2 vip2 sky130_fd_pr__cap_mim_m3_1 W=8 L=8 MF=6 m=6
XC6 venp2 vim2 sky130_fd_pr__cap_mim_m3_1 W=8 L=8 MF=6 m=6
XC5 venp1 vop1 sky130_fd_pr__cap_mim_m3_1 W=8 L=8 MF=4 m=4
XC7 vim2 vop1 sky130_fd_pr__cap_mim_m3_1 W=8 L=8 MF=4 m=4
XC3 vip2 vom1 sky130_fd_pr__cap_mim_m3_1 W=8 L=8 MF=4 m=4
XC8 venm1 vom1 sky130_fd_pr__cap_mim_m3_1 W=8 L=8 MF=4 m=4
XC9 vom1 vip1 sky130_fd_pr__cap_mim_m3_1 W=8 L=8 MF=4 m=4
XC10 vip1 vhpf sky130_fd_pr__cap_mim_m3_1 W=8 L=8 MF=4 m=4
XC11 vim1 vincm sky130_fd_pr__cap_mim_m3_1 W=8 L=8 MF=4 m=4
XC12 vop1 vim1 sky130_fd_pr__cap_mim_m3_1 W=8 L=8 MF=4 m=4
XC13 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=12 L=2 MF=20 m=20
XC14 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=8 L=2 MF=22 m=22
XC15 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=2 L=8 MF=24 m=24
x1 vom1 vop1 vip1 vim1 vocm VDD VSS ibiasn1 diff_fold_casc_ota_lvs
x2 vom vop vip2 vim2 vocm VDD VSS ibiasn2 diff_fold_casc_ota_lvs
x3 VDD rst VSS vincm vim1 txgate_lvs
x4 rst_n rst VDD VSS inv1
x9 VDD rst VSS vincm vip1 txgate_lvs
x10 VDD rst VSS vop1 vim2 txgate_lvs
x11 VDD rst VSS vom1 vip2 txgate_lvs
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/biquad_gm_c_filter_lvs.sym # of pins=13
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/biquad_gm_c_filter_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/biquad_gm_c_filter_lvs.sch
.subckt biquad_gm_c_filter_lvs  VDD VSS vip vim ibiasn1 ibiasn2 ibiasn3 ibiasn4 vocm vfiltp vfiltm
+ vintp vintm
*.ipin VDD
*.ipin VSS
*.ipin vip
*.ipin vim
*.ipin ibiasn1
*.ipin vocm
*.opin vfiltp
*.opin vfiltm
*.opin vintp
*.opin vintm
*.ipin ibiasn2
*.ipin ibiasn3
*.ipin ibiasn4
x1 vintp vintm vip vim vocm VDD VSS ibiasn1 gm_c_stage_lvs Itail=0.01u Wp=0.5 Wn_diff=8 Wpcm=0.5
+ Wncm=8 Wn_bias=1 Lp=1 Ln_diff=1 Lpcm=1 Lncm=1 Ln_bias=4
x4 vintm vintp vfiltp vfiltm vocm VDD VSS ibiasn4 gm_c_stage_lvs Itail=0.01u Wp=0.5 Wn_diff=8
+ Wpcm=0.5 Wncm=8 Wn_bias=1 Lp=1 Ln_diff=1 Lpcm=1 Lncm=1 Ln_bias=4
x2 vfiltm vfiltp vintm vintp vocm VDD VSS ibiasn3 gm_c_stage_lvs Itail=0.01u Wp=0.5 Wn_diff=8
+ Wpcm=0.5 Wncm=8 Wn_bias=1 Lp=1 Ln_diff=1 Lpcm=1 Lncm=1 Ln_bias=4
x3 vintm vintp vintm vintp vocm VDD VSS ibiasn2 gm_c_stage_lvs Itail=0.01u Wp=0.5 Wn_diff=8 Wpcm=0.5
+ Wncm=8 Wn_bias=1 Lp=1 Ln_diff=1 Lpcm=1 Lncm=1 Ln_bias=4
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/diff_to_se_converter_lvs.sym # of pins=8
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/diff_to_se_converter_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/diff_to_se_converter_lvs.sch
.subckt diff_to_se_converter_lvs  vocm VDD VSS vdiffp vse ibiasn vdiffm rst_n
*.ipin vdiffp
*.ipin vdiffm
*.ipin VDD
*.ipin VSS
*.ipin vocm
*.opin vse
*.ipin ibiasn
*.ipin rst_n
x1 VSS vse vip vim ibiasn VDD se_fold_casc_wide_swing_ota_lvs
XC13 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=12 L=2 MF=8 m=8
XC14 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=8 L=2 MF=8 m=8
XC15 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=2 L=8 MF=8 m=8
XC1 vse vim sky130_fd_pr__cap_mim_m3_1 W=8 L=8 MF=4 m=4
XC2 vim vdiffm sky130_fd_pr__cap_mim_m3_1 W=8 L=8 MF=4 m=4
XC3 vip vdiffp sky130_fd_pr__cap_mim_m3_1 W=8 L=8 MF=4 m=4
XC4 vip vocm sky130_fd_pr__cap_mim_m3_1 W=8 L=8 MF=4 m=4
x2 VDD rst VSS vim vdiffm txgate_lvs
x3 rst_n rst VDD VSS inv1
x4 VDD rst VSS vip vdiffp txgate_lvs
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/bias_current_distribution_lvs.sym # of pins=21
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/bias_current_distribution_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/bias_current_distribution_lvs.sch
.subckt bias_current_distribution_lvs  VDD VSS dac_8bit_ibiasp_B dac_8bit_ibiasp_A vbiasp vbiasn
+ peak_detector_ibiasn1 dac_8bit_ibiasn_B diff_to_se_converter_ibiasn sample_and_hold_ibiasn_B dac_8bit_ibiasn_A
+ comparator_ibiasn biquad_gm_c_filter_ibiasn1 biquad_gm_c_filter_ibiasn2 low_freq_pll_ibiasn sample_and_hold_ibiasn_A
+ biquad_gm_c_filter_ibiasn4 biquad_gm_c_filter_ibiasn3 peak_detector_ibiasn2 input_amplifier_ibiasn2 input_amplifier_ibiasn1
*.ipin VDD
*.ipin VSS
*.ipin vbiasp
*.opin input_amplifier_ibiasn1
*.opin input_amplifier_ibiasn2
*.opin diff_to_se_converter_ibiasn
*.opin peak_detector_ibiasn1
*.opin peak_detector_ibiasn2
*.opin sample_and_hold_ibiasn_A
*.opin dac_8bit_ibiasn_A
*.opin sample_and_hold_ibiasn_B
*.opin dac_8bit_ibiasn_B
*.opin comparator_ibiasn
*.opin biquad_gm_c_filter_ibiasn1
*.opin biquad_gm_c_filter_ibiasn2
*.opin biquad_gm_c_filter_ibiasn3
*.opin biquad_gm_c_filter_ibiasn4
*.opin low_freq_pll_ibiasn
*.ipin vbiasn
*.opin dac_8bit_ibiasp_A
*.opin dac_8bit_ibiasp_B
XM1 input_amplifier_ibiasn1 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM2 input_amplifier_ibiasn2 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM3 diff_to_se_converter_ibiasn vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM4 peak_detector_ibiasn1 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM5 peak_detector_ibiasn2 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM6 sample_and_hold_ibiasn_A vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM7 dac_8bit_ibiasn_A vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM8 sample_and_hold_ibiasn_B vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM9 dac_8bit_ibiasn_B vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM10 comparator_ibiasn vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM11 biquad_gm_c_filter_ibiasn1 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM12 biquad_gm_c_filter_ibiasn2 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM13 biquad_gm_c_filter_ibiasn3 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM14 biquad_gm_c_filter_ibiasn4 vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM15 low_freq_pll_ibiasn vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM16 dac_8bit_ibiasp_A vbiasn VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM17 dac_8bit_ibiasp_B vbiasn VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM18 dac_8bit_ibiasp_A VSS VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM19 dac_8bit_ibiasp_B VSS VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM20 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=10 m=10 
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/comparator_lvs.sym # of pins=6
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/comparator_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/comparator_lvs.sch
.subckt comparator_lvs  vip vim vo ibiasn VDD VSS
*.ipin vip
*.ipin vim
*.opin vo
*.ipin ibiasn
*.ipin VDD
*.ipin VSS
XM6 vcompp vcompp VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM3 vcompm vcompm VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM2 vtail ibiasn VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM14 ibiasn ibiasn VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM4 vcompm vip vtail VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM1 vcompp vim vtail VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM5 vcompp vcompm VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM7 vcompm vcompp VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM8 vo1 vcompp VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM9 vo1 vmirror VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM10 vmirror vcompm VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM11 vmirror vmirror VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM13 vo vo1 VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM15 vo vo1 VDD VDD sky130_fd_pr__pfet_01v8_hvt L=1 W=4 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM12 vtail vtail vtail VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM16 ibiasn ibiasn ibiasn VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM18 vo1 vo1 vo1 VSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM19 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM20 vo1 vo1 vo1 VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM21 vmirror vmirror vmirror VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM17 vcompm vcompm vcompm VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/peak_detector_lvs.sym # of pins=8
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/peak_detector_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/peak_detector_lvs.sch
.subckt peak_detector_lvs  VDD VSS vin ibiasn1 vpeakh vpeak_out ibiasn2 rst
*.ipin vin
*.ipin ibiasn1
*.opin vpeak_out
*.ipin VDD
*.ipin VSS
*.opin vpeakh
*.ipin rst
*.ipin ibiasn2
XM3 vpeakh verr VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM4 verr verr VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM2 vpeakh rst VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
x2 VSS vpeak_out vpeakh vpeak_out ibiasn2 VDD se_fold_casc_wide_swing_ota_lvs
x1 VSS verr vpeak_out vin ibiasn1 VDD se_fold_casc_wide_swing_ota_lvs
XM1 vpeakh VDD VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XC3 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=31 L=2 MF=4 m=4
XC4 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=4 L=29 MF=4 m=4
XC5 VSS VSS sky130_fd_pr__cap_mim_m3_2 W=29 L=4 MF=4 m=4
XC6 VSS VSS sky130_fd_pr__cap_mim_m3_2 W=2 L=31 MF=4 m=4
XC1 vpeakh VSS sky130_fd_pr__cap_mim_m3_1 W=26 L=24 MF=4 m=4
XC7 VSS vpeakh sky130_fd_pr__cap_mim_m3_2 W=24 L=26 MF=4 m=4
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/sample_and_hold_lvs.sym # of pins=7
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/sample_and_hold_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/sample_and_hold_lvs.sch
.subckt sample_and_hold_lvs  VDD clk VSS vhold vin vout ibiasn
*.ipin vin
*.ipin clk
*.ipin VDD
*.ipin VSS
*.ipin ibiasn
*.opin vout
*.opin vhold
XM1 vhold clk vin VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM2 vholdm clk vout VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=8 m=8 
x1 VSS vout vhold vholdm ibiasn VDD se_fold_casc_wide_swing_ota_lvs
XC1 vhold VSS sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=4 m=4
XC2 vholdm vout sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=4 m=4
XC3 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=14 L=2 MF=4 m=4
XC4 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=2 L=12 MF=4 m=4
XC5 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=2 L=10 MF=4 m=4
XM3 vhold VSS VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM4 vholdm VSS VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM5 vin VSS VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM6 vout VSS VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/low_freq_pll_block_lvs.sym # of pins=5
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/low_freq_pll_block_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/low_freq_pll_block_lvs.sch
.subckt low_freq_pll_block_lvs  vcp VDD VSS vsigin ibiasn
*.ipin VDD
*.ipin VSS
*.ipin vsigin
*.ipin ibiasn
*.opin vcp
x1 VDD VSS net1 net3 vcp cs_ring_osc_lvs
x2 VDD VSS net1 net2 freq_div_lvs
x3 VDD VSS vsigin ibiasn vcp net2 pfd_cp_lpf_lvs
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/dac_8bit_lvs.sym # of pins=20
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/dac_8bit_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/dac_8bit_lvs.sch
.subckt dac_8bit_lvs  vcom VDD sample ibiasn comp_outm VSS comp_out adc_clk ibiasp vin q0 q1 q2 q7
+ q3 q4 q5 q6 vref vlow
*.ipin sample
*.ipin VDD
*.ipin VSS
*.ipin vlow
*.ipin vref
*.ipin vin
*.ipin q7
*.ipin q6
*.ipin q5
*.ipin q4
*.ipin q3
*.ipin q2
*.ipin q1
*.ipin q0
*.ipin ibiasn
*.ipin ibiasp
*.ipin adc_clk
*.opin comp_out
*.opin comp_outm
*.opin vcom
XM7 vcom adc_run vlow VDD sky130_fd_pr__pfet_01v8_hvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM8 vlow sample vcom VSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
x3 sample adc_run VDD VSS inv1
x2 VSS vcom_buf vcom vcom_buf ibiasn VDD se_fold_casc_wide_swing_ota_lvs
x1 vcom_buf vlow comp_out comp_outm ibiasp VDD VSS adc_clk latched_comparator_folded_lvs
x4 VSS vref net9 vlow VDD VSS amux_2to1_lvs
x5 q0 vref net8 vlow VDD VSS amux_2to1_lvs
x6 q1 vref net7 vlow VDD VSS amux_2to1_lvs
x7 q2 vref net6 vlow VDD VSS amux_2to1_lvs
x8 q3 vref net5 vlow VDD VSS amux_2to1_lvs
x9 q4 vref net4 vlow VDD VSS amux_2to1_lvs
x10 q5 vref net3 vlow VDD VSS amux_2to1_lvs
x11 q6 vref net2 vlow VDD VSS amux_2to1_lvs
x12 q7 vref net1 vlow VDD VSS amux_2to1_lvs
x13 sample vin cdumm net9 VDD VSS amux_2to1_lvs
x14 sample vin c0m net8 VDD VSS amux_2to1_lvs
x15 sample vin c1m net7 VDD VSS amux_2to1_lvs
x16 sample vin c2m net6 VDD VSS amux_2to1_lvs
x17 sample vin c3m net5 VDD VSS amux_2to1_lvs
x18 sample vin c4m net4 VDD VSS amux_2to1_lvs
x19 sample vin c5m net3 VDD VSS amux_2to1_lvs
x20 sample vin c6m net2 VDD VSS amux_2to1_lvs
x21 sample vin c7m net1 VDD VSS amux_2to1_lvs
XC1 vcom cdumm sky130_fd_pr__cap_mim_m3_1 W=7 L=7 MF=1 m=1
XC2 vcom c0m sky130_fd_pr__cap_mim_m3_1 W=7 L=7 MF=1 m=1
XC3 vcom c1m sky130_fd_pr__cap_mim_m3_1 W=7 L=7 MF=2 m=2
XC4 vcom c2m sky130_fd_pr__cap_mim_m3_1 W=7 L=7 MF=4 m=4
XC5 vcom c3m sky130_fd_pr__cap_mim_m3_1 W=7 L=7 MF=8 m=8
XC6 vcom c4m sky130_fd_pr__cap_mim_m3_1 W=7 L=7 MF=16 m=16
XC7 vcom c5m sky130_fd_pr__cap_mim_m3_1 W=7 L=7 MF=32 m=32
XC8 vcom c6m sky130_fd_pr__cap_mim_m3_1 W=7 L=7 MF=64 m=64
XC9 vcom c7m sky130_fd_pr__cap_mim_m3_1 W=7 L=7 MF=128 m=128
XC10 vcom vcom sky130_fd_pr__cap_mim_m3_1 W=7 L=7 MF=68 m=68
XM1 vcom VSS VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM2 VDD VDD vcom VDD sky130_fd_pr__pfet_01v8_hvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/pulse_generator_lvs.sym # of pins=5
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/pulse_generator_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/pulse_generator_lvs.sch
.subckt pulse_generator_lvs  VDD VSS trigb pulse clk
*.ipin trigb
*.ipin VDD
*.ipin VSS
*.ipin clk
*.opin pulse
x1 net4 net2 clk net6 VDD VSS dff_stdcell
x2 trigb trig VDD VSS inv1
x3 net2 net7 clk net3 VDD VSS dff_stdcell
x4 net3 net1 clk net5 VDD VSS dff_stdcell
x5 trig net4 clk net8 VDD VSS dff_stdcell
x6 net2 pulse net1 VDD VSS and2 M=1
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/txgate_lvs.sym # of pins=5
* sym_path: /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/txgate_lvs.sym
* sch_path: /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/txgate_lvs.sch
.subckt txgate_lvs  VDD tx VSS out in
*.ipin in
*.opin out
*.ipin VDD
*.ipin VSS
*.ipin tx
XM7 in txb out VDD sky130_fd_pr__pfet_01v8_hvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM8 out tx in VSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM1 out VSS VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM2 VDD VDD out VDD sky130_fd_pr__pfet_01v8_hvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
x1 tx txb VDD VSS inv1
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/diff_fold_casc_ota_lvs.sym # of pins=8
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/diff_fold_casc_ota_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/diff_fold_casc_ota_lvs.sch
.subckt diff_fold_casc_ota_lvs  vom vop vip vim vocm VDD VSS ibiasn
*.opin vop
*.opin vom
*.ipin vip
*.ipin vim
*.ipin vocm
*.ipin ibiasn
*.ipin VDD
*.ipin VSS
XM41 M3d M3d vbias3 VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=50 m=50 
XM42 vbias3 M3d vbias4 VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM43 vbias4 vbias3 net1 VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=18 m=18 
XM44 net1 vbias4 VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=18 m=18 
XM45 M13d M13d VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM46 vcmn_casc_tail1 ibiasn VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM47 vcmn_casc_tail2 ibiasn VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM48 vcmcn2_casc vcmcn2_casc VDD VDD sky130_fd_pr__pfet_01v8 L=0.8 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=8 m=8 
XM49 vcmcn_casc vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 L=0.8 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=8 m=8 
XM50 ibiasn ibiasn VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM56 vcmc_casc vcmcn_casc VDD VDD sky130_fd_pr__pfet_01v8 L=0.8 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=8 m=8 
XM57 vcmcn1_casc vcmcn1_casc VDD VDD sky130_fd_pr__pfet_01v8 L=0.8 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=8 m=8 
XM1 M1d vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM5 vtail_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=18 m=18 
XM8 vfoldm vip vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt L=1.2 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=18 m=18 
XM3 M3d vbias2 M2d VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM2 M2d vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM6 M6d vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM4 vbias1 vbias2 M1d VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM13 M13d vbias2 M6d VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM7 vtail_casc vbias4 VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=18 m=18 
XM10 vcascnm vbias4 VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=18 m=18 
XM14 vcascnp vbias4 VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=18 m=18 
XM11 vom vbias3 vcascnm VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=18 m=18 
XM16 vop vbias3 vcascnp VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=18 m=18 
XM12 vom vbias2 vfoldm VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM17 vop vbias2 vfoldp VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM15 vfoldm vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=12 m=12 
XM18 vfoldp vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=12 m=12 
XM19 vcmc_casc vcmc_casc VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=18 m=18 
XM20 vcmcn_casc vom vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8_lvt L=0.8 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM21 vcmcn2_casc vocm vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8_lvt L=0.8 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM22 vcmcn_casc vop vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.8 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM23 vcmcn1_casc vocm vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.8 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM9 vfoldp vim vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt L=1.2 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=18 m=18 
XM26 vbias2 ibiasn VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM27 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=56 m=56 
XM24 vbias1 VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM25 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=10 m=10 
XM28 M3d VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM29 vfoldm VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM30 vfoldp VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM31 M13d VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM32 M6d VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM33 vcmc_casc VSS VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM34 M3d VSS VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM35 vbias4 VSS VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM36 M1d M1d M1d VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM37 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=9 m=9 
XM38 vop vop vop VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM40 M2d M2d M2d VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM51 vop vop vop VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM52 vom vom vom VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM53 vom vom vom VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM54 M2d M2d M2d VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM55 M1d M1d M1d VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM39 M6d M6d M6d VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM58 vtail_casc vtail_casc vtail_casc VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM59 vbias4 vbias4 vbias4 VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM60 vtail_casc vtail_casc vtail_casc VSS sky130_fd_pr__nfet_01v8_lvt L=1.2 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM61 vfoldm vfoldm vfoldm VSS sky130_fd_pr__nfet_01v8_lvt L=1.2 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM62 vfoldp vfoldp vfoldp VSS sky130_fd_pr__nfet_01v8_lvt L=1.2 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM63 vcmn_casc_tail2 vcmn_casc_tail2 vcmn_casc_tail2 VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM64 vcmn_casc_tail1 vcmn_casc_tail1 vcmn_casc_tail1 VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM65 ibiasn ibiasn ibiasn VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM66 vbias2 vbias2 vbias2 VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM67 vbias2 vbias2 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=8 m=8 
XM68 vbias1 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=8 m=8 
XM69 vcmcn_casc vcmcn_casc vcmcn_casc VSS sky130_fd_pr__nfet_01v8_lvt L=0.8 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM70 vcmcn_casc vcmcn_casc vcmcn_casc VDD sky130_fd_pr__pfet_01v8 L=0.8 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM71 vcmcn2_casc vcmcn2_casc vcmcn2_casc VDD sky130_fd_pr__pfet_01v8 L=0.8 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM72 vcmc_casc vcmc_casc vcmc_casc VDD sky130_fd_pr__pfet_01v8 L=0.8 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM73 vcmcn1_casc vcmcn1_casc vcmcn1_casc VDD sky130_fd_pr__pfet_01v8 L=0.8 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XC1 vop VSS sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=8 m=8
XC2 vom VSS sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=8 m=8
XC3 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=10 L=2 MF=8 m=8
XC4 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=2 L=10 MF=8 m=8
XC5 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=2 L=2 MF=4 m=4
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/inv1.sym # of pins=4
* sym_path: /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/inv1.sym
* sch_path: /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/inv1.sch
.subckt inv1  A Y VDD VSS
*.ipin A
*.opin Y
*.ipin VDD
*.ipin VSS
XM2 Y A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM1 Y A VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/gm_c_stage_lvs.sym # of pins=8
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/gm_c_stage_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/gm_c_stage_lvs.sch
.subckt gm_c_stage_lvs  vom vop vip vim vocm VDD VSS ibiasn   Itail=0.01u Wp=0.5 Wn_diff=8 Wpcm=0.5
+ Wncm=8 Wn_bias=1 Lp=1 Ln_diff=1 Lpcm=1 Lncm=1 Ln_bias=4
*.ipin vip
*.ipin vim
*.ipin vocm
*.opin vop
*.opin vom
*.ipin ibiasn
*.ipin VDD
*.ipin VSS
XM10 vcmn_tail2 ibiasn VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM12 ibiasn ibiasn VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=10 m=10 
XM8 vbiasp vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM9 vom vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM11 vop vbiasp VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM16 vcmcn vop vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM1 vom vip vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM2 vop vim vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM6 vcmcn vcmcn VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM20 vcmc vcmcn VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 vcmcn2 vcmcn2 VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 vcmcn1 vcmcn1 VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM17 vcmcn2 vocm vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM18 vcmcn1 vocm vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM19 vcmcn vom vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM3 vtail_diff ibiasn VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7 vtail_diff vcmc VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM13 vcmc vcmc VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM14 vbiasp ibiasn VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM15 vcmn_tail1 ibiasn VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM21 vbiasp VSS VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM22 vtail_diff VSS VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM23 vcmc VSS VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM24 vcmn_tail1 VSS VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM25 vcmn_tail2 VSS VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM26 ibiasn VSS VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM27 vcmcn VSS VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM28 vcmcn2 VSS VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM29 vom VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM30 vbiasp VDD VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM31 vom VDD VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM32 vop VDD VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM33 vcmcn VDD VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM34 vcmcn1 VDD VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM35 vcmcn2 VDD VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM36 vcmc VDD VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/se_fold_casc_wide_swing_ota_lvs.sym # of pins=6
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/se_fold_casc_wide_swing_ota_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/se_fold_casc_wide_swing_ota_lvs.sch
.subckt se_fold_casc_wide_swing_ota_lvs  VSS vo vip vim ibiasn VDD
*.ipin vip
*.ipin vim
*.opin vo
*.ipin ibiasn
*.ipin VDD
*.ipin VSS
XM11 vmirror vbias3 vcascnm VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=18 m=18 
XM12 vmirror vbias2 vcascpm VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=7 m=7 
XM5 vtail_cascn vbias4 VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=36 m=36 
XM6 vtail_cascp vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=12 m=12 
XM3 vcascnm vip vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM1 vcascpm vip vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=18 m=18 
XM7 M7d vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM8 M8d vbias2 M9d VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM9 M9d vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM13 M13d vbias1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=6 m=6 
XM14 vbias1 vbias2 M7d VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM16 M16d vbias2 M13d VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM26 vbias2 ibiasn VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM17 vbias1 vbias1 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=56 m=56 
XM10 vcascnp vbias4 VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=36 m=36 
XM18 vcascnm vbias4 VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=36 m=36 
XM4 vcascpp vim vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=18 m=18 
XM2 vcascnp vim vtail_cascp VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM15 vcascpp vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=12 m=12 
XM19 vcascpm vmirror VDD VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=12 m=12 
XM20 M21d vbias4 VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=18 m=18 
XM21 vbias4 vbias3 M21d VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=18 m=18 
XM22 M8d M8d vbias3 VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=40 m=40 
XM23 vbias3 M8d vbias4 VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM24 vo vbias3 vcascnp VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=18 m=18 
XM25 ibiasn ibiasn VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM27 M16d M16d VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM28 vo vbias2 vcascpp VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=7 m=7 
XM29 vbias1 VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM31 M8d VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM32 vcascpp VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=3 m=3 
XM33 vcascpm VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=3 m=3 
XM34 M16d VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM35 M13d VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM39 M7d M7d M7d VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM40 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=5 m=5 
XM41 vo vo vo VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM42 M9d M9d M9d VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM51 vo vo vo VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM52 vmirror vmirror vmirror VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM53 vmirror vmirror vmirror VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM54 M9d M9d M9d VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM55 M7d M7d M7d VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM43 M13d M13d M13d VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM58 vtail_cascn vtail_cascn vtail_cascn VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM60 vtail_cascn vtail_cascn vtail_cascn VSS sky130_fd_pr__nfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM61 vcascpm vcascpm vcascpm VSS sky130_fd_pr__nfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM62 vcascpp vcascpp vcascpp VSS sky130_fd_pr__nfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM66 ibiasn ibiasn ibiasn VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM67 vbias2 vbias2 vbias2 VSS sky130_fd_pr__nfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=8 m=8 
XM68 vbias1 vbias1 vbias1 VSS sky130_fd_pr__nfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=8 m=8 
XC3 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=31 L=2 MF=4 m=4
XC4 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=4 L=29 MF=4 m=4
XC1 vo VSS sky130_fd_pr__cap_mim_m3_1 W=26 L=24 MF=4 m=4
XM44 vcascpm vcascpm vcascpm VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM45 vcascpp vcascpp vcascpp VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM46 vo VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM47 vmirror VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM48 vcascnm vcascnm vcascnm VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM49 vcascnp vcascnp vcascnp VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM36 vcascnp vcascnp vcascnp VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM50 vcascnm vcascnm vcascnm VSS sky130_fd_pr__nfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM37 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM30 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=4.8 W=3 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=12 m=12 
XC2 VSS vo sky130_fd_pr__cap_mim_m3_2 W=24 L=26 MF=4 m=4
XC5 VSS VSS sky130_fd_pr__cap_mim_m3_2 W=29 L=4 MF=4 m=4
XC6 VSS VSS sky130_fd_pr__cap_mim_m3_2 W=2 L=31 MF=4 m=4
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/cs_ring_osc_lvs.sym # of pins=5
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/cs_ring_osc_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/cs_ring_osc_lvs.sch
.subckt cs_ring_osc_lvs  VDD VSS voscbuf vosc vctrl
*.ipin VDD
*.ipin VSS
*.ipin vctrl
*.opin voscbuf
*.opin vosc
XM7 vosc2 vosc VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM8 vosc2 vosc VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM9 voscbuf vosc2 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
XM10 voscbuf vosc2 VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=4 m=4 
x1 VDD vpbias net1 vosc vctrl VSS cs_ring_osc_stage_lvs_exp
x2 VDD vpbias net2 net1 vctrl VSS cs_ring_osc_stage_lvs_exp
x3 VDD vpbias net3 net2 vctrl VSS cs_ring_osc_stage_lvs_exp
x4 VDD vpbias net4 net3 vctrl VSS cs_ring_osc_stage_lvs_exp
x5 VDD vpbias net5 net4 vctrl VSS cs_ring_osc_stage_lvs_exp
x6 VDD vpbias net6 net5 vctrl VSS cs_ring_osc_stage_lvs_exp
XM3 vpbias vpbias net7 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM6 net7 vpbias net8 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM11 net8 vpbias net9 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM12 net9 vpbias net10 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM13 net10 vpbias net11 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM14 net11 vpbias net12 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM15 net12 vpbias net13 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM16 net13 vpbias VDD VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM37 vpbias vctrl net14 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM38 net14 vctrl net15 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM39 net15 vctrl net16 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM40 net16 vctrl net17 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM41 net17 vctrl net18 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM42 net18 vctrl net19 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM43 net19 vctrl net20 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM44 net20 vctrl VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM22 vosc net6 net21 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM23 net21 net6 net22 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM24 net22 net6 net23 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM25 net23 net6 net24 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM26 net24 net6 net25 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM27 net25 net6 net26 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM28 net26 net6 net27 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM29 net27 net6 VDD VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM45 vosc net6 net28 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM46 net28 net6 net29 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM47 net29 net6 net30 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM48 net30 net6 net31 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM49 net31 net6 net32 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM50 net32 net6 net33 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM51 net33 net6 net34 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM52 net34 net6 VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM1 vpbias VSS VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 vosc VSS VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM5 vosc VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM17 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM18 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/freq_div_lvs.sym # of pins=4
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/freq_div_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/freq_div_lvs.sch
.subckt freq_div_lvs  VDD VSS vin vout
*.ipin vin
*.opin vout
*.ipin VDD
*.ipin VSS
x1 net1 vdff1 vin net2 VDD VSS dff_stdcell
x2 net3 vdff2 vdff1 net4 VDD VSS dff_stdcell
x3 vdff3D vdff3 vdff2 vdff3QB VDD VSS dff_stdcell
x4 net5 vdff4 vdff3 net6 VDD VSS dff_stdcell
x5 net13 net15 vdff7 net14 VDD VSS dff_stdcell
x6 net11 vdff7 vdff6 net12 VDD VSS dff_stdcell
x7 net9 vdff6 vdff5 net10 VDD VSS dff_stdcell
x8 net7 vdff5 vdff4 net8 VDD VSS dff_stdcell
x31 net16 net18 net15 net17 VDD VSS dff_stdcell
x32 net19 net21 net18 net20 VDD VSS dff_stdcell
x33 net22 vout net21 net23 VDD VSS dff_stdcell
x15 net2 net24 VDD VSS inv1
x16 net24 net1 VDD VSS inv4
x9 net4 net25 VDD VSS inv1
x10 net25 net3 VDD VSS inv4
x11 vdff3QB net26 VDD VSS inv1
x12 net26 vdff3D VDD VSS inv4
x13 net6 net27 VDD VSS inv1
x14 net27 net5 VDD VSS inv4
x17 net8 net28 VDD VSS inv1
x18 net28 net7 VDD VSS inv4
x19 net10 net29 VDD VSS inv1
x20 net29 net9 VDD VSS inv4
x21 net12 net30 VDD VSS inv1
x22 net30 net11 VDD VSS inv4
x23 net14 net31 VDD VSS inv1
x24 net31 net13 VDD VSS inv4
x25 net17 net32 VDD VSS inv1
x26 net32 net16 VDD VSS inv4
x27 net20 net33 VDD VSS inv1
x28 net33 net19 VDD VSS inv4
x29 net23 net34 VDD VSS inv1
x30 net34 net22 VDD VSS inv4
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/pfd_cp_lpf_lvs.sym # of pins=6
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/pfd_cp_lpf_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/pfd_cp_lpf_lvs.sch
.subckt pfd_cp_lpf_lvs  VDD VSS vsig_in ibiasn vcp vin_div
*.ipin VDD
*.ipin VSS
*.ipin vin_div
*.ipin vsig_in
*.opin vcp
*.ipin ibiasn
XM1 ibiasn ibiasn VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=10 m=10 
XM2 vpbias ibiasn VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 vswitchl ibiasn VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 vcp vQB vswitchl VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 vcp vQAb vswitchh VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM6 vswitchh vpbias VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM20 vpbias vpbias VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM21 vndiode vndiode VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM22 vndiode vQA vswitchh VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM23 vpdiode vpdiode VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM24 vpdiode vQBb vswitchl VSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
x7 vQA vQAb VDD VSS inv M=1
x8 vQB vQBb VDD VSS inv M=1
x12 vQA vRSTN vQB VDD VSS nand2 M=1
x1 vRSTN VDD vQA vsig_in net2 VDD VSS dffr_stdcell
x2 vRSTN VDD vQB vin_div net1 VDD VSS dffr_stdcell
XM7 vpbias VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM8 vswitchh VDD VDD VDD sky130_fd_pr__pfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM9 vswitchh VDD VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM11 vswitchh VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM10 vcp VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM12 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM13 vswitchl VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM14 vcp VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM15 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM17 ibiasn VSS VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM18 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM19 vpdiode VDD VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM25 vndiode VDD VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM26 vndiode VSS VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM27 vswitchl VSS VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM28 vpbias VSS VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM29 vswitchl VSS VSS VSS sky130_fd_pr__nfet_01v8 L=4 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM30 vpdiode VSS VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/latched_comparator_folded_lvs.sym # of pins=8
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/latched_comparator_folded_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/latched_comparator_folded_lvs.sch
.subckt latched_comparator_folded_lvs  vim vip vop vom ibiasp VDD VSS clk
*.ipin vip
*.ipin vim
*.opin vop
*.opin vom
*.ipin clk
*.ipin ibiasp
*.ipin VDD
*.ipin VSS
XM5 vcompm vcompp VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM11 vcompmb vcompm VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM13 vcomppb vcompp VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM15 vcomppb vcompp VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM6 vcompp vcompm VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM14 vlatchm vlatchp VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM3 vcompm clk VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7 vcompp clk VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM8 vop vcompm_buf VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM9 vop vom VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM18 nandm vcompm_buf VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM19 vop vom nandm VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM20 vom vop VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM21 vom vcompp_buf VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM22 nandp vcompp_buf VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM23 vom vop nandp VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM25 vcompm_buf vcompmb VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM26 vcompp_buf vcomppb VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM27 vcompp_buf vcomppb VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM4 ibiasp ibiasp VDD VDD sky130_fd_pr__pfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM2 vlatchm vip vtailp VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=8 m=8 
XM1 vlatchp vim vtailp VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=8 m=8 
XM32 vlatchp clk vlatchm VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=7 m=7 
XM16 vtailp ibiasp VDD VDD sky130_fd_pr__pfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM12 vlatchp vlatchm VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XM17 vcompp clk vlatchp VSS sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM28 vcompm clk vlatchm VSS sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM24 vcompm_buf vcompmb VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM10 vcompmb vcompm VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM29 vcompm VDD VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM30 vcompp VDD VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM31 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM33 vlatchp VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM34 vlatchm VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM35 vlatchp VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM36 vlatchm VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM37 vtailp vtailp vtailp VDD sky130_fd_pr__pfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM38 vlatchp VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM39 vlatchm VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/amux_2to1_lvs.sym # of pins=6
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/amux_2to1_lvs.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/amux_2to1_lvs.sch
.subckt amux_2to1_lvs  SEL A Y B VDD VSS
*.ipin A
*.ipin B
*.ipin SEL
*.opin Y
*.ipin VDD
*.ipin VSS
XM7 Y SELB A VDD sky130_fd_pr__pfet_01v8_hvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM8 A SEL Y VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM1 Y SEL B VDD sky130_fd_pr__pfet_01v8_hvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM2 B SELB Y VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
x1 SEL SELB VDD VSS inv1
XM3 B VSS VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM4 B VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM5 A VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt L=1 W=2 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/dff_stdcell.sym # of pins=6
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/dff_stdcell.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/dff_stdcell.sch
.subckt dff_stdcell  D Q CLK QB VDD VSS
*.ipin D
*.ipin CLK
*.opin Q
*.opin QB
*.ipin VDD
*.ipin VSS
x12 CLK D VSS VSS VDD VDD Q QB sky130_fd_sc_hd__dfxbp_1
**** begin user architecture code

.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/dfxbp/sky130_fd_sc_hd__dfxbp_1.spice

**** end user architecture code
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/and2.sym # of pins=5
* sym_path: /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/and2.sym
* sch_path: /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/and2.sch
.subckt and2  A Y B VDD VSS   M=1
*.ipin A
*.ipin B
*.opin Y
*.ipin VDD
*.ipin VSS
x1 A net1 B VDD VSS nand2 M=M
x2 net1 Y VDD VSS inv M=M
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/cs_ring_osc_stage_lvs_exp.sym # of pins=6
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/cs_ring_osc_stage_lvs_exp.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/cs_ring_osc_stage_lvs_exp.sch
.subckt cs_ring_osc_stage_lvs_exp  VDD vbiasp vout vin vbiasn VSS
*.opin vout
*.ipin vin
*.ipin vbiasn
*.ipin vbiasp
*.ipin VDD
*.ipin VSS
XM5 voutcs vin net1 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM1 csinvp vbiasp net2 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=2 m=2 
XC1 vout VSS sky130_fd_pr__cap_mim_m3_1 W=2 L=2 MF=9 m=9
XM3 net2 vbiasp net3 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM6 net3 vbiasp net4 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM9 net4 vbiasp net5 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM10 net5 vbiasp net6 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM11 net6 vbiasp net7 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM12 net7 vbiasp net8 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM13 net8 vbiasp VDD VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM14 voutcs vin net9 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM15 net9 vin net10 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM16 net10 vin net11 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM17 net11 vin net12 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM18 net12 vin net13 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM19 net13 vin net14 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM20 net14 vin net15 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM21 net15 vin csinvp VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM22 vout voutcs net16 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM23 net16 voutcs net17 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM24 net17 voutcs net18 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM25 net18 voutcs net19 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM26 net19 voutcs net20 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM27 net20 voutcs net21 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM28 net21 voutcs net22 VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29'
+ as='((3)/2) * 2 * 0.29' pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)'
+ nrd='1' nrs='1' sa=0 sb=0 sd=0 mult=1 m=1 
XM29 net22 voutcs VDD VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM30 net1 vin net23 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM31 net23 vin net24 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM32 net24 vin net25 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM33 net25 vin net26 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM34 net26 vin net27 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM35 net27 vin net28 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM36 net28 vin csinvn VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM37 csinvn vbiasn net29 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM38 net29 vbiasn net30 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM39 net30 vbiasn net31 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM40 net31 vbiasn net32 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM41 net32 vbiasn net33 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM42 net33 vbiasn net34 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM43 net34 vbiasn net35 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM44 net35 vbiasn VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM45 vout voutcs net36 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM46 net36 voutcs net37 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM47 net37 voutcs net38 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM48 net38 voutcs net39 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM49 net39 voutcs net40 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM50 net40 voutcs net41 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM51 net41 voutcs net42 VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM52 net42 voutcs VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XC2 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=2 L=2 MF=16 m=16
XM7 csinvn VSS VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM8 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM2 voutcs VSS VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM56 vout VSS VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 csinvp VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM53 voutcs VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM54 vout VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM55 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=6 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM57 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt L=2 W=8 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=2 m=2 
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/inv4.sym # of pins=4
* sym_path: /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/inv4.sym
* sch_path: /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/inv4.sch
.subckt inv4  A Y VDD VSS
*.ipin A
*.opin Y
*.ipin VDD
*.ipin VSS
XM2 Y A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM1 Y A VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=4 m=4 
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/inv.sym # of pins=4
* sym_path: /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/inv.sym
* sch_path: /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/inv.sch
.subckt inv  A Y VDD VSS   M=1
*.ipin A
*.opin Y
*.ipin VDD
*.ipin VSS
XM2 Y A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=M m=M 
XM1 Y A VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=M m=M 
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/nand2.sym # of pins=5
* sym_path: /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/nand2.sym
* sch_path: /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/nand2.sch
.subckt nand2  A Y B VDD VSS   M=1
*.ipin A
*.ipin B
*.opin Y
*.ipin VDD
*.ipin VSS
XM2 Y A net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=M m=M 
XM1 Y A VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=M m=M 
XM3 net1 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=M m=M 
XM4 Y B VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='((2)/2) * 2 * 0.29' as='((3)/2) * 2 * 0.29'
+ pd='2*((2)/2) * (2 + 0.29)' ps='2*((3)/2) * (2 + 0.29)' nrd='1' nrs='1'
+ sa=0 sb=0 sd=0 mult=M m=M 
.ends


* expanding   symbol:
*+  /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/dffr_stdcell.sym # of pins=7
* sym_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/dffr_stdcell.sym
* sch_path:
*+ /home/users/nhpoole/ee272b/ee272b_mixed_signal_mmwave_accelerator/designs/dffr_stdcell.sch
.subckt dffr_stdcell  RN D Q CLK QB VDD VSS
*.ipin D
*.ipin CLK
*.opin Q
*.opin QB
*.ipin RN
*.ipin VDD
*.ipin VSS
x1 CLK D RN VSS VSS VDD VDD Q QB sky130_fd_sc_hd__dfrbp_1
**** begin user architecture code

.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/dfrbp/sky130_fd_sc_hd__dfrbp_1.spice

**** end user architecture code
.ends

** flattened .save nodes
.end
