magic
tech sky130A
magscale 1 2
timestamp 1620680478
<< pwell >>
rect -3221 -510 3221 510
<< nmos >>
rect -3025 -300 -2065 300
rect -2007 -300 -1047 300
rect -989 -300 -29 300
rect 29 -300 989 300
rect 1047 -300 2007 300
rect 2065 -300 3025 300
<< ndiff >>
rect -3083 288 -3025 300
rect -3083 -288 -3071 288
rect -3037 -288 -3025 288
rect -3083 -300 -3025 -288
rect -2065 288 -2007 300
rect -2065 -288 -2053 288
rect -2019 -288 -2007 288
rect -2065 -300 -2007 -288
rect -1047 288 -989 300
rect -1047 -288 -1035 288
rect -1001 -288 -989 288
rect -1047 -300 -989 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 989 288 1047 300
rect 989 -288 1001 288
rect 1035 -288 1047 288
rect 989 -300 1047 -288
rect 2007 288 2065 300
rect 2007 -288 2019 288
rect 2053 -288 2065 288
rect 2007 -300 2065 -288
rect 3025 288 3083 300
rect 3025 -288 3037 288
rect 3071 -288 3083 288
rect 3025 -300 3083 -288
<< ndiffc >>
rect -3071 -288 -3037 288
rect -2053 -288 -2019 288
rect -1035 -288 -1001 288
rect -17 -288 17 288
rect 1001 -288 1035 288
rect 2019 -288 2053 288
rect 3037 -288 3071 288
<< psubdiff >>
rect -3185 440 -3089 474
rect 3089 440 3185 474
rect -3185 378 -3151 440
rect 3151 378 3185 440
rect -3185 -440 -3151 -378
rect 3151 -440 3185 -378
rect -3185 -474 -3089 -440
rect 3089 -474 3185 -440
<< psubdiffcont >>
rect -3089 440 3089 474
rect -3185 -378 -3151 378
rect 3151 -378 3185 378
rect -3089 -474 3089 -440
<< poly >>
rect -2839 372 -2251 388
rect -2839 355 -2823 372
rect -3025 338 -2823 355
rect -2267 355 -2251 372
rect -1821 372 -1233 388
rect -1821 355 -1805 372
rect -2267 338 -2065 355
rect -3025 300 -2065 338
rect -2007 338 -1805 355
rect -1249 355 -1233 372
rect -803 372 -215 388
rect -803 355 -787 372
rect -1249 338 -1047 355
rect -2007 300 -1047 338
rect -989 338 -787 355
rect -231 355 -215 372
rect 215 372 803 388
rect 215 355 231 372
rect -231 338 -29 355
rect -989 300 -29 338
rect 29 338 231 355
rect 787 355 803 372
rect 1233 372 1821 388
rect 1233 355 1249 372
rect 787 338 989 355
rect 29 300 989 338
rect 1047 338 1249 355
rect 1805 355 1821 372
rect 2251 372 2839 388
rect 2251 355 2267 372
rect 1805 338 2007 355
rect 1047 300 2007 338
rect 2065 338 2267 355
rect 2823 355 2839 372
rect 2823 338 3025 355
rect 2065 300 3025 338
rect -3025 -338 -2065 -300
rect -3025 -355 -2823 -338
rect -2839 -372 -2823 -355
rect -2267 -355 -2065 -338
rect -2007 -338 -1047 -300
rect -2007 -355 -1805 -338
rect -2267 -372 -2251 -355
rect -2839 -388 -2251 -372
rect -1821 -372 -1805 -355
rect -1249 -355 -1047 -338
rect -989 -338 -29 -300
rect -989 -355 -787 -338
rect -1249 -372 -1233 -355
rect -1821 -388 -1233 -372
rect -803 -372 -787 -355
rect -231 -355 -29 -338
rect 29 -338 989 -300
rect 29 -355 231 -338
rect -231 -372 -215 -355
rect -803 -388 -215 -372
rect 215 -372 231 -355
rect 787 -355 989 -338
rect 1047 -338 2007 -300
rect 1047 -355 1249 -338
rect 787 -372 803 -355
rect 215 -388 803 -372
rect 1233 -372 1249 -355
rect 1805 -355 2007 -338
rect 2065 -338 3025 -300
rect 2065 -355 2267 -338
rect 1805 -372 1821 -355
rect 1233 -388 1821 -372
rect 2251 -372 2267 -355
rect 2823 -355 3025 -338
rect 2823 -372 2839 -355
rect 2251 -388 2839 -372
<< polycont >>
rect -2823 338 -2267 372
rect -1805 338 -1249 372
rect -787 338 -231 372
rect 231 338 787 372
rect 1249 338 1805 372
rect 2267 338 2823 372
rect -2823 -372 -2267 -338
rect -1805 -372 -1249 -338
rect -787 -372 -231 -338
rect 231 -372 787 -338
rect 1249 -372 1805 -338
rect 2267 -372 2823 -338
<< locali >>
rect -3185 440 -3089 474
rect 3089 440 3185 474
rect -3185 378 -3151 440
rect 3151 378 3185 440
rect -2839 338 -2823 372
rect -2267 338 -2251 372
rect -1821 338 -1805 372
rect -1249 338 -1233 372
rect -803 338 -787 372
rect -231 338 -215 372
rect 215 338 231 372
rect 787 338 803 372
rect 1233 338 1249 372
rect 1805 338 1821 372
rect 2251 338 2267 372
rect 2823 338 2839 372
rect -3071 288 -3037 304
rect -3071 -304 -3037 -288
rect -2053 288 -2019 304
rect -2053 -304 -2019 -288
rect -1035 288 -1001 304
rect -1035 -304 -1001 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 1001 288 1035 304
rect 1001 -304 1035 -288
rect 2019 288 2053 304
rect 2019 -304 2053 -288
rect 3037 288 3071 304
rect 3037 -304 3071 -288
rect -2839 -372 -2823 -338
rect -2267 -372 -2251 -338
rect -1821 -372 -1805 -338
rect -1249 -372 -1233 -338
rect -803 -372 -787 -338
rect -231 -372 -215 -338
rect 215 -372 231 -338
rect 787 -372 803 -338
rect 1233 -372 1249 -338
rect 1805 -372 1821 -338
rect 2251 -372 2267 -338
rect 2823 -372 2839 -338
rect -3185 -440 -3151 -378
rect 3151 -440 3185 -378
rect -3185 -474 -3089 -440
rect 3089 -474 3185 -440
<< viali >>
rect -2777 338 -2313 372
rect -1759 338 -1295 372
rect -741 338 -277 372
rect 277 338 741 372
rect 1295 338 1759 372
rect 2313 338 2777 372
rect -3071 -288 -3037 288
rect -2053 -288 -2019 288
rect -1035 -288 -1001 288
rect -17 -288 17 288
rect 1001 -288 1035 288
rect 2019 -288 2053 288
rect 3037 -288 3071 288
rect -2777 -372 -2313 -338
rect -1759 -372 -1295 -338
rect -741 -372 -277 -338
rect 277 -372 741 -338
rect 1295 -372 1759 -338
rect 2313 -372 2777 -338
<< metal1 >>
rect -2789 372 -2301 378
rect -2789 338 -2777 372
rect -2313 338 -2301 372
rect -2789 332 -2301 338
rect -1771 372 -1283 378
rect -1771 338 -1759 372
rect -1295 338 -1283 372
rect -1771 332 -1283 338
rect -753 372 -265 378
rect -753 338 -741 372
rect -277 338 -265 372
rect -753 332 -265 338
rect 265 372 753 378
rect 265 338 277 372
rect 741 338 753 372
rect 265 332 753 338
rect 1283 372 1771 378
rect 1283 338 1295 372
rect 1759 338 1771 372
rect 1283 332 1771 338
rect 2301 372 2789 378
rect 2301 338 2313 372
rect 2777 338 2789 372
rect 2301 332 2789 338
rect -3077 288 -3031 300
rect -3077 -288 -3071 288
rect -3037 -288 -3031 288
rect -3077 -300 -3031 -288
rect -2059 288 -2013 300
rect -2059 -288 -2053 288
rect -2019 -288 -2013 288
rect -2059 -300 -2013 -288
rect -1041 288 -995 300
rect -1041 -288 -1035 288
rect -1001 -288 -995 288
rect -1041 -300 -995 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 995 288 1041 300
rect 995 -288 1001 288
rect 1035 -288 1041 288
rect 995 -300 1041 -288
rect 2013 288 2059 300
rect 2013 -288 2019 288
rect 2053 -288 2059 288
rect 2013 -300 2059 -288
rect 3031 288 3077 300
rect 3031 -288 3037 288
rect 3071 -288 3077 288
rect 3031 -300 3077 -288
rect -2789 -338 -2301 -332
rect -2789 -372 -2777 -338
rect -2313 -372 -2301 -338
rect -2789 -378 -2301 -372
rect -1771 -338 -1283 -332
rect -1771 -372 -1759 -338
rect -1295 -372 -1283 -338
rect -1771 -378 -1283 -372
rect -753 -338 -265 -332
rect -753 -372 -741 -338
rect -277 -372 -265 -338
rect -753 -378 -265 -372
rect 265 -338 753 -332
rect 265 -372 277 -338
rect 741 -372 753 -338
rect 265 -378 753 -372
rect 1283 -338 1771 -332
rect 1283 -372 1295 -338
rect 1759 -372 1771 -338
rect 1283 -378 1771 -372
rect 2301 -338 2789 -332
rect 2301 -372 2313 -338
rect 2777 -372 2789 -338
rect 2301 -378 2789 -372
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -3168 -457 3168 457
string parameters w 3 l 4.8 m 1 nf 6 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
