magic
tech sky130A
magscale 1 2
timestamp 1623661481
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 29 -17 63 17
<< locali >>
rect 21 199 89 391
rect 359 324 431 475
rect 467 357 527 475
rect 359 199 393 324
rect 467 290 505 357
rect 679 325 729 493
rect 847 325 897 493
rect 439 199 505 290
rect 551 289 638 323
rect 679 291 993 325
rect 551 199 585 289
rect 945 181 993 291
rect 687 145 993 181
rect 687 51 737 145
rect 839 51 905 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 17 427 73 527
rect 119 413 157 491
rect 123 265 157 413
rect 207 349 273 490
rect 207 315 325 349
rect 123 199 243 265
rect 123 181 157 199
rect 17 17 69 165
rect 119 87 157 181
rect 291 165 325 315
rect 584 359 634 527
rect 763 359 813 527
rect 931 359 981 527
rect 619 215 911 249
rect 619 165 653 215
rect 291 131 653 165
rect 207 17 257 117
rect 323 61 357 131
rect 397 17 463 97
rect 497 61 531 131
rect 575 17 651 97
rect 771 17 805 111
rect 939 17 973 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel locali s 551 289 638 323 6 A
port 1 nsew signal input
rlabel locali s 551 199 585 289 6 A
port 1 nsew signal input
rlabel locali s 467 357 527 475 6 B
port 2 nsew signal input
rlabel locali s 467 290 505 357 6 B
port 2 nsew signal input
rlabel locali s 439 199 505 290 6 B
port 2 nsew signal input
rlabel locali s 359 324 431 475 6 C
port 3 nsew signal input
rlabel locali s 359 199 393 324 6 C
port 3 nsew signal input
rlabel locali s 21 199 89 391 6 D_N
port 4 nsew signal input
rlabel locali s 945 181 993 291 6 X
port 5 nsew signal output
rlabel locali s 847 325 897 493 6 X
port 5 nsew signal output
rlabel locali s 839 51 905 145 6 X
port 5 nsew signal output
rlabel locali s 687 145 993 181 6 X
port 5 nsew signal output
rlabel locali s 687 51 737 145 6 X
port 5 nsew signal output
rlabel locali s 679 325 729 493 6 X
port 5 nsew signal output
rlabel locali s 679 291 993 325 6 X
port 5 nsew signal output
rlabel metal1 s 0 -48 1012 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 1050 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 1012 592 6 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
