magic
tech sky130A
magscale 1 2
timestamp 1621486730
<< pwell >>
rect -1457 -310 1457 310
<< nmos >>
rect -1261 -100 -1061 100
rect -1003 -100 -803 100
rect -745 -100 -545 100
rect -487 -100 -287 100
rect -229 -100 -29 100
rect 29 -100 229 100
rect 287 -100 487 100
rect 545 -100 745 100
rect 803 -100 1003 100
rect 1061 -100 1261 100
<< ndiff >>
rect -1319 88 -1261 100
rect -1319 -88 -1307 88
rect -1273 -88 -1261 88
rect -1319 -100 -1261 -88
rect -1061 88 -1003 100
rect -1061 -88 -1049 88
rect -1015 -88 -1003 88
rect -1061 -100 -1003 -88
rect -803 88 -745 100
rect -803 -88 -791 88
rect -757 -88 -745 88
rect -803 -100 -745 -88
rect -545 88 -487 100
rect -545 -88 -533 88
rect -499 -88 -487 88
rect -545 -100 -487 -88
rect -287 88 -229 100
rect -287 -88 -275 88
rect -241 -88 -229 88
rect -287 -100 -229 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 229 88 287 100
rect 229 -88 241 88
rect 275 -88 287 88
rect 229 -100 287 -88
rect 487 88 545 100
rect 487 -88 499 88
rect 533 -88 545 88
rect 487 -100 545 -88
rect 745 88 803 100
rect 745 -88 757 88
rect 791 -88 803 88
rect 745 -100 803 -88
rect 1003 88 1061 100
rect 1003 -88 1015 88
rect 1049 -88 1061 88
rect 1003 -100 1061 -88
rect 1261 88 1319 100
rect 1261 -88 1273 88
rect 1307 -88 1319 88
rect 1261 -100 1319 -88
<< ndiffc >>
rect -1307 -88 -1273 88
rect -1049 -88 -1015 88
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
rect 1015 -88 1049 88
rect 1273 -88 1307 88
<< psubdiff >>
rect -1421 240 -1325 274
rect 1325 240 1421 274
rect -1421 178 -1387 240
rect 1387 178 1421 240
rect -1421 -240 -1387 -178
rect 1387 -240 1421 -178
rect -1421 -274 -1325 -240
rect 1325 -274 1421 -240
<< psubdiffcont >>
rect -1325 240 1325 274
rect -1421 -178 -1387 178
rect 1387 -178 1421 178
rect -1325 -274 1325 -240
<< poly >>
rect -1227 172 -1095 188
rect -1227 155 -1211 172
rect -1261 138 -1211 155
rect -1111 155 -1095 172
rect -969 172 -837 188
rect -969 155 -953 172
rect -1111 138 -1061 155
rect -1261 100 -1061 138
rect -1003 138 -953 155
rect -853 155 -837 172
rect -711 172 -579 188
rect -711 155 -695 172
rect -853 138 -803 155
rect -1003 100 -803 138
rect -745 138 -695 155
rect -595 155 -579 172
rect -453 172 -321 188
rect -453 155 -437 172
rect -595 138 -545 155
rect -745 100 -545 138
rect -487 138 -437 155
rect -337 155 -321 172
rect -195 172 -63 188
rect -195 155 -179 172
rect -337 138 -287 155
rect -487 100 -287 138
rect -229 138 -179 155
rect -79 155 -63 172
rect 63 172 195 188
rect 63 155 79 172
rect -79 138 -29 155
rect -229 100 -29 138
rect 29 138 79 155
rect 179 155 195 172
rect 321 172 453 188
rect 321 155 337 172
rect 179 138 229 155
rect 29 100 229 138
rect 287 138 337 155
rect 437 155 453 172
rect 579 172 711 188
rect 579 155 595 172
rect 437 138 487 155
rect 287 100 487 138
rect 545 138 595 155
rect 695 155 711 172
rect 837 172 969 188
rect 837 155 853 172
rect 695 138 745 155
rect 545 100 745 138
rect 803 138 853 155
rect 953 155 969 172
rect 1095 172 1227 188
rect 1095 155 1111 172
rect 953 138 1003 155
rect 803 100 1003 138
rect 1061 138 1111 155
rect 1211 155 1227 172
rect 1211 138 1261 155
rect 1061 100 1261 138
rect -1261 -138 -1061 -100
rect -1261 -155 -1211 -138
rect -1227 -172 -1211 -155
rect -1111 -155 -1061 -138
rect -1003 -138 -803 -100
rect -1003 -155 -953 -138
rect -1111 -172 -1095 -155
rect -1227 -188 -1095 -172
rect -969 -172 -953 -155
rect -853 -155 -803 -138
rect -745 -138 -545 -100
rect -745 -155 -695 -138
rect -853 -172 -837 -155
rect -969 -188 -837 -172
rect -711 -172 -695 -155
rect -595 -155 -545 -138
rect -487 -138 -287 -100
rect -487 -155 -437 -138
rect -595 -172 -579 -155
rect -711 -188 -579 -172
rect -453 -172 -437 -155
rect -337 -155 -287 -138
rect -229 -138 -29 -100
rect -229 -155 -179 -138
rect -337 -172 -321 -155
rect -453 -188 -321 -172
rect -195 -172 -179 -155
rect -79 -155 -29 -138
rect 29 -138 229 -100
rect 29 -155 79 -138
rect -79 -172 -63 -155
rect -195 -188 -63 -172
rect 63 -172 79 -155
rect 179 -155 229 -138
rect 287 -138 487 -100
rect 287 -155 337 -138
rect 179 -172 195 -155
rect 63 -188 195 -172
rect 321 -172 337 -155
rect 437 -155 487 -138
rect 545 -138 745 -100
rect 545 -155 595 -138
rect 437 -172 453 -155
rect 321 -188 453 -172
rect 579 -172 595 -155
rect 695 -155 745 -138
rect 803 -138 1003 -100
rect 803 -155 853 -138
rect 695 -172 711 -155
rect 579 -188 711 -172
rect 837 -172 853 -155
rect 953 -155 1003 -138
rect 1061 -138 1261 -100
rect 1061 -155 1111 -138
rect 953 -172 969 -155
rect 837 -188 969 -172
rect 1095 -172 1111 -155
rect 1211 -155 1261 -138
rect 1211 -172 1227 -155
rect 1095 -188 1227 -172
<< polycont >>
rect -1211 138 -1111 172
rect -953 138 -853 172
rect -695 138 -595 172
rect -437 138 -337 172
rect -179 138 -79 172
rect 79 138 179 172
rect 337 138 437 172
rect 595 138 695 172
rect 853 138 953 172
rect 1111 138 1211 172
rect -1211 -172 -1111 -138
rect -953 -172 -853 -138
rect -695 -172 -595 -138
rect -437 -172 -337 -138
rect -179 -172 -79 -138
rect 79 -172 179 -138
rect 337 -172 437 -138
rect 595 -172 695 -138
rect 853 -172 953 -138
rect 1111 -172 1211 -138
<< locali >>
rect -1421 240 -1325 274
rect 1325 240 1421 274
rect -1421 178 -1387 240
rect 1387 178 1421 240
rect -1227 138 -1211 172
rect -1111 138 -1095 172
rect -969 138 -953 172
rect -853 138 -837 172
rect -711 138 -695 172
rect -595 138 -579 172
rect -453 138 -437 172
rect -337 138 -321 172
rect -195 138 -179 172
rect -79 138 -63 172
rect 63 138 79 172
rect 179 138 195 172
rect 321 138 337 172
rect 437 138 453 172
rect 579 138 595 172
rect 695 138 711 172
rect 837 138 853 172
rect 953 138 969 172
rect 1095 138 1111 172
rect 1211 138 1227 172
rect -1307 88 -1273 104
rect -1307 -104 -1273 -88
rect -1049 88 -1015 104
rect -1049 -104 -1015 -88
rect -791 88 -757 104
rect -791 -104 -757 -88
rect -533 88 -499 104
rect -533 -104 -499 -88
rect -275 88 -241 104
rect -275 -104 -241 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 241 88 275 104
rect 241 -104 275 -88
rect 499 88 533 104
rect 499 -104 533 -88
rect 757 88 791 104
rect 757 -104 791 -88
rect 1015 88 1049 104
rect 1015 -104 1049 -88
rect 1273 88 1307 104
rect 1273 -104 1307 -88
rect -1227 -172 -1211 -138
rect -1111 -172 -1095 -138
rect -969 -172 -953 -138
rect -853 -172 -837 -138
rect -711 -172 -695 -138
rect -595 -172 -579 -138
rect -453 -172 -437 -138
rect -337 -172 -321 -138
rect -195 -172 -179 -138
rect -79 -172 -63 -138
rect 63 -172 79 -138
rect 179 -172 195 -138
rect 321 -172 337 -138
rect 437 -172 453 -138
rect 579 -172 595 -138
rect 695 -172 711 -138
rect 837 -172 853 -138
rect 953 -172 969 -138
rect 1095 -172 1111 -138
rect 1211 -172 1227 -138
rect -1421 -240 -1387 -178
rect 1387 -240 1421 -178
rect -1421 -274 -1325 -240
rect 1325 -274 1421 -240
<< viali >>
rect -1203 138 -1119 172
rect -945 138 -861 172
rect -687 138 -603 172
rect -429 138 -345 172
rect -171 138 -87 172
rect 87 138 171 172
rect 345 138 429 172
rect 603 138 687 172
rect 861 138 945 172
rect 1119 138 1203 172
rect -1307 -88 -1273 88
rect -1049 -88 -1015 88
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
rect 1015 -88 1049 88
rect 1273 -88 1307 88
rect -1203 -172 -1119 -138
rect -945 -172 -861 -138
rect -687 -172 -603 -138
rect -429 -172 -345 -138
rect -171 -172 -87 -138
rect 87 -172 171 -138
rect 345 -172 429 -138
rect 603 -172 687 -138
rect 861 -172 945 -138
rect 1119 -172 1203 -138
<< metal1 >>
rect -1215 172 -1107 178
rect -1215 138 -1203 172
rect -1119 138 -1107 172
rect -1215 132 -1107 138
rect -957 172 -849 178
rect -957 138 -945 172
rect -861 138 -849 172
rect -957 132 -849 138
rect -699 172 -591 178
rect -699 138 -687 172
rect -603 138 -591 172
rect -699 132 -591 138
rect -441 172 -333 178
rect -441 138 -429 172
rect -345 138 -333 172
rect -441 132 -333 138
rect -183 172 -75 178
rect -183 138 -171 172
rect -87 138 -75 172
rect -183 132 -75 138
rect 75 172 183 178
rect 75 138 87 172
rect 171 138 183 172
rect 75 132 183 138
rect 333 172 441 178
rect 333 138 345 172
rect 429 138 441 172
rect 333 132 441 138
rect 591 172 699 178
rect 591 138 603 172
rect 687 138 699 172
rect 591 132 699 138
rect 849 172 957 178
rect 849 138 861 172
rect 945 138 957 172
rect 849 132 957 138
rect 1107 172 1215 178
rect 1107 138 1119 172
rect 1203 138 1215 172
rect 1107 132 1215 138
rect -1313 88 -1267 100
rect -1313 -88 -1307 88
rect -1273 -88 -1267 88
rect -1313 -100 -1267 -88
rect -1055 88 -1009 100
rect -1055 -88 -1049 88
rect -1015 -88 -1009 88
rect -1055 -100 -1009 -88
rect -797 88 -751 100
rect -797 -88 -791 88
rect -757 -88 -751 88
rect -797 -100 -751 -88
rect -539 88 -493 100
rect -539 -88 -533 88
rect -499 -88 -493 88
rect -539 -100 -493 -88
rect -281 88 -235 100
rect -281 -88 -275 88
rect -241 -88 -235 88
rect -281 -100 -235 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 235 88 281 100
rect 235 -88 241 88
rect 275 -88 281 88
rect 235 -100 281 -88
rect 493 88 539 100
rect 493 -88 499 88
rect 533 -88 539 88
rect 493 -100 539 -88
rect 751 88 797 100
rect 751 -88 757 88
rect 791 -88 797 88
rect 751 -100 797 -88
rect 1009 88 1055 100
rect 1009 -88 1015 88
rect 1049 -88 1055 88
rect 1009 -100 1055 -88
rect 1267 88 1313 100
rect 1267 -88 1273 88
rect 1307 -88 1313 88
rect 1267 -100 1313 -88
rect -1215 -138 -1107 -132
rect -1215 -172 -1203 -138
rect -1119 -172 -1107 -138
rect -1215 -178 -1107 -172
rect -957 -138 -849 -132
rect -957 -172 -945 -138
rect -861 -172 -849 -138
rect -957 -178 -849 -172
rect -699 -138 -591 -132
rect -699 -172 -687 -138
rect -603 -172 -591 -138
rect -699 -178 -591 -172
rect -441 -138 -333 -132
rect -441 -172 -429 -138
rect -345 -172 -333 -138
rect -441 -178 -333 -172
rect -183 -138 -75 -132
rect -183 -172 -171 -138
rect -87 -172 -75 -138
rect -183 -178 -75 -172
rect 75 -138 183 -132
rect 75 -172 87 -138
rect 171 -172 183 -138
rect 75 -178 183 -172
rect 333 -138 441 -132
rect 333 -172 345 -138
rect 429 -172 441 -138
rect 333 -178 441 -172
rect 591 -138 699 -132
rect 591 -172 603 -138
rect 687 -172 699 -138
rect 591 -178 699 -172
rect 849 -138 957 -132
rect 849 -172 861 -138
rect 945 -172 957 -138
rect 849 -178 957 -172
rect 1107 -138 1215 -132
rect 1107 -172 1119 -138
rect 1203 -172 1215 -138
rect 1107 -178 1215 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1404 -257 1404 257
string parameters w 1 l 1 m 1 nf 10 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
