magic
tech sky130A
timestamp 1625948044
<< metal1 >>
rect -61 13 61 24
rect -35 -13 -29 13
rect -3 -13 3 13
rect 29 -13 35 13
rect -61 -24 61 -13
<< via1 >>
rect -61 -13 -35 13
rect -29 -13 -3 13
rect 3 -13 29 13
rect 35 -13 61 13
<< metal2 >>
rect -61 13 61 24
rect -35 -13 -29 13
rect -3 -13 3 13
rect 29 -13 35 13
rect -61 -24 61 -13
<< end >>
