magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -3889 -1657 3889 1657
<< pwell >>
rect -2629 -335 2629 335
<< nmos >>
rect -2545 109 -1745 309
rect -1687 109 -887 309
rect -829 109 -29 309
rect 29 109 829 309
rect 887 109 1687 309
rect 1745 109 2545 309
rect -2545 -309 -1745 -109
rect -1687 -309 -887 -109
rect -829 -309 -29 -109
rect 29 -309 829 -109
rect 887 -309 1687 -109
rect 1745 -309 2545 -109
<< ndiff >>
rect -2603 294 -2545 309
rect -2603 260 -2591 294
rect -2557 260 -2545 294
rect -2603 226 -2545 260
rect -2603 192 -2591 226
rect -2557 192 -2545 226
rect -2603 158 -2545 192
rect -2603 124 -2591 158
rect -2557 124 -2545 158
rect -2603 109 -2545 124
rect -1745 294 -1687 309
rect -1745 260 -1733 294
rect -1699 260 -1687 294
rect -1745 226 -1687 260
rect -1745 192 -1733 226
rect -1699 192 -1687 226
rect -1745 158 -1687 192
rect -1745 124 -1733 158
rect -1699 124 -1687 158
rect -1745 109 -1687 124
rect -887 294 -829 309
rect -887 260 -875 294
rect -841 260 -829 294
rect -887 226 -829 260
rect -887 192 -875 226
rect -841 192 -829 226
rect -887 158 -829 192
rect -887 124 -875 158
rect -841 124 -829 158
rect -887 109 -829 124
rect -29 294 29 309
rect -29 260 -17 294
rect 17 260 29 294
rect -29 226 29 260
rect -29 192 -17 226
rect 17 192 29 226
rect -29 158 29 192
rect -29 124 -17 158
rect 17 124 29 158
rect -29 109 29 124
rect 829 294 887 309
rect 829 260 841 294
rect 875 260 887 294
rect 829 226 887 260
rect 829 192 841 226
rect 875 192 887 226
rect 829 158 887 192
rect 829 124 841 158
rect 875 124 887 158
rect 829 109 887 124
rect 1687 294 1745 309
rect 1687 260 1699 294
rect 1733 260 1745 294
rect 1687 226 1745 260
rect 1687 192 1699 226
rect 1733 192 1745 226
rect 1687 158 1745 192
rect 1687 124 1699 158
rect 1733 124 1745 158
rect 1687 109 1745 124
rect 2545 294 2603 309
rect 2545 260 2557 294
rect 2591 260 2603 294
rect 2545 226 2603 260
rect 2545 192 2557 226
rect 2591 192 2603 226
rect 2545 158 2603 192
rect 2545 124 2557 158
rect 2591 124 2603 158
rect 2545 109 2603 124
rect -2603 -124 -2545 -109
rect -2603 -158 -2591 -124
rect -2557 -158 -2545 -124
rect -2603 -192 -2545 -158
rect -2603 -226 -2591 -192
rect -2557 -226 -2545 -192
rect -2603 -260 -2545 -226
rect -2603 -294 -2591 -260
rect -2557 -294 -2545 -260
rect -2603 -309 -2545 -294
rect -1745 -124 -1687 -109
rect -1745 -158 -1733 -124
rect -1699 -158 -1687 -124
rect -1745 -192 -1687 -158
rect -1745 -226 -1733 -192
rect -1699 -226 -1687 -192
rect -1745 -260 -1687 -226
rect -1745 -294 -1733 -260
rect -1699 -294 -1687 -260
rect -1745 -309 -1687 -294
rect -887 -124 -829 -109
rect -887 -158 -875 -124
rect -841 -158 -829 -124
rect -887 -192 -829 -158
rect -887 -226 -875 -192
rect -841 -226 -829 -192
rect -887 -260 -829 -226
rect -887 -294 -875 -260
rect -841 -294 -829 -260
rect -887 -309 -829 -294
rect -29 -124 29 -109
rect -29 -158 -17 -124
rect 17 -158 29 -124
rect -29 -192 29 -158
rect -29 -226 -17 -192
rect 17 -226 29 -192
rect -29 -260 29 -226
rect -29 -294 -17 -260
rect 17 -294 29 -260
rect -29 -309 29 -294
rect 829 -124 887 -109
rect 829 -158 841 -124
rect 875 -158 887 -124
rect 829 -192 887 -158
rect 829 -226 841 -192
rect 875 -226 887 -192
rect 829 -260 887 -226
rect 829 -294 841 -260
rect 875 -294 887 -260
rect 829 -309 887 -294
rect 1687 -124 1745 -109
rect 1687 -158 1699 -124
rect 1733 -158 1745 -124
rect 1687 -192 1745 -158
rect 1687 -226 1699 -192
rect 1733 -226 1745 -192
rect 1687 -260 1745 -226
rect 1687 -294 1699 -260
rect 1733 -294 1745 -260
rect 1687 -309 1745 -294
rect 2545 -124 2603 -109
rect 2545 -158 2557 -124
rect 2591 -158 2603 -124
rect 2545 -192 2603 -158
rect 2545 -226 2557 -192
rect 2591 -226 2603 -192
rect 2545 -260 2603 -226
rect 2545 -294 2557 -260
rect 2591 -294 2603 -260
rect 2545 -309 2603 -294
<< ndiffc >>
rect -2591 260 -2557 294
rect -2591 192 -2557 226
rect -2591 124 -2557 158
rect -1733 260 -1699 294
rect -1733 192 -1699 226
rect -1733 124 -1699 158
rect -875 260 -841 294
rect -875 192 -841 226
rect -875 124 -841 158
rect -17 260 17 294
rect -17 192 17 226
rect -17 124 17 158
rect 841 260 875 294
rect 841 192 875 226
rect 841 124 875 158
rect 1699 260 1733 294
rect 1699 192 1733 226
rect 1699 124 1733 158
rect 2557 260 2591 294
rect 2557 192 2591 226
rect 2557 124 2591 158
rect -2591 -158 -2557 -124
rect -2591 -226 -2557 -192
rect -2591 -294 -2557 -260
rect -1733 -158 -1699 -124
rect -1733 -226 -1699 -192
rect -1733 -294 -1699 -260
rect -875 -158 -841 -124
rect -875 -226 -841 -192
rect -875 -294 -841 -260
rect -17 -158 17 -124
rect -17 -226 17 -192
rect -17 -294 17 -260
rect 841 -158 875 -124
rect 841 -226 875 -192
rect 841 -294 875 -260
rect 1699 -158 1733 -124
rect 1699 -226 1733 -192
rect 1699 -294 1733 -260
rect 2557 -158 2591 -124
rect 2557 -226 2591 -192
rect 2557 -294 2591 -260
<< poly >>
rect -2391 381 -1899 397
rect -2391 364 -2366 381
rect -2545 347 -2366 364
rect -2332 347 -2298 381
rect -2264 347 -2230 381
rect -2196 347 -2162 381
rect -2128 347 -2094 381
rect -2060 347 -2026 381
rect -1992 347 -1958 381
rect -1924 364 -1899 381
rect -1533 381 -1041 397
rect -1533 364 -1508 381
rect -1924 347 -1745 364
rect -2545 309 -1745 347
rect -1687 347 -1508 364
rect -1474 347 -1440 381
rect -1406 347 -1372 381
rect -1338 347 -1304 381
rect -1270 347 -1236 381
rect -1202 347 -1168 381
rect -1134 347 -1100 381
rect -1066 364 -1041 381
rect -675 381 -183 397
rect -675 364 -650 381
rect -1066 347 -887 364
rect -1687 309 -887 347
rect -829 347 -650 364
rect -616 347 -582 381
rect -548 347 -514 381
rect -480 347 -446 381
rect -412 347 -378 381
rect -344 347 -310 381
rect -276 347 -242 381
rect -208 364 -183 381
rect 183 381 675 397
rect 183 364 208 381
rect -208 347 -29 364
rect -829 309 -29 347
rect 29 347 208 364
rect 242 347 276 381
rect 310 347 344 381
rect 378 347 412 381
rect 446 347 480 381
rect 514 347 548 381
rect 582 347 616 381
rect 650 364 675 381
rect 1041 381 1533 397
rect 1041 364 1066 381
rect 650 347 829 364
rect 29 309 829 347
rect 887 347 1066 364
rect 1100 347 1134 381
rect 1168 347 1202 381
rect 1236 347 1270 381
rect 1304 347 1338 381
rect 1372 347 1406 381
rect 1440 347 1474 381
rect 1508 364 1533 381
rect 1899 381 2391 397
rect 1899 364 1924 381
rect 1508 347 1687 364
rect 887 309 1687 347
rect 1745 347 1924 364
rect 1958 347 1992 381
rect 2026 347 2060 381
rect 2094 347 2128 381
rect 2162 347 2196 381
rect 2230 347 2264 381
rect 2298 347 2332 381
rect 2366 364 2391 381
rect 2366 347 2545 364
rect 1745 309 2545 347
rect -2545 71 -1745 109
rect -2545 54 -2366 71
rect -2391 37 -2366 54
rect -2332 37 -2298 71
rect -2264 37 -2230 71
rect -2196 37 -2162 71
rect -2128 37 -2094 71
rect -2060 37 -2026 71
rect -1992 37 -1958 71
rect -1924 54 -1745 71
rect -1687 71 -887 109
rect -1687 54 -1508 71
rect -1924 37 -1899 54
rect -2391 21 -1899 37
rect -1533 37 -1508 54
rect -1474 37 -1440 71
rect -1406 37 -1372 71
rect -1338 37 -1304 71
rect -1270 37 -1236 71
rect -1202 37 -1168 71
rect -1134 37 -1100 71
rect -1066 54 -887 71
rect -829 71 -29 109
rect -829 54 -650 71
rect -1066 37 -1041 54
rect -1533 21 -1041 37
rect -675 37 -650 54
rect -616 37 -582 71
rect -548 37 -514 71
rect -480 37 -446 71
rect -412 37 -378 71
rect -344 37 -310 71
rect -276 37 -242 71
rect -208 54 -29 71
rect 29 71 829 109
rect 29 54 208 71
rect -208 37 -183 54
rect -675 21 -183 37
rect 183 37 208 54
rect 242 37 276 71
rect 310 37 344 71
rect 378 37 412 71
rect 446 37 480 71
rect 514 37 548 71
rect 582 37 616 71
rect 650 54 829 71
rect 887 71 1687 109
rect 887 54 1066 71
rect 650 37 675 54
rect 183 21 675 37
rect 1041 37 1066 54
rect 1100 37 1134 71
rect 1168 37 1202 71
rect 1236 37 1270 71
rect 1304 37 1338 71
rect 1372 37 1406 71
rect 1440 37 1474 71
rect 1508 54 1687 71
rect 1745 71 2545 109
rect 1745 54 1924 71
rect 1508 37 1533 54
rect 1041 21 1533 37
rect 1899 37 1924 54
rect 1958 37 1992 71
rect 2026 37 2060 71
rect 2094 37 2128 71
rect 2162 37 2196 71
rect 2230 37 2264 71
rect 2298 37 2332 71
rect 2366 54 2545 71
rect 2366 37 2391 54
rect 1899 21 2391 37
rect -2391 -37 -1899 -21
rect -2391 -54 -2366 -37
rect -2545 -71 -2366 -54
rect -2332 -71 -2298 -37
rect -2264 -71 -2230 -37
rect -2196 -71 -2162 -37
rect -2128 -71 -2094 -37
rect -2060 -71 -2026 -37
rect -1992 -71 -1958 -37
rect -1924 -54 -1899 -37
rect -1533 -37 -1041 -21
rect -1533 -54 -1508 -37
rect -1924 -71 -1745 -54
rect -2545 -109 -1745 -71
rect -1687 -71 -1508 -54
rect -1474 -71 -1440 -37
rect -1406 -71 -1372 -37
rect -1338 -71 -1304 -37
rect -1270 -71 -1236 -37
rect -1202 -71 -1168 -37
rect -1134 -71 -1100 -37
rect -1066 -54 -1041 -37
rect -675 -37 -183 -21
rect -675 -54 -650 -37
rect -1066 -71 -887 -54
rect -1687 -109 -887 -71
rect -829 -71 -650 -54
rect -616 -71 -582 -37
rect -548 -71 -514 -37
rect -480 -71 -446 -37
rect -412 -71 -378 -37
rect -344 -71 -310 -37
rect -276 -71 -242 -37
rect -208 -54 -183 -37
rect 183 -37 675 -21
rect 183 -54 208 -37
rect -208 -71 -29 -54
rect -829 -109 -29 -71
rect 29 -71 208 -54
rect 242 -71 276 -37
rect 310 -71 344 -37
rect 378 -71 412 -37
rect 446 -71 480 -37
rect 514 -71 548 -37
rect 582 -71 616 -37
rect 650 -54 675 -37
rect 1041 -37 1533 -21
rect 1041 -54 1066 -37
rect 650 -71 829 -54
rect 29 -109 829 -71
rect 887 -71 1066 -54
rect 1100 -71 1134 -37
rect 1168 -71 1202 -37
rect 1236 -71 1270 -37
rect 1304 -71 1338 -37
rect 1372 -71 1406 -37
rect 1440 -71 1474 -37
rect 1508 -54 1533 -37
rect 1899 -37 2391 -21
rect 1899 -54 1924 -37
rect 1508 -71 1687 -54
rect 887 -109 1687 -71
rect 1745 -71 1924 -54
rect 1958 -71 1992 -37
rect 2026 -71 2060 -37
rect 2094 -71 2128 -37
rect 2162 -71 2196 -37
rect 2230 -71 2264 -37
rect 2298 -71 2332 -37
rect 2366 -54 2391 -37
rect 2366 -71 2545 -54
rect 1745 -109 2545 -71
rect -2545 -347 -1745 -309
rect -2545 -364 -2366 -347
rect -2391 -381 -2366 -364
rect -2332 -381 -2298 -347
rect -2264 -381 -2230 -347
rect -2196 -381 -2162 -347
rect -2128 -381 -2094 -347
rect -2060 -381 -2026 -347
rect -1992 -381 -1958 -347
rect -1924 -364 -1745 -347
rect -1687 -347 -887 -309
rect -1687 -364 -1508 -347
rect -1924 -381 -1899 -364
rect -2391 -397 -1899 -381
rect -1533 -381 -1508 -364
rect -1474 -381 -1440 -347
rect -1406 -381 -1372 -347
rect -1338 -381 -1304 -347
rect -1270 -381 -1236 -347
rect -1202 -381 -1168 -347
rect -1134 -381 -1100 -347
rect -1066 -364 -887 -347
rect -829 -347 -29 -309
rect -829 -364 -650 -347
rect -1066 -381 -1041 -364
rect -1533 -397 -1041 -381
rect -675 -381 -650 -364
rect -616 -381 -582 -347
rect -548 -381 -514 -347
rect -480 -381 -446 -347
rect -412 -381 -378 -347
rect -344 -381 -310 -347
rect -276 -381 -242 -347
rect -208 -364 -29 -347
rect 29 -347 829 -309
rect 29 -364 208 -347
rect -208 -381 -183 -364
rect -675 -397 -183 -381
rect 183 -381 208 -364
rect 242 -381 276 -347
rect 310 -381 344 -347
rect 378 -381 412 -347
rect 446 -381 480 -347
rect 514 -381 548 -347
rect 582 -381 616 -347
rect 650 -364 829 -347
rect 887 -347 1687 -309
rect 887 -364 1066 -347
rect 650 -381 675 -364
rect 183 -397 675 -381
rect 1041 -381 1066 -364
rect 1100 -381 1134 -347
rect 1168 -381 1202 -347
rect 1236 -381 1270 -347
rect 1304 -381 1338 -347
rect 1372 -381 1406 -347
rect 1440 -381 1474 -347
rect 1508 -364 1687 -347
rect 1745 -347 2545 -309
rect 1745 -364 1924 -347
rect 1508 -381 1533 -364
rect 1041 -397 1533 -381
rect 1899 -381 1924 -364
rect 1958 -381 1992 -347
rect 2026 -381 2060 -347
rect 2094 -381 2128 -347
rect 2162 -381 2196 -347
rect 2230 -381 2264 -347
rect 2298 -381 2332 -347
rect 2366 -364 2545 -347
rect 2366 -381 2391 -364
rect 1899 -397 2391 -381
<< polycont >>
rect -2366 347 -2332 381
rect -2298 347 -2264 381
rect -2230 347 -2196 381
rect -2162 347 -2128 381
rect -2094 347 -2060 381
rect -2026 347 -1992 381
rect -1958 347 -1924 381
rect -1508 347 -1474 381
rect -1440 347 -1406 381
rect -1372 347 -1338 381
rect -1304 347 -1270 381
rect -1236 347 -1202 381
rect -1168 347 -1134 381
rect -1100 347 -1066 381
rect -650 347 -616 381
rect -582 347 -548 381
rect -514 347 -480 381
rect -446 347 -412 381
rect -378 347 -344 381
rect -310 347 -276 381
rect -242 347 -208 381
rect 208 347 242 381
rect 276 347 310 381
rect 344 347 378 381
rect 412 347 446 381
rect 480 347 514 381
rect 548 347 582 381
rect 616 347 650 381
rect 1066 347 1100 381
rect 1134 347 1168 381
rect 1202 347 1236 381
rect 1270 347 1304 381
rect 1338 347 1372 381
rect 1406 347 1440 381
rect 1474 347 1508 381
rect 1924 347 1958 381
rect 1992 347 2026 381
rect 2060 347 2094 381
rect 2128 347 2162 381
rect 2196 347 2230 381
rect 2264 347 2298 381
rect 2332 347 2366 381
rect -2366 37 -2332 71
rect -2298 37 -2264 71
rect -2230 37 -2196 71
rect -2162 37 -2128 71
rect -2094 37 -2060 71
rect -2026 37 -1992 71
rect -1958 37 -1924 71
rect -1508 37 -1474 71
rect -1440 37 -1406 71
rect -1372 37 -1338 71
rect -1304 37 -1270 71
rect -1236 37 -1202 71
rect -1168 37 -1134 71
rect -1100 37 -1066 71
rect -650 37 -616 71
rect -582 37 -548 71
rect -514 37 -480 71
rect -446 37 -412 71
rect -378 37 -344 71
rect -310 37 -276 71
rect -242 37 -208 71
rect 208 37 242 71
rect 276 37 310 71
rect 344 37 378 71
rect 412 37 446 71
rect 480 37 514 71
rect 548 37 582 71
rect 616 37 650 71
rect 1066 37 1100 71
rect 1134 37 1168 71
rect 1202 37 1236 71
rect 1270 37 1304 71
rect 1338 37 1372 71
rect 1406 37 1440 71
rect 1474 37 1508 71
rect 1924 37 1958 71
rect 1992 37 2026 71
rect 2060 37 2094 71
rect 2128 37 2162 71
rect 2196 37 2230 71
rect 2264 37 2298 71
rect 2332 37 2366 71
rect -2366 -71 -2332 -37
rect -2298 -71 -2264 -37
rect -2230 -71 -2196 -37
rect -2162 -71 -2128 -37
rect -2094 -71 -2060 -37
rect -2026 -71 -1992 -37
rect -1958 -71 -1924 -37
rect -1508 -71 -1474 -37
rect -1440 -71 -1406 -37
rect -1372 -71 -1338 -37
rect -1304 -71 -1270 -37
rect -1236 -71 -1202 -37
rect -1168 -71 -1134 -37
rect -1100 -71 -1066 -37
rect -650 -71 -616 -37
rect -582 -71 -548 -37
rect -514 -71 -480 -37
rect -446 -71 -412 -37
rect -378 -71 -344 -37
rect -310 -71 -276 -37
rect -242 -71 -208 -37
rect 208 -71 242 -37
rect 276 -71 310 -37
rect 344 -71 378 -37
rect 412 -71 446 -37
rect 480 -71 514 -37
rect 548 -71 582 -37
rect 616 -71 650 -37
rect 1066 -71 1100 -37
rect 1134 -71 1168 -37
rect 1202 -71 1236 -37
rect 1270 -71 1304 -37
rect 1338 -71 1372 -37
rect 1406 -71 1440 -37
rect 1474 -71 1508 -37
rect 1924 -71 1958 -37
rect 1992 -71 2026 -37
rect 2060 -71 2094 -37
rect 2128 -71 2162 -37
rect 2196 -71 2230 -37
rect 2264 -71 2298 -37
rect 2332 -71 2366 -37
rect -2366 -381 -2332 -347
rect -2298 -381 -2264 -347
rect -2230 -381 -2196 -347
rect -2162 -381 -2128 -347
rect -2094 -381 -2060 -347
rect -2026 -381 -1992 -347
rect -1958 -381 -1924 -347
rect -1508 -381 -1474 -347
rect -1440 -381 -1406 -347
rect -1372 -381 -1338 -347
rect -1304 -381 -1270 -347
rect -1236 -381 -1202 -347
rect -1168 -381 -1134 -347
rect -1100 -381 -1066 -347
rect -650 -381 -616 -347
rect -582 -381 -548 -347
rect -514 -381 -480 -347
rect -446 -381 -412 -347
rect -378 -381 -344 -347
rect -310 -381 -276 -347
rect -242 -381 -208 -347
rect 208 -381 242 -347
rect 276 -381 310 -347
rect 344 -381 378 -347
rect 412 -381 446 -347
rect 480 -381 514 -347
rect 548 -381 582 -347
rect 616 -381 650 -347
rect 1066 -381 1100 -347
rect 1134 -381 1168 -347
rect 1202 -381 1236 -347
rect 1270 -381 1304 -347
rect 1338 -381 1372 -347
rect 1406 -381 1440 -347
rect 1474 -381 1508 -347
rect 1924 -381 1958 -347
rect 1992 -381 2026 -347
rect 2060 -381 2094 -347
rect 2128 -381 2162 -347
rect 2196 -381 2230 -347
rect 2264 -381 2298 -347
rect 2332 -381 2366 -347
<< locali >>
rect -2391 347 -2366 381
rect -2332 347 -2306 381
rect -2264 347 -2234 381
rect -2196 347 -2162 381
rect -2128 347 -2094 381
rect -2056 347 -2026 381
rect -1984 347 -1958 381
rect -1924 347 -1899 381
rect -1533 347 -1508 381
rect -1474 347 -1448 381
rect -1406 347 -1376 381
rect -1338 347 -1304 381
rect -1270 347 -1236 381
rect -1198 347 -1168 381
rect -1126 347 -1100 381
rect -1066 347 -1041 381
rect -675 347 -650 381
rect -616 347 -590 381
rect -548 347 -518 381
rect -480 347 -446 381
rect -412 347 -378 381
rect -340 347 -310 381
rect -268 347 -242 381
rect -208 347 -183 381
rect 183 347 208 381
rect 242 347 268 381
rect 310 347 340 381
rect 378 347 412 381
rect 446 347 480 381
rect 518 347 548 381
rect 590 347 616 381
rect 650 347 675 381
rect 1041 347 1066 381
rect 1100 347 1126 381
rect 1168 347 1198 381
rect 1236 347 1270 381
rect 1304 347 1338 381
rect 1376 347 1406 381
rect 1448 347 1474 381
rect 1508 347 1533 381
rect 1899 347 1924 381
rect 1958 347 1984 381
rect 2026 347 2056 381
rect 2094 347 2128 381
rect 2162 347 2196 381
rect 2234 347 2264 381
rect 2306 347 2332 381
rect 2366 347 2391 381
rect -2591 294 -2557 313
rect -2591 226 -2557 228
rect -2591 190 -2557 192
rect -2591 105 -2557 124
rect -1733 294 -1699 313
rect -1733 226 -1699 228
rect -1733 190 -1699 192
rect -1733 105 -1699 124
rect -875 294 -841 313
rect -875 226 -841 228
rect -875 190 -841 192
rect -875 105 -841 124
rect -17 294 17 313
rect -17 226 17 228
rect -17 190 17 192
rect -17 105 17 124
rect 841 294 875 313
rect 841 226 875 228
rect 841 190 875 192
rect 841 105 875 124
rect 1699 294 1733 313
rect 1699 226 1733 228
rect 1699 190 1733 192
rect 1699 105 1733 124
rect 2557 294 2591 313
rect 2557 226 2591 228
rect 2557 190 2591 192
rect 2557 105 2591 124
rect -2391 37 -2366 71
rect -2332 37 -2306 71
rect -2264 37 -2234 71
rect -2196 37 -2162 71
rect -2128 37 -2094 71
rect -2056 37 -2026 71
rect -1984 37 -1958 71
rect -1924 37 -1899 71
rect -1533 37 -1508 71
rect -1474 37 -1448 71
rect -1406 37 -1376 71
rect -1338 37 -1304 71
rect -1270 37 -1236 71
rect -1198 37 -1168 71
rect -1126 37 -1100 71
rect -1066 37 -1041 71
rect -675 37 -650 71
rect -616 37 -590 71
rect -548 37 -518 71
rect -480 37 -446 71
rect -412 37 -378 71
rect -340 37 -310 71
rect -268 37 -242 71
rect -208 37 -183 71
rect 183 37 208 71
rect 242 37 268 71
rect 310 37 340 71
rect 378 37 412 71
rect 446 37 480 71
rect 518 37 548 71
rect 590 37 616 71
rect 650 37 675 71
rect 1041 37 1066 71
rect 1100 37 1126 71
rect 1168 37 1198 71
rect 1236 37 1270 71
rect 1304 37 1338 71
rect 1376 37 1406 71
rect 1448 37 1474 71
rect 1508 37 1533 71
rect 1899 37 1924 71
rect 1958 37 1984 71
rect 2026 37 2056 71
rect 2094 37 2128 71
rect 2162 37 2196 71
rect 2234 37 2264 71
rect 2306 37 2332 71
rect 2366 37 2391 71
rect -2391 -71 -2366 -37
rect -2332 -71 -2306 -37
rect -2264 -71 -2234 -37
rect -2196 -71 -2162 -37
rect -2128 -71 -2094 -37
rect -2056 -71 -2026 -37
rect -1984 -71 -1958 -37
rect -1924 -71 -1899 -37
rect -1533 -71 -1508 -37
rect -1474 -71 -1448 -37
rect -1406 -71 -1376 -37
rect -1338 -71 -1304 -37
rect -1270 -71 -1236 -37
rect -1198 -71 -1168 -37
rect -1126 -71 -1100 -37
rect -1066 -71 -1041 -37
rect -675 -71 -650 -37
rect -616 -71 -590 -37
rect -548 -71 -518 -37
rect -480 -71 -446 -37
rect -412 -71 -378 -37
rect -340 -71 -310 -37
rect -268 -71 -242 -37
rect -208 -71 -183 -37
rect 183 -71 208 -37
rect 242 -71 268 -37
rect 310 -71 340 -37
rect 378 -71 412 -37
rect 446 -71 480 -37
rect 518 -71 548 -37
rect 590 -71 616 -37
rect 650 -71 675 -37
rect 1041 -71 1066 -37
rect 1100 -71 1126 -37
rect 1168 -71 1198 -37
rect 1236 -71 1270 -37
rect 1304 -71 1338 -37
rect 1376 -71 1406 -37
rect 1448 -71 1474 -37
rect 1508 -71 1533 -37
rect 1899 -71 1924 -37
rect 1958 -71 1984 -37
rect 2026 -71 2056 -37
rect 2094 -71 2128 -37
rect 2162 -71 2196 -37
rect 2234 -71 2264 -37
rect 2306 -71 2332 -37
rect 2366 -71 2391 -37
rect -2591 -124 -2557 -105
rect -2591 -192 -2557 -190
rect -2591 -228 -2557 -226
rect -2591 -313 -2557 -294
rect -1733 -124 -1699 -105
rect -1733 -192 -1699 -190
rect -1733 -228 -1699 -226
rect -1733 -313 -1699 -294
rect -875 -124 -841 -105
rect -875 -192 -841 -190
rect -875 -228 -841 -226
rect -875 -313 -841 -294
rect -17 -124 17 -105
rect -17 -192 17 -190
rect -17 -228 17 -226
rect -17 -313 17 -294
rect 841 -124 875 -105
rect 841 -192 875 -190
rect 841 -228 875 -226
rect 841 -313 875 -294
rect 1699 -124 1733 -105
rect 1699 -192 1733 -190
rect 1699 -228 1733 -226
rect 1699 -313 1733 -294
rect 2557 -124 2591 -105
rect 2557 -192 2591 -190
rect 2557 -228 2591 -226
rect 2557 -313 2591 -294
rect -2391 -381 -2366 -347
rect -2332 -381 -2306 -347
rect -2264 -381 -2234 -347
rect -2196 -381 -2162 -347
rect -2128 -381 -2094 -347
rect -2056 -381 -2026 -347
rect -1984 -381 -1958 -347
rect -1924 -381 -1899 -347
rect -1533 -381 -1508 -347
rect -1474 -381 -1448 -347
rect -1406 -381 -1376 -347
rect -1338 -381 -1304 -347
rect -1270 -381 -1236 -347
rect -1198 -381 -1168 -347
rect -1126 -381 -1100 -347
rect -1066 -381 -1041 -347
rect -675 -381 -650 -347
rect -616 -381 -590 -347
rect -548 -381 -518 -347
rect -480 -381 -446 -347
rect -412 -381 -378 -347
rect -340 -381 -310 -347
rect -268 -381 -242 -347
rect -208 -381 -183 -347
rect 183 -381 208 -347
rect 242 -381 268 -347
rect 310 -381 340 -347
rect 378 -381 412 -347
rect 446 -381 480 -347
rect 518 -381 548 -347
rect 590 -381 616 -347
rect 650 -381 675 -347
rect 1041 -381 1066 -347
rect 1100 -381 1126 -347
rect 1168 -381 1198 -347
rect 1236 -381 1270 -347
rect 1304 -381 1338 -347
rect 1376 -381 1406 -347
rect 1448 -381 1474 -347
rect 1508 -381 1533 -347
rect 1899 -381 1924 -347
rect 1958 -381 1984 -347
rect 2026 -381 2056 -347
rect 2094 -381 2128 -347
rect 2162 -381 2196 -347
rect 2234 -381 2264 -347
rect 2306 -381 2332 -347
rect 2366 -381 2391 -347
<< viali >>
rect -2306 347 -2298 381
rect -2298 347 -2272 381
rect -2234 347 -2230 381
rect -2230 347 -2200 381
rect -2162 347 -2128 381
rect -2090 347 -2060 381
rect -2060 347 -2056 381
rect -2018 347 -1992 381
rect -1992 347 -1984 381
rect -1448 347 -1440 381
rect -1440 347 -1414 381
rect -1376 347 -1372 381
rect -1372 347 -1342 381
rect -1304 347 -1270 381
rect -1232 347 -1202 381
rect -1202 347 -1198 381
rect -1160 347 -1134 381
rect -1134 347 -1126 381
rect -590 347 -582 381
rect -582 347 -556 381
rect -518 347 -514 381
rect -514 347 -484 381
rect -446 347 -412 381
rect -374 347 -344 381
rect -344 347 -340 381
rect -302 347 -276 381
rect -276 347 -268 381
rect 268 347 276 381
rect 276 347 302 381
rect 340 347 344 381
rect 344 347 374 381
rect 412 347 446 381
rect 484 347 514 381
rect 514 347 518 381
rect 556 347 582 381
rect 582 347 590 381
rect 1126 347 1134 381
rect 1134 347 1160 381
rect 1198 347 1202 381
rect 1202 347 1232 381
rect 1270 347 1304 381
rect 1342 347 1372 381
rect 1372 347 1376 381
rect 1414 347 1440 381
rect 1440 347 1448 381
rect 1984 347 1992 381
rect 1992 347 2018 381
rect 2056 347 2060 381
rect 2060 347 2090 381
rect 2128 347 2162 381
rect 2200 347 2230 381
rect 2230 347 2234 381
rect 2272 347 2298 381
rect 2298 347 2306 381
rect -2591 260 -2557 262
rect -2591 228 -2557 260
rect -2591 158 -2557 190
rect -2591 156 -2557 158
rect -1733 260 -1699 262
rect -1733 228 -1699 260
rect -1733 158 -1699 190
rect -1733 156 -1699 158
rect -875 260 -841 262
rect -875 228 -841 260
rect -875 158 -841 190
rect -875 156 -841 158
rect -17 260 17 262
rect -17 228 17 260
rect -17 158 17 190
rect -17 156 17 158
rect 841 260 875 262
rect 841 228 875 260
rect 841 158 875 190
rect 841 156 875 158
rect 1699 260 1733 262
rect 1699 228 1733 260
rect 1699 158 1733 190
rect 1699 156 1733 158
rect 2557 260 2591 262
rect 2557 228 2591 260
rect 2557 158 2591 190
rect 2557 156 2591 158
rect -2306 37 -2298 71
rect -2298 37 -2272 71
rect -2234 37 -2230 71
rect -2230 37 -2200 71
rect -2162 37 -2128 71
rect -2090 37 -2060 71
rect -2060 37 -2056 71
rect -2018 37 -1992 71
rect -1992 37 -1984 71
rect -1448 37 -1440 71
rect -1440 37 -1414 71
rect -1376 37 -1372 71
rect -1372 37 -1342 71
rect -1304 37 -1270 71
rect -1232 37 -1202 71
rect -1202 37 -1198 71
rect -1160 37 -1134 71
rect -1134 37 -1126 71
rect -590 37 -582 71
rect -582 37 -556 71
rect -518 37 -514 71
rect -514 37 -484 71
rect -446 37 -412 71
rect -374 37 -344 71
rect -344 37 -340 71
rect -302 37 -276 71
rect -276 37 -268 71
rect 268 37 276 71
rect 276 37 302 71
rect 340 37 344 71
rect 344 37 374 71
rect 412 37 446 71
rect 484 37 514 71
rect 514 37 518 71
rect 556 37 582 71
rect 582 37 590 71
rect 1126 37 1134 71
rect 1134 37 1160 71
rect 1198 37 1202 71
rect 1202 37 1232 71
rect 1270 37 1304 71
rect 1342 37 1372 71
rect 1372 37 1376 71
rect 1414 37 1440 71
rect 1440 37 1448 71
rect 1984 37 1992 71
rect 1992 37 2018 71
rect 2056 37 2060 71
rect 2060 37 2090 71
rect 2128 37 2162 71
rect 2200 37 2230 71
rect 2230 37 2234 71
rect 2272 37 2298 71
rect 2298 37 2306 71
rect -2306 -71 -2298 -37
rect -2298 -71 -2272 -37
rect -2234 -71 -2230 -37
rect -2230 -71 -2200 -37
rect -2162 -71 -2128 -37
rect -2090 -71 -2060 -37
rect -2060 -71 -2056 -37
rect -2018 -71 -1992 -37
rect -1992 -71 -1984 -37
rect -1448 -71 -1440 -37
rect -1440 -71 -1414 -37
rect -1376 -71 -1372 -37
rect -1372 -71 -1342 -37
rect -1304 -71 -1270 -37
rect -1232 -71 -1202 -37
rect -1202 -71 -1198 -37
rect -1160 -71 -1134 -37
rect -1134 -71 -1126 -37
rect -590 -71 -582 -37
rect -582 -71 -556 -37
rect -518 -71 -514 -37
rect -514 -71 -484 -37
rect -446 -71 -412 -37
rect -374 -71 -344 -37
rect -344 -71 -340 -37
rect -302 -71 -276 -37
rect -276 -71 -268 -37
rect 268 -71 276 -37
rect 276 -71 302 -37
rect 340 -71 344 -37
rect 344 -71 374 -37
rect 412 -71 446 -37
rect 484 -71 514 -37
rect 514 -71 518 -37
rect 556 -71 582 -37
rect 582 -71 590 -37
rect 1126 -71 1134 -37
rect 1134 -71 1160 -37
rect 1198 -71 1202 -37
rect 1202 -71 1232 -37
rect 1270 -71 1304 -37
rect 1342 -71 1372 -37
rect 1372 -71 1376 -37
rect 1414 -71 1440 -37
rect 1440 -71 1448 -37
rect 1984 -71 1992 -37
rect 1992 -71 2018 -37
rect 2056 -71 2060 -37
rect 2060 -71 2090 -37
rect 2128 -71 2162 -37
rect 2200 -71 2230 -37
rect 2230 -71 2234 -37
rect 2272 -71 2298 -37
rect 2298 -71 2306 -37
rect -2591 -158 -2557 -156
rect -2591 -190 -2557 -158
rect -2591 -260 -2557 -228
rect -2591 -262 -2557 -260
rect -1733 -158 -1699 -156
rect -1733 -190 -1699 -158
rect -1733 -260 -1699 -228
rect -1733 -262 -1699 -260
rect -875 -158 -841 -156
rect -875 -190 -841 -158
rect -875 -260 -841 -228
rect -875 -262 -841 -260
rect -17 -158 17 -156
rect -17 -190 17 -158
rect -17 -260 17 -228
rect -17 -262 17 -260
rect 841 -158 875 -156
rect 841 -190 875 -158
rect 841 -260 875 -228
rect 841 -262 875 -260
rect 1699 -158 1733 -156
rect 1699 -190 1733 -158
rect 1699 -260 1733 -228
rect 1699 -262 1733 -260
rect 2557 -158 2591 -156
rect 2557 -190 2591 -158
rect 2557 -260 2591 -228
rect 2557 -262 2591 -260
rect -2306 -381 -2298 -347
rect -2298 -381 -2272 -347
rect -2234 -381 -2230 -347
rect -2230 -381 -2200 -347
rect -2162 -381 -2128 -347
rect -2090 -381 -2060 -347
rect -2060 -381 -2056 -347
rect -2018 -381 -1992 -347
rect -1992 -381 -1984 -347
rect -1448 -381 -1440 -347
rect -1440 -381 -1414 -347
rect -1376 -381 -1372 -347
rect -1372 -381 -1342 -347
rect -1304 -381 -1270 -347
rect -1232 -381 -1202 -347
rect -1202 -381 -1198 -347
rect -1160 -381 -1134 -347
rect -1134 -381 -1126 -347
rect -590 -381 -582 -347
rect -582 -381 -556 -347
rect -518 -381 -514 -347
rect -514 -381 -484 -347
rect -446 -381 -412 -347
rect -374 -381 -344 -347
rect -344 -381 -340 -347
rect -302 -381 -276 -347
rect -276 -381 -268 -347
rect 268 -381 276 -347
rect 276 -381 302 -347
rect 340 -381 344 -347
rect 344 -381 374 -347
rect 412 -381 446 -347
rect 484 -381 514 -347
rect 514 -381 518 -347
rect 556 -381 582 -347
rect 582 -381 590 -347
rect 1126 -381 1134 -347
rect 1134 -381 1160 -347
rect 1198 -381 1202 -347
rect 1202 -381 1232 -347
rect 1270 -381 1304 -347
rect 1342 -381 1372 -347
rect 1372 -381 1376 -347
rect 1414 -381 1440 -347
rect 1440 -381 1448 -347
rect 1984 -381 1992 -347
rect 1992 -381 2018 -347
rect 2056 -381 2060 -347
rect 2060 -381 2090 -347
rect 2128 -381 2162 -347
rect 2200 -381 2230 -347
rect 2230 -381 2234 -347
rect 2272 -381 2298 -347
rect 2298 -381 2306 -347
<< metal1 >>
rect -2349 381 -1941 387
rect -2349 347 -2306 381
rect -2272 347 -2234 381
rect -2200 347 -2162 381
rect -2128 347 -2090 381
rect -2056 347 -2018 381
rect -1984 347 -1941 381
rect -2349 341 -1941 347
rect -1491 381 -1083 387
rect -1491 347 -1448 381
rect -1414 347 -1376 381
rect -1342 347 -1304 381
rect -1270 347 -1232 381
rect -1198 347 -1160 381
rect -1126 347 -1083 381
rect -1491 341 -1083 347
rect -633 381 -225 387
rect -633 347 -590 381
rect -556 347 -518 381
rect -484 347 -446 381
rect -412 347 -374 381
rect -340 347 -302 381
rect -268 347 -225 381
rect -633 341 -225 347
rect 225 381 633 387
rect 225 347 268 381
rect 302 347 340 381
rect 374 347 412 381
rect 446 347 484 381
rect 518 347 556 381
rect 590 347 633 381
rect 225 341 633 347
rect 1083 381 1491 387
rect 1083 347 1126 381
rect 1160 347 1198 381
rect 1232 347 1270 381
rect 1304 347 1342 381
rect 1376 347 1414 381
rect 1448 347 1491 381
rect 1083 341 1491 347
rect 1941 381 2349 387
rect 1941 347 1984 381
rect 2018 347 2056 381
rect 2090 347 2128 381
rect 2162 347 2200 381
rect 2234 347 2272 381
rect 2306 347 2349 381
rect 1941 341 2349 347
rect -2597 262 -2551 309
rect -2597 228 -2591 262
rect -2557 228 -2551 262
rect -2597 190 -2551 228
rect -2597 156 -2591 190
rect -2557 156 -2551 190
rect -2597 109 -2551 156
rect -1739 262 -1693 309
rect -1739 228 -1733 262
rect -1699 228 -1693 262
rect -1739 190 -1693 228
rect -1739 156 -1733 190
rect -1699 156 -1693 190
rect -1739 109 -1693 156
rect -881 262 -835 309
rect -881 228 -875 262
rect -841 228 -835 262
rect -881 190 -835 228
rect -881 156 -875 190
rect -841 156 -835 190
rect -881 109 -835 156
rect -23 262 23 309
rect -23 228 -17 262
rect 17 228 23 262
rect -23 190 23 228
rect -23 156 -17 190
rect 17 156 23 190
rect -23 109 23 156
rect 835 262 881 309
rect 835 228 841 262
rect 875 228 881 262
rect 835 190 881 228
rect 835 156 841 190
rect 875 156 881 190
rect 835 109 881 156
rect 1693 262 1739 309
rect 1693 228 1699 262
rect 1733 228 1739 262
rect 1693 190 1739 228
rect 1693 156 1699 190
rect 1733 156 1739 190
rect 1693 109 1739 156
rect 2551 262 2597 309
rect 2551 228 2557 262
rect 2591 228 2597 262
rect 2551 190 2597 228
rect 2551 156 2557 190
rect 2591 156 2597 190
rect 2551 109 2597 156
rect -2349 71 -1941 77
rect -2349 37 -2306 71
rect -2272 37 -2234 71
rect -2200 37 -2162 71
rect -2128 37 -2090 71
rect -2056 37 -2018 71
rect -1984 37 -1941 71
rect -2349 31 -1941 37
rect -1491 71 -1083 77
rect -1491 37 -1448 71
rect -1414 37 -1376 71
rect -1342 37 -1304 71
rect -1270 37 -1232 71
rect -1198 37 -1160 71
rect -1126 37 -1083 71
rect -1491 31 -1083 37
rect -633 71 -225 77
rect -633 37 -590 71
rect -556 37 -518 71
rect -484 37 -446 71
rect -412 37 -374 71
rect -340 37 -302 71
rect -268 37 -225 71
rect -633 31 -225 37
rect 225 71 633 77
rect 225 37 268 71
rect 302 37 340 71
rect 374 37 412 71
rect 446 37 484 71
rect 518 37 556 71
rect 590 37 633 71
rect 225 31 633 37
rect 1083 71 1491 77
rect 1083 37 1126 71
rect 1160 37 1198 71
rect 1232 37 1270 71
rect 1304 37 1342 71
rect 1376 37 1414 71
rect 1448 37 1491 71
rect 1083 31 1491 37
rect 1941 71 2349 77
rect 1941 37 1984 71
rect 2018 37 2056 71
rect 2090 37 2128 71
rect 2162 37 2200 71
rect 2234 37 2272 71
rect 2306 37 2349 71
rect 1941 31 2349 37
rect -2349 -37 -1941 -31
rect -2349 -71 -2306 -37
rect -2272 -71 -2234 -37
rect -2200 -71 -2162 -37
rect -2128 -71 -2090 -37
rect -2056 -71 -2018 -37
rect -1984 -71 -1941 -37
rect -2349 -77 -1941 -71
rect -1491 -37 -1083 -31
rect -1491 -71 -1448 -37
rect -1414 -71 -1376 -37
rect -1342 -71 -1304 -37
rect -1270 -71 -1232 -37
rect -1198 -71 -1160 -37
rect -1126 -71 -1083 -37
rect -1491 -77 -1083 -71
rect -633 -37 -225 -31
rect -633 -71 -590 -37
rect -556 -71 -518 -37
rect -484 -71 -446 -37
rect -412 -71 -374 -37
rect -340 -71 -302 -37
rect -268 -71 -225 -37
rect -633 -77 -225 -71
rect 225 -37 633 -31
rect 225 -71 268 -37
rect 302 -71 340 -37
rect 374 -71 412 -37
rect 446 -71 484 -37
rect 518 -71 556 -37
rect 590 -71 633 -37
rect 225 -77 633 -71
rect 1083 -37 1491 -31
rect 1083 -71 1126 -37
rect 1160 -71 1198 -37
rect 1232 -71 1270 -37
rect 1304 -71 1342 -37
rect 1376 -71 1414 -37
rect 1448 -71 1491 -37
rect 1083 -77 1491 -71
rect 1941 -37 2349 -31
rect 1941 -71 1984 -37
rect 2018 -71 2056 -37
rect 2090 -71 2128 -37
rect 2162 -71 2200 -37
rect 2234 -71 2272 -37
rect 2306 -71 2349 -37
rect 1941 -77 2349 -71
rect -2597 -156 -2551 -109
rect -2597 -190 -2591 -156
rect -2557 -190 -2551 -156
rect -2597 -228 -2551 -190
rect -2597 -262 -2591 -228
rect -2557 -262 -2551 -228
rect -2597 -309 -2551 -262
rect -1739 -156 -1693 -109
rect -1739 -190 -1733 -156
rect -1699 -190 -1693 -156
rect -1739 -228 -1693 -190
rect -1739 -262 -1733 -228
rect -1699 -262 -1693 -228
rect -1739 -309 -1693 -262
rect -881 -156 -835 -109
rect -881 -190 -875 -156
rect -841 -190 -835 -156
rect -881 -228 -835 -190
rect -881 -262 -875 -228
rect -841 -262 -835 -228
rect -881 -309 -835 -262
rect -23 -156 23 -109
rect -23 -190 -17 -156
rect 17 -190 23 -156
rect -23 -228 23 -190
rect -23 -262 -17 -228
rect 17 -262 23 -228
rect -23 -309 23 -262
rect 835 -156 881 -109
rect 835 -190 841 -156
rect 875 -190 881 -156
rect 835 -228 881 -190
rect 835 -262 841 -228
rect 875 -262 881 -228
rect 835 -309 881 -262
rect 1693 -156 1739 -109
rect 1693 -190 1699 -156
rect 1733 -190 1739 -156
rect 1693 -228 1739 -190
rect 1693 -262 1699 -228
rect 1733 -262 1739 -228
rect 1693 -309 1739 -262
rect 2551 -156 2597 -109
rect 2551 -190 2557 -156
rect 2591 -190 2597 -156
rect 2551 -228 2597 -190
rect 2551 -262 2557 -228
rect 2591 -262 2597 -228
rect 2551 -309 2597 -262
rect -2349 -347 -1941 -341
rect -2349 -381 -2306 -347
rect -2272 -381 -2234 -347
rect -2200 -381 -2162 -347
rect -2128 -381 -2090 -347
rect -2056 -381 -2018 -347
rect -1984 -381 -1941 -347
rect -2349 -387 -1941 -381
rect -1491 -347 -1083 -341
rect -1491 -381 -1448 -347
rect -1414 -381 -1376 -347
rect -1342 -381 -1304 -347
rect -1270 -381 -1232 -347
rect -1198 -381 -1160 -347
rect -1126 -381 -1083 -347
rect -1491 -387 -1083 -381
rect -633 -347 -225 -341
rect -633 -381 -590 -347
rect -556 -381 -518 -347
rect -484 -381 -446 -347
rect -412 -381 -374 -347
rect -340 -381 -302 -347
rect -268 -381 -225 -347
rect -633 -387 -225 -381
rect 225 -347 633 -341
rect 225 -381 268 -347
rect 302 -381 340 -347
rect 374 -381 412 -347
rect 446 -381 484 -347
rect 518 -381 556 -347
rect 590 -381 633 -347
rect 225 -387 633 -381
rect 1083 -347 1491 -341
rect 1083 -381 1126 -347
rect 1160 -381 1198 -347
rect 1232 -381 1270 -347
rect 1304 -381 1342 -347
rect 1376 -381 1414 -347
rect 1448 -381 1491 -347
rect 1083 -387 1491 -381
rect 1941 -347 2349 -341
rect 1941 -381 1984 -347
rect 2018 -381 2056 -347
rect 2090 -381 2128 -347
rect 2162 -381 2200 -347
rect 2234 -381 2272 -347
rect 2306 -381 2349 -347
rect 1941 -387 2349 -381
<< end >>
