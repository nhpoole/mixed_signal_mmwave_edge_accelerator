magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< error_p >>
rect -1645 566 1645 600
rect -1675 -566 1675 566
rect -1645 -600 1645 -566
<< nwell >>
rect -1645 -600 1645 600
<< mvpmos >>
rect -1551 -500 -1451 500
rect -1393 -500 -1293 500
rect -1235 -500 -1135 500
rect -1077 -500 -977 500
rect -919 -500 -819 500
rect -761 -500 -661 500
rect -603 -500 -503 500
rect -445 -500 -345 500
rect -287 -500 -187 500
rect -129 -500 -29 500
rect 29 -500 129 500
rect 187 -500 287 500
rect 345 -500 445 500
rect 503 -500 603 500
rect 661 -500 761 500
rect 819 -500 919 500
rect 977 -500 1077 500
rect 1135 -500 1235 500
rect 1293 -500 1393 500
rect 1451 -500 1551 500
<< mvpdiff >>
rect -1609 488 -1551 500
rect -1609 -488 -1597 488
rect -1563 -488 -1551 488
rect -1609 -500 -1551 -488
rect -1451 488 -1393 500
rect -1451 -488 -1439 488
rect -1405 -488 -1393 488
rect -1451 -500 -1393 -488
rect -1293 488 -1235 500
rect -1293 -488 -1281 488
rect -1247 -488 -1235 488
rect -1293 -500 -1235 -488
rect -1135 488 -1077 500
rect -1135 -488 -1123 488
rect -1089 -488 -1077 488
rect -1135 -500 -1077 -488
rect -977 488 -919 500
rect -977 -488 -965 488
rect -931 -488 -919 488
rect -977 -500 -919 -488
rect -819 488 -761 500
rect -819 -488 -807 488
rect -773 -488 -761 488
rect -819 -500 -761 -488
rect -661 488 -603 500
rect -661 -488 -649 488
rect -615 -488 -603 488
rect -661 -500 -603 -488
rect -503 488 -445 500
rect -503 -488 -491 488
rect -457 -488 -445 488
rect -503 -500 -445 -488
rect -345 488 -287 500
rect -345 -488 -333 488
rect -299 -488 -287 488
rect -345 -500 -287 -488
rect -187 488 -129 500
rect -187 -488 -175 488
rect -141 -488 -129 488
rect -187 -500 -129 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 129 488 187 500
rect 129 -488 141 488
rect 175 -488 187 488
rect 129 -500 187 -488
rect 287 488 345 500
rect 287 -488 299 488
rect 333 -488 345 488
rect 287 -500 345 -488
rect 445 488 503 500
rect 445 -488 457 488
rect 491 -488 503 488
rect 445 -500 503 -488
rect 603 488 661 500
rect 603 -488 615 488
rect 649 -488 661 488
rect 603 -500 661 -488
rect 761 488 819 500
rect 761 -488 773 488
rect 807 -488 819 488
rect 761 -500 819 -488
rect 919 488 977 500
rect 919 -488 931 488
rect 965 -488 977 488
rect 919 -500 977 -488
rect 1077 488 1135 500
rect 1077 -488 1089 488
rect 1123 -488 1135 488
rect 1077 -500 1135 -488
rect 1235 488 1293 500
rect 1235 -488 1247 488
rect 1281 -488 1293 488
rect 1235 -500 1293 -488
rect 1393 488 1451 500
rect 1393 -488 1405 488
rect 1439 -488 1451 488
rect 1393 -500 1451 -488
rect 1551 488 1609 500
rect 1551 -488 1563 488
rect 1597 -488 1609 488
rect 1551 -500 1609 -488
<< mvpdiffc >>
rect -1597 -488 -1563 488
rect -1439 -488 -1405 488
rect -1281 -488 -1247 488
rect -1123 -488 -1089 488
rect -965 -488 -931 488
rect -807 -488 -773 488
rect -649 -488 -615 488
rect -491 -488 -457 488
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
rect 457 -488 491 488
rect 615 -488 649 488
rect 773 -488 807 488
rect 931 -488 965 488
rect 1089 -488 1123 488
rect 1247 -488 1281 488
rect 1405 -488 1439 488
rect 1563 -488 1597 488
<< poly >>
rect -1537 581 -1465 597
rect -1537 564 -1521 581
rect -1551 547 -1521 564
rect -1481 564 -1465 581
rect -1379 581 -1307 597
rect -1379 564 -1363 581
rect -1481 547 -1451 564
rect -1551 500 -1451 547
rect -1393 547 -1363 564
rect -1323 564 -1307 581
rect -1221 581 -1149 597
rect -1221 564 -1205 581
rect -1323 547 -1293 564
rect -1393 500 -1293 547
rect -1235 547 -1205 564
rect -1165 564 -1149 581
rect -1063 581 -991 597
rect -1063 564 -1047 581
rect -1165 547 -1135 564
rect -1235 500 -1135 547
rect -1077 547 -1047 564
rect -1007 564 -991 581
rect -905 581 -833 597
rect -905 564 -889 581
rect -1007 547 -977 564
rect -1077 500 -977 547
rect -919 547 -889 564
rect -849 564 -833 581
rect -747 581 -675 597
rect -747 564 -731 581
rect -849 547 -819 564
rect -919 500 -819 547
rect -761 547 -731 564
rect -691 564 -675 581
rect -589 581 -517 597
rect -589 564 -573 581
rect -691 547 -661 564
rect -761 500 -661 547
rect -603 547 -573 564
rect -533 564 -517 581
rect -431 581 -359 597
rect -431 564 -415 581
rect -533 547 -503 564
rect -603 500 -503 547
rect -445 547 -415 564
rect -375 564 -359 581
rect -273 581 -201 597
rect -273 564 -257 581
rect -375 547 -345 564
rect -445 500 -345 547
rect -287 547 -257 564
rect -217 564 -201 581
rect -115 581 -43 597
rect -115 564 -99 581
rect -217 547 -187 564
rect -287 500 -187 547
rect -129 547 -99 564
rect -59 564 -43 581
rect 43 581 115 597
rect 43 564 59 581
rect -59 547 -29 564
rect -129 500 -29 547
rect 29 547 59 564
rect 99 564 115 581
rect 201 581 273 597
rect 201 564 217 581
rect 99 547 129 564
rect 29 500 129 547
rect 187 547 217 564
rect 257 564 273 581
rect 359 581 431 597
rect 359 564 375 581
rect 257 547 287 564
rect 187 500 287 547
rect 345 547 375 564
rect 415 564 431 581
rect 517 581 589 597
rect 517 564 533 581
rect 415 547 445 564
rect 345 500 445 547
rect 503 547 533 564
rect 573 564 589 581
rect 675 581 747 597
rect 675 564 691 581
rect 573 547 603 564
rect 503 500 603 547
rect 661 547 691 564
rect 731 564 747 581
rect 833 581 905 597
rect 833 564 849 581
rect 731 547 761 564
rect 661 500 761 547
rect 819 547 849 564
rect 889 564 905 581
rect 991 581 1063 597
rect 991 564 1007 581
rect 889 547 919 564
rect 819 500 919 547
rect 977 547 1007 564
rect 1047 564 1063 581
rect 1149 581 1221 597
rect 1149 564 1165 581
rect 1047 547 1077 564
rect 977 500 1077 547
rect 1135 547 1165 564
rect 1205 564 1221 581
rect 1307 581 1379 597
rect 1307 564 1323 581
rect 1205 547 1235 564
rect 1135 500 1235 547
rect 1293 547 1323 564
rect 1363 564 1379 581
rect 1465 581 1537 597
rect 1465 564 1481 581
rect 1363 547 1393 564
rect 1293 500 1393 547
rect 1451 547 1481 564
rect 1521 564 1537 581
rect 1521 547 1551 564
rect 1451 500 1551 547
rect -1551 -547 -1451 -500
rect -1551 -564 -1521 -547
rect -1537 -581 -1521 -564
rect -1481 -564 -1451 -547
rect -1393 -547 -1293 -500
rect -1393 -564 -1363 -547
rect -1481 -581 -1465 -564
rect -1537 -597 -1465 -581
rect -1379 -581 -1363 -564
rect -1323 -564 -1293 -547
rect -1235 -547 -1135 -500
rect -1235 -564 -1205 -547
rect -1323 -581 -1307 -564
rect -1379 -597 -1307 -581
rect -1221 -581 -1205 -564
rect -1165 -564 -1135 -547
rect -1077 -547 -977 -500
rect -1077 -564 -1047 -547
rect -1165 -581 -1149 -564
rect -1221 -597 -1149 -581
rect -1063 -581 -1047 -564
rect -1007 -564 -977 -547
rect -919 -547 -819 -500
rect -919 -564 -889 -547
rect -1007 -581 -991 -564
rect -1063 -597 -991 -581
rect -905 -581 -889 -564
rect -849 -564 -819 -547
rect -761 -547 -661 -500
rect -761 -564 -731 -547
rect -849 -581 -833 -564
rect -905 -597 -833 -581
rect -747 -581 -731 -564
rect -691 -564 -661 -547
rect -603 -547 -503 -500
rect -603 -564 -573 -547
rect -691 -581 -675 -564
rect -747 -597 -675 -581
rect -589 -581 -573 -564
rect -533 -564 -503 -547
rect -445 -547 -345 -500
rect -445 -564 -415 -547
rect -533 -581 -517 -564
rect -589 -597 -517 -581
rect -431 -581 -415 -564
rect -375 -564 -345 -547
rect -287 -547 -187 -500
rect -287 -564 -257 -547
rect -375 -581 -359 -564
rect -431 -597 -359 -581
rect -273 -581 -257 -564
rect -217 -564 -187 -547
rect -129 -547 -29 -500
rect -129 -564 -99 -547
rect -217 -581 -201 -564
rect -273 -597 -201 -581
rect -115 -581 -99 -564
rect -59 -564 -29 -547
rect 29 -547 129 -500
rect 29 -564 59 -547
rect -59 -581 -43 -564
rect -115 -597 -43 -581
rect 43 -581 59 -564
rect 99 -564 129 -547
rect 187 -547 287 -500
rect 187 -564 217 -547
rect 99 -581 115 -564
rect 43 -597 115 -581
rect 201 -581 217 -564
rect 257 -564 287 -547
rect 345 -547 445 -500
rect 345 -564 375 -547
rect 257 -581 273 -564
rect 201 -597 273 -581
rect 359 -581 375 -564
rect 415 -564 445 -547
rect 503 -547 603 -500
rect 503 -564 533 -547
rect 415 -581 431 -564
rect 359 -597 431 -581
rect 517 -581 533 -564
rect 573 -564 603 -547
rect 661 -547 761 -500
rect 661 -564 691 -547
rect 573 -581 589 -564
rect 517 -597 589 -581
rect 675 -581 691 -564
rect 731 -564 761 -547
rect 819 -547 919 -500
rect 819 -564 849 -547
rect 731 -581 747 -564
rect 675 -597 747 -581
rect 833 -581 849 -564
rect 889 -564 919 -547
rect 977 -547 1077 -500
rect 977 -564 1007 -547
rect 889 -581 905 -564
rect 833 -597 905 -581
rect 991 -581 1007 -564
rect 1047 -564 1077 -547
rect 1135 -547 1235 -500
rect 1135 -564 1165 -547
rect 1047 -581 1063 -564
rect 991 -597 1063 -581
rect 1149 -581 1165 -564
rect 1205 -564 1235 -547
rect 1293 -547 1393 -500
rect 1293 -564 1323 -547
rect 1205 -581 1221 -564
rect 1149 -597 1221 -581
rect 1307 -581 1323 -564
rect 1363 -564 1393 -547
rect 1451 -547 1551 -500
rect 1451 -564 1481 -547
rect 1363 -581 1379 -564
rect 1307 -597 1379 -581
rect 1465 -581 1481 -564
rect 1521 -564 1551 -547
rect 1521 -581 1537 -564
rect 1465 -597 1537 -581
<< polycont >>
rect -1521 547 -1481 581
rect -1363 547 -1323 581
rect -1205 547 -1165 581
rect -1047 547 -1007 581
rect -889 547 -849 581
rect -731 547 -691 581
rect -573 547 -533 581
rect -415 547 -375 581
rect -257 547 -217 581
rect -99 547 -59 581
rect 59 547 99 581
rect 217 547 257 581
rect 375 547 415 581
rect 533 547 573 581
rect 691 547 731 581
rect 849 547 889 581
rect 1007 547 1047 581
rect 1165 547 1205 581
rect 1323 547 1363 581
rect 1481 547 1521 581
rect -1521 -581 -1481 -547
rect -1363 -581 -1323 -547
rect -1205 -581 -1165 -547
rect -1047 -581 -1007 -547
rect -889 -581 -849 -547
rect -731 -581 -691 -547
rect -573 -581 -533 -547
rect -415 -581 -375 -547
rect -257 -581 -217 -547
rect -99 -581 -59 -547
rect 59 -581 99 -547
rect 217 -581 257 -547
rect 375 -581 415 -547
rect 533 -581 573 -547
rect 691 -581 731 -547
rect 849 -581 889 -547
rect 1007 -581 1047 -547
rect 1165 -581 1205 -547
rect 1323 -581 1363 -547
rect 1481 -581 1521 -547
<< locali >>
rect -1537 547 -1521 581
rect -1481 547 -1465 581
rect -1379 547 -1363 581
rect -1323 547 -1307 581
rect -1221 547 -1205 581
rect -1165 547 -1149 581
rect -1063 547 -1047 581
rect -1007 547 -991 581
rect -905 547 -889 581
rect -849 547 -833 581
rect -747 547 -731 581
rect -691 547 -675 581
rect -589 547 -573 581
rect -533 547 -517 581
rect -431 547 -415 581
rect -375 547 -359 581
rect -273 547 -257 581
rect -217 547 -201 581
rect -115 547 -99 581
rect -59 547 -43 581
rect 43 547 59 581
rect 99 547 115 581
rect 201 547 217 581
rect 257 547 273 581
rect 359 547 375 581
rect 415 547 431 581
rect 517 547 533 581
rect 573 547 589 581
rect 675 547 691 581
rect 731 547 747 581
rect 833 547 849 581
rect 889 547 905 581
rect 991 547 1007 581
rect 1047 547 1063 581
rect 1149 547 1165 581
rect 1205 547 1221 581
rect 1307 547 1323 581
rect 1363 547 1379 581
rect 1465 547 1481 581
rect 1521 547 1537 581
rect -1597 488 -1563 504
rect -1597 -504 -1563 -488
rect -1439 488 -1405 504
rect -1439 -504 -1405 -488
rect -1281 488 -1247 504
rect -1281 -504 -1247 -488
rect -1123 488 -1089 504
rect -1123 -504 -1089 -488
rect -965 488 -931 504
rect -965 -504 -931 -488
rect -807 488 -773 504
rect -807 -504 -773 -488
rect -649 488 -615 504
rect -649 -504 -615 -488
rect -491 488 -457 504
rect -491 -504 -457 -488
rect -333 488 -299 504
rect -333 -504 -299 -488
rect -175 488 -141 504
rect -175 -504 -141 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 141 488 175 504
rect 141 -504 175 -488
rect 299 488 333 504
rect 299 -504 333 -488
rect 457 488 491 504
rect 457 -504 491 -488
rect 615 488 649 504
rect 615 -504 649 -488
rect 773 488 807 504
rect 773 -504 807 -488
rect 931 488 965 504
rect 931 -504 965 -488
rect 1089 488 1123 504
rect 1089 -504 1123 -488
rect 1247 488 1281 504
rect 1247 -504 1281 -488
rect 1405 488 1439 504
rect 1405 -504 1439 -488
rect 1563 488 1597 504
rect 1563 -504 1597 -488
rect -1537 -581 -1521 -547
rect -1481 -581 -1465 -547
rect -1379 -581 -1363 -547
rect -1323 -581 -1307 -547
rect -1221 -581 -1205 -547
rect -1165 -581 -1149 -547
rect -1063 -581 -1047 -547
rect -1007 -581 -991 -547
rect -905 -581 -889 -547
rect -849 -581 -833 -547
rect -747 -581 -731 -547
rect -691 -581 -675 -547
rect -589 -581 -573 -547
rect -533 -581 -517 -547
rect -431 -581 -415 -547
rect -375 -581 -359 -547
rect -273 -581 -257 -547
rect -217 -581 -201 -547
rect -115 -581 -99 -547
rect -59 -581 -43 -547
rect 43 -581 59 -547
rect 99 -581 115 -547
rect 201 -581 217 -547
rect 257 -581 273 -547
rect 359 -581 375 -547
rect 415 -581 431 -547
rect 517 -581 533 -547
rect 573 -581 589 -547
rect 675 -581 691 -547
rect 731 -581 747 -547
rect 833 -581 849 -547
rect 889 -581 905 -547
rect 991 -581 1007 -547
rect 1047 -581 1063 -547
rect 1149 -581 1165 -547
rect 1205 -581 1221 -547
rect 1307 -581 1323 -547
rect 1363 -581 1379 -547
rect 1465 -581 1481 -547
rect 1521 -581 1537 -547
<< viali >>
rect -1597 -488 -1563 488
rect -1439 -488 -1405 488
rect -1281 -488 -1247 488
rect -1123 -488 -1089 488
rect -965 -488 -931 488
rect -807 -488 -773 488
rect -649 -488 -615 488
rect -491 -488 -457 488
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
rect 457 -488 491 488
rect 615 -488 649 488
rect 773 -488 807 488
rect 931 -488 965 488
rect 1089 -488 1123 488
rect 1247 -488 1281 488
rect 1405 -488 1439 488
rect 1563 -488 1597 488
<< metal1 >>
rect -1603 488 -1557 500
rect -1603 -488 -1597 488
rect -1563 -488 -1557 488
rect -1603 -500 -1557 -488
rect -1445 488 -1399 500
rect -1445 -488 -1439 488
rect -1405 -488 -1399 488
rect -1445 -500 -1399 -488
rect -1287 488 -1241 500
rect -1287 -488 -1281 488
rect -1247 -488 -1241 488
rect -1287 -500 -1241 -488
rect -1129 488 -1083 500
rect -1129 -488 -1123 488
rect -1089 -488 -1083 488
rect -1129 -500 -1083 -488
rect -971 488 -925 500
rect -971 -488 -965 488
rect -931 -488 -925 488
rect -971 -500 -925 -488
rect -813 488 -767 500
rect -813 -488 -807 488
rect -773 -488 -767 488
rect -813 -500 -767 -488
rect -655 488 -609 500
rect -655 -488 -649 488
rect -615 -488 -609 488
rect -655 -500 -609 -488
rect -497 488 -451 500
rect -497 -488 -491 488
rect -457 -488 -451 488
rect -497 -500 -451 -488
rect -339 488 -293 500
rect -339 -488 -333 488
rect -299 -488 -293 488
rect -339 -500 -293 -488
rect -181 488 -135 500
rect -181 -488 -175 488
rect -141 -488 -135 488
rect -181 -500 -135 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 135 488 181 500
rect 135 -488 141 488
rect 175 -488 181 488
rect 135 -500 181 -488
rect 293 488 339 500
rect 293 -488 299 488
rect 333 -488 339 488
rect 293 -500 339 -488
rect 451 488 497 500
rect 451 -488 457 488
rect 491 -488 497 488
rect 451 -500 497 -488
rect 609 488 655 500
rect 609 -488 615 488
rect 649 -488 655 488
rect 609 -500 655 -488
rect 767 488 813 500
rect 767 -488 773 488
rect 807 -488 813 488
rect 767 -500 813 -488
rect 925 488 971 500
rect 925 -488 931 488
rect 965 -488 971 488
rect 925 -500 971 -488
rect 1083 488 1129 500
rect 1083 -488 1089 488
rect 1123 -488 1129 488
rect 1083 -500 1129 -488
rect 1241 488 1287 500
rect 1241 -488 1247 488
rect 1281 -488 1287 488
rect 1241 -500 1287 -488
rect 1399 488 1445 500
rect 1399 -488 1405 488
rect 1439 -488 1445 488
rect 1399 -500 1445 -488
rect 1557 488 1603 500
rect 1557 -488 1563 488
rect 1597 -488 1603 488
rect 1557 -500 1603 -488
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string parameters w 5 l 0.5 m 1 nf 20 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
