magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< error_p >>
rect -1668 -300 -1610 300
rect -1370 -300 -1312 300
rect -1072 -300 -1014 300
rect -774 -300 -716 300
rect -476 -300 -418 300
rect -178 -300 -120 300
rect 120 -300 178 300
rect 418 -300 476 300
rect 716 -300 774 300
rect 1014 -300 1072 300
rect 1312 -300 1370 300
rect 1610 -300 1668 300
<< nmoslvt >>
rect -1610 -300 -1370 300
rect -1312 -300 -1072 300
rect -1014 -300 -774 300
rect -716 -300 -476 300
rect -418 -300 -178 300
rect -120 -300 120 300
rect 178 -300 418 300
rect 476 -300 716 300
rect 774 -300 1014 300
rect 1072 -300 1312 300
rect 1370 -300 1610 300
<< ndiff >>
rect -1668 288 -1610 300
rect -1668 -288 -1656 288
rect -1622 -288 -1610 288
rect -1668 -300 -1610 -288
rect -1370 288 -1312 300
rect -1370 -288 -1358 288
rect -1324 -288 -1312 288
rect -1370 -300 -1312 -288
rect -1072 288 -1014 300
rect -1072 -288 -1060 288
rect -1026 -288 -1014 288
rect -1072 -300 -1014 -288
rect -774 288 -716 300
rect -774 -288 -762 288
rect -728 -288 -716 288
rect -774 -300 -716 -288
rect -476 288 -418 300
rect -476 -288 -464 288
rect -430 -288 -418 288
rect -476 -300 -418 -288
rect -178 288 -120 300
rect -178 -288 -166 288
rect -132 -288 -120 288
rect -178 -300 -120 -288
rect 120 288 178 300
rect 120 -288 132 288
rect 166 -288 178 288
rect 120 -300 178 -288
rect 418 288 476 300
rect 418 -288 430 288
rect 464 -288 476 288
rect 418 -300 476 -288
rect 716 288 774 300
rect 716 -288 728 288
rect 762 -288 774 288
rect 716 -300 774 -288
rect 1014 288 1072 300
rect 1014 -288 1026 288
rect 1060 -288 1072 288
rect 1014 -300 1072 -288
rect 1312 288 1370 300
rect 1312 -288 1324 288
rect 1358 -288 1370 288
rect 1312 -300 1370 -288
rect 1610 288 1668 300
rect 1610 -288 1622 288
rect 1656 -288 1668 288
rect 1610 -300 1668 -288
<< ndiffc >>
rect -1656 -288 -1622 288
rect -1358 -288 -1324 288
rect -1060 -288 -1026 288
rect -762 -288 -728 288
rect -464 -288 -430 288
rect -166 -288 -132 288
rect 132 -288 166 288
rect 430 -288 464 288
rect 728 -288 762 288
rect 1026 -288 1060 288
rect 1324 -288 1358 288
rect 1622 -288 1656 288
<< poly >>
rect -1568 372 -1412 388
rect -1568 355 -1552 372
rect -1610 338 -1552 355
rect -1428 355 -1412 372
rect -1270 372 -1114 388
rect -1270 355 -1254 372
rect -1428 338 -1370 355
rect -1610 300 -1370 338
rect -1312 338 -1254 355
rect -1130 355 -1114 372
rect -972 372 -816 388
rect -972 355 -956 372
rect -1130 338 -1072 355
rect -1312 300 -1072 338
rect -1014 338 -956 355
rect -832 355 -816 372
rect -674 372 -518 388
rect -674 355 -658 372
rect -832 338 -774 355
rect -1014 300 -774 338
rect -716 338 -658 355
rect -534 355 -518 372
rect -376 372 -220 388
rect -376 355 -360 372
rect -534 338 -476 355
rect -716 300 -476 338
rect -418 338 -360 355
rect -236 355 -220 372
rect -78 372 78 388
rect -78 355 -62 372
rect -236 338 -178 355
rect -418 300 -178 338
rect -120 338 -62 355
rect 62 355 78 372
rect 220 372 376 388
rect 220 355 236 372
rect 62 338 120 355
rect -120 300 120 338
rect 178 338 236 355
rect 360 355 376 372
rect 518 372 674 388
rect 518 355 534 372
rect 360 338 418 355
rect 178 300 418 338
rect 476 338 534 355
rect 658 355 674 372
rect 816 372 972 388
rect 816 355 832 372
rect 658 338 716 355
rect 476 300 716 338
rect 774 338 832 355
rect 956 355 972 372
rect 1114 372 1270 388
rect 1114 355 1130 372
rect 956 338 1014 355
rect 774 300 1014 338
rect 1072 338 1130 355
rect 1254 355 1270 372
rect 1412 372 1568 388
rect 1412 355 1428 372
rect 1254 338 1312 355
rect 1072 300 1312 338
rect 1370 338 1428 355
rect 1552 355 1568 372
rect 1552 338 1610 355
rect 1370 300 1610 338
rect -1610 -338 -1370 -300
rect -1610 -355 -1552 -338
rect -1568 -372 -1552 -355
rect -1428 -355 -1370 -338
rect -1312 -338 -1072 -300
rect -1312 -355 -1254 -338
rect -1428 -372 -1412 -355
rect -1568 -388 -1412 -372
rect -1270 -372 -1254 -355
rect -1130 -355 -1072 -338
rect -1014 -338 -774 -300
rect -1014 -355 -956 -338
rect -1130 -372 -1114 -355
rect -1270 -388 -1114 -372
rect -972 -372 -956 -355
rect -832 -355 -774 -338
rect -716 -338 -476 -300
rect -716 -355 -658 -338
rect -832 -372 -816 -355
rect -972 -388 -816 -372
rect -674 -372 -658 -355
rect -534 -355 -476 -338
rect -418 -338 -178 -300
rect -418 -355 -360 -338
rect -534 -372 -518 -355
rect -674 -388 -518 -372
rect -376 -372 -360 -355
rect -236 -355 -178 -338
rect -120 -338 120 -300
rect -120 -355 -62 -338
rect -236 -372 -220 -355
rect -376 -388 -220 -372
rect -78 -372 -62 -355
rect 62 -355 120 -338
rect 178 -338 418 -300
rect 178 -355 236 -338
rect 62 -372 78 -355
rect -78 -388 78 -372
rect 220 -372 236 -355
rect 360 -355 418 -338
rect 476 -338 716 -300
rect 476 -355 534 -338
rect 360 -372 376 -355
rect 220 -388 376 -372
rect 518 -372 534 -355
rect 658 -355 716 -338
rect 774 -338 1014 -300
rect 774 -355 832 -338
rect 658 -372 674 -355
rect 518 -388 674 -372
rect 816 -372 832 -355
rect 956 -355 1014 -338
rect 1072 -338 1312 -300
rect 1072 -355 1130 -338
rect 956 -372 972 -355
rect 816 -388 972 -372
rect 1114 -372 1130 -355
rect 1254 -355 1312 -338
rect 1370 -338 1610 -300
rect 1370 -355 1428 -338
rect 1254 -372 1270 -355
rect 1114 -388 1270 -372
rect 1412 -372 1428 -355
rect 1552 -355 1610 -338
rect 1552 -372 1568 -355
rect 1412 -388 1568 -372
<< polycont >>
rect -1552 338 -1428 372
rect -1254 338 -1130 372
rect -956 338 -832 372
rect -658 338 -534 372
rect -360 338 -236 372
rect -62 338 62 372
rect 236 338 360 372
rect 534 338 658 372
rect 832 338 956 372
rect 1130 338 1254 372
rect 1428 338 1552 372
rect -1552 -372 -1428 -338
rect -1254 -372 -1130 -338
rect -956 -372 -832 -338
rect -658 -372 -534 -338
rect -360 -372 -236 -338
rect -62 -372 62 -338
rect 236 -372 360 -338
rect 534 -372 658 -338
rect 832 -372 956 -338
rect 1130 -372 1254 -338
rect 1428 -372 1552 -338
<< locali >>
rect -1568 338 -1552 372
rect -1428 338 -1412 372
rect -1270 338 -1254 372
rect -1130 338 -1114 372
rect -972 338 -956 372
rect -832 338 -816 372
rect -674 338 -658 372
rect -534 338 -518 372
rect -376 338 -360 372
rect -236 338 -220 372
rect -78 338 -62 372
rect 62 338 78 372
rect 220 338 236 372
rect 360 338 376 372
rect 518 338 534 372
rect 658 338 674 372
rect 816 338 832 372
rect 956 338 972 372
rect 1114 338 1130 372
rect 1254 338 1270 372
rect 1412 338 1428 372
rect 1552 338 1568 372
rect -1656 288 -1622 304
rect -1656 -304 -1622 -288
rect -1358 288 -1324 304
rect -1358 -304 -1324 -288
rect -1060 288 -1026 304
rect -1060 -304 -1026 -288
rect -762 288 -728 304
rect -762 -304 -728 -288
rect -464 288 -430 304
rect -464 -304 -430 -288
rect -166 288 -132 304
rect -166 -304 -132 -288
rect 132 288 166 304
rect 132 -304 166 -288
rect 430 288 464 304
rect 430 -304 464 -288
rect 728 288 762 304
rect 728 -304 762 -288
rect 1026 288 1060 304
rect 1026 -304 1060 -288
rect 1324 288 1358 304
rect 1324 -304 1358 -288
rect 1622 288 1656 304
rect 1622 -304 1656 -288
rect -1568 -372 -1552 -338
rect -1428 -372 -1412 -338
rect -1270 -372 -1254 -338
rect -1130 -372 -1114 -338
rect -972 -372 -956 -338
rect -832 -372 -816 -338
rect -674 -372 -658 -338
rect -534 -372 -518 -338
rect -376 -372 -360 -338
rect -236 -372 -220 -338
rect -78 -372 -62 -338
rect 62 -372 78 -338
rect 220 -372 236 -338
rect 360 -372 376 -338
rect 518 -372 534 -338
rect 658 -372 674 -338
rect 816 -372 832 -338
rect 956 -372 972 -338
rect 1114 -372 1130 -338
rect 1254 -372 1270 -338
rect 1412 -372 1428 -338
rect 1552 -372 1568 -338
<< viali >>
rect -1542 338 -1438 372
rect -1244 338 -1140 372
rect -946 338 -842 372
rect -648 338 -544 372
rect -350 338 -246 372
rect -52 338 52 372
rect 246 338 350 372
rect 544 338 648 372
rect 842 338 946 372
rect 1140 338 1244 372
rect 1438 338 1542 372
rect -1656 -288 -1622 288
rect -1358 -288 -1324 288
rect -1060 -288 -1026 288
rect -762 -288 -728 288
rect -464 -288 -430 288
rect -166 -288 -132 288
rect 132 -288 166 288
rect 430 -288 464 288
rect 728 -288 762 288
rect 1026 -288 1060 288
rect 1324 -288 1358 288
rect 1622 -288 1656 288
rect -1542 -372 -1438 -338
rect -1244 -372 -1140 -338
rect -946 -372 -842 -338
rect -648 -372 -544 -338
rect -350 -372 -246 -338
rect -52 -372 52 -338
rect 246 -372 350 -338
rect 544 -372 648 -338
rect 842 -372 946 -338
rect 1140 -372 1244 -338
rect 1438 -372 1542 -338
<< metal1 >>
rect -1554 372 -1426 378
rect -1554 338 -1542 372
rect -1438 338 -1426 372
rect -1554 332 -1426 338
rect -1256 372 -1128 378
rect -1256 338 -1244 372
rect -1140 338 -1128 372
rect -1256 332 -1128 338
rect -958 372 -830 378
rect -958 338 -946 372
rect -842 338 -830 372
rect -958 332 -830 338
rect -660 372 -532 378
rect -660 338 -648 372
rect -544 338 -532 372
rect -660 332 -532 338
rect -362 372 -234 378
rect -362 338 -350 372
rect -246 338 -234 372
rect -362 332 -234 338
rect -64 372 64 378
rect -64 338 -52 372
rect 52 338 64 372
rect -64 332 64 338
rect 234 372 362 378
rect 234 338 246 372
rect 350 338 362 372
rect 234 332 362 338
rect 532 372 660 378
rect 532 338 544 372
rect 648 338 660 372
rect 532 332 660 338
rect 830 372 958 378
rect 830 338 842 372
rect 946 338 958 372
rect 830 332 958 338
rect 1128 372 1256 378
rect 1128 338 1140 372
rect 1244 338 1256 372
rect 1128 332 1256 338
rect 1426 372 1554 378
rect 1426 338 1438 372
rect 1542 338 1554 372
rect 1426 332 1554 338
rect -1662 288 -1616 300
rect -1662 -288 -1656 288
rect -1622 -288 -1616 288
rect -1662 -300 -1616 -288
rect -1364 288 -1318 300
rect -1364 -288 -1358 288
rect -1324 -288 -1318 288
rect -1364 -300 -1318 -288
rect -1066 288 -1020 300
rect -1066 -288 -1060 288
rect -1026 -288 -1020 288
rect -1066 -300 -1020 -288
rect -768 288 -722 300
rect -768 -288 -762 288
rect -728 -288 -722 288
rect -768 -300 -722 -288
rect -470 288 -424 300
rect -470 -288 -464 288
rect -430 -288 -424 288
rect -470 -300 -424 -288
rect -172 288 -126 300
rect -172 -288 -166 288
rect -132 -288 -126 288
rect -172 -300 -126 -288
rect 126 288 172 300
rect 126 -288 132 288
rect 166 -288 172 288
rect 126 -300 172 -288
rect 424 288 470 300
rect 424 -288 430 288
rect 464 -288 470 288
rect 424 -300 470 -288
rect 722 288 768 300
rect 722 -288 728 288
rect 762 -288 768 288
rect 722 -300 768 -288
rect 1020 288 1066 300
rect 1020 -288 1026 288
rect 1060 -288 1066 288
rect 1020 -300 1066 -288
rect 1318 288 1364 300
rect 1318 -288 1324 288
rect 1358 -288 1364 288
rect 1318 -300 1364 -288
rect 1616 288 1662 300
rect 1616 -288 1622 288
rect 1656 -288 1662 288
rect 1616 -300 1662 -288
rect -1554 -338 -1426 -332
rect -1554 -372 -1542 -338
rect -1438 -372 -1426 -338
rect -1554 -378 -1426 -372
rect -1256 -338 -1128 -332
rect -1256 -372 -1244 -338
rect -1140 -372 -1128 -338
rect -1256 -378 -1128 -372
rect -958 -338 -830 -332
rect -958 -372 -946 -338
rect -842 -372 -830 -338
rect -958 -378 -830 -372
rect -660 -338 -532 -332
rect -660 -372 -648 -338
rect -544 -372 -532 -338
rect -660 -378 -532 -372
rect -362 -338 -234 -332
rect -362 -372 -350 -338
rect -246 -372 -234 -338
rect -362 -378 -234 -372
rect -64 -338 64 -332
rect -64 -372 -52 -338
rect 52 -372 64 -338
rect -64 -378 64 -372
rect 234 -338 362 -332
rect 234 -372 246 -338
rect 350 -372 362 -338
rect 234 -378 362 -372
rect 532 -338 660 -332
rect 532 -372 544 -338
rect 648 -372 660 -338
rect 532 -378 660 -372
rect 830 -338 958 -332
rect 830 -372 842 -338
rect 946 -372 958 -338
rect 830 -378 958 -372
rect 1128 -338 1256 -332
rect 1128 -372 1140 -338
rect 1244 -372 1256 -338
rect 1128 -378 1256 -372
rect 1426 -338 1554 -332
rect 1426 -372 1438 -338
rect 1542 -372 1554 -338
rect 1426 -378 1554 -372
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string parameters w 3 l 1.2 m 1 nf 11 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
