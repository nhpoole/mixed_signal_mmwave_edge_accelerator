../../6-sram/outputs/sky130_sram_2kbyte_1rw1r_32x512_8.lef