magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -5176 -1448 5176 1448
<< pwell >>
rect -3916 -126 3916 126
<< nmos >>
rect -3832 -100 -3032 100
rect -2974 -100 -2174 100
rect -2116 -100 -1316 100
rect -1258 -100 -458 100
rect -400 -100 400 100
rect 458 -100 1258 100
rect 1316 -100 2116 100
rect 2174 -100 2974 100
rect 3032 -100 3832 100
<< ndiff >>
rect -3890 85 -3832 100
rect -3890 51 -3878 85
rect -3844 51 -3832 85
rect -3890 17 -3832 51
rect -3890 -17 -3878 17
rect -3844 -17 -3832 17
rect -3890 -51 -3832 -17
rect -3890 -85 -3878 -51
rect -3844 -85 -3832 -51
rect -3890 -100 -3832 -85
rect -3032 85 -2974 100
rect -3032 51 -3020 85
rect -2986 51 -2974 85
rect -3032 17 -2974 51
rect -3032 -17 -3020 17
rect -2986 -17 -2974 17
rect -3032 -51 -2974 -17
rect -3032 -85 -3020 -51
rect -2986 -85 -2974 -51
rect -3032 -100 -2974 -85
rect -2174 85 -2116 100
rect -2174 51 -2162 85
rect -2128 51 -2116 85
rect -2174 17 -2116 51
rect -2174 -17 -2162 17
rect -2128 -17 -2116 17
rect -2174 -51 -2116 -17
rect -2174 -85 -2162 -51
rect -2128 -85 -2116 -51
rect -2174 -100 -2116 -85
rect -1316 85 -1258 100
rect -1316 51 -1304 85
rect -1270 51 -1258 85
rect -1316 17 -1258 51
rect -1316 -17 -1304 17
rect -1270 -17 -1258 17
rect -1316 -51 -1258 -17
rect -1316 -85 -1304 -51
rect -1270 -85 -1258 -51
rect -1316 -100 -1258 -85
rect -458 85 -400 100
rect -458 51 -446 85
rect -412 51 -400 85
rect -458 17 -400 51
rect -458 -17 -446 17
rect -412 -17 -400 17
rect -458 -51 -400 -17
rect -458 -85 -446 -51
rect -412 -85 -400 -51
rect -458 -100 -400 -85
rect 400 85 458 100
rect 400 51 412 85
rect 446 51 458 85
rect 400 17 458 51
rect 400 -17 412 17
rect 446 -17 458 17
rect 400 -51 458 -17
rect 400 -85 412 -51
rect 446 -85 458 -51
rect 400 -100 458 -85
rect 1258 85 1316 100
rect 1258 51 1270 85
rect 1304 51 1316 85
rect 1258 17 1316 51
rect 1258 -17 1270 17
rect 1304 -17 1316 17
rect 1258 -51 1316 -17
rect 1258 -85 1270 -51
rect 1304 -85 1316 -51
rect 1258 -100 1316 -85
rect 2116 85 2174 100
rect 2116 51 2128 85
rect 2162 51 2174 85
rect 2116 17 2174 51
rect 2116 -17 2128 17
rect 2162 -17 2174 17
rect 2116 -51 2174 -17
rect 2116 -85 2128 -51
rect 2162 -85 2174 -51
rect 2116 -100 2174 -85
rect 2974 85 3032 100
rect 2974 51 2986 85
rect 3020 51 3032 85
rect 2974 17 3032 51
rect 2974 -17 2986 17
rect 3020 -17 3032 17
rect 2974 -51 3032 -17
rect 2974 -85 2986 -51
rect 3020 -85 3032 -51
rect 2974 -100 3032 -85
rect 3832 85 3890 100
rect 3832 51 3844 85
rect 3878 51 3890 85
rect 3832 17 3890 51
rect 3832 -17 3844 17
rect 3878 -17 3890 17
rect 3832 -51 3890 -17
rect 3832 -85 3844 -51
rect 3878 -85 3890 -51
rect 3832 -100 3890 -85
<< ndiffc >>
rect -3878 51 -3844 85
rect -3878 -17 -3844 17
rect -3878 -85 -3844 -51
rect -3020 51 -2986 85
rect -3020 -17 -2986 17
rect -3020 -85 -2986 -51
rect -2162 51 -2128 85
rect -2162 -17 -2128 17
rect -2162 -85 -2128 -51
rect -1304 51 -1270 85
rect -1304 -17 -1270 17
rect -1304 -85 -1270 -51
rect -446 51 -412 85
rect -446 -17 -412 17
rect -446 -85 -412 -51
rect 412 51 446 85
rect 412 -17 446 17
rect 412 -85 446 -51
rect 1270 51 1304 85
rect 1270 -17 1304 17
rect 1270 -85 1304 -51
rect 2128 51 2162 85
rect 2128 -17 2162 17
rect 2128 -85 2162 -51
rect 2986 51 3020 85
rect 2986 -17 3020 17
rect 2986 -85 3020 -51
rect 3844 51 3878 85
rect 3844 -17 3878 17
rect 3844 -85 3878 -51
<< poly >>
rect -3678 172 -3186 188
rect -3678 155 -3653 172
rect -3832 138 -3653 155
rect -3619 138 -3585 172
rect -3551 138 -3517 172
rect -3483 138 -3449 172
rect -3415 138 -3381 172
rect -3347 138 -3313 172
rect -3279 138 -3245 172
rect -3211 155 -3186 172
rect -2820 172 -2328 188
rect -2820 155 -2795 172
rect -3211 138 -3032 155
rect -3832 100 -3032 138
rect -2974 138 -2795 155
rect -2761 138 -2727 172
rect -2693 138 -2659 172
rect -2625 138 -2591 172
rect -2557 138 -2523 172
rect -2489 138 -2455 172
rect -2421 138 -2387 172
rect -2353 155 -2328 172
rect -1962 172 -1470 188
rect -1962 155 -1937 172
rect -2353 138 -2174 155
rect -2974 100 -2174 138
rect -2116 138 -1937 155
rect -1903 138 -1869 172
rect -1835 138 -1801 172
rect -1767 138 -1733 172
rect -1699 138 -1665 172
rect -1631 138 -1597 172
rect -1563 138 -1529 172
rect -1495 155 -1470 172
rect -1104 172 -612 188
rect -1104 155 -1079 172
rect -1495 138 -1316 155
rect -2116 100 -1316 138
rect -1258 138 -1079 155
rect -1045 138 -1011 172
rect -977 138 -943 172
rect -909 138 -875 172
rect -841 138 -807 172
rect -773 138 -739 172
rect -705 138 -671 172
rect -637 155 -612 172
rect -246 172 246 188
rect -246 155 -221 172
rect -637 138 -458 155
rect -1258 100 -458 138
rect -400 138 -221 155
rect -187 138 -153 172
rect -119 138 -85 172
rect -51 138 -17 172
rect 17 138 51 172
rect 85 138 119 172
rect 153 138 187 172
rect 221 155 246 172
rect 612 172 1104 188
rect 612 155 637 172
rect 221 138 400 155
rect -400 100 400 138
rect 458 138 637 155
rect 671 138 705 172
rect 739 138 773 172
rect 807 138 841 172
rect 875 138 909 172
rect 943 138 977 172
rect 1011 138 1045 172
rect 1079 155 1104 172
rect 1470 172 1962 188
rect 1470 155 1495 172
rect 1079 138 1258 155
rect 458 100 1258 138
rect 1316 138 1495 155
rect 1529 138 1563 172
rect 1597 138 1631 172
rect 1665 138 1699 172
rect 1733 138 1767 172
rect 1801 138 1835 172
rect 1869 138 1903 172
rect 1937 155 1962 172
rect 2328 172 2820 188
rect 2328 155 2353 172
rect 1937 138 2116 155
rect 1316 100 2116 138
rect 2174 138 2353 155
rect 2387 138 2421 172
rect 2455 138 2489 172
rect 2523 138 2557 172
rect 2591 138 2625 172
rect 2659 138 2693 172
rect 2727 138 2761 172
rect 2795 155 2820 172
rect 3186 172 3678 188
rect 3186 155 3211 172
rect 2795 138 2974 155
rect 2174 100 2974 138
rect 3032 138 3211 155
rect 3245 138 3279 172
rect 3313 138 3347 172
rect 3381 138 3415 172
rect 3449 138 3483 172
rect 3517 138 3551 172
rect 3585 138 3619 172
rect 3653 155 3678 172
rect 3653 138 3832 155
rect 3032 100 3832 138
rect -3832 -138 -3032 -100
rect -3832 -155 -3653 -138
rect -3678 -172 -3653 -155
rect -3619 -172 -3585 -138
rect -3551 -172 -3517 -138
rect -3483 -172 -3449 -138
rect -3415 -172 -3381 -138
rect -3347 -172 -3313 -138
rect -3279 -172 -3245 -138
rect -3211 -155 -3032 -138
rect -2974 -138 -2174 -100
rect -2974 -155 -2795 -138
rect -3211 -172 -3186 -155
rect -3678 -188 -3186 -172
rect -2820 -172 -2795 -155
rect -2761 -172 -2727 -138
rect -2693 -172 -2659 -138
rect -2625 -172 -2591 -138
rect -2557 -172 -2523 -138
rect -2489 -172 -2455 -138
rect -2421 -172 -2387 -138
rect -2353 -155 -2174 -138
rect -2116 -138 -1316 -100
rect -2116 -155 -1937 -138
rect -2353 -172 -2328 -155
rect -2820 -188 -2328 -172
rect -1962 -172 -1937 -155
rect -1903 -172 -1869 -138
rect -1835 -172 -1801 -138
rect -1767 -172 -1733 -138
rect -1699 -172 -1665 -138
rect -1631 -172 -1597 -138
rect -1563 -172 -1529 -138
rect -1495 -155 -1316 -138
rect -1258 -138 -458 -100
rect -1258 -155 -1079 -138
rect -1495 -172 -1470 -155
rect -1962 -188 -1470 -172
rect -1104 -172 -1079 -155
rect -1045 -172 -1011 -138
rect -977 -172 -943 -138
rect -909 -172 -875 -138
rect -841 -172 -807 -138
rect -773 -172 -739 -138
rect -705 -172 -671 -138
rect -637 -155 -458 -138
rect -400 -138 400 -100
rect -400 -155 -221 -138
rect -637 -172 -612 -155
rect -1104 -188 -612 -172
rect -246 -172 -221 -155
rect -187 -172 -153 -138
rect -119 -172 -85 -138
rect -51 -172 -17 -138
rect 17 -172 51 -138
rect 85 -172 119 -138
rect 153 -172 187 -138
rect 221 -155 400 -138
rect 458 -138 1258 -100
rect 458 -155 637 -138
rect 221 -172 246 -155
rect -246 -188 246 -172
rect 612 -172 637 -155
rect 671 -172 705 -138
rect 739 -172 773 -138
rect 807 -172 841 -138
rect 875 -172 909 -138
rect 943 -172 977 -138
rect 1011 -172 1045 -138
rect 1079 -155 1258 -138
rect 1316 -138 2116 -100
rect 1316 -155 1495 -138
rect 1079 -172 1104 -155
rect 612 -188 1104 -172
rect 1470 -172 1495 -155
rect 1529 -172 1563 -138
rect 1597 -172 1631 -138
rect 1665 -172 1699 -138
rect 1733 -172 1767 -138
rect 1801 -172 1835 -138
rect 1869 -172 1903 -138
rect 1937 -155 2116 -138
rect 2174 -138 2974 -100
rect 2174 -155 2353 -138
rect 1937 -172 1962 -155
rect 1470 -188 1962 -172
rect 2328 -172 2353 -155
rect 2387 -172 2421 -138
rect 2455 -172 2489 -138
rect 2523 -172 2557 -138
rect 2591 -172 2625 -138
rect 2659 -172 2693 -138
rect 2727 -172 2761 -138
rect 2795 -155 2974 -138
rect 3032 -138 3832 -100
rect 3032 -155 3211 -138
rect 2795 -172 2820 -155
rect 2328 -188 2820 -172
rect 3186 -172 3211 -155
rect 3245 -172 3279 -138
rect 3313 -172 3347 -138
rect 3381 -172 3415 -138
rect 3449 -172 3483 -138
rect 3517 -172 3551 -138
rect 3585 -172 3619 -138
rect 3653 -155 3832 -138
rect 3653 -172 3678 -155
rect 3186 -188 3678 -172
<< polycont >>
rect -3653 138 -3619 172
rect -3585 138 -3551 172
rect -3517 138 -3483 172
rect -3449 138 -3415 172
rect -3381 138 -3347 172
rect -3313 138 -3279 172
rect -3245 138 -3211 172
rect -2795 138 -2761 172
rect -2727 138 -2693 172
rect -2659 138 -2625 172
rect -2591 138 -2557 172
rect -2523 138 -2489 172
rect -2455 138 -2421 172
rect -2387 138 -2353 172
rect -1937 138 -1903 172
rect -1869 138 -1835 172
rect -1801 138 -1767 172
rect -1733 138 -1699 172
rect -1665 138 -1631 172
rect -1597 138 -1563 172
rect -1529 138 -1495 172
rect -1079 138 -1045 172
rect -1011 138 -977 172
rect -943 138 -909 172
rect -875 138 -841 172
rect -807 138 -773 172
rect -739 138 -705 172
rect -671 138 -637 172
rect -221 138 -187 172
rect -153 138 -119 172
rect -85 138 -51 172
rect -17 138 17 172
rect 51 138 85 172
rect 119 138 153 172
rect 187 138 221 172
rect 637 138 671 172
rect 705 138 739 172
rect 773 138 807 172
rect 841 138 875 172
rect 909 138 943 172
rect 977 138 1011 172
rect 1045 138 1079 172
rect 1495 138 1529 172
rect 1563 138 1597 172
rect 1631 138 1665 172
rect 1699 138 1733 172
rect 1767 138 1801 172
rect 1835 138 1869 172
rect 1903 138 1937 172
rect 2353 138 2387 172
rect 2421 138 2455 172
rect 2489 138 2523 172
rect 2557 138 2591 172
rect 2625 138 2659 172
rect 2693 138 2727 172
rect 2761 138 2795 172
rect 3211 138 3245 172
rect 3279 138 3313 172
rect 3347 138 3381 172
rect 3415 138 3449 172
rect 3483 138 3517 172
rect 3551 138 3585 172
rect 3619 138 3653 172
rect -3653 -172 -3619 -138
rect -3585 -172 -3551 -138
rect -3517 -172 -3483 -138
rect -3449 -172 -3415 -138
rect -3381 -172 -3347 -138
rect -3313 -172 -3279 -138
rect -3245 -172 -3211 -138
rect -2795 -172 -2761 -138
rect -2727 -172 -2693 -138
rect -2659 -172 -2625 -138
rect -2591 -172 -2557 -138
rect -2523 -172 -2489 -138
rect -2455 -172 -2421 -138
rect -2387 -172 -2353 -138
rect -1937 -172 -1903 -138
rect -1869 -172 -1835 -138
rect -1801 -172 -1767 -138
rect -1733 -172 -1699 -138
rect -1665 -172 -1631 -138
rect -1597 -172 -1563 -138
rect -1529 -172 -1495 -138
rect -1079 -172 -1045 -138
rect -1011 -172 -977 -138
rect -943 -172 -909 -138
rect -875 -172 -841 -138
rect -807 -172 -773 -138
rect -739 -172 -705 -138
rect -671 -172 -637 -138
rect -221 -172 -187 -138
rect -153 -172 -119 -138
rect -85 -172 -51 -138
rect -17 -172 17 -138
rect 51 -172 85 -138
rect 119 -172 153 -138
rect 187 -172 221 -138
rect 637 -172 671 -138
rect 705 -172 739 -138
rect 773 -172 807 -138
rect 841 -172 875 -138
rect 909 -172 943 -138
rect 977 -172 1011 -138
rect 1045 -172 1079 -138
rect 1495 -172 1529 -138
rect 1563 -172 1597 -138
rect 1631 -172 1665 -138
rect 1699 -172 1733 -138
rect 1767 -172 1801 -138
rect 1835 -172 1869 -138
rect 1903 -172 1937 -138
rect 2353 -172 2387 -138
rect 2421 -172 2455 -138
rect 2489 -172 2523 -138
rect 2557 -172 2591 -138
rect 2625 -172 2659 -138
rect 2693 -172 2727 -138
rect 2761 -172 2795 -138
rect 3211 -172 3245 -138
rect 3279 -172 3313 -138
rect 3347 -172 3381 -138
rect 3415 -172 3449 -138
rect 3483 -172 3517 -138
rect 3551 -172 3585 -138
rect 3619 -172 3653 -138
<< locali >>
rect -3678 138 -3653 172
rect -3619 138 -3593 172
rect -3551 138 -3521 172
rect -3483 138 -3449 172
rect -3415 138 -3381 172
rect -3343 138 -3313 172
rect -3271 138 -3245 172
rect -3211 138 -3186 172
rect -2820 138 -2795 172
rect -2761 138 -2735 172
rect -2693 138 -2663 172
rect -2625 138 -2591 172
rect -2557 138 -2523 172
rect -2485 138 -2455 172
rect -2413 138 -2387 172
rect -2353 138 -2328 172
rect -1962 138 -1937 172
rect -1903 138 -1877 172
rect -1835 138 -1805 172
rect -1767 138 -1733 172
rect -1699 138 -1665 172
rect -1627 138 -1597 172
rect -1555 138 -1529 172
rect -1495 138 -1470 172
rect -1104 138 -1079 172
rect -1045 138 -1019 172
rect -977 138 -947 172
rect -909 138 -875 172
rect -841 138 -807 172
rect -769 138 -739 172
rect -697 138 -671 172
rect -637 138 -612 172
rect -246 138 -221 172
rect -187 138 -161 172
rect -119 138 -89 172
rect -51 138 -17 172
rect 17 138 51 172
rect 89 138 119 172
rect 161 138 187 172
rect 221 138 246 172
rect 612 138 637 172
rect 671 138 697 172
rect 739 138 769 172
rect 807 138 841 172
rect 875 138 909 172
rect 947 138 977 172
rect 1019 138 1045 172
rect 1079 138 1104 172
rect 1470 138 1495 172
rect 1529 138 1555 172
rect 1597 138 1627 172
rect 1665 138 1699 172
rect 1733 138 1767 172
rect 1805 138 1835 172
rect 1877 138 1903 172
rect 1937 138 1962 172
rect 2328 138 2353 172
rect 2387 138 2413 172
rect 2455 138 2485 172
rect 2523 138 2557 172
rect 2591 138 2625 172
rect 2663 138 2693 172
rect 2735 138 2761 172
rect 2795 138 2820 172
rect 3186 138 3211 172
rect 3245 138 3271 172
rect 3313 138 3343 172
rect 3381 138 3415 172
rect 3449 138 3483 172
rect 3521 138 3551 172
rect 3593 138 3619 172
rect 3653 138 3678 172
rect -3878 85 -3844 104
rect -3878 17 -3844 19
rect -3878 -19 -3844 -17
rect -3878 -104 -3844 -85
rect -3020 85 -2986 104
rect -3020 17 -2986 19
rect -3020 -19 -2986 -17
rect -3020 -104 -2986 -85
rect -2162 85 -2128 104
rect -2162 17 -2128 19
rect -2162 -19 -2128 -17
rect -2162 -104 -2128 -85
rect -1304 85 -1270 104
rect -1304 17 -1270 19
rect -1304 -19 -1270 -17
rect -1304 -104 -1270 -85
rect -446 85 -412 104
rect -446 17 -412 19
rect -446 -19 -412 -17
rect -446 -104 -412 -85
rect 412 85 446 104
rect 412 17 446 19
rect 412 -19 446 -17
rect 412 -104 446 -85
rect 1270 85 1304 104
rect 1270 17 1304 19
rect 1270 -19 1304 -17
rect 1270 -104 1304 -85
rect 2128 85 2162 104
rect 2128 17 2162 19
rect 2128 -19 2162 -17
rect 2128 -104 2162 -85
rect 2986 85 3020 104
rect 2986 17 3020 19
rect 2986 -19 3020 -17
rect 2986 -104 3020 -85
rect 3844 85 3878 104
rect 3844 17 3878 19
rect 3844 -19 3878 -17
rect 3844 -104 3878 -85
rect -3678 -172 -3653 -138
rect -3619 -172 -3593 -138
rect -3551 -172 -3521 -138
rect -3483 -172 -3449 -138
rect -3415 -172 -3381 -138
rect -3343 -172 -3313 -138
rect -3271 -172 -3245 -138
rect -3211 -172 -3186 -138
rect -2820 -172 -2795 -138
rect -2761 -172 -2735 -138
rect -2693 -172 -2663 -138
rect -2625 -172 -2591 -138
rect -2557 -172 -2523 -138
rect -2485 -172 -2455 -138
rect -2413 -172 -2387 -138
rect -2353 -172 -2328 -138
rect -1962 -172 -1937 -138
rect -1903 -172 -1877 -138
rect -1835 -172 -1805 -138
rect -1767 -172 -1733 -138
rect -1699 -172 -1665 -138
rect -1627 -172 -1597 -138
rect -1555 -172 -1529 -138
rect -1495 -172 -1470 -138
rect -1104 -172 -1079 -138
rect -1045 -172 -1019 -138
rect -977 -172 -947 -138
rect -909 -172 -875 -138
rect -841 -172 -807 -138
rect -769 -172 -739 -138
rect -697 -172 -671 -138
rect -637 -172 -612 -138
rect -246 -172 -221 -138
rect -187 -172 -161 -138
rect -119 -172 -89 -138
rect -51 -172 -17 -138
rect 17 -172 51 -138
rect 89 -172 119 -138
rect 161 -172 187 -138
rect 221 -172 246 -138
rect 612 -172 637 -138
rect 671 -172 697 -138
rect 739 -172 769 -138
rect 807 -172 841 -138
rect 875 -172 909 -138
rect 947 -172 977 -138
rect 1019 -172 1045 -138
rect 1079 -172 1104 -138
rect 1470 -172 1495 -138
rect 1529 -172 1555 -138
rect 1597 -172 1627 -138
rect 1665 -172 1699 -138
rect 1733 -172 1767 -138
rect 1805 -172 1835 -138
rect 1877 -172 1903 -138
rect 1937 -172 1962 -138
rect 2328 -172 2353 -138
rect 2387 -172 2413 -138
rect 2455 -172 2485 -138
rect 2523 -172 2557 -138
rect 2591 -172 2625 -138
rect 2663 -172 2693 -138
rect 2735 -172 2761 -138
rect 2795 -172 2820 -138
rect 3186 -172 3211 -138
rect 3245 -172 3271 -138
rect 3313 -172 3343 -138
rect 3381 -172 3415 -138
rect 3449 -172 3483 -138
rect 3521 -172 3551 -138
rect 3593 -172 3619 -138
rect 3653 -172 3678 -138
<< viali >>
rect -3593 138 -3585 172
rect -3585 138 -3559 172
rect -3521 138 -3517 172
rect -3517 138 -3487 172
rect -3449 138 -3415 172
rect -3377 138 -3347 172
rect -3347 138 -3343 172
rect -3305 138 -3279 172
rect -3279 138 -3271 172
rect -2735 138 -2727 172
rect -2727 138 -2701 172
rect -2663 138 -2659 172
rect -2659 138 -2629 172
rect -2591 138 -2557 172
rect -2519 138 -2489 172
rect -2489 138 -2485 172
rect -2447 138 -2421 172
rect -2421 138 -2413 172
rect -1877 138 -1869 172
rect -1869 138 -1843 172
rect -1805 138 -1801 172
rect -1801 138 -1771 172
rect -1733 138 -1699 172
rect -1661 138 -1631 172
rect -1631 138 -1627 172
rect -1589 138 -1563 172
rect -1563 138 -1555 172
rect -1019 138 -1011 172
rect -1011 138 -985 172
rect -947 138 -943 172
rect -943 138 -913 172
rect -875 138 -841 172
rect -803 138 -773 172
rect -773 138 -769 172
rect -731 138 -705 172
rect -705 138 -697 172
rect -161 138 -153 172
rect -153 138 -127 172
rect -89 138 -85 172
rect -85 138 -55 172
rect -17 138 17 172
rect 55 138 85 172
rect 85 138 89 172
rect 127 138 153 172
rect 153 138 161 172
rect 697 138 705 172
rect 705 138 731 172
rect 769 138 773 172
rect 773 138 803 172
rect 841 138 875 172
rect 913 138 943 172
rect 943 138 947 172
rect 985 138 1011 172
rect 1011 138 1019 172
rect 1555 138 1563 172
rect 1563 138 1589 172
rect 1627 138 1631 172
rect 1631 138 1661 172
rect 1699 138 1733 172
rect 1771 138 1801 172
rect 1801 138 1805 172
rect 1843 138 1869 172
rect 1869 138 1877 172
rect 2413 138 2421 172
rect 2421 138 2447 172
rect 2485 138 2489 172
rect 2489 138 2519 172
rect 2557 138 2591 172
rect 2629 138 2659 172
rect 2659 138 2663 172
rect 2701 138 2727 172
rect 2727 138 2735 172
rect 3271 138 3279 172
rect 3279 138 3305 172
rect 3343 138 3347 172
rect 3347 138 3377 172
rect 3415 138 3449 172
rect 3487 138 3517 172
rect 3517 138 3521 172
rect 3559 138 3585 172
rect 3585 138 3593 172
rect -3878 51 -3844 53
rect -3878 19 -3844 51
rect -3878 -51 -3844 -19
rect -3878 -53 -3844 -51
rect -3020 51 -2986 53
rect -3020 19 -2986 51
rect -3020 -51 -2986 -19
rect -3020 -53 -2986 -51
rect -2162 51 -2128 53
rect -2162 19 -2128 51
rect -2162 -51 -2128 -19
rect -2162 -53 -2128 -51
rect -1304 51 -1270 53
rect -1304 19 -1270 51
rect -1304 -51 -1270 -19
rect -1304 -53 -1270 -51
rect -446 51 -412 53
rect -446 19 -412 51
rect -446 -51 -412 -19
rect -446 -53 -412 -51
rect 412 51 446 53
rect 412 19 446 51
rect 412 -51 446 -19
rect 412 -53 446 -51
rect 1270 51 1304 53
rect 1270 19 1304 51
rect 1270 -51 1304 -19
rect 1270 -53 1304 -51
rect 2128 51 2162 53
rect 2128 19 2162 51
rect 2128 -51 2162 -19
rect 2128 -53 2162 -51
rect 2986 51 3020 53
rect 2986 19 3020 51
rect 2986 -51 3020 -19
rect 2986 -53 3020 -51
rect 3844 51 3878 53
rect 3844 19 3878 51
rect 3844 -51 3878 -19
rect 3844 -53 3878 -51
rect -3593 -172 -3585 -138
rect -3585 -172 -3559 -138
rect -3521 -172 -3517 -138
rect -3517 -172 -3487 -138
rect -3449 -172 -3415 -138
rect -3377 -172 -3347 -138
rect -3347 -172 -3343 -138
rect -3305 -172 -3279 -138
rect -3279 -172 -3271 -138
rect -2735 -172 -2727 -138
rect -2727 -172 -2701 -138
rect -2663 -172 -2659 -138
rect -2659 -172 -2629 -138
rect -2591 -172 -2557 -138
rect -2519 -172 -2489 -138
rect -2489 -172 -2485 -138
rect -2447 -172 -2421 -138
rect -2421 -172 -2413 -138
rect -1877 -172 -1869 -138
rect -1869 -172 -1843 -138
rect -1805 -172 -1801 -138
rect -1801 -172 -1771 -138
rect -1733 -172 -1699 -138
rect -1661 -172 -1631 -138
rect -1631 -172 -1627 -138
rect -1589 -172 -1563 -138
rect -1563 -172 -1555 -138
rect -1019 -172 -1011 -138
rect -1011 -172 -985 -138
rect -947 -172 -943 -138
rect -943 -172 -913 -138
rect -875 -172 -841 -138
rect -803 -172 -773 -138
rect -773 -172 -769 -138
rect -731 -172 -705 -138
rect -705 -172 -697 -138
rect -161 -172 -153 -138
rect -153 -172 -127 -138
rect -89 -172 -85 -138
rect -85 -172 -55 -138
rect -17 -172 17 -138
rect 55 -172 85 -138
rect 85 -172 89 -138
rect 127 -172 153 -138
rect 153 -172 161 -138
rect 697 -172 705 -138
rect 705 -172 731 -138
rect 769 -172 773 -138
rect 773 -172 803 -138
rect 841 -172 875 -138
rect 913 -172 943 -138
rect 943 -172 947 -138
rect 985 -172 1011 -138
rect 1011 -172 1019 -138
rect 1555 -172 1563 -138
rect 1563 -172 1589 -138
rect 1627 -172 1631 -138
rect 1631 -172 1661 -138
rect 1699 -172 1733 -138
rect 1771 -172 1801 -138
rect 1801 -172 1805 -138
rect 1843 -172 1869 -138
rect 1869 -172 1877 -138
rect 2413 -172 2421 -138
rect 2421 -172 2447 -138
rect 2485 -172 2489 -138
rect 2489 -172 2519 -138
rect 2557 -172 2591 -138
rect 2629 -172 2659 -138
rect 2659 -172 2663 -138
rect 2701 -172 2727 -138
rect 2727 -172 2735 -138
rect 3271 -172 3279 -138
rect 3279 -172 3305 -138
rect 3343 -172 3347 -138
rect 3347 -172 3377 -138
rect 3415 -172 3449 -138
rect 3487 -172 3517 -138
rect 3517 -172 3521 -138
rect 3559 -172 3585 -138
rect 3585 -172 3593 -138
<< metal1 >>
rect -3636 172 -3228 178
rect -3636 138 -3593 172
rect -3559 138 -3521 172
rect -3487 138 -3449 172
rect -3415 138 -3377 172
rect -3343 138 -3305 172
rect -3271 138 -3228 172
rect -3636 132 -3228 138
rect -2778 172 -2370 178
rect -2778 138 -2735 172
rect -2701 138 -2663 172
rect -2629 138 -2591 172
rect -2557 138 -2519 172
rect -2485 138 -2447 172
rect -2413 138 -2370 172
rect -2778 132 -2370 138
rect -1920 172 -1512 178
rect -1920 138 -1877 172
rect -1843 138 -1805 172
rect -1771 138 -1733 172
rect -1699 138 -1661 172
rect -1627 138 -1589 172
rect -1555 138 -1512 172
rect -1920 132 -1512 138
rect -1062 172 -654 178
rect -1062 138 -1019 172
rect -985 138 -947 172
rect -913 138 -875 172
rect -841 138 -803 172
rect -769 138 -731 172
rect -697 138 -654 172
rect -1062 132 -654 138
rect -204 172 204 178
rect -204 138 -161 172
rect -127 138 -89 172
rect -55 138 -17 172
rect 17 138 55 172
rect 89 138 127 172
rect 161 138 204 172
rect -204 132 204 138
rect 654 172 1062 178
rect 654 138 697 172
rect 731 138 769 172
rect 803 138 841 172
rect 875 138 913 172
rect 947 138 985 172
rect 1019 138 1062 172
rect 654 132 1062 138
rect 1512 172 1920 178
rect 1512 138 1555 172
rect 1589 138 1627 172
rect 1661 138 1699 172
rect 1733 138 1771 172
rect 1805 138 1843 172
rect 1877 138 1920 172
rect 1512 132 1920 138
rect 2370 172 2778 178
rect 2370 138 2413 172
rect 2447 138 2485 172
rect 2519 138 2557 172
rect 2591 138 2629 172
rect 2663 138 2701 172
rect 2735 138 2778 172
rect 2370 132 2778 138
rect 3228 172 3636 178
rect 3228 138 3271 172
rect 3305 138 3343 172
rect 3377 138 3415 172
rect 3449 138 3487 172
rect 3521 138 3559 172
rect 3593 138 3636 172
rect 3228 132 3636 138
rect -3884 53 -3838 100
rect -3884 19 -3878 53
rect -3844 19 -3838 53
rect -3884 -19 -3838 19
rect -3884 -53 -3878 -19
rect -3844 -53 -3838 -19
rect -3884 -100 -3838 -53
rect -3026 53 -2980 100
rect -3026 19 -3020 53
rect -2986 19 -2980 53
rect -3026 -19 -2980 19
rect -3026 -53 -3020 -19
rect -2986 -53 -2980 -19
rect -3026 -100 -2980 -53
rect -2168 53 -2122 100
rect -2168 19 -2162 53
rect -2128 19 -2122 53
rect -2168 -19 -2122 19
rect -2168 -53 -2162 -19
rect -2128 -53 -2122 -19
rect -2168 -100 -2122 -53
rect -1310 53 -1264 100
rect -1310 19 -1304 53
rect -1270 19 -1264 53
rect -1310 -19 -1264 19
rect -1310 -53 -1304 -19
rect -1270 -53 -1264 -19
rect -1310 -100 -1264 -53
rect -452 53 -406 100
rect -452 19 -446 53
rect -412 19 -406 53
rect -452 -19 -406 19
rect -452 -53 -446 -19
rect -412 -53 -406 -19
rect -452 -100 -406 -53
rect 406 53 452 100
rect 406 19 412 53
rect 446 19 452 53
rect 406 -19 452 19
rect 406 -53 412 -19
rect 446 -53 452 -19
rect 406 -100 452 -53
rect 1264 53 1310 100
rect 1264 19 1270 53
rect 1304 19 1310 53
rect 1264 -19 1310 19
rect 1264 -53 1270 -19
rect 1304 -53 1310 -19
rect 1264 -100 1310 -53
rect 2122 53 2168 100
rect 2122 19 2128 53
rect 2162 19 2168 53
rect 2122 -19 2168 19
rect 2122 -53 2128 -19
rect 2162 -53 2168 -19
rect 2122 -100 2168 -53
rect 2980 53 3026 100
rect 2980 19 2986 53
rect 3020 19 3026 53
rect 2980 -19 3026 19
rect 2980 -53 2986 -19
rect 3020 -53 3026 -19
rect 2980 -100 3026 -53
rect 3838 53 3884 100
rect 3838 19 3844 53
rect 3878 19 3884 53
rect 3838 -19 3884 19
rect 3838 -53 3844 -19
rect 3878 -53 3884 -19
rect 3838 -100 3884 -53
rect -3636 -138 -3228 -132
rect -3636 -172 -3593 -138
rect -3559 -172 -3521 -138
rect -3487 -172 -3449 -138
rect -3415 -172 -3377 -138
rect -3343 -172 -3305 -138
rect -3271 -172 -3228 -138
rect -3636 -178 -3228 -172
rect -2778 -138 -2370 -132
rect -2778 -172 -2735 -138
rect -2701 -172 -2663 -138
rect -2629 -172 -2591 -138
rect -2557 -172 -2519 -138
rect -2485 -172 -2447 -138
rect -2413 -172 -2370 -138
rect -2778 -178 -2370 -172
rect -1920 -138 -1512 -132
rect -1920 -172 -1877 -138
rect -1843 -172 -1805 -138
rect -1771 -172 -1733 -138
rect -1699 -172 -1661 -138
rect -1627 -172 -1589 -138
rect -1555 -172 -1512 -138
rect -1920 -178 -1512 -172
rect -1062 -138 -654 -132
rect -1062 -172 -1019 -138
rect -985 -172 -947 -138
rect -913 -172 -875 -138
rect -841 -172 -803 -138
rect -769 -172 -731 -138
rect -697 -172 -654 -138
rect -1062 -178 -654 -172
rect -204 -138 204 -132
rect -204 -172 -161 -138
rect -127 -172 -89 -138
rect -55 -172 -17 -138
rect 17 -172 55 -138
rect 89 -172 127 -138
rect 161 -172 204 -138
rect -204 -178 204 -172
rect 654 -138 1062 -132
rect 654 -172 697 -138
rect 731 -172 769 -138
rect 803 -172 841 -138
rect 875 -172 913 -138
rect 947 -172 985 -138
rect 1019 -172 1062 -138
rect 654 -178 1062 -172
rect 1512 -138 1920 -132
rect 1512 -172 1555 -138
rect 1589 -172 1627 -138
rect 1661 -172 1699 -138
rect 1733 -172 1771 -138
rect 1805 -172 1843 -138
rect 1877 -172 1920 -138
rect 1512 -178 1920 -172
rect 2370 -138 2778 -132
rect 2370 -172 2413 -138
rect 2447 -172 2485 -138
rect 2519 -172 2557 -138
rect 2591 -172 2629 -138
rect 2663 -172 2701 -138
rect 2735 -172 2778 -138
rect 2370 -178 2778 -172
rect 3228 -138 3636 -132
rect 3228 -172 3271 -138
rect 3305 -172 3343 -138
rect 3377 -172 3415 -138
rect 3449 -172 3487 -138
rect 3521 -172 3559 -138
rect 3593 -172 3636 -138
rect 3228 -178 3636 -172
<< end >>
