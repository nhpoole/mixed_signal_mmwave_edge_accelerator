magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1260 -1272 82506 2028
<< metal1 >>
rect 816 0 844 754
rect 1280 0 1308 754
rect 1440 0 1468 754
rect 1904 0 1932 754
rect 2064 0 2092 754
rect 2528 0 2556 754
rect 2688 0 2716 754
rect 3152 0 3180 754
rect 3312 0 3340 754
rect 3776 0 3804 754
rect 3936 0 3964 754
rect 4400 0 4428 754
rect 4560 0 4588 754
rect 5024 0 5052 754
rect 5184 0 5212 754
rect 5648 0 5676 754
rect 5808 0 5836 754
rect 6272 0 6300 754
rect 6432 0 6460 754
rect 6896 0 6924 754
rect 7056 0 7084 754
rect 7520 0 7548 754
rect 7680 0 7708 754
rect 8144 0 8172 754
rect 8304 0 8332 754
rect 8768 0 8796 754
rect 8928 0 8956 754
rect 9392 0 9420 754
rect 9552 0 9580 754
rect 10016 0 10044 754
rect 10176 0 10204 754
rect 10640 0 10668 754
rect 10800 0 10828 754
rect 11264 0 11292 754
rect 11424 0 11452 754
rect 11888 0 11916 754
rect 12048 0 12076 754
rect 12512 0 12540 754
rect 12672 0 12700 754
rect 13136 0 13164 754
rect 13296 0 13324 754
rect 13760 0 13788 754
rect 13920 0 13948 754
rect 14384 0 14412 754
rect 14544 0 14572 754
rect 15008 0 15036 754
rect 15168 0 15196 754
rect 15632 0 15660 754
rect 15792 0 15820 754
rect 16256 0 16284 754
rect 16416 0 16444 754
rect 16880 0 16908 754
rect 17040 0 17068 754
rect 17504 0 17532 754
rect 17664 0 17692 754
rect 18128 0 18156 754
rect 18288 0 18316 754
rect 18752 0 18780 754
rect 18912 0 18940 754
rect 19376 0 19404 754
rect 19536 0 19564 754
rect 20000 0 20028 754
rect 20160 0 20188 754
rect 20624 0 20652 754
rect 20784 0 20812 754
rect 21248 0 21276 754
rect 21408 0 21436 754
rect 21872 0 21900 754
rect 22032 0 22060 754
rect 22496 0 22524 754
rect 22656 0 22684 754
rect 23120 0 23148 754
rect 23280 0 23308 754
rect 23744 0 23772 754
rect 23904 0 23932 754
rect 24368 0 24396 754
rect 24528 0 24556 754
rect 24992 0 25020 754
rect 25152 0 25180 754
rect 25616 0 25644 754
rect 25776 0 25804 754
rect 26240 0 26268 754
rect 26400 0 26428 754
rect 26864 0 26892 754
rect 27024 0 27052 754
rect 27488 0 27516 754
rect 27648 0 27676 754
rect 28112 0 28140 754
rect 28272 0 28300 754
rect 28736 0 28764 754
rect 28896 0 28924 754
rect 29360 0 29388 754
rect 29520 0 29548 754
rect 29984 0 30012 754
rect 30144 0 30172 754
rect 30608 0 30636 754
rect 30768 0 30796 754
rect 31232 0 31260 754
rect 31392 0 31420 754
rect 31856 0 31884 754
rect 32016 0 32044 754
rect 32480 0 32508 754
rect 32640 0 32668 754
rect 33104 0 33132 754
rect 33264 0 33292 754
rect 33728 0 33756 754
rect 33888 0 33916 754
rect 34352 0 34380 754
rect 34512 0 34540 754
rect 34976 0 35004 754
rect 35136 0 35164 754
rect 35600 0 35628 754
rect 35760 0 35788 754
rect 36224 0 36252 754
rect 36384 0 36412 754
rect 36848 0 36876 754
rect 37008 0 37036 754
rect 37472 0 37500 754
rect 37632 0 37660 754
rect 38096 0 38124 754
rect 38256 0 38284 754
rect 38720 0 38748 754
rect 38880 0 38908 754
rect 39344 0 39372 754
rect 39504 0 39532 754
rect 39968 0 39996 754
rect 40128 0 40156 754
rect 40592 0 40620 754
rect 40752 0 40780 754
rect 41216 0 41244 754
rect 41376 0 41404 754
rect 41840 0 41868 754
rect 42000 0 42028 754
rect 42464 0 42492 754
rect 42624 0 42652 754
rect 43088 0 43116 754
rect 43248 0 43276 754
rect 43712 0 43740 754
rect 43872 0 43900 754
rect 44336 0 44364 754
rect 44496 0 44524 754
rect 44960 0 44988 754
rect 45120 0 45148 754
rect 45584 0 45612 754
rect 45744 0 45772 754
rect 46208 0 46236 754
rect 46368 0 46396 754
rect 46832 0 46860 754
rect 46992 0 47020 754
rect 47456 0 47484 754
rect 47616 0 47644 754
rect 48080 0 48108 754
rect 48240 0 48268 754
rect 48704 0 48732 754
rect 48864 0 48892 754
rect 49328 0 49356 754
rect 49488 0 49516 754
rect 49952 0 49980 754
rect 50112 0 50140 754
rect 50576 0 50604 754
rect 50736 0 50764 754
rect 51200 0 51228 754
rect 51360 0 51388 754
rect 51824 0 51852 754
rect 51984 0 52012 754
rect 52448 0 52476 754
rect 52608 0 52636 754
rect 53072 0 53100 754
rect 53232 0 53260 754
rect 53696 0 53724 754
rect 53856 0 53884 754
rect 54320 0 54348 754
rect 54480 0 54508 754
rect 54944 0 54972 754
rect 55104 0 55132 754
rect 55568 0 55596 754
rect 55728 0 55756 754
rect 56192 0 56220 754
rect 56352 0 56380 754
rect 56816 0 56844 754
rect 56976 0 57004 754
rect 57440 0 57468 754
rect 57600 0 57628 754
rect 58064 0 58092 754
rect 58224 0 58252 754
rect 58688 0 58716 754
rect 58848 0 58876 754
rect 59312 0 59340 754
rect 59472 0 59500 754
rect 59936 0 59964 754
rect 60096 0 60124 754
rect 60560 0 60588 754
rect 60720 0 60748 754
rect 61184 0 61212 754
rect 61344 0 61372 754
rect 61808 0 61836 754
rect 61968 0 61996 754
rect 62432 0 62460 754
rect 62592 0 62620 754
rect 63056 0 63084 754
rect 63216 0 63244 754
rect 63680 0 63708 754
rect 63840 0 63868 754
rect 64304 0 64332 754
rect 64464 0 64492 754
rect 64928 0 64956 754
rect 65088 0 65116 754
rect 65552 0 65580 754
rect 65712 0 65740 754
rect 66176 0 66204 754
rect 66336 0 66364 754
rect 66800 0 66828 754
rect 66960 0 66988 754
rect 67424 0 67452 754
rect 67584 0 67612 754
rect 68048 0 68076 754
rect 68208 0 68236 754
rect 68672 0 68700 754
rect 68832 0 68860 754
rect 69296 0 69324 754
rect 69456 0 69484 754
rect 69920 0 69948 754
rect 70080 0 70108 754
rect 70544 0 70572 754
rect 70704 0 70732 754
rect 71168 0 71196 754
rect 71328 0 71356 754
rect 71792 0 71820 754
rect 71952 0 71980 754
rect 72416 0 72444 754
rect 72576 0 72604 754
rect 73040 0 73068 754
rect 73200 0 73228 754
rect 73664 0 73692 754
rect 73824 0 73852 754
rect 74288 0 74316 754
rect 74448 0 74476 754
rect 74912 0 74940 754
rect 75072 0 75100 754
rect 75536 0 75564 754
rect 75696 0 75724 754
rect 76160 0 76188 754
rect 76320 0 76348 754
rect 76784 0 76812 754
rect 76944 0 76972 754
rect 77408 0 77436 754
rect 77568 0 77596 754
rect 78032 0 78060 754
rect 78192 0 78220 754
rect 78656 0 78684 754
rect 78816 0 78844 754
rect 79280 0 79308 754
rect 79440 0 79468 754
rect 79904 0 79932 754
rect 80064 0 80092 754
rect 80528 0 80556 754
rect 80688 0 80716 754
rect 81152 0 81180 754
<< metal3 >>
rect 1132 595 1230 693
rect 1518 595 1616 693
rect 2380 595 2478 693
rect 2766 595 2864 693
rect 3628 595 3726 693
rect 4014 595 4112 693
rect 4876 595 4974 693
rect 5262 595 5360 693
rect 6124 595 6222 693
rect 6510 595 6608 693
rect 7372 595 7470 693
rect 7758 595 7856 693
rect 8620 595 8718 693
rect 9006 595 9104 693
rect 9868 595 9966 693
rect 10254 595 10352 693
rect 11116 595 11214 693
rect 11502 595 11600 693
rect 12364 595 12462 693
rect 12750 595 12848 693
rect 13612 595 13710 693
rect 13998 595 14096 693
rect 14860 595 14958 693
rect 15246 595 15344 693
rect 16108 595 16206 693
rect 16494 595 16592 693
rect 17356 595 17454 693
rect 17742 595 17840 693
rect 18604 595 18702 693
rect 18990 595 19088 693
rect 19852 595 19950 693
rect 20238 595 20336 693
rect 21100 595 21198 693
rect 21486 595 21584 693
rect 22348 595 22446 693
rect 22734 595 22832 693
rect 23596 595 23694 693
rect 23982 595 24080 693
rect 24844 595 24942 693
rect 25230 595 25328 693
rect 26092 595 26190 693
rect 26478 595 26576 693
rect 27340 595 27438 693
rect 27726 595 27824 693
rect 28588 595 28686 693
rect 28974 595 29072 693
rect 29836 595 29934 693
rect 30222 595 30320 693
rect 31084 595 31182 693
rect 31470 595 31568 693
rect 32332 595 32430 693
rect 32718 595 32816 693
rect 33580 595 33678 693
rect 33966 595 34064 693
rect 34828 595 34926 693
rect 35214 595 35312 693
rect 36076 595 36174 693
rect 36462 595 36560 693
rect 37324 595 37422 693
rect 37710 595 37808 693
rect 38572 595 38670 693
rect 38958 595 39056 693
rect 39820 595 39918 693
rect 40206 595 40304 693
rect 41068 595 41166 693
rect 41454 595 41552 693
rect 42316 595 42414 693
rect 42702 595 42800 693
rect 43564 595 43662 693
rect 43950 595 44048 693
rect 44812 595 44910 693
rect 45198 595 45296 693
rect 46060 595 46158 693
rect 46446 595 46544 693
rect 47308 595 47406 693
rect 47694 595 47792 693
rect 48556 595 48654 693
rect 48942 595 49040 693
rect 49804 595 49902 693
rect 50190 595 50288 693
rect 51052 595 51150 693
rect 51438 595 51536 693
rect 52300 595 52398 693
rect 52686 595 52784 693
rect 53548 595 53646 693
rect 53934 595 54032 693
rect 54796 595 54894 693
rect 55182 595 55280 693
rect 56044 595 56142 693
rect 56430 595 56528 693
rect 57292 595 57390 693
rect 57678 595 57776 693
rect 58540 595 58638 693
rect 58926 595 59024 693
rect 59788 595 59886 693
rect 60174 595 60272 693
rect 61036 595 61134 693
rect 61422 595 61520 693
rect 62284 595 62382 693
rect 62670 595 62768 693
rect 63532 595 63630 693
rect 63918 595 64016 693
rect 64780 595 64878 693
rect 65166 595 65264 693
rect 66028 595 66126 693
rect 66414 595 66512 693
rect 67276 595 67374 693
rect 67662 595 67760 693
rect 68524 595 68622 693
rect 68910 595 69008 693
rect 69772 595 69870 693
rect 70158 595 70256 693
rect 71020 595 71118 693
rect 71406 595 71504 693
rect 72268 595 72366 693
rect 72654 595 72752 693
rect 73516 595 73614 693
rect 73902 595 74000 693
rect 74764 595 74862 693
rect 75150 595 75248 693
rect 76012 595 76110 693
rect 76398 595 76496 693
rect 77260 595 77358 693
rect 77646 595 77744 693
rect 78508 595 78606 693
rect 78894 595 78992 693
rect 79756 595 79854 693
rect 80142 595 80240 693
rect 81004 595 81102 693
rect 0 -5 81246 55
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_128
timestamp 1626065694
transform -1 0 41310 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_127
timestamp 1626065694
transform -1 0 61278 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_126
timestamp 1626065694
transform 1 0 61278 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_125
timestamp 1626065694
transform -1 0 62526 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_124
timestamp 1626065694
transform 1 0 62526 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_123
timestamp 1626065694
transform -1 0 63774 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_122
timestamp 1626065694
transform 1 0 63774 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_121
timestamp 1626065694
transform -1 0 65022 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_120
timestamp 1626065694
transform 1 0 65022 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_119
timestamp 1626065694
transform -1 0 66270 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_118
timestamp 1626065694
transform 1 0 66270 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_117
timestamp 1626065694
transform -1 0 67518 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_116
timestamp 1626065694
transform 1 0 67518 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_115
timestamp 1626065694
transform -1 0 68766 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_114
timestamp 1626065694
transform 1 0 68766 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_113
timestamp 1626065694
transform -1 0 70014 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_112
timestamp 1626065694
transform 1 0 70014 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_111
timestamp 1626065694
transform -1 0 71262 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_110
timestamp 1626065694
transform 1 0 71262 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_109
timestamp 1626065694
transform -1 0 72510 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_108
timestamp 1626065694
transform 1 0 72510 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_107
timestamp 1626065694
transform -1 0 73758 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_106
timestamp 1626065694
transform 1 0 73758 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_105
timestamp 1626065694
transform -1 0 75006 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_104
timestamp 1626065694
transform 1 0 75006 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_103
timestamp 1626065694
transform -1 0 76254 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_102
timestamp 1626065694
transform 1 0 76254 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_101
timestamp 1626065694
transform -1 0 77502 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_100
timestamp 1626065694
transform 1 0 77502 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_99
timestamp 1626065694
transform -1 0 78750 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_98
timestamp 1626065694
transform 1 0 78750 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_97
timestamp 1626065694
transform -1 0 79998 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_96
timestamp 1626065694
transform 1 0 79998 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_95
timestamp 1626065694
transform -1 0 81246 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_94
timestamp 1626065694
transform 1 0 43806 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_93
timestamp 1626065694
transform -1 0 45054 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_92
timestamp 1626065694
transform 1 0 45054 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_91
timestamp 1626065694
transform -1 0 46302 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_90
timestamp 1626065694
transform 1 0 46302 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_89
timestamp 1626065694
transform -1 0 47550 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_88
timestamp 1626065694
transform 1 0 47550 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_87
timestamp 1626065694
transform -1 0 48798 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_86
timestamp 1626065694
transform 1 0 48798 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_85
timestamp 1626065694
transform -1 0 50046 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_84
timestamp 1626065694
transform 1 0 50046 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_83
timestamp 1626065694
transform -1 0 51294 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_82
timestamp 1626065694
transform 1 0 51294 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_81
timestamp 1626065694
transform -1 0 52542 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_80
timestamp 1626065694
transform 1 0 52542 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_79
timestamp 1626065694
transform -1 0 53790 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_78
timestamp 1626065694
transform 1 0 53790 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_77
timestamp 1626065694
transform -1 0 55038 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_76
timestamp 1626065694
transform 1 0 55038 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_75
timestamp 1626065694
transform -1 0 56286 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_74
timestamp 1626065694
transform 1 0 56286 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_73
timestamp 1626065694
transform -1 0 57534 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_72
timestamp 1626065694
transform 1 0 57534 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_71
timestamp 1626065694
transform -1 0 58782 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_70
timestamp 1626065694
transform 1 0 58782 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_69
timestamp 1626065694
transform -1 0 60030 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_68
timestamp 1626065694
transform 1 0 60030 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_67
timestamp 1626065694
transform -1 0 42558 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_66
timestamp 1626065694
transform 1 0 42558 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_65
timestamp 1626065694
transform -1 0 43806 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_64
timestamp 1626065694
transform 1 0 41310 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_63
timestamp 1626065694
transform -1 0 21342 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_62
timestamp 1626065694
transform 1 0 21342 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_61
timestamp 1626065694
transform -1 0 22590 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_60
timestamp 1626065694
transform 1 0 22590 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_59
timestamp 1626065694
transform -1 0 23838 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_58
timestamp 1626065694
transform 1 0 23838 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_57
timestamp 1626065694
transform -1 0 25086 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_56
timestamp 1626065694
transform 1 0 25086 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_55
timestamp 1626065694
transform -1 0 26334 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_54
timestamp 1626065694
transform 1 0 26334 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_53
timestamp 1626065694
transform -1 0 27582 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_52
timestamp 1626065694
transform 1 0 27582 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_51
timestamp 1626065694
transform -1 0 28830 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_50
timestamp 1626065694
transform 1 0 28830 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_49
timestamp 1626065694
transform -1 0 30078 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_48
timestamp 1626065694
transform 1 0 30078 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_47
timestamp 1626065694
transform -1 0 31326 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_46
timestamp 1626065694
transform 1 0 31326 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_45
timestamp 1626065694
transform -1 0 32574 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_44
timestamp 1626065694
transform 1 0 32574 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_43
timestamp 1626065694
transform -1 0 33822 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_42
timestamp 1626065694
transform 1 0 33822 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_41
timestamp 1626065694
transform -1 0 35070 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_40
timestamp 1626065694
transform 1 0 35070 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_39
timestamp 1626065694
transform -1 0 36318 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_38
timestamp 1626065694
transform 1 0 36318 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_37
timestamp 1626065694
transform -1 0 37566 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_36
timestamp 1626065694
transform 1 0 37566 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_35
timestamp 1626065694
transform -1 0 38814 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_34
timestamp 1626065694
transform 1 0 38814 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_33
timestamp 1626065694
transform -1 0 40062 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_32
timestamp 1626065694
transform 1 0 40062 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_31
timestamp 1626065694
transform -1 0 2622 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_30
timestamp 1626065694
transform 1 0 2622 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_29
timestamp 1626065694
transform -1 0 3870 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_28
timestamp 1626065694
transform 1 0 3870 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_27
timestamp 1626065694
transform -1 0 5118 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_26
timestamp 1626065694
transform 1 0 5118 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_25
timestamp 1626065694
transform -1 0 6366 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_24
timestamp 1626065694
transform 1 0 6366 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_23
timestamp 1626065694
transform -1 0 7614 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_22
timestamp 1626065694
transform 1 0 7614 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_21
timestamp 1626065694
transform -1 0 8862 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_20
timestamp 1626065694
transform 1 0 8862 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_19
timestamp 1626065694
transform -1 0 10110 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_18
timestamp 1626065694
transform 1 0 10110 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_17
timestamp 1626065694
transform -1 0 11358 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_16
timestamp 1626065694
transform 1 0 11358 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_15
timestamp 1626065694
transform -1 0 12606 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_14
timestamp 1626065694
transform 1 0 12606 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_13
timestamp 1626065694
transform -1 0 13854 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_12
timestamp 1626065694
transform 1 0 13854 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_11
timestamp 1626065694
transform -1 0 15102 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_10
timestamp 1626065694
transform 1 0 15102 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_9
timestamp 1626065694
transform -1 0 16350 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_8
timestamp 1626065694
transform 1 0 16350 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_7
timestamp 1626065694
transform -1 0 17598 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_6
timestamp 1626065694
transform 1 0 17598 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_5
timestamp 1626065694
transform -1 0 18846 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_4
timestamp 1626065694
transform 1 0 18846 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_3
timestamp 1626065694
transform -1 0 20094 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_2
timestamp 1626065694
transform 1 0 20094 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_1
timestamp 1626065694
transform 1 0 1374 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0  sky130_sram_2kbyte_1rw1r_32x512_8_precharge_0_0
timestamp 1626065694
transform -1 0 1374 0 1 0
box 0 -8 624 768
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1626065694
transform 1 0 1029 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1626065694
transform 1 0 1653 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_2
timestamp 1626065694
transform 1 0 20373 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_3
timestamp 1626065694
transform 1 0 19749 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_4
timestamp 1626065694
transform 1 0 19125 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_5
timestamp 1626065694
transform 1 0 18501 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_6
timestamp 1626065694
transform 1 0 17877 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_7
timestamp 1626065694
transform 1 0 17253 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_8
timestamp 1626065694
transform 1 0 16629 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_9
timestamp 1626065694
transform 1 0 16005 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_10
timestamp 1626065694
transform 1 0 15381 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_11
timestamp 1626065694
transform 1 0 14757 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_12
timestamp 1626065694
transform 1 0 14133 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_13
timestamp 1626065694
transform 1 0 13509 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_14
timestamp 1626065694
transform 1 0 12885 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_15
timestamp 1626065694
transform 1 0 12261 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_16
timestamp 1626065694
transform 1 0 11637 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_17
timestamp 1626065694
transform 1 0 11013 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_18
timestamp 1626065694
transform 1 0 10389 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_19
timestamp 1626065694
transform 1 0 9765 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_20
timestamp 1626065694
transform 1 0 9141 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_21
timestamp 1626065694
transform 1 0 8517 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_22
timestamp 1626065694
transform 1 0 7893 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_23
timestamp 1626065694
transform 1 0 7269 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_24
timestamp 1626065694
transform 1 0 6645 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_25
timestamp 1626065694
transform 1 0 6021 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_26
timestamp 1626065694
transform 1 0 5397 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_27
timestamp 1626065694
transform 1 0 4773 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_28
timestamp 1626065694
transform 1 0 4149 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_29
timestamp 1626065694
transform 1 0 3525 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_30
timestamp 1626065694
transform 1 0 2901 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_31
timestamp 1626065694
transform 1 0 2277 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_32
timestamp 1626065694
transform 1 0 20997 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_33
timestamp 1626065694
transform 1 0 40341 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_34
timestamp 1626065694
transform 1 0 39717 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_35
timestamp 1626065694
transform 1 0 39093 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_36
timestamp 1626065694
transform 1 0 38469 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_37
timestamp 1626065694
transform 1 0 37845 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_38
timestamp 1626065694
transform 1 0 37221 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_39
timestamp 1626065694
transform 1 0 36597 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_40
timestamp 1626065694
transform 1 0 35973 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_41
timestamp 1626065694
transform 1 0 35349 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_42
timestamp 1626065694
transform 1 0 34725 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_43
timestamp 1626065694
transform 1 0 34101 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_44
timestamp 1626065694
transform 1 0 33477 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_45
timestamp 1626065694
transform 1 0 32853 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_46
timestamp 1626065694
transform 1 0 32229 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_47
timestamp 1626065694
transform 1 0 31605 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_48
timestamp 1626065694
transform 1 0 30981 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_49
timestamp 1626065694
transform 1 0 30357 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_50
timestamp 1626065694
transform 1 0 29733 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_51
timestamp 1626065694
transform 1 0 29109 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_52
timestamp 1626065694
transform 1 0 28485 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_53
timestamp 1626065694
transform 1 0 27861 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_54
timestamp 1626065694
transform 1 0 27237 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_55
timestamp 1626065694
transform 1 0 26613 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_56
timestamp 1626065694
transform 1 0 25989 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_57
timestamp 1626065694
transform 1 0 25365 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_58
timestamp 1626065694
transform 1 0 24741 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_59
timestamp 1626065694
transform 1 0 24117 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_60
timestamp 1626065694
transform 1 0 23493 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_61
timestamp 1626065694
transform 1 0 22869 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_62
timestamp 1626065694
transform 1 0 22245 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_63
timestamp 1626065694
transform 1 0 21621 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_64
timestamp 1626065694
transform 1 0 41589 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_65
timestamp 1626065694
transform 1 0 60933 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_66
timestamp 1626065694
transform 1 0 60309 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_67
timestamp 1626065694
transform 1 0 59685 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_68
timestamp 1626065694
transform 1 0 59061 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_69
timestamp 1626065694
transform 1 0 58437 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_70
timestamp 1626065694
transform 1 0 57813 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_71
timestamp 1626065694
transform 1 0 57189 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_72
timestamp 1626065694
transform 1 0 56565 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_73
timestamp 1626065694
transform 1 0 55941 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_74
timestamp 1626065694
transform 1 0 55317 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_75
timestamp 1626065694
transform 1 0 54693 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_76
timestamp 1626065694
transform 1 0 54069 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_77
timestamp 1626065694
transform 1 0 53445 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_78
timestamp 1626065694
transform 1 0 52821 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_79
timestamp 1626065694
transform 1 0 52197 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_80
timestamp 1626065694
transform 1 0 51573 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_81
timestamp 1626065694
transform 1 0 50949 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_82
timestamp 1626065694
transform 1 0 50325 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_83
timestamp 1626065694
transform 1 0 49701 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_84
timestamp 1626065694
transform 1 0 49077 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_85
timestamp 1626065694
transform 1 0 48453 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_86
timestamp 1626065694
transform 1 0 47829 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_87
timestamp 1626065694
transform 1 0 47205 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_88
timestamp 1626065694
transform 1 0 46581 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_89
timestamp 1626065694
transform 1 0 45957 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_90
timestamp 1626065694
transform 1 0 45333 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_91
timestamp 1626065694
transform 1 0 44709 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_92
timestamp 1626065694
transform 1 0 44085 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_93
timestamp 1626065694
transform 1 0 43461 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_94
timestamp 1626065694
transform 1 0 42837 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_95
timestamp 1626065694
transform 1 0 42213 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_96
timestamp 1626065694
transform 1 0 80901 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_97
timestamp 1626065694
transform 1 0 80277 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_98
timestamp 1626065694
transform 1 0 79653 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_99
timestamp 1626065694
transform 1 0 79029 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_100
timestamp 1626065694
transform 1 0 78405 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_101
timestamp 1626065694
transform 1 0 77781 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_102
timestamp 1626065694
transform 1 0 77157 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_103
timestamp 1626065694
transform 1 0 76533 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_104
timestamp 1626065694
transform 1 0 75909 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_105
timestamp 1626065694
transform 1 0 75285 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_106
timestamp 1626065694
transform 1 0 74661 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_107
timestamp 1626065694
transform 1 0 74037 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_108
timestamp 1626065694
transform 1 0 73413 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_109
timestamp 1626065694
transform 1 0 72789 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_110
timestamp 1626065694
transform 1 0 72165 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_111
timestamp 1626065694
transform 1 0 71541 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_112
timestamp 1626065694
transform 1 0 70917 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_113
timestamp 1626065694
transform 1 0 70293 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_114
timestamp 1626065694
transform 1 0 69669 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_115
timestamp 1626065694
transform 1 0 69045 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_116
timestamp 1626065694
transform 1 0 68421 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_117
timestamp 1626065694
transform 1 0 67797 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_118
timestamp 1626065694
transform 1 0 67173 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_119
timestamp 1626065694
transform 1 0 66549 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_120
timestamp 1626065694
transform 1 0 65925 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_121
timestamp 1626065694
transform 1 0 65301 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_122
timestamp 1626065694
transform 1 0 64677 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_123
timestamp 1626065694
transform 1 0 64053 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_124
timestamp 1626065694
transform 1 0 63429 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_125
timestamp 1626065694
transform 1 0 62805 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_126
timestamp 1626065694
transform 1 0 62181 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_127
timestamp 1626065694
transform 1 0 61557 0 1 -12
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_128
timestamp 1626065694
transform 1 0 40965 0 1 -12
box 0 0 66 74
<< labels >>
rlabel metal3 s 48556 595 48654 693 4 vdd
rlabel metal3 s 66028 595 66126 693 4 vdd
rlabel metal3 s 81004 595 81102 693 4 vdd
rlabel metal3 s 45198 595 45296 693 4 vdd
rlabel metal3 s 46060 595 46158 693 4 vdd
rlabel metal3 s 71020 595 71118 693 4 vdd
rlabel metal3 s 43564 595 43662 693 4 vdd
rlabel metal3 s 62670 595 62768 693 4 vdd
rlabel metal3 s 66414 595 66512 693 4 vdd
rlabel metal3 s 55182 595 55280 693 4 vdd
rlabel metal3 s 75150 595 75248 693 4 vdd
rlabel metal3 s 48942 595 49040 693 4 vdd
rlabel metal3 s 63918 595 64016 693 4 vdd
rlabel metal3 s 69772 595 69870 693 4 vdd
rlabel metal3 s 78508 595 78606 693 4 vdd
rlabel metal3 s 65166 595 65264 693 4 vdd
rlabel metal3 s 68910 595 69008 693 4 vdd
rlabel metal3 s 46446 595 46544 693 4 vdd
rlabel metal3 s 52300 595 52398 693 4 vdd
rlabel metal3 s 63532 595 63630 693 4 vdd
rlabel metal3 s 49804 595 49902 693 4 vdd
rlabel metal3 s 44812 595 44910 693 4 vdd
rlabel metal3 s 64780 595 64878 693 4 vdd
rlabel metal3 s 77260 595 77358 693 4 vdd
rlabel metal3 s 67662 595 67760 693 4 vdd
rlabel metal3 s 68524 595 68622 693 4 vdd
rlabel metal3 s 42702 595 42800 693 4 vdd
rlabel metal3 s 56430 595 56528 693 4 vdd
rlabel metal3 s 76398 595 76496 693 4 vdd
rlabel metal3 s 71406 595 71504 693 4 vdd
rlabel metal3 s 53934 595 54032 693 4 vdd
rlabel metal3 s 42316 595 42414 693 4 vdd
rlabel metal3 s 77646 595 77744 693 4 vdd
rlabel metal3 s 58540 595 58638 693 4 vdd
rlabel metal3 s 61422 595 61520 693 4 vdd
rlabel metal3 s 54796 595 54894 693 4 vdd
rlabel metal3 s 53548 595 53646 693 4 vdd
rlabel metal3 s 80142 595 80240 693 4 vdd
rlabel metal3 s 41454 595 41552 693 4 vdd
rlabel metal3 s 70158 595 70256 693 4 vdd
rlabel metal3 s 60174 595 60272 693 4 vdd
rlabel metal3 s 57678 595 57776 693 4 vdd
rlabel metal3 s 61036 595 61134 693 4 vdd
rlabel metal3 s 74764 595 74862 693 4 vdd
rlabel metal3 s 73516 595 73614 693 4 vdd
rlabel metal3 s 47308 595 47406 693 4 vdd
rlabel metal3 s 50190 595 50288 693 4 vdd
rlabel metal3 s 51052 595 51150 693 4 vdd
rlabel metal3 s 73902 595 74000 693 4 vdd
rlabel metal3 s 72654 595 72752 693 4 vdd
rlabel metal3 s 43950 595 44048 693 4 vdd
rlabel metal3 s 78894 595 78992 693 4 vdd
rlabel metal3 s 47694 595 47792 693 4 vdd
rlabel metal3 s 57292 595 57390 693 4 vdd
rlabel metal3 s 67276 595 67374 693 4 vdd
rlabel metal3 s 52686 595 52784 693 4 vdd
rlabel metal3 s 58926 595 59024 693 4 vdd
rlabel metal3 s 79756 595 79854 693 4 vdd
rlabel metal3 s 51438 595 51536 693 4 vdd
rlabel metal3 s 62284 595 62382 693 4 vdd
rlabel metal3 s 56044 595 56142 693 4 vdd
rlabel metal3 s 59788 595 59886 693 4 vdd
rlabel metal3 s 72268 595 72366 693 4 vdd
rlabel metal3 s 76012 595 76110 693 4 vdd
rlabel metal3 s 23596 595 23694 693 4 vdd
rlabel metal3 s 23982 595 24080 693 4 vdd
rlabel metal3 s 1132 595 1230 693 4 vdd
rlabel metal3 s 28974 595 29072 693 4 vdd
rlabel metal3 s 31470 595 31568 693 4 vdd
rlabel metal3 s 38572 595 38670 693 4 vdd
rlabel metal3 s 16494 595 16592 693 4 vdd
rlabel metal3 s 2380 595 2478 693 4 vdd
rlabel metal3 s 9006 595 9104 693 4 vdd
rlabel metal3 s 21486 595 21584 693 4 vdd
rlabel metal3 s 38958 595 39056 693 4 vdd
rlabel metal3 s 12750 595 12848 693 4 vdd
rlabel metal3 s 17742 595 17840 693 4 vdd
rlabel metal3 s 26478 595 26576 693 4 vdd
rlabel metal3 s 21100 595 21198 693 4 vdd
rlabel metal3 s 27726 595 27824 693 4 vdd
rlabel metal3 s 19852 595 19950 693 4 vdd
rlabel metal3 s 26092 595 26190 693 4 vdd
rlabel metal3 s 2766 595 2864 693 4 vdd
rlabel metal3 s 33580 595 33678 693 4 vdd
rlabel metal3 s 10254 595 10352 693 4 vdd
rlabel metal3 s 4014 595 4112 693 4 vdd
rlabel metal3 s 6124 595 6222 693 4 vdd
rlabel metal3 s 17356 595 17454 693 4 vdd
rlabel metal3 s 18604 595 18702 693 4 vdd
rlabel metal3 s 12364 595 12462 693 4 vdd
rlabel metal3 s 36462 595 36560 693 4 vdd
rlabel metal3 s 13612 595 13710 693 4 vdd
rlabel metal3 s 15246 595 15344 693 4 vdd
rlabel metal3 s 28588 595 28686 693 4 vdd
rlabel metal3 s 27340 595 27438 693 4 vdd
rlabel metal3 s 35214 595 35312 693 4 vdd
rlabel metal3 s 9868 595 9966 693 4 vdd
rlabel metal3 s 14860 595 14958 693 4 vdd
rlabel metal3 s 39820 595 39918 693 4 vdd
rlabel metal3 s 5262 595 5360 693 4 vdd
rlabel metal3 s 7372 595 7470 693 4 vdd
rlabel metal3 s 11502 595 11600 693 4 vdd
rlabel metal3 s 18990 595 19088 693 4 vdd
rlabel metal3 s 34828 595 34926 693 4 vdd
rlabel metal3 s 8620 595 8718 693 4 vdd
rlabel metal3 s 7758 595 7856 693 4 vdd
rlabel metal3 s 11116 595 11214 693 4 vdd
rlabel metal3 s 22348 595 22446 693 4 vdd
rlabel metal3 s 22734 595 22832 693 4 vdd
rlabel metal3 s 32718 595 32816 693 4 vdd
rlabel metal3 s 25230 595 25328 693 4 vdd
rlabel metal3 s 40206 595 40304 693 4 vdd
rlabel metal3 s 37324 595 37422 693 4 vdd
rlabel metal3 s 41068 595 41166 693 4 vdd
rlabel metal3 s 32332 595 32430 693 4 vdd
rlabel metal3 s 36076 595 36174 693 4 vdd
rlabel metal3 s 4876 595 4974 693 4 vdd
rlabel metal3 s 16108 595 16206 693 4 vdd
rlabel metal3 s 24844 595 24942 693 4 vdd
rlabel metal3 s 37710 595 37808 693 4 vdd
rlabel metal3 s 6510 595 6608 693 4 vdd
rlabel metal3 s 13998 595 14096 693 4 vdd
rlabel metal3 s 1518 595 1616 693 4 vdd
rlabel metal3 s 3628 595 3726 693 4 vdd
rlabel metal3 s 30222 595 30320 693 4 vdd
rlabel metal3 s 29836 595 29934 693 4 vdd
rlabel metal3 s 31084 595 31182 693 4 vdd
rlabel metal3 s 20238 595 20336 693 4 vdd
rlabel metal3 s 33966 595 34064 693 4 vdd
rlabel metal3 s 0 -5 81246 55 4 en_bar
rlabel metal1 s 1280 0 1308 754 4 bl_0
rlabel metal1 s 816 0 844 754 4 br_0
rlabel metal1 s 1440 0 1468 754 4 bl_1
rlabel metal1 s 1904 0 1932 754 4 br_1
rlabel metal1 s 2528 0 2556 754 4 bl_2
rlabel metal1 s 2064 0 2092 754 4 br_2
rlabel metal1 s 2688 0 2716 754 4 bl_3
rlabel metal1 s 3152 0 3180 754 4 br_3
rlabel metal1 s 3776 0 3804 754 4 bl_4
rlabel metal1 s 3312 0 3340 754 4 br_4
rlabel metal1 s 3936 0 3964 754 4 bl_5
rlabel metal1 s 4400 0 4428 754 4 br_5
rlabel metal1 s 5024 0 5052 754 4 bl_6
rlabel metal1 s 4560 0 4588 754 4 br_6
rlabel metal1 s 5184 0 5212 754 4 bl_7
rlabel metal1 s 5648 0 5676 754 4 br_7
rlabel metal1 s 6272 0 6300 754 4 bl_8
rlabel metal1 s 5808 0 5836 754 4 br_8
rlabel metal1 s 6432 0 6460 754 4 bl_9
rlabel metal1 s 6896 0 6924 754 4 br_9
rlabel metal1 s 7520 0 7548 754 4 bl_10
rlabel metal1 s 7056 0 7084 754 4 br_10
rlabel metal1 s 7680 0 7708 754 4 bl_11
rlabel metal1 s 8144 0 8172 754 4 br_11
rlabel metal1 s 8768 0 8796 754 4 bl_12
rlabel metal1 s 8304 0 8332 754 4 br_12
rlabel metal1 s 8928 0 8956 754 4 bl_13
rlabel metal1 s 9392 0 9420 754 4 br_13
rlabel metal1 s 10016 0 10044 754 4 bl_14
rlabel metal1 s 9552 0 9580 754 4 br_14
rlabel metal1 s 10176 0 10204 754 4 bl_15
rlabel metal1 s 10640 0 10668 754 4 br_15
rlabel metal1 s 11264 0 11292 754 4 bl_16
rlabel metal1 s 10800 0 10828 754 4 br_16
rlabel metal1 s 11424 0 11452 754 4 bl_17
rlabel metal1 s 11888 0 11916 754 4 br_17
rlabel metal1 s 12512 0 12540 754 4 bl_18
rlabel metal1 s 12048 0 12076 754 4 br_18
rlabel metal1 s 12672 0 12700 754 4 bl_19
rlabel metal1 s 13136 0 13164 754 4 br_19
rlabel metal1 s 13760 0 13788 754 4 bl_20
rlabel metal1 s 13296 0 13324 754 4 br_20
rlabel metal1 s 13920 0 13948 754 4 bl_21
rlabel metal1 s 14384 0 14412 754 4 br_21
rlabel metal1 s 15008 0 15036 754 4 bl_22
rlabel metal1 s 14544 0 14572 754 4 br_22
rlabel metal1 s 15168 0 15196 754 4 bl_23
rlabel metal1 s 15632 0 15660 754 4 br_23
rlabel metal1 s 16256 0 16284 754 4 bl_24
rlabel metal1 s 15792 0 15820 754 4 br_24
rlabel metal1 s 16416 0 16444 754 4 bl_25
rlabel metal1 s 16880 0 16908 754 4 br_25
rlabel metal1 s 17504 0 17532 754 4 bl_26
rlabel metal1 s 17040 0 17068 754 4 br_26
rlabel metal1 s 17664 0 17692 754 4 bl_27
rlabel metal1 s 18128 0 18156 754 4 br_27
rlabel metal1 s 18752 0 18780 754 4 bl_28
rlabel metal1 s 18288 0 18316 754 4 br_28
rlabel metal1 s 18912 0 18940 754 4 bl_29
rlabel metal1 s 19376 0 19404 754 4 br_29
rlabel metal1 s 20000 0 20028 754 4 bl_30
rlabel metal1 s 19536 0 19564 754 4 br_30
rlabel metal1 s 20160 0 20188 754 4 bl_31
rlabel metal1 s 20624 0 20652 754 4 br_31
rlabel metal1 s 20784 0 20812 754 4 br_32
rlabel metal1 s 21248 0 21276 754 4 bl_32
rlabel metal1 s 21408 0 21436 754 4 bl_33
rlabel metal1 s 21872 0 21900 754 4 br_33
rlabel metal1 s 22496 0 22524 754 4 bl_34
rlabel metal1 s 22032 0 22060 754 4 br_34
rlabel metal1 s 22656 0 22684 754 4 bl_35
rlabel metal1 s 23120 0 23148 754 4 br_35
rlabel metal1 s 23744 0 23772 754 4 bl_36
rlabel metal1 s 23280 0 23308 754 4 br_36
rlabel metal1 s 23904 0 23932 754 4 bl_37
rlabel metal1 s 24368 0 24396 754 4 br_37
rlabel metal1 s 24992 0 25020 754 4 bl_38
rlabel metal1 s 24528 0 24556 754 4 br_38
rlabel metal1 s 25152 0 25180 754 4 bl_39
rlabel metal1 s 25616 0 25644 754 4 br_39
rlabel metal1 s 26240 0 26268 754 4 bl_40
rlabel metal1 s 25776 0 25804 754 4 br_40
rlabel metal1 s 26400 0 26428 754 4 bl_41
rlabel metal1 s 26864 0 26892 754 4 br_41
rlabel metal1 s 27488 0 27516 754 4 bl_42
rlabel metal1 s 27024 0 27052 754 4 br_42
rlabel metal1 s 27648 0 27676 754 4 bl_43
rlabel metal1 s 28112 0 28140 754 4 br_43
rlabel metal1 s 28736 0 28764 754 4 bl_44
rlabel metal1 s 28272 0 28300 754 4 br_44
rlabel metal1 s 28896 0 28924 754 4 bl_45
rlabel metal1 s 29360 0 29388 754 4 br_45
rlabel metal1 s 29984 0 30012 754 4 bl_46
rlabel metal1 s 29520 0 29548 754 4 br_46
rlabel metal1 s 30144 0 30172 754 4 bl_47
rlabel metal1 s 30608 0 30636 754 4 br_47
rlabel metal1 s 31232 0 31260 754 4 bl_48
rlabel metal1 s 30768 0 30796 754 4 br_48
rlabel metal1 s 31392 0 31420 754 4 bl_49
rlabel metal1 s 31856 0 31884 754 4 br_49
rlabel metal1 s 32480 0 32508 754 4 bl_50
rlabel metal1 s 32016 0 32044 754 4 br_50
rlabel metal1 s 32640 0 32668 754 4 bl_51
rlabel metal1 s 33104 0 33132 754 4 br_51
rlabel metal1 s 33728 0 33756 754 4 bl_52
rlabel metal1 s 33264 0 33292 754 4 br_52
rlabel metal1 s 33888 0 33916 754 4 bl_53
rlabel metal1 s 34352 0 34380 754 4 br_53
rlabel metal1 s 34976 0 35004 754 4 bl_54
rlabel metal1 s 34512 0 34540 754 4 br_54
rlabel metal1 s 35136 0 35164 754 4 bl_55
rlabel metal1 s 35600 0 35628 754 4 br_55
rlabel metal1 s 36224 0 36252 754 4 bl_56
rlabel metal1 s 35760 0 35788 754 4 br_56
rlabel metal1 s 36384 0 36412 754 4 bl_57
rlabel metal1 s 36848 0 36876 754 4 br_57
rlabel metal1 s 37472 0 37500 754 4 bl_58
rlabel metal1 s 37008 0 37036 754 4 br_58
rlabel metal1 s 37632 0 37660 754 4 bl_59
rlabel metal1 s 38096 0 38124 754 4 br_59
rlabel metal1 s 38720 0 38748 754 4 bl_60
rlabel metal1 s 38256 0 38284 754 4 br_60
rlabel metal1 s 38880 0 38908 754 4 bl_61
rlabel metal1 s 39344 0 39372 754 4 br_61
rlabel metal1 s 39968 0 39996 754 4 bl_62
rlabel metal1 s 39504 0 39532 754 4 br_62
rlabel metal1 s 40128 0 40156 754 4 bl_63
rlabel metal1 s 40592 0 40620 754 4 br_63
rlabel metal1 s 40752 0 40780 754 4 br_64
rlabel metal1 s 41216 0 41244 754 4 bl_64
rlabel metal1 s 41376 0 41404 754 4 bl_65
rlabel metal1 s 41840 0 41868 754 4 br_65
rlabel metal1 s 42464 0 42492 754 4 bl_66
rlabel metal1 s 42000 0 42028 754 4 br_66
rlabel metal1 s 42624 0 42652 754 4 bl_67
rlabel metal1 s 43088 0 43116 754 4 br_67
rlabel metal1 s 43712 0 43740 754 4 bl_68
rlabel metal1 s 43248 0 43276 754 4 br_68
rlabel metal1 s 43872 0 43900 754 4 bl_69
rlabel metal1 s 44336 0 44364 754 4 br_69
rlabel metal1 s 44960 0 44988 754 4 bl_70
rlabel metal1 s 44496 0 44524 754 4 br_70
rlabel metal1 s 45120 0 45148 754 4 bl_71
rlabel metal1 s 45584 0 45612 754 4 br_71
rlabel metal1 s 46208 0 46236 754 4 bl_72
rlabel metal1 s 45744 0 45772 754 4 br_72
rlabel metal1 s 46368 0 46396 754 4 bl_73
rlabel metal1 s 46832 0 46860 754 4 br_73
rlabel metal1 s 47456 0 47484 754 4 bl_74
rlabel metal1 s 46992 0 47020 754 4 br_74
rlabel metal1 s 47616 0 47644 754 4 bl_75
rlabel metal1 s 48080 0 48108 754 4 br_75
rlabel metal1 s 48704 0 48732 754 4 bl_76
rlabel metal1 s 48240 0 48268 754 4 br_76
rlabel metal1 s 48864 0 48892 754 4 bl_77
rlabel metal1 s 49328 0 49356 754 4 br_77
rlabel metal1 s 49952 0 49980 754 4 bl_78
rlabel metal1 s 49488 0 49516 754 4 br_78
rlabel metal1 s 50112 0 50140 754 4 bl_79
rlabel metal1 s 50576 0 50604 754 4 br_79
rlabel metal1 s 51200 0 51228 754 4 bl_80
rlabel metal1 s 50736 0 50764 754 4 br_80
rlabel metal1 s 51360 0 51388 754 4 bl_81
rlabel metal1 s 51824 0 51852 754 4 br_81
rlabel metal1 s 52448 0 52476 754 4 bl_82
rlabel metal1 s 51984 0 52012 754 4 br_82
rlabel metal1 s 52608 0 52636 754 4 bl_83
rlabel metal1 s 53072 0 53100 754 4 br_83
rlabel metal1 s 53696 0 53724 754 4 bl_84
rlabel metal1 s 53232 0 53260 754 4 br_84
rlabel metal1 s 53856 0 53884 754 4 bl_85
rlabel metal1 s 54320 0 54348 754 4 br_85
rlabel metal1 s 54944 0 54972 754 4 bl_86
rlabel metal1 s 54480 0 54508 754 4 br_86
rlabel metal1 s 55104 0 55132 754 4 bl_87
rlabel metal1 s 55568 0 55596 754 4 br_87
rlabel metal1 s 56192 0 56220 754 4 bl_88
rlabel metal1 s 55728 0 55756 754 4 br_88
rlabel metal1 s 56352 0 56380 754 4 bl_89
rlabel metal1 s 56816 0 56844 754 4 br_89
rlabel metal1 s 57440 0 57468 754 4 bl_90
rlabel metal1 s 56976 0 57004 754 4 br_90
rlabel metal1 s 57600 0 57628 754 4 bl_91
rlabel metal1 s 58064 0 58092 754 4 br_91
rlabel metal1 s 58688 0 58716 754 4 bl_92
rlabel metal1 s 58224 0 58252 754 4 br_92
rlabel metal1 s 58848 0 58876 754 4 bl_93
rlabel metal1 s 59312 0 59340 754 4 br_93
rlabel metal1 s 59936 0 59964 754 4 bl_94
rlabel metal1 s 59472 0 59500 754 4 br_94
rlabel metal1 s 60096 0 60124 754 4 bl_95
rlabel metal1 s 60560 0 60588 754 4 br_95
rlabel metal1 s 60720 0 60748 754 4 br_96
rlabel metal1 s 61184 0 61212 754 4 bl_96
rlabel metal1 s 61344 0 61372 754 4 bl_97
rlabel metal1 s 61808 0 61836 754 4 br_97
rlabel metal1 s 62432 0 62460 754 4 bl_98
rlabel metal1 s 61968 0 61996 754 4 br_98
rlabel metal1 s 62592 0 62620 754 4 bl_99
rlabel metal1 s 63056 0 63084 754 4 br_99
rlabel metal1 s 63680 0 63708 754 4 bl_100
rlabel metal1 s 63216 0 63244 754 4 br_100
rlabel metal1 s 63840 0 63868 754 4 bl_101
rlabel metal1 s 64304 0 64332 754 4 br_101
rlabel metal1 s 64928 0 64956 754 4 bl_102
rlabel metal1 s 64464 0 64492 754 4 br_102
rlabel metal1 s 65088 0 65116 754 4 bl_103
rlabel metal1 s 65552 0 65580 754 4 br_103
rlabel metal1 s 66176 0 66204 754 4 bl_104
rlabel metal1 s 65712 0 65740 754 4 br_104
rlabel metal1 s 66336 0 66364 754 4 bl_105
rlabel metal1 s 66800 0 66828 754 4 br_105
rlabel metal1 s 67424 0 67452 754 4 bl_106
rlabel metal1 s 66960 0 66988 754 4 br_106
rlabel metal1 s 67584 0 67612 754 4 bl_107
rlabel metal1 s 68048 0 68076 754 4 br_107
rlabel metal1 s 68672 0 68700 754 4 bl_108
rlabel metal1 s 68208 0 68236 754 4 br_108
rlabel metal1 s 68832 0 68860 754 4 bl_109
rlabel metal1 s 69296 0 69324 754 4 br_109
rlabel metal1 s 69920 0 69948 754 4 bl_110
rlabel metal1 s 69456 0 69484 754 4 br_110
rlabel metal1 s 70080 0 70108 754 4 bl_111
rlabel metal1 s 70544 0 70572 754 4 br_111
rlabel metal1 s 71168 0 71196 754 4 bl_112
rlabel metal1 s 70704 0 70732 754 4 br_112
rlabel metal1 s 71328 0 71356 754 4 bl_113
rlabel metal1 s 71792 0 71820 754 4 br_113
rlabel metal1 s 72416 0 72444 754 4 bl_114
rlabel metal1 s 71952 0 71980 754 4 br_114
rlabel metal1 s 72576 0 72604 754 4 bl_115
rlabel metal1 s 73040 0 73068 754 4 br_115
rlabel metal1 s 73664 0 73692 754 4 bl_116
rlabel metal1 s 73200 0 73228 754 4 br_116
rlabel metal1 s 73824 0 73852 754 4 bl_117
rlabel metal1 s 74288 0 74316 754 4 br_117
rlabel metal1 s 74912 0 74940 754 4 bl_118
rlabel metal1 s 74448 0 74476 754 4 br_118
rlabel metal1 s 75072 0 75100 754 4 bl_119
rlabel metal1 s 75536 0 75564 754 4 br_119
rlabel metal1 s 76160 0 76188 754 4 bl_120
rlabel metal1 s 75696 0 75724 754 4 br_120
rlabel metal1 s 76320 0 76348 754 4 bl_121
rlabel metal1 s 76784 0 76812 754 4 br_121
rlabel metal1 s 77408 0 77436 754 4 bl_122
rlabel metal1 s 76944 0 76972 754 4 br_122
rlabel metal1 s 77568 0 77596 754 4 bl_123
rlabel metal1 s 78032 0 78060 754 4 br_123
rlabel metal1 s 78656 0 78684 754 4 bl_124
rlabel metal1 s 78192 0 78220 754 4 br_124
rlabel metal1 s 78816 0 78844 754 4 bl_125
rlabel metal1 s 79280 0 79308 754 4 br_125
rlabel metal1 s 79904 0 79932 754 4 bl_126
rlabel metal1 s 79440 0 79468 754 4 br_126
rlabel metal1 s 80064 0 80092 754 4 bl_127
rlabel metal1 s 80528 0 80556 754 4 br_127
rlabel metal1 s 81152 0 81180 754 4 bl_128
rlabel metal1 s 80688 0 80716 754 4 br_128
<< properties >>
string FIXED_BBOX 0 0 81246 754
<< end >>
