* NGSPICE file created from freq_div_flat.ext - technology: sky130A

.subckt freq_div_flat vin vout VDD VSS
X0 VSS a_1515_n911# a_1473_n1179# VSS sky130_fd_pr__nfet_01v8 ad=1.78827e+13p pd=1.9096e+08u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X1 a_n1351_n813# a_n2049_n1179# a_n1608_n1067# VSS sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=1.978e+11p ps=1.99e+06u w=360000u l=150000u
X2 a_n1776_n813# a_n2215_n1179# a_n1861_n1179# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=1.626e+11p ps=1.66e+06u w=360000u l=150000u
X3 sky130_fd_sc_hd__dfxbp_1_7/Q a_1515_n911# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4 sky130_fd_sc_hd__inv_4_7/A sky130_fd_sc_hd__inv_1_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.61695e+13p ps=2.4618e+08u w=1e+06u l=150000u
X5 VSS a_n1183_n1999# a_n1225_n2267# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X6 a_n1776_n1723# a_n2049_n1717# a_n1861_n1723# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X7 VDD sky130_fd_sc_hd__dfxbp_1_4/Q a_n2215_n2805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X8 VDD a_1090_n661# a_1017_n635# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X9 a_n1650_n2433# a_n2049_n2805# a_n1776_n2811# VSS sky130_fd_pr__nfet_01v8 ad=1.392e+11p pd=1.53e+06u as=1.242e+11p ps=1.41e+06u w=360000u l=150000u
X10 a_n1351_n1723# a_n2215_n1717# a_n1608_n1749# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=2.19e+11p ps=2.15e+06u w=420000u l=150000u
X11 a_n1681_n813# a_n2215_n1179# a_n1776_n813# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X12 a_922_n635# a_649_n629# a_837_n635# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X13 sky130_fd_sc_hd__inv_1_2/A a_n752_n1723# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X14 VDD a_n1183_n2837# a_n752_n2811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X15 VSS sky130_fd_sc_hd__inv_4_7/A sky130_fd_sc_hd__inv_4_7/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X16 VSS a_1347_n635# a_1515_n661# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X17 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__inv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X18 VSS a_n1183_n1749# a_n1225_n1345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X19 sky130_fd_sc_hd__inv_1_8/A a_1946_n1723# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X20 a_n1650_n91# a_n2049_n91# a_n1776_275# VSS sky130_fd_pr__nfet_01v8 ad=1.392e+11p pd=1.53e+06u as=1.242e+11p ps=1.41e+06u w=360000u l=150000u
X21 VSS a_1347_n813# a_1515_n911# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22 VSS sky130_fd_sc_hd__inv_4_4/A sky130_fd_sc_hd__inv_4_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X23 VSS a_n1183_177# a_n1225_n91# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X24 a_n1861_n635# sky130_fd_sc_hd__inv_4_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X25 a_n2049_n2805# a_n2215_n2805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X26 VDD sky130_fd_sc_hd__inv_4_4/A sky130_fd_sc_hd__inv_4_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X27 VDD a_n1183_n911# a_n752_n857# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X28 a_n1267_n1723# a_n2049_n1717# a_n1351_n1723# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=0p ps=0u w=420000u l=150000u
X29 a_n1608_21# a_n1776_275# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X30 sky130_fd_sc_hd__inv_4_4/A sky130_fd_sc_hd__inv_1_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X31 a_n1650_n2267# a_n2049_n2267# a_n1776_n1901# VSS sky130_fd_pr__nfet_01v8 ad=1.392e+11p pd=1.53e+06u as=1.242e+11p ps=1.41e+06u w=360000u l=150000u
X32 VSS sky130_fd_sc_hd__inv_4_8/A sky130_fd_sc_hd__inv_4_8/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X33 a_n1225_n1345# a_n2215_n1717# a_n1351_n1723# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.368e+11p ps=1.48e+06u w=360000u l=150000u
X34 sky130_fd_sc_hd__inv_4_4/A sky130_fd_sc_hd__inv_1_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X35 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__inv_4_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 a_1090_n2837# a_922_n2811# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X37 a_n1861_n2267# sky130_fd_sc_hd__inv_4_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.626e+11p pd=1.66e+06u as=0p ps=0u w=420000u l=150000u
X38 sky130_fd_sc_hd__inv_4_8/A sky130_fd_sc_hd__inv_1_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X39 VDD a_n1183_177# a_n752_231# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X40 sky130_fd_sc_hd__inv_1_1/A a_n752_n635# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X41 sky130_fd_sc_hd__dfxbp_1_8/Q a_1515_n1749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X42 a_1017_n813# a_483_n1179# a_922_n813# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X43 a_n1608_n1749# a_n1776_n1723# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.978e+11p pd=1.99e+06u as=0p ps=0u w=640000u l=150000u
X44 a_1090_n661# a_922_n635# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X45 VDD a_n1608_21# a_n1681_275# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X46 VSS a_n1183_n1999# a_n752_n1945# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X47 sky130_fd_sc_hd__inv_4_2/Y sky130_fd_sc_hd__inv_4_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X48 VDD a_1515_n1999# a_1946_n1945# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X49 sky130_fd_sc_hd__inv_4_8/Y sky130_fd_sc_hd__inv_4_8/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X50 a_837_n2267# sky130_fd_sc_hd__inv_4_9/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.626e+11p pd=1.66e+06u as=0p ps=0u w=420000u l=150000u
X51 a_n1861_n1723# sky130_fd_sc_hd__inv_4_2/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.626e+11p pd=1.66e+06u as=0p ps=0u w=420000u l=150000u
X52 sky130_fd_sc_hd__dfxbp_1_1/Q a_n1183_n661# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X53 a_n2049_n629# a_n2215_n629# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X54 a_n1225_n257# a_n2215_n629# a_n1351_n635# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=1.368e+11p ps=1.48e+06u w=360000u l=150000u
X55 a_n1225_n1179# a_n2215_n1179# a_n1351_n813# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X56 VDD a_n1351_n1901# a_n1183_n1999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X57 sky130_fd_sc_hd__inv_4_0/Y sky130_fd_sc_hd__inv_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X58 a_922_n2811# a_483_n2805# a_837_n2811# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=1.626e+11p ps=1.66e+06u w=360000u l=150000u
X59 VSS a_1090_n1067# a_1048_n1179# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+11p ps=1.53e+06u w=420000u l=150000u
X60 sky130_fd_sc_hd__inv_1_9/A a_1946_n1945# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X61 VSS a_1515_n2837# a_1946_n2811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X62 a_1090_n2155# a_922_n1901# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.978e+11p pd=1.99e+06u as=0p ps=0u w=640000u l=150000u
X63 VSS a_n1183_n1749# a_n752_n1723# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X64 VSS sky130_fd_sc_hd__dfxbp_1_4/Q a_n2215_n2805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X65 VDD a_1347_n1723# a_1515_n1749# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X66 a_n1776_275# a_n2049_n91# a_n1861_n91# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X67 sky130_fd_sc_hd__inv_1_9/A a_1946_n1945# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X68 VDD sky130_fd_sc_hd__dfxbp_1_9/Q a_483_n1717# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X69 sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__inv_1_1/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X70 a_1048_n2433# a_649_n2805# a_922_n2811# VSS sky130_fd_pr__nfet_01v8 ad=1.392e+11p pd=1.53e+06u as=0p ps=0u w=360000u l=150000u
X71 a_837_n1723# sky130_fd_sc_hd__inv_4_8/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.626e+11p pd=1.66e+06u as=0p ps=0u w=420000u l=150000u
X72 VDD a_1515_n2837# a_1431_n2811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.764e+11p ps=1.68e+06u w=420000u l=150000u
X73 VSS sky130_fd_sc_hd__inv_4_9/A sky130_fd_sc_hd__inv_4_9/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X74 VDD a_1090_n2837# a_1017_n2811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X75 sky130_fd_sc_hd__inv_4_1/Y sky130_fd_sc_hd__inv_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X76 VDD sky130_fd_sc_hd__inv_4_9/A sky130_fd_sc_hd__inv_4_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X77 sky130_fd_sc_hd__dfxbp_1_8/Q a_1515_n1749# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X78 VSS a_1090_n661# a_1048_n257# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+11p ps=1.53e+06u w=420000u l=150000u
X79 a_n1608_n2155# a_n1776_n1901# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X80 a_649_n1179# a_483_n1179# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X81 VDD a_n1183_n1999# a_n752_n1945# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X82 sky130_fd_sc_hd__dfxbp_1_4/Q a_n1183_n1999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X83 VSS sky130_fd_sc_hd__inv_4_3/A sky130_fd_sc_hd__inv_4_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X84 sky130_fd_sc_hd__inv_4_2/Y sky130_fd_sc_hd__inv_4_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X85 a_922_n1901# a_483_n2267# a_837_n2267# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=0p ps=0u w=360000u l=150000u
X86 sky130_fd_sc_hd__dfxbp_1_5/Q a_n1183_n2837# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X87 VDD a_1515_n1999# a_1431_n1901# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.764e+11p ps=1.68e+06u w=420000u l=150000u
X88 sky130_fd_sc_hd__dfxbp_1_7/Q a_1515_n911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X89 VDD a_1090_n2155# a_1017_n1901# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X90 a_1347_n813# a_483_n1179# a_1090_n1067# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=2.19e+11p ps=2.15e+06u w=420000u l=150000u
X91 a_n2049_n2805# a_n2215_n2805# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X92 a_1473_n257# a_483_n629# a_1347_n635# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=1.368e+11p ps=1.48e+06u w=360000u l=150000u
X93 a_1048_n2267# a_649_n2267# a_922_n1901# VSS sky130_fd_pr__nfet_01v8 ad=1.392e+11p pd=1.53e+06u as=0p ps=0u w=360000u l=150000u
X94 VSS sky130_fd_sc_hd__inv_4_8/A sky130_fd_sc_hd__inv_4_8/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X95 sky130_fd_sc_hd__inv_4_3/A sky130_fd_sc_hd__inv_1_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X96 a_n1776_n2811# a_n2215_n2805# a_n1861_n2811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.626e+11p ps=1.66e+06u w=360000u l=150000u
X97 sky130_fd_sc_hd__inv_1_5/A a_n752_n2811# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X98 sky130_fd_sc_hd__inv_4_9/Y sky130_fd_sc_hd__inv_4_9/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X99 a_n1351_n2811# a_n2049_n2805# a_n1608_n2837# VSS sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=1.978e+11p ps=1.99e+06u w=360000u l=150000u
X100 sky130_fd_sc_hd__inv_4_6/Y sky130_fd_sc_hd__inv_4_6/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X101 VDD a_1515_n911# a_1946_n857# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X102 VDD a_1515_n911# a_1431_n813# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.764e+11p ps=1.68e+06u w=420000u l=150000u
X103 sky130_fd_sc_hd__inv_4_0/Y sky130_fd_sc_hd__inv_4_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X104 VSS sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__inv_4_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X105 sky130_fd_sc_hd__inv_4_9/Y sky130_fd_sc_hd__inv_4_9/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X106 VSS a_1347_n1723# a_1515_n1749# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X107 a_837_n635# sky130_fd_sc_hd__inv_4_6/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.626e+11p pd=1.66e+06u as=0p ps=0u w=420000u l=150000u
X108 VSS a_n1183_177# a_n752_231# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X109 a_n2049_n1179# a_n2215_n1179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X110 sky130_fd_sc_hd__inv_4_6/A sky130_fd_sc_hd__inv_1_6/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X111 VSS sky130_fd_sc_hd__dfxbp_1_10/Q a_483_n2267# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X112 sky130_fd_sc_hd__inv_4_8/Y sky130_fd_sc_hd__inv_4_8/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X113 VSS a_1515_n1999# a_1473_n2267# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X114 VDD a_n1351_n813# a_n1183_n911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X115 a_n2049_n629# a_n2215_n629# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X116 VDD sky130_fd_sc_hd__dfxbp_1_10/Q a_483_n2267# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X117 a_n1776_n1901# a_n2215_n2267# a_n1861_n2267# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X118 VDD sky130_fd_sc_hd__inv_4_2/A sky130_fd_sc_hd__inv_4_2/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X119 a_n1351_n1901# a_n2049_n2267# a_n1608_n2155# VSS sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=1.978e+11p ps=1.99e+06u w=360000u l=150000u
X120 a_1473_n1345# a_483_n1717# a_1347_n1723# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=1.368e+11p ps=1.48e+06u w=360000u l=150000u
X121 a_n1650_n257# a_n2049_n629# a_n1776_n635# VSS sky130_fd_pr__nfet_01v8 ad=1.392e+11p pd=1.53e+06u as=1.242e+11p ps=1.41e+06u w=360000u l=150000u
X122 sky130_fd_sc_hd__dfxbp_1_9/Q a_1515_n1999# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X123 a_n1776_n2811# a_n2049_n2805# a_n1861_n2811# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X124 sky130_fd_sc_hd__inv_4_2/A sky130_fd_sc_hd__inv_1_2/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X125 VDD sky130_fd_sc_hd__inv_4_3/A sky130_fd_sc_hd__inv_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X126 a_n1776_n635# a_n2215_n629# a_n1861_n635# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.626e+11p ps=1.66e+06u w=360000u l=150000u
X127 a_n1351_n2811# a_n2215_n2805# a_n1608_n2837# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=2.19e+11p ps=2.15e+06u w=420000u l=150000u
X128 sky130_fd_sc_hd__inv_4_10/A sky130_fd_sc_hd__inv_1_10/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X129 a_n1267_n813# a_n2049_n1179# a_n1351_n813# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X130 sky130_fd_sc_hd__inv_4_6/Y sky130_fd_sc_hd__inv_4_6/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X131 sky130_fd_sc_hd__inv_1_5/A a_n752_n2811# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X132 VSS sky130_fd_sc_hd__dfxbp_1_9/Q a_483_n1717# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X133 sky130_fd_sc_hd__inv_4_1/Y sky130_fd_sc_hd__inv_4_1/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X134 VSS vin a_n2215_n91# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X135 VSS a_1515_n1749# a_1473_n1345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X136 a_n1681_275# a_n2215_n91# a_n1776_275# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X137 VSS sky130_fd_sc_hd__inv_4_9/A sky130_fd_sc_hd__inv_4_9/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X138 a_1017_n1723# a_483_n1717# a_922_n1723# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X139 a_n1861_n1723# sky130_fd_sc_hd__inv_4_2/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X140 sky130_fd_sc_hd__inv_4_5/Y sky130_fd_sc_hd__inv_4_5/A VSS VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X141 a_1090_n2155# a_922_n1901# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X142 sky130_fd_sc_hd__inv_1_6/A a_1946_n635# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X143 a_n1776_n1901# a_n2049_n2267# a_n1861_n2267# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X144 VSS a_n1608_n1067# a_n1650_n1179# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+11p ps=1.53e+06u w=420000u l=150000u
X145 VSS a_n1183_n2837# a_n1225_n2433# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X146 VDD sky130_fd_sc_hd__inv_4_9/A sky130_fd_sc_hd__inv_4_9/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X147 VDD a_1090_n1067# a_1017_n813# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X148 a_922_n813# a_649_n1179# a_837_n1179# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X149 a_n1861_n91# sky130_fd_sc_hd__inv_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.626e+11p pd=1.66e+06u as=0p ps=0u w=420000u l=150000u
X150 a_n1351_n1901# a_n2215_n2267# a_n1608_n2155# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X151 a_1473_n1179# a_483_n1179# a_1347_n813# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.368e+11p ps=1.48e+06u w=360000u l=150000u
X152 VSS a_1347_n1901# a_1515_n1999# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X153 a_n1608_n2837# a_n1776_n2811# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X154 VDD a_n1351_n1723# a_n1183_n1749# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X155 a_n1267_n2811# a_n2049_n2805# a_n1351_n2811# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=0p ps=0u w=420000u l=150000u
X156 a_837_n1723# sky130_fd_sc_hd__inv_4_8/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X157 a_n1608_n661# a_n1776_n635# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X158 VSS sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__inv_4_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X159 a_n1681_n1723# a_n2215_n1717# a_n1776_n1723# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X160 a_649_n1717# a_483_n1717# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X161 VSS a_1515_n661# a_1473_n257# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X162 a_n1225_n2433# a_n2215_n2805# a_n1351_n2811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X163 a_1090_n1749# a_922_n1723# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.978e+11p pd=1.99e+06u as=0p ps=0u w=640000u l=150000u
X164 sky130_fd_sc_hd__inv_4_3/Y sky130_fd_sc_hd__inv_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X165 sky130_fd_sc_hd__inv_4_9/Y sky130_fd_sc_hd__inv_4_9/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X166 sky130_fd_sc_hd__inv_1_8/A a_1946_n1723# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X167 VSS sky130_fd_sc_hd__inv_4_2/A sky130_fd_sc_hd__inv_4_2/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X168 a_n1861_n1179# sky130_fd_sc_hd__inv_4_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X169 sky130_fd_sc_hd__inv_4_10/A sky130_fd_sc_hd__inv_1_10/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X170 sky130_fd_sc_hd__inv_4_9/Y sky130_fd_sc_hd__inv_4_9/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X171 sky130_fd_sc_hd__inv_1_7/A a_1946_n857# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X172 a_n1267_n1901# a_n2049_n2267# a_n1351_n1901# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=0p ps=0u w=420000u l=150000u
X173 sky130_fd_sc_hd__dfxbp_1_10/Q a_1515_n2837# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X174 VDD sky130_fd_sc_hd__inv_4_8/A sky130_fd_sc_hd__inv_4_8/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X175 VSS a_n1351_n2811# a_n1183_n2837# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X176 sky130_fd_sc_hd__inv_4_5/Y sky130_fd_sc_hd__inv_4_5/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X177 sky130_fd_sc_hd__dfxbp_1_2/Q a_n1183_n1749# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X178 sky130_fd_sc_hd__inv_4_5/Y sky130_fd_sc_hd__inv_4_5/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X179 a_n1861_n2811# sky130_fd_sc_hd__inv_4_5/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X180 a_1431_n1723# a_649_n1717# a_1347_n1723# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X181 VDD sky130_fd_sc_hd__inv_4_3/A sky130_fd_sc_hd__inv_4_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X182 a_n1225_n2267# a_n2215_n2267# a_n1351_n1901# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X183 a_1347_n1723# a_649_n1717# a_1090_n1749# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X184 a_n2049_n91# a_n2215_n91# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X185 VSS a_1090_n2155# a_1048_n2267# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X186 VSS a_1515_n661# a_1946_n635# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X187 a_837_n635# sky130_fd_sc_hd__inv_4_6/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X188 VSS a_n1183_n2837# a_n752_n2811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X189 VDD sky130_fd_sc_hd__dfxbp_1_7/Q a_483_n629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X190 VDD a_1347_n2811# a_1515_n2837# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X191 VDD sky130_fd_sc_hd__dfxbp_1_5/Q a_483_n2805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X192 a_837_n2811# sky130_fd_sc_hd__inv_4_10/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X193 sky130_fd_sc_hd__inv_4_8/Y sky130_fd_sc_hd__inv_4_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X194 VDD a_n1608_n661# a_n1681_n635# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.533e+11p ps=1.57e+06u w=420000u l=150000u
X195 VSS a_1090_n1749# a_1048_n1345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+11p ps=1.53e+06u w=420000u l=150000u
X196 vout a_1515_n661# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X197 VSS a_n1351_n635# a_n1183_n661# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X198 a_1347_n1723# a_483_n1717# a_1090_n1749# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.19e+11p ps=2.15e+06u w=420000u l=150000u
X199 VSS a_n1183_n661# a_n1225_n257# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X200 a_649_n2267# a_483_n2267# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X201 VSS a_n1351_275# a_n1183_177# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X202 a_1347_n813# a_649_n1179# a_1090_n1067# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.978e+11p ps=1.99e+06u w=360000u l=150000u
X203 VDD vin a_n2215_n91# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X204 a_649_n2267# a_483_n2267# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X205 a_n1776_n635# a_n2049_n629# a_n1861_n635# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X206 a_n1608_21# a_n1776_275# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.978e+11p pd=1.99e+06u as=0p ps=0u w=640000u l=150000u
X207 VSS sky130_fd_sc_hd__inv_4_4/A sky130_fd_sc_hd__inv_4_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X208 sky130_fd_sc_hd__inv_4_5/Y sky130_fd_sc_hd__inv_4_5/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X209 a_1431_n635# a_649_n629# a_1347_n635# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X210 VSS sky130_fd_sc_hd__inv_4_5/A sky130_fd_sc_hd__inv_4_5/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X211 sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__inv_1_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X212 VSS a_n1608_21# a_n1650_n91# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X213 VDD sky130_fd_sc_hd__inv_4_4/A sky130_fd_sc_hd__inv_4_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X214 sky130_fd_sc_hd__dfxbp_1_3/Q a_n1183_n911# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X215 sky130_fd_sc_hd__inv_4_5/A sky130_fd_sc_hd__inv_1_5/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X216 VSS sky130_fd_sc_hd__inv_4_6/A sky130_fd_sc_hd__inv_4_6/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X217 a_649_n1717# a_483_n1717# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X218 sky130_fd_sc_hd__inv_1_3/A a_n752_n857# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X219 VDD sky130_fd_sc_hd__inv_4_0/A sky130_fd_sc_hd__inv_4_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X220 VDD a_n1351_n635# a_n1183_n661# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X221 VDD sky130_fd_sc_hd__inv_4_8/A sky130_fd_sc_hd__inv_4_8/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X222 VSS a_1515_n911# a_1946_n857# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X223 sky130_fd_sc_hd__dfxbp_1_0/Q a_n1183_177# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X224 VDD a_n1183_n661# a_n1267_n635# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.764e+11p ps=1.68e+06u w=420000u l=150000u
X225 VDD sky130_fd_sc_hd__dfxbp_1_8/Q a_483_n1179# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X226 VDD sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__inv_4_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X227 VDD sky130_fd_sc_hd__inv_4_7/A sky130_fd_sc_hd__inv_4_7/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X228 VSS sky130_fd_sc_hd__dfxbp_1_1/Q a_n2215_n1179# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X229 VDD sky130_fd_sc_hd__inv_4_5/A sky130_fd_sc_hd__inv_4_5/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X230 a_1473_n2433# a_483_n2805# a_1347_n2811# VSS sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=1.368e+11p ps=1.48e+06u w=360000u l=150000u
X231 sky130_fd_sc_hd__inv_1_0/A a_n752_231# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X232 a_n1776_275# a_n2215_n91# a_n1861_n91# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X233 sky130_fd_sc_hd__inv_1_10/A a_1946_n2811# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X234 VSS sky130_fd_sc_hd__inv_4_6/A sky130_fd_sc_hd__inv_4_6/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X235 sky130_fd_sc_hd__inv_4_5/A sky130_fd_sc_hd__inv_1_5/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X236 a_n1351_n635# a_n2215_n629# a_n1608_n661# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X237 VSS sky130_fd_sc_hd__dfxbp_1_7/Q a_483_n629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X238 a_n2049_n91# a_n2215_n91# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X239 VSS sky130_fd_sc_hd__dfxbp_1_5/Q a_483_n2805# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X240 sky130_fd_sc_hd__inv_4_7/A sky130_fd_sc_hd__inv_1_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X241 VSS a_1515_n2837# a_1473_n2433# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X242 sky130_fd_sc_hd__inv_4_8/Y sky130_fd_sc_hd__inv_4_8/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X243 VDD a_n1608_n1749# a_n1681_n1723# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X244 a_1090_n2837# a_922_n2811# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.978e+11p pd=1.99e+06u as=0p ps=0u w=640000u l=150000u
X245 VSS sky130_fd_sc_hd__inv_4_10/A sky130_fd_sc_hd__inv_4_10/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X246 a_n1351_275# a_n2049_n91# a_n1608_21# VSS sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=0p ps=0u w=360000u l=150000u
X247 a_1017_n2811# a_483_n2805# a_922_n2811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X248 VDD a_n1183_n1749# a_n1267_n1723# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X249 a_n1861_n2811# sky130_fd_sc_hd__inv_4_5/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X250 a_n1608_n1067# a_n1776_n813# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X251 a_n2049_n1179# a_n2215_n1179# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X252 VSS a_n1608_n2155# a_n1650_n2267# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X253 VDD a_1347_n813# a_1515_n911# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X254 sky130_fd_sc_hd__inv_4_3/Y sky130_fd_sc_hd__inv_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X255 a_n1351_n635# a_n2049_n629# a_n1608_n661# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.978e+11p ps=1.99e+06u w=360000u l=150000u
X256 VDD a_n1183_n661# a_n752_n635# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X257 VSS sky130_fd_sc_hd__inv_4_0/A sky130_fd_sc_hd__inv_4_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X258 a_1473_n2267# a_483_n2267# a_1347_n1901# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.368e+11p ps=1.48e+06u w=360000u l=150000u
X259 sky130_fd_sc_hd__inv_4_0/Y sky130_fd_sc_hd__inv_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X260 a_1090_n1067# a_922_n813# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X261 sky130_fd_sc_hd__inv_4_1/Y sky130_fd_sc_hd__inv_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X262 VDD a_n1351_n2811# a_n1183_n2837# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X263 vout a_1515_n661# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X264 VDD sky130_fd_sc_hd__inv_4_7/A sky130_fd_sc_hd__inv_4_7/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X265 a_837_n2811# sky130_fd_sc_hd__inv_4_10/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X266 a_1017_n1901# a_483_n2267# a_922_n1901# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X267 a_n1861_n2267# sky130_fd_sc_hd__inv_4_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X268 a_n1681_n2811# a_n2215_n2805# a_n1776_n2811# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X269 a_649_n2805# a_483_n2805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X270 VSS a_n1608_n1749# a_n1650_n1345# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+11p ps=1.53e+06u w=420000u l=150000u
X271 sky130_fd_sc_hd__inv_1_6/A a_1946_n635# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X272 sky130_fd_sc_hd__inv_4_10/Y sky130_fd_sc_hd__inv_4_10/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X273 sky130_fd_sc_hd__inv_1_10/A a_1946_n2811# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X274 sky130_fd_sc_hd__inv_1_0/A a_n752_231# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X275 a_922_n1723# a_649_n1717# a_837_n1723# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X276 VDD sky130_fd_sc_hd__inv_4_0/A sky130_fd_sc_hd__inv_4_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X277 VDD a_n1183_177# a_n1267_275# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.764e+11p ps=1.68e+06u w=420000u l=150000u
X278 a_837_n2267# sky130_fd_sc_hd__inv_4_9/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X279 a_n1681_n1901# a_n2215_n2267# a_n1776_n1901# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X280 a_n1608_n1749# a_n1776_n1723# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X281 VDD sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__inv_4_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X282 a_n1608_n661# a_n1776_n635# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X283 VDD a_1515_n1749# a_1946_n1723# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X284 sky130_fd_sc_hd__dfxbp_1_2/Q a_n1183_n1749# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X285 VDD sky130_fd_sc_hd__inv_4_10/A sky130_fd_sc_hd__inv_4_10/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X286 sky130_fd_sc_hd__dfxbp_1_5/Q a_n1183_n2837# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X287 sky130_fd_sc_hd__dfxbp_1_3/Q a_n1183_n911# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X288 sky130_fd_sc_hd__inv_4_3/Y sky130_fd_sc_hd__inv_4_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X289 VSS a_n1351_n813# a_n1183_n911# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X290 a_1431_n2811# a_649_n2805# a_1347_n2811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X291 a_n1681_n635# a_n2215_n629# a_n1776_n635# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X292 VDD sky130_fd_sc_hd__inv_4_2/A sky130_fd_sc_hd__inv_4_2/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X293 sky130_fd_sc_hd__inv_1_2/A a_n752_n1723# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X294 VDD a_n1351_275# a_n1183_177# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X295 a_1347_n2811# a_649_n2805# a_1090_n2837# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X296 sky130_fd_sc_hd__dfxbp_1_10/Q a_1515_n2837# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X297 sky130_fd_sc_hd__inv_4_0/Y sky130_fd_sc_hd__inv_4_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X298 a_n1351_275# a_n2215_n91# a_n1608_21# VDD sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X299 VDD sky130_fd_sc_hd__dfxbp_1_0/Q a_n2215_n629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X300 VSS a_n1183_n911# a_n1225_n1179# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X301 VDD sky130_fd_sc_hd__dfxbp_1_3/Q a_n2215_n1717# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X302 a_1347_n635# a_649_n629# a_1090_n661# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.978e+11p ps=1.99e+06u w=360000u l=150000u
X303 sky130_fd_sc_hd__inv_4_10/Y sky130_fd_sc_hd__inv_4_10/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X304 a_1431_n1901# a_649_n2267# a_1347_n1901# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X305 a_n1650_n1345# a_n2049_n1717# a_n1776_n1723# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.242e+11p ps=1.41e+06u w=360000u l=150000u
X306 VSS a_1090_n2837# a_1048_n2433# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X307 VDD a_n1183_n1749# a_n752_n1723# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X308 VSS sky130_fd_sc_hd__inv_4_10/A sky130_fd_sc_hd__inv_4_10/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X309 a_837_n1179# sky130_fd_sc_hd__inv_4_7/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X310 a_1347_n2811# a_483_n2805# a_1090_n2837# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X311 VSS sky130_fd_sc_hd__inv_4_0/A sky130_fd_sc_hd__inv_4_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X312 a_1347_n1901# a_649_n2267# a_1090_n2155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X313 VSS a_1347_n2811# a_1515_n2837# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X314 VDD a_n1608_n1067# a_n1681_n813# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X315 a_649_n629# a_483_n629# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X316 VSS sky130_fd_sc_hd__inv_4_3/A sky130_fd_sc_hd__inv_4_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X317 sky130_fd_sc_hd__dfxbp_1_4/Q a_n1183_n1999# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X318 sky130_fd_sc_hd__inv_4_8/A sky130_fd_sc_hd__inv_1_8/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X319 sky130_fd_sc_hd__inv_1_1/A a_n752_n635# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X320 a_n2049_n1717# a_n2215_n1717# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X321 VDD a_1515_n661# a_1946_n635# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X322 a_1347_n1901# a_483_n2267# a_1090_n2155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X323 a_649_n2805# a_483_n2805# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X324 sky130_fd_sc_hd__inv_4_3/A sky130_fd_sc_hd__inv_1_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X325 a_n1650_n1179# a_n2049_n1179# a_n1776_n813# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X326 a_1090_n661# a_922_n635# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X327 a_n1776_n813# a_n2049_n1179# a_n1861_n1179# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X328 a_1017_n635# a_483_n629# a_922_n635# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X329 sky130_fd_sc_hd__inv_4_10/Y sky130_fd_sc_hd__inv_4_10/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X330 sky130_fd_sc_hd__inv_1_4/A a_n752_n1945# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X331 sky130_fd_sc_hd__inv_4_2/Y sky130_fd_sc_hd__inv_4_2/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X332 a_1431_n813# a_649_n1179# a_1347_n813# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X333 a_1048_n257# a_649_n629# a_922_n635# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.242e+11p ps=1.41e+06u w=360000u l=150000u
X334 a_1090_n1749# a_922_n1723# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X335 sky130_fd_sc_hd__inv_1_4/A a_n752_n1945# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X336 a_n1861_n1179# sky130_fd_sc_hd__inv_4_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X337 a_922_n635# a_483_n629# a_837_n635# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X338 sky130_fd_sc_hd__dfxbp_1_0/Q a_n1183_177# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X339 VDD sky130_fd_sc_hd__inv_4_6/A sky130_fd_sc_hd__inv_4_6/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X340 VDD sky130_fd_sc_hd__inv_4_10/A sky130_fd_sc_hd__inv_4_10/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X341 a_n1267_275# a_n2049_n91# a_n1351_275# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X342 VSS a_1515_n1999# a_1946_n1945# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X343 VSS a_n1183_n911# a_n752_n857# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X344 VSS sky130_fd_sc_hd__dfxbp_1_2/Q a_n2215_n2267# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X345 sky130_fd_sc_hd__inv_1_3/A a_n752_n857# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X346 VDD sky130_fd_sc_hd__dfxbp_1_1/Q a_n2215_n1179# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X347 a_837_n1179# sky130_fd_sc_hd__inv_4_7/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.626e+11p pd=1.66e+06u as=0p ps=0u w=420000u l=150000u
X348 VDD sky130_fd_sc_hd__dfxbp_1_2/Q a_n2215_n2267# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X349 sky130_fd_sc_hd__inv_4_0/A sky130_fd_sc_hd__inv_1_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X350 a_922_n1723# a_483_n1717# a_837_n1723# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=0p ps=0u w=360000u l=150000u
X351 a_1090_n1067# a_922_n813# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X352 sky130_fd_sc_hd__inv_4_1/Y sky130_fd_sc_hd__inv_4_1/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X353 VSS a_1515_n1749# a_1946_n1723# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X354 sky130_fd_sc_hd__inv_1_7/A a_1946_n857# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X355 a_n1225_n91# a_n2215_n91# a_n1351_275# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X356 a_n1608_n1067# a_n1776_n813# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X357 VDD a_n1183_n911# a_n1267_n813# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X358 VSS sky130_fd_sc_hd__dfxbp_1_0/Q a_n2215_n629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X359 a_n1861_n635# sky130_fd_sc_hd__inv_4_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X360 sky130_fd_sc_hd__inv_4_9/A sky130_fd_sc_hd__inv_1_9/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X361 sky130_fd_sc_hd__inv_4_2/Y sky130_fd_sc_hd__inv_4_2/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X362 VSS a_n1351_n1723# a_n1183_n1749# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X363 VSS sky130_fd_sc_hd__dfxbp_1_3/Q a_n2215_n1717# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X364 VDD a_1347_n635# a_1515_n661# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X365 VDD a_n1608_n2837# a_n1681_n2811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X366 sky130_fd_sc_hd__inv_4_10/Y sky130_fd_sc_hd__inv_4_10/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X367 a_1048_n1345# a_649_n1717# a_922_n1723# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X368 VDD a_1515_n1749# a_1431_n1723# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X369 VDD a_n1183_n2837# a_n1267_n2811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X370 sky130_fd_sc_hd__inv_4_9/A sky130_fd_sc_hd__inv_1_9/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X371 VSS sky130_fd_sc_hd__inv_4_7/A sky130_fd_sc_hd__inv_4_7/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X372 a_649_n1179# a_483_n1179# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X373 a_n1608_n2155# a_n1776_n1901# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X374 VDD a_1090_n1749# a_1017_n1723# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X375 a_1347_n635# a_483_n629# a_1090_n661# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X376 a_n2049_n2267# a_n2215_n2267# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X377 a_n1351_n813# a_n2215_n1179# a_n1608_n1067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X378 sky130_fd_sc_hd__dfxbp_1_9/Q a_1515_n1999# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X379 sky130_fd_sc_hd__inv_4_4/Y sky130_fd_sc_hd__inv_4_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X380 VDD sky130_fd_sc_hd__inv_4_6/A sky130_fd_sc_hd__inv_4_6/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X381 a_n2049_n2267# a_n2215_n2267# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X382 VSS sky130_fd_sc_hd__inv_4_5/A sky130_fd_sc_hd__inv_4_5/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X383 VSS a_n1608_n661# a_n1650_n257# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X384 sky130_fd_sc_hd__inv_4_6/Y sky130_fd_sc_hd__inv_4_6/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X385 sky130_fd_sc_hd__inv_4_4/Y sky130_fd_sc_hd__inv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X386 VDD a_n1608_n2155# a_n1681_n1901# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X387 a_922_n813# a_483_n1179# a_837_n1179# VSS sky130_fd_pr__nfet_01v8 ad=1.242e+11p pd=1.41e+06u as=0p ps=0u w=360000u l=150000u
X388 VDD a_1515_n661# a_1431_n635# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X389 a_649_n629# a_483_n629# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X390 VDD a_n1183_n1999# a_n1267_n1901# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X391 sky130_fd_sc_hd__inv_4_3/Y sky130_fd_sc_hd__inv_4_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X392 a_n2049_n1717# a_n2215_n1717# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X393 VSS a_n1608_n2837# a_n1650_n2433# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X394 a_1048_n1179# a_649_n1179# a_922_n813# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X395 a_n1351_n1723# a_n2049_n1717# a_n1608_n1749# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X396 a_n1776_n1723# a_n2215_n1717# a_n1861_n1723# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X397 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__inv_4_7/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X398 VSS a_n1183_n661# a_n752_n635# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X399 sky130_fd_sc_hd__inv_4_0/A sky130_fd_sc_hd__inv_1_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X400 sky130_fd_sc_hd__dfxbp_1_1/Q a_n1183_n661# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X401 a_922_n2811# a_649_n2805# a_837_n2811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X402 sky130_fd_sc_hd__inv_4_6/A sky130_fd_sc_hd__inv_1_6/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X403 VDD a_1347_n1901# a_1515_n1999# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X404 a_n1608_n2837# a_n1776_n2811# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X405 VSS sky130_fd_sc_hd__inv_4_2/A sky130_fd_sc_hd__inv_4_2/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X406 VDD a_1515_n2837# a_1946_n2811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X407 a_n1861_n91# sky130_fd_sc_hd__inv_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X408 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__inv_4_7/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X409 sky130_fd_sc_hd__inv_4_4/Y sky130_fd_sc_hd__inv_4_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X410 sky130_fd_sc_hd__inv_4_2/A sky130_fd_sc_hd__inv_1_2/A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X411 VSS a_n1351_n1901# a_n1183_n1999# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X412 a_922_n1901# a_649_n2267# a_837_n2267# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X413 sky130_fd_sc_hd__inv_4_6/Y sky130_fd_sc_hd__inv_4_6/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X414 VDD sky130_fd_sc_hd__inv_4_5/A sky130_fd_sc_hd__inv_4_5/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X415 sky130_fd_sc_hd__inv_4_4/Y sky130_fd_sc_hd__inv_4_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X416 a_n1267_n635# a_n2049_n629# a_n1351_n635# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X417 VSS sky130_fd_sc_hd__dfxbp_1_8/Q a_483_n1179# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
C0 a_n2049_n2267# sky130_fd_sc_hd__inv_4_4/Y 0.61fF
C1 VDD vin 0.16fF
C2 a_649_n1179# sky130_fd_sc_hd__dfxbp_1_7/Q 0.03fF
C3 a_n1861_n1179# sky130_fd_sc_hd__inv_4_3/Y 0.38fF
C4 a_n2215_n2267# a_n2215_n1717# 0.20fF
C5 a_n1776_n635# a_n1183_n661# 0.02fF
C6 a_n1861_n2267# a_n2215_n2267# 0.21fF
C7 sky130_fd_sc_hd__dfxbp_1_10/Q sky130_fd_sc_hd__inv_1_10/A 0.07fF
C8 VDD sky130_fd_sc_hd__inv_4_8/A 0.62fF
C9 a_1515_n1999# VDD 0.45fF
C10 a_483_n629# a_1090_n661# 0.37fF
C11 sky130_fd_sc_hd__dfxbp_1_9/Q sky130_fd_sc_hd__inv_1_9/A 0.07fF
C12 VDD a_n752_n635# 0.37fF
C13 a_483_n1717# a_837_n1723# 0.21fF
C14 VDD a_n2049_n629# 0.43fF
C15 a_922_n813# a_483_n1179# 0.63fF
C16 sky130_fd_sc_hd__inv_4_10/Y a_1515_n2837# 0.17fF
C17 a_n1861_n91# a_n2049_n91# 0.26fF
C18 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__dfxbp_1_8/Q 0.42fF
C19 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_4_7/Y 0.27fF
C20 sky130_fd_sc_hd__dfxbp_1_1/Q VDD 2.18fF
C21 sky130_fd_sc_hd__inv_1_1/A a_n752_n635# 0.25fF
C22 a_922_n813# a_1017_n813# 0.04fF
C23 a_1946_n857# a_1946_n1723# 0.04fF
C24 a_n1776_n813# sky130_fd_sc_hd__inv_4_3/Y 0.16fF
C25 VDD a_n2049_n91# 0.43fF
C26 a_n752_231# a_n1183_177# 0.31fF
C27 a_1515_n661# a_649_n629# 0.11fF
C28 sky130_fd_sc_hd__dfxbp_1_1/Q sky130_fd_sc_hd__inv_1_1/A 0.07fF
C29 a_n1351_n1901# a_n1267_n1901# 0.05fF
C30 a_n1351_n1901# sky130_fd_sc_hd__inv_4_4/Y 0.14fF
C31 a_1515_n1999# sky130_fd_sc_hd__inv_1_9/A 0.04fF
C32 a_1515_n661# a_1515_n911# 0.09fF
C33 VDD a_n752_n2811# 0.37fF
C34 a_n1351_n2811# sky130_fd_sc_hd__dfxbp_1_5/Q 0.04fF
C35 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__inv_4_7/A 1.64fF
C36 a_n1776_n1901# a_n1776_n2811# 0.05fF
C37 sky130_fd_sc_hd__dfxbp_1_9/Q a_837_n1723# 0.02fF
C38 a_1515_n1749# a_1946_n1723# 0.31fF
C39 a_n1776_275# a_n2049_n91# 0.38fF
C40 sky130_fd_sc_hd__inv_4_5/Y a_n1861_n2811# 0.38fF
C41 a_1515_n1749# a_922_n1723# 0.02fF
C42 a_n1183_n1999# sky130_fd_sc_hd__dfxbp_1_2/Q 0.02fF
C43 VDD a_1017_n1901# 0.02fF
C44 a_n1183_n661# a_n752_n635# 0.31fF
C45 a_n1608_n1749# a_n1351_n1723# 0.11fF
C46 sky130_fd_sc_hd__inv_4_10/Y sky130_fd_sc_hd__inv_4_9/Y 0.13fF
C47 a_n2049_n2267# a_n1351_n2811# 0.01fF
C48 a_837_n2267# a_649_n2267# 0.26fF
C49 sky130_fd_sc_hd__inv_4_0/A sky130_fd_sc_hd__inv_4_0/Y 1.64fF
C50 a_1347_n813# a_649_n1717# 0.01fF
C51 a_n1351_n813# a_n2049_n1179# 0.44fF
C52 VDD a_n2215_n629# 0.79fF
C53 a_1946_n857# a_1515_n911# 0.31fF
C54 a_n1183_n661# a_n2049_n629# 0.11fF
C55 a_n1351_n2811# a_n1183_n2837# 0.67fF
C56 VDD a_1347_n813# 0.22fF
C57 a_n1861_n2811# a_n1776_n2811# 0.11fF
C58 a_n1351_275# a_n2049_n629# 0.01fF
C59 VDD sky130_fd_sc_hd__dfxbp_1_2/Q 2.18fF
C60 sky130_fd_sc_hd__dfxbp_1_1/Q a_n1183_n661# 0.39fF
C61 a_837_n2267# sky130_fd_sc_hd__inv_4_9/Y 0.38fF
C62 a_n2215_n2805# a_n1351_n2811# 0.09fF
C63 a_n1608_n661# sky130_fd_sc_hd__inv_4_1/Y 0.15fF
C64 a_649_n2267# sky130_fd_sc_hd__inv_4_9/Y 0.61fF
C65 sky130_fd_sc_hd__dfxbp_1_8/Q a_483_n1717# 0.03fF
C66 sky130_fd_sc_hd__dfxbp_1_0/Q a_n1183_177# 0.39fF
C67 a_922_n1901# a_1090_n2155# 0.59fF
C68 a_n752_n1945# a_n1351_n1901# 0.02fF
C69 VDD a_483_n2805# 0.78fF
C70 sky130_fd_sc_hd__dfxbp_1_3/Q a_n752_n857# 0.37fF
C71 a_n1351_275# a_n2049_n91# 0.44fF
C72 sky130_fd_sc_hd__inv_4_5/Y a_n2049_n2805# 0.61fF
C73 a_483_n629# a_922_n635# 0.63fF
C74 sky130_fd_sc_hd__dfxbp_1_3/Q sky130_fd_sc_hd__inv_4_3/Y 0.41fF
C75 a_n1776_275# a_n2215_n629# 0.01fF
C76 a_1090_n1749# a_649_n1717# 0.28fF
C77 a_n2049_n1717# a_n1351_n1723# 0.44fF
C78 a_n1183_177# a_n1608_21# 0.04fF
C79 a_483_n2805# a_1347_n2811# 0.09fF
C80 a_483_n2267# a_649_n2805# 0.02fF
C81 a_n2049_n2805# a_n1776_n2811# 0.38fF
C82 a_1515_n1749# a_1515_n911# 0.09fF
C83 VDD a_1090_n1749# 0.23fF
C84 a_n1608_n1067# a_n1608_n1749# 0.05fF
C85 a_n2049_n1717# a_n2049_n2267# 0.05fF
C86 a_n2215_n1179# VDD 0.79fF
C87 VDD a_n2215_n1717# 0.79fF
C88 a_n1776_n1723# a_n1608_n1749# 0.59fF
C89 VDD a_1090_n1067# 0.23fF
C90 VDD a_n1861_n2267# 0.15fF
C91 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_4/A 0.04fF
C92 a_n1351_n2811# a_n1608_n2837# 0.11fF
C93 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__dfxbp_1_7/Q 0.29fF
C94 a_n752_n857# sky130_fd_sc_hd__inv_4_3/Y 0.11fF
C95 sky130_fd_sc_hd__inv_4_2/Y sky130_fd_sc_hd__inv_4_4/Y 0.06fF
C96 a_n1183_n1749# sky130_fd_sc_hd__dfxbp_1_3/Q 0.02fF
C97 a_n1776_n813# a_n1351_n813# 0.03fF
C98 a_n1351_n1901# a_n1351_n2811# 0.07fF
C99 sky130_fd_sc_hd__inv_4_2/A sky130_fd_sc_hd__inv_1_2/A 0.35fF
C100 a_483_n2267# a_1090_n2155# 0.37fF
C101 sky130_fd_sc_hd__dfxbp_1_9/Q sky130_fd_sc_hd__dfxbp_1_8/Q 0.08fF
C102 a_n2215_n629# a_n1183_n661# 0.11fF
C103 VDD a_837_n2811# 0.15fF
C104 a_1048_n2433# a_922_n2811# 0.02fF
C105 a_922_n1901# a_1347_n1901# 0.03fF
C106 a_n2049_n2267# a_n1608_n2155# 0.28fF
C107 sky130_fd_sc_hd__inv_4_0/Y vin 0.05fF
C108 a_1515_n661# a_1946_n635# 0.31fF
C109 a_649_n2805# sky130_fd_sc_hd__dfxbp_1_5/Q 0.06fF
C110 a_n752_n857# sky130_fd_sc_hd__inv_4_3/A 0.05fF
C111 a_1515_n661# a_1347_n635# 0.67fF
C112 a_1473_n2433# a_1347_n2811# 0.04fF
C113 sky130_fd_sc_hd__dfxbp_1_4/Q sky130_fd_sc_hd__dfxbp_1_2/Q 0.08fF
C114 sky130_fd_sc_hd__inv_4_3/Y sky130_fd_sc_hd__inv_4_3/A 1.64fF
C115 sky130_fd_sc_hd__inv_1_2/A VDD 0.48fF
C116 a_n1351_275# a_n1225_n91# 0.04fF
C117 a_n1776_n1723# a_n1681_n1723# 0.04fF
C118 a_n1776_n1723# a_n2049_n1717# 0.38fF
C119 VDD a_1946_n1945# 0.37fF
C120 VDD sky130_fd_sc_hd__inv_4_1/A 0.62fF
C121 a_n2215_n91# a_n1776_n635# 0.01fF
C122 a_1347_n1723# a_649_n1717# 0.44fF
C123 VDD a_922_n813# 0.36fF
C124 VDD a_1347_n1723# 0.22fF
C125 VDD sky130_fd_sc_hd__dfxbp_1_10/Q 0.38fF
C126 a_1347_n1901# a_483_n2267# 0.09fF
C127 a_649_n2805# a_1090_n2837# 0.28fF
C128 sky130_fd_sc_hd__dfxbp_1_10/Q sky130_fd_sc_hd__inv_4_4/A 0.02fF
C129 sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__inv_1_1/A 0.35fF
C130 a_1946_n857# a_1946_n635# 0.04fF
C131 VDD sky130_fd_sc_hd__inv_1_10/A 0.48fF
C132 sky130_fd_sc_hd__inv_4_10/Y sky130_fd_sc_hd__inv_4_10/A 1.64fF
C133 VDD a_n1681_275# 0.02fF
C134 sky130_fd_sc_hd__inv_4_0/Y a_n2049_n91# 0.61fF
C135 a_922_n1723# a_1017_n1723# 0.04fF
C136 sky130_fd_sc_hd__dfxbp_1_10/Q a_1347_n2811# 0.05fF
C137 a_1515_n661# sky130_fd_sc_hd__inv_1_6/A 0.04fF
C138 a_483_n1179# a_649_n1717# 0.02fF
C139 a_922_n2811# a_649_n2805# 0.38fF
C140 a_n1608_n2155# a_n1608_n2837# 0.05fF
C141 sky130_fd_sc_hd__inv_1_9/A a_1946_n1945# 0.25fF
C142 a_1515_n661# a_1090_n661# 0.04fF
C143 a_n1351_n1901# a_n1608_n2155# 0.11fF
C144 sky130_fd_sc_hd__inv_4_0/A sky130_fd_sc_hd__inv_4_1/Y 0.03fF
C145 a_1090_n2155# a_1090_n2837# 0.05fF
C146 VDD a_483_n1179# 0.78fF
C147 a_1090_n1749# a_837_n1723# 0.04fF
C148 a_n1608_n661# a_n1608_21# 0.05fF
C149 sky130_fd_sc_hd__inv_4_7/A sky130_fd_sc_hd__inv_4_8/A 0.10fF
C150 a_n1267_n2811# a_n1351_n2811# 0.05fF
C151 VDD a_n1183_n911# 0.45fF
C152 a_n1351_n813# sky130_fd_sc_hd__dfxbp_1_3/Q 0.05fF
C153 VDD a_1017_n813# 0.02fF
C154 a_n1861_n1723# a_n1608_n1749# 0.04fF
C155 sky130_fd_sc_hd__inv_4_9/Y sky130_fd_sc_hd__inv_4_10/A 0.03fF
C156 a_n2049_n1179# a_n1351_n1723# 0.01fF
C157 sky130_fd_sc_hd__inv_4_2/Y a_n1608_n1749# 0.15fF
C158 a_n1776_n635# sky130_fd_sc_hd__inv_4_1/Y 0.16fF
C159 a_n2215_n91# vin 0.41fF
C160 sky130_fd_sc_hd__inv_1_9/A sky130_fd_sc_hd__inv_1_10/A 0.04fF
C161 a_n1776_275# a_n1681_275# 0.04fF
C162 sky130_fd_sc_hd__inv_4_6/Y a_837_n635# 0.38fF
C163 sky130_fd_sc_hd__inv_4_6/A sky130_fd_sc_hd__inv_4_6/Y 1.64fF
C164 a_n1351_n813# a_n1267_n813# 0.05fF
C165 a_n1183_n1999# a_n2215_n2267# 0.11fF
C166 a_n1351_n813# a_n752_n857# 0.02fF
C167 VDD a_n2215_n2267# 0.79fF
C168 sky130_fd_sc_hd__dfxbp_1_2/Q sky130_fd_sc_hd__inv_4_4/Y 0.30fF
C169 VDD a_837_n635# 0.15fF
C170 sky130_fd_sc_hd__inv_4_6/A VDD 0.62fF
C171 a_n1351_n813# sky130_fd_sc_hd__inv_4_3/Y 0.14fF
C172 sky130_fd_sc_hd__inv_4_0/A a_n752_231# 0.05fF
C173 a_n2215_n91# a_n2049_n629# 0.02fF
C174 a_n1225_n1179# a_n1351_n813# 0.04fF
C175 sky130_fd_sc_hd__inv_4_5/Y sky130_fd_sc_hd__dfxbp_1_5/Q 0.66fF
C176 VDD sky130_fd_sc_hd__inv_4_5/A 0.62fF
C177 a_922_n1901# a_922_n1723# 0.08fF
C178 sky130_fd_sc_hd__inv_4_4/A sky130_fd_sc_hd__inv_4_5/A 0.10fF
C179 a_n1861_n1723# a_n2049_n1717# 0.26fF
C180 a_n752_n1945# a_n752_n2811# 0.04fF
C181 a_1347_n635# a_649_n629# 0.44fF
C182 a_922_n1901# a_837_n2267# 0.11fF
C183 a_n1608_n661# a_n1861_n635# 0.04fF
C184 a_1347_n1723# a_1473_n1345# 0.04fF
C185 sky130_fd_sc_hd__inv_4_8/Y a_1946_n1723# 0.11fF
C186 a_n1861_n2811# a_n2049_n2805# 0.26fF
C187 sky130_fd_sc_hd__inv_1_5/A sky130_fd_sc_hd__dfxbp_1_5/Q 0.15fF
C188 a_922_n1901# a_649_n2267# 0.38fF
C189 a_n1608_n1067# a_n2049_n1179# 0.28fF
C190 sky130_fd_sc_hd__inv_4_2/Y a_n2049_n1717# 0.61fF
C191 sky130_fd_sc_hd__inv_4_8/Y a_922_n1723# 0.16fF
C192 a_n2049_n91# a_n2215_n91# 2.23fF
C193 a_649_n1179# a_649_n629# 0.05fF
C194 sky130_fd_sc_hd__inv_4_6/Y vout 0.10fF
C195 a_922_n1901# sky130_fd_sc_hd__inv_4_9/Y 0.16fF
C196 a_1515_n1749# sky130_fd_sc_hd__inv_4_8/Y 0.17fF
C197 VDD sky130_fd_sc_hd__inv_1_0/A 0.48fF
C198 a_649_n1179# a_1515_n911# 0.11fF
C199 a_n1183_n911# a_n1183_n661# 0.09fF
C200 a_n1351_n813# a_n1351_n635# 0.05fF
C201 a_n1861_n2267# sky130_fd_sc_hd__inv_4_4/Y 0.38fF
C202 sky130_fd_sc_hd__inv_4_5/Y a_n1183_n2837# 0.17fF
C203 a_n1861_n1179# a_n1608_n1067# 0.04fF
C204 VDD vout 0.30fF
C205 sky130_fd_sc_hd__inv_4_8/Y sky130_fd_sc_hd__inv_4_9/Y 0.06fF
C206 sky130_fd_sc_hd__inv_4_5/Y a_n2215_n2805# 0.35fF
C207 sky130_fd_sc_hd__inv_1_5/A a_n1183_n2837# 0.04fF
C208 a_n752_n2811# a_n1351_n2811# 0.02fF
C209 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_0/A 0.04fF
C210 a_922_n1723# a_483_n2267# 0.02fF
C211 a_837_n2267# a_483_n2267# 0.21fF
C212 a_n1776_n2811# a_n1183_n2837# 0.02fF
C213 VDD a_n1681_n2811# 0.02fF
C214 sky130_fd_sc_hd__inv_4_1/Y a_n752_n635# 0.11fF
C215 a_483_n2267# a_649_n2267# 2.23fF
C216 a_n752_n857# a_n752_n1723# 0.04fF
C217 sky130_fd_sc_hd__inv_4_1/Y a_n2049_n629# 0.61fF
C218 a_n1776_n2811# a_n2215_n2805# 0.63fF
C219 a_1515_n661# a_922_n635# 0.02fF
C220 a_483_n2267# sky130_fd_sc_hd__inv_4_9/Y 0.35fF
C221 a_1090_n661# a_649_n629# 0.28fF
C222 a_n2215_n629# a_n2215_n91# 0.08fF
C223 sky130_fd_sc_hd__dfxbp_1_1/Q sky130_fd_sc_hd__inv_4_1/Y 0.29fF
C224 sky130_fd_sc_hd__dfxbp_1_4/Q a_n2215_n2267# 0.03fF
C225 a_n1776_n813# a_n1608_n1067# 0.59fF
C226 sky130_fd_sc_hd__inv_4_10/Y sky130_fd_sc_hd__dfxbp_1_5/Q 0.08fF
C227 sky130_fd_sc_hd__inv_1_8/A a_1946_n1723# 0.25fF
C228 a_n1776_n813# a_n1776_n1723# 0.05fF
C229 a_1090_n2837# a_1515_n2837# 0.04fF
C230 sky130_fd_sc_hd__inv_1_4/A a_n1183_n1999# 0.04fF
C231 sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__inv_4_0/Y 0.03fF
C232 a_n1183_n1749# a_n752_n1723# 0.31fF
C233 sky130_fd_sc_hd__inv_4_5/Y a_n1608_n2837# 0.15fF
C234 a_1515_n1749# sky130_fd_sc_hd__inv_1_8/A 0.04fF
C235 a_n1681_n813# a_n1776_n813# 0.04fF
C236 sky130_fd_sc_hd__inv_1_4/A VDD 0.48fF
C237 a_n752_n635# a_n752_231# 0.04fF
C238 a_1946_n857# sky130_fd_sc_hd__inv_4_7/Y 0.11fF
C239 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_4_4/A 0.35fF
C240 a_n1267_n635# VDD 0.02fF
C241 sky130_fd_sc_hd__dfxbp_1_10/Q sky130_fd_sc_hd__inv_4_4/Y 0.04fF
C242 a_922_n2811# a_1515_n2837# 0.02fF
C243 a_n1776_n2811# a_n1608_n2837# 0.59fF
C244 a_1946_n2811# a_1946_n1945# 0.04fF
C245 sky130_fd_sc_hd__inv_4_2/A VDD 0.62fF
C246 sky130_fd_sc_hd__inv_4_2/A sky130_fd_sc_hd__inv_4_4/A 0.09fF
C247 sky130_fd_sc_hd__dfxbp_1_8/Q a_1347_n1723# 0.05fF
C248 sky130_fd_sc_hd__inv_4_10/Y a_1090_n2837# 0.15fF
C249 VDD a_n1861_n91# 0.15fF
C250 VDD sky130_fd_sc_hd__inv_4_6/Y 0.93fF
C251 VDD a_1431_n2811# 0.02fF
C252 VDD a_n1183_n1999# 0.45fF
C253 sky130_fd_sc_hd__dfxbp_1_10/Q a_1946_n2811# 0.37fF
C254 VDD a_649_n1717# 0.43fF
C255 sky130_fd_sc_hd__dfxbp_1_3/Q sky130_fd_sc_hd__inv_1_3/A 0.07fF
C256 a_n2215_n629# sky130_fd_sc_hd__inv_4_1/Y 0.35fF
C257 sky130_fd_sc_hd__dfxbp_1_7/Q a_1347_n813# 0.05fF
C258 a_1431_n2811# a_1347_n2811# 0.05fF
C259 a_1946_n2811# sky130_fd_sc_hd__inv_1_10/A 0.25fF
C260 sky130_fd_sc_hd__inv_4_10/Y a_922_n2811# 0.16fF
C261 VDD sky130_fd_sc_hd__inv_4_4/A 0.62fF
C262 a_n1608_n1749# a_n2215_n1717# 0.37fF
C263 a_1515_n1999# a_1090_n2155# 0.04fF
C264 a_1347_n635# a_1946_n635# 0.02fF
C265 a_n2049_n1717# sky130_fd_sc_hd__dfxbp_1_2/Q 0.03fF
C266 VDD a_n1681_n635# 0.02fF
C267 sky130_fd_sc_hd__dfxbp_1_8/Q a_483_n1179# 0.49fF
C268 a_n1861_n1723# a_n1861_n1179# 0.02fF
C269 sky130_fd_sc_hd__dfxbp_1_0/Q vin 0.04fF
C270 VDD a_1347_n2811# 0.22fF
C271 sky130_fd_sc_hd__inv_1_3/A a_n752_n857# 0.25fF
C272 sky130_fd_sc_hd__dfxbp_1_9/Q a_1347_n1901# 0.05fF
C273 a_n1776_n813# a_n1776_n635# 0.08fF
C274 VDD sky130_fd_sc_hd__inv_1_1/A 0.48fF
C275 a_n1861_n91# a_n1776_275# 0.11fF
C276 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_4_3/Y 0.27fF
C277 a_n1861_n635# a_n1776_n635# 0.11fF
C278 a_n1608_n661# a_n1351_n635# 0.11fF
C279 a_n2215_n2267# sky130_fd_sc_hd__inv_4_4/Y 0.35fF
C280 VDD a_n1776_275# 0.36fF
C281 sky130_fd_sc_hd__dfxbp_1_0/Q a_n2049_n629# 0.08fF
C282 a_n1183_n1749# a_n1351_n1723# 0.67fF
C283 a_n2049_n2267# a_n1776_n1901# 0.38fF
C284 a_n2049_n1179# a_n2049_n629# 0.05fF
C285 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfxbp_1_4/Q 0.07fF
C286 VDD sky130_fd_sc_hd__inv_1_9/A 0.48fF
C287 a_922_n635# a_649_n629# 0.38fF
C288 a_n2215_n1179# a_n2049_n1717# 0.02fF
C289 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_4_3/A 0.35fF
C290 a_1017_n2811# a_922_n2811# 0.04fF
C291 a_649_n1179# a_837_n1179# 0.26fF
C292 a_n2049_n1717# a_n2215_n1717# 2.23fF
C293 sky130_fd_sc_hd__dfxbp_1_1/Q sky130_fd_sc_hd__dfxbp_1_0/Q 0.07fF
C294 sky130_fd_sc_hd__inv_4_5/A sky130_fd_sc_hd__inv_4_4/Y 0.03fF
C295 sky130_fd_sc_hd__inv_1_6/A a_1946_n635# 0.25fF
C296 sky130_fd_sc_hd__inv_4_7/Y a_1515_n911# 0.17fF
C297 VDD a_1431_n635# 0.02fF
C298 sky130_fd_sc_hd__dfxbp_1_1/Q a_n2049_n1179# 0.09fF
C299 a_n1776_n1901# a_n2215_n2805# 0.01fF
C300 a_1347_n1901# a_1515_n1999# 0.67fF
C301 sky130_fd_sc_hd__dfxbp_1_0/Q a_n2049_n91# 0.03fF
C302 a_1431_n813# a_1347_n813# 0.05fF
C303 a_n1183_n1999# sky130_fd_sc_hd__dfxbp_1_4/Q 0.39fF
C304 a_1347_n635# a_1090_n661# 0.11fF
C305 a_n1608_n1067# sky130_fd_sc_hd__inv_4_3/Y 0.15fF
C306 VDD a_n1183_n661# 0.45fF
C307 a_483_n629# a_922_n813# 0.02fF
C308 sky130_fd_sc_hd__inv_4_0/Y sky130_fd_sc_hd__inv_1_0/A 0.27fF
C309 sky130_fd_sc_hd__dfxbp_1_1/Q a_n1861_n1179# 0.02fF
C310 VDD a_n1351_275# 0.22fF
C311 VDD sky130_fd_sc_hd__dfxbp_1_4/Q 0.38fF
C312 a_n2049_n91# a_n1608_21# 0.28fF
C313 a_n2049_n2805# sky130_fd_sc_hd__dfxbp_1_5/Q 0.01fF
C314 a_n1861_n2267# a_n1608_n2155# 0.04fF
C315 a_n1861_n2811# a_n2215_n2805# 0.21fF
C316 a_922_n1723# a_483_n1717# 0.63fF
C317 sky130_fd_sc_hd__inv_1_1/A a_n1183_n661# 0.04fF
C318 a_483_n2805# a_649_n2805# 2.23fF
C319 sky130_fd_sc_hd__inv_4_10/Y sky130_fd_sc_hd__inv_4_9/A 0.03fF
C320 a_1515_n1749# a_483_n1717# 0.11fF
C321 a_n1776_n1723# a_n1776_n1901# 0.08fF
C322 a_837_n1723# a_649_n1717# 0.26fF
C323 sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__dfxbp_1_7/Q 0.02fF
C324 sky130_fd_sc_hd__inv_4_6/A sky130_fd_sc_hd__inv_4_7/A 0.09fF
C325 a_483_n1717# a_649_n2267# 0.09fF
C326 a_n1183_n1749# a_n1776_n1723# 0.02fF
C327 sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__inv_4_1/Y 1.66fF
C328 VDD a_837_n1723# 0.15fF
C329 a_n1776_n1723# a_n1650_n1345# 0.02fF
C330 a_483_n629# a_483_n1179# 0.20fF
C331 a_n1351_n1901# a_n1776_n1901# 0.03fF
C332 sky130_fd_sc_hd__dfxbp_1_0/Q a_n2215_n629# 0.49fF
C333 a_n2049_n2805# a_n2049_n2267# 0.06fF
C334 a_n1351_n1901# a_n1225_n2267# 0.04fF
C335 a_1347_n635# a_1473_n257# 0.04fF
C336 a_n2049_n1179# a_n2215_n629# 0.09fF
C337 a_n1776_275# a_n1351_275# 0.03fF
C338 a_n1861_n635# a_n2049_n629# 0.26fF
C339 a_n2049_n2805# a_n1183_n2837# 0.11fF
C340 sky130_fd_sc_hd__inv_4_9/A sky130_fd_sc_hd__inv_4_9/Y 1.66fF
C341 a_n2049_n2805# a_n2215_n2805# 2.23fF
C342 a_922_n1901# a_483_n2267# 0.63fF
C343 a_n1861_n2811# a_n1608_n2837# 0.04fF
C344 a_1090_n1749# a_1090_n2155# 0.03fF
C345 a_1515_n1999# a_1515_n2837# 0.09fF
C346 sky130_fd_sc_hd__dfxbp_1_7/Q a_483_n1179# 0.03fF
C347 a_n1351_n813# a_n1351_n1723# 0.07fF
C348 a_837_n2811# a_649_n2805# 0.26fF
C349 sky130_fd_sc_hd__inv_4_5/Y a_n752_n2811# 0.11fF
C350 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_4_4/Y 0.27fF
C351 sky130_fd_sc_hd__dfxbp_1_9/Q a_1515_n1749# 0.02fF
C352 a_n1861_n1723# sky130_fd_sc_hd__dfxbp_1_3/Q 0.02fF
C353 sky130_fd_sc_hd__dfxbp_1_9/Q a_649_n2267# 0.03fF
C354 sky130_fd_sc_hd__inv_1_5/A a_n752_n2811# 0.25fF
C355 a_483_n629# a_837_n635# 0.21fF
C356 sky130_fd_sc_hd__inv_4_2/A sky130_fd_sc_hd__inv_4_4/Y 0.01fF
C357 sky130_fd_sc_hd__inv_4_2/Y sky130_fd_sc_hd__dfxbp_1_3/Q 0.42fF
C358 sky130_fd_sc_hd__dfxbp_1_9/Q sky130_fd_sc_hd__inv_4_9/Y 0.29fF
C359 a_n1861_n91# sky130_fd_sc_hd__inv_4_0/Y 0.38fF
C360 a_n1183_n1999# sky130_fd_sc_hd__inv_4_4/Y 0.17fF
C361 a_n2215_n1179# a_n2049_n1179# 2.23fF
C362 a_n2049_n1179# a_n2215_n1717# 0.02fF
C363 a_1946_n1723# sky130_fd_sc_hd__inv_4_8/A 0.05fF
C364 a_n2049_n2805# a_n1608_n2837# 0.28fF
C365 VDD a_n1267_n1901# 0.02fF
C366 a_n2049_n2805# a_n1351_n1901# 0.01fF
C367 a_n1776_n813# a_n2215_n629# 0.02fF
C368 VDD sky130_fd_sc_hd__inv_4_4/Y 0.91fF
C369 VDD sky130_fd_sc_hd__inv_4_0/Y 0.96fF
C370 a_n1650_n2267# a_n1776_n1901# 0.02fF
C371 sky130_fd_sc_hd__dfxbp_1_10/Q a_649_n2805# 0.03fF
C372 sky130_fd_sc_hd__inv_4_8/Y sky130_fd_sc_hd__inv_1_8/A 0.27fF
C373 sky130_fd_sc_hd__dfxbp_1_7/Q a_837_n635# 0.02fF
C374 sky130_fd_sc_hd__inv_4_4/A sky130_fd_sc_hd__inv_4_4/Y 1.64fF
C375 a_1347_n635# a_922_n635# 0.03fF
C376 a_n1776_n635# a_n1351_n635# 0.03fF
C377 sky130_fd_sc_hd__dfxbp_1_8/Q a_649_n1717# 0.03fF
C378 a_1515_n1749# a_1515_n1999# 0.09fF
C379 a_n1608_n1067# a_n1351_n813# 0.11fF
C380 a_n2049_n1717# a_n2215_n2267# 0.09fF
C381 a_n1861_n1179# a_n2215_n1179# 0.21fF
C382 a_1515_n1999# a_649_n2267# 0.11fF
C383 sky130_fd_sc_hd__inv_4_2/Y sky130_fd_sc_hd__inv_4_3/Y 0.13fF
C384 a_n2215_n629# a_n1861_n635# 0.21fF
C385 a_649_n1179# sky130_fd_sc_hd__inv_4_7/Y 0.61fF
C386 VDD sky130_fd_sc_hd__dfxbp_1_8/Q 0.38fF
C387 sky130_fd_sc_hd__inv_4_9/Y sky130_fd_sc_hd__inv_4_8/A 0.01fF
C388 VDD sky130_fd_sc_hd__inv_1_7/A 0.48fF
C389 a_1515_n1999# sky130_fd_sc_hd__inv_4_9/Y 0.17fF
C390 VDD a_n1681_n1901# 0.02fF
C391 VDD a_1946_n2811# 0.37fF
C392 sky130_fd_sc_hd__inv_1_4/A a_n752_n1945# 0.25fF
C393 sky130_fd_sc_hd__inv_4_7/Y a_837_n1179# 0.38fF
C394 sky130_fd_sc_hd__inv_4_5/Y a_483_n2805# 0.04fF
C395 a_n752_n1723# a_n1351_n1723# 0.02fF
C396 sky130_fd_sc_hd__inv_4_2/Y sky130_fd_sc_hd__inv_4_3/A 0.03fF
C397 a_n1183_n1749# sky130_fd_sc_hd__inv_4_2/Y 0.17fF
C398 sky130_fd_sc_hd__dfxbp_1_1/Q sky130_fd_sc_hd__dfxbp_1_3/Q 0.08fF
C399 a_1946_n2811# a_1347_n2811# 0.02fF
C400 a_n752_n857# a_n752_n635# 0.04fF
C401 a_n1776_275# sky130_fd_sc_hd__inv_4_0/Y 0.16fF
C402 a_n1225_n1345# a_n1351_n1723# 0.04fF
C403 sky130_fd_sc_hd__inv_4_6/Y sky130_fd_sc_hd__inv_4_7/A 0.01fF
C404 a_n1608_n2155# a_n2215_n2267# 0.37fF
C405 a_922_n1901# a_922_n2811# 0.05fF
C406 sky130_fd_sc_hd__dfxbp_1_7/Q vout 0.03fF
C407 a_n1776_n813# a_n2215_n1179# 0.63fF
C408 a_n752_n1945# a_n1183_n1999# 0.31fF
C409 sky130_fd_sc_hd__inv_4_8/Y sky130_fd_sc_hd__inv_4_7/Y 0.13fF
C410 a_n1776_n813# a_n2215_n1717# 0.01fF
C411 a_1946_n857# a_1347_n813# 0.02fF
C412 VDD sky130_fd_sc_hd__inv_4_7/A 0.62fF
C413 a_1347_n1901# a_1946_n1945# 0.02fF
C414 a_922_n635# a_1090_n661# 0.59fF
C415 VDD a_n752_n1945# 0.37fF
C416 a_n752_n1945# sky130_fd_sc_hd__inv_4_4/A 0.05fF
C417 sky130_fd_sc_hd__dfxbp_1_1/Q sky130_fd_sc_hd__inv_4_3/Y 0.30fF
C418 a_483_n2805# a_1515_n2837# 0.11fF
C419 a_n1861_n91# a_n2215_n91# 0.21fF
C420 sky130_fd_sc_hd__inv_4_9/A sky130_fd_sc_hd__inv_4_10/A 0.10fF
C421 a_1347_n1901# a_1347_n1723# 0.05fF
C422 a_n1351_275# sky130_fd_sc_hd__inv_4_0/Y 0.14fF
C423 sky130_fd_sc_hd__dfxbp_1_4/Q sky130_fd_sc_hd__inv_4_4/Y 0.42fF
C424 a_n752_n635# a_n1351_n635# 0.02fF
C425 VDD a_n2215_n91# 0.79fF
C426 sky130_fd_sc_hd__inv_1_0/A a_n752_231# 0.25fF
C427 a_483_n2267# a_922_n2811# 0.01fF
C428 a_n2049_n1179# a_n1183_n911# 0.11fF
C429 a_n2049_n629# a_n1351_n635# 0.44fF
C430 a_483_n629# sky130_fd_sc_hd__inv_4_6/Y 0.35fF
C431 a_649_n1179# a_483_n1717# 0.02fF
C432 VDD a_n1351_n2811# 0.22fF
C433 sky130_fd_sc_hd__inv_4_10/Y a_483_n2805# 0.35fF
C434 VDD a_n1608_n1749# 0.23fF
C435 sky130_fd_sc_hd__dfxbp_1_3/Q sky130_fd_sc_hd__dfxbp_1_2/Q 0.08fF
C436 sky130_fd_sc_hd__dfxbp_1_1/Q a_n1351_n635# 0.05fF
C437 a_n1183_n2837# sky130_fd_sc_hd__dfxbp_1_5/Q 0.38fF
C438 a_n1351_n2811# a_n1225_n2433# 0.04fF
C439 a_483_n629# VDD 0.78fF
C440 a_n2049_n91# a_n1351_n635# 0.01fF
C441 a_483_n2805# a_649_n2267# 0.02fF
C442 a_922_n1901# a_483_n1717# 0.02fF
C443 sky130_fd_sc_hd__inv_4_6/Y sky130_fd_sc_hd__dfxbp_1_7/Q 0.30fF
C444 a_n1776_275# a_n2215_n91# 0.63fF
C445 a_922_n1723# a_1090_n1749# 0.59fF
C446 a_1515_n1749# a_1090_n1749# 0.04fF
C447 sky130_fd_sc_hd__inv_4_8/Y a_483_n1717# 0.35fF
C448 a_n1608_n1067# a_n1608_n661# 0.03fF
C449 a_n2049_n2267# a_n2215_n2805# 0.02fF
C450 VDD sky130_fd_sc_hd__dfxbp_1_7/Q 2.23fF
C451 a_1347_n813# a_1515_n911# 0.67fF
C452 a_n2215_n1179# sky130_fd_sc_hd__dfxbp_1_3/Q 0.03fF
C453 a_922_n813# a_1048_n1179# 0.02fF
C454 a_n752_n1945# sky130_fd_sc_hd__dfxbp_1_4/Q 0.37fF
C455 sky130_fd_sc_hd__dfxbp_1_3/Q a_n2215_n1717# 0.49fF
C456 VDD sky130_fd_sc_hd__inv_4_1/Y 0.91fF
C457 a_837_n2811# sky130_fd_sc_hd__inv_4_10/Y 0.38fF
C458 VDD a_n1681_n1723# 0.02fF
C459 a_n2049_n1717# VDD 0.43fF
C460 a_n2215_n2805# a_n1183_n2837# 0.11fF
C461 sky130_fd_sc_hd__inv_4_8/Y sky130_fd_sc_hd__inv_4_9/A 0.01fF
C462 a_n1650_n257# a_n1776_n635# 0.02fF
C463 a_n1776_n813# a_n1183_n911# 0.02fF
C464 sky130_fd_sc_hd__dfxbp_1_10/Q a_1515_n2837# 0.39fF
C465 a_n1183_n1749# sky130_fd_sc_hd__dfxbp_1_2/Q 0.39fF
C466 sky130_fd_sc_hd__dfxbp_1_0/Q sky130_fd_sc_hd__inv_1_0/A 0.07fF
C467 a_837_n2811# a_837_n2267# 0.02fF
C468 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_4_1/Y 0.27fF
C469 a_n2215_n629# a_n1351_n635# 0.09fF
C470 a_1515_n2837# sky130_fd_sc_hd__inv_1_10/A 0.04fF
C471 a_483_n1717# a_483_n2267# 0.20fF
C472 a_n1351_275# a_n2215_n91# 0.09fF
C473 a_922_n2811# a_1090_n2837# 0.59fF
C474 a_n1183_n1999# a_n1608_n2155# 0.04fF
C475 a_n1776_n1723# a_n1351_n1723# 0.03fF
C476 a_n2215_n1179# sky130_fd_sc_hd__inv_4_3/Y 0.35fF
C477 a_1946_n1723# a_1946_n1945# 0.04fF
C478 a_n1351_n1723# a_n1267_n1723# 0.05fF
C479 VDD a_n1608_n2155# 0.23fF
C480 sky130_fd_sc_hd__dfxbp_1_9/Q sky130_fd_sc_hd__inv_4_8/Y 0.30fF
C481 a_n1351_n1901# a_n1351_n1723# 0.05fF
C482 a_1515_n911# a_1090_n1067# 0.04fF
C483 a_1473_n1179# a_1347_n813# 0.04fF
C484 a_1946_n1723# a_1347_n1723# 0.02fF
C485 sky130_fd_sc_hd__dfxbp_1_10/Q sky130_fd_sc_hd__inv_4_10/Y 0.42fF
C486 VDD a_n752_231# 0.37fF
C487 a_n1351_n1901# a_n2049_n2267# 0.44fF
C488 a_922_n1723# a_1048_n1345# 0.02fF
C489 a_n1183_n2837# a_n1608_n2837# 0.04fF
C490 a_n1776_n1901# a_n1861_n2267# 0.11fF
C491 a_n1776_n1901# a_n2215_n1717# 0.02fF
C492 sky130_fd_sc_hd__inv_4_10/Y sky130_fd_sc_hd__inv_1_10/A 0.27fF
C493 a_922_n1723# a_922_n813# 0.05fF
C494 sky130_fd_sc_hd__inv_4_5/Y sky130_fd_sc_hd__inv_4_5/A 1.64fF
C495 a_n1183_n1749# a_n2215_n1717# 0.11fF
C496 a_n1776_n2811# a_n2215_n2267# 0.01fF
C497 sky130_fd_sc_hd__inv_4_2/Y a_n752_n1723# 0.11fF
C498 a_922_n1723# a_1347_n1723# 0.03fF
C499 a_n2215_n2805# a_n1608_n2837# 0.37fF
C500 a_1946_n1945# sky130_fd_sc_hd__inv_4_9/Y 0.11fF
C501 sky130_fd_sc_hd__dfxbp_1_10/Q a_837_n2267# 0.02fF
C502 a_1515_n1749# a_1347_n1723# 0.67fF
C503 VDD a_1431_n813# 0.02fF
C504 sky130_fd_sc_hd__inv_4_5/A sky130_fd_sc_hd__inv_1_5/A 0.35fF
C505 sky130_fd_sc_hd__dfxbp_1_10/Q a_649_n2267# 0.08fF
C506 VDD a_649_n2805# 0.43fF
C507 a_922_n635# a_1048_n257# 0.02fF
C508 a_922_n1901# a_1515_n1999# 0.02fF
C509 sky130_fd_sc_hd__dfxbp_1_9/Q a_483_n2267# 0.03fF
C510 a_n1608_n661# a_n1776_n635# 0.59fF
C511 a_n2049_n91# a_n1183_177# 0.11fF
C512 sky130_fd_sc_hd__inv_4_1/Y a_n1183_n661# 0.17fF
C513 sky130_fd_sc_hd__dfxbp_1_10/Q sky130_fd_sc_hd__inv_4_9/Y 0.42fF
C514 sky130_fd_sc_hd__inv_4_8/Y sky130_fd_sc_hd__inv_4_8/A 1.64fF
C515 a_n1861_n2811# a_n1861_n2267# 0.02fF
C516 a_649_n2805# a_1347_n2811# 0.44fF
C517 sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__inv_4_3/Y 0.01fF
C518 a_922_n1723# a_483_n1179# 0.01fF
C519 VDD a_1090_n2155# 0.23fF
C520 a_n752_n1945# sky130_fd_sc_hd__inv_4_4/Y 0.11fF
C521 a_1515_n661# vout 0.38fF
C522 sky130_fd_sc_hd__inv_1_2/A a_n1183_n1749# 0.04fF
C523 a_922_n813# a_1515_n911# 0.02fF
C524 sky130_fd_sc_hd__dfxbp_1_3/Q a_n1183_n911# 0.39fF
C525 sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__inv_4_3/A 0.09fF
C526 a_1515_n1999# a_483_n2267# 0.11fF
C527 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_4_7/A 0.35fF
C528 a_922_n635# a_1017_n635# 0.04fF
C529 a_n1776_n2811# a_n1681_n2811# 0.04fF
C530 VDD sky130_fd_sc_hd__dfxbp_1_0/Q 0.38fF
C531 a_n1861_n91# a_n1608_21# 0.04fF
C532 VDD a_n2049_n1179# 0.43fF
C533 a_1347_n635# a_1347_n813# 0.05fF
C534 sky130_fd_sc_hd__inv_4_0/Y a_n2215_n91# 0.35fF
C535 a_n1351_275# a_n752_231# 0.02fF
C536 a_649_n629# a_483_n1179# 0.09fF
C537 sky130_fd_sc_hd__inv_4_3/Y a_483_n1179# 0.04fF
C538 a_n752_n857# a_n1183_n911# 0.31fF
C539 a_649_n1179# a_1347_n813# 0.44fF
C540 a_1515_n911# a_483_n1179# 0.11fF
C541 VDD a_n1608_21# 0.23fF
C542 sky130_fd_sc_hd__inv_4_3/Y a_n1183_n911# 0.17fF
C543 sky130_fd_sc_hd__inv_4_2/Y a_n1351_n1723# 0.14fF
C544 a_1347_n1901# VDD 0.22fF
C545 a_n1861_n1179# VDD 0.15fF
C546 a_n1351_n813# a_n2215_n1179# 0.09fF
C547 sky130_fd_sc_hd__inv_1_8/A sky130_fd_sc_hd__inv_4_8/A 0.35fF
C548 a_922_n1901# a_1017_n1901# 0.04fF
C549 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_5/A 0.04fF
C550 a_n1608_n661# a_n2049_n629# 0.28fF
C551 a_1347_n1901# a_1347_n2811# 0.07fF
C552 a_n1183_n1749# a_n1183_n911# 0.09fF
C553 a_649_n629# a_837_n635# 0.26fF
C554 a_1515_n661# sky130_fd_sc_hd__inv_4_6/Y 0.17fF
C555 a_n1861_n91# a_n1861_n635# 0.02fF
C556 a_649_n1179# a_1090_n1067# 0.28fF
C557 a_n1776_275# a_n1608_21# 0.59fF
C558 sky130_fd_sc_hd__inv_4_0/Y sky130_fd_sc_hd__inv_4_1/Y 0.13fF
C559 a_922_n1901# a_483_n2805# 0.01fF
C560 sky130_fd_sc_hd__dfxbp_1_2/Q a_n752_n1723# 0.37fF
C561 sky130_fd_sc_hd__inv_4_5/Y VDD 0.91fF
C562 a_n1776_n813# VDD 0.36fF
C563 sky130_fd_sc_hd__inv_4_5/Y sky130_fd_sc_hd__inv_4_4/A 0.03fF
C564 a_n1861_n1723# a_n1776_n1723# 0.11fF
C565 a_n1776_n1901# a_n2215_n2267# 0.63fF
C566 sky130_fd_sc_hd__dfxbp_1_0/Q a_n1183_n661# 0.02fF
C567 sky130_fd_sc_hd__dfxbp_1_8/Q sky130_fd_sc_hd__dfxbp_1_7/Q 0.08fF
C568 a_1515_n661# VDD 0.45fF
C569 a_837_n1179# a_1090_n1067# 0.04fF
C570 VDD sky130_fd_sc_hd__inv_1_5/A 0.48fF
C571 sky130_fd_sc_hd__dfxbp_1_0/Q a_n1351_275# 0.05fF
C572 VDD a_n1861_n635# 0.15fF
C573 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__dfxbp_1_7/Q 0.07fF
C574 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__inv_4_8/A 0.03fF
C575 a_n1776_n1723# sky130_fd_sc_hd__inv_4_2/Y 0.16fF
C576 VDD a_n1776_n2811# 0.36fF
C577 a_n752_n2811# sky130_fd_sc_hd__dfxbp_1_5/Q 0.45fF
C578 a_649_n629# vout 0.01fF
C579 sky130_fd_sc_hd__inv_4_8/Y a_1090_n1749# 0.15fF
C580 a_n1351_275# a_n1608_21# 0.11fF
C581 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__inv_4_10/A 0.35fF
C582 a_n1608_n2155# sky130_fd_sc_hd__inv_4_4/Y 0.15fF
C583 a_483_n2805# a_483_n2267# 0.08fF
C584 a_1090_n661# a_1090_n1067# 0.03fF
C585 VDD a_1515_n2837# 0.45fF
C586 sky130_fd_sc_hd__inv_4_0/Y a_n752_231# 0.11fF
C587 VDD a_1431_n1901# 0.02fF
C588 a_1946_n857# VDD 0.37fF
C589 a_n1608_n661# a_n2215_n629# 0.37fF
C590 a_n752_n2811# a_n1183_n2837# 0.31fF
C591 a_1347_n2811# a_1515_n2837# 0.67fF
C592 a_649_n1179# a_922_n813# 0.38fF
C593 a_649_n1179# a_1347_n1723# 0.01fF
C594 sky130_fd_sc_hd__dfxbp_1_9/Q a_483_n1717# 0.51fF
C595 sky130_fd_sc_hd__inv_4_2/Y a_483_n1717# 0.04fF
C596 a_922_n813# a_837_n1179# 0.11fF
C597 a_n1351_n813# a_n1183_n911# 0.67fF
C598 a_n2049_n2805# a_n2215_n2267# 0.02fF
C599 VDD sky130_fd_sc_hd__inv_4_10/Y 0.93fF
C600 VDD a_1946_n1723# 0.37fF
C601 a_922_n1723# a_649_n1717# 0.38fF
C602 sky130_fd_sc_hd__inv_4_5/Y sky130_fd_sc_hd__dfxbp_1_4/Q 0.42fF
C603 a_483_n2805# sky130_fd_sc_hd__dfxbp_1_5/Q 0.41fF
C604 sky130_fd_sc_hd__inv_1_2/A a_n752_n1723# 0.25fF
C605 a_1515_n1749# a_649_n1717# 0.11fF
C606 a_649_n2267# a_649_n1717# 0.05fF
C607 sky130_fd_sc_hd__dfxbp_1_2/Q a_n1351_n1723# 0.05fF
C608 VDD a_922_n1723# 0.36fF
C609 sky130_fd_sc_hd__inv_4_10/Y a_1347_n2811# 0.14fF
C610 VDD a_837_n2267# 0.15fF
C611 a_n2049_n2267# sky130_fd_sc_hd__dfxbp_1_2/Q 0.09fF
C612 a_649_n1179# a_483_n1179# 2.23fF
C613 a_1515_n1749# VDD 0.45fF
C614 VDD a_649_n2267# 0.43fF
C615 VDD sky130_fd_sc_hd__dfxbp_1_3/Q 0.38fF
C616 sky130_fd_sc_hd__inv_4_8/Y a_1347_n1723# 0.14fF
C617 sky130_fd_sc_hd__inv_4_2/A sky130_fd_sc_hd__inv_4_3/Y 0.03fF
C618 a_483_n629# sky130_fd_sc_hd__dfxbp_1_7/Q 0.51fF
C619 a_n2049_n1717# a_n1608_n1749# 0.28fF
C620 a_837_n1179# a_483_n1179# 0.21fF
C621 VDD sky130_fd_sc_hd__inv_4_9/Y 0.93fF
C622 sky130_fd_sc_hd__inv_4_7/Y a_1347_n813# 0.14fF
C623 a_483_n629# sky130_fd_sc_hd__inv_4_1/Y 0.04fF
C624 a_649_n2267# a_1347_n2811# 0.01fF
C625 a_649_n629# sky130_fd_sc_hd__inv_4_6/Y 0.61fF
C626 a_n1267_n813# VDD 0.02fF
C627 sky130_fd_sc_hd__dfxbp_1_0/Q sky130_fd_sc_hd__inv_4_0/Y 0.42fF
C628 sky130_fd_sc_hd__inv_4_9/A sky130_fd_sc_hd__inv_4_8/A 0.09fF
C629 sky130_fd_sc_hd__inv_4_6/A a_1946_n635# 0.05fF
C630 VDD a_n752_n857# 0.37fF
C631 a_n1861_n1723# sky130_fd_sc_hd__inv_4_2/Y 0.38fF
C632 a_483_n2805# a_1090_n2837# 0.37fF
C633 sky130_fd_sc_hd__dfxbp_1_9/Q sky130_fd_sc_hd__inv_4_2/Y 0.02fF
C634 VDD a_1017_n2811# 0.02fF
C635 sky130_fd_sc_hd__inv_4_2/A sky130_fd_sc_hd__inv_4_3/A 0.10fF
C636 VDD a_649_n629# 0.43fF
C637 a_837_n2811# sky130_fd_sc_hd__dfxbp_1_5/Q 0.02fF
C638 VDD sky130_fd_sc_hd__inv_4_3/Y 0.91fF
C639 a_n2215_n1717# a_n1351_n1723# 0.09fF
C640 a_n1776_n635# a_n2049_n629# 0.38fF
C641 sky130_fd_sc_hd__dfxbp_1_10/Q a_483_n2267# 0.49fF
C642 a_n2049_n2267# a_n1861_n2267# 0.26fF
C643 a_n1776_n1901# a_n1183_n1999# 0.02fF
C644 a_n2049_n2267# a_n2215_n1717# 0.09fF
C645 a_n1267_n635# a_n1351_n635# 0.05fF
C646 sky130_fd_sc_hd__inv_4_0/Y a_n1608_21# 0.15fF
C647 a_n1183_n1749# a_n1183_n1999# 0.09fF
C648 a_n1608_n2155# a_n1608_n1749# 0.03fF
C649 VDD a_1515_n911# 0.45fF
C650 sky130_fd_sc_hd__dfxbp_1_7/Q sky130_fd_sc_hd__inv_4_1/Y 0.02fF
C651 a_483_n2805# a_922_n2811# 0.63fF
C652 VDD a_n1776_n1901# 0.36fF
C653 a_837_n635# a_837_n1179# 0.02fF
C654 a_n1183_n1749# VDD 0.45fF
C655 sky130_fd_sc_hd__inv_1_9/A sky130_fd_sc_hd__inv_4_9/Y 0.27fF
C656 sky130_fd_sc_hd__inv_4_7/Y a_1090_n1067# 0.15fF
C657 VDD sky130_fd_sc_hd__inv_4_3/A 0.62fF
C658 sky130_fd_sc_hd__dfxbp_1_9/Q a_1515_n1999# 0.39fF
C659 vout a_1946_n635# 0.37fF
C660 a_837_n2811# a_1090_n2837# 0.04fF
C661 VDD a_n1351_n635# 0.22fF
C662 a_1347_n635# vout 0.04fF
C663 sky130_fd_sc_hd__inv_4_6/A sky130_fd_sc_hd__inv_1_6/A 0.35fF
C664 sky130_fd_sc_hd__inv_1_0/A a_n1183_177# 0.04fF
C665 sky130_fd_sc_hd__dfxbp_1_10/Q sky130_fd_sc_hd__dfxbp_1_5/Q 0.06fF
C666 a_n1608_n1067# a_n2215_n1179# 0.37fF
C667 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_3/A 0.04fF
C668 a_n1861_n2811# VDD 0.15fF
C669 sky130_fd_sc_hd__inv_4_5/Y sky130_fd_sc_hd__inv_4_4/Y 0.13fF
C670 a_n1776_n1723# a_n2215_n1179# 0.01fF
C671 a_1090_n661# a_837_n635# 0.04fF
C672 a_n1776_n1723# a_n2215_n1717# 0.63fF
C673 a_837_n2811# a_922_n2811# 0.11fF
C674 a_1347_n1723# a_1431_n1723# 0.05fF
C675 a_922_n1723# a_837_n1723# 0.11fF
C676 a_837_n2267# a_837_n1723# 0.02fF
C677 sky130_fd_sc_hd__dfxbp_1_0/Q a_n2215_n91# 0.03fF
C678 a_n2215_n629# a_n1776_n635# 0.63fF
C679 a_n1776_n2811# a_n1650_n2433# 0.02fF
C680 sky130_fd_sc_hd__inv_4_7/Y a_922_n813# 0.16fF
C681 sky130_fd_sc_hd__inv_1_6/A vout 0.07fF
C682 a_n2049_n2805# VDD 0.43fF
C683 a_n2049_n91# vin 0.06fF
C684 a_922_n635# a_922_n813# 0.08fF
C685 a_n2215_n91# a_n1608_21# 0.37fF
C686 sky130_fd_sc_hd__dfxbp_1_1/Q a_n752_n635# 0.37fF
C687 VDD a_1017_n1723# 0.02fF
C688 sky130_fd_sc_hd__dfxbp_1_1/Q a_n2049_n629# 0.03fF
C689 a_1090_n1749# a_483_n1717# 0.37fF
C690 VDD sky130_fd_sc_hd__inv_4_10/A 0.62fF
C691 sky130_fd_sc_hd__inv_1_3/A a_n1183_n911# 0.04fF
C692 a_n1183_n661# a_n1351_n635# 0.67fF
C693 sky130_fd_sc_hd__inv_4_6/Y a_1946_n635# 0.11fF
C694 a_n2049_n91# a_n2049_n629# 0.06fF
C695 a_1946_n2811# a_1515_n2837# 0.31fF
C696 a_1347_n635# sky130_fd_sc_hd__inv_4_6/Y 0.14fF
C697 a_n1351_275# a_n1351_n635# 0.07fF
C698 a_n1351_n813# VDD 0.22fF
C699 sky130_fd_sc_hd__inv_4_7/Y a_483_n1179# 0.35fF
C700 a_n2215_n1179# a_n1776_n635# 0.02fF
C701 a_1946_n857# sky130_fd_sc_hd__inv_1_7/A 0.25fF
C702 a_922_n635# a_483_n1179# 0.02fF
C703 sky130_fd_sc_hd__inv_4_5/A sky130_fd_sc_hd__dfxbp_1_5/Q 0.14fF
C704 sky130_fd_sc_hd__inv_4_2/Y sky130_fd_sc_hd__dfxbp_1_2/Q 0.29fF
C705 a_n1861_n2811# sky130_fd_sc_hd__dfxbp_1_4/Q 0.02fF
C706 VDD a_1946_n635# 0.37fF
C707 sky130_fd_sc_hd__dfxbp_1_0/Q sky130_fd_sc_hd__inv_4_1/Y 0.42fF
C708 VDD a_1347_n635# 0.22fF
C709 a_649_n1179# a_649_n1717# 0.06fF
C710 a_n2049_n1717# a_n2049_n1179# 0.06fF
C711 a_n2049_n2267# a_n2215_n2267# 2.23fF
C712 a_1946_n1723# sky130_fd_sc_hd__dfxbp_1_8/Q 0.37fF
C713 VDD a_n1183_177# 0.45fF
C714 a_649_n1179# VDD 0.43fF
C715 sky130_fd_sc_hd__inv_4_5/Y a_n1351_n2811# 0.14fF
C716 sky130_fd_sc_hd__inv_4_10/Y a_1946_n2811# 0.11fF
C717 a_n1608_n1067# a_n1183_n911# 0.04fF
C718 a_n2215_n2805# a_n2215_n2267# 0.08fF
C719 a_1515_n1749# sky130_fd_sc_hd__dfxbp_1_8/Q 0.39fF
C720 sky130_fd_sc_hd__inv_4_1/A sky130_fd_sc_hd__inv_4_0/A 0.10fF
C721 a_1946_n857# sky130_fd_sc_hd__inv_4_7/A 0.05fF
C722 a_n1861_n1723# a_n2215_n1717# 0.21fF
C723 VDD a_837_n1179# 0.15fF
C724 a_n1861_n1723# a_n1861_n2267# 0.02fF
C725 a_n2215_n629# a_n2049_n629# 2.23fF
C726 sky130_fd_sc_hd__inv_4_6/A sky130_fd_sc_hd__inv_4_7/Y 0.01fF
C727 sky130_fd_sc_hd__inv_1_6/A sky130_fd_sc_hd__inv_4_6/Y 0.27fF
C728 a_n1776_n2811# a_n1351_n2811# 0.03fF
C729 a_922_n635# a_837_n635# 0.11fF
C730 sky130_fd_sc_hd__inv_4_2/A a_n752_n1723# 0.05fF
C731 a_n2049_n2805# sky130_fd_sc_hd__dfxbp_1_4/Q 0.08fF
C732 sky130_fd_sc_hd__inv_4_2/Y a_n2215_n1717# 0.35fF
C733 a_483_n1717# a_922_n813# 0.01fF
C734 a_922_n1901# VDD 0.36fF
C735 a_1515_n661# a_483_n629# 0.11fF
C736 sky130_fd_sc_hd__inv_4_9/A a_1946_n1945# 0.05fF
C737 a_483_n1717# a_1347_n1723# 0.09fF
C738 a_1090_n661# sky130_fd_sc_hd__inv_4_6/Y 0.15fF
C739 sky130_fd_sc_hd__dfxbp_1_1/Q a_n2215_n629# 0.03fF
C740 sky130_fd_sc_hd__dfxbp_1_0/Q a_n752_231# 0.37fF
C741 sky130_fd_sc_hd__inv_4_8/Y a_649_n1717# 0.61fF
C742 VDD sky130_fd_sc_hd__inv_1_6/A 0.48fF
C743 a_n1776_275# a_n1183_177# 0.02fF
C744 a_n2215_n629# a_n2049_n91# 0.02fF
C745 sky130_fd_sc_hd__inv_4_8/Y VDD 0.93fF
C746 a_1347_n635# a_1431_n635# 0.05fF
C747 a_n1776_n1723# a_n2215_n2267# 0.02fF
C748 VDD a_n752_n1723# 0.37fF
C749 a_n1650_n91# a_n1776_275# 0.02fF
C750 VDD a_1090_n661# 0.23fF
C751 sky130_fd_sc_hd__inv_4_3/Y sky130_fd_sc_hd__dfxbp_1_8/Q 0.04fF
C752 a_n1776_n1901# sky130_fd_sc_hd__inv_4_4/Y 0.16fF
C753 a_1515_n661# sky130_fd_sc_hd__dfxbp_1_7/Q 0.02fF
C754 sky130_fd_sc_hd__dfxbp_1_8/Q a_1515_n911# 0.02fF
C755 a_483_n1717# a_483_n1179# 0.08fF
C756 a_n1351_n1901# a_n2215_n2267# 0.09fF
C757 a_483_n2267# a_649_n1717# 0.09fF
C758 sky130_fd_sc_hd__dfxbp_1_9/Q a_1946_n1945# 0.37fF
C759 sky130_fd_sc_hd__inv_1_7/A a_1515_n911# 0.04fF
C760 a_n1861_n635# sky130_fd_sc_hd__inv_4_1/Y 0.38fF
C761 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_4_2/Y 0.27fF
C762 a_n2215_n1179# a_n2049_n629# 0.09fF
C763 VDD a_483_n2267# 0.78fF
C764 a_n1183_n661# a_n1183_177# 0.09fF
C765 sky130_fd_sc_hd__dfxbp_1_8/Q sky130_fd_sc_hd__inv_4_3/A 0.02fF
C766 a_n1681_n1901# a_n1776_n1901# 0.04fF
C767 sky130_fd_sc_hd__dfxbp_1_1/Q a_n2215_n1179# 0.51fF
C768 a_n1351_275# a_n1183_177# 0.67fF
C769 sky130_fd_sc_hd__dfxbp_1_9/Q sky130_fd_sc_hd__dfxbp_1_10/Q 0.07fF
C770 a_1347_n1901# a_649_n2805# 0.01fF
C771 a_1946_n857# sky130_fd_sc_hd__dfxbp_1_7/Q 0.37fF
C772 a_1515_n1999# a_1946_n1945# 0.31fF
C773 VDD a_n1608_n661# 0.23fF
C774 a_1347_n1901# a_1090_n2155# 0.11fF
C775 VDD sky130_fd_sc_hd__inv_1_8/A 0.48fF
C776 VDD sky130_fd_sc_hd__dfxbp_1_5/Q 1.02fF
C777 a_n1776_n813# a_n1650_n1179# 0.02fF
C778 sky130_fd_sc_hd__inv_4_1/A a_n752_n635# 0.05fF
C779 a_837_n1723# a_837_n1179# 0.02fF
C780 a_n2049_n2267# a_n1183_n1999# 0.11fF
C781 a_1515_n1999# sky130_fd_sc_hd__dfxbp_1_10/Q 0.02fF
C782 VDD a_1431_n1723# 0.02fF
C783 a_n1183_n1999# a_n1183_n2837# 0.09fF
C784 VDD a_n1351_n1723# 0.22fF
C785 a_n1861_n1179# a_n2049_n1179# 0.26fF
C786 sky130_fd_sc_hd__inv_4_0/A sky130_fd_sc_hd__inv_1_0/A 0.35fF
C787 VDD a_n2049_n2267# 0.43fF
C788 VDD sky130_fd_sc_hd__inv_1_3/A 0.48fF
C789 a_n2215_n1179# a_n2215_n629# 0.20fF
C790 sky130_fd_sc_hd__inv_4_7/Y sky130_fd_sc_hd__inv_4_6/Y 0.06fF
C791 sky130_fd_sc_hd__inv_4_8/Y a_837_n1723# 0.38fF
C792 a_922_n635# sky130_fd_sc_hd__inv_4_6/Y 0.16fF
C793 VDD a_n1183_n2837# 0.45fF
C794 a_483_n629# a_649_n629# 2.23fF
C795 a_1347_n813# a_1090_n1067# 0.11fF
C796 VDD a_1090_n2837# 0.23fF
C797 a_n2215_n1717# sky130_fd_sc_hd__dfxbp_1_2/Q 0.03fF
C798 a_n1861_n2267# sky130_fd_sc_hd__dfxbp_1_2/Q 0.02fF
C799 VDD a_n2215_n2805# 0.79fF
C800 a_n2049_n1717# sky130_fd_sc_hd__dfxbp_1_3/Q 0.08fF
C801 sky130_fd_sc_hd__inv_1_8/A sky130_fd_sc_hd__inv_1_9/A 0.04fF
C802 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_1/A 0.04fF
C803 VDD sky130_fd_sc_hd__inv_4_7/Y 0.93fF
C804 a_n1183_n1749# a_n1608_n1749# 0.04fF
C805 a_1347_n2811# a_1090_n2837# 0.11fF
C806 a_649_n2805# a_1515_n2837# 0.11fF
C807 VDD a_922_n635# 0.36fF
C808 a_1946_n2811# sky130_fd_sc_hd__inv_4_10/A 0.05fF
C809 VDD a_922_n2811# 0.36fF
C810 a_n1776_n813# a_n2049_n1179# 0.38fF
C811 a_n1267_275# VDD 0.02fF
C812 a_649_n629# sky130_fd_sc_hd__dfxbp_1_7/Q 0.09fF
C813 sky130_fd_sc_hd__inv_4_0/Y a_n1183_177# 0.17fF
C814 a_n1608_n661# a_n1183_n661# 0.04fF
C815 sky130_fd_sc_hd__dfxbp_1_0/Q a_n1861_n635# 0.02fF
C816 sky130_fd_sc_hd__inv_4_3/Y sky130_fd_sc_hd__inv_4_1/Y 0.06fF
C817 a_922_n2811# a_1347_n2811# 0.03fF
C818 a_n1608_n1067# VDD 0.23fF
C819 sky130_fd_sc_hd__dfxbp_1_1/Q a_n1183_n911# 0.02fF
C820 a_1090_n1749# a_1090_n1067# 0.05fF
C821 sky130_fd_sc_hd__dfxbp_1_7/Q a_1515_n911# 0.39fF
C822 a_n1776_n1723# VDD 0.36fF
C823 a_n1351_n1901# a_n1183_n1999# 0.67fF
C824 a_n2215_n1179# a_n2215_n1717# 0.08fF
C825 sky130_fd_sc_hd__dfxbp_1_4/Q sky130_fd_sc_hd__dfxbp_1_5/Q 0.04fF
C826 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__dfxbp_1_2/Q 0.07fF
C827 VDD a_n1267_n1723# 0.02fF
C828 a_837_n2811# a_483_n2805# 0.21fF
C829 a_649_n1179# sky130_fd_sc_hd__dfxbp_1_8/Q 0.08fF
C830 sky130_fd_sc_hd__inv_4_10/Y a_649_n2805# 0.61fF
C831 a_n1776_n813# a_n1861_n1179# 0.11fF
C832 a_1347_n1901# a_1473_n2267# 0.04fF
C833 VDD a_n1608_n2837# 0.23fF
C834 a_n1681_n813# VDD 0.02fF
C835 VDD a_n1351_n1901# 0.22fF
C836 sky130_fd_sc_hd__inv_4_1/Y sky130_fd_sc_hd__inv_4_3/A 0.01fF
C837 a_n1183_n1749# a_n2049_n1717# 0.11fF
C838 a_n1861_n1179# a_n1861_n635# 0.02fF
C839 a_922_n813# a_1347_n813# 0.03fF
C840 sky130_fd_sc_hd__dfxbp_1_8/Q a_837_n1179# 0.02fF
C841 a_1347_n813# a_1347_n1723# 0.07fF
C842 a_649_n2267# a_649_n2805# 0.06fF
C843 a_n2049_n2267# sky130_fd_sc_hd__dfxbp_1_4/Q 0.03fF
C844 sky130_fd_sc_hd__inv_4_1/Y a_n1351_n635# 0.14fF
C845 a_n2049_n2805# a_n1351_n2811# 0.44fF
C846 sky130_fd_sc_hd__dfxbp_1_4/Q a_n1183_n2837# 0.02fF
C847 a_922_n1901# a_1048_n2267# 0.02fF
C848 sky130_fd_sc_hd__dfxbp_1_4/Q a_n2215_n2805# 0.49fF
C849 sky130_fd_sc_hd__inv_4_8/Y sky130_fd_sc_hd__dfxbp_1_8/Q 0.41fF
C850 a_837_n2267# a_1090_n2155# 0.04fF
C851 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_6/A 0.04fF
C852 a_483_n1717# a_649_n1717# 2.23fF
C853 sky130_fd_sc_hd__dfxbp_1_10/Q a_483_n2805# 0.03fF
C854 a_n1776_n1901# a_n1608_n2155# 0.59fF
C855 VDD sky130_fd_sc_hd__inv_4_0/A 0.62fF
C856 a_649_n2267# a_1090_n2155# 0.28fF
C857 a_1347_n813# a_483_n1179# 0.09fF
C858 VDD a_483_n1717# 0.78fF
C859 sky130_fd_sc_hd__inv_4_5/Y sky130_fd_sc_hd__inv_1_5/A 0.27fF
C860 VDD a_1017_n635# 0.02fF
C861 a_1347_n1901# a_1431_n1901# 0.05fF
C862 a_483_n2267# sky130_fd_sc_hd__inv_4_4/Y 0.04fF
C863 sky130_fd_sc_hd__inv_4_5/Y a_n1776_n2811# 0.16fF
C864 a_1090_n2155# sky130_fd_sc_hd__inv_4_9/Y 0.15fF
C865 a_1090_n1749# a_1347_n1723# 0.11fF
C866 a_922_n813# a_1090_n1067# 0.59fF
C867 sky130_fd_sc_hd__inv_4_5/A a_n752_n2811# 0.05fF
C868 a_n1267_275# a_n1351_275# 0.05fF
C869 VDD a_n1776_n635# 0.36fF
C870 VDD sky130_fd_sc_hd__inv_4_9/A 0.62fF
C871 a_n2215_n91# a_n1183_177# 0.11fF
C872 a_n1681_n635# a_n1776_n635# 0.04fF
C873 sky130_fd_sc_hd__dfxbp_1_9/Q sky130_fd_sc_hd__inv_4_2/A 0.02fF
C874 sky130_fd_sc_hd__dfxbp_1_3/Q a_n2049_n1179# 0.03fF
C875 sky130_fd_sc_hd__inv_4_2/A sky130_fd_sc_hd__inv_4_2/Y 1.64fF
C876 sky130_fd_sc_hd__inv_4_8/Y sky130_fd_sc_hd__inv_4_7/A 0.03fF
C877 a_483_n629# a_1347_n635# 0.09fF
C878 a_n1351_n1901# sky130_fd_sc_hd__dfxbp_1_4/Q 0.05fF
C879 sky130_fd_sc_hd__dfxbp_1_9/Q a_649_n1717# 0.09fF
C880 a_1090_n1067# a_483_n1179# 0.37fF
C881 a_n752_n1945# a_n752_n1723# 0.04fF
C882 a_n2215_n2267# sky130_fd_sc_hd__dfxbp_1_2/Q 0.51fF
C883 a_1347_n1901# a_649_n2267# 0.44fF
C884 a_649_n1179# a_483_n629# 0.09fF
C885 a_n1267_n2811# VDD 0.02fF
C886 a_n2215_n1179# a_n1183_n911# 0.11fF
C887 sky130_fd_sc_hd__dfxbp_1_9/Q VDD 2.23fF
C888 a_n1861_n1723# VDD 0.15fF
C889 a_n1776_275# a_n1776_n635# 0.05fF
C890 a_n2049_n1179# sky130_fd_sc_hd__inv_4_3/Y 0.61fF
C891 a_n1351_n813# a_n2049_n1717# 0.01fF
C892 sky130_fd_sc_hd__inv_4_2/Y VDD 0.91fF
C893 sky130_fd_sc_hd__inv_1_8/A sky130_fd_sc_hd__dfxbp_1_8/Q 0.07fF
C894 sky130_fd_sc_hd__inv_4_9/A sky130_fd_sc_hd__inv_1_9/A 0.35fF
C895 a_1347_n1901# sky130_fd_sc_hd__inv_4_9/Y 0.14fF
C896 a_n1861_n91# vin 0.02fF
C897 sky130_fd_sc_hd__inv_4_2/Y sky130_fd_sc_hd__inv_4_4/A 0.01fF
C898 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_8/A 0.04fF
C899 a_n1225_n257# a_n1351_n635# 0.04fF
C900 a_1473_n2433# VSS 0.01fF
C901 a_1048_n2433# VSS 0.01fF
C902 a_837_n2811# VSS 0.20fF
C903 a_n1225_n2433# VSS 0.01fF
C904 a_n1650_n2433# VSS 0.01fF
C905 a_n1861_n2811# VSS 0.20fF
C906 sky130_fd_sc_hd__inv_4_10/A VSS 0.89fF
C907 sky130_fd_sc_hd__inv_1_10/A VSS 0.41fF
C908 a_1946_n2811# VSS 0.31fF
C909 a_1347_n2811# VSS 0.60fF
C910 a_1515_n2837# VSS 1.13fF
C911 a_922_n2811# VSS 0.49fF
C912 a_1090_n2837# VSS 0.61fF
C913 a_649_n2805# VSS 0.16fF
C914 sky130_fd_sc_hd__inv_4_10/Y VSS 0.25fF
C915 a_483_n2805# VSS 0.34fF
C916 sky130_fd_sc_hd__dfxbp_1_5/Q VSS 0.74fF
C917 sky130_fd_sc_hd__inv_4_5/A VSS 0.82fF
C918 sky130_fd_sc_hd__inv_1_5/A VSS 0.41fF
C919 a_n752_n2811# VSS 0.31fF
C920 a_n1351_n2811# VSS 0.60fF
C921 a_n1183_n2837# VSS 1.13fF
C922 a_n1776_n2811# VSS 0.49fF
C923 a_n1608_n2837# VSS 0.61fF
C924 a_n2049_n2805# VSS 0.16fF
C925 sky130_fd_sc_hd__inv_4_5/Y VSS 0.25fF
C926 a_n2215_n2805# VSS 0.34fF
C927 a_1473_n2267# VSS 0.01fF
C928 a_1048_n2267# VSS 0.01fF
C929 a_n1225_n2267# VSS 0.01fF
C930 a_837_n2267# VSS 0.20fF
C931 sky130_fd_sc_hd__inv_4_9/A VSS 0.89fF
C932 sky130_fd_sc_hd__inv_1_9/A VSS 0.41fF
C933 a_1946_n1945# VSS 0.31fF
C934 a_1347_n1901# VSS 0.60fF
C935 a_1515_n1999# VSS 1.13fF
C936 a_922_n1901# VSS 0.49fF
C937 a_1090_n2155# VSS 0.61fF
C938 a_649_n2267# VSS 0.16fF
C939 sky130_fd_sc_hd__inv_4_9/Y VSS 0.25fF
C940 a_483_n2267# VSS 0.34fF
C941 sky130_fd_sc_hd__dfxbp_1_10/Q VSS 0.30fF
C942 sky130_fd_sc_hd__dfxbp_1_4/Q VSS 0.30fF
C943 a_n1650_n2267# VSS 0.01fF
C944 a_n1861_n2267# VSS 0.20fF
C945 sky130_fd_sc_hd__inv_4_4/A VSS 0.82fF
C946 sky130_fd_sc_hd__inv_1_4/A VSS 0.41fF
C947 a_n752_n1945# VSS 0.31fF
C948 a_n1351_n1901# VSS 0.60fF
C949 a_n1183_n1999# VSS 1.13fF
C950 a_n1776_n1901# VSS 0.49fF
C951 a_n1608_n2155# VSS 0.61fF
C952 a_n2049_n2267# VSS 0.16fF
C953 sky130_fd_sc_hd__inv_4_4/Y VSS 0.25fF
C954 a_n2215_n2267# VSS 0.34fF
C955 a_1473_n1345# VSS 0.01fF
C956 a_1048_n1345# VSS 0.01fF
C957 a_837_n1723# VSS 0.20fF
C958 sky130_fd_sc_hd__dfxbp_1_2/Q VSS 0.39fF
C959 a_n1225_n1345# VSS 0.01fF
C960 a_n1650_n1345# VSS 0.01fF
C961 a_n1861_n1723# VSS 0.20fF
C962 sky130_fd_sc_hd__inv_4_8/A VSS 0.08fF
C963 sky130_fd_sc_hd__inv_1_8/A VSS 0.08fF
C964 a_1946_n1723# VSS 0.08fF
C965 a_1347_n1723# VSS 0.60fF
C966 a_1515_n1749# VSS 1.13fF
C967 a_922_n1723# VSS 0.49fF
C968 a_1090_n1749# VSS 0.61fF
C969 a_649_n1717# VSS 0.08fF
C970 sky130_fd_sc_hd__inv_4_8/Y VSS 0.10fF
C971 a_483_n1717# VSS 0.09fF
C972 sky130_fd_sc_hd__dfxbp_1_9/Q VSS 0.43fF
C973 sky130_fd_sc_hd__inv_4_2/A VSS 0.08fF
C974 sky130_fd_sc_hd__inv_1_2/A VSS 0.08fF
C975 a_n752_n1723# VSS 0.08fF
C976 a_n1351_n1723# VSS 0.60fF
C977 a_n1183_n1749# VSS 1.13fF
C978 a_n1776_n1723# VSS 0.49fF
C979 a_n1608_n1749# VSS 0.61fF
C980 a_n2049_n1717# VSS 1.17fF
C981 sky130_fd_sc_hd__inv_4_2/Y VSS 1.30fF
C982 a_n2215_n1717# VSS 1.52fF
C983 a_1473_n1179# VSS 0.01fF
C984 a_1048_n1179# VSS 0.01fF
C985 a_n1225_n1179# VSS 0.01fF
C986 a_837_n1179# VSS 0.20fF
C987 sky130_fd_sc_hd__inv_4_7/A VSS 0.89fF
C988 sky130_fd_sc_hd__inv_1_7/A VSS 0.41fF
C989 a_1946_n857# VSS 0.31fF
C990 a_1347_n813# VSS 0.60fF
C991 a_1515_n911# VSS 1.13fF
C992 a_922_n813# VSS 0.49fF
C993 a_1090_n1067# VSS 0.61fF
C994 a_649_n1179# VSS 0.16fF
C995 sky130_fd_sc_hd__inv_4_7/Y VSS 0.25fF
C996 a_483_n1179# VSS 0.34fF
C997 sky130_fd_sc_hd__dfxbp_1_8/Q VSS 0.30fF
C998 sky130_fd_sc_hd__dfxbp_1_3/Q VSS 2.29fF
C999 a_n1650_n1179# VSS 0.01fF
C1000 a_n1861_n1179# VSS 0.20fF
C1001 sky130_fd_sc_hd__inv_4_3/A VSS 0.82fF
C1002 sky130_fd_sc_hd__inv_1_3/A VSS 0.41fF
C1003 a_n752_n857# VSS 0.31fF
C1004 a_n1351_n813# VSS 0.60fF
C1005 a_n1183_n911# VSS 1.13fF
C1006 a_n1776_n813# VSS 0.49fF
C1007 a_n1608_n1067# VSS 0.61fF
C1008 a_n2049_n1179# VSS 0.16fF
C1009 sky130_fd_sc_hd__inv_4_3/Y VSS 0.25fF
C1010 a_n2215_n1179# VSS 0.34fF
C1011 vout VSS 0.58fF
C1012 a_1473_n257# VSS 0.01fF
C1013 a_1048_n257# VSS 0.01fF
C1014 a_837_n635# VSS 0.20fF
C1015 sky130_fd_sc_hd__dfxbp_1_1/Q VSS 0.30fF
C1016 a_n1225_n257# VSS 0.01fF
C1017 a_n1650_n257# VSS 0.01fF
C1018 a_n1861_n635# VSS 0.20fF
C1019 sky130_fd_sc_hd__inv_4_6/A VSS 0.89fF
C1020 sky130_fd_sc_hd__inv_1_6/A VSS 0.41fF
C1021 a_1946_n635# VSS 0.31fF
C1022 a_1347_n635# VSS 0.60fF
C1023 a_1515_n661# VSS 1.13fF
C1024 a_922_n635# VSS 0.49fF
C1025 a_1090_n661# VSS 0.61fF
C1026 a_649_n629# VSS 0.16fF
C1027 sky130_fd_sc_hd__inv_4_6/Y VSS 0.25fF
C1028 a_483_n629# VSS 0.34fF
C1029 sky130_fd_sc_hd__dfxbp_1_7/Q VSS 0.30fF
C1030 sky130_fd_sc_hd__inv_4_1/A VSS 0.82fF
C1031 sky130_fd_sc_hd__inv_1_1/A VSS 0.41fF
C1032 a_n752_n635# VSS 0.31fF
C1033 a_n1351_n635# VSS 0.60fF
C1034 a_n1183_n661# VSS 1.13fF
C1035 a_n1776_n635# VSS 0.49fF
C1036 a_n1608_n661# VSS 0.61fF
C1037 a_n2049_n629# VSS 0.16fF
C1038 sky130_fd_sc_hd__inv_4_1/Y VSS 0.25fF
C1039 a_n2215_n629# VSS 0.34fF
C1040 a_n1225_n91# VSS 0.01fF
C1041 sky130_fd_sc_hd__dfxbp_1_0/Q VSS 0.40fF
C1042 a_n1650_n91# VSS 0.01fF
C1043 a_n1861_n91# VSS 0.20fF
C1044 sky130_fd_sc_hd__inv_4_0/A VSS 1.38fF
C1045 sky130_fd_sc_hd__inv_1_0/A VSS 0.71fF
C1046 a_n752_231# VSS 0.29fF
C1047 a_n1351_275# VSS 0.60fF
C1048 a_n1183_177# VSS 1.13fF
C1049 a_n1776_275# VSS 0.49fF
C1050 a_n1608_21# VSS 0.61fF
C1051 a_n2049_n91# VSS 1.17fF
C1052 sky130_fd_sc_hd__inv_4_0/Y VSS 0.19fF
C1053 a_n2215_n91# VSS 1.52fF
C1054 vin VSS 0.75fF
C1055 VDD VSS 53.58fF
.ends

