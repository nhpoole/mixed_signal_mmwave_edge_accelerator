magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< locali >>
rect 8134 101294 8374 101328
rect 9976 101223 12393 101257
rect 8240 100983 8299 101017
rect 12365 100983 12393 101017
rect 8265 100838 8299 100983
rect 8265 100804 8358 100838
rect 8265 100612 8358 100646
rect 8265 100467 8299 100612
rect 8240 100433 8299 100467
rect 12365 100433 12393 100467
rect 8240 100193 8299 100227
rect 12365 100193 12393 100227
rect 8265 100048 8299 100193
rect 8265 100014 8358 100048
rect 8265 99822 8358 99856
rect 8265 99677 8299 99822
rect 8240 99643 8299 99677
rect 12365 99643 12393 99677
rect 8240 99403 8299 99437
rect 12365 99403 12393 99437
rect 8265 99258 8299 99403
rect 8265 99224 8358 99258
rect 8265 99032 8358 99066
rect 8265 98887 8299 99032
rect 8240 98853 8299 98887
rect 12365 98853 12393 98887
rect 8240 98613 8299 98647
rect 12365 98613 12393 98647
rect 8265 98468 8299 98613
rect 8265 98434 8358 98468
rect 8265 98242 8358 98276
rect 8265 98097 8299 98242
rect 8240 98063 8299 98097
rect 12365 98063 12393 98097
rect 8240 97823 8299 97857
rect 12365 97823 12393 97857
rect 8265 97678 8299 97823
rect 8265 97644 8358 97678
rect 8265 97452 8358 97486
rect 8265 97307 8299 97452
rect 8240 97273 8299 97307
rect 12365 97273 12393 97307
rect 8240 97033 8299 97067
rect 12365 97033 12393 97067
rect 8265 96888 8299 97033
rect 8265 96854 8358 96888
rect 8265 96662 8358 96696
rect 8265 96517 8299 96662
rect 8240 96483 8299 96517
rect 12365 96483 12393 96517
rect 8240 96243 8299 96277
rect 12365 96243 12393 96277
rect 8265 96098 8299 96243
rect 8265 96064 8358 96098
rect 8265 95872 8358 95906
rect 8265 95727 8299 95872
rect 8240 95693 8299 95727
rect 12365 95693 12393 95727
rect 8240 95453 8299 95487
rect 12365 95453 12393 95487
rect 8265 95308 8299 95453
rect 8265 95274 8358 95308
rect 8265 95082 8358 95116
rect 8265 94937 8299 95082
rect 8240 94903 8299 94937
rect 12365 94903 12393 94937
rect 8240 94663 8299 94697
rect 12365 94663 12393 94697
rect 8265 94518 8299 94663
rect 8265 94484 8358 94518
rect 8265 94292 8358 94326
rect 8265 94147 8299 94292
rect 8240 94113 8299 94147
rect 12365 94113 12393 94147
rect 8240 93873 8299 93907
rect 12365 93873 12393 93907
rect 8265 93728 8299 93873
rect 8265 93694 8358 93728
rect 8265 93502 8358 93536
rect 8265 93357 8299 93502
rect 8240 93323 8299 93357
rect 12365 93323 12393 93357
rect 8240 93083 8299 93117
rect 12365 93083 12393 93117
rect 8265 92938 8299 93083
rect 8265 92904 8358 92938
rect 8265 92712 8358 92746
rect 8265 92567 8299 92712
rect 8240 92533 8299 92567
rect 12365 92533 12393 92567
rect 8240 92293 8299 92327
rect 12365 92293 12393 92327
rect 8265 92148 8299 92293
rect 8265 92114 8358 92148
rect 8265 91922 8358 91956
rect 8265 91777 8299 91922
rect 8240 91743 8299 91777
rect 12365 91743 12393 91777
rect 8240 91503 8299 91537
rect 12365 91503 12393 91537
rect 8265 91358 8299 91503
rect 8265 91324 8358 91358
rect 8265 91132 8358 91166
rect 8265 90987 8299 91132
rect 8240 90953 8299 90987
rect 12365 90953 12393 90987
rect 8240 90713 8299 90747
rect 12365 90713 12393 90747
rect 8265 90568 8299 90713
rect 8265 90534 8358 90568
rect 8265 90342 8358 90376
rect 8265 90197 8299 90342
rect 8240 90163 8299 90197
rect 12365 90163 12393 90197
rect 8240 89923 8299 89957
rect 12365 89923 12393 89957
rect 8265 89778 8299 89923
rect 8265 89744 8358 89778
rect 8265 89552 8358 89586
rect 8265 89407 8299 89552
rect 8240 89373 8299 89407
rect 12365 89373 12393 89407
rect 8240 89133 8299 89167
rect 12365 89133 12393 89167
rect 8265 88988 8299 89133
rect 8265 88954 8358 88988
rect 8265 88762 8358 88796
rect 8265 88617 8299 88762
rect 8240 88583 8299 88617
rect 12365 88583 12393 88617
rect 8240 88343 8299 88377
rect 12365 88343 12393 88377
rect 8265 88198 8299 88343
rect 8265 88164 8358 88198
rect 8265 87972 8358 88006
rect 8265 87827 8299 87972
rect 8240 87793 8299 87827
rect 12365 87793 12393 87827
rect 8240 87553 8299 87587
rect 12365 87553 12393 87587
rect 8265 87408 8299 87553
rect 8265 87374 8358 87408
rect 8265 87182 8358 87216
rect 8265 87037 8299 87182
rect 8240 87003 8299 87037
rect 12365 87003 12393 87037
rect 8240 86763 8299 86797
rect 12365 86763 12393 86797
rect 8265 86618 8299 86763
rect 8265 86584 8358 86618
rect 8265 86392 8358 86426
rect 8265 86247 8299 86392
rect 8240 86213 8299 86247
rect 12365 86213 12393 86247
rect 8240 85973 8299 86007
rect 12365 85973 12393 86007
rect 8265 85828 8299 85973
rect 8265 85794 8358 85828
rect 8265 85602 8358 85636
rect 8265 85457 8299 85602
rect 8240 85423 8299 85457
rect 12365 85423 12393 85457
rect 8240 85183 8299 85217
rect 12365 85183 12393 85217
rect 8265 85038 8299 85183
rect 8265 85004 8358 85038
rect 8265 84812 8358 84846
rect 8265 84667 8299 84812
rect 8240 84633 8299 84667
rect 12365 84633 12393 84667
rect 8240 84393 8299 84427
rect 12365 84393 12393 84427
rect 8265 84248 8299 84393
rect 8265 84214 8358 84248
rect 8265 84022 8358 84056
rect 8265 83877 8299 84022
rect 8240 83843 8299 83877
rect 12365 83843 12393 83877
rect 8240 83603 8299 83637
rect 12365 83603 12393 83637
rect 8265 83458 8299 83603
rect 8265 83424 8358 83458
rect 8265 83232 8358 83266
rect 8265 83087 8299 83232
rect 8240 83053 8299 83087
rect 12365 83053 12393 83087
rect 8240 82813 8299 82847
rect 12365 82813 12393 82847
rect 8265 82668 8299 82813
rect 8265 82634 8358 82668
rect 8265 82442 8358 82476
rect 8265 82297 8299 82442
rect 8240 82263 8299 82297
rect 12365 82263 12393 82297
rect 8240 82023 8299 82057
rect 12365 82023 12393 82057
rect 8265 81878 8299 82023
rect 8265 81844 8358 81878
rect 8265 81652 8358 81686
rect 8265 81507 8299 81652
rect 8240 81473 8299 81507
rect 12365 81473 12393 81507
rect 8240 81233 8299 81267
rect 12365 81233 12393 81267
rect 8265 81088 8299 81233
rect 8265 81054 8358 81088
rect 8265 80862 8358 80896
rect 8265 80717 8299 80862
rect 8240 80683 8299 80717
rect 12365 80683 12393 80717
rect 8240 80443 8299 80477
rect 12365 80443 12393 80477
rect 8265 80298 8299 80443
rect 8265 80264 8358 80298
rect 8265 80072 8358 80106
rect 8265 79927 8299 80072
rect 8240 79893 8299 79927
rect 12365 79893 12393 79927
rect 8240 79653 8299 79687
rect 12365 79653 12393 79687
rect 8265 79508 8299 79653
rect 8265 79474 8358 79508
rect 8265 79282 8358 79316
rect 8265 79137 8299 79282
rect 8240 79103 8299 79137
rect 12365 79103 12393 79137
rect 8240 78863 8299 78897
rect 12365 78863 12393 78897
rect 8265 78718 8299 78863
rect 8265 78684 8358 78718
rect 8265 78492 8358 78526
rect 8265 78347 8299 78492
rect 8240 78313 8299 78347
rect 12365 78313 12393 78347
rect 8240 78073 8299 78107
rect 12365 78073 12393 78107
rect 8265 77928 8299 78073
rect 8265 77894 8358 77928
rect 8265 77702 8358 77736
rect 8265 77557 8299 77702
rect 8240 77523 8299 77557
rect 12365 77523 12393 77557
rect 8240 77283 8299 77317
rect 12365 77283 12393 77317
rect 8265 77138 8299 77283
rect 8265 77104 8358 77138
rect 8265 76912 8358 76946
rect 8265 76767 8299 76912
rect 8240 76733 8299 76767
rect 12365 76733 12393 76767
rect 8240 76493 8299 76527
rect 12365 76493 12393 76527
rect 8265 76348 8299 76493
rect 8265 76314 8358 76348
rect 8265 76122 8358 76156
rect 8265 75977 8299 76122
rect 8240 75943 8299 75977
rect 12365 75943 12393 75977
rect 8240 75703 8299 75737
rect 12365 75703 12393 75737
rect 8265 75558 8299 75703
rect 8265 75524 8358 75558
rect 8265 75332 8358 75366
rect 8265 75187 8299 75332
rect 8240 75153 8299 75187
rect 12365 75153 12393 75187
rect 8240 74913 8299 74947
rect 12365 74913 12393 74947
rect 8265 74768 8299 74913
rect 8265 74734 8358 74768
rect 8265 74542 8358 74576
rect 8265 74397 8299 74542
rect 8240 74363 8299 74397
rect 12365 74363 12393 74397
rect 8240 74123 8299 74157
rect 12365 74123 12393 74157
rect 8265 73978 8299 74123
rect 8265 73944 8358 73978
rect 8265 73752 8358 73786
rect 8265 73607 8299 73752
rect 8240 73573 8299 73607
rect 12365 73573 12393 73607
rect 8240 73333 8299 73367
rect 12365 73333 12393 73367
rect 8265 73188 8299 73333
rect 8265 73154 8358 73188
rect 8265 72962 8358 72996
rect 8265 72817 8299 72962
rect 8240 72783 8299 72817
rect 12365 72783 12393 72817
rect 8240 72543 8299 72577
rect 12365 72543 12393 72577
rect 8265 72398 8299 72543
rect 8265 72364 8358 72398
rect 8265 72172 8358 72206
rect 8265 72027 8299 72172
rect 8240 71993 8299 72027
rect 12365 71993 12393 72027
rect 8240 71753 8299 71787
rect 12365 71753 12393 71787
rect 8265 71608 8299 71753
rect 8265 71574 8358 71608
rect 8265 71382 8358 71416
rect 8265 71237 8299 71382
rect 8240 71203 8299 71237
rect 12365 71203 12393 71237
rect 8240 70963 8299 70997
rect 12365 70963 12393 70997
rect 8265 70818 8299 70963
rect 8265 70784 8358 70818
rect 8265 70592 8358 70626
rect 8265 70447 8299 70592
rect 8240 70413 8299 70447
rect 12365 70413 12393 70447
rect 8240 70173 8299 70207
rect 12365 70173 12393 70207
rect 8265 70028 8299 70173
rect 8265 69994 8358 70028
rect 8265 69802 8358 69836
rect 8265 69657 8299 69802
rect 8240 69623 8299 69657
rect 12365 69623 12393 69657
rect 8240 69383 8299 69417
rect 12365 69383 12393 69417
rect 8265 69238 8299 69383
rect 8265 69204 8358 69238
rect 8265 69012 8358 69046
rect 8265 68867 8299 69012
rect 8240 68833 8299 68867
rect 12365 68833 12393 68867
rect 8240 68593 8299 68627
rect 12365 68593 12393 68627
rect 8265 68448 8299 68593
rect 8265 68414 8358 68448
rect 8265 68222 8358 68256
rect 8265 68077 8299 68222
rect 8240 68043 8299 68077
rect 12365 68043 12393 68077
rect 8240 67803 8299 67837
rect 12365 67803 12393 67837
rect 8265 67658 8299 67803
rect 8265 67624 8358 67658
rect 8265 67432 8358 67466
rect 8265 67287 8299 67432
rect 8240 67253 8299 67287
rect 12365 67253 12393 67287
rect 8240 67013 8299 67047
rect 12365 67013 12393 67047
rect 8265 66868 8299 67013
rect 8265 66834 8358 66868
rect 8265 66642 8358 66676
rect 8265 66497 8299 66642
rect 8240 66463 8299 66497
rect 12365 66463 12393 66497
rect 8240 66223 8299 66257
rect 12365 66223 12393 66257
rect 8265 66078 8299 66223
rect 8265 66044 8358 66078
rect 8265 65852 8358 65886
rect 8265 65707 8299 65852
rect 8240 65673 8299 65707
rect 12365 65673 12393 65707
rect 8240 65433 8299 65467
rect 12365 65433 12393 65467
rect 8265 65288 8299 65433
rect 8265 65254 8358 65288
rect 8265 65062 8358 65096
rect 8265 64917 8299 65062
rect 8240 64883 8299 64917
rect 12365 64883 12393 64917
rect 8240 64643 8299 64677
rect 12365 64643 12393 64677
rect 8265 64498 8299 64643
rect 8265 64464 8358 64498
rect 8265 64272 8358 64306
rect 8265 64127 8299 64272
rect 8240 64093 8299 64127
rect 12365 64093 12393 64127
rect 8240 63853 8299 63887
rect 12365 63853 12393 63887
rect 8265 63708 8299 63853
rect 8265 63674 8358 63708
rect 8265 63482 8358 63516
rect 8265 63337 8299 63482
rect 8240 63303 8299 63337
rect 12365 63303 12393 63337
rect 8240 63063 8299 63097
rect 12365 63063 12393 63097
rect 8265 62918 8299 63063
rect 8265 62884 8358 62918
rect 8265 62692 8358 62726
rect 8265 62547 8299 62692
rect 8240 62513 8299 62547
rect 12365 62513 12393 62547
rect 8240 62273 8299 62307
rect 12365 62273 12393 62307
rect 8265 62128 8299 62273
rect 8265 62094 8358 62128
rect 8265 61902 8358 61936
rect 8265 61757 8299 61902
rect 8240 61723 8299 61757
rect 12365 61723 12393 61757
rect 8240 61483 8299 61517
rect 12365 61483 12393 61517
rect 8265 61338 8299 61483
rect 8265 61304 8358 61338
rect 8265 61112 8358 61146
rect 8265 60967 8299 61112
rect 8240 60933 8299 60967
rect 12365 60933 12393 60967
rect 8240 60693 8299 60727
rect 12365 60693 12393 60727
rect 8265 60548 8299 60693
rect 8265 60514 8358 60548
rect 8265 60322 8358 60356
rect 8265 60177 8299 60322
rect 8240 60143 8299 60177
rect 12365 60143 12393 60177
rect 8240 59903 8299 59937
rect 12365 59903 12393 59937
rect 8265 59758 8299 59903
rect 8265 59724 8358 59758
rect 8265 59532 8358 59566
rect 8265 59387 8299 59532
rect 8240 59353 8299 59387
rect 12365 59353 12393 59387
rect 8240 59113 8299 59147
rect 12365 59113 12393 59147
rect 8265 58968 8299 59113
rect 8265 58934 8358 58968
rect 8265 58742 8358 58776
rect 8265 58597 8299 58742
rect 8240 58563 8299 58597
rect 12365 58563 12393 58597
rect 8240 58323 8299 58357
rect 12365 58323 12393 58357
rect 8265 58178 8299 58323
rect 8265 58144 8358 58178
rect 8265 57952 8358 57986
rect 8265 57807 8299 57952
rect 8240 57773 8299 57807
rect 12365 57773 12393 57807
rect 8240 57533 8299 57567
rect 12365 57533 12393 57567
rect 8265 57388 8299 57533
rect 8265 57354 8358 57388
rect 8265 57162 8358 57196
rect 8265 57017 8299 57162
rect 8240 56983 8299 57017
rect 12365 56983 12393 57017
rect 8240 56743 8299 56777
rect 12365 56743 12393 56777
rect 8265 56598 8299 56743
rect 8265 56564 8358 56598
rect 8265 56372 8358 56406
rect 8265 56227 8299 56372
rect 8240 56193 8299 56227
rect 12365 56193 12393 56227
rect 8240 55953 8299 55987
rect 12365 55953 12393 55987
rect 8265 55808 8299 55953
rect 8265 55774 8358 55808
rect 8265 55582 8358 55616
rect 8265 55437 8299 55582
rect 8240 55403 8299 55437
rect 12365 55403 12393 55437
rect 8240 55163 8299 55197
rect 12365 55163 12393 55197
rect 8265 55018 8299 55163
rect 8265 54984 8358 55018
rect 8265 54792 8358 54826
rect 8265 54647 8299 54792
rect 8240 54613 8299 54647
rect 12365 54613 12393 54647
rect 8240 54373 8299 54407
rect 12365 54373 12393 54407
rect 8265 54228 8299 54373
rect 8265 54194 8358 54228
rect 8265 54002 8358 54036
rect 8265 53857 8299 54002
rect 8240 53823 8299 53857
rect 12365 53823 12393 53857
rect 8240 53583 8299 53617
rect 12365 53583 12393 53617
rect 8265 53438 8299 53583
rect 8265 53404 8358 53438
rect 8265 53212 8358 53246
rect 8265 53067 8299 53212
rect 8240 53033 8299 53067
rect 12365 53033 12393 53067
rect 8240 52793 8299 52827
rect 12365 52793 12393 52827
rect 8265 52648 8299 52793
rect 8265 52614 8358 52648
rect 8265 52422 8358 52456
rect 8265 52277 8299 52422
rect 8240 52243 8299 52277
rect 12365 52243 12393 52277
rect 8240 52003 8299 52037
rect 12365 52003 12393 52037
rect 8265 51858 8299 52003
rect 8265 51824 8358 51858
rect 8265 51632 8358 51666
rect 8265 51487 8299 51632
rect 8240 51453 8299 51487
rect 12365 51453 12393 51487
rect 8240 51213 8299 51247
rect 12365 51213 12393 51247
rect 8265 51068 8299 51213
rect 8265 51034 8358 51068
rect 8265 50842 8358 50876
rect 8265 50697 8299 50842
rect 8240 50663 8299 50697
rect 12365 50663 12393 50697
rect 8240 50423 8299 50457
rect 12365 50423 12393 50457
rect 8265 50278 8299 50423
rect 8265 50244 8358 50278
rect 8265 50052 8358 50086
rect 8265 49907 8299 50052
rect 8240 49873 8299 49907
rect 12365 49873 12393 49907
rect 8240 49633 8299 49667
rect 12365 49633 12393 49667
rect 8265 49488 8299 49633
rect 8265 49454 8358 49488
rect 8265 49262 8358 49296
rect 8265 49117 8299 49262
rect 8240 49083 8299 49117
rect 12365 49083 12393 49117
rect 8240 48843 8299 48877
rect 12365 48843 12393 48877
rect 8265 48698 8299 48843
rect 8265 48664 8358 48698
rect 8265 48472 8358 48506
rect 8265 48327 8299 48472
rect 8240 48293 8299 48327
rect 12365 48293 12393 48327
rect 8240 48053 8299 48087
rect 12365 48053 12393 48087
rect 8265 47908 8299 48053
rect 8265 47874 8358 47908
rect 8265 47682 8358 47716
rect 8265 47537 8299 47682
rect 8240 47503 8299 47537
rect 12365 47503 12393 47537
rect 8240 47263 8299 47297
rect 12365 47263 12393 47297
rect 8265 47118 8299 47263
rect 8265 47084 8358 47118
rect 8265 46892 8358 46926
rect 8265 46747 8299 46892
rect 8240 46713 8299 46747
rect 12365 46713 12393 46747
rect 8240 46473 8299 46507
rect 12365 46473 12393 46507
rect 8265 46328 8299 46473
rect 8265 46294 8358 46328
rect 8265 46102 8358 46136
rect 8265 45957 8299 46102
rect 8240 45923 8299 45957
rect 12365 45923 12393 45957
rect 8240 45683 8299 45717
rect 12365 45683 12393 45717
rect 8265 45538 8299 45683
rect 8265 45504 8358 45538
rect 8265 45312 8358 45346
rect 8265 45167 8299 45312
rect 8240 45133 8299 45167
rect 12365 45133 12393 45167
rect 8240 44893 8299 44927
rect 12365 44893 12393 44927
rect 8265 44748 8299 44893
rect 8265 44714 8358 44748
rect 8265 44522 8358 44556
rect 8265 44377 8299 44522
rect 8240 44343 8299 44377
rect 12365 44343 12393 44377
rect 8240 44103 8299 44137
rect 12365 44103 12393 44137
rect 8265 43958 8299 44103
rect 8265 43924 8358 43958
rect 8265 43732 8358 43766
rect 8265 43587 8299 43732
rect 8240 43553 8299 43587
rect 12365 43553 12393 43587
rect 8240 43313 8299 43347
rect 12365 43313 12393 43347
rect 8265 43168 8299 43313
rect 8265 43134 8358 43168
rect 8265 42942 8358 42976
rect 8265 42797 8299 42942
rect 8240 42763 8299 42797
rect 12365 42763 12393 42797
rect 8240 42523 8299 42557
rect 12365 42523 12393 42557
rect 8265 42378 8299 42523
rect 8265 42344 8358 42378
rect 8265 42152 8358 42186
rect 8265 42007 8299 42152
rect 8240 41973 8299 42007
rect 12365 41973 12393 42007
rect 8240 41733 8299 41767
rect 12365 41733 12393 41767
rect 8265 41588 8299 41733
rect 8265 41554 8358 41588
rect 8265 41362 8358 41396
rect 8265 41217 8299 41362
rect 8240 41183 8299 41217
rect 12365 41183 12393 41217
rect 8240 40943 8299 40977
rect 12365 40943 12393 40977
rect 8265 40798 8299 40943
rect 8265 40764 8358 40798
rect 8265 40572 8358 40606
rect 8265 40427 8299 40572
rect 8240 40393 8299 40427
rect 12365 40393 12393 40427
rect 8240 40153 8299 40187
rect 12365 40153 12393 40187
rect 8265 40008 8299 40153
rect 8265 39974 8358 40008
rect 8265 39782 8358 39816
rect 8265 39637 8299 39782
rect 8240 39603 8299 39637
rect 12365 39603 12393 39637
rect 8240 39363 8299 39397
rect 12365 39363 12393 39397
rect 8265 39218 8299 39363
rect 8265 39184 8358 39218
rect 8265 38992 8358 39026
rect 8265 38847 8299 38992
rect 8240 38813 8299 38847
rect 12365 38813 12393 38847
rect 8240 38573 8299 38607
rect 12365 38573 12393 38607
rect 8265 38428 8299 38573
rect 8265 38394 8358 38428
rect 8265 38202 8358 38236
rect 8265 38057 8299 38202
rect 8240 38023 8299 38057
rect 12365 38023 12393 38057
rect 8240 37783 8299 37817
rect 12365 37783 12393 37817
rect 8265 37638 8299 37783
rect 8265 37604 8358 37638
rect 8265 37412 8358 37446
rect 8265 37267 8299 37412
rect 8240 37233 8299 37267
rect 12365 37233 12393 37267
rect 8240 36993 8299 37027
rect 12365 36993 12393 37027
rect 8265 36848 8299 36993
rect 8265 36814 8358 36848
rect 8265 36622 8358 36656
rect 8265 36477 8299 36622
rect 8240 36443 8299 36477
rect 12365 36443 12393 36477
rect 8240 36203 8299 36237
rect 12365 36203 12393 36237
rect 8265 36058 8299 36203
rect 8265 36024 8358 36058
rect 8265 35832 8358 35866
rect 8265 35687 8299 35832
rect 8240 35653 8299 35687
rect 12365 35653 12393 35687
rect 8240 35413 8299 35447
rect 12365 35413 12393 35447
rect 8265 35268 8299 35413
rect 8265 35234 8358 35268
rect 8265 35042 8358 35076
rect 8265 34897 8299 35042
rect 8240 34863 8299 34897
rect 12365 34863 12393 34897
rect 8240 34623 8299 34657
rect 12365 34623 12393 34657
rect 8265 34478 8299 34623
rect 8265 34444 8358 34478
rect 8265 34252 8358 34286
rect 8265 34107 8299 34252
rect 8240 34073 8299 34107
rect 12365 34073 12393 34107
rect 8240 33833 8299 33867
rect 12365 33833 12393 33867
rect 8265 33688 8299 33833
rect 8265 33654 8358 33688
rect 8265 33462 8358 33496
rect 8265 33317 8299 33462
rect 8240 33283 8299 33317
rect 12365 33283 12393 33317
rect 8240 33043 8299 33077
rect 12365 33043 12393 33077
rect 8265 32898 8299 33043
rect 8265 32864 8358 32898
rect 8265 32672 8358 32706
rect 8265 32527 8299 32672
rect 8240 32493 8299 32527
rect 12365 32493 12393 32527
rect 8240 32253 8299 32287
rect 12365 32253 12393 32287
rect 8265 32108 8299 32253
rect 8265 32074 8358 32108
rect 8265 31882 8358 31916
rect 8265 31737 8299 31882
rect 8240 31703 8299 31737
rect 12365 31703 12393 31737
rect 8240 31463 8299 31497
rect 12365 31463 12393 31497
rect 8265 31318 8299 31463
rect 8265 31284 8358 31318
rect 8265 31092 8358 31126
rect 8265 30947 8299 31092
rect 8240 30913 8299 30947
rect 12365 30913 12393 30947
rect 8240 30673 8299 30707
rect 12365 30673 12393 30707
rect 8265 30528 8299 30673
rect 8265 30494 8358 30528
rect 8265 30302 8358 30336
rect 8265 30157 8299 30302
rect 8240 30123 8299 30157
rect 12365 30123 12393 30157
rect 8240 29883 8299 29917
rect 12365 29883 12393 29917
rect 8265 29738 8299 29883
rect 8265 29704 8358 29738
rect 8265 29512 8358 29546
rect 8265 29367 8299 29512
rect 8240 29333 8299 29367
rect 12365 29333 12393 29367
rect 8240 29093 8299 29127
rect 12365 29093 12393 29127
rect 8265 28948 8299 29093
rect 8265 28914 8358 28948
rect 8265 28722 8358 28756
rect 8265 28577 8299 28722
rect 8240 28543 8299 28577
rect 12365 28543 12393 28577
rect 8240 28303 8299 28337
rect 12365 28303 12393 28337
rect 8265 28158 8299 28303
rect 8265 28124 8358 28158
rect 8265 27932 8358 27966
rect 8265 27787 8299 27932
rect 8240 27753 8299 27787
rect 12365 27753 12393 27787
rect 8240 27513 8299 27547
rect 12365 27513 12393 27547
rect 8265 27368 8299 27513
rect 8265 27334 8358 27368
rect 8265 27142 8358 27176
rect 8265 26997 8299 27142
rect 8240 26963 8299 26997
rect 12365 26963 12393 26997
rect 8240 26723 8299 26757
rect 12365 26723 12393 26757
rect 8265 26578 8299 26723
rect 8265 26544 8358 26578
rect 8265 26352 8358 26386
rect 8265 26207 8299 26352
rect 8240 26173 8299 26207
rect 12365 26173 12393 26207
rect 8240 25933 8299 25967
rect 12365 25933 12393 25967
rect 8265 25788 8299 25933
rect 8265 25754 8358 25788
rect 8265 25562 8358 25596
rect 8265 25417 8299 25562
rect 8240 25383 8299 25417
rect 12365 25383 12393 25417
rect 8240 25143 8299 25177
rect 12365 25143 12393 25177
rect 8265 24998 8299 25143
rect 8265 24964 8358 24998
rect 8265 24772 8358 24806
rect 8265 24627 8299 24772
rect 8240 24593 8299 24627
rect 12365 24593 12393 24627
rect 8240 24353 8299 24387
rect 12365 24353 12393 24387
rect 8265 24208 8299 24353
rect 8265 24174 8358 24208
rect 8265 23982 8358 24016
rect 8265 23837 8299 23982
rect 8240 23803 8299 23837
rect 12365 23803 12393 23837
rect 8240 23563 8299 23597
rect 12365 23563 12393 23597
rect 8265 23418 8299 23563
rect 8265 23384 8358 23418
rect 8265 23192 8358 23226
rect 8265 23047 8299 23192
rect 8240 23013 8299 23047
rect 12365 23013 12393 23047
rect 8240 22773 8299 22807
rect 12365 22773 12393 22807
rect 8265 22628 8299 22773
rect 8265 22594 8358 22628
rect 8265 22402 8358 22436
rect 8265 22257 8299 22402
rect 8240 22223 8299 22257
rect 12365 22223 12393 22257
rect 8240 21983 8299 22017
rect 12365 21983 12393 22017
rect 8265 21838 8299 21983
rect 8265 21804 8358 21838
rect 8265 21612 8358 21646
rect 8265 21467 8299 21612
rect 8240 21433 8299 21467
rect 12365 21433 12393 21467
rect 8240 21193 8299 21227
rect 12365 21193 12393 21227
rect 8265 21048 8299 21193
rect 8265 21014 8358 21048
rect 8265 20822 8358 20856
rect 8265 20677 8299 20822
rect 8240 20643 8299 20677
rect 12365 20643 12393 20677
rect 8240 20403 8299 20437
rect 12365 20403 12393 20437
rect 8265 20258 8299 20403
rect 8265 20224 8358 20258
rect 8265 20032 8358 20066
rect 8265 19887 8299 20032
rect 8240 19853 8299 19887
rect 12365 19853 12393 19887
rect 8240 19613 8299 19647
rect 12365 19613 12393 19647
rect 8265 19468 8299 19613
rect 8265 19434 8358 19468
rect 8265 19242 8358 19276
rect 8265 19097 8299 19242
rect 8240 19063 8299 19097
rect 12365 19063 12393 19097
rect 8240 18823 8299 18857
rect 12365 18823 12393 18857
rect 8265 18678 8299 18823
rect 8265 18644 8358 18678
rect 8265 18452 8358 18486
rect 8265 18307 8299 18452
rect 8240 18273 8299 18307
rect 12365 18273 12393 18307
rect 8240 18033 8299 18067
rect 12365 18033 12393 18067
rect 8265 17888 8299 18033
rect 8265 17854 8358 17888
rect 8265 17662 8358 17696
rect 8265 17517 8299 17662
rect 8240 17483 8299 17517
rect 12365 17483 12393 17517
rect 8240 17243 8299 17277
rect 12365 17243 12393 17277
rect 8265 17098 8299 17243
rect 8265 17064 8358 17098
rect 8265 16872 8358 16906
rect 8265 16727 8299 16872
rect 8240 16693 8299 16727
rect 12365 16693 12393 16727
rect 8240 16453 8299 16487
rect 12365 16453 12393 16487
rect 8265 16308 8299 16453
rect 8265 16274 8358 16308
rect 8265 16082 8358 16116
rect 8265 15937 8299 16082
rect 8240 15903 8299 15937
rect 12365 15903 12393 15937
rect 8240 15663 8299 15697
rect 12365 15663 12393 15697
rect 8265 15518 8299 15663
rect 8265 15484 8358 15518
rect 8265 15292 8358 15326
rect 8265 15147 8299 15292
rect 8240 15113 8299 15147
rect 12365 15113 12393 15147
rect 8240 14873 8299 14907
rect 12365 14873 12393 14907
rect 8265 14728 8299 14873
rect 8265 14694 8358 14728
rect 8265 14502 8358 14536
rect 8265 14357 8299 14502
rect 8240 14323 8299 14357
rect 12365 14323 12393 14357
rect 8240 14083 8299 14117
rect 12365 14083 12393 14117
rect 8265 13938 8299 14083
rect 8265 13904 8358 13938
rect 8265 13712 8358 13746
rect 8265 13567 8299 13712
rect 8240 13533 8299 13567
rect 12365 13533 12393 13567
rect 8240 13293 8299 13327
rect 12365 13293 12393 13327
rect 8265 13148 8299 13293
rect 8265 13114 8358 13148
rect 8265 12922 8358 12956
rect 8265 12777 8299 12922
rect 8240 12743 8299 12777
rect 12365 12743 12393 12777
rect 8240 12503 8299 12537
rect 12365 12503 12393 12537
rect 8265 12358 8299 12503
rect 8265 12324 8358 12358
rect 8265 12132 8358 12166
rect 8265 11987 8299 12132
rect 8240 11953 8299 11987
rect 12365 11953 12393 11987
rect 8240 11713 8299 11747
rect 12365 11713 12393 11747
rect 8265 11568 8299 11713
rect 8265 11534 8358 11568
rect 8265 11342 8358 11376
rect 8265 11197 8299 11342
rect 8240 11163 8299 11197
rect 12365 11163 12393 11197
rect 8240 10923 8299 10957
rect 12365 10923 12393 10957
rect 8265 10778 8299 10923
rect 8265 10744 8358 10778
rect 8265 10552 8358 10586
rect 8265 10407 8299 10552
rect 8240 10373 8299 10407
rect 12365 10373 12393 10407
rect 8240 10133 8299 10167
rect 12365 10133 12393 10167
rect 8265 9988 8299 10133
rect 8265 9954 8358 9988
rect 8265 9762 8358 9796
rect 8265 9617 8299 9762
rect 8240 9583 8299 9617
rect 12365 9583 12393 9617
rect 8240 9343 8299 9377
rect 12365 9343 12393 9377
rect 8265 9198 8299 9343
rect 8265 9164 8358 9198
rect 8265 8972 8358 9006
rect 8265 8827 8299 8972
rect 8240 8793 8299 8827
rect 12365 8793 12393 8827
rect 8240 8553 8299 8587
rect 12365 8553 12393 8587
rect 8265 8408 8299 8553
rect 8265 8374 8358 8408
rect 8265 8182 8358 8216
rect 8265 8037 8299 8182
rect 8240 8003 8299 8037
rect 12365 8003 12393 8037
rect 8240 7763 8299 7797
rect 12365 7763 12393 7797
rect 8265 7618 8299 7763
rect 8265 7584 8358 7618
rect 8265 7392 8358 7426
rect 8265 7247 8299 7392
rect 8240 7213 8299 7247
rect 12365 7213 12393 7247
rect 8240 6973 8299 7007
rect 12365 6973 12393 7007
rect 8265 6828 8299 6973
rect 8265 6794 8358 6828
rect 8265 6602 8358 6636
rect 8265 6457 8299 6602
rect 8240 6423 8299 6457
rect 12365 6423 12393 6457
rect 8240 6183 8299 6217
rect 12365 6183 12393 6217
rect 8265 6038 8299 6183
rect 8265 6004 8358 6038
rect 8265 5812 8358 5846
rect 8265 5667 8299 5812
rect 8240 5633 8299 5667
rect 12365 5633 12393 5667
rect 8240 5393 8299 5427
rect 12365 5393 12393 5427
rect 8265 5248 8299 5393
rect 8265 5214 8358 5248
rect 8265 5022 8358 5056
rect 8265 4877 8299 5022
rect 8240 4843 8299 4877
rect 12365 4843 12393 4877
rect 8240 4603 8299 4637
rect 12365 4603 12393 4637
rect 8265 4458 8299 4603
rect 8265 4424 8358 4458
rect 8265 4232 8358 4266
rect 8265 4087 8299 4232
rect 8240 4053 8299 4087
rect 12365 4053 12393 4087
rect 8240 3813 8299 3847
rect 12365 3813 12393 3847
rect 8265 3668 8299 3813
rect 8265 3634 8358 3668
rect 8265 3442 8358 3476
rect 8265 3297 8299 3442
rect 8240 3263 8299 3297
rect 12365 3263 12393 3297
rect 8240 3023 8299 3057
rect 12365 3023 12393 3057
rect 8265 2878 8299 3023
rect 8265 2844 8358 2878
rect 8265 2652 8358 2686
rect 8265 2507 8299 2652
rect 8240 2473 8299 2507
rect 12365 2473 12393 2507
rect 8240 2233 8299 2267
rect 12365 2233 12393 2267
rect 8265 2088 8299 2233
rect 8265 2054 8358 2088
rect 8265 1862 8358 1896
rect 8265 1717 8299 1862
rect 8240 1683 8299 1717
rect 12365 1683 12393 1717
rect 8240 1443 8299 1477
rect 12365 1443 12393 1477
rect 8265 1298 8299 1443
rect 8265 1264 8358 1298
rect 8265 1072 8358 1106
rect 8265 927 8299 1072
rect 8240 893 8299 927
rect 12365 893 12393 927
rect 8240 653 8299 687
rect 12365 653 12393 687
rect 8265 508 8299 653
rect 8265 474 8358 508
rect 8265 282 8358 316
rect 8265 137 8299 282
rect 8240 103 8299 137
rect 12365 103 12393 137
<< metal1 >>
rect 8342 101393 8406 101445
rect 8102 101285 8166 101337
rect 19 0 47 9480
rect 99 0 127 9480
rect 179 0 207 9480
rect 259 0 287 9480
rect 339 0 367 9480
rect 419 0 447 9480
rect 499 0 527 9480
rect 579 0 607 9480
<< metal2 >>
rect 8106 101287 8162 101335
rect 8360 101284 8388 101433
rect 8341 101256 8388 101284
rect 8938 101281 8994 101329
rect 11629 101293 11685 101341
rect 8341 101120 8369 101256
rect 8513 50521 8569 50569
rect 8938 50520 8994 50568
rect 9981 50536 10037 50584
rect 11629 50536 11685 50584
<< metal3 >>
rect 8085 101262 8183 101360
rect 8917 101256 9015 101354
rect 11608 101268 11706 101366
rect 6425 100699 6523 100797
rect 6850 100699 6948 100797
rect 7282 100699 7380 100797
rect 7664 100676 7762 100774
rect 8060 100676 8158 100774
rect 6425 100325 6523 100423
rect 6850 100267 6948 100365
rect 7282 100267 7380 100365
rect 7664 100281 7762 100379
rect 8060 100281 8158 100379
rect 6425 99909 6523 100007
rect 6850 99909 6948 100007
rect 7282 99909 7380 100007
rect 7664 99886 7762 99984
rect 8060 99886 8158 99984
rect 6425 99535 6523 99633
rect 6850 99477 6948 99575
rect 7282 99477 7380 99575
rect 7664 99491 7762 99589
rect 8060 99491 8158 99589
rect 6425 99119 6523 99217
rect 6850 99119 6948 99217
rect 7282 99119 7380 99217
rect 7664 99096 7762 99194
rect 8060 99096 8158 99194
rect 6425 98745 6523 98843
rect 6850 98687 6948 98785
rect 7282 98687 7380 98785
rect 7664 98701 7762 98799
rect 8060 98701 8158 98799
rect 6425 98329 6523 98427
rect 6850 98329 6948 98427
rect 7282 98329 7380 98427
rect 7664 98306 7762 98404
rect 8060 98306 8158 98404
rect 6425 97955 6523 98053
rect 6850 97897 6948 97995
rect 7282 97897 7380 97995
rect 7664 97911 7762 98009
rect 8060 97911 8158 98009
rect 6425 97539 6523 97637
rect 6850 97539 6948 97637
rect 7282 97539 7380 97637
rect 7664 97516 7762 97614
rect 8060 97516 8158 97614
rect 6425 97165 6523 97263
rect 6850 97107 6948 97205
rect 7282 97107 7380 97205
rect 7664 97121 7762 97219
rect 8060 97121 8158 97219
rect 6425 96749 6523 96847
rect 6850 96749 6948 96847
rect 7282 96749 7380 96847
rect 7664 96726 7762 96824
rect 8060 96726 8158 96824
rect 6425 96375 6523 96473
rect 6850 96317 6948 96415
rect 7282 96317 7380 96415
rect 7664 96331 7762 96429
rect 8060 96331 8158 96429
rect 6425 95959 6523 96057
rect 6850 95959 6948 96057
rect 7282 95959 7380 96057
rect 7664 95936 7762 96034
rect 8060 95936 8158 96034
rect 6425 95585 6523 95683
rect 6850 95527 6948 95625
rect 7282 95527 7380 95625
rect 7664 95541 7762 95639
rect 8060 95541 8158 95639
rect 6425 95169 6523 95267
rect 6850 95169 6948 95267
rect 7282 95169 7380 95267
rect 7664 95146 7762 95244
rect 8060 95146 8158 95244
rect 6425 94795 6523 94893
rect 6850 94737 6948 94835
rect 7282 94737 7380 94835
rect 7664 94751 7762 94849
rect 8060 94751 8158 94849
rect 6425 94379 6523 94477
rect 6850 94379 6948 94477
rect 7282 94379 7380 94477
rect 7664 94356 7762 94454
rect 8060 94356 8158 94454
rect 6425 94005 6523 94103
rect 6850 93947 6948 94045
rect 7282 93947 7380 94045
rect 7664 93961 7762 94059
rect 8060 93961 8158 94059
rect 6425 93589 6523 93687
rect 6850 93589 6948 93687
rect 7282 93589 7380 93687
rect 7664 93566 7762 93664
rect 8060 93566 8158 93664
rect 6425 93215 6523 93313
rect 6850 93157 6948 93255
rect 7282 93157 7380 93255
rect 7664 93171 7762 93269
rect 8060 93171 8158 93269
rect 6425 92799 6523 92897
rect 6850 92799 6948 92897
rect 7282 92799 7380 92897
rect 7664 92776 7762 92874
rect 8060 92776 8158 92874
rect 6425 92425 6523 92523
rect 6850 92367 6948 92465
rect 7282 92367 7380 92465
rect 7664 92381 7762 92479
rect 8060 92381 8158 92479
rect 6425 92009 6523 92107
rect 6850 92009 6948 92107
rect 7282 92009 7380 92107
rect 7664 91986 7762 92084
rect 8060 91986 8158 92084
rect 6425 91635 6523 91733
rect 6850 91577 6948 91675
rect 7282 91577 7380 91675
rect 7664 91591 7762 91689
rect 8060 91591 8158 91689
rect 6425 91219 6523 91317
rect 6850 91219 6948 91317
rect 7282 91219 7380 91317
rect 7664 91196 7762 91294
rect 8060 91196 8158 91294
rect 6425 90845 6523 90943
rect 6850 90787 6948 90885
rect 7282 90787 7380 90885
rect 7664 90801 7762 90899
rect 8060 90801 8158 90899
rect 6425 90429 6523 90527
rect 6850 90429 6948 90527
rect 7282 90429 7380 90527
rect 7664 90406 7762 90504
rect 8060 90406 8158 90504
rect 6425 90055 6523 90153
rect 6850 89997 6948 90095
rect 7282 89997 7380 90095
rect 7664 90011 7762 90109
rect 8060 90011 8158 90109
rect 6425 89639 6523 89737
rect 6850 89639 6948 89737
rect 7282 89639 7380 89737
rect 7664 89616 7762 89714
rect 8060 89616 8158 89714
rect 6425 89265 6523 89363
rect 6850 89207 6948 89305
rect 7282 89207 7380 89305
rect 7664 89221 7762 89319
rect 8060 89221 8158 89319
rect 6425 88849 6523 88947
rect 6850 88849 6948 88947
rect 7282 88849 7380 88947
rect 7664 88826 7762 88924
rect 8060 88826 8158 88924
rect 6425 88475 6523 88573
rect 6850 88417 6948 88515
rect 7282 88417 7380 88515
rect 7664 88431 7762 88529
rect 8060 88431 8158 88529
rect 6425 88059 6523 88157
rect 6850 88059 6948 88157
rect 7282 88059 7380 88157
rect 7664 88036 7762 88134
rect 8060 88036 8158 88134
rect 6425 87685 6523 87783
rect 6850 87627 6948 87725
rect 7282 87627 7380 87725
rect 7664 87641 7762 87739
rect 8060 87641 8158 87739
rect 6425 87269 6523 87367
rect 6850 87269 6948 87367
rect 7282 87269 7380 87367
rect 7664 87246 7762 87344
rect 8060 87246 8158 87344
rect 6425 86895 6523 86993
rect 6850 86837 6948 86935
rect 7282 86837 7380 86935
rect 7664 86851 7762 86949
rect 8060 86851 8158 86949
rect 6425 86479 6523 86577
rect 6850 86479 6948 86577
rect 7282 86479 7380 86577
rect 7664 86456 7762 86554
rect 8060 86456 8158 86554
rect 6425 86105 6523 86203
rect 6850 86047 6948 86145
rect 7282 86047 7380 86145
rect 7664 86061 7762 86159
rect 8060 86061 8158 86159
rect 6425 85689 6523 85787
rect 6850 85689 6948 85787
rect 7282 85689 7380 85787
rect 7664 85666 7762 85764
rect 8060 85666 8158 85764
rect 6425 85315 6523 85413
rect 6850 85257 6948 85355
rect 7282 85257 7380 85355
rect 7664 85271 7762 85369
rect 8060 85271 8158 85369
rect 6425 84899 6523 84997
rect 6850 84899 6948 84997
rect 7282 84899 7380 84997
rect 7664 84876 7762 84974
rect 8060 84876 8158 84974
rect 6425 84525 6523 84623
rect 6850 84467 6948 84565
rect 7282 84467 7380 84565
rect 7664 84481 7762 84579
rect 8060 84481 8158 84579
rect 6425 84109 6523 84207
rect 6850 84109 6948 84207
rect 7282 84109 7380 84207
rect 7664 84086 7762 84184
rect 8060 84086 8158 84184
rect 6425 83735 6523 83833
rect 6850 83677 6948 83775
rect 7282 83677 7380 83775
rect 7664 83691 7762 83789
rect 8060 83691 8158 83789
rect 6425 83319 6523 83417
rect 6850 83319 6948 83417
rect 7282 83319 7380 83417
rect 7664 83296 7762 83394
rect 8060 83296 8158 83394
rect 6425 82945 6523 83043
rect 6850 82887 6948 82985
rect 7282 82887 7380 82985
rect 7664 82901 7762 82999
rect 8060 82901 8158 82999
rect 6425 82529 6523 82627
rect 6850 82529 6948 82627
rect 7282 82529 7380 82627
rect 7664 82506 7762 82604
rect 8060 82506 8158 82604
rect 6425 82155 6523 82253
rect 6850 82097 6948 82195
rect 7282 82097 7380 82195
rect 7664 82111 7762 82209
rect 8060 82111 8158 82209
rect 6425 81739 6523 81837
rect 6850 81739 6948 81837
rect 7282 81739 7380 81837
rect 7664 81716 7762 81814
rect 8060 81716 8158 81814
rect 6425 81365 6523 81463
rect 6850 81307 6948 81405
rect 7282 81307 7380 81405
rect 7664 81321 7762 81419
rect 8060 81321 8158 81419
rect 6425 80949 6523 81047
rect 6850 80949 6948 81047
rect 7282 80949 7380 81047
rect 7664 80926 7762 81024
rect 8060 80926 8158 81024
rect 6425 80575 6523 80673
rect 6850 80517 6948 80615
rect 7282 80517 7380 80615
rect 7664 80531 7762 80629
rect 8060 80531 8158 80629
rect 6425 80159 6523 80257
rect 6850 80159 6948 80257
rect 7282 80159 7380 80257
rect 7664 80136 7762 80234
rect 8060 80136 8158 80234
rect 6425 79785 6523 79883
rect 6850 79727 6948 79825
rect 7282 79727 7380 79825
rect 7664 79741 7762 79839
rect 8060 79741 8158 79839
rect 6425 79369 6523 79467
rect 6850 79369 6948 79467
rect 7282 79369 7380 79467
rect 7664 79346 7762 79444
rect 8060 79346 8158 79444
rect 6425 78995 6523 79093
rect 6850 78937 6948 79035
rect 7282 78937 7380 79035
rect 7664 78951 7762 79049
rect 8060 78951 8158 79049
rect 6425 78579 6523 78677
rect 6850 78579 6948 78677
rect 7282 78579 7380 78677
rect 7664 78556 7762 78654
rect 8060 78556 8158 78654
rect 6425 78205 6523 78303
rect 6850 78147 6948 78245
rect 7282 78147 7380 78245
rect 7664 78161 7762 78259
rect 8060 78161 8158 78259
rect 6425 77789 6523 77887
rect 6850 77789 6948 77887
rect 7282 77789 7380 77887
rect 7664 77766 7762 77864
rect 8060 77766 8158 77864
rect 6425 77415 6523 77513
rect 6850 77357 6948 77455
rect 7282 77357 7380 77455
rect 7664 77371 7762 77469
rect 8060 77371 8158 77469
rect 6425 76999 6523 77097
rect 6850 76999 6948 77097
rect 7282 76999 7380 77097
rect 7664 76976 7762 77074
rect 8060 76976 8158 77074
rect 6425 76625 6523 76723
rect 6850 76567 6948 76665
rect 7282 76567 7380 76665
rect 7664 76581 7762 76679
rect 8060 76581 8158 76679
rect 6425 76209 6523 76307
rect 6850 76209 6948 76307
rect 7282 76209 7380 76307
rect 7664 76186 7762 76284
rect 8060 76186 8158 76284
rect 6425 75835 6523 75933
rect 6850 75777 6948 75875
rect 7282 75777 7380 75875
rect 7664 75791 7762 75889
rect 8060 75791 8158 75889
rect 6425 75419 6523 75517
rect 6850 75419 6948 75517
rect 7282 75419 7380 75517
rect 7664 75396 7762 75494
rect 8060 75396 8158 75494
rect 6425 75045 6523 75143
rect 6850 74987 6948 75085
rect 7282 74987 7380 75085
rect 7664 75001 7762 75099
rect 8060 75001 8158 75099
rect 6425 74629 6523 74727
rect 6850 74629 6948 74727
rect 7282 74629 7380 74727
rect 7664 74606 7762 74704
rect 8060 74606 8158 74704
rect 6425 74255 6523 74353
rect 6850 74197 6948 74295
rect 7282 74197 7380 74295
rect 7664 74211 7762 74309
rect 8060 74211 8158 74309
rect 6425 73839 6523 73937
rect 6850 73839 6948 73937
rect 7282 73839 7380 73937
rect 7664 73816 7762 73914
rect 8060 73816 8158 73914
rect 6425 73465 6523 73563
rect 6850 73407 6948 73505
rect 7282 73407 7380 73505
rect 7664 73421 7762 73519
rect 8060 73421 8158 73519
rect 6425 73049 6523 73147
rect 6850 73049 6948 73147
rect 7282 73049 7380 73147
rect 7664 73026 7762 73124
rect 8060 73026 8158 73124
rect 6425 72675 6523 72773
rect 6850 72617 6948 72715
rect 7282 72617 7380 72715
rect 7664 72631 7762 72729
rect 8060 72631 8158 72729
rect 6425 72259 6523 72357
rect 6850 72259 6948 72357
rect 7282 72259 7380 72357
rect 7664 72236 7762 72334
rect 8060 72236 8158 72334
rect 6425 71885 6523 71983
rect 6850 71827 6948 71925
rect 7282 71827 7380 71925
rect 7664 71841 7762 71939
rect 8060 71841 8158 71939
rect 6425 71469 6523 71567
rect 6850 71469 6948 71567
rect 7282 71469 7380 71567
rect 7664 71446 7762 71544
rect 8060 71446 8158 71544
rect 6425 71095 6523 71193
rect 6850 71037 6948 71135
rect 7282 71037 7380 71135
rect 7664 71051 7762 71149
rect 8060 71051 8158 71149
rect 6425 70679 6523 70777
rect 6850 70679 6948 70777
rect 7282 70679 7380 70777
rect 7664 70656 7762 70754
rect 8060 70656 8158 70754
rect 6425 70305 6523 70403
rect 6850 70247 6948 70345
rect 7282 70247 7380 70345
rect 7664 70261 7762 70359
rect 8060 70261 8158 70359
rect 6425 69889 6523 69987
rect 6850 69889 6948 69987
rect 7282 69889 7380 69987
rect 7664 69866 7762 69964
rect 8060 69866 8158 69964
rect 6425 69515 6523 69613
rect 6850 69457 6948 69555
rect 7282 69457 7380 69555
rect 7664 69471 7762 69569
rect 8060 69471 8158 69569
rect 6425 69099 6523 69197
rect 6850 69099 6948 69197
rect 7282 69099 7380 69197
rect 7664 69076 7762 69174
rect 8060 69076 8158 69174
rect 6425 68725 6523 68823
rect 6850 68667 6948 68765
rect 7282 68667 7380 68765
rect 7664 68681 7762 68779
rect 8060 68681 8158 68779
rect 6425 68309 6523 68407
rect 6850 68309 6948 68407
rect 7282 68309 7380 68407
rect 7664 68286 7762 68384
rect 8060 68286 8158 68384
rect 6425 67935 6523 68033
rect 6850 67877 6948 67975
rect 7282 67877 7380 67975
rect 7664 67891 7762 67989
rect 8060 67891 8158 67989
rect 6425 67519 6523 67617
rect 6850 67519 6948 67617
rect 7282 67519 7380 67617
rect 7664 67496 7762 67594
rect 8060 67496 8158 67594
rect 6425 67145 6523 67243
rect 6850 67087 6948 67185
rect 7282 67087 7380 67185
rect 7664 67101 7762 67199
rect 8060 67101 8158 67199
rect 6425 66729 6523 66827
rect 6850 66729 6948 66827
rect 7282 66729 7380 66827
rect 7664 66706 7762 66804
rect 8060 66706 8158 66804
rect 6425 66355 6523 66453
rect 6850 66297 6948 66395
rect 7282 66297 7380 66395
rect 7664 66311 7762 66409
rect 8060 66311 8158 66409
rect 6425 65939 6523 66037
rect 6850 65939 6948 66037
rect 7282 65939 7380 66037
rect 7664 65916 7762 66014
rect 8060 65916 8158 66014
rect 6425 65565 6523 65663
rect 6850 65507 6948 65605
rect 7282 65507 7380 65605
rect 7664 65521 7762 65619
rect 8060 65521 8158 65619
rect 6425 65149 6523 65247
rect 6850 65149 6948 65247
rect 7282 65149 7380 65247
rect 7664 65126 7762 65224
rect 8060 65126 8158 65224
rect 6425 64775 6523 64873
rect 6850 64717 6948 64815
rect 7282 64717 7380 64815
rect 7664 64731 7762 64829
rect 8060 64731 8158 64829
rect 6425 64359 6523 64457
rect 6850 64359 6948 64457
rect 7282 64359 7380 64457
rect 7664 64336 7762 64434
rect 8060 64336 8158 64434
rect 6425 63985 6523 64083
rect 6850 63927 6948 64025
rect 7282 63927 7380 64025
rect 7664 63941 7762 64039
rect 8060 63941 8158 64039
rect 6425 63569 6523 63667
rect 6850 63569 6948 63667
rect 7282 63569 7380 63667
rect 7664 63546 7762 63644
rect 8060 63546 8158 63644
rect 6425 63195 6523 63293
rect 6850 63137 6948 63235
rect 7282 63137 7380 63235
rect 7664 63151 7762 63249
rect 8060 63151 8158 63249
rect 6425 62779 6523 62877
rect 6850 62779 6948 62877
rect 7282 62779 7380 62877
rect 7664 62756 7762 62854
rect 8060 62756 8158 62854
rect 6425 62405 6523 62503
rect 6850 62347 6948 62445
rect 7282 62347 7380 62445
rect 7664 62361 7762 62459
rect 8060 62361 8158 62459
rect 6425 61989 6523 62087
rect 6850 61989 6948 62087
rect 7282 61989 7380 62087
rect 7664 61966 7762 62064
rect 8060 61966 8158 62064
rect 6425 61615 6523 61713
rect 6850 61557 6948 61655
rect 7282 61557 7380 61655
rect 7664 61571 7762 61669
rect 8060 61571 8158 61669
rect 6425 61199 6523 61297
rect 6850 61199 6948 61297
rect 7282 61199 7380 61297
rect 7664 61176 7762 61274
rect 8060 61176 8158 61274
rect 6425 60825 6523 60923
rect 6850 60767 6948 60865
rect 7282 60767 7380 60865
rect 7664 60781 7762 60879
rect 8060 60781 8158 60879
rect 6425 60409 6523 60507
rect 6850 60409 6948 60507
rect 7282 60409 7380 60507
rect 7664 60386 7762 60484
rect 8060 60386 8158 60484
rect 6425 60035 6523 60133
rect 6850 59977 6948 60075
rect 7282 59977 7380 60075
rect 7664 59991 7762 60089
rect 8060 59991 8158 60089
rect 6425 59619 6523 59717
rect 6850 59619 6948 59717
rect 7282 59619 7380 59717
rect 7664 59596 7762 59694
rect 8060 59596 8158 59694
rect 6425 59245 6523 59343
rect 6850 59187 6948 59285
rect 7282 59187 7380 59285
rect 7664 59201 7762 59299
rect 8060 59201 8158 59299
rect 6425 58829 6523 58927
rect 6850 58829 6948 58927
rect 7282 58829 7380 58927
rect 7664 58806 7762 58904
rect 8060 58806 8158 58904
rect 6425 58455 6523 58553
rect 6850 58397 6948 58495
rect 7282 58397 7380 58495
rect 7664 58411 7762 58509
rect 8060 58411 8158 58509
rect 6425 58039 6523 58137
rect 6850 58039 6948 58137
rect 7282 58039 7380 58137
rect 7664 58016 7762 58114
rect 8060 58016 8158 58114
rect 6425 57665 6523 57763
rect 6850 57607 6948 57705
rect 7282 57607 7380 57705
rect 7664 57621 7762 57719
rect 8060 57621 8158 57719
rect 6425 57249 6523 57347
rect 6850 57249 6948 57347
rect 7282 57249 7380 57347
rect 7664 57226 7762 57324
rect 8060 57226 8158 57324
rect 6425 56875 6523 56973
rect 6850 56817 6948 56915
rect 7282 56817 7380 56915
rect 7664 56831 7762 56929
rect 8060 56831 8158 56929
rect 6425 56459 6523 56557
rect 6850 56459 6948 56557
rect 7282 56459 7380 56557
rect 7664 56436 7762 56534
rect 8060 56436 8158 56534
rect 6425 56085 6523 56183
rect 6850 56027 6948 56125
rect 7282 56027 7380 56125
rect 7664 56041 7762 56139
rect 8060 56041 8158 56139
rect 6425 55669 6523 55767
rect 6850 55669 6948 55767
rect 7282 55669 7380 55767
rect 7664 55646 7762 55744
rect 8060 55646 8158 55744
rect 6425 55295 6523 55393
rect 6850 55237 6948 55335
rect 7282 55237 7380 55335
rect 7664 55251 7762 55349
rect 8060 55251 8158 55349
rect 6425 54879 6523 54977
rect 6850 54879 6948 54977
rect 7282 54879 7380 54977
rect 7664 54856 7762 54954
rect 8060 54856 8158 54954
rect 6425 54505 6523 54603
rect 6850 54447 6948 54545
rect 7282 54447 7380 54545
rect 7664 54461 7762 54559
rect 8060 54461 8158 54559
rect 6425 54089 6523 54187
rect 6850 54089 6948 54187
rect 7282 54089 7380 54187
rect 7664 54066 7762 54164
rect 8060 54066 8158 54164
rect 6425 53715 6523 53813
rect 6850 53657 6948 53755
rect 7282 53657 7380 53755
rect 7664 53671 7762 53769
rect 8060 53671 8158 53769
rect 6425 53299 6523 53397
rect 6850 53299 6948 53397
rect 7282 53299 7380 53397
rect 7664 53276 7762 53374
rect 8060 53276 8158 53374
rect 6425 52925 6523 53023
rect 6850 52867 6948 52965
rect 7282 52867 7380 52965
rect 7664 52881 7762 52979
rect 8060 52881 8158 52979
rect 6425 52509 6523 52607
rect 6850 52509 6948 52607
rect 7282 52509 7380 52607
rect 7664 52486 7762 52584
rect 8060 52486 8158 52584
rect 6425 52135 6523 52233
rect 6850 52077 6948 52175
rect 7282 52077 7380 52175
rect 7664 52091 7762 52189
rect 8060 52091 8158 52189
rect 6425 51719 6523 51817
rect 6850 51719 6948 51817
rect 7282 51719 7380 51817
rect 7664 51696 7762 51794
rect 8060 51696 8158 51794
rect 6425 51345 6523 51443
rect 6850 51287 6948 51385
rect 7282 51287 7380 51385
rect 7664 51301 7762 51399
rect 8060 51301 8158 51399
rect 6425 50929 6523 51027
rect 6850 50929 6948 51027
rect 7282 50929 7380 51027
rect 7664 50906 7762 51004
rect 8060 50906 8158 51004
rect 6425 50555 6523 50653
rect 6850 50497 6948 50595
rect 7282 50497 7380 50595
rect 7664 50511 7762 50609
rect 8060 50511 8158 50609
rect 8492 50496 8590 50594
rect 8917 50495 9015 50593
rect 9960 50511 10058 50609
rect 11608 50511 11706 50609
rect 6425 50139 6523 50237
rect 6850 50139 6948 50237
rect 7282 50139 7380 50237
rect 7664 50116 7762 50214
rect 8060 50116 8158 50214
rect 6425 49765 6523 49863
rect 6850 49707 6948 49805
rect 7282 49707 7380 49805
rect 7664 49721 7762 49819
rect 8060 49721 8158 49819
rect 6425 49349 6523 49447
rect 6850 49349 6948 49447
rect 7282 49349 7380 49447
rect 7664 49326 7762 49424
rect 8060 49326 8158 49424
rect 6425 48975 6523 49073
rect 6850 48917 6948 49015
rect 7282 48917 7380 49015
rect 7664 48931 7762 49029
rect 8060 48931 8158 49029
rect 6425 48559 6523 48657
rect 6850 48559 6948 48657
rect 7282 48559 7380 48657
rect 7664 48536 7762 48634
rect 8060 48536 8158 48634
rect 6425 48185 6523 48283
rect 6850 48127 6948 48225
rect 7282 48127 7380 48225
rect 7664 48141 7762 48239
rect 8060 48141 8158 48239
rect 6425 47769 6523 47867
rect 6850 47769 6948 47867
rect 7282 47769 7380 47867
rect 7664 47746 7762 47844
rect 8060 47746 8158 47844
rect 6425 47395 6523 47493
rect 6850 47337 6948 47435
rect 7282 47337 7380 47435
rect 7664 47351 7762 47449
rect 8060 47351 8158 47449
rect 6425 46979 6523 47077
rect 6850 46979 6948 47077
rect 7282 46979 7380 47077
rect 7664 46956 7762 47054
rect 8060 46956 8158 47054
rect 6425 46605 6523 46703
rect 6850 46547 6948 46645
rect 7282 46547 7380 46645
rect 7664 46561 7762 46659
rect 8060 46561 8158 46659
rect 6425 46189 6523 46287
rect 6850 46189 6948 46287
rect 7282 46189 7380 46287
rect 7664 46166 7762 46264
rect 8060 46166 8158 46264
rect 6425 45815 6523 45913
rect 6850 45757 6948 45855
rect 7282 45757 7380 45855
rect 7664 45771 7762 45869
rect 8060 45771 8158 45869
rect 6425 45399 6523 45497
rect 6850 45399 6948 45497
rect 7282 45399 7380 45497
rect 7664 45376 7762 45474
rect 8060 45376 8158 45474
rect 6425 45025 6523 45123
rect 6850 44967 6948 45065
rect 7282 44967 7380 45065
rect 7664 44981 7762 45079
rect 8060 44981 8158 45079
rect 6425 44609 6523 44707
rect 6850 44609 6948 44707
rect 7282 44609 7380 44707
rect 7664 44586 7762 44684
rect 8060 44586 8158 44684
rect 6425 44235 6523 44333
rect 6850 44177 6948 44275
rect 7282 44177 7380 44275
rect 7664 44191 7762 44289
rect 8060 44191 8158 44289
rect 6425 43819 6523 43917
rect 6850 43819 6948 43917
rect 7282 43819 7380 43917
rect 7664 43796 7762 43894
rect 8060 43796 8158 43894
rect 6425 43445 6523 43543
rect 6850 43387 6948 43485
rect 7282 43387 7380 43485
rect 7664 43401 7762 43499
rect 8060 43401 8158 43499
rect 6425 43029 6523 43127
rect 6850 43029 6948 43127
rect 7282 43029 7380 43127
rect 7664 43006 7762 43104
rect 8060 43006 8158 43104
rect 6425 42655 6523 42753
rect 6850 42597 6948 42695
rect 7282 42597 7380 42695
rect 7664 42611 7762 42709
rect 8060 42611 8158 42709
rect 6425 42239 6523 42337
rect 6850 42239 6948 42337
rect 7282 42239 7380 42337
rect 7664 42216 7762 42314
rect 8060 42216 8158 42314
rect 6425 41865 6523 41963
rect 6850 41807 6948 41905
rect 7282 41807 7380 41905
rect 7664 41821 7762 41919
rect 8060 41821 8158 41919
rect 6425 41449 6523 41547
rect 6850 41449 6948 41547
rect 7282 41449 7380 41547
rect 7664 41426 7762 41524
rect 8060 41426 8158 41524
rect 6425 41075 6523 41173
rect 6850 41017 6948 41115
rect 7282 41017 7380 41115
rect 7664 41031 7762 41129
rect 8060 41031 8158 41129
rect 6425 40659 6523 40757
rect 6850 40659 6948 40757
rect 7282 40659 7380 40757
rect 7664 40636 7762 40734
rect 8060 40636 8158 40734
rect 6425 40285 6523 40383
rect 6850 40227 6948 40325
rect 7282 40227 7380 40325
rect 7664 40241 7762 40339
rect 8060 40241 8158 40339
rect 6425 39869 6523 39967
rect 6850 39869 6948 39967
rect 7282 39869 7380 39967
rect 7664 39846 7762 39944
rect 8060 39846 8158 39944
rect 6425 39495 6523 39593
rect 6850 39437 6948 39535
rect 7282 39437 7380 39535
rect 7664 39451 7762 39549
rect 8060 39451 8158 39549
rect 6425 39079 6523 39177
rect 6850 39079 6948 39177
rect 7282 39079 7380 39177
rect 7664 39056 7762 39154
rect 8060 39056 8158 39154
rect 6425 38705 6523 38803
rect 6850 38647 6948 38745
rect 7282 38647 7380 38745
rect 7664 38661 7762 38759
rect 8060 38661 8158 38759
rect 6425 38289 6523 38387
rect 6850 38289 6948 38387
rect 7282 38289 7380 38387
rect 7664 38266 7762 38364
rect 8060 38266 8158 38364
rect 6425 37915 6523 38013
rect 6850 37857 6948 37955
rect 7282 37857 7380 37955
rect 7664 37871 7762 37969
rect 8060 37871 8158 37969
rect 6425 37499 6523 37597
rect 6850 37499 6948 37597
rect 7282 37499 7380 37597
rect 7664 37476 7762 37574
rect 8060 37476 8158 37574
rect 6425 37125 6523 37223
rect 6850 37067 6948 37165
rect 7282 37067 7380 37165
rect 7664 37081 7762 37179
rect 8060 37081 8158 37179
rect 6425 36709 6523 36807
rect 6850 36709 6948 36807
rect 7282 36709 7380 36807
rect 7664 36686 7762 36784
rect 8060 36686 8158 36784
rect 6425 36335 6523 36433
rect 6850 36277 6948 36375
rect 7282 36277 7380 36375
rect 7664 36291 7762 36389
rect 8060 36291 8158 36389
rect 6425 35919 6523 36017
rect 6850 35919 6948 36017
rect 7282 35919 7380 36017
rect 7664 35896 7762 35994
rect 8060 35896 8158 35994
rect 6425 35545 6523 35643
rect 6850 35487 6948 35585
rect 7282 35487 7380 35585
rect 7664 35501 7762 35599
rect 8060 35501 8158 35599
rect 6425 35129 6523 35227
rect 6850 35129 6948 35227
rect 7282 35129 7380 35227
rect 7664 35106 7762 35204
rect 8060 35106 8158 35204
rect 6425 34755 6523 34853
rect 6850 34697 6948 34795
rect 7282 34697 7380 34795
rect 7664 34711 7762 34809
rect 8060 34711 8158 34809
rect 6425 34339 6523 34437
rect 6850 34339 6948 34437
rect 7282 34339 7380 34437
rect 7664 34316 7762 34414
rect 8060 34316 8158 34414
rect 6425 33965 6523 34063
rect 6850 33907 6948 34005
rect 7282 33907 7380 34005
rect 7664 33921 7762 34019
rect 8060 33921 8158 34019
rect 6425 33549 6523 33647
rect 6850 33549 6948 33647
rect 7282 33549 7380 33647
rect 7664 33526 7762 33624
rect 8060 33526 8158 33624
rect 6425 33175 6523 33273
rect 6850 33117 6948 33215
rect 7282 33117 7380 33215
rect 7664 33131 7762 33229
rect 8060 33131 8158 33229
rect 6425 32759 6523 32857
rect 6850 32759 6948 32857
rect 7282 32759 7380 32857
rect 7664 32736 7762 32834
rect 8060 32736 8158 32834
rect 6425 32385 6523 32483
rect 6850 32327 6948 32425
rect 7282 32327 7380 32425
rect 7664 32341 7762 32439
rect 8060 32341 8158 32439
rect 6425 31969 6523 32067
rect 6850 31969 6948 32067
rect 7282 31969 7380 32067
rect 7664 31946 7762 32044
rect 8060 31946 8158 32044
rect 6425 31595 6523 31693
rect 6850 31537 6948 31635
rect 7282 31537 7380 31635
rect 7664 31551 7762 31649
rect 8060 31551 8158 31649
rect 6425 31179 6523 31277
rect 6850 31179 6948 31277
rect 7282 31179 7380 31277
rect 7664 31156 7762 31254
rect 8060 31156 8158 31254
rect 6425 30805 6523 30903
rect 6850 30747 6948 30845
rect 7282 30747 7380 30845
rect 7664 30761 7762 30859
rect 8060 30761 8158 30859
rect 6425 30389 6523 30487
rect 6850 30389 6948 30487
rect 7282 30389 7380 30487
rect 7664 30366 7762 30464
rect 8060 30366 8158 30464
rect 6425 30015 6523 30113
rect 6850 29957 6948 30055
rect 7282 29957 7380 30055
rect 7664 29971 7762 30069
rect 8060 29971 8158 30069
rect 6425 29599 6523 29697
rect 6850 29599 6948 29697
rect 7282 29599 7380 29697
rect 7664 29576 7762 29674
rect 8060 29576 8158 29674
rect 6425 29225 6523 29323
rect 6850 29167 6948 29265
rect 7282 29167 7380 29265
rect 7664 29181 7762 29279
rect 8060 29181 8158 29279
rect 6425 28809 6523 28907
rect 6850 28809 6948 28907
rect 7282 28809 7380 28907
rect 7664 28786 7762 28884
rect 8060 28786 8158 28884
rect 6425 28435 6523 28533
rect 6850 28377 6948 28475
rect 7282 28377 7380 28475
rect 7664 28391 7762 28489
rect 8060 28391 8158 28489
rect 6425 28019 6523 28117
rect 6850 28019 6948 28117
rect 7282 28019 7380 28117
rect 7664 27996 7762 28094
rect 8060 27996 8158 28094
rect 6425 27645 6523 27743
rect 6850 27587 6948 27685
rect 7282 27587 7380 27685
rect 7664 27601 7762 27699
rect 8060 27601 8158 27699
rect 6425 27229 6523 27327
rect 6850 27229 6948 27327
rect 7282 27229 7380 27327
rect 7664 27206 7762 27304
rect 8060 27206 8158 27304
rect 6425 26855 6523 26953
rect 6850 26797 6948 26895
rect 7282 26797 7380 26895
rect 7664 26811 7762 26909
rect 8060 26811 8158 26909
rect 6425 26439 6523 26537
rect 6850 26439 6948 26537
rect 7282 26439 7380 26537
rect 7664 26416 7762 26514
rect 8060 26416 8158 26514
rect 6425 26065 6523 26163
rect 6850 26007 6948 26105
rect 7282 26007 7380 26105
rect 7664 26021 7762 26119
rect 8060 26021 8158 26119
rect 6425 25649 6523 25747
rect 6850 25649 6948 25747
rect 7282 25649 7380 25747
rect 7664 25626 7762 25724
rect 8060 25626 8158 25724
rect 6425 25275 6523 25373
rect 6850 25217 6948 25315
rect 7282 25217 7380 25315
rect 7664 25231 7762 25329
rect 8060 25231 8158 25329
rect 6425 24859 6523 24957
rect 6850 24859 6948 24957
rect 7282 24859 7380 24957
rect 7664 24836 7762 24934
rect 8060 24836 8158 24934
rect 6425 24485 6523 24583
rect 6850 24427 6948 24525
rect 7282 24427 7380 24525
rect 7664 24441 7762 24539
rect 8060 24441 8158 24539
rect 6425 24069 6523 24167
rect 6850 24069 6948 24167
rect 7282 24069 7380 24167
rect 7664 24046 7762 24144
rect 8060 24046 8158 24144
rect 6425 23695 6523 23793
rect 6850 23637 6948 23735
rect 7282 23637 7380 23735
rect 7664 23651 7762 23749
rect 8060 23651 8158 23749
rect 6425 23279 6523 23377
rect 6850 23279 6948 23377
rect 7282 23279 7380 23377
rect 7664 23256 7762 23354
rect 8060 23256 8158 23354
rect 6425 22905 6523 23003
rect 6850 22847 6948 22945
rect 7282 22847 7380 22945
rect 7664 22861 7762 22959
rect 8060 22861 8158 22959
rect 6425 22489 6523 22587
rect 6850 22489 6948 22587
rect 7282 22489 7380 22587
rect 7664 22466 7762 22564
rect 8060 22466 8158 22564
rect 6425 22115 6523 22213
rect 6850 22057 6948 22155
rect 7282 22057 7380 22155
rect 7664 22071 7762 22169
rect 8060 22071 8158 22169
rect 6425 21699 6523 21797
rect 6850 21699 6948 21797
rect 7282 21699 7380 21797
rect 7664 21676 7762 21774
rect 8060 21676 8158 21774
rect 6425 21325 6523 21423
rect 6850 21267 6948 21365
rect 7282 21267 7380 21365
rect 7664 21281 7762 21379
rect 8060 21281 8158 21379
rect 6425 20909 6523 21007
rect 6850 20909 6948 21007
rect 7282 20909 7380 21007
rect 7664 20886 7762 20984
rect 8060 20886 8158 20984
rect 6425 20535 6523 20633
rect 6850 20477 6948 20575
rect 7282 20477 7380 20575
rect 7664 20491 7762 20589
rect 8060 20491 8158 20589
rect 6425 20119 6523 20217
rect 6850 20119 6948 20217
rect 7282 20119 7380 20217
rect 7664 20096 7762 20194
rect 8060 20096 8158 20194
rect 6425 19745 6523 19843
rect 6850 19687 6948 19785
rect 7282 19687 7380 19785
rect 7664 19701 7762 19799
rect 8060 19701 8158 19799
rect 6425 19329 6523 19427
rect 6850 19329 6948 19427
rect 7282 19329 7380 19427
rect 7664 19306 7762 19404
rect 8060 19306 8158 19404
rect 6425 18955 6523 19053
rect 6850 18897 6948 18995
rect 7282 18897 7380 18995
rect 7664 18911 7762 19009
rect 8060 18911 8158 19009
rect 6425 18539 6523 18637
rect 6850 18539 6948 18637
rect 7282 18539 7380 18637
rect 7664 18516 7762 18614
rect 8060 18516 8158 18614
rect 6425 18165 6523 18263
rect 6850 18107 6948 18205
rect 7282 18107 7380 18205
rect 7664 18121 7762 18219
rect 8060 18121 8158 18219
rect 6425 17749 6523 17847
rect 6850 17749 6948 17847
rect 7282 17749 7380 17847
rect 7664 17726 7762 17824
rect 8060 17726 8158 17824
rect 6425 17375 6523 17473
rect 6850 17317 6948 17415
rect 7282 17317 7380 17415
rect 7664 17331 7762 17429
rect 8060 17331 8158 17429
rect 6425 16959 6523 17057
rect 6850 16959 6948 17057
rect 7282 16959 7380 17057
rect 7664 16936 7762 17034
rect 8060 16936 8158 17034
rect 6425 16585 6523 16683
rect 6850 16527 6948 16625
rect 7282 16527 7380 16625
rect 7664 16541 7762 16639
rect 8060 16541 8158 16639
rect 6425 16169 6523 16267
rect 6850 16169 6948 16267
rect 7282 16169 7380 16267
rect 7664 16146 7762 16244
rect 8060 16146 8158 16244
rect 6425 15795 6523 15893
rect 6850 15737 6948 15835
rect 7282 15737 7380 15835
rect 7664 15751 7762 15849
rect 8060 15751 8158 15849
rect 6425 15379 6523 15477
rect 6850 15379 6948 15477
rect 7282 15379 7380 15477
rect 7664 15356 7762 15454
rect 8060 15356 8158 15454
rect 6425 15005 6523 15103
rect 6850 14947 6948 15045
rect 7282 14947 7380 15045
rect 7664 14961 7762 15059
rect 8060 14961 8158 15059
rect 6425 14589 6523 14687
rect 6850 14589 6948 14687
rect 7282 14589 7380 14687
rect 7664 14566 7762 14664
rect 8060 14566 8158 14664
rect 6425 14215 6523 14313
rect 6850 14157 6948 14255
rect 7282 14157 7380 14255
rect 7664 14171 7762 14269
rect 8060 14171 8158 14269
rect 6425 13799 6523 13897
rect 6850 13799 6948 13897
rect 7282 13799 7380 13897
rect 7664 13776 7762 13874
rect 8060 13776 8158 13874
rect 6425 13425 6523 13523
rect 6850 13367 6948 13465
rect 7282 13367 7380 13465
rect 7664 13381 7762 13479
rect 8060 13381 8158 13479
rect 6425 13009 6523 13107
rect 6850 13009 6948 13107
rect 7282 13009 7380 13107
rect 7664 12986 7762 13084
rect 8060 12986 8158 13084
rect 6425 12635 6523 12733
rect 6850 12577 6948 12675
rect 7282 12577 7380 12675
rect 7664 12591 7762 12689
rect 8060 12591 8158 12689
rect 6425 12219 6523 12317
rect 6850 12219 6948 12317
rect 7282 12219 7380 12317
rect 7664 12196 7762 12294
rect 8060 12196 8158 12294
rect 6425 11845 6523 11943
rect 6850 11787 6948 11885
rect 7282 11787 7380 11885
rect 7664 11801 7762 11899
rect 8060 11801 8158 11899
rect 6425 11429 6523 11527
rect 6850 11429 6948 11527
rect 7282 11429 7380 11527
rect 7664 11406 7762 11504
rect 8060 11406 8158 11504
rect 6425 11055 6523 11153
rect 6850 10997 6948 11095
rect 7282 10997 7380 11095
rect 7664 11011 7762 11109
rect 8060 11011 8158 11109
rect 6425 10639 6523 10737
rect 6850 10639 6948 10737
rect 7282 10639 7380 10737
rect 7664 10616 7762 10714
rect 8060 10616 8158 10714
rect 6425 10265 6523 10363
rect 6850 10207 6948 10305
rect 7282 10207 7380 10305
rect 7664 10221 7762 10319
rect 8060 10221 8158 10319
rect 6425 9849 6523 9947
rect 6850 9849 6948 9947
rect 7282 9849 7380 9947
rect 7664 9826 7762 9924
rect 8060 9826 8158 9924
rect 6425 9475 6523 9573
rect 6850 9417 6948 9515
rect 7282 9417 7380 9515
rect 7664 9431 7762 9529
rect 8060 9431 8158 9529
rect 2691 9059 2789 9157
rect 3116 9059 3214 9157
rect 3548 9059 3646 9157
rect 3930 9036 4028 9134
rect 4326 9036 4424 9134
rect 6425 9059 6523 9157
rect 6850 9059 6948 9157
rect 7282 9059 7380 9157
rect 7664 9036 7762 9134
rect 8060 9036 8158 9134
rect 6425 8685 6523 8783
rect 6850 8627 6948 8725
rect 7282 8627 7380 8725
rect 7664 8641 7762 8739
rect 8060 8641 8158 8739
rect 2691 8269 2789 8367
rect 3116 8269 3214 8367
rect 3548 8269 3646 8367
rect 3930 8246 4028 8344
rect 4326 8246 4424 8344
rect 6425 8269 6523 8367
rect 6850 8269 6948 8367
rect 7282 8269 7380 8367
rect 7664 8246 7762 8344
rect 8060 8246 8158 8344
rect 6425 7895 6523 7993
rect 6850 7837 6948 7935
rect 7282 7837 7380 7935
rect 7664 7851 7762 7949
rect 8060 7851 8158 7949
rect 2691 7479 2789 7577
rect 3116 7479 3214 7577
rect 3548 7479 3646 7577
rect 3930 7456 4028 7554
rect 4326 7456 4424 7554
rect 6425 7479 6523 7577
rect 6850 7479 6948 7577
rect 7282 7479 7380 7577
rect 7664 7456 7762 7554
rect 8060 7456 8158 7554
rect 6425 7105 6523 7203
rect 6850 7047 6948 7145
rect 7282 7047 7380 7145
rect 7664 7061 7762 7159
rect 8060 7061 8158 7159
rect 1236 6666 1334 6764
rect 1632 6666 1730 6764
rect 2691 6689 2789 6787
rect 3116 6689 3214 6787
rect 3548 6689 3646 6787
rect 3930 6666 4028 6764
rect 4326 6666 4424 6764
rect 6425 6689 6523 6787
rect 6850 6689 6948 6787
rect 7282 6689 7380 6787
rect 7664 6666 7762 6764
rect 8060 6666 8158 6764
rect 6425 6315 6523 6413
rect 6850 6257 6948 6355
rect 7282 6257 7380 6355
rect 7664 6271 7762 6369
rect 8060 6271 8158 6369
rect 6425 5899 6523 5997
rect 6850 5899 6948 5997
rect 7282 5899 7380 5997
rect 7664 5876 7762 5974
rect 8060 5876 8158 5974
rect 6425 5525 6523 5623
rect 6850 5467 6948 5565
rect 7282 5467 7380 5565
rect 7664 5481 7762 5579
rect 8060 5481 8158 5579
rect 2691 5109 2789 5207
rect 3116 5109 3214 5207
rect 3548 5109 3646 5207
rect 3930 5086 4028 5184
rect 4326 5086 4424 5184
rect 6425 5109 6523 5207
rect 6850 5109 6948 5207
rect 7282 5109 7380 5207
rect 7664 5086 7762 5184
rect 8060 5086 8158 5184
rect 6425 4735 6523 4833
rect 6850 4677 6948 4775
rect 7282 4677 7380 4775
rect 7664 4691 7762 4789
rect 8060 4691 8158 4789
rect 2691 4319 2789 4417
rect 3116 4319 3214 4417
rect 3548 4319 3646 4417
rect 3930 4296 4028 4394
rect 4326 4296 4424 4394
rect 6425 4319 6523 4417
rect 6850 4319 6948 4417
rect 7282 4319 7380 4417
rect 7664 4296 7762 4394
rect 8060 4296 8158 4394
rect 6425 3945 6523 4043
rect 6850 3887 6948 3985
rect 7282 3887 7380 3985
rect 7664 3901 7762 3999
rect 8060 3901 8158 3999
rect 2691 3529 2789 3627
rect 3116 3529 3214 3627
rect 3548 3529 3646 3627
rect 3930 3506 4028 3604
rect 4326 3506 4424 3604
rect 6425 3529 6523 3627
rect 6850 3529 6948 3627
rect 7282 3529 7380 3627
rect 7664 3506 7762 3604
rect 8060 3506 8158 3604
rect 6425 3155 6523 3253
rect 6850 3097 6948 3195
rect 7282 3097 7380 3195
rect 7664 3111 7762 3209
rect 8060 3111 8158 3209
rect 1236 2716 1334 2814
rect 1632 2716 1730 2814
rect 2691 2739 2789 2837
rect 3116 2739 3214 2837
rect 3548 2739 3646 2837
rect 3930 2716 4028 2814
rect 4326 2716 4424 2814
rect 6425 2739 6523 2837
rect 6850 2739 6948 2837
rect 7282 2739 7380 2837
rect 7664 2716 7762 2814
rect 8060 2716 8158 2814
rect 6425 2365 6523 2463
rect 6850 2307 6948 2405
rect 7282 2307 7380 2405
rect 7664 2321 7762 2419
rect 8060 2321 8158 2419
rect 6425 1949 6523 2047
rect 6850 1949 6948 2047
rect 7282 1949 7380 2047
rect 7664 1926 7762 2024
rect 8060 1926 8158 2024
rect 6425 1575 6523 1673
rect 6850 1517 6948 1615
rect 7282 1517 7380 1615
rect 7664 1531 7762 1629
rect 8060 1531 8158 1629
rect 3126 1143 3224 1241
rect 3551 1143 3649 1241
rect 3930 1136 4028 1234
rect 4326 1136 4424 1234
rect 6425 1159 6523 1257
rect 6850 1159 6948 1257
rect 7282 1159 7380 1257
rect 7664 1136 7762 1234
rect 8060 1136 8158 1234
rect 6425 785 6523 883
rect 6850 727 6948 825
rect 7282 727 7380 825
rect 7664 741 7762 839
rect 8060 741 8158 839
rect 1832 346 1930 444
rect 2228 346 2326 444
rect 3126 353 3224 451
rect 3551 353 3649 451
rect 3930 346 4028 444
rect 4326 346 4424 444
rect 6425 369 6523 467
rect 6850 369 6948 467
rect 7282 369 7380 467
rect 7664 346 7762 444
rect 8060 346 8158 444
use contact_9  contact_9_3
timestamp 1624494425
transform 1 0 9976 0 1 50523
box 0 0 66 74
use contact_8  contact_8_3
timestamp 1624494425
transform 1 0 9977 0 1 50528
box 0 0 64 64
use contact_9  contact_9_4
timestamp 1624494425
transform 1 0 8508 0 1 50508
box 0 0 66 74
use contact_8  contact_8_4
timestamp 1624494425
transform 1 0 8509 0 1 50513
box 0 0 64 64
use contact_9  contact_9_5
timestamp 1624494425
transform 1 0 11624 0 1 50523
box 0 0 66 74
use contact_8  contact_8_5
timestamp 1624494425
transform 1 0 11625 0 1 50528
box 0 0 64 64
use contact_9  contact_9_6
timestamp 1624494425
transform 1 0 8933 0 1 50507
box 0 0 66 74
use contact_8  contact_8_6
timestamp 1624494425
transform 1 0 8934 0 1 50512
box 0 0 64 64
use contact_7  contact_7_1
timestamp 1624494425
transform 1 0 8345 0 1 101386
box 0 0 58 66
use contact_8  contact_8_7
timestamp 1624494425
transform 1 0 8342 0 1 101387
box 0 0 64 64
use contact_8  contact_8_2
timestamp 1624494425
transform 1 0 8934 0 1 101273
box 0 0 64 64
use contact_9  contact_9_2
timestamp 1624494425
transform 1 0 8933 0 1 101268
box 0 0 66 74
use contact_8  contact_8_1
timestamp 1624494425
transform 1 0 11625 0 1 101286
box 0 0 64 64
use contact_9  contact_9_1
timestamp 1624494425
transform 1 0 11624 0 1 101280
box 0 0 66 74
use contact_7  contact_7_0
timestamp 1624494425
transform 1 0 8105 0 1 101278
box 0 0 58 66
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 8102 0 1 101279
box 0 0 64 64
use contact_9  contact_9_0
timestamp 1624494425
transform 1 0 8101 0 1 101274
box 0 0 66 74
use and2_dec_0  and2_dec_0_0
timestamp 1624494425
transform 1 0 8271 0 1 101120
box 70 -56 4140 490
use wordline_driver_array  wordline_driver_array_0
timestamp 1624494425
transform 1 0 8271 0 1 0
box 70 -56 4140 101176
use hierarchical_decoder  hierarchical_decoder_0
timestamp 1624494425
transform 1 0 0 0 1 0
box 0 -60 8275 101180
<< labels >>
rlabel metal1 s 19 0 47 9480 4 addr_0
rlabel metal1 s 99 0 127 9480 4 addr_1
rlabel metal1 s 179 0 207 9480 4 addr_2
rlabel metal1 s 259 0 287 9480 4 addr_3
rlabel metal1 s 339 0 367 9480 4 addr_4
rlabel metal1 s 419 0 447 9480 4 addr_5
rlabel metal1 s 499 0 527 9480 4 addr_6
rlabel metal1 s 579 0 607 9480 4 addr_7
rlabel locali s 12379 120 12379 120 4 wl_0
rlabel locali s 12379 670 12379 670 4 wl_1
rlabel locali s 12379 910 12379 910 4 wl_2
rlabel locali s 12379 1460 12379 1460 4 wl_3
rlabel locali s 12379 1700 12379 1700 4 wl_4
rlabel locali s 12379 2250 12379 2250 4 wl_5
rlabel locali s 12379 2490 12379 2490 4 wl_6
rlabel locali s 12379 3040 12379 3040 4 wl_7
rlabel locali s 12379 3280 12379 3280 4 wl_8
rlabel locali s 12379 3830 12379 3830 4 wl_9
rlabel locali s 12379 4070 12379 4070 4 wl_10
rlabel locali s 12379 4620 12379 4620 4 wl_11
rlabel locali s 12379 4860 12379 4860 4 wl_12
rlabel locali s 12379 5410 12379 5410 4 wl_13
rlabel locali s 12379 5650 12379 5650 4 wl_14
rlabel locali s 12379 6200 12379 6200 4 wl_15
rlabel locali s 12379 6440 12379 6440 4 wl_16
rlabel locali s 12379 6990 12379 6990 4 wl_17
rlabel locali s 12379 7230 12379 7230 4 wl_18
rlabel locali s 12379 7780 12379 7780 4 wl_19
rlabel locali s 12379 8020 12379 8020 4 wl_20
rlabel locali s 12379 8570 12379 8570 4 wl_21
rlabel locali s 12379 8810 12379 8810 4 wl_22
rlabel locali s 12379 9360 12379 9360 4 wl_23
rlabel locali s 12379 9600 12379 9600 4 wl_24
rlabel locali s 12379 10150 12379 10150 4 wl_25
rlabel locali s 12379 10390 12379 10390 4 wl_26
rlabel locali s 12379 10940 12379 10940 4 wl_27
rlabel locali s 12379 11180 12379 11180 4 wl_28
rlabel locali s 12379 11730 12379 11730 4 wl_29
rlabel locali s 12379 11970 12379 11970 4 wl_30
rlabel locali s 12379 12520 12379 12520 4 wl_31
rlabel locali s 12379 12760 12379 12760 4 wl_32
rlabel locali s 12379 13310 12379 13310 4 wl_33
rlabel locali s 12379 13550 12379 13550 4 wl_34
rlabel locali s 12379 14100 12379 14100 4 wl_35
rlabel locali s 12379 14340 12379 14340 4 wl_36
rlabel locali s 12379 14890 12379 14890 4 wl_37
rlabel locali s 12379 15130 12379 15130 4 wl_38
rlabel locali s 12379 15680 12379 15680 4 wl_39
rlabel locali s 12379 15920 12379 15920 4 wl_40
rlabel locali s 12379 16470 12379 16470 4 wl_41
rlabel locali s 12379 16710 12379 16710 4 wl_42
rlabel locali s 12379 17260 12379 17260 4 wl_43
rlabel locali s 12379 17500 12379 17500 4 wl_44
rlabel locali s 12379 18050 12379 18050 4 wl_45
rlabel locali s 12379 18290 12379 18290 4 wl_46
rlabel locali s 12379 18840 12379 18840 4 wl_47
rlabel locali s 12379 19080 12379 19080 4 wl_48
rlabel locali s 12379 19630 12379 19630 4 wl_49
rlabel locali s 12379 19870 12379 19870 4 wl_50
rlabel locali s 12379 20420 12379 20420 4 wl_51
rlabel locali s 12379 20660 12379 20660 4 wl_52
rlabel locali s 12379 21210 12379 21210 4 wl_53
rlabel locali s 12379 21450 12379 21450 4 wl_54
rlabel locali s 12379 22000 12379 22000 4 wl_55
rlabel locali s 12379 22240 12379 22240 4 wl_56
rlabel locali s 12379 22790 12379 22790 4 wl_57
rlabel locali s 12379 23030 12379 23030 4 wl_58
rlabel locali s 12379 23580 12379 23580 4 wl_59
rlabel locali s 12379 23820 12379 23820 4 wl_60
rlabel locali s 12379 24370 12379 24370 4 wl_61
rlabel locali s 12379 24610 12379 24610 4 wl_62
rlabel locali s 12379 25160 12379 25160 4 wl_63
rlabel locali s 12379 25400 12379 25400 4 wl_64
rlabel locali s 12379 25950 12379 25950 4 wl_65
rlabel locali s 12379 26190 12379 26190 4 wl_66
rlabel locali s 12379 26740 12379 26740 4 wl_67
rlabel locali s 12379 26980 12379 26980 4 wl_68
rlabel locali s 12379 27530 12379 27530 4 wl_69
rlabel locali s 12379 27770 12379 27770 4 wl_70
rlabel locali s 12379 28320 12379 28320 4 wl_71
rlabel locali s 12379 28560 12379 28560 4 wl_72
rlabel locali s 12379 29110 12379 29110 4 wl_73
rlabel locali s 12379 29350 12379 29350 4 wl_74
rlabel locali s 12379 29900 12379 29900 4 wl_75
rlabel locali s 12379 30140 12379 30140 4 wl_76
rlabel locali s 12379 30690 12379 30690 4 wl_77
rlabel locali s 12379 30930 12379 30930 4 wl_78
rlabel locali s 12379 31480 12379 31480 4 wl_79
rlabel locali s 12379 31720 12379 31720 4 wl_80
rlabel locali s 12379 32270 12379 32270 4 wl_81
rlabel locali s 12379 32510 12379 32510 4 wl_82
rlabel locali s 12379 33060 12379 33060 4 wl_83
rlabel locali s 12379 33300 12379 33300 4 wl_84
rlabel locali s 12379 33850 12379 33850 4 wl_85
rlabel locali s 12379 34090 12379 34090 4 wl_86
rlabel locali s 12379 34640 12379 34640 4 wl_87
rlabel locali s 12379 34880 12379 34880 4 wl_88
rlabel locali s 12379 35430 12379 35430 4 wl_89
rlabel locali s 12379 35670 12379 35670 4 wl_90
rlabel locali s 12379 36220 12379 36220 4 wl_91
rlabel locali s 12379 36460 12379 36460 4 wl_92
rlabel locali s 12379 37010 12379 37010 4 wl_93
rlabel locali s 12379 37250 12379 37250 4 wl_94
rlabel locali s 12379 37800 12379 37800 4 wl_95
rlabel locali s 12379 38040 12379 38040 4 wl_96
rlabel locali s 12379 38590 12379 38590 4 wl_97
rlabel locali s 12379 38830 12379 38830 4 wl_98
rlabel locali s 12379 39380 12379 39380 4 wl_99
rlabel locali s 12379 39620 12379 39620 4 wl_100
rlabel locali s 12379 40170 12379 40170 4 wl_101
rlabel locali s 12379 40410 12379 40410 4 wl_102
rlabel locali s 12379 40960 12379 40960 4 wl_103
rlabel locali s 12379 41200 12379 41200 4 wl_104
rlabel locali s 12379 41750 12379 41750 4 wl_105
rlabel locali s 12379 41990 12379 41990 4 wl_106
rlabel locali s 12379 42540 12379 42540 4 wl_107
rlabel locali s 12379 42780 12379 42780 4 wl_108
rlabel locali s 12379 43330 12379 43330 4 wl_109
rlabel locali s 12379 43570 12379 43570 4 wl_110
rlabel locali s 12379 44120 12379 44120 4 wl_111
rlabel locali s 12379 44360 12379 44360 4 wl_112
rlabel locali s 12379 44910 12379 44910 4 wl_113
rlabel locali s 12379 45150 12379 45150 4 wl_114
rlabel locali s 12379 45700 12379 45700 4 wl_115
rlabel locali s 12379 45940 12379 45940 4 wl_116
rlabel locali s 12379 46490 12379 46490 4 wl_117
rlabel locali s 12379 46730 12379 46730 4 wl_118
rlabel locali s 12379 47280 12379 47280 4 wl_119
rlabel locali s 12379 47520 12379 47520 4 wl_120
rlabel locali s 12379 48070 12379 48070 4 wl_121
rlabel locali s 12379 48310 12379 48310 4 wl_122
rlabel locali s 12379 48860 12379 48860 4 wl_123
rlabel locali s 12379 49100 12379 49100 4 wl_124
rlabel locali s 12379 49650 12379 49650 4 wl_125
rlabel locali s 12379 49890 12379 49890 4 wl_126
rlabel locali s 12379 50440 12379 50440 4 wl_127
rlabel locali s 12379 50680 12379 50680 4 wl_128
rlabel locali s 12379 51230 12379 51230 4 wl_129
rlabel locali s 12379 51470 12379 51470 4 wl_130
rlabel locali s 12379 52020 12379 52020 4 wl_131
rlabel locali s 12379 52260 12379 52260 4 wl_132
rlabel locali s 12379 52810 12379 52810 4 wl_133
rlabel locali s 12379 53050 12379 53050 4 wl_134
rlabel locali s 12379 53600 12379 53600 4 wl_135
rlabel locali s 12379 53840 12379 53840 4 wl_136
rlabel locali s 12379 54390 12379 54390 4 wl_137
rlabel locali s 12379 54630 12379 54630 4 wl_138
rlabel locali s 12379 55180 12379 55180 4 wl_139
rlabel locali s 12379 55420 12379 55420 4 wl_140
rlabel locali s 12379 55970 12379 55970 4 wl_141
rlabel locali s 12379 56210 12379 56210 4 wl_142
rlabel locali s 12379 56760 12379 56760 4 wl_143
rlabel locali s 12379 57000 12379 57000 4 wl_144
rlabel locali s 12379 57550 12379 57550 4 wl_145
rlabel locali s 12379 57790 12379 57790 4 wl_146
rlabel locali s 12379 58340 12379 58340 4 wl_147
rlabel locali s 12379 58580 12379 58580 4 wl_148
rlabel locali s 12379 59130 12379 59130 4 wl_149
rlabel locali s 12379 59370 12379 59370 4 wl_150
rlabel locali s 12379 59920 12379 59920 4 wl_151
rlabel locali s 12379 60160 12379 60160 4 wl_152
rlabel locali s 12379 60710 12379 60710 4 wl_153
rlabel locali s 12379 60950 12379 60950 4 wl_154
rlabel locali s 12379 61500 12379 61500 4 wl_155
rlabel locali s 12379 61740 12379 61740 4 wl_156
rlabel locali s 12379 62290 12379 62290 4 wl_157
rlabel locali s 12379 62530 12379 62530 4 wl_158
rlabel locali s 12379 63080 12379 63080 4 wl_159
rlabel locali s 12379 63320 12379 63320 4 wl_160
rlabel locali s 12379 63870 12379 63870 4 wl_161
rlabel locali s 12379 64110 12379 64110 4 wl_162
rlabel locali s 12379 64660 12379 64660 4 wl_163
rlabel locali s 12379 64900 12379 64900 4 wl_164
rlabel locali s 12379 65450 12379 65450 4 wl_165
rlabel locali s 12379 65690 12379 65690 4 wl_166
rlabel locali s 12379 66240 12379 66240 4 wl_167
rlabel locali s 12379 66480 12379 66480 4 wl_168
rlabel locali s 12379 67030 12379 67030 4 wl_169
rlabel locali s 12379 67270 12379 67270 4 wl_170
rlabel locali s 12379 67820 12379 67820 4 wl_171
rlabel locali s 12379 68060 12379 68060 4 wl_172
rlabel locali s 12379 68610 12379 68610 4 wl_173
rlabel locali s 12379 68850 12379 68850 4 wl_174
rlabel locali s 12379 69400 12379 69400 4 wl_175
rlabel locali s 12379 69640 12379 69640 4 wl_176
rlabel locali s 12379 70190 12379 70190 4 wl_177
rlabel locali s 12379 70430 12379 70430 4 wl_178
rlabel locali s 12379 70980 12379 70980 4 wl_179
rlabel locali s 12379 71220 12379 71220 4 wl_180
rlabel locali s 12379 71770 12379 71770 4 wl_181
rlabel locali s 12379 72010 12379 72010 4 wl_182
rlabel locali s 12379 72560 12379 72560 4 wl_183
rlabel locali s 12379 72800 12379 72800 4 wl_184
rlabel locali s 12379 73350 12379 73350 4 wl_185
rlabel locali s 12379 73590 12379 73590 4 wl_186
rlabel locali s 12379 74140 12379 74140 4 wl_187
rlabel locali s 12379 74380 12379 74380 4 wl_188
rlabel locali s 12379 74930 12379 74930 4 wl_189
rlabel locali s 12379 75170 12379 75170 4 wl_190
rlabel locali s 12379 75720 12379 75720 4 wl_191
rlabel locali s 12379 75960 12379 75960 4 wl_192
rlabel locali s 12379 76510 12379 76510 4 wl_193
rlabel locali s 12379 76750 12379 76750 4 wl_194
rlabel locali s 12379 77300 12379 77300 4 wl_195
rlabel locali s 12379 77540 12379 77540 4 wl_196
rlabel locali s 12379 78090 12379 78090 4 wl_197
rlabel locali s 12379 78330 12379 78330 4 wl_198
rlabel locali s 12379 78880 12379 78880 4 wl_199
rlabel locali s 12379 79120 12379 79120 4 wl_200
rlabel locali s 12379 79670 12379 79670 4 wl_201
rlabel locali s 12379 79910 12379 79910 4 wl_202
rlabel locali s 12379 80460 12379 80460 4 wl_203
rlabel locali s 12379 80700 12379 80700 4 wl_204
rlabel locali s 12379 81250 12379 81250 4 wl_205
rlabel locali s 12379 81490 12379 81490 4 wl_206
rlabel locali s 12379 82040 12379 82040 4 wl_207
rlabel locali s 12379 82280 12379 82280 4 wl_208
rlabel locali s 12379 82830 12379 82830 4 wl_209
rlabel locali s 12379 83070 12379 83070 4 wl_210
rlabel locali s 12379 83620 12379 83620 4 wl_211
rlabel locali s 12379 83860 12379 83860 4 wl_212
rlabel locali s 12379 84410 12379 84410 4 wl_213
rlabel locali s 12379 84650 12379 84650 4 wl_214
rlabel locali s 12379 85200 12379 85200 4 wl_215
rlabel locali s 12379 85440 12379 85440 4 wl_216
rlabel locali s 12379 85990 12379 85990 4 wl_217
rlabel locali s 12379 86230 12379 86230 4 wl_218
rlabel locali s 12379 86780 12379 86780 4 wl_219
rlabel locali s 12379 87020 12379 87020 4 wl_220
rlabel locali s 12379 87570 12379 87570 4 wl_221
rlabel locali s 12379 87810 12379 87810 4 wl_222
rlabel locali s 12379 88360 12379 88360 4 wl_223
rlabel locali s 12379 88600 12379 88600 4 wl_224
rlabel locali s 12379 89150 12379 89150 4 wl_225
rlabel locali s 12379 89390 12379 89390 4 wl_226
rlabel locali s 12379 89940 12379 89940 4 wl_227
rlabel locali s 12379 90180 12379 90180 4 wl_228
rlabel locali s 12379 90730 12379 90730 4 wl_229
rlabel locali s 12379 90970 12379 90970 4 wl_230
rlabel locali s 12379 91520 12379 91520 4 wl_231
rlabel locali s 12379 91760 12379 91760 4 wl_232
rlabel locali s 12379 92310 12379 92310 4 wl_233
rlabel locali s 12379 92550 12379 92550 4 wl_234
rlabel locali s 12379 93100 12379 93100 4 wl_235
rlabel locali s 12379 93340 12379 93340 4 wl_236
rlabel locali s 12379 93890 12379 93890 4 wl_237
rlabel locali s 12379 94130 12379 94130 4 wl_238
rlabel locali s 12379 94680 12379 94680 4 wl_239
rlabel locali s 12379 94920 12379 94920 4 wl_240
rlabel locali s 12379 95470 12379 95470 4 wl_241
rlabel locali s 12379 95710 12379 95710 4 wl_242
rlabel locali s 12379 96260 12379 96260 4 wl_243
rlabel locali s 12379 96500 12379 96500 4 wl_244
rlabel locali s 12379 97050 12379 97050 4 wl_245
rlabel locali s 12379 97290 12379 97290 4 wl_246
rlabel locali s 12379 97840 12379 97840 4 wl_247
rlabel locali s 12379 98080 12379 98080 4 wl_248
rlabel locali s 12379 98630 12379 98630 4 wl_249
rlabel locali s 12379 98870 12379 98870 4 wl_250
rlabel locali s 12379 99420 12379 99420 4 wl_251
rlabel locali s 12379 99660 12379 99660 4 wl_252
rlabel locali s 12379 100210 12379 100210 4 wl_253
rlabel locali s 12379 100450 12379 100450 4 wl_254
rlabel locali s 12379 101000 12379 101000 4 wl_255
rlabel locali s 11184 101240 11184 101240 4 rbl_wl
rlabel metal2 s 8360 101405 8388 101433 4 wl_en
rlabel metal3 s 8060 98701 8158 98799 4 vdd
rlabel metal3 s 7282 52077 7380 52175 4 vdd
rlabel metal3 s 6850 32327 6948 32425 4 vdd
rlabel metal3 s 8060 67891 8158 67989 4 vdd
rlabel metal3 s 6850 20119 6948 20217 4 vdd
rlabel metal3 s 6850 40227 6948 40325 4 vdd
rlabel metal3 s 3548 8269 3646 8367 4 vdd
rlabel metal3 s 8060 2716 8158 2814 4 vdd
rlabel metal3 s 6850 90787 6948 90885 4 vdd
rlabel metal3 s 8060 67101 8158 67199 4 vdd
rlabel metal3 s 6850 98329 6948 98427 4 vdd
rlabel metal3 s 7282 93947 7380 94045 4 vdd
rlabel metal3 s 7282 81307 7380 81405 4 vdd
rlabel metal3 s 7282 66297 7380 66395 4 vdd
rlabel metal3 s 8060 100676 8158 100774 4 vdd
rlabel metal3 s 8060 5086 8158 5184 4 vdd
rlabel metal3 s 4326 9036 4424 9134 4 vdd
rlabel metal3 s 6850 63927 6948 64025 4 vdd
rlabel metal3 s 8060 35896 8158 35994 4 vdd
rlabel metal3 s 8060 57621 8158 57719 4 vdd
rlabel metal3 s 6850 14947 6948 15045 4 vdd
rlabel metal3 s 4326 1136 4424 1234 4 vdd
rlabel metal3 s 8060 33526 8158 33624 4 vdd
rlabel metal3 s 7282 53657 7380 53755 4 vdd
rlabel metal3 s 6850 23637 6948 23735 4 vdd
rlabel metal3 s 3116 6689 3214 6787 4 vdd
rlabel metal3 s 7282 7837 7380 7935 4 vdd
rlabel metal3 s 8060 8246 8158 8344 4 vdd
rlabel metal3 s 7282 60767 7380 60865 4 vdd
rlabel metal3 s 8060 59596 8158 59694 4 vdd
rlabel metal3 s 7282 44609 7380 44707 4 vdd
rlabel metal3 s 7282 23637 7380 23735 4 vdd
rlabel metal3 s 7282 84109 7380 84207 4 vdd
rlabel metal3 s 7282 26439 7380 26537 4 vdd
rlabel metal3 s 6850 97897 6948 97995 4 vdd
rlabel metal3 s 8060 78556 8158 78654 4 vdd
rlabel metal3 s 6850 6257 6948 6355 4 vdd
rlabel metal3 s 6850 88849 6948 88947 4 vdd
rlabel metal3 s 6850 38289 6948 38387 4 vdd
rlabel metal3 s 7282 92799 7380 92897 4 vdd
rlabel metal3 s 6850 85257 6948 85355 4 vdd
rlabel metal3 s 6850 83677 6948 83775 4 vdd
rlabel metal3 s 7282 3529 7380 3627 4 vdd
rlabel metal3 s 7282 57607 7380 57705 4 vdd
rlabel metal3 s 6850 4677 6948 4775 4 vdd
rlabel metal3 s 8060 79346 8158 79444 4 vdd
rlabel metal3 s 6850 54447 6948 54545 4 vdd
rlabel metal3 s 7282 69889 7380 69987 4 vdd
rlabel metal3 s 7282 52867 7380 52965 4 vdd
rlabel metal3 s 8060 58016 8158 58114 4 vdd
rlabel metal3 s 7282 67087 7380 67185 4 vdd
rlabel metal3 s 8060 51301 8158 51399 4 vdd
rlabel metal3 s 7282 35487 7380 35585 4 vdd
rlabel metal3 s 6850 31537 6948 31635 4 vdd
rlabel metal3 s 6850 1517 6948 1615 4 vdd
rlabel metal3 s 7282 90787 7380 90885 4 vdd
rlabel metal3 s 6850 26007 6948 26105 4 vdd
rlabel metal3 s 8060 31946 8158 32044 4 vdd
rlabel metal3 s 6850 39869 6948 39967 4 vdd
rlabel metal3 s 6850 50497 6948 50595 4 vdd
rlabel metal3 s 6850 22847 6948 22945 4 vdd
rlabel metal3 s 7282 68667 7380 68765 4 vdd
rlabel metal3 s 8060 48141 8158 48239 4 vdd
rlabel metal3 s 7282 20909 7380 21007 4 vdd
rlabel metal3 s 6850 67087 6948 67185 4 vdd
rlabel metal3 s 8060 26416 8158 26514 4 vdd
rlabel metal3 s 8060 54856 8158 54954 4 vdd
rlabel metal3 s 7282 56027 7380 56125 4 vdd
rlabel metal3 s 7282 56817 7380 56915 4 vdd
rlabel metal3 s 6850 37067 6948 37165 4 vdd
rlabel metal3 s 7282 85257 7380 85355 4 vdd
rlabel metal3 s 8060 82111 8158 82209 4 vdd
rlabel metal3 s 8060 35501 8158 35599 4 vdd
rlabel metal3 s 7282 21699 7380 21797 4 vdd
rlabel metal3 s 6850 99477 6948 99575 4 vdd
rlabel metal3 s 8060 99096 8158 99194 4 vdd
rlabel metal3 s 8060 54066 8158 54164 4 vdd
rlabel metal3 s 8060 18121 8158 18219 4 vdd
rlabel metal3 s 7282 26797 7380 26895 4 vdd
rlabel metal3 s 7282 39437 7380 39535 4 vdd
rlabel metal3 s 8060 73816 8158 73914 4 vdd
rlabel metal3 s 4326 346 4424 444 4 vdd
rlabel metal3 s 8060 80926 8158 81024 4 vdd
rlabel metal3 s 8060 28786 8158 28884 4 vdd
rlabel metal3 s 6850 21699 6948 21797 4 vdd
rlabel metal3 s 7282 24427 7380 24525 4 vdd
rlabel metal3 s 8060 58411 8158 58509 4 vdd
rlabel metal3 s 6850 63569 6948 63667 4 vdd
rlabel metal3 s 6850 49707 6948 49805 4 vdd
rlabel metal3 s 6850 65507 6948 65605 4 vdd
rlabel metal3 s 8060 71446 8158 71544 4 vdd
rlabel metal3 s 7282 86837 7380 86935 4 vdd
rlabel metal3 s 7282 98329 7380 98427 4 vdd
rlabel metal3 s 7282 56459 7380 56557 4 vdd
rlabel metal3 s 7282 76567 7380 76665 4 vdd
rlabel metal3 s 6850 3887 6948 3985 4 vdd
rlabel metal3 s 6850 79727 6948 79825 4 vdd
rlabel metal3 s 8060 76581 8158 76679 4 vdd
rlabel metal3 s 8060 64336 8158 64434 4 vdd
rlabel metal3 s 8060 68681 8158 68779 4 vdd
rlabel metal3 s 7282 18107 7380 18205 4 vdd
rlabel metal3 s 6850 48559 6948 48657 4 vdd
rlabel metal3 s 7282 65149 7380 65247 4 vdd
rlabel metal3 s 8060 85666 8158 85764 4 vdd
rlabel metal3 s 6850 24859 6948 24957 4 vdd
rlabel metal3 s 6850 58039 6948 58137 4 vdd
rlabel metal3 s 6850 91219 6948 91317 4 vdd
rlabel metal3 s 6850 2307 6948 2405 4 vdd
rlabel metal3 s 6850 13009 6948 13107 4 vdd
rlabel metal3 s 7282 60409 7380 60507 4 vdd
rlabel metal3 s 8060 45771 8158 45869 4 vdd
rlabel metal3 s 7282 10639 7380 10737 4 vdd
rlabel metal3 s 8060 85271 8158 85369 4 vdd
rlabel metal3 s 7282 14589 7380 14687 4 vdd
rlabel metal3 s 6850 77789 6948 77887 4 vdd
rlabel metal3 s 7282 12577 7380 12675 4 vdd
rlabel metal3 s 7282 41017 7380 41115 4 vdd
rlabel metal3 s 6850 64717 6948 64815 4 vdd
rlabel metal3 s 7282 38289 7380 38387 4 vdd
rlabel metal3 s 7282 16959 7380 17057 4 vdd
rlabel metal3 s 7282 95527 7380 95625 4 vdd
rlabel metal3 s 8060 66706 8158 66804 4 vdd
rlabel metal3 s 7282 46189 7380 46287 4 vdd
rlabel metal3 s 6850 42597 6948 42695 4 vdd
rlabel metal3 s 6850 100267 6948 100365 4 vdd
rlabel metal3 s 7282 13367 7380 13465 4 vdd
rlabel metal3 s 6850 19687 6948 19785 4 vdd
rlabel metal3 s 6850 84899 6948 84997 4 vdd
rlabel metal3 s 6850 50929 6948 51027 4 vdd
rlabel metal3 s 7282 54447 7380 54545 4 vdd
rlabel metal3 s 8060 18516 8158 18614 4 vdd
rlabel metal3 s 8060 24441 8158 24539 4 vdd
rlabel metal3 s 7282 98687 7380 98785 4 vdd
rlabel metal3 s 8060 55251 8158 55349 4 vdd
rlabel metal3 s 6850 82887 6948 82985 4 vdd
rlabel metal3 s 8060 86851 8158 86949 4 vdd
rlabel metal3 s 3116 9059 3214 9157 4 vdd
rlabel metal3 s 3548 4319 3646 4417 4 vdd
rlabel metal3 s 6850 54879 6948 54977 4 vdd
rlabel metal3 s 7282 94379 7380 94477 4 vdd
rlabel metal3 s 7282 50497 7380 50595 4 vdd
rlabel metal3 s 7282 9849 7380 9947 4 vdd
rlabel metal3 s 4326 8246 4424 8344 4 vdd
rlabel metal3 s 8060 3506 8158 3604 4 vdd
rlabel metal3 s 6850 87627 6948 87725 4 vdd
rlabel metal3 s 8060 25231 8158 25329 4 vdd
rlabel metal3 s 8060 80136 8158 80234 4 vdd
rlabel metal3 s 7282 16527 7380 16625 4 vdd
rlabel metal3 s 4326 6666 4424 6764 4 vdd
rlabel metal3 s 8060 36291 8158 36389 4 vdd
rlabel metal3 s 6850 24427 6948 24525 4 vdd
rlabel metal3 s 7282 70247 7380 70345 4 vdd
rlabel metal3 s 8917 50495 9015 50593 4 vdd
rlabel metal3 s 8060 64731 8158 64829 4 vdd
rlabel metal3 s 7282 55669 7380 55767 4 vdd
rlabel metal3 s 6850 42239 6948 42337 4 vdd
rlabel metal3 s 8060 53276 8158 53374 4 vdd
rlabel metal3 s 6850 7479 6948 7577 4 vdd
rlabel metal3 s 8060 54461 8158 54559 4 vdd
rlabel metal3 s 6850 16959 6948 17057 4 vdd
rlabel metal3 s 3548 9059 3646 9157 4 vdd
rlabel metal3 s 7282 36709 7380 36807 4 vdd
rlabel metal3 s 8060 97516 8158 97614 4 vdd
rlabel metal3 s 7282 70679 7380 70777 4 vdd
rlabel metal3 s 7282 19687 7380 19785 4 vdd
rlabel metal3 s 6850 65149 6948 65247 4 vdd
rlabel metal3 s 6850 97107 6948 97205 4 vdd
rlabel metal3 s 8060 63151 8158 63249 4 vdd
rlabel metal3 s 7282 95169 7380 95267 4 vdd
rlabel metal3 s 6850 83319 6948 83417 4 vdd
rlabel metal3 s 6850 3529 6948 3627 4 vdd
rlabel metal3 s 8060 4296 8158 4394 4 vdd
rlabel metal3 s 8060 87246 8158 87344 4 vdd
rlabel metal3 s 6850 38647 6948 38745 4 vdd
rlabel metal3 s 6850 26439 6948 26537 4 vdd
rlabel metal3 s 6850 76999 6948 77097 4 vdd
rlabel metal3 s 7282 32759 7380 32857 4 vdd
rlabel metal3 s 6850 12577 6948 12675 4 vdd
rlabel metal3 s 8060 72631 8158 72729 4 vdd
rlabel metal3 s 7282 54879 7380 54977 4 vdd
rlabel metal3 s 8060 32341 8158 32439 4 vdd
rlabel metal3 s 8060 19306 8158 19404 4 vdd
rlabel metal3 s 7282 99477 7380 99575 4 vdd
rlabel metal3 s 7282 61199 7380 61297 4 vdd
rlabel metal3 s 8060 31156 8158 31254 4 vdd
rlabel metal3 s 8060 57226 8158 57324 4 vdd
rlabel metal3 s 6850 93589 6948 93687 4 vdd
rlabel metal3 s 8060 90011 8158 90109 4 vdd
rlabel metal3 s 8060 69076 8158 69174 4 vdd
rlabel metal3 s 7282 58039 7380 58137 4 vdd
rlabel metal3 s 6850 43387 6948 43485 4 vdd
rlabel metal3 s 6850 27587 6948 27685 4 vdd
rlabel metal3 s 6850 61199 6948 61297 4 vdd
rlabel metal3 s 6850 31969 6948 32067 4 vdd
rlabel metal3 s 6850 18107 6948 18205 4 vdd
rlabel metal3 s 8060 81716 8158 81814 4 vdd
rlabel metal3 s 6850 5467 6948 5565 4 vdd
rlabel metal3 s 7282 1517 7380 1615 4 vdd
rlabel metal3 s 8060 16936 8158 17034 4 vdd
rlabel metal3 s 6850 17749 6948 17847 4 vdd
rlabel metal3 s 1632 2716 1730 2814 4 vdd
rlabel metal3 s 8060 77371 8158 77469 4 vdd
rlabel metal3 s 6850 52509 6948 52607 4 vdd
rlabel metal3 s 8060 96331 8158 96429 4 vdd
rlabel metal3 s 7282 86047 7380 86145 4 vdd
rlabel metal3 s 7282 28377 7380 28475 4 vdd
rlabel metal3 s 8060 14961 8158 15059 4 vdd
rlabel metal3 s 7282 92009 7380 92107 4 vdd
rlabel metal3 s 8060 56041 8158 56139 4 vdd
rlabel metal3 s 7282 37067 7380 37165 4 vdd
rlabel metal3 s 7282 62779 7380 62877 4 vdd
rlabel metal3 s 6850 15737 6948 15835 4 vdd
rlabel metal3 s 7282 11787 7380 11885 4 vdd
rlabel metal3 s 7282 29599 7380 29697 4 vdd
rlabel metal3 s 8060 65126 8158 65224 4 vdd
rlabel metal3 s 7282 79369 7380 79467 4 vdd
rlabel metal3 s 6850 44177 6948 44275 4 vdd
rlabel metal3 s 8060 7061 8158 7159 4 vdd
rlabel metal3 s 7282 22057 7380 22155 4 vdd
rlabel metal3 s 6850 62347 6948 62445 4 vdd
rlabel metal3 s 6850 369 6948 467 4 vdd
rlabel metal3 s 8060 51696 8158 51794 4 vdd
rlabel metal3 s 7282 4677 7380 4775 4 vdd
rlabel metal3 s 7282 8269 7380 8367 4 vdd
rlabel metal3 s 8060 70261 8158 70359 4 vdd
rlabel metal3 s 7282 46979 7380 47077 4 vdd
rlabel metal3 s 6850 14157 6948 14255 4 vdd
rlabel metal3 s 7282 59977 7380 60075 4 vdd
rlabel metal3 s 7282 1949 7380 2047 4 vdd
rlabel metal3 s 8060 55646 8158 55744 4 vdd
rlabel metal3 s 6850 58829 6948 58927 4 vdd
rlabel metal3 s 6850 89639 6948 89737 4 vdd
rlabel metal3 s 6850 88059 6948 88157 4 vdd
rlabel metal3 s 6850 20909 6948 21007 4 vdd
rlabel metal3 s 7282 84899 7380 84997 4 vdd
rlabel metal3 s 6850 89207 6948 89305 4 vdd
rlabel metal3 s 8060 89616 8158 89714 4 vdd
rlabel metal3 s 8060 72236 8158 72334 4 vdd
rlabel metal3 s 6850 80517 6948 80615 4 vdd
rlabel metal3 s 6850 8627 6948 8725 4 vdd
rlabel metal3 s 6850 73407 6948 73505 4 vdd
rlabel metal3 s 8060 52486 8158 52584 4 vdd
rlabel metal3 s 6850 92799 6948 92897 4 vdd
rlabel metal3 s 6850 37857 6948 37955 4 vdd
rlabel metal3 s 6850 48127 6948 48225 4 vdd
rlabel metal3 s 8060 44191 8158 44289 4 vdd
rlabel metal3 s 8060 41031 8158 41129 4 vdd
rlabel metal3 s 8060 93171 8158 93269 4 vdd
rlabel metal3 s 7282 100699 7380 100797 4 vdd
rlabel metal3 s 8060 94751 8158 94849 4 vdd
rlabel metal3 s 8060 38661 8158 38759 4 vdd
rlabel metal3 s 7282 71827 7380 71925 4 vdd
rlabel metal3 s 7282 80949 7380 81047 4 vdd
rlabel metal3 s 8060 53671 8158 53769 4 vdd
rlabel metal3 s 6850 34697 6948 34795 4 vdd
rlabel metal3 s 8060 15751 8158 15849 4 vdd
rlabel metal3 s 6850 36277 6948 36375 4 vdd
rlabel metal3 s 7282 55237 7380 55335 4 vdd
rlabel metal3 s 8060 62361 8158 62459 4 vdd
rlabel metal3 s 6850 51287 6948 51385 4 vdd
rlabel metal3 s 8060 77766 8158 77864 4 vdd
rlabel metal3 s 7282 65939 7380 66037 4 vdd
rlabel metal3 s 8060 71841 8158 71939 4 vdd
rlabel metal3 s 11608 50511 11706 50609 4 vdd
rlabel metal3 s 8060 90406 8158 90504 4 vdd
rlabel metal3 s 7282 63569 7380 63667 4 vdd
rlabel metal3 s 8060 36686 8158 36784 4 vdd
rlabel metal3 s 6850 61989 6948 62087 4 vdd
rlabel metal3 s 6850 95169 6948 95267 4 vdd
rlabel metal3 s 7282 84467 7380 84565 4 vdd
rlabel metal3 s 8060 83691 8158 83789 4 vdd
rlabel metal3 s 7282 22847 7380 22945 4 vdd
rlabel metal3 s 6850 24069 6948 24167 4 vdd
rlabel metal3 s 8060 46166 8158 46264 4 vdd
rlabel metal3 s 3116 8269 3214 8367 4 vdd
rlabel metal3 s 7282 49349 7380 49447 4 vdd
rlabel metal3 s 8060 39846 8158 39944 4 vdd
rlabel metal3 s 7282 21267 7380 21365 4 vdd
rlabel metal3 s 7282 78937 7380 79035 4 vdd
rlabel metal3 s 8060 44981 8158 45079 4 vdd
rlabel metal3 s 7282 47769 7380 47867 4 vdd
rlabel metal3 s 7282 42597 7380 42695 4 vdd
rlabel metal3 s 7282 39869 7380 39967 4 vdd
rlabel metal3 s 7282 71469 7380 71567 4 vdd
rlabel metal3 s 7282 50139 7380 50237 4 vdd
rlabel metal3 s 6850 10997 6948 11095 4 vdd
rlabel metal3 s 6850 47337 6948 47435 4 vdd
rlabel metal3 s 7282 5899 7380 5997 4 vdd
rlabel metal3 s 8060 91986 8158 92084 4 vdd
rlabel metal3 s 7282 69457 7380 69555 4 vdd
rlabel metal3 s 6850 72617 6948 72715 4 vdd
rlabel metal3 s 8060 11011 8158 11109 4 vdd
rlabel metal3 s 6850 32759 6948 32857 4 vdd
rlabel metal3 s 8060 41426 8158 41524 4 vdd
rlabel metal3 s 7282 727 7380 825 4 vdd
rlabel metal3 s 8060 12196 8158 12294 4 vdd
rlabel metal3 s 6850 86837 6948 86935 4 vdd
rlabel metal3 s 7282 63927 7380 64025 4 vdd
rlabel metal3 s 8060 11406 8158 11504 4 vdd
rlabel metal3 s 6850 33549 6948 33647 4 vdd
rlabel metal3 s 7282 24859 7380 24957 4 vdd
rlabel metal3 s 8917 101256 9015 101354 4 vdd
rlabel metal3 s 7282 36277 7380 36375 4 vdd
rlabel metal3 s 7282 40227 7380 40325 4 vdd
rlabel metal3 s 6850 34339 6948 34437 4 vdd
rlabel metal3 s 6850 8269 6948 8367 4 vdd
rlabel metal3 s 6850 36709 6948 36807 4 vdd
rlabel metal3 s 7282 31179 7380 31277 4 vdd
rlabel metal3 s 8060 93961 8158 94059 4 vdd
rlabel metal3 s 7282 96317 7380 96415 4 vdd
rlabel metal3 s 6850 47769 6948 47867 4 vdd
rlabel metal3 s 7282 48917 7380 49015 4 vdd
rlabel metal3 s 6850 76209 6948 76307 4 vdd
rlabel metal3 s 7282 76209 7380 76307 4 vdd
rlabel metal3 s 7282 51719 7380 51817 4 vdd
rlabel metal3 s 7282 34339 7380 34437 4 vdd
rlabel metal3 s 8060 98306 8158 98404 4 vdd
rlabel metal3 s 7282 2307 7380 2405 4 vdd
rlabel metal3 s 6850 96749 6948 96847 4 vdd
rlabel metal3 s 6850 43029 6948 43127 4 vdd
rlabel metal3 s 8060 6271 8158 6369 4 vdd
rlabel metal3 s 7282 99909 7380 100007 4 vdd
rlabel metal3 s 7282 7047 7380 7145 4 vdd
rlabel metal3 s 8060 8641 8158 8739 4 vdd
rlabel metal3 s 6850 9059 6948 9157 4 vdd
rlabel metal3 s 7282 369 7380 467 4 vdd
rlabel metal3 s 6850 91577 6948 91675 4 vdd
rlabel metal3 s 6850 78937 6948 79035 4 vdd
rlabel metal3 s 6850 41449 6948 41547 4 vdd
rlabel metal3 s 6850 99119 6948 99217 4 vdd
rlabel metal3 s 8060 11801 8158 11899 4 vdd
rlabel metal3 s 7282 28809 7380 28907 4 vdd
rlabel metal3 s 7282 27229 7380 27327 4 vdd
rlabel metal3 s 7282 87269 7380 87367 4 vdd
rlabel metal3 s 7282 38647 7380 38745 4 vdd
rlabel metal3 s 7282 44177 7380 44275 4 vdd
rlabel metal3 s 3548 7479 3646 7577 4 vdd
rlabel metal3 s 7282 19329 7380 19427 4 vdd
rlabel metal3 s 6850 6689 6948 6787 4 vdd
rlabel metal3 s 8060 42216 8158 42314 4 vdd
rlabel metal3 s 7282 50929 7380 51027 4 vdd
rlabel metal3 s 7282 13799 7380 13897 4 vdd
rlabel metal3 s 6850 28019 6948 28117 4 vdd
rlabel metal3 s 8060 56436 8158 56534 4 vdd
rlabel metal3 s 8060 22466 8158 22564 4 vdd
rlabel metal3 s 6850 77357 6948 77455 4 vdd
rlabel metal3 s 11608 101268 11706 101366 4 vdd
rlabel metal3 s 6850 59977 6948 60075 4 vdd
rlabel metal3 s 6850 49349 6948 49447 4 vdd
rlabel metal3 s 6850 63137 6948 63235 4 vdd
rlabel metal3 s 7282 90429 7380 90527 4 vdd
rlabel metal3 s 7282 17749 7380 17847 4 vdd
rlabel metal3 s 6850 25649 6948 25747 4 vdd
rlabel metal3 s 7282 81739 7380 81837 4 vdd
rlabel metal3 s 8060 27601 8158 27699 4 vdd
rlabel metal3 s 7282 34697 7380 34795 4 vdd
rlabel metal3 s 7282 5467 7380 5565 4 vdd
rlabel metal3 s 7282 87627 7380 87725 4 vdd
rlabel metal3 s 7282 5109 7380 5207 4 vdd
rlabel metal3 s 6850 93157 6948 93255 4 vdd
rlabel metal3 s 8060 34711 8158 34809 4 vdd
rlabel metal3 s 8060 67496 8158 67594 4 vdd
rlabel metal3 s 6850 5899 6948 5997 4 vdd
rlabel metal3 s 7282 44967 7380 45065 4 vdd
rlabel metal3 s 8060 39056 8158 39154 4 vdd
rlabel metal3 s 6850 18539 6948 18637 4 vdd
rlabel metal3 s 8060 21676 8158 21774 4 vdd
rlabel metal3 s 6850 4319 6948 4417 4 vdd
rlabel metal3 s 6850 56459 6948 56557 4 vdd
rlabel metal3 s 7282 18897 7380 18995 4 vdd
rlabel metal3 s 7282 89997 7380 90095 4 vdd
rlabel metal3 s 8060 81321 8158 81419 4 vdd
rlabel metal3 s 7282 47337 7380 47435 4 vdd
rlabel metal3 s 8060 48931 8158 49029 4 vdd
rlabel metal3 s 7282 78147 7380 78245 4 vdd
rlabel metal3 s 7282 88849 7380 88947 4 vdd
rlabel metal3 s 4326 7456 4424 7554 4 vdd
rlabel metal3 s 8060 20886 8158 20984 4 vdd
rlabel metal3 s 7282 14947 7380 15045 4 vdd
rlabel metal3 s 8060 37081 8158 37179 4 vdd
rlabel metal3 s 8060 10616 8158 10714 4 vdd
rlabel metal3 s 6850 41017 6948 41115 4 vdd
rlabel metal3 s 6850 9417 6948 9515 4 vdd
rlabel metal3 s 8060 49326 8158 49424 4 vdd
rlabel metal3 s 8060 5876 8158 5974 4 vdd
rlabel metal3 s 7282 58397 7380 58495 4 vdd
rlabel metal3 s 7282 83319 7380 83417 4 vdd
rlabel metal3 s 8060 50906 8158 51004 4 vdd
rlabel metal3 s 6850 89997 6948 90095 4 vdd
rlabel metal3 s 6850 43819 6948 43917 4 vdd
rlabel metal3 s 7282 41807 7380 41905 4 vdd
rlabel metal3 s 7282 64359 7380 64457 4 vdd
rlabel metal3 s 6850 22489 6948 22587 4 vdd
rlabel metal3 s 8060 49721 8158 49819 4 vdd
rlabel metal3 s 6850 28809 6948 28907 4 vdd
rlabel metal3 s 6850 1159 6948 1257 4 vdd
rlabel metal3 s 6850 11787 6948 11885 4 vdd
rlabel metal3 s 7282 74987 7380 75085 4 vdd
rlabel metal3 s 6850 73839 6948 73937 4 vdd
rlabel metal3 s 8060 29576 8158 29674 4 vdd
rlabel metal3 s 6850 93947 6948 94045 4 vdd
rlabel metal3 s 6850 96317 6948 96415 4 vdd
rlabel metal3 s 7282 72259 7380 72357 4 vdd
rlabel metal3 s 7282 35129 7380 35227 4 vdd
rlabel metal3 s 6850 69889 6948 69987 4 vdd
rlabel metal3 s 7282 61557 7380 61655 4 vdd
rlabel metal3 s 8085 101262 8183 101360 4 vdd
rlabel metal3 s 6850 66729 6948 66827 4 vdd
rlabel metal3 s 8060 99491 8158 99589 4 vdd
rlabel metal3 s 8060 12591 8158 12689 4 vdd
rlabel metal3 s 8060 34316 8158 34414 4 vdd
rlabel metal3 s 3548 6689 3646 6787 4 vdd
rlabel metal3 s 6850 35129 6948 35227 4 vdd
rlabel metal3 s 6850 64359 6948 64457 4 vdd
rlabel metal3 s 8060 90801 8158 90899 4 vdd
rlabel metal3 s 6850 58397 6948 58495 4 vdd
rlabel metal3 s 8060 65916 8158 66014 4 vdd
rlabel metal3 s 6850 53299 6948 53397 4 vdd
rlabel metal3 s 7282 30747 7380 30845 4 vdd
rlabel metal3 s 6850 94737 6948 94835 4 vdd
rlabel metal3 s 8060 20491 8158 20589 4 vdd
rlabel metal3 s 6850 82529 6948 82627 4 vdd
rlabel metal3 s 7282 23279 7380 23377 4 vdd
rlabel metal3 s 7282 89207 7380 89305 4 vdd
rlabel metal3 s 8060 61176 8158 61274 4 vdd
rlabel metal3 s 6850 59619 6948 59717 4 vdd
rlabel metal3 s 7282 53299 7380 53397 4 vdd
rlabel metal3 s 8060 19701 8158 19799 4 vdd
rlabel metal3 s 8060 69866 8158 69964 4 vdd
rlabel metal3 s 3116 4319 3214 4417 4 vdd
rlabel metal3 s 6850 14589 6948 14687 4 vdd
rlabel metal3 s 6850 76567 6948 76665 4 vdd
rlabel metal3 s 7282 3097 7380 3195 4 vdd
rlabel metal3 s 7282 6257 7380 6355 4 vdd
rlabel metal3 s 8060 38266 8158 38364 4 vdd
rlabel metal3 s 8060 16541 8158 16639 4 vdd
rlabel metal3 s 6850 68309 6948 68407 4 vdd
rlabel metal3 s 7282 61989 7380 62087 4 vdd
rlabel metal3 s 7282 18539 7380 18637 4 vdd
rlabel metal3 s 8060 1926 8158 2024 4 vdd
rlabel metal3 s 8060 58806 8158 58904 4 vdd
rlabel metal3 s 6850 73049 6948 73147 4 vdd
rlabel metal3 s 6850 44609 6948 44707 4 vdd
rlabel metal3 s 8060 9431 8158 9529 4 vdd
rlabel metal3 s 8060 43401 8158 43499 4 vdd
rlabel metal3 s 8060 66311 8158 66409 4 vdd
rlabel metal3 s 6850 39079 6948 39177 4 vdd
rlabel metal3 s 8060 88826 8158 88924 4 vdd
rlabel metal3 s 8060 21281 8158 21379 4 vdd
rlabel metal3 s 6850 27229 6948 27327 4 vdd
rlabel metal3 s 8060 3901 8158 3999 4 vdd
rlabel metal3 s 8060 37871 8158 37969 4 vdd
rlabel metal3 s 7282 67877 7380 67975 4 vdd
rlabel metal3 s 8060 84876 8158 84974 4 vdd
rlabel metal3 s 7282 48559 7380 48657 4 vdd
rlabel metal3 s 8060 78161 8158 78259 4 vdd
rlabel metal3 s 7282 33117 7380 33215 4 vdd
rlabel metal3 s 8060 86061 8158 86159 4 vdd
rlabel metal3 s 7282 15737 7380 15835 4 vdd
rlabel metal3 s 7282 3887 7380 3985 4 vdd
rlabel metal3 s 8060 75791 8158 75889 4 vdd
rlabel metal3 s 8060 74606 8158 74704 4 vdd
rlabel metal3 s 6850 20477 6948 20575 4 vdd
rlabel metal3 s 8060 6666 8158 6764 4 vdd
rlabel metal3 s 6850 51719 6948 51817 4 vdd
rlabel metal3 s 6850 21267 6948 21365 4 vdd
rlabel metal3 s 8060 24046 8158 24144 4 vdd
rlabel metal3 s 6850 66297 6948 66395 4 vdd
rlabel metal3 s 8060 41821 8158 41919 4 vdd
rlabel metal3 s 8060 46561 8158 46659 4 vdd
rlabel metal3 s 7282 93157 7380 93255 4 vdd
rlabel metal3 s 8060 44586 8158 44684 4 vdd
rlabel metal3 s 7282 22489 7380 22587 4 vdd
rlabel metal3 s 8060 86456 8158 86554 4 vdd
rlabel metal3 s 7282 62347 7380 62445 4 vdd
rlabel metal3 s 8060 17726 8158 17824 4 vdd
rlabel metal3 s 6850 71827 6948 71925 4 vdd
rlabel metal3 s 8060 94356 8158 94454 4 vdd
rlabel metal3 s 7282 37857 7380 37955 4 vdd
rlabel metal3 s 6850 48917 6948 49015 4 vdd
rlabel metal3 s 6850 37499 6948 37597 4 vdd
rlabel metal3 s 8060 63941 8158 64039 4 vdd
rlabel metal3 s 7282 51287 7380 51385 4 vdd
rlabel metal3 s 7282 73407 7380 73505 4 vdd
rlabel metal3 s 6850 13367 6948 13465 4 vdd
rlabel metal3 s 8060 3111 8158 3209 4 vdd
rlabel metal3 s 8060 40241 8158 40339 4 vdd
rlabel metal3 s 6850 29957 6948 30055 4 vdd
rlabel metal3 s 7282 10997 7380 11095 4 vdd
rlabel metal3 s 8060 16146 8158 16244 4 vdd
rlabel metal3 s 6850 80949 6948 81047 4 vdd
rlabel metal3 s 7282 83677 7380 83775 4 vdd
rlabel metal3 s 7282 91577 7380 91675 4 vdd
rlabel metal3 s 7282 77357 7380 77455 4 vdd
rlabel metal3 s 6850 35919 6948 36017 4 vdd
rlabel metal3 s 6850 60767 6948 60865 4 vdd
rlabel metal3 s 6850 44967 6948 45065 4 vdd
rlabel metal3 s 7282 39079 7380 39177 4 vdd
rlabel metal3 s 7282 30389 7380 30487 4 vdd
rlabel metal3 s 8060 62756 8158 62854 4 vdd
rlabel metal3 s 7282 77789 7380 77887 4 vdd
rlabel metal3 s 8060 28391 8158 28489 4 vdd
rlabel metal3 s 7282 11429 7380 11527 4 vdd
rlabel metal3 s 8060 10221 8158 10319 4 vdd
rlabel metal3 s 8060 741 8158 839 4 vdd
rlabel metal3 s 8060 22861 8158 22959 4 vdd
rlabel metal3 s 7282 67519 7380 67617 4 vdd
rlabel metal3 s 8060 35106 8158 35204 4 vdd
rlabel metal3 s 6850 41807 6948 41905 4 vdd
rlabel metal3 s 6850 78579 6948 78677 4 vdd
rlabel metal3 s 8060 95146 8158 95244 4 vdd
rlabel metal3 s 8060 88431 8158 88529 4 vdd
rlabel metal3 s 6850 46547 6948 46645 4 vdd
rlabel metal3 s 8060 46956 8158 47054 4 vdd
rlabel metal3 s 7282 26007 7380 26105 4 vdd
rlabel metal3 s 6850 78147 6948 78245 4 vdd
rlabel metal3 s 6850 68667 6948 68765 4 vdd
rlabel metal3 s 4326 4296 4424 4394 4 vdd
rlabel metal3 s 7282 94737 7380 94835 4 vdd
rlabel metal3 s 6850 100699 6948 100797 4 vdd
rlabel metal3 s 7282 100267 7380 100365 4 vdd
rlabel metal3 s 6850 23279 6948 23377 4 vdd
rlabel metal3 s 6850 69457 6948 69555 4 vdd
rlabel metal3 s 7282 59619 7380 59717 4 vdd
rlabel metal3 s 7282 57249 7380 57347 4 vdd
rlabel metal3 s 8060 65521 8158 65619 4 vdd
rlabel metal3 s 8060 52881 8158 52979 4 vdd
rlabel metal3 s 6850 59187 6948 59285 4 vdd
rlabel metal3 s 6850 29599 6948 29697 4 vdd
rlabel metal3 s 7282 75777 7380 75875 4 vdd
rlabel metal3 s 7282 29957 7380 30055 4 vdd
rlabel metal3 s 7282 13009 7380 13107 4 vdd
rlabel metal3 s 8060 50511 8158 50609 4 vdd
rlabel metal3 s 8060 346 8158 444 4 vdd
rlabel metal3 s 8060 12986 8158 13084 4 vdd
rlabel metal3 s 8060 14171 8158 14269 4 vdd
rlabel metal3 s 6850 74197 6948 74295 4 vdd
rlabel metal3 s 7282 8627 7380 8725 4 vdd
rlabel metal3 s 6850 65939 6948 66037 4 vdd
rlabel metal3 s 8060 48536 8158 48634 4 vdd
rlabel metal3 s 7282 12219 7380 12317 4 vdd
rlabel metal3 s 7282 29167 7380 29265 4 vdd
rlabel metal3 s 8060 73026 8158 73124 4 vdd
rlabel metal3 s 6850 30747 6948 30845 4 vdd
rlabel metal3 s 6850 97539 6948 97637 4 vdd
rlabel metal3 s 7282 28019 7380 28117 4 vdd
rlabel metal3 s 8060 1531 8158 1629 4 vdd
rlabel metal3 s 7282 15379 7380 15477 4 vdd
rlabel metal3 s 7282 33549 7380 33647 4 vdd
rlabel metal3 s 8060 2321 8158 2419 4 vdd
rlabel metal3 s 6850 7837 6948 7935 4 vdd
rlabel metal3 s 3548 5109 3646 5207 4 vdd
rlabel metal3 s 8060 73421 8158 73519 4 vdd
rlabel metal3 s 7282 75419 7380 75517 4 vdd
rlabel metal3 s 7282 82097 7380 82195 4 vdd
rlabel metal3 s 7282 27587 7380 27685 4 vdd
rlabel metal3 s 6850 46979 6948 47077 4 vdd
rlabel metal3 s 6850 67877 6948 67975 4 vdd
rlabel metal3 s 7282 6689 7380 6787 4 vdd
rlabel metal3 s 6850 81739 6948 81837 4 vdd
rlabel metal3 s 8060 13776 8158 13874 4 vdd
rlabel metal3 s 6850 10639 6948 10737 4 vdd
rlabel metal3 s 6850 85689 6948 85787 4 vdd
rlabel metal3 s 7282 25649 7380 25747 4 vdd
rlabel metal3 s 7282 17317 7380 17415 4 vdd
rlabel metal3 s 7282 14157 7380 14255 4 vdd
rlabel metal3 s 6850 30389 6948 30487 4 vdd
rlabel metal3 s 6850 79369 6948 79467 4 vdd
rlabel metal3 s 6850 75777 6948 75875 4 vdd
rlabel metal3 s 8060 22071 8158 22169 4 vdd
rlabel metal3 s 8060 31551 8158 31649 4 vdd
rlabel metal3 s 6850 25217 6948 25315 4 vdd
rlabel metal3 s 8060 79741 8158 79839 4 vdd
rlabel metal3 s 6850 74987 6948 75085 4 vdd
rlabel metal3 s 6850 98687 6948 98785 4 vdd
rlabel metal3 s 7282 92367 7380 92465 4 vdd
rlabel metal3 s 8060 13381 8158 13479 4 vdd
rlabel metal3 s 7282 89639 7380 89737 4 vdd
rlabel metal3 s 8060 29181 8158 29279 4 vdd
rlabel metal3 s 7282 32327 7380 32425 4 vdd
rlabel metal3 s 6850 12219 6948 12317 4 vdd
rlabel metal3 s 7282 93589 7380 93687 4 vdd
rlabel metal3 s 8060 100281 8158 100379 4 vdd
rlabel metal3 s 7282 74629 7380 74727 4 vdd
rlabel metal3 s 8060 69471 8158 69569 4 vdd
rlabel metal3 s 7282 88417 7380 88515 4 vdd
rlabel metal3 s 8060 39451 8158 39549 4 vdd
rlabel metal3 s 7282 58829 7380 58927 4 vdd
rlabel metal3 s 8060 43796 8158 43894 4 vdd
rlabel metal3 s 7282 99119 7380 99217 4 vdd
rlabel metal3 s 3116 3529 3214 3627 4 vdd
rlabel metal3 s 8060 47351 8158 47449 4 vdd
rlabel metal3 s 6850 45399 6948 45497 4 vdd
rlabel metal3 s 7282 88059 7380 88157 4 vdd
rlabel metal3 s 8060 76976 8158 77074 4 vdd
rlabel metal3 s 7282 97897 7380 97995 4 vdd
rlabel metal3 s 7282 54089 7380 54187 4 vdd
rlabel metal3 s 6850 13799 6948 13897 4 vdd
rlabel metal3 s 6850 33117 6948 33215 4 vdd
rlabel metal3 s 7282 74197 7380 74295 4 vdd
rlabel metal3 s 8060 70656 8158 70754 4 vdd
rlabel metal3 s 8060 74211 8158 74309 4 vdd
rlabel metal3 s 6850 3097 6948 3195 4 vdd
rlabel metal3 s 6850 62779 6948 62877 4 vdd
rlabel metal3 s 7282 65507 7380 65605 4 vdd
rlabel metal3 s 8060 75396 8158 75494 4 vdd
rlabel metal3 s 6850 29167 6948 29265 4 vdd
rlabel metal3 s 7282 43387 7380 43485 4 vdd
rlabel metal3 s 7282 46547 7380 46645 4 vdd
rlabel metal3 s 7282 25217 7380 25315 4 vdd
rlabel metal3 s 8060 88036 8158 88134 4 vdd
rlabel metal3 s 7282 20119 7380 20217 4 vdd
rlabel metal3 s 8060 92381 8158 92479 4 vdd
rlabel metal3 s 7282 80159 7380 80257 4 vdd
rlabel metal3 s 8060 45376 8158 45474 4 vdd
rlabel metal3 s 8060 47746 8158 47844 4 vdd
rlabel metal3 s 7282 20477 7380 20575 4 vdd
rlabel metal3 s 3116 5109 3214 5207 4 vdd
rlabel metal3 s 7282 48127 7380 48225 4 vdd
rlabel metal3 s 8060 17331 8158 17429 4 vdd
rlabel metal3 s 6850 74629 6948 74727 4 vdd
rlabel metal3 s 6850 99909 6948 100007 4 vdd
rlabel metal3 s 8060 97121 8158 97219 4 vdd
rlabel metal3 s 8060 99886 8158 99984 4 vdd
rlabel metal3 s 7282 2739 7380 2837 4 vdd
rlabel metal3 s 4326 3506 4424 3604 4 vdd
rlabel metal3 s 8060 5481 8158 5579 4 vdd
rlabel metal3 s 8060 84481 8158 84579 4 vdd
rlabel metal3 s 8060 78951 8158 79049 4 vdd
rlabel metal3 s 8060 95936 8158 96034 4 vdd
rlabel metal3 s 3551 353 3649 451 4 vdd
rlabel metal3 s 7282 7479 7380 7577 4 vdd
rlabel metal3 s 6850 55669 6948 55767 4 vdd
rlabel metal3 s 6850 69099 6948 69197 4 vdd
rlabel metal3 s 8060 68286 8158 68384 4 vdd
rlabel metal3 s 6850 52077 6948 52175 4 vdd
rlabel metal3 s 8060 56831 8158 56929 4 vdd
rlabel metal3 s 4326 5086 4424 5184 4 vdd
rlabel metal3 s 8060 32736 8158 32834 4 vdd
rlabel metal3 s 8060 25626 8158 25724 4 vdd
rlabel metal3 s 6850 92009 6948 92107 4 vdd
rlabel metal3 s 8060 26811 8158 26909 4 vdd
rlabel metal3 s 6850 71469 6948 71567 4 vdd
rlabel metal3 s 6850 72259 6948 72357 4 vdd
rlabel metal3 s 7282 33907 7380 34005 4 vdd
rlabel metal3 s 7282 82887 7380 82985 4 vdd
rlabel metal3 s 7282 71037 7380 71135 4 vdd
rlabel metal3 s 6850 81307 6948 81405 4 vdd
rlabel metal3 s 8060 24836 8158 24934 4 vdd
rlabel metal3 s 8060 23651 8158 23749 4 vdd
rlabel metal3 s 7282 31969 7380 32067 4 vdd
rlabel metal3 s 6850 95527 6948 95625 4 vdd
rlabel metal3 s 8060 60781 8158 60879 4 vdd
rlabel metal3 s 8060 75001 8158 75099 4 vdd
rlabel metal3 s 8060 14566 8158 14664 4 vdd
rlabel metal3 s 6850 71037 6948 71135 4 vdd
rlabel metal3 s 7282 82529 7380 82627 4 vdd
rlabel metal3 s 6850 52867 6948 52965 4 vdd
rlabel metal3 s 6850 5109 6948 5207 4 vdd
rlabel metal3 s 8060 23256 8158 23354 4 vdd
rlabel metal3 s 6850 18897 6948 18995 4 vdd
rlabel metal3 s 7282 68309 7380 68407 4 vdd
rlabel metal3 s 8060 59991 8158 60089 4 vdd
rlabel metal3 s 8060 89221 8158 89319 4 vdd
rlabel metal3 s 7282 45399 7380 45497 4 vdd
rlabel metal3 s 6850 80159 6948 80257 4 vdd
rlabel metal3 s 8060 27206 8158 27304 4 vdd
rlabel metal3 s 8060 84086 8158 84184 4 vdd
rlabel metal3 s 8060 9036 8158 9134 4 vdd
rlabel metal3 s 6850 90429 6948 90527 4 vdd
rlabel metal3 s 7282 79727 7380 79825 4 vdd
rlabel metal3 s 6850 87269 6948 87367 4 vdd
rlabel metal3 s 8060 82901 8158 82999 4 vdd
rlabel metal3 s 6850 95959 6948 96057 4 vdd
rlabel metal3 s 1632 6666 1730 6764 4 vdd
rlabel metal3 s 8060 96726 8158 96824 4 vdd
rlabel metal3 s 7282 49707 7380 49805 4 vdd
rlabel metal3 s 8060 83296 8158 83394 4 vdd
rlabel metal3 s 7282 31537 7380 31635 4 vdd
rlabel metal3 s 6850 57607 6948 57705 4 vdd
rlabel metal3 s 8060 33131 8158 33229 4 vdd
rlabel metal3 s 8060 76186 8158 76284 4 vdd
rlabel metal3 s 7282 42239 7380 42337 4 vdd
rlabel metal3 s 7282 24069 7380 24167 4 vdd
rlabel metal3 s 6850 11429 6948 11527 4 vdd
rlabel metal3 s 7282 64717 7380 64815 4 vdd
rlabel metal3 s 6850 50139 6948 50237 4 vdd
rlabel metal3 s 6850 9849 6948 9947 4 vdd
rlabel metal3 s 6850 54089 6948 54187 4 vdd
rlabel metal3 s 8060 7456 8158 7554 4 vdd
rlabel metal3 s 7282 91219 7380 91317 4 vdd
rlabel metal3 s 8060 60386 8158 60484 4 vdd
rlabel metal3 s 7282 45757 7380 45855 4 vdd
rlabel metal3 s 4326 2716 4424 2814 4 vdd
rlabel metal3 s 6850 55237 6948 55335 4 vdd
rlabel metal3 s 8060 40636 8158 40734 4 vdd
rlabel metal3 s 8060 15356 8158 15454 4 vdd
rlabel metal3 s 8060 29971 8158 30069 4 vdd
rlabel metal3 s 3551 1143 3649 1241 4 vdd
rlabel metal3 s 3548 3529 3646 3627 4 vdd
rlabel metal3 s 8060 82506 8158 82604 4 vdd
rlabel metal3 s 6850 2739 6948 2837 4 vdd
rlabel metal3 s 7282 78579 7380 78677 4 vdd
rlabel metal3 s 6850 86047 6948 86145 4 vdd
rlabel metal3 s 6850 45757 6948 45855 4 vdd
rlabel metal3 s 6850 28377 6948 28475 4 vdd
rlabel metal3 s 3116 2739 3214 2837 4 vdd
rlabel metal3 s 6850 88417 6948 88515 4 vdd
rlabel metal3 s 8060 7851 8158 7949 4 vdd
rlabel metal3 s 6850 16169 6948 16267 4 vdd
rlabel metal3 s 8060 20096 8158 20194 4 vdd
rlabel metal3 s 7282 85689 7380 85787 4 vdd
rlabel metal3 s 7282 95959 7380 96057 4 vdd
rlabel metal3 s 6850 84109 6948 84207 4 vdd
rlabel metal3 s 6850 82097 6948 82195 4 vdd
rlabel metal3 s 7282 97107 7380 97205 4 vdd
rlabel metal3 s 8060 61966 8158 62064 4 vdd
rlabel metal3 s 7282 41449 7380 41547 4 vdd
rlabel metal3 s 8060 97911 8158 98009 4 vdd
rlabel metal3 s 7282 16169 7380 16267 4 vdd
rlabel metal3 s 8060 61571 8158 61669 4 vdd
rlabel metal3 s 8060 92776 8158 92874 4 vdd
rlabel metal3 s 7282 59187 7380 59285 4 vdd
rlabel metal3 s 7282 63137 7380 63235 4 vdd
rlabel metal3 s 6850 84467 6948 84565 4 vdd
rlabel metal3 s 6850 26797 6948 26895 4 vdd
rlabel metal3 s 7282 76999 7380 77097 4 vdd
rlabel metal3 s 8060 87641 8158 87739 4 vdd
rlabel metal3 s 6850 70247 6948 70345 4 vdd
rlabel metal3 s 6850 46189 6948 46287 4 vdd
rlabel metal3 s 6850 19329 6948 19427 4 vdd
rlabel metal3 s 6850 57249 6948 57347 4 vdd
rlabel metal3 s 6850 15379 6948 15477 4 vdd
rlabel metal3 s 6850 16527 6948 16625 4 vdd
rlabel metal3 s 6850 1949 6948 2047 4 vdd
rlabel metal3 s 6850 727 6948 825 4 vdd
rlabel metal3 s 8060 1136 8158 1234 4 vdd
rlabel metal3 s 7282 40659 7380 40757 4 vdd
rlabel metal3 s 8060 9826 8158 9924 4 vdd
rlabel metal3 s 3548 2739 3646 2837 4 vdd
rlabel metal3 s 7282 72617 7380 72715 4 vdd
rlabel metal3 s 8060 33921 8158 34019 4 vdd
rlabel metal3 s 8060 26021 8158 26119 4 vdd
rlabel metal3 s 6850 70679 6948 70777 4 vdd
rlabel metal3 s 7282 37499 7380 37597 4 vdd
rlabel metal3 s 8060 43006 8158 43104 4 vdd
rlabel metal3 s 7282 9417 7380 9515 4 vdd
rlabel metal3 s 8060 30761 8158 30859 4 vdd
rlabel metal3 s 7282 52509 7380 52607 4 vdd
rlabel metal3 s 7282 80517 7380 80615 4 vdd
rlabel metal3 s 6850 39437 6948 39535 4 vdd
rlabel metal3 s 6850 56027 6948 56125 4 vdd
rlabel metal3 s 8060 52091 8158 52189 4 vdd
rlabel metal3 s 8060 37476 8158 37574 4 vdd
rlabel metal3 s 7282 66729 7380 66827 4 vdd
rlabel metal3 s 7282 35919 7380 36017 4 vdd
rlabel metal3 s 7282 69099 7380 69197 4 vdd
rlabel metal3 s 8060 27996 8158 28094 4 vdd
rlabel metal3 s 6850 31179 6948 31277 4 vdd
rlabel metal3 s 6850 35487 6948 35585 4 vdd
rlabel metal3 s 6850 75419 6948 75517 4 vdd
rlabel metal3 s 8060 63546 8158 63644 4 vdd
rlabel metal3 s 3116 7479 3214 7577 4 vdd
rlabel metal3 s 7282 73839 7380 73937 4 vdd
rlabel metal3 s 6850 33907 6948 34005 4 vdd
rlabel metal3 s 6850 92367 6948 92465 4 vdd
rlabel metal3 s 8060 71051 8158 71149 4 vdd
rlabel metal3 s 8060 93566 8158 93664 4 vdd
rlabel metal3 s 7282 1159 7380 1257 4 vdd
rlabel metal3 s 8060 91591 8158 91689 4 vdd
rlabel metal3 s 6850 53657 6948 53755 4 vdd
rlabel metal3 s 6850 7047 6948 7145 4 vdd
rlabel metal3 s 7282 86479 7380 86577 4 vdd
rlabel metal3 s 8060 59201 8158 59299 4 vdd
rlabel metal3 s 8060 4691 8158 4789 4 vdd
rlabel metal3 s 8060 30366 8158 30464 4 vdd
rlabel metal3 s 8060 95541 8158 95639 4 vdd
rlabel metal3 s 7282 73049 7380 73147 4 vdd
rlabel metal3 s 6850 86479 6948 86577 4 vdd
rlabel metal3 s 8060 18911 8158 19009 4 vdd
rlabel metal3 s 6850 40659 6948 40757 4 vdd
rlabel metal3 s 8060 42611 8158 42709 4 vdd
rlabel metal3 s 7282 4319 7380 4417 4 vdd
rlabel metal3 s 6850 10207 6948 10305 4 vdd
rlabel metal3 s 7282 10207 7380 10305 4 vdd
rlabel metal3 s 7282 43029 7380 43127 4 vdd
rlabel metal3 s 7282 9059 7380 9157 4 vdd
rlabel metal3 s 6850 61557 6948 61655 4 vdd
rlabel metal3 s 6850 67519 6948 67617 4 vdd
rlabel metal3 s 7282 43819 7380 43917 4 vdd
rlabel metal3 s 8060 80531 8158 80629 4 vdd
rlabel metal3 s 6850 22057 6948 22155 4 vdd
rlabel metal3 s 6850 60409 6948 60507 4 vdd
rlabel metal3 s 6850 17317 6948 17415 4 vdd
rlabel metal3 s 6850 94379 6948 94477 4 vdd
rlabel metal3 s 8060 91196 8158 91294 4 vdd
rlabel metal3 s 8060 50116 8158 50214 4 vdd
rlabel metal3 s 7282 97539 7380 97637 4 vdd
rlabel metal3 s 2228 346 2326 444 4 vdd
rlabel metal3 s 6850 56817 6948 56915 4 vdd
rlabel metal3 s 7282 96749 7380 96847 4 vdd
rlabel metal3 s 7664 99491 7762 99589 4 gnd
rlabel metal3 s 7664 90801 7762 90899 4 gnd
rlabel metal3 s 7664 82506 7762 82604 4 gnd
rlabel metal3 s 6425 8685 6523 8783 4 gnd
rlabel metal3 s 6425 20535 6523 20633 4 gnd
rlabel metal3 s 6425 86895 6523 86993 4 gnd
rlabel metal3 s 7664 72631 7762 72729 4 gnd
rlabel metal3 s 6425 58829 6523 58927 4 gnd
rlabel metal3 s 6425 10265 6523 10363 4 gnd
rlabel metal3 s 6425 30389 6523 30487 4 gnd
rlabel metal3 s 6425 16959 6523 17057 4 gnd
rlabel metal3 s 7664 2716 7762 2814 4 gnd
rlabel metal3 s 6425 62405 6523 62503 4 gnd
rlabel metal3 s 6425 42239 6523 42337 4 gnd
rlabel metal3 s 3930 6666 4028 6764 4 gnd
rlabel metal3 s 6425 8269 6523 8367 4 gnd
rlabel metal3 s 6425 93589 6523 93687 4 gnd
rlabel metal3 s 6425 61615 6523 61713 4 gnd
rlabel metal3 s 7664 10616 7762 10714 4 gnd
rlabel metal3 s 6425 50139 6523 50237 4 gnd
rlabel metal3 s 7664 58806 7762 58904 4 gnd
rlabel metal3 s 6425 75045 6523 75143 4 gnd
rlabel metal3 s 6425 89639 6523 89737 4 gnd
rlabel metal3 s 1236 6666 1334 6764 4 gnd
rlabel metal3 s 6425 95169 6523 95267 4 gnd
rlabel metal3 s 7664 99096 7762 99194 4 gnd
rlabel metal3 s 7664 12196 7762 12294 4 gnd
rlabel metal3 s 6425 31595 6523 31693 4 gnd
rlabel metal3 s 6425 62779 6523 62877 4 gnd
rlabel metal3 s 3930 8246 4028 8344 4 gnd
rlabel metal3 s 7664 36291 7762 36389 4 gnd
rlabel metal3 s 6425 83735 6523 83833 4 gnd
rlabel metal3 s 7664 86456 7762 86554 4 gnd
rlabel metal3 s 6425 33965 6523 34063 4 gnd
rlabel metal3 s 6425 79785 6523 79883 4 gnd
rlabel metal3 s 7664 33526 7762 33624 4 gnd
rlabel metal3 s 7664 37476 7762 37574 4 gnd
rlabel metal3 s 6425 3945 6523 4043 4 gnd
rlabel metal3 s 6425 56875 6523 56973 4 gnd
rlabel metal3 s 7664 80926 7762 81024 4 gnd
rlabel metal3 s 6425 96749 6523 96847 4 gnd
rlabel metal3 s 7664 27206 7762 27304 4 gnd
rlabel metal3 s 6425 13009 6523 13107 4 gnd
rlabel metal3 s 6425 9475 6523 9573 4 gnd
rlabel metal3 s 7664 3111 7762 3209 4 gnd
rlabel metal3 s 6425 11429 6523 11527 4 gnd
rlabel metal3 s 6425 72259 6523 72357 4 gnd
rlabel metal3 s 6425 92425 6523 92523 4 gnd
rlabel metal3 s 7664 82901 7762 82999 4 gnd
rlabel metal3 s 7664 93566 7762 93664 4 gnd
rlabel metal3 s 6425 35545 6523 35643 4 gnd
rlabel metal3 s 6425 49349 6523 49447 4 gnd
rlabel metal3 s 6425 55669 6523 55767 4 gnd
rlabel metal3 s 7664 22861 7762 22959 4 gnd
rlabel metal3 s 7664 26021 7762 26119 4 gnd
rlabel metal3 s 6425 75419 6523 75517 4 gnd
rlabel metal3 s 7664 11406 7762 11504 4 gnd
rlabel metal3 s 6425 1575 6523 1673 4 gnd
rlabel metal3 s 6425 52135 6523 52233 4 gnd
rlabel metal3 s 6425 84525 6523 84623 4 gnd
rlabel metal3 s 6425 34339 6523 34437 4 gnd
rlabel metal3 s 6425 28435 6523 28533 4 gnd
rlabel metal3 s 7664 99886 7762 99984 4 gnd
rlabel metal3 s 7664 33131 7762 33229 4 gnd
rlabel metal3 s 6425 52509 6523 52607 4 gnd
rlabel metal3 s 6425 34755 6523 34853 4 gnd
rlabel metal3 s 6425 40659 6523 40757 4 gnd
rlabel metal3 s 7664 30366 7762 30464 4 gnd
rlabel metal3 s 7664 31156 7762 31254 4 gnd
rlabel metal3 s 6425 36709 6523 36807 4 gnd
rlabel metal3 s 7664 43006 7762 43104 4 gnd
rlabel metal3 s 7664 7851 7762 7949 4 gnd
rlabel metal3 s 7664 12986 7762 13084 4 gnd
rlabel metal3 s 6425 23279 6523 23377 4 gnd
rlabel metal3 s 6425 39869 6523 39967 4 gnd
rlabel metal3 s 6425 73465 6523 73563 4 gnd
rlabel metal3 s 7664 18911 7762 19009 4 gnd
rlabel metal3 s 6425 72675 6523 72773 4 gnd
rlabel metal3 s 6425 48559 6523 48657 4 gnd
rlabel metal3 s 7664 61176 7762 61274 4 gnd
rlabel metal3 s 6425 28809 6523 28907 4 gnd
rlabel metal3 s 6425 73049 6523 73147 4 gnd
rlabel metal3 s 6425 71885 6523 71983 4 gnd
rlabel metal3 s 6425 80949 6523 81047 4 gnd
rlabel metal3 s 6425 17375 6523 17473 4 gnd
rlabel metal3 s 6425 21699 6523 21797 4 gnd
rlabel metal3 s 7664 11801 7762 11899 4 gnd
rlabel metal3 s 7664 78161 7762 78259 4 gnd
rlabel metal3 s 7664 24441 7762 24539 4 gnd
rlabel metal3 s 7664 17726 7762 17824 4 gnd
rlabel metal3 s 7664 76186 7762 76284 4 gnd
rlabel metal3 s 7664 27996 7762 28094 4 gnd
rlabel metal3 s 6425 91219 6523 91317 4 gnd
rlabel metal3 s 7664 14961 7762 15059 4 gnd
rlabel metal3 s 7664 21676 7762 21774 4 gnd
rlabel metal3 s 6425 99119 6523 99217 4 gnd
rlabel metal3 s 6425 95959 6523 96057 4 gnd
rlabel metal3 s 2691 4319 2789 4417 4 gnd
rlabel metal3 s 6425 67935 6523 68033 4 gnd
rlabel metal3 s 7664 44191 7762 44289 4 gnd
rlabel metal3 s 7664 41821 7762 41919 4 gnd
rlabel metal3 s 7664 56831 7762 56929 4 gnd
rlabel metal3 s 6425 64775 6523 64873 4 gnd
rlabel metal3 s 6425 22115 6523 22213 4 gnd
rlabel metal3 s 6425 88849 6523 88947 4 gnd
rlabel metal3 s 7664 77371 7762 77469 4 gnd
rlabel metal3 s 6425 41449 6523 41547 4 gnd
rlabel metal3 s 3930 346 4028 444 4 gnd
rlabel metal3 s 7664 53276 7762 53374 4 gnd
rlabel metal3 s 6425 45399 6523 45497 4 gnd
rlabel metal3 s 6425 1949 6523 2047 4 gnd
rlabel metal3 s 7664 53671 7762 53769 4 gnd
rlabel metal3 s 6425 35919 6523 36017 4 gnd
rlabel metal3 s 6425 55295 6523 55393 4 gnd
rlabel metal3 s 7664 67496 7762 67594 4 gnd
rlabel metal3 s 7664 73816 7762 73914 4 gnd
rlabel metal3 s 7664 10221 7762 10319 4 gnd
rlabel metal3 s 6425 98745 6523 98843 4 gnd
rlabel metal3 s 6425 73839 6523 73937 4 gnd
rlabel metal3 s 6425 57249 6523 57347 4 gnd
rlabel metal3 s 7664 46166 7762 46264 4 gnd
rlabel metal3 s 7664 16146 7762 16244 4 gnd
rlabel metal3 s 6425 29225 6523 29323 4 gnd
rlabel metal3 s 6425 45815 6523 45913 4 gnd
rlabel metal3 s 6425 70305 6523 70403 4 gnd
rlabel metal3 s 6425 91635 6523 91733 4 gnd
rlabel metal3 s 7664 5876 7762 5974 4 gnd
rlabel metal3 s 7664 44586 7762 44684 4 gnd
rlabel metal3 s 7664 38266 7762 38364 4 gnd
rlabel metal3 s 6425 99909 6523 100007 4 gnd
rlabel metal3 s 7664 78556 7762 78654 4 gnd
rlabel metal3 s 6425 13425 6523 13523 4 gnd
rlabel metal3 s 7664 79741 7762 79839 4 gnd
rlabel metal3 s 6425 95585 6523 95683 4 gnd
rlabel metal3 s 6425 10639 6523 10737 4 gnd
rlabel metal3 s 7664 32736 7762 32834 4 gnd
rlabel metal3 s 7664 50511 7762 50609 4 gnd
rlabel metal3 s 6425 88059 6523 88157 4 gnd
rlabel metal3 s 7664 64731 7762 64829 4 gnd
rlabel metal3 s 7664 91591 7762 91689 4 gnd
rlabel metal3 s 7664 48931 7762 49029 4 gnd
rlabel metal3 s 7664 9826 7762 9924 4 gnd
rlabel metal3 s 6425 44235 6523 44333 4 gnd
rlabel metal3 s 7664 90011 7762 90109 4 gnd
rlabel metal3 s 7664 55251 7762 55349 4 gnd
rlabel metal3 s 7664 89616 7762 89714 4 gnd
rlabel metal3 s 6425 4735 6523 4833 4 gnd
rlabel metal3 s 6425 25649 6523 25747 4 gnd
rlabel metal3 s 7664 52091 7762 52189 4 gnd
rlabel metal3 s 7664 61571 7762 61669 4 gnd
rlabel metal3 s 7664 47746 7762 47844 4 gnd
rlabel metal3 s 7664 56041 7762 56139 4 gnd
rlabel metal3 s 7664 23256 7762 23354 4 gnd
rlabel metal3 s 6425 43445 6523 43543 4 gnd
rlabel metal3 s 7664 95541 7762 95639 4 gnd
rlabel metal3 s 7664 33921 7762 34019 4 gnd
rlabel metal3 s 6425 2739 6523 2837 4 gnd
rlabel metal3 s 6425 30805 6523 30903 4 gnd
rlabel metal3 s 7664 60386 7762 60484 4 gnd
rlabel metal3 s 7664 20096 7762 20194 4 gnd
rlabel metal3 s 6425 48185 6523 48283 4 gnd
rlabel metal3 s 7664 58411 7762 58509 4 gnd
rlabel metal3 s 7664 68681 7762 68779 4 gnd
rlabel metal3 s 6425 7479 6523 7577 4 gnd
rlabel metal3 s 7664 20886 7762 20984 4 gnd
rlabel metal3 s 7664 17331 7762 17429 4 gnd
rlabel metal3 s 7664 90406 7762 90504 4 gnd
rlabel metal3 s 6425 51345 6523 51443 4 gnd
rlabel metal3 s 6425 64359 6523 64457 4 gnd
rlabel metal3 s 3930 4296 4028 4394 4 gnd
rlabel metal3 s 6425 68309 6523 68407 4 gnd
rlabel metal3 s 6425 92799 6523 92897 4 gnd
rlabel metal3 s 6425 14215 6523 14313 4 gnd
rlabel metal3 s 7664 30761 7762 30859 4 gnd
rlabel metal3 s 7664 79346 7762 79444 4 gnd
rlabel metal3 s 7664 84086 7762 84184 4 gnd
rlabel metal3 s 7664 67101 7762 67199 4 gnd
rlabel metal3 s 6425 54879 6523 54977 4 gnd
rlabel metal3 s 2691 2739 2789 2837 4 gnd
rlabel metal3 s 7664 62756 7762 62854 4 gnd
rlabel metal3 s 7664 69076 7762 69174 4 gnd
rlabel metal3 s 6425 94795 6523 94893 4 gnd
rlabel metal3 s 2691 3529 2789 3627 4 gnd
rlabel metal3 s 7664 66311 7762 66409 4 gnd
rlabel metal3 s 6425 85689 6523 85787 4 gnd
rlabel metal3 s 7664 51696 7762 51794 4 gnd
rlabel metal3 s 7664 50116 7762 50214 4 gnd
rlabel metal3 s 7664 76976 7762 77074 4 gnd
rlabel metal3 s 6425 21325 6523 21423 4 gnd
rlabel metal3 s 6425 38705 6523 38803 4 gnd
rlabel metal3 s 7664 24046 7762 24144 4 gnd
rlabel metal3 s 6425 14589 6523 14687 4 gnd
rlabel metal3 s 6425 785 6523 883 4 gnd
rlabel metal3 s 6425 5899 6523 5997 4 gnd
rlabel metal3 s 6425 69099 6523 69197 4 gnd
rlabel metal3 s 7664 78951 7762 79049 4 gnd
rlabel metal3 s 7664 44981 7762 45079 4 gnd
rlabel metal3 s 7664 50906 7762 51004 4 gnd
rlabel metal3 s 6425 60825 6523 60923 4 gnd
rlabel metal3 s 7664 95146 7762 95244 4 gnd
rlabel metal3 s 6425 32759 6523 32857 4 gnd
rlabel metal3 s 6425 48975 6523 49073 4 gnd
rlabel metal3 s 7664 11011 7762 11109 4 gnd
rlabel metal3 s 7664 49326 7762 49424 4 gnd
rlabel metal3 s 6425 30015 6523 30113 4 gnd
rlabel metal3 s 6425 51719 6523 51817 4 gnd
rlabel metal3 s 3930 3506 4028 3604 4 gnd
rlabel metal3 s 7664 85666 7762 85764 4 gnd
rlabel metal3 s 6425 58039 6523 58137 4 gnd
rlabel metal3 s 6425 86479 6523 86577 4 gnd
rlabel metal3 s 6425 22489 6523 22587 4 gnd
rlabel metal3 s 7664 21281 7762 21379 4 gnd
rlabel metal3 s 6425 13799 6523 13897 4 gnd
rlabel metal3 s 7664 75001 7762 75099 4 gnd
rlabel metal3 s 7664 45376 7762 45474 4 gnd
rlabel metal3 s 6425 2365 6523 2463 4 gnd
rlabel metal3 s 7664 39846 7762 39944 4 gnd
rlabel metal3 s 6425 65939 6523 66037 4 gnd
rlabel metal3 s 6425 33175 6523 33273 4 gnd
rlabel metal3 s 7664 88826 7762 88924 4 gnd
rlabel metal3 s 6425 69889 6523 69987 4 gnd
rlabel metal3 s 7664 59596 7762 59694 4 gnd
rlabel metal3 s 7664 14566 7762 14664 4 gnd
rlabel metal3 s 6425 92009 6523 92107 4 gnd
rlabel metal3 s 6425 61989 6523 62087 4 gnd
rlabel metal3 s 6425 90429 6523 90527 4 gnd
rlabel metal3 s 6425 59619 6523 59717 4 gnd
rlabel metal3 s 6425 43029 6523 43127 4 gnd
rlabel metal3 s 6425 4319 6523 4417 4 gnd
rlabel metal3 s 7664 7061 7762 7159 4 gnd
rlabel metal3 s 7664 71446 7762 71544 4 gnd
rlabel metal3 s 7664 94356 7762 94454 4 gnd
rlabel metal3 s 6425 41865 6523 41963 4 gnd
rlabel metal3 s 6425 16169 6523 16267 4 gnd
rlabel metal3 s 7664 15751 7762 15849 4 gnd
rlabel metal3 s 7664 73026 7762 73124 4 gnd
rlabel metal3 s 7664 81716 7762 81814 4 gnd
rlabel metal3 s 6425 75835 6523 75933 4 gnd
rlabel metal3 s 6425 40285 6523 40383 4 gnd
rlabel metal3 s 6425 49765 6523 49863 4 gnd
rlabel metal3 s 6425 63569 6523 63667 4 gnd
rlabel metal3 s 7664 74606 7762 74704 4 gnd
rlabel metal3 s 7664 45771 7762 45869 4 gnd
rlabel metal3 s 6425 36335 6523 36433 4 gnd
rlabel metal3 s 6425 53299 6523 53397 4 gnd
rlabel metal3 s 7664 96331 7762 96429 4 gnd
rlabel metal3 s 6425 100325 6523 100423 4 gnd
rlabel metal3 s 3930 2716 4028 2814 4 gnd
rlabel metal3 s 6425 97165 6523 97263 4 gnd
rlabel metal3 s 7664 1531 7762 1629 4 gnd
rlabel metal3 s 6425 50555 6523 50653 4 gnd
rlabel metal3 s 7664 65126 7762 65224 4 gnd
rlabel metal3 s 7664 29181 7762 29279 4 gnd
rlabel metal3 s 6425 15795 6523 15893 4 gnd
rlabel metal3 s 6425 76209 6523 76307 4 gnd
rlabel metal3 s 7664 37871 7762 37969 4 gnd
rlabel metal3 s 6425 15379 6523 15477 4 gnd
rlabel metal3 s 6425 37125 6523 37223 4 gnd
rlabel metal3 s 7664 35501 7762 35599 4 gnd
rlabel metal3 s 6425 65149 6523 65247 4 gnd
rlabel metal3 s 7664 94751 7762 94849 4 gnd
rlabel metal3 s 6425 71095 6523 71193 4 gnd
rlabel metal3 s 7664 86061 7762 86159 4 gnd
rlabel metal3 s 7664 92381 7762 92479 4 gnd
rlabel metal3 s 6425 74629 6523 74727 4 gnd
rlabel metal3 s 6425 94005 6523 94103 4 gnd
rlabel metal3 s 6425 67145 6523 67243 4 gnd
rlabel metal3 s 7664 5086 7762 5184 4 gnd
rlabel metal3 s 7664 67891 7762 67989 4 gnd
rlabel metal3 s 7664 71051 7762 71149 4 gnd
rlabel metal3 s 7664 84876 7762 84974 4 gnd
rlabel metal3 s 6425 3529 6523 3627 4 gnd
rlabel metal3 s 6425 41075 6523 41173 4 gnd
rlabel metal3 s 7664 98701 7762 98799 4 gnd
rlabel metal3 s 6425 31969 6523 32067 4 gnd
rlabel metal3 s 7664 31551 7762 31649 4 gnd
rlabel metal3 s 6425 59245 6523 59343 4 gnd
rlabel metal3 s 7664 76581 7762 76679 4 gnd
rlabel metal3 s 7664 82111 7762 82209 4 gnd
rlabel metal3 s 7664 4296 7762 4394 4 gnd
rlabel metal3 s 7664 65521 7762 65619 4 gnd
rlabel metal3 s 2691 8269 2789 8367 4 gnd
rlabel metal3 s 6425 20119 6523 20217 4 gnd
rlabel metal3 s 6425 84109 6523 84207 4 gnd
rlabel metal3 s 6425 29599 6523 29697 4 gnd
rlabel metal3 s 2691 9059 2789 9157 4 gnd
rlabel metal3 s 6425 89265 6523 89363 4 gnd
rlabel metal3 s 7664 26811 7762 26909 4 gnd
rlabel metal3 s 6425 97955 6523 98053 4 gnd
rlabel metal3 s 6425 52925 6523 53023 4 gnd
rlabel metal3 s 6425 26439 6523 26537 4 gnd
rlabel metal3 s 2691 5109 2789 5207 4 gnd
rlabel metal3 s 6425 78205 6523 78303 4 gnd
rlabel metal3 s 6425 99535 6523 99633 4 gnd
rlabel metal3 s 6425 78579 6523 78677 4 gnd
rlabel metal3 s 6425 58455 6523 58553 4 gnd
rlabel metal3 s 7664 69866 7762 69964 4 gnd
rlabel metal3 s 7664 75791 7762 75889 4 gnd
rlabel metal3 s 6425 88475 6523 88573 4 gnd
rlabel metal3 s 6425 45025 6523 45123 4 gnd
rlabel metal3 s 6425 86105 6523 86203 4 gnd
rlabel metal3 s 7664 65916 7762 66014 4 gnd
rlabel metal3 s 6425 90055 6523 90153 4 gnd
rlabel metal3 s 1236 2716 1334 2814 4 gnd
rlabel metal3 s 7664 75396 7762 75494 4 gnd
rlabel metal3 s 7664 64336 7762 64434 4 gnd
rlabel metal3 s 7664 97121 7762 97219 4 gnd
rlabel metal3 s 6425 39495 6523 39593 4 gnd
rlabel metal3 s 7664 7456 7762 7554 4 gnd
rlabel metal3 s 7664 100281 7762 100379 4 gnd
rlabel metal3 s 9960 50511 10058 50609 4 gnd
rlabel metal3 s 6425 77415 6523 77513 4 gnd
rlabel metal3 s 7664 93171 7762 93269 4 gnd
rlabel metal3 s 6425 24069 6523 24167 4 gnd
rlabel metal3 s 6425 63195 6523 63293 4 gnd
rlabel metal3 s 7664 93961 7762 94059 4 gnd
rlabel metal3 s 6425 1159 6523 1257 4 gnd
rlabel metal3 s 7664 28786 7762 28884 4 gnd
rlabel metal3 s 7664 87246 7762 87344 4 gnd
rlabel metal3 s 6425 87269 6523 87367 4 gnd
rlabel metal3 s 6425 87685 6523 87783 4 gnd
rlabel metal3 s 6425 46189 6523 46287 4 gnd
rlabel metal3 s 6425 98329 6523 98427 4 gnd
rlabel metal3 s 1832 346 1930 444 4 gnd
rlabel metal3 s 6425 100699 6523 100797 4 gnd
rlabel metal3 s 7664 13776 7762 13874 4 gnd
rlabel metal3 s 7664 73421 7762 73519 4 gnd
rlabel metal3 s 7664 38661 7762 38759 4 gnd
rlabel metal3 s 6425 76625 6523 76723 4 gnd
rlabel metal3 s 6425 90845 6523 90943 4 gnd
rlabel metal3 s 6425 85315 6523 85413 4 gnd
rlabel metal3 s 6425 5525 6523 5623 4 gnd
rlabel metal3 s 6425 3155 6523 3253 4 gnd
rlabel metal3 s 6425 82529 6523 82627 4 gnd
rlabel metal3 s 7664 72236 7762 72334 4 gnd
rlabel metal3 s 6425 18955 6523 19053 4 gnd
rlabel metal3 s 7664 14171 7762 14269 4 gnd
rlabel metal3 s 6425 9849 6523 9947 4 gnd
rlabel metal3 s 7664 51301 7762 51399 4 gnd
rlabel metal3 s 7664 91196 7762 91294 4 gnd
rlabel metal3 s 7664 41031 7762 41129 4 gnd
rlabel metal3 s 6425 16585 6523 16683 4 gnd
rlabel metal3 s 6425 28019 6523 28117 4 gnd
rlabel metal3 s 7664 34711 7762 34809 4 gnd
rlabel metal3 s 6425 97539 6523 97637 4 gnd
rlabel metal3 s 6425 53715 6523 53813 4 gnd
rlabel metal3 s 6425 80159 6523 80257 4 gnd
rlabel metal3 s 7664 5481 7762 5579 4 gnd
rlabel metal3 s 7664 54461 7762 54559 4 gnd
rlabel metal3 s 6425 5109 6523 5207 4 gnd
rlabel metal3 s 6425 65565 6523 65663 4 gnd
rlabel metal3 s 7664 1136 7762 1234 4 gnd
rlabel metal3 s 7664 54856 7762 54954 4 gnd
rlabel metal3 s 7664 95936 7762 96034 4 gnd
rlabel metal3 s 6425 77789 6523 77887 4 gnd
rlabel metal3 s 6425 47769 6523 47867 4 gnd
rlabel metal3 s 8492 50496 8590 50594 4 gnd
rlabel metal3 s 6425 18165 6523 18263 4 gnd
rlabel metal3 s 7664 32341 7762 32439 4 gnd
rlabel metal3 s 6425 26065 6523 26163 4 gnd
rlabel metal3 s 7664 81321 7762 81419 4 gnd
rlabel metal3 s 6425 54505 6523 54603 4 gnd
rlabel metal3 s 7664 97911 7762 98009 4 gnd
rlabel metal3 s 6425 19745 6523 19843 4 gnd
rlabel metal3 s 6425 76999 6523 77097 4 gnd
rlabel metal3 s 7664 42216 7762 42314 4 gnd
rlabel metal3 s 7664 43796 7762 43894 4 gnd
rlabel metal3 s 6425 74255 6523 74353 4 gnd
rlabel metal3 s 3126 1143 3224 1241 4 gnd
rlabel metal3 s 7664 35106 7762 35204 4 gnd
rlabel metal3 s 7664 97516 7762 97614 4 gnd
rlabel metal3 s 7664 69471 7762 69569 4 gnd
rlabel metal3 s 7664 8246 7762 8344 4 gnd
rlabel metal3 s 6425 24485 6523 24583 4 gnd
rlabel metal3 s 6425 27229 6523 27327 4 gnd
rlabel metal3 s 7664 31946 7762 32044 4 gnd
rlabel metal3 s 6425 61199 6523 61297 4 gnd
rlabel metal3 s 7664 1926 7762 2024 4 gnd
rlabel metal3 s 7664 346 7762 444 4 gnd
rlabel metal3 s 7664 9431 7762 9529 4 gnd
rlabel metal3 s 6425 60035 6523 60133 4 gnd
rlabel metal3 s 7664 80531 7762 80629 4 gnd
rlabel metal3 s 7664 40241 7762 40339 4 gnd
rlabel metal3 s 6425 71469 6523 71567 4 gnd
rlabel metal3 s 7664 55646 7762 55744 4 gnd
rlabel metal3 s 7664 48141 7762 48239 4 gnd
rlabel metal3 s 6425 27645 6523 27743 4 gnd
rlabel metal3 s 7664 27601 7762 27699 4 gnd
rlabel metal3 s 7664 70656 7762 70754 4 gnd
rlabel metal3 s 7664 98306 7762 98404 4 gnd
rlabel metal3 s 7664 61966 7762 62064 4 gnd
rlabel metal3 s 6425 26855 6523 26953 4 gnd
rlabel metal3 s 6425 69515 6523 69613 4 gnd
rlabel metal3 s 7664 88431 7762 88529 4 gnd
rlabel metal3 s 6425 6689 6523 6787 4 gnd
rlabel metal3 s 6425 32385 6523 32483 4 gnd
rlabel metal3 s 7664 36686 7762 36784 4 gnd
rlabel metal3 s 6425 23695 6523 23793 4 gnd
rlabel metal3 s 7664 42611 7762 42709 4 gnd
rlabel metal3 s 7664 89221 7762 89319 4 gnd
rlabel metal3 s 6425 20909 6523 21007 4 gnd
rlabel metal3 s 6425 31179 6523 31277 4 gnd
rlabel metal3 s 6425 42655 6523 42753 4 gnd
rlabel metal3 s 7664 83691 7762 83789 4 gnd
rlabel metal3 s 7664 83296 7762 83394 4 gnd
rlabel metal3 s 7664 57226 7762 57324 4 gnd
rlabel metal3 s 7664 22071 7762 22169 4 gnd
rlabel metal3 s 7664 40636 7762 40734 4 gnd
rlabel metal3 s 6425 93215 6523 93313 4 gnd
rlabel metal3 s 7664 3901 7762 3999 4 gnd
rlabel metal3 s 7664 48536 7762 48634 4 gnd
rlabel metal3 s 7664 15356 7762 15454 4 gnd
rlabel metal3 s 7664 39056 7762 39154 4 gnd
rlabel metal3 s 2691 7479 2789 7577 4 gnd
rlabel metal3 s 7664 88036 7762 88134 4 gnd
rlabel metal3 s 6425 82155 6523 82253 4 gnd
rlabel metal3 s 7664 741 7762 839 4 gnd
rlabel metal3 s 6425 17749 6523 17847 4 gnd
rlabel metal3 s 6425 50929 6523 51027 4 gnd
rlabel metal3 s 7664 52486 7762 52584 4 gnd
rlabel metal3 s 7664 29576 7762 29674 4 gnd
rlabel metal3 s 6425 83319 6523 83417 4 gnd
rlabel metal3 s 6425 46605 6523 46703 4 gnd
rlabel metal3 s 6425 60409 6523 60507 4 gnd
rlabel metal3 s 7664 59991 7762 60089 4 gnd
rlabel metal3 s 7664 18516 7762 18614 4 gnd
rlabel metal3 s 7664 23651 7762 23749 4 gnd
rlabel metal3 s 7664 54066 7762 54164 4 gnd
rlabel metal3 s 7664 56436 7762 56534 4 gnd
rlabel metal3 s 7664 2321 7762 2419 4 gnd
rlabel metal3 s 7664 87641 7762 87739 4 gnd
rlabel metal3 s 7664 19701 7762 19799 4 gnd
rlabel metal3 s 7664 6271 7762 6369 4 gnd
rlabel metal3 s 7664 52881 7762 52979 4 gnd
rlabel metal3 s 6425 84899 6523 84997 4 gnd
rlabel metal3 s 7664 63151 7762 63249 4 gnd
rlabel metal3 s 7664 28391 7762 28489 4 gnd
rlabel metal3 s 7664 46561 7762 46659 4 gnd
rlabel metal3 s 6425 7105 6523 7203 4 gnd
rlabel metal3 s 7664 39451 7762 39549 4 gnd
rlabel metal3 s 6425 22905 6523 23003 4 gnd
rlabel metal3 s 7664 41426 7762 41524 4 gnd
rlabel metal3 s 6425 81739 6523 81837 4 gnd
rlabel metal3 s 7664 19306 7762 19404 4 gnd
rlabel metal3 s 6425 57665 6523 57763 4 gnd
rlabel metal3 s 7664 84481 7762 84579 4 gnd
rlabel metal3 s 6425 66355 6523 66453 4 gnd
rlabel metal3 s 7664 60781 7762 60879 4 gnd
rlabel metal3 s 6425 12635 6523 12733 4 gnd
rlabel metal3 s 7664 62361 7762 62459 4 gnd
rlabel metal3 s 7664 26416 7762 26514 4 gnd
rlabel metal3 s 7664 35896 7762 35994 4 gnd
rlabel metal3 s 6425 56459 6523 56557 4 gnd
rlabel metal3 s 7664 49721 7762 49819 4 gnd
rlabel metal3 s 6425 39079 6523 39177 4 gnd
rlabel metal3 s 7664 63546 7762 63644 4 gnd
rlabel metal3 s 7664 86851 7762 86949 4 gnd
rlabel metal3 s 6425 80575 6523 80673 4 gnd
rlabel metal3 s 7664 43401 7762 43499 4 gnd
rlabel metal3 s 7664 20491 7762 20589 4 gnd
rlabel metal3 s 6425 19329 6523 19427 4 gnd
rlabel metal3 s 2691 6689 2789 6787 4 gnd
rlabel metal3 s 7664 13381 7762 13479 4 gnd
rlabel metal3 s 7664 37081 7762 37179 4 gnd
rlabel metal3 s 7664 9036 7762 9134 4 gnd
rlabel metal3 s 7664 29971 7762 30069 4 gnd
rlabel metal3 s 7664 16936 7762 17034 4 gnd
rlabel metal3 s 7664 63941 7762 64039 4 gnd
rlabel metal3 s 7664 58016 7762 58114 4 gnd
rlabel metal3 s 6425 81365 6523 81463 4 gnd
rlabel metal3 s 7664 8641 7762 8739 4 gnd
rlabel metal3 s 3930 1136 4028 1234 4 gnd
rlabel metal3 s 7664 46956 7762 47054 4 gnd
rlabel metal3 s 7664 71841 7762 71939 4 gnd
rlabel metal3 s 3930 5086 4028 5184 4 gnd
rlabel metal3 s 7664 85271 7762 85369 4 gnd
rlabel metal3 s 7664 24836 7762 24934 4 gnd
rlabel metal3 s 6425 54089 6523 54187 4 gnd
rlabel metal3 s 6425 47395 6523 47493 4 gnd
rlabel metal3 s 7664 3506 7762 3604 4 gnd
rlabel metal3 s 7664 100676 7762 100774 4 gnd
rlabel metal3 s 7664 18121 7762 18219 4 gnd
rlabel metal3 s 3930 7456 4028 7554 4 gnd
rlabel metal3 s 6425 68725 6523 68823 4 gnd
rlabel metal3 s 6425 11055 6523 11153 4 gnd
rlabel metal3 s 7664 12591 7762 12689 4 gnd
rlabel metal3 s 6425 44609 6523 44707 4 gnd
rlabel metal3 s 6425 78995 6523 79093 4 gnd
rlabel metal3 s 6425 38289 6523 38387 4 gnd
rlabel metal3 s 7664 25626 7762 25724 4 gnd
rlabel metal3 s 6425 9059 6523 9157 4 gnd
rlabel metal3 s 6425 67519 6523 67617 4 gnd
rlabel metal3 s 6425 79369 6523 79467 4 gnd
rlabel metal3 s 6425 63985 6523 64083 4 gnd
rlabel metal3 s 7664 59201 7762 59299 4 gnd
rlabel metal3 s 6425 66729 6523 66827 4 gnd
rlabel metal3 s 6425 82945 6523 83043 4 gnd
rlabel metal3 s 7664 70261 7762 70359 4 gnd
rlabel metal3 s 7664 74211 7762 74309 4 gnd
rlabel metal3 s 7664 57621 7762 57719 4 gnd
rlabel metal3 s 6425 96375 6523 96473 4 gnd
rlabel metal3 s 6425 7895 6523 7993 4 gnd
rlabel metal3 s 7664 16541 7762 16639 4 gnd
rlabel metal3 s 6425 15005 6523 15103 4 gnd
rlabel metal3 s 7664 96726 7762 96824 4 gnd
rlabel metal3 s 6425 18539 6523 18637 4 gnd
rlabel metal3 s 6425 35129 6523 35227 4 gnd
rlabel metal3 s 6425 37499 6523 37597 4 gnd
rlabel metal3 s 6425 46979 6523 47077 4 gnd
rlabel metal3 s 6425 24859 6523 24957 4 gnd
rlabel metal3 s 6425 25275 6523 25373 4 gnd
rlabel metal3 s 6425 11845 6523 11943 4 gnd
rlabel metal3 s 7664 68286 7762 68384 4 gnd
rlabel metal3 s 6425 33549 6523 33647 4 gnd
rlabel metal3 s 7664 66706 7762 66804 4 gnd
rlabel metal3 s 6425 37915 6523 38013 4 gnd
rlabel metal3 s 7664 91986 7762 92084 4 gnd
rlabel metal3 s 7664 77766 7762 77864 4 gnd
rlabel metal3 s 6425 94379 6523 94477 4 gnd
rlabel metal3 s 7664 25231 7762 25329 4 gnd
rlabel metal3 s 6425 56085 6523 56183 4 gnd
rlabel metal3 s 6425 6315 6523 6413 4 gnd
rlabel metal3 s 7664 6666 7762 6764 4 gnd
rlabel metal3 s 7664 47351 7762 47449 4 gnd
rlabel metal3 s 7664 92776 7762 92874 4 gnd
rlabel metal3 s 3126 353 3224 451 4 gnd
rlabel metal3 s 6425 12219 6523 12317 4 gnd
rlabel metal3 s 3930 9036 4028 9134 4 gnd
rlabel metal3 s 7664 4691 7762 4789 4 gnd
rlabel metal3 s 6425 43819 6523 43917 4 gnd
rlabel metal3 s 7664 34316 7762 34414 4 gnd
rlabel metal3 s 7664 22466 7762 22564 4 gnd
rlabel metal3 s 6425 369 6523 467 4 gnd
rlabel metal3 s 7664 80136 7762 80234 4 gnd
rlabel metal3 s 6425 70679 6523 70777 4 gnd
<< properties >>
string FIXED_BBOX 0 0 12429 101148
<< end >>
