magic
tech sky130A
magscale 1 2
timestamp 1621059499
<< nwell >>
rect -101 261 314 582
rect 696 420 1118 1058
<< pwell >>
rect 29 -17 63 17
rect 698 -140 1120 410
<< nmos >>
rect 894 70 924 200
<< scnmos >>
rect 120 47 150 177
<< scpmoshvt >>
rect 120 297 150 497
<< pmoshvt >>
rect 892 639 922 839
<< ndiff >>
rect 68 165 120 177
rect 68 131 76 165
rect 110 131 120 165
rect 68 97 120 131
rect 68 63 76 97
rect 110 63 120 97
rect 68 47 120 63
rect 150 165 202 177
rect 150 131 160 165
rect 194 131 202 165
rect 150 97 202 131
rect 150 63 160 97
rect 194 63 202 97
rect 150 47 202 63
rect 836 188 894 200
rect 836 82 848 188
rect 882 82 894 188
rect 836 70 894 82
rect 924 188 982 200
rect 924 82 936 188
rect 970 82 982 188
rect 924 70 982 82
<< pdiff >>
rect 834 827 892 839
rect 834 651 846 827
rect 880 651 892 827
rect 834 639 892 651
rect 922 827 980 839
rect 922 651 934 827
rect 968 651 980 827
rect 922 639 980 651
rect 68 485 120 497
rect 68 451 76 485
rect 110 451 120 485
rect 68 417 120 451
rect 68 383 76 417
rect 110 383 120 417
rect 68 349 120 383
rect 68 315 76 349
rect 110 315 120 349
rect 68 297 120 315
rect 150 485 202 497
rect 150 451 160 485
rect 194 451 202 485
rect 150 417 202 451
rect 150 383 160 417
rect 194 383 202 417
rect 150 349 202 383
rect 150 315 160 349
rect 194 315 202 349
rect 150 297 202 315
<< ndiffc >>
rect 76 131 110 165
rect 76 63 110 97
rect 160 131 194 165
rect 160 63 194 97
rect 848 82 882 188
rect 936 82 970 188
<< pdiffc >>
rect 846 651 880 827
rect 934 651 968 827
rect 76 451 110 485
rect 76 383 110 417
rect 76 315 110 349
rect 160 451 194 485
rect 160 383 194 417
rect 160 315 194 349
<< psubdiff >>
rect 734 340 830 374
rect 988 340 1084 374
rect -64 160 14 190
rect 734 278 768 340
rect -64 81 -51 160
rect 1 81 14 160
rect -64 55 14 81
rect 1050 278 1084 340
rect 734 -70 768 -8
rect 1050 -70 1084 -8
rect 734 -104 830 -70
rect 988 -104 1084 -70
<< nsubdiff >>
rect 732 988 828 1022
rect 986 988 1082 1022
rect 732 926 766 988
rect 1048 926 1082 988
rect -64 448 14 479
rect -64 385 -51 448
rect 3 385 14 448
rect -64 336 14 385
rect 732 490 766 552
rect 1048 490 1082 552
rect 732 456 828 490
rect 986 456 1082 490
<< psubdiffcont >>
rect 830 340 988 374
rect -51 81 1 160
rect 734 -8 768 278
rect 1050 -8 1084 278
rect 830 -104 988 -70
<< nsubdiffcont >>
rect 828 988 986 1022
rect 732 552 766 926
rect -51 385 3 448
rect 1048 552 1082 926
rect 828 456 986 490
<< poly >>
rect 874 920 940 936
rect 874 886 890 920
rect 924 886 940 920
rect 874 870 940 886
rect 892 839 922 870
rect 892 608 922 639
rect 120 497 150 523
rect 874 592 940 608
rect 874 558 890 592
rect 924 558 940 592
rect 874 542 940 558
rect 120 265 150 297
rect 64 249 150 265
rect 64 215 80 249
rect 114 215 150 249
rect 64 199 150 215
rect 120 177 150 199
rect 120 21 150 47
rect 876 272 942 288
rect 876 238 892 272
rect 926 238 942 272
rect 876 222 942 238
rect 894 200 924 222
rect 894 48 924 70
rect 876 32 942 48
rect 876 -2 892 32
rect 926 -2 942 32
rect 876 -18 942 -2
<< polycont >>
rect 890 886 924 920
rect 890 558 924 592
rect 80 215 114 249
rect 892 238 926 272
rect 892 -2 926 32
<< locali >>
rect 732 988 828 1022
rect 986 988 1082 1022
rect 732 926 766 988
rect 668 780 732 798
rect 1048 926 1082 988
rect 874 886 890 920
rect 924 886 940 920
rect 846 827 880 843
rect 766 780 800 798
rect 668 694 718 780
rect 780 694 800 780
rect 668 682 732 694
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 766 682 800 694
rect 846 635 880 651
rect 934 827 968 843
rect 934 635 968 651
rect 874 558 890 592
rect 924 558 940 592
rect 68 485 110 527
rect 68 466 76 485
rect -64 451 76 466
rect -64 448 110 451
rect -64 385 -51 448
rect 3 417 110 448
rect 3 385 76 417
rect -64 383 76 385
rect -64 359 110 383
rect 68 349 110 359
rect 68 315 76 349
rect 68 299 110 315
rect 144 485 210 493
rect 144 451 160 485
rect 194 451 210 485
rect 732 490 766 552
rect 1048 490 1082 552
rect 732 456 828 490
rect 986 456 1082 490
rect 144 417 210 451
rect 144 383 160 417
rect 194 383 210 417
rect 144 349 210 383
rect 144 315 160 349
rect 194 315 210 349
rect 144 297 210 315
rect 164 263 210 297
rect 734 340 830 374
rect 988 340 1084 374
rect 734 278 768 340
rect -101 215 -98 263
rect -50 249 130 263
rect -50 215 80 249
rect 114 215 130 249
rect 164 215 246 263
rect 294 215 314 263
rect -64 165 110 181
rect 164 177 210 215
rect -64 160 76 165
rect -64 81 -51 160
rect 1 131 76 160
rect 1 97 110 131
rect 1 81 76 97
rect -64 63 76 81
rect -64 62 110 63
rect 64 17 110 62
rect 144 165 210 177
rect 144 131 160 165
rect 194 131 210 165
rect 144 97 210 131
rect 144 63 160 97
rect 194 63 210 97
rect 144 51 210 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
rect 1050 278 1084 340
rect 876 238 892 272
rect 926 238 942 272
rect 848 188 882 204
rect 848 66 882 82
rect 936 188 970 204
rect 936 66 970 82
rect 876 -2 892 32
rect 926 -2 942 32
rect 734 -70 768 -8
rect 1050 -70 1084 -8
rect 734 -104 830 -70
rect 988 -104 1084 -70
<< viali >>
rect 890 886 924 920
rect 718 694 732 780
rect 732 694 766 780
rect 766 694 780 780
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 846 651 880 827
rect 934 651 968 827
rect 890 558 924 592
rect -98 215 -50 263
rect 246 215 294 263
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 892 238 926 272
rect 848 82 882 188
rect 936 82 970 188
rect 892 -2 926 32
<< metal1 >>
rect 864 922 1234 958
rect -234 920 1234 922
rect -234 886 890 920
rect 924 886 1234 920
rect -234 880 936 886
rect -234 874 934 880
rect -234 263 -186 874
rect 840 827 886 839
rect 668 780 800 798
rect 668 760 718 780
rect 98 712 718 760
rect 98 592 146 712
rect 668 694 718 712
rect 780 760 800 780
rect 840 760 846 827
rect 780 712 846 760
rect 780 694 800 712
rect 668 682 800 694
rect 840 651 846 712
rect 880 651 886 827
rect 840 639 886 651
rect 928 827 974 839
rect 928 651 934 827
rect 968 806 974 827
rect 968 754 988 806
rect 1062 754 1068 756
rect 968 706 1068 754
rect 968 672 988 706
rect 1062 704 1068 706
rect 1120 704 1126 756
rect 968 651 974 672
rect 928 639 974 651
rect 868 592 940 604
rect -101 561 314 592
rect -101 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 314 561
rect -101 496 314 527
rect 868 558 890 592
rect 924 578 940 592
rect 1162 578 1234 886
rect 924 558 1234 578
rect 868 506 1234 558
rect 620 352 626 404
rect 678 352 684 404
rect -104 263 -44 275
rect -234 215 -98 263
rect -50 215 -44 263
rect -104 203 -44 215
rect 240 263 300 275
rect 240 215 246 263
rect 294 215 418 263
rect 240 203 300 215
rect 628 162 676 352
rect 870 306 942 506
rect 870 272 1232 306
rect 870 238 892 272
rect 926 238 1232 272
rect 870 234 1232 238
rect 880 232 938 234
rect 842 188 888 200
rect 842 162 848 188
rect 628 114 848 162
rect 842 82 848 114
rect 882 82 888 188
rect 842 70 888 82
rect 930 188 976 200
rect 930 82 936 188
rect 970 158 976 188
rect 1062 158 1068 160
rect 970 110 1068 158
rect 970 82 976 110
rect 1062 108 1068 110
rect 1120 108 1126 160
rect 930 70 976 82
rect -101 17 314 48
rect 1160 42 1232 234
rect -101 4 29 17
rect -101 -48 -70 4
rect -18 -17 29 4
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 314 17
rect -18 -48 314 -17
rect 880 32 1232 42
rect 880 -2 892 32
rect 926 -2 1232 32
rect 880 -30 1232 -2
<< via1 >>
rect 1068 704 1120 756
rect 626 352 678 404
rect 1068 108 1120 160
rect -70 -48 -18 4
<< metal2 >>
rect 1068 756 1120 762
rect 1120 706 1330 754
rect 1068 698 1120 704
rect 626 404 678 410
rect 1282 402 1330 706
rect 678 354 1330 402
rect 626 346 678 352
rect 1068 160 1120 166
rect 1120 110 1370 158
rect 1068 102 1120 108
rect -70 4 -18 10
rect -70 -54 -18 -48
rect -68 -180 -20 -54
rect 1322 -180 1370 110
rect -68 -228 1370 -180
<< labels >>
flabel metal1 -214 658 -214 658 1 FreeSans 480 0 0 0 in
port 2 n
flabel metal2 1312 536 1312 536 1 FreeSans 480 0 0 0 out
port 4 n
flabel metal1 326 734 326 734 1 FreeSans 480 0 0 0 VDD
port 1 n power bidirectional
flabel metal2 512 -206 512 -206 1 FreeSans 480 0 0 0 VSS
port 3 n ground bidirectional
flabel metal1 392 236 392 236 1 FreeSans 480 0 0 0 out2
port 5 n
flabel locali 72 221 106 255 0 FreeSans 340 0 0 0 inv1_0/A
flabel locali 164 289 198 323 0 FreeSans 340 0 0 0 inv1_0/Y
flabel metal1 29 527 63 561 0 FreeSans 200 0 0 0 inv1_0/VPWR
flabel metal1 29 -17 63 17 0 FreeSans 200 0 0 0 inv1_0/VGND
rlabel comment 0 0 0 0 4 inv1_0/inv_1
<< end >>
