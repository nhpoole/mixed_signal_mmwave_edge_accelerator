magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< metal1 >>
rect -60 300 60 357
rect -60 -357 60 -300
<< rmetal1 >>
rect -60 -300 60 300
<< properties >>
string gencell sky130_fd_pr__res_generic_m1
string parameters w 0.6 l 3 m 1 nx 1 wmin 0.14 lmin 0.14 rho 0.125 val 625.0m dummy 0 dw 0.0 term 0.0 roverlap 0
string library sky130
<< end >>
