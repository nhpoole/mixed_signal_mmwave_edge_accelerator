magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -2895 -1848 2895 1848
<< pwell >>
rect -1635 -526 1635 526
<< mvnmos >>
rect -1551 -500 -1451 500
rect -1393 -500 -1293 500
rect -1235 -500 -1135 500
rect -1077 -500 -977 500
rect -919 -500 -819 500
rect -761 -500 -661 500
rect -603 -500 -503 500
rect -445 -500 -345 500
rect -287 -500 -187 500
rect -129 -500 -29 500
rect 29 -500 129 500
rect 187 -500 287 500
rect 345 -500 445 500
rect 503 -500 603 500
rect 661 -500 761 500
rect 819 -500 919 500
rect 977 -500 1077 500
rect 1135 -500 1235 500
rect 1293 -500 1393 500
rect 1451 -500 1551 500
<< mvndiff >>
rect -1609 459 -1551 500
rect -1609 425 -1597 459
rect -1563 425 -1551 459
rect -1609 391 -1551 425
rect -1609 357 -1597 391
rect -1563 357 -1551 391
rect -1609 323 -1551 357
rect -1609 289 -1597 323
rect -1563 289 -1551 323
rect -1609 255 -1551 289
rect -1609 221 -1597 255
rect -1563 221 -1551 255
rect -1609 187 -1551 221
rect -1609 153 -1597 187
rect -1563 153 -1551 187
rect -1609 119 -1551 153
rect -1609 85 -1597 119
rect -1563 85 -1551 119
rect -1609 51 -1551 85
rect -1609 17 -1597 51
rect -1563 17 -1551 51
rect -1609 -17 -1551 17
rect -1609 -51 -1597 -17
rect -1563 -51 -1551 -17
rect -1609 -85 -1551 -51
rect -1609 -119 -1597 -85
rect -1563 -119 -1551 -85
rect -1609 -153 -1551 -119
rect -1609 -187 -1597 -153
rect -1563 -187 -1551 -153
rect -1609 -221 -1551 -187
rect -1609 -255 -1597 -221
rect -1563 -255 -1551 -221
rect -1609 -289 -1551 -255
rect -1609 -323 -1597 -289
rect -1563 -323 -1551 -289
rect -1609 -357 -1551 -323
rect -1609 -391 -1597 -357
rect -1563 -391 -1551 -357
rect -1609 -425 -1551 -391
rect -1609 -459 -1597 -425
rect -1563 -459 -1551 -425
rect -1609 -500 -1551 -459
rect -1451 459 -1393 500
rect -1451 425 -1439 459
rect -1405 425 -1393 459
rect -1451 391 -1393 425
rect -1451 357 -1439 391
rect -1405 357 -1393 391
rect -1451 323 -1393 357
rect -1451 289 -1439 323
rect -1405 289 -1393 323
rect -1451 255 -1393 289
rect -1451 221 -1439 255
rect -1405 221 -1393 255
rect -1451 187 -1393 221
rect -1451 153 -1439 187
rect -1405 153 -1393 187
rect -1451 119 -1393 153
rect -1451 85 -1439 119
rect -1405 85 -1393 119
rect -1451 51 -1393 85
rect -1451 17 -1439 51
rect -1405 17 -1393 51
rect -1451 -17 -1393 17
rect -1451 -51 -1439 -17
rect -1405 -51 -1393 -17
rect -1451 -85 -1393 -51
rect -1451 -119 -1439 -85
rect -1405 -119 -1393 -85
rect -1451 -153 -1393 -119
rect -1451 -187 -1439 -153
rect -1405 -187 -1393 -153
rect -1451 -221 -1393 -187
rect -1451 -255 -1439 -221
rect -1405 -255 -1393 -221
rect -1451 -289 -1393 -255
rect -1451 -323 -1439 -289
rect -1405 -323 -1393 -289
rect -1451 -357 -1393 -323
rect -1451 -391 -1439 -357
rect -1405 -391 -1393 -357
rect -1451 -425 -1393 -391
rect -1451 -459 -1439 -425
rect -1405 -459 -1393 -425
rect -1451 -500 -1393 -459
rect -1293 459 -1235 500
rect -1293 425 -1281 459
rect -1247 425 -1235 459
rect -1293 391 -1235 425
rect -1293 357 -1281 391
rect -1247 357 -1235 391
rect -1293 323 -1235 357
rect -1293 289 -1281 323
rect -1247 289 -1235 323
rect -1293 255 -1235 289
rect -1293 221 -1281 255
rect -1247 221 -1235 255
rect -1293 187 -1235 221
rect -1293 153 -1281 187
rect -1247 153 -1235 187
rect -1293 119 -1235 153
rect -1293 85 -1281 119
rect -1247 85 -1235 119
rect -1293 51 -1235 85
rect -1293 17 -1281 51
rect -1247 17 -1235 51
rect -1293 -17 -1235 17
rect -1293 -51 -1281 -17
rect -1247 -51 -1235 -17
rect -1293 -85 -1235 -51
rect -1293 -119 -1281 -85
rect -1247 -119 -1235 -85
rect -1293 -153 -1235 -119
rect -1293 -187 -1281 -153
rect -1247 -187 -1235 -153
rect -1293 -221 -1235 -187
rect -1293 -255 -1281 -221
rect -1247 -255 -1235 -221
rect -1293 -289 -1235 -255
rect -1293 -323 -1281 -289
rect -1247 -323 -1235 -289
rect -1293 -357 -1235 -323
rect -1293 -391 -1281 -357
rect -1247 -391 -1235 -357
rect -1293 -425 -1235 -391
rect -1293 -459 -1281 -425
rect -1247 -459 -1235 -425
rect -1293 -500 -1235 -459
rect -1135 459 -1077 500
rect -1135 425 -1123 459
rect -1089 425 -1077 459
rect -1135 391 -1077 425
rect -1135 357 -1123 391
rect -1089 357 -1077 391
rect -1135 323 -1077 357
rect -1135 289 -1123 323
rect -1089 289 -1077 323
rect -1135 255 -1077 289
rect -1135 221 -1123 255
rect -1089 221 -1077 255
rect -1135 187 -1077 221
rect -1135 153 -1123 187
rect -1089 153 -1077 187
rect -1135 119 -1077 153
rect -1135 85 -1123 119
rect -1089 85 -1077 119
rect -1135 51 -1077 85
rect -1135 17 -1123 51
rect -1089 17 -1077 51
rect -1135 -17 -1077 17
rect -1135 -51 -1123 -17
rect -1089 -51 -1077 -17
rect -1135 -85 -1077 -51
rect -1135 -119 -1123 -85
rect -1089 -119 -1077 -85
rect -1135 -153 -1077 -119
rect -1135 -187 -1123 -153
rect -1089 -187 -1077 -153
rect -1135 -221 -1077 -187
rect -1135 -255 -1123 -221
rect -1089 -255 -1077 -221
rect -1135 -289 -1077 -255
rect -1135 -323 -1123 -289
rect -1089 -323 -1077 -289
rect -1135 -357 -1077 -323
rect -1135 -391 -1123 -357
rect -1089 -391 -1077 -357
rect -1135 -425 -1077 -391
rect -1135 -459 -1123 -425
rect -1089 -459 -1077 -425
rect -1135 -500 -1077 -459
rect -977 459 -919 500
rect -977 425 -965 459
rect -931 425 -919 459
rect -977 391 -919 425
rect -977 357 -965 391
rect -931 357 -919 391
rect -977 323 -919 357
rect -977 289 -965 323
rect -931 289 -919 323
rect -977 255 -919 289
rect -977 221 -965 255
rect -931 221 -919 255
rect -977 187 -919 221
rect -977 153 -965 187
rect -931 153 -919 187
rect -977 119 -919 153
rect -977 85 -965 119
rect -931 85 -919 119
rect -977 51 -919 85
rect -977 17 -965 51
rect -931 17 -919 51
rect -977 -17 -919 17
rect -977 -51 -965 -17
rect -931 -51 -919 -17
rect -977 -85 -919 -51
rect -977 -119 -965 -85
rect -931 -119 -919 -85
rect -977 -153 -919 -119
rect -977 -187 -965 -153
rect -931 -187 -919 -153
rect -977 -221 -919 -187
rect -977 -255 -965 -221
rect -931 -255 -919 -221
rect -977 -289 -919 -255
rect -977 -323 -965 -289
rect -931 -323 -919 -289
rect -977 -357 -919 -323
rect -977 -391 -965 -357
rect -931 -391 -919 -357
rect -977 -425 -919 -391
rect -977 -459 -965 -425
rect -931 -459 -919 -425
rect -977 -500 -919 -459
rect -819 459 -761 500
rect -819 425 -807 459
rect -773 425 -761 459
rect -819 391 -761 425
rect -819 357 -807 391
rect -773 357 -761 391
rect -819 323 -761 357
rect -819 289 -807 323
rect -773 289 -761 323
rect -819 255 -761 289
rect -819 221 -807 255
rect -773 221 -761 255
rect -819 187 -761 221
rect -819 153 -807 187
rect -773 153 -761 187
rect -819 119 -761 153
rect -819 85 -807 119
rect -773 85 -761 119
rect -819 51 -761 85
rect -819 17 -807 51
rect -773 17 -761 51
rect -819 -17 -761 17
rect -819 -51 -807 -17
rect -773 -51 -761 -17
rect -819 -85 -761 -51
rect -819 -119 -807 -85
rect -773 -119 -761 -85
rect -819 -153 -761 -119
rect -819 -187 -807 -153
rect -773 -187 -761 -153
rect -819 -221 -761 -187
rect -819 -255 -807 -221
rect -773 -255 -761 -221
rect -819 -289 -761 -255
rect -819 -323 -807 -289
rect -773 -323 -761 -289
rect -819 -357 -761 -323
rect -819 -391 -807 -357
rect -773 -391 -761 -357
rect -819 -425 -761 -391
rect -819 -459 -807 -425
rect -773 -459 -761 -425
rect -819 -500 -761 -459
rect -661 459 -603 500
rect -661 425 -649 459
rect -615 425 -603 459
rect -661 391 -603 425
rect -661 357 -649 391
rect -615 357 -603 391
rect -661 323 -603 357
rect -661 289 -649 323
rect -615 289 -603 323
rect -661 255 -603 289
rect -661 221 -649 255
rect -615 221 -603 255
rect -661 187 -603 221
rect -661 153 -649 187
rect -615 153 -603 187
rect -661 119 -603 153
rect -661 85 -649 119
rect -615 85 -603 119
rect -661 51 -603 85
rect -661 17 -649 51
rect -615 17 -603 51
rect -661 -17 -603 17
rect -661 -51 -649 -17
rect -615 -51 -603 -17
rect -661 -85 -603 -51
rect -661 -119 -649 -85
rect -615 -119 -603 -85
rect -661 -153 -603 -119
rect -661 -187 -649 -153
rect -615 -187 -603 -153
rect -661 -221 -603 -187
rect -661 -255 -649 -221
rect -615 -255 -603 -221
rect -661 -289 -603 -255
rect -661 -323 -649 -289
rect -615 -323 -603 -289
rect -661 -357 -603 -323
rect -661 -391 -649 -357
rect -615 -391 -603 -357
rect -661 -425 -603 -391
rect -661 -459 -649 -425
rect -615 -459 -603 -425
rect -661 -500 -603 -459
rect -503 459 -445 500
rect -503 425 -491 459
rect -457 425 -445 459
rect -503 391 -445 425
rect -503 357 -491 391
rect -457 357 -445 391
rect -503 323 -445 357
rect -503 289 -491 323
rect -457 289 -445 323
rect -503 255 -445 289
rect -503 221 -491 255
rect -457 221 -445 255
rect -503 187 -445 221
rect -503 153 -491 187
rect -457 153 -445 187
rect -503 119 -445 153
rect -503 85 -491 119
rect -457 85 -445 119
rect -503 51 -445 85
rect -503 17 -491 51
rect -457 17 -445 51
rect -503 -17 -445 17
rect -503 -51 -491 -17
rect -457 -51 -445 -17
rect -503 -85 -445 -51
rect -503 -119 -491 -85
rect -457 -119 -445 -85
rect -503 -153 -445 -119
rect -503 -187 -491 -153
rect -457 -187 -445 -153
rect -503 -221 -445 -187
rect -503 -255 -491 -221
rect -457 -255 -445 -221
rect -503 -289 -445 -255
rect -503 -323 -491 -289
rect -457 -323 -445 -289
rect -503 -357 -445 -323
rect -503 -391 -491 -357
rect -457 -391 -445 -357
rect -503 -425 -445 -391
rect -503 -459 -491 -425
rect -457 -459 -445 -425
rect -503 -500 -445 -459
rect -345 459 -287 500
rect -345 425 -333 459
rect -299 425 -287 459
rect -345 391 -287 425
rect -345 357 -333 391
rect -299 357 -287 391
rect -345 323 -287 357
rect -345 289 -333 323
rect -299 289 -287 323
rect -345 255 -287 289
rect -345 221 -333 255
rect -299 221 -287 255
rect -345 187 -287 221
rect -345 153 -333 187
rect -299 153 -287 187
rect -345 119 -287 153
rect -345 85 -333 119
rect -299 85 -287 119
rect -345 51 -287 85
rect -345 17 -333 51
rect -299 17 -287 51
rect -345 -17 -287 17
rect -345 -51 -333 -17
rect -299 -51 -287 -17
rect -345 -85 -287 -51
rect -345 -119 -333 -85
rect -299 -119 -287 -85
rect -345 -153 -287 -119
rect -345 -187 -333 -153
rect -299 -187 -287 -153
rect -345 -221 -287 -187
rect -345 -255 -333 -221
rect -299 -255 -287 -221
rect -345 -289 -287 -255
rect -345 -323 -333 -289
rect -299 -323 -287 -289
rect -345 -357 -287 -323
rect -345 -391 -333 -357
rect -299 -391 -287 -357
rect -345 -425 -287 -391
rect -345 -459 -333 -425
rect -299 -459 -287 -425
rect -345 -500 -287 -459
rect -187 459 -129 500
rect -187 425 -175 459
rect -141 425 -129 459
rect -187 391 -129 425
rect -187 357 -175 391
rect -141 357 -129 391
rect -187 323 -129 357
rect -187 289 -175 323
rect -141 289 -129 323
rect -187 255 -129 289
rect -187 221 -175 255
rect -141 221 -129 255
rect -187 187 -129 221
rect -187 153 -175 187
rect -141 153 -129 187
rect -187 119 -129 153
rect -187 85 -175 119
rect -141 85 -129 119
rect -187 51 -129 85
rect -187 17 -175 51
rect -141 17 -129 51
rect -187 -17 -129 17
rect -187 -51 -175 -17
rect -141 -51 -129 -17
rect -187 -85 -129 -51
rect -187 -119 -175 -85
rect -141 -119 -129 -85
rect -187 -153 -129 -119
rect -187 -187 -175 -153
rect -141 -187 -129 -153
rect -187 -221 -129 -187
rect -187 -255 -175 -221
rect -141 -255 -129 -221
rect -187 -289 -129 -255
rect -187 -323 -175 -289
rect -141 -323 -129 -289
rect -187 -357 -129 -323
rect -187 -391 -175 -357
rect -141 -391 -129 -357
rect -187 -425 -129 -391
rect -187 -459 -175 -425
rect -141 -459 -129 -425
rect -187 -500 -129 -459
rect -29 459 29 500
rect -29 425 -17 459
rect 17 425 29 459
rect -29 391 29 425
rect -29 357 -17 391
rect 17 357 29 391
rect -29 323 29 357
rect -29 289 -17 323
rect 17 289 29 323
rect -29 255 29 289
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -289 29 -255
rect -29 -323 -17 -289
rect 17 -323 29 -289
rect -29 -357 29 -323
rect -29 -391 -17 -357
rect 17 -391 29 -357
rect -29 -425 29 -391
rect -29 -459 -17 -425
rect 17 -459 29 -425
rect -29 -500 29 -459
rect 129 459 187 500
rect 129 425 141 459
rect 175 425 187 459
rect 129 391 187 425
rect 129 357 141 391
rect 175 357 187 391
rect 129 323 187 357
rect 129 289 141 323
rect 175 289 187 323
rect 129 255 187 289
rect 129 221 141 255
rect 175 221 187 255
rect 129 187 187 221
rect 129 153 141 187
rect 175 153 187 187
rect 129 119 187 153
rect 129 85 141 119
rect 175 85 187 119
rect 129 51 187 85
rect 129 17 141 51
rect 175 17 187 51
rect 129 -17 187 17
rect 129 -51 141 -17
rect 175 -51 187 -17
rect 129 -85 187 -51
rect 129 -119 141 -85
rect 175 -119 187 -85
rect 129 -153 187 -119
rect 129 -187 141 -153
rect 175 -187 187 -153
rect 129 -221 187 -187
rect 129 -255 141 -221
rect 175 -255 187 -221
rect 129 -289 187 -255
rect 129 -323 141 -289
rect 175 -323 187 -289
rect 129 -357 187 -323
rect 129 -391 141 -357
rect 175 -391 187 -357
rect 129 -425 187 -391
rect 129 -459 141 -425
rect 175 -459 187 -425
rect 129 -500 187 -459
rect 287 459 345 500
rect 287 425 299 459
rect 333 425 345 459
rect 287 391 345 425
rect 287 357 299 391
rect 333 357 345 391
rect 287 323 345 357
rect 287 289 299 323
rect 333 289 345 323
rect 287 255 345 289
rect 287 221 299 255
rect 333 221 345 255
rect 287 187 345 221
rect 287 153 299 187
rect 333 153 345 187
rect 287 119 345 153
rect 287 85 299 119
rect 333 85 345 119
rect 287 51 345 85
rect 287 17 299 51
rect 333 17 345 51
rect 287 -17 345 17
rect 287 -51 299 -17
rect 333 -51 345 -17
rect 287 -85 345 -51
rect 287 -119 299 -85
rect 333 -119 345 -85
rect 287 -153 345 -119
rect 287 -187 299 -153
rect 333 -187 345 -153
rect 287 -221 345 -187
rect 287 -255 299 -221
rect 333 -255 345 -221
rect 287 -289 345 -255
rect 287 -323 299 -289
rect 333 -323 345 -289
rect 287 -357 345 -323
rect 287 -391 299 -357
rect 333 -391 345 -357
rect 287 -425 345 -391
rect 287 -459 299 -425
rect 333 -459 345 -425
rect 287 -500 345 -459
rect 445 459 503 500
rect 445 425 457 459
rect 491 425 503 459
rect 445 391 503 425
rect 445 357 457 391
rect 491 357 503 391
rect 445 323 503 357
rect 445 289 457 323
rect 491 289 503 323
rect 445 255 503 289
rect 445 221 457 255
rect 491 221 503 255
rect 445 187 503 221
rect 445 153 457 187
rect 491 153 503 187
rect 445 119 503 153
rect 445 85 457 119
rect 491 85 503 119
rect 445 51 503 85
rect 445 17 457 51
rect 491 17 503 51
rect 445 -17 503 17
rect 445 -51 457 -17
rect 491 -51 503 -17
rect 445 -85 503 -51
rect 445 -119 457 -85
rect 491 -119 503 -85
rect 445 -153 503 -119
rect 445 -187 457 -153
rect 491 -187 503 -153
rect 445 -221 503 -187
rect 445 -255 457 -221
rect 491 -255 503 -221
rect 445 -289 503 -255
rect 445 -323 457 -289
rect 491 -323 503 -289
rect 445 -357 503 -323
rect 445 -391 457 -357
rect 491 -391 503 -357
rect 445 -425 503 -391
rect 445 -459 457 -425
rect 491 -459 503 -425
rect 445 -500 503 -459
rect 603 459 661 500
rect 603 425 615 459
rect 649 425 661 459
rect 603 391 661 425
rect 603 357 615 391
rect 649 357 661 391
rect 603 323 661 357
rect 603 289 615 323
rect 649 289 661 323
rect 603 255 661 289
rect 603 221 615 255
rect 649 221 661 255
rect 603 187 661 221
rect 603 153 615 187
rect 649 153 661 187
rect 603 119 661 153
rect 603 85 615 119
rect 649 85 661 119
rect 603 51 661 85
rect 603 17 615 51
rect 649 17 661 51
rect 603 -17 661 17
rect 603 -51 615 -17
rect 649 -51 661 -17
rect 603 -85 661 -51
rect 603 -119 615 -85
rect 649 -119 661 -85
rect 603 -153 661 -119
rect 603 -187 615 -153
rect 649 -187 661 -153
rect 603 -221 661 -187
rect 603 -255 615 -221
rect 649 -255 661 -221
rect 603 -289 661 -255
rect 603 -323 615 -289
rect 649 -323 661 -289
rect 603 -357 661 -323
rect 603 -391 615 -357
rect 649 -391 661 -357
rect 603 -425 661 -391
rect 603 -459 615 -425
rect 649 -459 661 -425
rect 603 -500 661 -459
rect 761 459 819 500
rect 761 425 773 459
rect 807 425 819 459
rect 761 391 819 425
rect 761 357 773 391
rect 807 357 819 391
rect 761 323 819 357
rect 761 289 773 323
rect 807 289 819 323
rect 761 255 819 289
rect 761 221 773 255
rect 807 221 819 255
rect 761 187 819 221
rect 761 153 773 187
rect 807 153 819 187
rect 761 119 819 153
rect 761 85 773 119
rect 807 85 819 119
rect 761 51 819 85
rect 761 17 773 51
rect 807 17 819 51
rect 761 -17 819 17
rect 761 -51 773 -17
rect 807 -51 819 -17
rect 761 -85 819 -51
rect 761 -119 773 -85
rect 807 -119 819 -85
rect 761 -153 819 -119
rect 761 -187 773 -153
rect 807 -187 819 -153
rect 761 -221 819 -187
rect 761 -255 773 -221
rect 807 -255 819 -221
rect 761 -289 819 -255
rect 761 -323 773 -289
rect 807 -323 819 -289
rect 761 -357 819 -323
rect 761 -391 773 -357
rect 807 -391 819 -357
rect 761 -425 819 -391
rect 761 -459 773 -425
rect 807 -459 819 -425
rect 761 -500 819 -459
rect 919 459 977 500
rect 919 425 931 459
rect 965 425 977 459
rect 919 391 977 425
rect 919 357 931 391
rect 965 357 977 391
rect 919 323 977 357
rect 919 289 931 323
rect 965 289 977 323
rect 919 255 977 289
rect 919 221 931 255
rect 965 221 977 255
rect 919 187 977 221
rect 919 153 931 187
rect 965 153 977 187
rect 919 119 977 153
rect 919 85 931 119
rect 965 85 977 119
rect 919 51 977 85
rect 919 17 931 51
rect 965 17 977 51
rect 919 -17 977 17
rect 919 -51 931 -17
rect 965 -51 977 -17
rect 919 -85 977 -51
rect 919 -119 931 -85
rect 965 -119 977 -85
rect 919 -153 977 -119
rect 919 -187 931 -153
rect 965 -187 977 -153
rect 919 -221 977 -187
rect 919 -255 931 -221
rect 965 -255 977 -221
rect 919 -289 977 -255
rect 919 -323 931 -289
rect 965 -323 977 -289
rect 919 -357 977 -323
rect 919 -391 931 -357
rect 965 -391 977 -357
rect 919 -425 977 -391
rect 919 -459 931 -425
rect 965 -459 977 -425
rect 919 -500 977 -459
rect 1077 459 1135 500
rect 1077 425 1089 459
rect 1123 425 1135 459
rect 1077 391 1135 425
rect 1077 357 1089 391
rect 1123 357 1135 391
rect 1077 323 1135 357
rect 1077 289 1089 323
rect 1123 289 1135 323
rect 1077 255 1135 289
rect 1077 221 1089 255
rect 1123 221 1135 255
rect 1077 187 1135 221
rect 1077 153 1089 187
rect 1123 153 1135 187
rect 1077 119 1135 153
rect 1077 85 1089 119
rect 1123 85 1135 119
rect 1077 51 1135 85
rect 1077 17 1089 51
rect 1123 17 1135 51
rect 1077 -17 1135 17
rect 1077 -51 1089 -17
rect 1123 -51 1135 -17
rect 1077 -85 1135 -51
rect 1077 -119 1089 -85
rect 1123 -119 1135 -85
rect 1077 -153 1135 -119
rect 1077 -187 1089 -153
rect 1123 -187 1135 -153
rect 1077 -221 1135 -187
rect 1077 -255 1089 -221
rect 1123 -255 1135 -221
rect 1077 -289 1135 -255
rect 1077 -323 1089 -289
rect 1123 -323 1135 -289
rect 1077 -357 1135 -323
rect 1077 -391 1089 -357
rect 1123 -391 1135 -357
rect 1077 -425 1135 -391
rect 1077 -459 1089 -425
rect 1123 -459 1135 -425
rect 1077 -500 1135 -459
rect 1235 459 1293 500
rect 1235 425 1247 459
rect 1281 425 1293 459
rect 1235 391 1293 425
rect 1235 357 1247 391
rect 1281 357 1293 391
rect 1235 323 1293 357
rect 1235 289 1247 323
rect 1281 289 1293 323
rect 1235 255 1293 289
rect 1235 221 1247 255
rect 1281 221 1293 255
rect 1235 187 1293 221
rect 1235 153 1247 187
rect 1281 153 1293 187
rect 1235 119 1293 153
rect 1235 85 1247 119
rect 1281 85 1293 119
rect 1235 51 1293 85
rect 1235 17 1247 51
rect 1281 17 1293 51
rect 1235 -17 1293 17
rect 1235 -51 1247 -17
rect 1281 -51 1293 -17
rect 1235 -85 1293 -51
rect 1235 -119 1247 -85
rect 1281 -119 1293 -85
rect 1235 -153 1293 -119
rect 1235 -187 1247 -153
rect 1281 -187 1293 -153
rect 1235 -221 1293 -187
rect 1235 -255 1247 -221
rect 1281 -255 1293 -221
rect 1235 -289 1293 -255
rect 1235 -323 1247 -289
rect 1281 -323 1293 -289
rect 1235 -357 1293 -323
rect 1235 -391 1247 -357
rect 1281 -391 1293 -357
rect 1235 -425 1293 -391
rect 1235 -459 1247 -425
rect 1281 -459 1293 -425
rect 1235 -500 1293 -459
rect 1393 459 1451 500
rect 1393 425 1405 459
rect 1439 425 1451 459
rect 1393 391 1451 425
rect 1393 357 1405 391
rect 1439 357 1451 391
rect 1393 323 1451 357
rect 1393 289 1405 323
rect 1439 289 1451 323
rect 1393 255 1451 289
rect 1393 221 1405 255
rect 1439 221 1451 255
rect 1393 187 1451 221
rect 1393 153 1405 187
rect 1439 153 1451 187
rect 1393 119 1451 153
rect 1393 85 1405 119
rect 1439 85 1451 119
rect 1393 51 1451 85
rect 1393 17 1405 51
rect 1439 17 1451 51
rect 1393 -17 1451 17
rect 1393 -51 1405 -17
rect 1439 -51 1451 -17
rect 1393 -85 1451 -51
rect 1393 -119 1405 -85
rect 1439 -119 1451 -85
rect 1393 -153 1451 -119
rect 1393 -187 1405 -153
rect 1439 -187 1451 -153
rect 1393 -221 1451 -187
rect 1393 -255 1405 -221
rect 1439 -255 1451 -221
rect 1393 -289 1451 -255
rect 1393 -323 1405 -289
rect 1439 -323 1451 -289
rect 1393 -357 1451 -323
rect 1393 -391 1405 -357
rect 1439 -391 1451 -357
rect 1393 -425 1451 -391
rect 1393 -459 1405 -425
rect 1439 -459 1451 -425
rect 1393 -500 1451 -459
rect 1551 459 1609 500
rect 1551 425 1563 459
rect 1597 425 1609 459
rect 1551 391 1609 425
rect 1551 357 1563 391
rect 1597 357 1609 391
rect 1551 323 1609 357
rect 1551 289 1563 323
rect 1597 289 1609 323
rect 1551 255 1609 289
rect 1551 221 1563 255
rect 1597 221 1609 255
rect 1551 187 1609 221
rect 1551 153 1563 187
rect 1597 153 1609 187
rect 1551 119 1609 153
rect 1551 85 1563 119
rect 1597 85 1609 119
rect 1551 51 1609 85
rect 1551 17 1563 51
rect 1597 17 1609 51
rect 1551 -17 1609 17
rect 1551 -51 1563 -17
rect 1597 -51 1609 -17
rect 1551 -85 1609 -51
rect 1551 -119 1563 -85
rect 1597 -119 1609 -85
rect 1551 -153 1609 -119
rect 1551 -187 1563 -153
rect 1597 -187 1609 -153
rect 1551 -221 1609 -187
rect 1551 -255 1563 -221
rect 1597 -255 1609 -221
rect 1551 -289 1609 -255
rect 1551 -323 1563 -289
rect 1597 -323 1609 -289
rect 1551 -357 1609 -323
rect 1551 -391 1563 -357
rect 1597 -391 1609 -357
rect 1551 -425 1609 -391
rect 1551 -459 1563 -425
rect 1597 -459 1609 -425
rect 1551 -500 1609 -459
<< mvndiffc >>
rect -1597 425 -1563 459
rect -1597 357 -1563 391
rect -1597 289 -1563 323
rect -1597 221 -1563 255
rect -1597 153 -1563 187
rect -1597 85 -1563 119
rect -1597 17 -1563 51
rect -1597 -51 -1563 -17
rect -1597 -119 -1563 -85
rect -1597 -187 -1563 -153
rect -1597 -255 -1563 -221
rect -1597 -323 -1563 -289
rect -1597 -391 -1563 -357
rect -1597 -459 -1563 -425
rect -1439 425 -1405 459
rect -1439 357 -1405 391
rect -1439 289 -1405 323
rect -1439 221 -1405 255
rect -1439 153 -1405 187
rect -1439 85 -1405 119
rect -1439 17 -1405 51
rect -1439 -51 -1405 -17
rect -1439 -119 -1405 -85
rect -1439 -187 -1405 -153
rect -1439 -255 -1405 -221
rect -1439 -323 -1405 -289
rect -1439 -391 -1405 -357
rect -1439 -459 -1405 -425
rect -1281 425 -1247 459
rect -1281 357 -1247 391
rect -1281 289 -1247 323
rect -1281 221 -1247 255
rect -1281 153 -1247 187
rect -1281 85 -1247 119
rect -1281 17 -1247 51
rect -1281 -51 -1247 -17
rect -1281 -119 -1247 -85
rect -1281 -187 -1247 -153
rect -1281 -255 -1247 -221
rect -1281 -323 -1247 -289
rect -1281 -391 -1247 -357
rect -1281 -459 -1247 -425
rect -1123 425 -1089 459
rect -1123 357 -1089 391
rect -1123 289 -1089 323
rect -1123 221 -1089 255
rect -1123 153 -1089 187
rect -1123 85 -1089 119
rect -1123 17 -1089 51
rect -1123 -51 -1089 -17
rect -1123 -119 -1089 -85
rect -1123 -187 -1089 -153
rect -1123 -255 -1089 -221
rect -1123 -323 -1089 -289
rect -1123 -391 -1089 -357
rect -1123 -459 -1089 -425
rect -965 425 -931 459
rect -965 357 -931 391
rect -965 289 -931 323
rect -965 221 -931 255
rect -965 153 -931 187
rect -965 85 -931 119
rect -965 17 -931 51
rect -965 -51 -931 -17
rect -965 -119 -931 -85
rect -965 -187 -931 -153
rect -965 -255 -931 -221
rect -965 -323 -931 -289
rect -965 -391 -931 -357
rect -965 -459 -931 -425
rect -807 425 -773 459
rect -807 357 -773 391
rect -807 289 -773 323
rect -807 221 -773 255
rect -807 153 -773 187
rect -807 85 -773 119
rect -807 17 -773 51
rect -807 -51 -773 -17
rect -807 -119 -773 -85
rect -807 -187 -773 -153
rect -807 -255 -773 -221
rect -807 -323 -773 -289
rect -807 -391 -773 -357
rect -807 -459 -773 -425
rect -649 425 -615 459
rect -649 357 -615 391
rect -649 289 -615 323
rect -649 221 -615 255
rect -649 153 -615 187
rect -649 85 -615 119
rect -649 17 -615 51
rect -649 -51 -615 -17
rect -649 -119 -615 -85
rect -649 -187 -615 -153
rect -649 -255 -615 -221
rect -649 -323 -615 -289
rect -649 -391 -615 -357
rect -649 -459 -615 -425
rect -491 425 -457 459
rect -491 357 -457 391
rect -491 289 -457 323
rect -491 221 -457 255
rect -491 153 -457 187
rect -491 85 -457 119
rect -491 17 -457 51
rect -491 -51 -457 -17
rect -491 -119 -457 -85
rect -491 -187 -457 -153
rect -491 -255 -457 -221
rect -491 -323 -457 -289
rect -491 -391 -457 -357
rect -491 -459 -457 -425
rect -333 425 -299 459
rect -333 357 -299 391
rect -333 289 -299 323
rect -333 221 -299 255
rect -333 153 -299 187
rect -333 85 -299 119
rect -333 17 -299 51
rect -333 -51 -299 -17
rect -333 -119 -299 -85
rect -333 -187 -299 -153
rect -333 -255 -299 -221
rect -333 -323 -299 -289
rect -333 -391 -299 -357
rect -333 -459 -299 -425
rect -175 425 -141 459
rect -175 357 -141 391
rect -175 289 -141 323
rect -175 221 -141 255
rect -175 153 -141 187
rect -175 85 -141 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -175 -119 -141 -85
rect -175 -187 -141 -153
rect -175 -255 -141 -221
rect -175 -323 -141 -289
rect -175 -391 -141 -357
rect -175 -459 -141 -425
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect 141 425 175 459
rect 141 357 175 391
rect 141 289 175 323
rect 141 221 175 255
rect 141 153 175 187
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect 141 -187 175 -153
rect 141 -255 175 -221
rect 141 -323 175 -289
rect 141 -391 175 -357
rect 141 -459 175 -425
rect 299 425 333 459
rect 299 357 333 391
rect 299 289 333 323
rect 299 221 333 255
rect 299 153 333 187
rect 299 85 333 119
rect 299 17 333 51
rect 299 -51 333 -17
rect 299 -119 333 -85
rect 299 -187 333 -153
rect 299 -255 333 -221
rect 299 -323 333 -289
rect 299 -391 333 -357
rect 299 -459 333 -425
rect 457 425 491 459
rect 457 357 491 391
rect 457 289 491 323
rect 457 221 491 255
rect 457 153 491 187
rect 457 85 491 119
rect 457 17 491 51
rect 457 -51 491 -17
rect 457 -119 491 -85
rect 457 -187 491 -153
rect 457 -255 491 -221
rect 457 -323 491 -289
rect 457 -391 491 -357
rect 457 -459 491 -425
rect 615 425 649 459
rect 615 357 649 391
rect 615 289 649 323
rect 615 221 649 255
rect 615 153 649 187
rect 615 85 649 119
rect 615 17 649 51
rect 615 -51 649 -17
rect 615 -119 649 -85
rect 615 -187 649 -153
rect 615 -255 649 -221
rect 615 -323 649 -289
rect 615 -391 649 -357
rect 615 -459 649 -425
rect 773 425 807 459
rect 773 357 807 391
rect 773 289 807 323
rect 773 221 807 255
rect 773 153 807 187
rect 773 85 807 119
rect 773 17 807 51
rect 773 -51 807 -17
rect 773 -119 807 -85
rect 773 -187 807 -153
rect 773 -255 807 -221
rect 773 -323 807 -289
rect 773 -391 807 -357
rect 773 -459 807 -425
rect 931 425 965 459
rect 931 357 965 391
rect 931 289 965 323
rect 931 221 965 255
rect 931 153 965 187
rect 931 85 965 119
rect 931 17 965 51
rect 931 -51 965 -17
rect 931 -119 965 -85
rect 931 -187 965 -153
rect 931 -255 965 -221
rect 931 -323 965 -289
rect 931 -391 965 -357
rect 931 -459 965 -425
rect 1089 425 1123 459
rect 1089 357 1123 391
rect 1089 289 1123 323
rect 1089 221 1123 255
rect 1089 153 1123 187
rect 1089 85 1123 119
rect 1089 17 1123 51
rect 1089 -51 1123 -17
rect 1089 -119 1123 -85
rect 1089 -187 1123 -153
rect 1089 -255 1123 -221
rect 1089 -323 1123 -289
rect 1089 -391 1123 -357
rect 1089 -459 1123 -425
rect 1247 425 1281 459
rect 1247 357 1281 391
rect 1247 289 1281 323
rect 1247 221 1281 255
rect 1247 153 1281 187
rect 1247 85 1281 119
rect 1247 17 1281 51
rect 1247 -51 1281 -17
rect 1247 -119 1281 -85
rect 1247 -187 1281 -153
rect 1247 -255 1281 -221
rect 1247 -323 1281 -289
rect 1247 -391 1281 -357
rect 1247 -459 1281 -425
rect 1405 425 1439 459
rect 1405 357 1439 391
rect 1405 289 1439 323
rect 1405 221 1439 255
rect 1405 153 1439 187
rect 1405 85 1439 119
rect 1405 17 1439 51
rect 1405 -51 1439 -17
rect 1405 -119 1439 -85
rect 1405 -187 1439 -153
rect 1405 -255 1439 -221
rect 1405 -323 1439 -289
rect 1405 -391 1439 -357
rect 1405 -459 1439 -425
rect 1563 425 1597 459
rect 1563 357 1597 391
rect 1563 289 1597 323
rect 1563 221 1597 255
rect 1563 153 1597 187
rect 1563 85 1597 119
rect 1563 17 1597 51
rect 1563 -51 1597 -17
rect 1563 -119 1597 -85
rect 1563 -187 1597 -153
rect 1563 -255 1597 -221
rect 1563 -323 1597 -289
rect 1563 -391 1597 -357
rect 1563 -459 1597 -425
<< poly >>
rect -1537 572 -1465 588
rect -1537 555 -1518 572
rect -1551 538 -1518 555
rect -1484 555 -1465 572
rect -1379 572 -1307 588
rect -1379 555 -1360 572
rect -1484 538 -1451 555
rect -1551 500 -1451 538
rect -1393 538 -1360 555
rect -1326 555 -1307 572
rect -1221 572 -1149 588
rect -1221 555 -1202 572
rect -1326 538 -1293 555
rect -1393 500 -1293 538
rect -1235 538 -1202 555
rect -1168 555 -1149 572
rect -1063 572 -991 588
rect -1063 555 -1044 572
rect -1168 538 -1135 555
rect -1235 500 -1135 538
rect -1077 538 -1044 555
rect -1010 555 -991 572
rect -905 572 -833 588
rect -905 555 -886 572
rect -1010 538 -977 555
rect -1077 500 -977 538
rect -919 538 -886 555
rect -852 555 -833 572
rect -747 572 -675 588
rect -747 555 -728 572
rect -852 538 -819 555
rect -919 500 -819 538
rect -761 538 -728 555
rect -694 555 -675 572
rect -589 572 -517 588
rect -589 555 -570 572
rect -694 538 -661 555
rect -761 500 -661 538
rect -603 538 -570 555
rect -536 555 -517 572
rect -431 572 -359 588
rect -431 555 -412 572
rect -536 538 -503 555
rect -603 500 -503 538
rect -445 538 -412 555
rect -378 555 -359 572
rect -273 572 -201 588
rect -273 555 -254 572
rect -378 538 -345 555
rect -445 500 -345 538
rect -287 538 -254 555
rect -220 555 -201 572
rect -115 572 -43 588
rect -115 555 -96 572
rect -220 538 -187 555
rect -287 500 -187 538
rect -129 538 -96 555
rect -62 555 -43 572
rect 43 572 115 588
rect 43 555 62 572
rect -62 538 -29 555
rect -129 500 -29 538
rect 29 538 62 555
rect 96 555 115 572
rect 201 572 273 588
rect 201 555 220 572
rect 96 538 129 555
rect 29 500 129 538
rect 187 538 220 555
rect 254 555 273 572
rect 359 572 431 588
rect 359 555 378 572
rect 254 538 287 555
rect 187 500 287 538
rect 345 538 378 555
rect 412 555 431 572
rect 517 572 589 588
rect 517 555 536 572
rect 412 538 445 555
rect 345 500 445 538
rect 503 538 536 555
rect 570 555 589 572
rect 675 572 747 588
rect 675 555 694 572
rect 570 538 603 555
rect 503 500 603 538
rect 661 538 694 555
rect 728 555 747 572
rect 833 572 905 588
rect 833 555 852 572
rect 728 538 761 555
rect 661 500 761 538
rect 819 538 852 555
rect 886 555 905 572
rect 991 572 1063 588
rect 991 555 1010 572
rect 886 538 919 555
rect 819 500 919 538
rect 977 538 1010 555
rect 1044 555 1063 572
rect 1149 572 1221 588
rect 1149 555 1168 572
rect 1044 538 1077 555
rect 977 500 1077 538
rect 1135 538 1168 555
rect 1202 555 1221 572
rect 1307 572 1379 588
rect 1307 555 1326 572
rect 1202 538 1235 555
rect 1135 500 1235 538
rect 1293 538 1326 555
rect 1360 555 1379 572
rect 1465 572 1537 588
rect 1465 555 1484 572
rect 1360 538 1393 555
rect 1293 500 1393 538
rect 1451 538 1484 555
rect 1518 555 1537 572
rect 1518 538 1551 555
rect 1451 500 1551 538
rect -1551 -538 -1451 -500
rect -1551 -555 -1518 -538
rect -1537 -572 -1518 -555
rect -1484 -555 -1451 -538
rect -1393 -538 -1293 -500
rect -1393 -555 -1360 -538
rect -1484 -572 -1465 -555
rect -1537 -588 -1465 -572
rect -1379 -572 -1360 -555
rect -1326 -555 -1293 -538
rect -1235 -538 -1135 -500
rect -1235 -555 -1202 -538
rect -1326 -572 -1307 -555
rect -1379 -588 -1307 -572
rect -1221 -572 -1202 -555
rect -1168 -555 -1135 -538
rect -1077 -538 -977 -500
rect -1077 -555 -1044 -538
rect -1168 -572 -1149 -555
rect -1221 -588 -1149 -572
rect -1063 -572 -1044 -555
rect -1010 -555 -977 -538
rect -919 -538 -819 -500
rect -919 -555 -886 -538
rect -1010 -572 -991 -555
rect -1063 -588 -991 -572
rect -905 -572 -886 -555
rect -852 -555 -819 -538
rect -761 -538 -661 -500
rect -761 -555 -728 -538
rect -852 -572 -833 -555
rect -905 -588 -833 -572
rect -747 -572 -728 -555
rect -694 -555 -661 -538
rect -603 -538 -503 -500
rect -603 -555 -570 -538
rect -694 -572 -675 -555
rect -747 -588 -675 -572
rect -589 -572 -570 -555
rect -536 -555 -503 -538
rect -445 -538 -345 -500
rect -445 -555 -412 -538
rect -536 -572 -517 -555
rect -589 -588 -517 -572
rect -431 -572 -412 -555
rect -378 -555 -345 -538
rect -287 -538 -187 -500
rect -287 -555 -254 -538
rect -378 -572 -359 -555
rect -431 -588 -359 -572
rect -273 -572 -254 -555
rect -220 -555 -187 -538
rect -129 -538 -29 -500
rect -129 -555 -96 -538
rect -220 -572 -201 -555
rect -273 -588 -201 -572
rect -115 -572 -96 -555
rect -62 -555 -29 -538
rect 29 -538 129 -500
rect 29 -555 62 -538
rect -62 -572 -43 -555
rect -115 -588 -43 -572
rect 43 -572 62 -555
rect 96 -555 129 -538
rect 187 -538 287 -500
rect 187 -555 220 -538
rect 96 -572 115 -555
rect 43 -588 115 -572
rect 201 -572 220 -555
rect 254 -555 287 -538
rect 345 -538 445 -500
rect 345 -555 378 -538
rect 254 -572 273 -555
rect 201 -588 273 -572
rect 359 -572 378 -555
rect 412 -555 445 -538
rect 503 -538 603 -500
rect 503 -555 536 -538
rect 412 -572 431 -555
rect 359 -588 431 -572
rect 517 -572 536 -555
rect 570 -555 603 -538
rect 661 -538 761 -500
rect 661 -555 694 -538
rect 570 -572 589 -555
rect 517 -588 589 -572
rect 675 -572 694 -555
rect 728 -555 761 -538
rect 819 -538 919 -500
rect 819 -555 852 -538
rect 728 -572 747 -555
rect 675 -588 747 -572
rect 833 -572 852 -555
rect 886 -555 919 -538
rect 977 -538 1077 -500
rect 977 -555 1010 -538
rect 886 -572 905 -555
rect 833 -588 905 -572
rect 991 -572 1010 -555
rect 1044 -555 1077 -538
rect 1135 -538 1235 -500
rect 1135 -555 1168 -538
rect 1044 -572 1063 -555
rect 991 -588 1063 -572
rect 1149 -572 1168 -555
rect 1202 -555 1235 -538
rect 1293 -538 1393 -500
rect 1293 -555 1326 -538
rect 1202 -572 1221 -555
rect 1149 -588 1221 -572
rect 1307 -572 1326 -555
rect 1360 -555 1393 -538
rect 1451 -538 1551 -500
rect 1451 -555 1484 -538
rect 1360 -572 1379 -555
rect 1307 -588 1379 -572
rect 1465 -572 1484 -555
rect 1518 -555 1551 -538
rect 1518 -572 1537 -555
rect 1465 -588 1537 -572
<< polycont >>
rect -1518 538 -1484 572
rect -1360 538 -1326 572
rect -1202 538 -1168 572
rect -1044 538 -1010 572
rect -886 538 -852 572
rect -728 538 -694 572
rect -570 538 -536 572
rect -412 538 -378 572
rect -254 538 -220 572
rect -96 538 -62 572
rect 62 538 96 572
rect 220 538 254 572
rect 378 538 412 572
rect 536 538 570 572
rect 694 538 728 572
rect 852 538 886 572
rect 1010 538 1044 572
rect 1168 538 1202 572
rect 1326 538 1360 572
rect 1484 538 1518 572
rect -1518 -572 -1484 -538
rect -1360 -572 -1326 -538
rect -1202 -572 -1168 -538
rect -1044 -572 -1010 -538
rect -886 -572 -852 -538
rect -728 -572 -694 -538
rect -570 -572 -536 -538
rect -412 -572 -378 -538
rect -254 -572 -220 -538
rect -96 -572 -62 -538
rect 62 -572 96 -538
rect 220 -572 254 -538
rect 378 -572 412 -538
rect 536 -572 570 -538
rect 694 -572 728 -538
rect 852 -572 886 -538
rect 1010 -572 1044 -538
rect 1168 -572 1202 -538
rect 1326 -572 1360 -538
rect 1484 -572 1518 -538
<< locali >>
rect -1537 538 -1518 572
rect -1484 538 -1465 572
rect -1379 538 -1360 572
rect -1326 538 -1307 572
rect -1221 538 -1202 572
rect -1168 538 -1149 572
rect -1063 538 -1044 572
rect -1010 538 -991 572
rect -905 538 -886 572
rect -852 538 -833 572
rect -747 538 -728 572
rect -694 538 -675 572
rect -589 538 -570 572
rect -536 538 -517 572
rect -431 538 -412 572
rect -378 538 -359 572
rect -273 538 -254 572
rect -220 538 -201 572
rect -115 538 -96 572
rect -62 538 -43 572
rect 43 538 62 572
rect 96 538 115 572
rect 201 538 220 572
rect 254 538 273 572
rect 359 538 378 572
rect 412 538 431 572
rect 517 538 536 572
rect 570 538 589 572
rect 675 538 694 572
rect 728 538 747 572
rect 833 538 852 572
rect 886 538 905 572
rect 991 538 1010 572
rect 1044 538 1063 572
rect 1149 538 1168 572
rect 1202 538 1221 572
rect 1307 538 1326 572
rect 1360 538 1379 572
rect 1465 538 1484 572
rect 1518 538 1537 572
rect -1597 485 -1563 504
rect -1597 413 -1563 425
rect -1597 341 -1563 357
rect -1597 269 -1563 289
rect -1597 197 -1563 221
rect -1597 125 -1563 153
rect -1597 53 -1563 85
rect -1597 -17 -1563 17
rect -1597 -85 -1563 -53
rect -1597 -153 -1563 -125
rect -1597 -221 -1563 -197
rect -1597 -289 -1563 -269
rect -1597 -357 -1563 -341
rect -1597 -425 -1563 -413
rect -1597 -504 -1563 -485
rect -1439 485 -1405 504
rect -1439 413 -1405 425
rect -1439 341 -1405 357
rect -1439 269 -1405 289
rect -1439 197 -1405 221
rect -1439 125 -1405 153
rect -1439 53 -1405 85
rect -1439 -17 -1405 17
rect -1439 -85 -1405 -53
rect -1439 -153 -1405 -125
rect -1439 -221 -1405 -197
rect -1439 -289 -1405 -269
rect -1439 -357 -1405 -341
rect -1439 -425 -1405 -413
rect -1439 -504 -1405 -485
rect -1281 485 -1247 504
rect -1281 413 -1247 425
rect -1281 341 -1247 357
rect -1281 269 -1247 289
rect -1281 197 -1247 221
rect -1281 125 -1247 153
rect -1281 53 -1247 85
rect -1281 -17 -1247 17
rect -1281 -85 -1247 -53
rect -1281 -153 -1247 -125
rect -1281 -221 -1247 -197
rect -1281 -289 -1247 -269
rect -1281 -357 -1247 -341
rect -1281 -425 -1247 -413
rect -1281 -504 -1247 -485
rect -1123 485 -1089 504
rect -1123 413 -1089 425
rect -1123 341 -1089 357
rect -1123 269 -1089 289
rect -1123 197 -1089 221
rect -1123 125 -1089 153
rect -1123 53 -1089 85
rect -1123 -17 -1089 17
rect -1123 -85 -1089 -53
rect -1123 -153 -1089 -125
rect -1123 -221 -1089 -197
rect -1123 -289 -1089 -269
rect -1123 -357 -1089 -341
rect -1123 -425 -1089 -413
rect -1123 -504 -1089 -485
rect -965 485 -931 504
rect -965 413 -931 425
rect -965 341 -931 357
rect -965 269 -931 289
rect -965 197 -931 221
rect -965 125 -931 153
rect -965 53 -931 85
rect -965 -17 -931 17
rect -965 -85 -931 -53
rect -965 -153 -931 -125
rect -965 -221 -931 -197
rect -965 -289 -931 -269
rect -965 -357 -931 -341
rect -965 -425 -931 -413
rect -965 -504 -931 -485
rect -807 485 -773 504
rect -807 413 -773 425
rect -807 341 -773 357
rect -807 269 -773 289
rect -807 197 -773 221
rect -807 125 -773 153
rect -807 53 -773 85
rect -807 -17 -773 17
rect -807 -85 -773 -53
rect -807 -153 -773 -125
rect -807 -221 -773 -197
rect -807 -289 -773 -269
rect -807 -357 -773 -341
rect -807 -425 -773 -413
rect -807 -504 -773 -485
rect -649 485 -615 504
rect -649 413 -615 425
rect -649 341 -615 357
rect -649 269 -615 289
rect -649 197 -615 221
rect -649 125 -615 153
rect -649 53 -615 85
rect -649 -17 -615 17
rect -649 -85 -615 -53
rect -649 -153 -615 -125
rect -649 -221 -615 -197
rect -649 -289 -615 -269
rect -649 -357 -615 -341
rect -649 -425 -615 -413
rect -649 -504 -615 -485
rect -491 485 -457 504
rect -491 413 -457 425
rect -491 341 -457 357
rect -491 269 -457 289
rect -491 197 -457 221
rect -491 125 -457 153
rect -491 53 -457 85
rect -491 -17 -457 17
rect -491 -85 -457 -53
rect -491 -153 -457 -125
rect -491 -221 -457 -197
rect -491 -289 -457 -269
rect -491 -357 -457 -341
rect -491 -425 -457 -413
rect -491 -504 -457 -485
rect -333 485 -299 504
rect -333 413 -299 425
rect -333 341 -299 357
rect -333 269 -299 289
rect -333 197 -299 221
rect -333 125 -299 153
rect -333 53 -299 85
rect -333 -17 -299 17
rect -333 -85 -299 -53
rect -333 -153 -299 -125
rect -333 -221 -299 -197
rect -333 -289 -299 -269
rect -333 -357 -299 -341
rect -333 -425 -299 -413
rect -333 -504 -299 -485
rect -175 485 -141 504
rect -175 413 -141 425
rect -175 341 -141 357
rect -175 269 -141 289
rect -175 197 -141 221
rect -175 125 -141 153
rect -175 53 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -53
rect -175 -153 -141 -125
rect -175 -221 -141 -197
rect -175 -289 -141 -269
rect -175 -357 -141 -341
rect -175 -425 -141 -413
rect -175 -504 -141 -485
rect -17 485 17 504
rect -17 413 17 425
rect -17 341 17 357
rect -17 269 17 289
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -289 17 -269
rect -17 -357 17 -341
rect -17 -425 17 -413
rect -17 -504 17 -485
rect 141 485 175 504
rect 141 413 175 425
rect 141 341 175 357
rect 141 269 175 289
rect 141 197 175 221
rect 141 125 175 153
rect 141 53 175 85
rect 141 -17 175 17
rect 141 -85 175 -53
rect 141 -153 175 -125
rect 141 -221 175 -197
rect 141 -289 175 -269
rect 141 -357 175 -341
rect 141 -425 175 -413
rect 141 -504 175 -485
rect 299 485 333 504
rect 299 413 333 425
rect 299 341 333 357
rect 299 269 333 289
rect 299 197 333 221
rect 299 125 333 153
rect 299 53 333 85
rect 299 -17 333 17
rect 299 -85 333 -53
rect 299 -153 333 -125
rect 299 -221 333 -197
rect 299 -289 333 -269
rect 299 -357 333 -341
rect 299 -425 333 -413
rect 299 -504 333 -485
rect 457 485 491 504
rect 457 413 491 425
rect 457 341 491 357
rect 457 269 491 289
rect 457 197 491 221
rect 457 125 491 153
rect 457 53 491 85
rect 457 -17 491 17
rect 457 -85 491 -53
rect 457 -153 491 -125
rect 457 -221 491 -197
rect 457 -289 491 -269
rect 457 -357 491 -341
rect 457 -425 491 -413
rect 457 -504 491 -485
rect 615 485 649 504
rect 615 413 649 425
rect 615 341 649 357
rect 615 269 649 289
rect 615 197 649 221
rect 615 125 649 153
rect 615 53 649 85
rect 615 -17 649 17
rect 615 -85 649 -53
rect 615 -153 649 -125
rect 615 -221 649 -197
rect 615 -289 649 -269
rect 615 -357 649 -341
rect 615 -425 649 -413
rect 615 -504 649 -485
rect 773 485 807 504
rect 773 413 807 425
rect 773 341 807 357
rect 773 269 807 289
rect 773 197 807 221
rect 773 125 807 153
rect 773 53 807 85
rect 773 -17 807 17
rect 773 -85 807 -53
rect 773 -153 807 -125
rect 773 -221 807 -197
rect 773 -289 807 -269
rect 773 -357 807 -341
rect 773 -425 807 -413
rect 773 -504 807 -485
rect 931 485 965 504
rect 931 413 965 425
rect 931 341 965 357
rect 931 269 965 289
rect 931 197 965 221
rect 931 125 965 153
rect 931 53 965 85
rect 931 -17 965 17
rect 931 -85 965 -53
rect 931 -153 965 -125
rect 931 -221 965 -197
rect 931 -289 965 -269
rect 931 -357 965 -341
rect 931 -425 965 -413
rect 931 -504 965 -485
rect 1089 485 1123 504
rect 1089 413 1123 425
rect 1089 341 1123 357
rect 1089 269 1123 289
rect 1089 197 1123 221
rect 1089 125 1123 153
rect 1089 53 1123 85
rect 1089 -17 1123 17
rect 1089 -85 1123 -53
rect 1089 -153 1123 -125
rect 1089 -221 1123 -197
rect 1089 -289 1123 -269
rect 1089 -357 1123 -341
rect 1089 -425 1123 -413
rect 1089 -504 1123 -485
rect 1247 485 1281 504
rect 1247 413 1281 425
rect 1247 341 1281 357
rect 1247 269 1281 289
rect 1247 197 1281 221
rect 1247 125 1281 153
rect 1247 53 1281 85
rect 1247 -17 1281 17
rect 1247 -85 1281 -53
rect 1247 -153 1281 -125
rect 1247 -221 1281 -197
rect 1247 -289 1281 -269
rect 1247 -357 1281 -341
rect 1247 -425 1281 -413
rect 1247 -504 1281 -485
rect 1405 485 1439 504
rect 1405 413 1439 425
rect 1405 341 1439 357
rect 1405 269 1439 289
rect 1405 197 1439 221
rect 1405 125 1439 153
rect 1405 53 1439 85
rect 1405 -17 1439 17
rect 1405 -85 1439 -53
rect 1405 -153 1439 -125
rect 1405 -221 1439 -197
rect 1405 -289 1439 -269
rect 1405 -357 1439 -341
rect 1405 -425 1439 -413
rect 1405 -504 1439 -485
rect 1563 485 1597 504
rect 1563 413 1597 425
rect 1563 341 1597 357
rect 1563 269 1597 289
rect 1563 197 1597 221
rect 1563 125 1597 153
rect 1563 53 1597 85
rect 1563 -17 1597 17
rect 1563 -85 1597 -53
rect 1563 -153 1597 -125
rect 1563 -221 1597 -197
rect 1563 -289 1597 -269
rect 1563 -357 1597 -341
rect 1563 -425 1597 -413
rect 1563 -504 1597 -485
rect -1537 -572 -1518 -538
rect -1484 -572 -1465 -538
rect -1379 -572 -1360 -538
rect -1326 -572 -1307 -538
rect -1221 -572 -1202 -538
rect -1168 -572 -1149 -538
rect -1063 -572 -1044 -538
rect -1010 -572 -991 -538
rect -905 -572 -886 -538
rect -852 -572 -833 -538
rect -747 -572 -728 -538
rect -694 -572 -675 -538
rect -589 -572 -570 -538
rect -536 -572 -517 -538
rect -431 -572 -412 -538
rect -378 -572 -359 -538
rect -273 -572 -254 -538
rect -220 -572 -201 -538
rect -115 -572 -96 -538
rect -62 -572 -43 -538
rect 43 -572 62 -538
rect 96 -572 115 -538
rect 201 -572 220 -538
rect 254 -572 273 -538
rect 359 -572 378 -538
rect 412 -572 431 -538
rect 517 -572 536 -538
rect 570 -572 589 -538
rect 675 -572 694 -538
rect 728 -572 747 -538
rect 833 -572 852 -538
rect 886 -572 905 -538
rect 991 -572 1010 -538
rect 1044 -572 1063 -538
rect 1149 -572 1168 -538
rect 1202 -572 1221 -538
rect 1307 -572 1326 -538
rect 1360 -572 1379 -538
rect 1465 -572 1484 -538
rect 1518 -572 1537 -538
<< viali >>
rect -1597 459 -1563 485
rect -1597 451 -1563 459
rect -1597 391 -1563 413
rect -1597 379 -1563 391
rect -1597 323 -1563 341
rect -1597 307 -1563 323
rect -1597 255 -1563 269
rect -1597 235 -1563 255
rect -1597 187 -1563 197
rect -1597 163 -1563 187
rect -1597 119 -1563 125
rect -1597 91 -1563 119
rect -1597 51 -1563 53
rect -1597 19 -1563 51
rect -1597 -51 -1563 -19
rect -1597 -53 -1563 -51
rect -1597 -119 -1563 -91
rect -1597 -125 -1563 -119
rect -1597 -187 -1563 -163
rect -1597 -197 -1563 -187
rect -1597 -255 -1563 -235
rect -1597 -269 -1563 -255
rect -1597 -323 -1563 -307
rect -1597 -341 -1563 -323
rect -1597 -391 -1563 -379
rect -1597 -413 -1563 -391
rect -1597 -459 -1563 -451
rect -1597 -485 -1563 -459
rect -1439 459 -1405 485
rect -1439 451 -1405 459
rect -1439 391 -1405 413
rect -1439 379 -1405 391
rect -1439 323 -1405 341
rect -1439 307 -1405 323
rect -1439 255 -1405 269
rect -1439 235 -1405 255
rect -1439 187 -1405 197
rect -1439 163 -1405 187
rect -1439 119 -1405 125
rect -1439 91 -1405 119
rect -1439 51 -1405 53
rect -1439 19 -1405 51
rect -1439 -51 -1405 -19
rect -1439 -53 -1405 -51
rect -1439 -119 -1405 -91
rect -1439 -125 -1405 -119
rect -1439 -187 -1405 -163
rect -1439 -197 -1405 -187
rect -1439 -255 -1405 -235
rect -1439 -269 -1405 -255
rect -1439 -323 -1405 -307
rect -1439 -341 -1405 -323
rect -1439 -391 -1405 -379
rect -1439 -413 -1405 -391
rect -1439 -459 -1405 -451
rect -1439 -485 -1405 -459
rect -1281 459 -1247 485
rect -1281 451 -1247 459
rect -1281 391 -1247 413
rect -1281 379 -1247 391
rect -1281 323 -1247 341
rect -1281 307 -1247 323
rect -1281 255 -1247 269
rect -1281 235 -1247 255
rect -1281 187 -1247 197
rect -1281 163 -1247 187
rect -1281 119 -1247 125
rect -1281 91 -1247 119
rect -1281 51 -1247 53
rect -1281 19 -1247 51
rect -1281 -51 -1247 -19
rect -1281 -53 -1247 -51
rect -1281 -119 -1247 -91
rect -1281 -125 -1247 -119
rect -1281 -187 -1247 -163
rect -1281 -197 -1247 -187
rect -1281 -255 -1247 -235
rect -1281 -269 -1247 -255
rect -1281 -323 -1247 -307
rect -1281 -341 -1247 -323
rect -1281 -391 -1247 -379
rect -1281 -413 -1247 -391
rect -1281 -459 -1247 -451
rect -1281 -485 -1247 -459
rect -1123 459 -1089 485
rect -1123 451 -1089 459
rect -1123 391 -1089 413
rect -1123 379 -1089 391
rect -1123 323 -1089 341
rect -1123 307 -1089 323
rect -1123 255 -1089 269
rect -1123 235 -1089 255
rect -1123 187 -1089 197
rect -1123 163 -1089 187
rect -1123 119 -1089 125
rect -1123 91 -1089 119
rect -1123 51 -1089 53
rect -1123 19 -1089 51
rect -1123 -51 -1089 -19
rect -1123 -53 -1089 -51
rect -1123 -119 -1089 -91
rect -1123 -125 -1089 -119
rect -1123 -187 -1089 -163
rect -1123 -197 -1089 -187
rect -1123 -255 -1089 -235
rect -1123 -269 -1089 -255
rect -1123 -323 -1089 -307
rect -1123 -341 -1089 -323
rect -1123 -391 -1089 -379
rect -1123 -413 -1089 -391
rect -1123 -459 -1089 -451
rect -1123 -485 -1089 -459
rect -965 459 -931 485
rect -965 451 -931 459
rect -965 391 -931 413
rect -965 379 -931 391
rect -965 323 -931 341
rect -965 307 -931 323
rect -965 255 -931 269
rect -965 235 -931 255
rect -965 187 -931 197
rect -965 163 -931 187
rect -965 119 -931 125
rect -965 91 -931 119
rect -965 51 -931 53
rect -965 19 -931 51
rect -965 -51 -931 -19
rect -965 -53 -931 -51
rect -965 -119 -931 -91
rect -965 -125 -931 -119
rect -965 -187 -931 -163
rect -965 -197 -931 -187
rect -965 -255 -931 -235
rect -965 -269 -931 -255
rect -965 -323 -931 -307
rect -965 -341 -931 -323
rect -965 -391 -931 -379
rect -965 -413 -931 -391
rect -965 -459 -931 -451
rect -965 -485 -931 -459
rect -807 459 -773 485
rect -807 451 -773 459
rect -807 391 -773 413
rect -807 379 -773 391
rect -807 323 -773 341
rect -807 307 -773 323
rect -807 255 -773 269
rect -807 235 -773 255
rect -807 187 -773 197
rect -807 163 -773 187
rect -807 119 -773 125
rect -807 91 -773 119
rect -807 51 -773 53
rect -807 19 -773 51
rect -807 -51 -773 -19
rect -807 -53 -773 -51
rect -807 -119 -773 -91
rect -807 -125 -773 -119
rect -807 -187 -773 -163
rect -807 -197 -773 -187
rect -807 -255 -773 -235
rect -807 -269 -773 -255
rect -807 -323 -773 -307
rect -807 -341 -773 -323
rect -807 -391 -773 -379
rect -807 -413 -773 -391
rect -807 -459 -773 -451
rect -807 -485 -773 -459
rect -649 459 -615 485
rect -649 451 -615 459
rect -649 391 -615 413
rect -649 379 -615 391
rect -649 323 -615 341
rect -649 307 -615 323
rect -649 255 -615 269
rect -649 235 -615 255
rect -649 187 -615 197
rect -649 163 -615 187
rect -649 119 -615 125
rect -649 91 -615 119
rect -649 51 -615 53
rect -649 19 -615 51
rect -649 -51 -615 -19
rect -649 -53 -615 -51
rect -649 -119 -615 -91
rect -649 -125 -615 -119
rect -649 -187 -615 -163
rect -649 -197 -615 -187
rect -649 -255 -615 -235
rect -649 -269 -615 -255
rect -649 -323 -615 -307
rect -649 -341 -615 -323
rect -649 -391 -615 -379
rect -649 -413 -615 -391
rect -649 -459 -615 -451
rect -649 -485 -615 -459
rect -491 459 -457 485
rect -491 451 -457 459
rect -491 391 -457 413
rect -491 379 -457 391
rect -491 323 -457 341
rect -491 307 -457 323
rect -491 255 -457 269
rect -491 235 -457 255
rect -491 187 -457 197
rect -491 163 -457 187
rect -491 119 -457 125
rect -491 91 -457 119
rect -491 51 -457 53
rect -491 19 -457 51
rect -491 -51 -457 -19
rect -491 -53 -457 -51
rect -491 -119 -457 -91
rect -491 -125 -457 -119
rect -491 -187 -457 -163
rect -491 -197 -457 -187
rect -491 -255 -457 -235
rect -491 -269 -457 -255
rect -491 -323 -457 -307
rect -491 -341 -457 -323
rect -491 -391 -457 -379
rect -491 -413 -457 -391
rect -491 -459 -457 -451
rect -491 -485 -457 -459
rect -333 459 -299 485
rect -333 451 -299 459
rect -333 391 -299 413
rect -333 379 -299 391
rect -333 323 -299 341
rect -333 307 -299 323
rect -333 255 -299 269
rect -333 235 -299 255
rect -333 187 -299 197
rect -333 163 -299 187
rect -333 119 -299 125
rect -333 91 -299 119
rect -333 51 -299 53
rect -333 19 -299 51
rect -333 -51 -299 -19
rect -333 -53 -299 -51
rect -333 -119 -299 -91
rect -333 -125 -299 -119
rect -333 -187 -299 -163
rect -333 -197 -299 -187
rect -333 -255 -299 -235
rect -333 -269 -299 -255
rect -333 -323 -299 -307
rect -333 -341 -299 -323
rect -333 -391 -299 -379
rect -333 -413 -299 -391
rect -333 -459 -299 -451
rect -333 -485 -299 -459
rect -175 459 -141 485
rect -175 451 -141 459
rect -175 391 -141 413
rect -175 379 -141 391
rect -175 323 -141 341
rect -175 307 -141 323
rect -175 255 -141 269
rect -175 235 -141 255
rect -175 187 -141 197
rect -175 163 -141 187
rect -175 119 -141 125
rect -175 91 -141 119
rect -175 51 -141 53
rect -175 19 -141 51
rect -175 -51 -141 -19
rect -175 -53 -141 -51
rect -175 -119 -141 -91
rect -175 -125 -141 -119
rect -175 -187 -141 -163
rect -175 -197 -141 -187
rect -175 -255 -141 -235
rect -175 -269 -141 -255
rect -175 -323 -141 -307
rect -175 -341 -141 -323
rect -175 -391 -141 -379
rect -175 -413 -141 -391
rect -175 -459 -141 -451
rect -175 -485 -141 -459
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect 141 459 175 485
rect 141 451 175 459
rect 141 391 175 413
rect 141 379 175 391
rect 141 323 175 341
rect 141 307 175 323
rect 141 255 175 269
rect 141 235 175 255
rect 141 187 175 197
rect 141 163 175 187
rect 141 119 175 125
rect 141 91 175 119
rect 141 51 175 53
rect 141 19 175 51
rect 141 -51 175 -19
rect 141 -53 175 -51
rect 141 -119 175 -91
rect 141 -125 175 -119
rect 141 -187 175 -163
rect 141 -197 175 -187
rect 141 -255 175 -235
rect 141 -269 175 -255
rect 141 -323 175 -307
rect 141 -341 175 -323
rect 141 -391 175 -379
rect 141 -413 175 -391
rect 141 -459 175 -451
rect 141 -485 175 -459
rect 299 459 333 485
rect 299 451 333 459
rect 299 391 333 413
rect 299 379 333 391
rect 299 323 333 341
rect 299 307 333 323
rect 299 255 333 269
rect 299 235 333 255
rect 299 187 333 197
rect 299 163 333 187
rect 299 119 333 125
rect 299 91 333 119
rect 299 51 333 53
rect 299 19 333 51
rect 299 -51 333 -19
rect 299 -53 333 -51
rect 299 -119 333 -91
rect 299 -125 333 -119
rect 299 -187 333 -163
rect 299 -197 333 -187
rect 299 -255 333 -235
rect 299 -269 333 -255
rect 299 -323 333 -307
rect 299 -341 333 -323
rect 299 -391 333 -379
rect 299 -413 333 -391
rect 299 -459 333 -451
rect 299 -485 333 -459
rect 457 459 491 485
rect 457 451 491 459
rect 457 391 491 413
rect 457 379 491 391
rect 457 323 491 341
rect 457 307 491 323
rect 457 255 491 269
rect 457 235 491 255
rect 457 187 491 197
rect 457 163 491 187
rect 457 119 491 125
rect 457 91 491 119
rect 457 51 491 53
rect 457 19 491 51
rect 457 -51 491 -19
rect 457 -53 491 -51
rect 457 -119 491 -91
rect 457 -125 491 -119
rect 457 -187 491 -163
rect 457 -197 491 -187
rect 457 -255 491 -235
rect 457 -269 491 -255
rect 457 -323 491 -307
rect 457 -341 491 -323
rect 457 -391 491 -379
rect 457 -413 491 -391
rect 457 -459 491 -451
rect 457 -485 491 -459
rect 615 459 649 485
rect 615 451 649 459
rect 615 391 649 413
rect 615 379 649 391
rect 615 323 649 341
rect 615 307 649 323
rect 615 255 649 269
rect 615 235 649 255
rect 615 187 649 197
rect 615 163 649 187
rect 615 119 649 125
rect 615 91 649 119
rect 615 51 649 53
rect 615 19 649 51
rect 615 -51 649 -19
rect 615 -53 649 -51
rect 615 -119 649 -91
rect 615 -125 649 -119
rect 615 -187 649 -163
rect 615 -197 649 -187
rect 615 -255 649 -235
rect 615 -269 649 -255
rect 615 -323 649 -307
rect 615 -341 649 -323
rect 615 -391 649 -379
rect 615 -413 649 -391
rect 615 -459 649 -451
rect 615 -485 649 -459
rect 773 459 807 485
rect 773 451 807 459
rect 773 391 807 413
rect 773 379 807 391
rect 773 323 807 341
rect 773 307 807 323
rect 773 255 807 269
rect 773 235 807 255
rect 773 187 807 197
rect 773 163 807 187
rect 773 119 807 125
rect 773 91 807 119
rect 773 51 807 53
rect 773 19 807 51
rect 773 -51 807 -19
rect 773 -53 807 -51
rect 773 -119 807 -91
rect 773 -125 807 -119
rect 773 -187 807 -163
rect 773 -197 807 -187
rect 773 -255 807 -235
rect 773 -269 807 -255
rect 773 -323 807 -307
rect 773 -341 807 -323
rect 773 -391 807 -379
rect 773 -413 807 -391
rect 773 -459 807 -451
rect 773 -485 807 -459
rect 931 459 965 485
rect 931 451 965 459
rect 931 391 965 413
rect 931 379 965 391
rect 931 323 965 341
rect 931 307 965 323
rect 931 255 965 269
rect 931 235 965 255
rect 931 187 965 197
rect 931 163 965 187
rect 931 119 965 125
rect 931 91 965 119
rect 931 51 965 53
rect 931 19 965 51
rect 931 -51 965 -19
rect 931 -53 965 -51
rect 931 -119 965 -91
rect 931 -125 965 -119
rect 931 -187 965 -163
rect 931 -197 965 -187
rect 931 -255 965 -235
rect 931 -269 965 -255
rect 931 -323 965 -307
rect 931 -341 965 -323
rect 931 -391 965 -379
rect 931 -413 965 -391
rect 931 -459 965 -451
rect 931 -485 965 -459
rect 1089 459 1123 485
rect 1089 451 1123 459
rect 1089 391 1123 413
rect 1089 379 1123 391
rect 1089 323 1123 341
rect 1089 307 1123 323
rect 1089 255 1123 269
rect 1089 235 1123 255
rect 1089 187 1123 197
rect 1089 163 1123 187
rect 1089 119 1123 125
rect 1089 91 1123 119
rect 1089 51 1123 53
rect 1089 19 1123 51
rect 1089 -51 1123 -19
rect 1089 -53 1123 -51
rect 1089 -119 1123 -91
rect 1089 -125 1123 -119
rect 1089 -187 1123 -163
rect 1089 -197 1123 -187
rect 1089 -255 1123 -235
rect 1089 -269 1123 -255
rect 1089 -323 1123 -307
rect 1089 -341 1123 -323
rect 1089 -391 1123 -379
rect 1089 -413 1123 -391
rect 1089 -459 1123 -451
rect 1089 -485 1123 -459
rect 1247 459 1281 485
rect 1247 451 1281 459
rect 1247 391 1281 413
rect 1247 379 1281 391
rect 1247 323 1281 341
rect 1247 307 1281 323
rect 1247 255 1281 269
rect 1247 235 1281 255
rect 1247 187 1281 197
rect 1247 163 1281 187
rect 1247 119 1281 125
rect 1247 91 1281 119
rect 1247 51 1281 53
rect 1247 19 1281 51
rect 1247 -51 1281 -19
rect 1247 -53 1281 -51
rect 1247 -119 1281 -91
rect 1247 -125 1281 -119
rect 1247 -187 1281 -163
rect 1247 -197 1281 -187
rect 1247 -255 1281 -235
rect 1247 -269 1281 -255
rect 1247 -323 1281 -307
rect 1247 -341 1281 -323
rect 1247 -391 1281 -379
rect 1247 -413 1281 -391
rect 1247 -459 1281 -451
rect 1247 -485 1281 -459
rect 1405 459 1439 485
rect 1405 451 1439 459
rect 1405 391 1439 413
rect 1405 379 1439 391
rect 1405 323 1439 341
rect 1405 307 1439 323
rect 1405 255 1439 269
rect 1405 235 1439 255
rect 1405 187 1439 197
rect 1405 163 1439 187
rect 1405 119 1439 125
rect 1405 91 1439 119
rect 1405 51 1439 53
rect 1405 19 1439 51
rect 1405 -51 1439 -19
rect 1405 -53 1439 -51
rect 1405 -119 1439 -91
rect 1405 -125 1439 -119
rect 1405 -187 1439 -163
rect 1405 -197 1439 -187
rect 1405 -255 1439 -235
rect 1405 -269 1439 -255
rect 1405 -323 1439 -307
rect 1405 -341 1439 -323
rect 1405 -391 1439 -379
rect 1405 -413 1439 -391
rect 1405 -459 1439 -451
rect 1405 -485 1439 -459
rect 1563 459 1597 485
rect 1563 451 1597 459
rect 1563 391 1597 413
rect 1563 379 1597 391
rect 1563 323 1597 341
rect 1563 307 1597 323
rect 1563 255 1597 269
rect 1563 235 1597 255
rect 1563 187 1597 197
rect 1563 163 1597 187
rect 1563 119 1597 125
rect 1563 91 1597 119
rect 1563 51 1597 53
rect 1563 19 1597 51
rect 1563 -51 1597 -19
rect 1563 -53 1597 -51
rect 1563 -119 1597 -91
rect 1563 -125 1597 -119
rect 1563 -187 1597 -163
rect 1563 -197 1597 -187
rect 1563 -255 1597 -235
rect 1563 -269 1597 -255
rect 1563 -323 1597 -307
rect 1563 -341 1597 -323
rect 1563 -391 1597 -379
rect 1563 -413 1597 -391
rect 1563 -459 1597 -451
rect 1563 -485 1597 -459
<< metal1 >>
rect -1603 485 -1557 500
rect -1603 451 -1597 485
rect -1563 451 -1557 485
rect -1603 413 -1557 451
rect -1603 379 -1597 413
rect -1563 379 -1557 413
rect -1603 341 -1557 379
rect -1603 307 -1597 341
rect -1563 307 -1557 341
rect -1603 269 -1557 307
rect -1603 235 -1597 269
rect -1563 235 -1557 269
rect -1603 197 -1557 235
rect -1603 163 -1597 197
rect -1563 163 -1557 197
rect -1603 125 -1557 163
rect -1603 91 -1597 125
rect -1563 91 -1557 125
rect -1603 53 -1557 91
rect -1603 19 -1597 53
rect -1563 19 -1557 53
rect -1603 -19 -1557 19
rect -1603 -53 -1597 -19
rect -1563 -53 -1557 -19
rect -1603 -91 -1557 -53
rect -1603 -125 -1597 -91
rect -1563 -125 -1557 -91
rect -1603 -163 -1557 -125
rect -1603 -197 -1597 -163
rect -1563 -197 -1557 -163
rect -1603 -235 -1557 -197
rect -1603 -269 -1597 -235
rect -1563 -269 -1557 -235
rect -1603 -307 -1557 -269
rect -1603 -341 -1597 -307
rect -1563 -341 -1557 -307
rect -1603 -379 -1557 -341
rect -1603 -413 -1597 -379
rect -1563 -413 -1557 -379
rect -1603 -451 -1557 -413
rect -1603 -485 -1597 -451
rect -1563 -485 -1557 -451
rect -1603 -500 -1557 -485
rect -1445 485 -1399 500
rect -1445 451 -1439 485
rect -1405 451 -1399 485
rect -1445 413 -1399 451
rect -1445 379 -1439 413
rect -1405 379 -1399 413
rect -1445 341 -1399 379
rect -1445 307 -1439 341
rect -1405 307 -1399 341
rect -1445 269 -1399 307
rect -1445 235 -1439 269
rect -1405 235 -1399 269
rect -1445 197 -1399 235
rect -1445 163 -1439 197
rect -1405 163 -1399 197
rect -1445 125 -1399 163
rect -1445 91 -1439 125
rect -1405 91 -1399 125
rect -1445 53 -1399 91
rect -1445 19 -1439 53
rect -1405 19 -1399 53
rect -1445 -19 -1399 19
rect -1445 -53 -1439 -19
rect -1405 -53 -1399 -19
rect -1445 -91 -1399 -53
rect -1445 -125 -1439 -91
rect -1405 -125 -1399 -91
rect -1445 -163 -1399 -125
rect -1445 -197 -1439 -163
rect -1405 -197 -1399 -163
rect -1445 -235 -1399 -197
rect -1445 -269 -1439 -235
rect -1405 -269 -1399 -235
rect -1445 -307 -1399 -269
rect -1445 -341 -1439 -307
rect -1405 -341 -1399 -307
rect -1445 -379 -1399 -341
rect -1445 -413 -1439 -379
rect -1405 -413 -1399 -379
rect -1445 -451 -1399 -413
rect -1445 -485 -1439 -451
rect -1405 -485 -1399 -451
rect -1445 -500 -1399 -485
rect -1287 485 -1241 500
rect -1287 451 -1281 485
rect -1247 451 -1241 485
rect -1287 413 -1241 451
rect -1287 379 -1281 413
rect -1247 379 -1241 413
rect -1287 341 -1241 379
rect -1287 307 -1281 341
rect -1247 307 -1241 341
rect -1287 269 -1241 307
rect -1287 235 -1281 269
rect -1247 235 -1241 269
rect -1287 197 -1241 235
rect -1287 163 -1281 197
rect -1247 163 -1241 197
rect -1287 125 -1241 163
rect -1287 91 -1281 125
rect -1247 91 -1241 125
rect -1287 53 -1241 91
rect -1287 19 -1281 53
rect -1247 19 -1241 53
rect -1287 -19 -1241 19
rect -1287 -53 -1281 -19
rect -1247 -53 -1241 -19
rect -1287 -91 -1241 -53
rect -1287 -125 -1281 -91
rect -1247 -125 -1241 -91
rect -1287 -163 -1241 -125
rect -1287 -197 -1281 -163
rect -1247 -197 -1241 -163
rect -1287 -235 -1241 -197
rect -1287 -269 -1281 -235
rect -1247 -269 -1241 -235
rect -1287 -307 -1241 -269
rect -1287 -341 -1281 -307
rect -1247 -341 -1241 -307
rect -1287 -379 -1241 -341
rect -1287 -413 -1281 -379
rect -1247 -413 -1241 -379
rect -1287 -451 -1241 -413
rect -1287 -485 -1281 -451
rect -1247 -485 -1241 -451
rect -1287 -500 -1241 -485
rect -1129 485 -1083 500
rect -1129 451 -1123 485
rect -1089 451 -1083 485
rect -1129 413 -1083 451
rect -1129 379 -1123 413
rect -1089 379 -1083 413
rect -1129 341 -1083 379
rect -1129 307 -1123 341
rect -1089 307 -1083 341
rect -1129 269 -1083 307
rect -1129 235 -1123 269
rect -1089 235 -1083 269
rect -1129 197 -1083 235
rect -1129 163 -1123 197
rect -1089 163 -1083 197
rect -1129 125 -1083 163
rect -1129 91 -1123 125
rect -1089 91 -1083 125
rect -1129 53 -1083 91
rect -1129 19 -1123 53
rect -1089 19 -1083 53
rect -1129 -19 -1083 19
rect -1129 -53 -1123 -19
rect -1089 -53 -1083 -19
rect -1129 -91 -1083 -53
rect -1129 -125 -1123 -91
rect -1089 -125 -1083 -91
rect -1129 -163 -1083 -125
rect -1129 -197 -1123 -163
rect -1089 -197 -1083 -163
rect -1129 -235 -1083 -197
rect -1129 -269 -1123 -235
rect -1089 -269 -1083 -235
rect -1129 -307 -1083 -269
rect -1129 -341 -1123 -307
rect -1089 -341 -1083 -307
rect -1129 -379 -1083 -341
rect -1129 -413 -1123 -379
rect -1089 -413 -1083 -379
rect -1129 -451 -1083 -413
rect -1129 -485 -1123 -451
rect -1089 -485 -1083 -451
rect -1129 -500 -1083 -485
rect -971 485 -925 500
rect -971 451 -965 485
rect -931 451 -925 485
rect -971 413 -925 451
rect -971 379 -965 413
rect -931 379 -925 413
rect -971 341 -925 379
rect -971 307 -965 341
rect -931 307 -925 341
rect -971 269 -925 307
rect -971 235 -965 269
rect -931 235 -925 269
rect -971 197 -925 235
rect -971 163 -965 197
rect -931 163 -925 197
rect -971 125 -925 163
rect -971 91 -965 125
rect -931 91 -925 125
rect -971 53 -925 91
rect -971 19 -965 53
rect -931 19 -925 53
rect -971 -19 -925 19
rect -971 -53 -965 -19
rect -931 -53 -925 -19
rect -971 -91 -925 -53
rect -971 -125 -965 -91
rect -931 -125 -925 -91
rect -971 -163 -925 -125
rect -971 -197 -965 -163
rect -931 -197 -925 -163
rect -971 -235 -925 -197
rect -971 -269 -965 -235
rect -931 -269 -925 -235
rect -971 -307 -925 -269
rect -971 -341 -965 -307
rect -931 -341 -925 -307
rect -971 -379 -925 -341
rect -971 -413 -965 -379
rect -931 -413 -925 -379
rect -971 -451 -925 -413
rect -971 -485 -965 -451
rect -931 -485 -925 -451
rect -971 -500 -925 -485
rect -813 485 -767 500
rect -813 451 -807 485
rect -773 451 -767 485
rect -813 413 -767 451
rect -813 379 -807 413
rect -773 379 -767 413
rect -813 341 -767 379
rect -813 307 -807 341
rect -773 307 -767 341
rect -813 269 -767 307
rect -813 235 -807 269
rect -773 235 -767 269
rect -813 197 -767 235
rect -813 163 -807 197
rect -773 163 -767 197
rect -813 125 -767 163
rect -813 91 -807 125
rect -773 91 -767 125
rect -813 53 -767 91
rect -813 19 -807 53
rect -773 19 -767 53
rect -813 -19 -767 19
rect -813 -53 -807 -19
rect -773 -53 -767 -19
rect -813 -91 -767 -53
rect -813 -125 -807 -91
rect -773 -125 -767 -91
rect -813 -163 -767 -125
rect -813 -197 -807 -163
rect -773 -197 -767 -163
rect -813 -235 -767 -197
rect -813 -269 -807 -235
rect -773 -269 -767 -235
rect -813 -307 -767 -269
rect -813 -341 -807 -307
rect -773 -341 -767 -307
rect -813 -379 -767 -341
rect -813 -413 -807 -379
rect -773 -413 -767 -379
rect -813 -451 -767 -413
rect -813 -485 -807 -451
rect -773 -485 -767 -451
rect -813 -500 -767 -485
rect -655 485 -609 500
rect -655 451 -649 485
rect -615 451 -609 485
rect -655 413 -609 451
rect -655 379 -649 413
rect -615 379 -609 413
rect -655 341 -609 379
rect -655 307 -649 341
rect -615 307 -609 341
rect -655 269 -609 307
rect -655 235 -649 269
rect -615 235 -609 269
rect -655 197 -609 235
rect -655 163 -649 197
rect -615 163 -609 197
rect -655 125 -609 163
rect -655 91 -649 125
rect -615 91 -609 125
rect -655 53 -609 91
rect -655 19 -649 53
rect -615 19 -609 53
rect -655 -19 -609 19
rect -655 -53 -649 -19
rect -615 -53 -609 -19
rect -655 -91 -609 -53
rect -655 -125 -649 -91
rect -615 -125 -609 -91
rect -655 -163 -609 -125
rect -655 -197 -649 -163
rect -615 -197 -609 -163
rect -655 -235 -609 -197
rect -655 -269 -649 -235
rect -615 -269 -609 -235
rect -655 -307 -609 -269
rect -655 -341 -649 -307
rect -615 -341 -609 -307
rect -655 -379 -609 -341
rect -655 -413 -649 -379
rect -615 -413 -609 -379
rect -655 -451 -609 -413
rect -655 -485 -649 -451
rect -615 -485 -609 -451
rect -655 -500 -609 -485
rect -497 485 -451 500
rect -497 451 -491 485
rect -457 451 -451 485
rect -497 413 -451 451
rect -497 379 -491 413
rect -457 379 -451 413
rect -497 341 -451 379
rect -497 307 -491 341
rect -457 307 -451 341
rect -497 269 -451 307
rect -497 235 -491 269
rect -457 235 -451 269
rect -497 197 -451 235
rect -497 163 -491 197
rect -457 163 -451 197
rect -497 125 -451 163
rect -497 91 -491 125
rect -457 91 -451 125
rect -497 53 -451 91
rect -497 19 -491 53
rect -457 19 -451 53
rect -497 -19 -451 19
rect -497 -53 -491 -19
rect -457 -53 -451 -19
rect -497 -91 -451 -53
rect -497 -125 -491 -91
rect -457 -125 -451 -91
rect -497 -163 -451 -125
rect -497 -197 -491 -163
rect -457 -197 -451 -163
rect -497 -235 -451 -197
rect -497 -269 -491 -235
rect -457 -269 -451 -235
rect -497 -307 -451 -269
rect -497 -341 -491 -307
rect -457 -341 -451 -307
rect -497 -379 -451 -341
rect -497 -413 -491 -379
rect -457 -413 -451 -379
rect -497 -451 -451 -413
rect -497 -485 -491 -451
rect -457 -485 -451 -451
rect -497 -500 -451 -485
rect -339 485 -293 500
rect -339 451 -333 485
rect -299 451 -293 485
rect -339 413 -293 451
rect -339 379 -333 413
rect -299 379 -293 413
rect -339 341 -293 379
rect -339 307 -333 341
rect -299 307 -293 341
rect -339 269 -293 307
rect -339 235 -333 269
rect -299 235 -293 269
rect -339 197 -293 235
rect -339 163 -333 197
rect -299 163 -293 197
rect -339 125 -293 163
rect -339 91 -333 125
rect -299 91 -293 125
rect -339 53 -293 91
rect -339 19 -333 53
rect -299 19 -293 53
rect -339 -19 -293 19
rect -339 -53 -333 -19
rect -299 -53 -293 -19
rect -339 -91 -293 -53
rect -339 -125 -333 -91
rect -299 -125 -293 -91
rect -339 -163 -293 -125
rect -339 -197 -333 -163
rect -299 -197 -293 -163
rect -339 -235 -293 -197
rect -339 -269 -333 -235
rect -299 -269 -293 -235
rect -339 -307 -293 -269
rect -339 -341 -333 -307
rect -299 -341 -293 -307
rect -339 -379 -293 -341
rect -339 -413 -333 -379
rect -299 -413 -293 -379
rect -339 -451 -293 -413
rect -339 -485 -333 -451
rect -299 -485 -293 -451
rect -339 -500 -293 -485
rect -181 485 -135 500
rect -181 451 -175 485
rect -141 451 -135 485
rect -181 413 -135 451
rect -181 379 -175 413
rect -141 379 -135 413
rect -181 341 -135 379
rect -181 307 -175 341
rect -141 307 -135 341
rect -181 269 -135 307
rect -181 235 -175 269
rect -141 235 -135 269
rect -181 197 -135 235
rect -181 163 -175 197
rect -141 163 -135 197
rect -181 125 -135 163
rect -181 91 -175 125
rect -141 91 -135 125
rect -181 53 -135 91
rect -181 19 -175 53
rect -141 19 -135 53
rect -181 -19 -135 19
rect -181 -53 -175 -19
rect -141 -53 -135 -19
rect -181 -91 -135 -53
rect -181 -125 -175 -91
rect -141 -125 -135 -91
rect -181 -163 -135 -125
rect -181 -197 -175 -163
rect -141 -197 -135 -163
rect -181 -235 -135 -197
rect -181 -269 -175 -235
rect -141 -269 -135 -235
rect -181 -307 -135 -269
rect -181 -341 -175 -307
rect -141 -341 -135 -307
rect -181 -379 -135 -341
rect -181 -413 -175 -379
rect -141 -413 -135 -379
rect -181 -451 -135 -413
rect -181 -485 -175 -451
rect -141 -485 -135 -451
rect -181 -500 -135 -485
rect -23 485 23 500
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -500 23 -485
rect 135 485 181 500
rect 135 451 141 485
rect 175 451 181 485
rect 135 413 181 451
rect 135 379 141 413
rect 175 379 181 413
rect 135 341 181 379
rect 135 307 141 341
rect 175 307 181 341
rect 135 269 181 307
rect 135 235 141 269
rect 175 235 181 269
rect 135 197 181 235
rect 135 163 141 197
rect 175 163 181 197
rect 135 125 181 163
rect 135 91 141 125
rect 175 91 181 125
rect 135 53 181 91
rect 135 19 141 53
rect 175 19 181 53
rect 135 -19 181 19
rect 135 -53 141 -19
rect 175 -53 181 -19
rect 135 -91 181 -53
rect 135 -125 141 -91
rect 175 -125 181 -91
rect 135 -163 181 -125
rect 135 -197 141 -163
rect 175 -197 181 -163
rect 135 -235 181 -197
rect 135 -269 141 -235
rect 175 -269 181 -235
rect 135 -307 181 -269
rect 135 -341 141 -307
rect 175 -341 181 -307
rect 135 -379 181 -341
rect 135 -413 141 -379
rect 175 -413 181 -379
rect 135 -451 181 -413
rect 135 -485 141 -451
rect 175 -485 181 -451
rect 135 -500 181 -485
rect 293 485 339 500
rect 293 451 299 485
rect 333 451 339 485
rect 293 413 339 451
rect 293 379 299 413
rect 333 379 339 413
rect 293 341 339 379
rect 293 307 299 341
rect 333 307 339 341
rect 293 269 339 307
rect 293 235 299 269
rect 333 235 339 269
rect 293 197 339 235
rect 293 163 299 197
rect 333 163 339 197
rect 293 125 339 163
rect 293 91 299 125
rect 333 91 339 125
rect 293 53 339 91
rect 293 19 299 53
rect 333 19 339 53
rect 293 -19 339 19
rect 293 -53 299 -19
rect 333 -53 339 -19
rect 293 -91 339 -53
rect 293 -125 299 -91
rect 333 -125 339 -91
rect 293 -163 339 -125
rect 293 -197 299 -163
rect 333 -197 339 -163
rect 293 -235 339 -197
rect 293 -269 299 -235
rect 333 -269 339 -235
rect 293 -307 339 -269
rect 293 -341 299 -307
rect 333 -341 339 -307
rect 293 -379 339 -341
rect 293 -413 299 -379
rect 333 -413 339 -379
rect 293 -451 339 -413
rect 293 -485 299 -451
rect 333 -485 339 -451
rect 293 -500 339 -485
rect 451 485 497 500
rect 451 451 457 485
rect 491 451 497 485
rect 451 413 497 451
rect 451 379 457 413
rect 491 379 497 413
rect 451 341 497 379
rect 451 307 457 341
rect 491 307 497 341
rect 451 269 497 307
rect 451 235 457 269
rect 491 235 497 269
rect 451 197 497 235
rect 451 163 457 197
rect 491 163 497 197
rect 451 125 497 163
rect 451 91 457 125
rect 491 91 497 125
rect 451 53 497 91
rect 451 19 457 53
rect 491 19 497 53
rect 451 -19 497 19
rect 451 -53 457 -19
rect 491 -53 497 -19
rect 451 -91 497 -53
rect 451 -125 457 -91
rect 491 -125 497 -91
rect 451 -163 497 -125
rect 451 -197 457 -163
rect 491 -197 497 -163
rect 451 -235 497 -197
rect 451 -269 457 -235
rect 491 -269 497 -235
rect 451 -307 497 -269
rect 451 -341 457 -307
rect 491 -341 497 -307
rect 451 -379 497 -341
rect 451 -413 457 -379
rect 491 -413 497 -379
rect 451 -451 497 -413
rect 451 -485 457 -451
rect 491 -485 497 -451
rect 451 -500 497 -485
rect 609 485 655 500
rect 609 451 615 485
rect 649 451 655 485
rect 609 413 655 451
rect 609 379 615 413
rect 649 379 655 413
rect 609 341 655 379
rect 609 307 615 341
rect 649 307 655 341
rect 609 269 655 307
rect 609 235 615 269
rect 649 235 655 269
rect 609 197 655 235
rect 609 163 615 197
rect 649 163 655 197
rect 609 125 655 163
rect 609 91 615 125
rect 649 91 655 125
rect 609 53 655 91
rect 609 19 615 53
rect 649 19 655 53
rect 609 -19 655 19
rect 609 -53 615 -19
rect 649 -53 655 -19
rect 609 -91 655 -53
rect 609 -125 615 -91
rect 649 -125 655 -91
rect 609 -163 655 -125
rect 609 -197 615 -163
rect 649 -197 655 -163
rect 609 -235 655 -197
rect 609 -269 615 -235
rect 649 -269 655 -235
rect 609 -307 655 -269
rect 609 -341 615 -307
rect 649 -341 655 -307
rect 609 -379 655 -341
rect 609 -413 615 -379
rect 649 -413 655 -379
rect 609 -451 655 -413
rect 609 -485 615 -451
rect 649 -485 655 -451
rect 609 -500 655 -485
rect 767 485 813 500
rect 767 451 773 485
rect 807 451 813 485
rect 767 413 813 451
rect 767 379 773 413
rect 807 379 813 413
rect 767 341 813 379
rect 767 307 773 341
rect 807 307 813 341
rect 767 269 813 307
rect 767 235 773 269
rect 807 235 813 269
rect 767 197 813 235
rect 767 163 773 197
rect 807 163 813 197
rect 767 125 813 163
rect 767 91 773 125
rect 807 91 813 125
rect 767 53 813 91
rect 767 19 773 53
rect 807 19 813 53
rect 767 -19 813 19
rect 767 -53 773 -19
rect 807 -53 813 -19
rect 767 -91 813 -53
rect 767 -125 773 -91
rect 807 -125 813 -91
rect 767 -163 813 -125
rect 767 -197 773 -163
rect 807 -197 813 -163
rect 767 -235 813 -197
rect 767 -269 773 -235
rect 807 -269 813 -235
rect 767 -307 813 -269
rect 767 -341 773 -307
rect 807 -341 813 -307
rect 767 -379 813 -341
rect 767 -413 773 -379
rect 807 -413 813 -379
rect 767 -451 813 -413
rect 767 -485 773 -451
rect 807 -485 813 -451
rect 767 -500 813 -485
rect 925 485 971 500
rect 925 451 931 485
rect 965 451 971 485
rect 925 413 971 451
rect 925 379 931 413
rect 965 379 971 413
rect 925 341 971 379
rect 925 307 931 341
rect 965 307 971 341
rect 925 269 971 307
rect 925 235 931 269
rect 965 235 971 269
rect 925 197 971 235
rect 925 163 931 197
rect 965 163 971 197
rect 925 125 971 163
rect 925 91 931 125
rect 965 91 971 125
rect 925 53 971 91
rect 925 19 931 53
rect 965 19 971 53
rect 925 -19 971 19
rect 925 -53 931 -19
rect 965 -53 971 -19
rect 925 -91 971 -53
rect 925 -125 931 -91
rect 965 -125 971 -91
rect 925 -163 971 -125
rect 925 -197 931 -163
rect 965 -197 971 -163
rect 925 -235 971 -197
rect 925 -269 931 -235
rect 965 -269 971 -235
rect 925 -307 971 -269
rect 925 -341 931 -307
rect 965 -341 971 -307
rect 925 -379 971 -341
rect 925 -413 931 -379
rect 965 -413 971 -379
rect 925 -451 971 -413
rect 925 -485 931 -451
rect 965 -485 971 -451
rect 925 -500 971 -485
rect 1083 485 1129 500
rect 1083 451 1089 485
rect 1123 451 1129 485
rect 1083 413 1129 451
rect 1083 379 1089 413
rect 1123 379 1129 413
rect 1083 341 1129 379
rect 1083 307 1089 341
rect 1123 307 1129 341
rect 1083 269 1129 307
rect 1083 235 1089 269
rect 1123 235 1129 269
rect 1083 197 1129 235
rect 1083 163 1089 197
rect 1123 163 1129 197
rect 1083 125 1129 163
rect 1083 91 1089 125
rect 1123 91 1129 125
rect 1083 53 1129 91
rect 1083 19 1089 53
rect 1123 19 1129 53
rect 1083 -19 1129 19
rect 1083 -53 1089 -19
rect 1123 -53 1129 -19
rect 1083 -91 1129 -53
rect 1083 -125 1089 -91
rect 1123 -125 1129 -91
rect 1083 -163 1129 -125
rect 1083 -197 1089 -163
rect 1123 -197 1129 -163
rect 1083 -235 1129 -197
rect 1083 -269 1089 -235
rect 1123 -269 1129 -235
rect 1083 -307 1129 -269
rect 1083 -341 1089 -307
rect 1123 -341 1129 -307
rect 1083 -379 1129 -341
rect 1083 -413 1089 -379
rect 1123 -413 1129 -379
rect 1083 -451 1129 -413
rect 1083 -485 1089 -451
rect 1123 -485 1129 -451
rect 1083 -500 1129 -485
rect 1241 485 1287 500
rect 1241 451 1247 485
rect 1281 451 1287 485
rect 1241 413 1287 451
rect 1241 379 1247 413
rect 1281 379 1287 413
rect 1241 341 1287 379
rect 1241 307 1247 341
rect 1281 307 1287 341
rect 1241 269 1287 307
rect 1241 235 1247 269
rect 1281 235 1287 269
rect 1241 197 1287 235
rect 1241 163 1247 197
rect 1281 163 1287 197
rect 1241 125 1287 163
rect 1241 91 1247 125
rect 1281 91 1287 125
rect 1241 53 1287 91
rect 1241 19 1247 53
rect 1281 19 1287 53
rect 1241 -19 1287 19
rect 1241 -53 1247 -19
rect 1281 -53 1287 -19
rect 1241 -91 1287 -53
rect 1241 -125 1247 -91
rect 1281 -125 1287 -91
rect 1241 -163 1287 -125
rect 1241 -197 1247 -163
rect 1281 -197 1287 -163
rect 1241 -235 1287 -197
rect 1241 -269 1247 -235
rect 1281 -269 1287 -235
rect 1241 -307 1287 -269
rect 1241 -341 1247 -307
rect 1281 -341 1287 -307
rect 1241 -379 1287 -341
rect 1241 -413 1247 -379
rect 1281 -413 1287 -379
rect 1241 -451 1287 -413
rect 1241 -485 1247 -451
rect 1281 -485 1287 -451
rect 1241 -500 1287 -485
rect 1399 485 1445 500
rect 1399 451 1405 485
rect 1439 451 1445 485
rect 1399 413 1445 451
rect 1399 379 1405 413
rect 1439 379 1445 413
rect 1399 341 1445 379
rect 1399 307 1405 341
rect 1439 307 1445 341
rect 1399 269 1445 307
rect 1399 235 1405 269
rect 1439 235 1445 269
rect 1399 197 1445 235
rect 1399 163 1405 197
rect 1439 163 1445 197
rect 1399 125 1445 163
rect 1399 91 1405 125
rect 1439 91 1445 125
rect 1399 53 1445 91
rect 1399 19 1405 53
rect 1439 19 1445 53
rect 1399 -19 1445 19
rect 1399 -53 1405 -19
rect 1439 -53 1445 -19
rect 1399 -91 1445 -53
rect 1399 -125 1405 -91
rect 1439 -125 1445 -91
rect 1399 -163 1445 -125
rect 1399 -197 1405 -163
rect 1439 -197 1445 -163
rect 1399 -235 1445 -197
rect 1399 -269 1405 -235
rect 1439 -269 1445 -235
rect 1399 -307 1445 -269
rect 1399 -341 1405 -307
rect 1439 -341 1445 -307
rect 1399 -379 1445 -341
rect 1399 -413 1405 -379
rect 1439 -413 1445 -379
rect 1399 -451 1445 -413
rect 1399 -485 1405 -451
rect 1439 -485 1445 -451
rect 1399 -500 1445 -485
rect 1557 485 1603 500
rect 1557 451 1563 485
rect 1597 451 1603 485
rect 1557 413 1603 451
rect 1557 379 1563 413
rect 1597 379 1603 413
rect 1557 341 1603 379
rect 1557 307 1563 341
rect 1597 307 1603 341
rect 1557 269 1603 307
rect 1557 235 1563 269
rect 1597 235 1603 269
rect 1557 197 1603 235
rect 1557 163 1563 197
rect 1597 163 1603 197
rect 1557 125 1603 163
rect 1557 91 1563 125
rect 1597 91 1603 125
rect 1557 53 1603 91
rect 1557 19 1563 53
rect 1597 19 1603 53
rect 1557 -19 1603 19
rect 1557 -53 1563 -19
rect 1597 -53 1603 -19
rect 1557 -91 1603 -53
rect 1557 -125 1563 -91
rect 1597 -125 1603 -91
rect 1557 -163 1603 -125
rect 1557 -197 1563 -163
rect 1597 -197 1603 -163
rect 1557 -235 1603 -197
rect 1557 -269 1563 -235
rect 1597 -269 1603 -235
rect 1557 -307 1603 -269
rect 1557 -341 1563 -307
rect 1597 -341 1603 -307
rect 1557 -379 1603 -341
rect 1557 -413 1563 -379
rect 1597 -413 1603 -379
rect 1557 -451 1603 -413
rect 1557 -485 1563 -451
rect 1597 -485 1603 -451
rect 1557 -500 1603 -485
<< end >>
