magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< locali >>
rect -43 652 81 686
<< metal1 >>
rect 624 12700 688 12752
rect 1360 12700 1424 12752
rect 49 11955 113 12007
rect 164 11955 228 12007
rect 417 11955 481 12007
rect 785 11955 849 12007
rect 1153 11955 1217 12007
rect 1521 11955 1585 12007
rect 624 11286 688 11338
rect 1360 11286 1424 11338
rect 49 10617 113 10669
rect 164 10617 228 10669
rect 417 10617 481 10669
rect 785 10617 849 10669
rect 1153 10617 1217 10669
rect 1521 10617 1585 10669
rect 624 9872 688 9924
rect 1360 9872 1424 9924
rect 49 9127 113 9179
rect 164 9127 228 9179
rect 417 9127 481 9179
rect 785 9127 849 9179
rect 1153 9127 1217 9179
rect 1521 9127 1585 9179
rect 624 8458 688 8510
rect 1360 8458 1424 8510
rect 49 7789 113 7841
rect 164 7789 228 7841
rect 417 7789 481 7841
rect 785 7789 849 7841
rect 1153 7789 1217 7841
rect 1521 7789 1585 7841
rect 624 7044 688 7096
rect 1360 7044 1424 7096
rect 49 6299 113 6351
rect 164 6299 228 6351
rect 417 6299 481 6351
rect 785 6299 849 6351
rect 1153 6299 1217 6351
rect 1521 6299 1585 6351
rect 624 5630 688 5682
rect 1360 5630 1424 5682
rect 49 4961 113 5013
rect 164 4961 228 5013
rect 417 4961 481 5013
rect 785 4961 849 5013
rect 1153 4961 1217 5013
rect 1521 4961 1585 5013
rect 624 4216 688 4268
rect 1360 4216 1424 4268
rect 49 3471 113 3523
rect 164 3471 228 3523
rect 417 3471 481 3523
rect 785 3471 849 3523
rect 1153 3471 1217 3523
rect 1521 3471 1585 3523
rect 624 2802 688 2854
rect 1360 2802 1424 2854
rect 49 2133 113 2185
rect 164 2133 228 2185
rect 417 2133 481 2185
rect 785 2133 849 2185
rect 1153 2133 1217 2185
rect 1521 2133 1585 2185
rect 624 1388 688 1440
rect 1360 1388 1424 1440
rect -75 643 -11 695
rect 49 643 113 695
rect 164 643 228 695
rect 417 643 481 695
rect 785 643 849 695
rect 1153 643 1217 695
rect 1521 643 1585 695
rect 624 -26 688 26
rect 1360 -26 1424 26
<< metal2 >>
rect 628 12702 684 12750
rect 1364 12702 1420 12750
rect 67 11326 95 11981
rect 168 11957 224 12005
rect 421 11957 477 12005
rect 789 11957 845 12005
rect 1157 11957 1213 12005
rect 1525 11957 1581 12005
rect 67 11298 210 11326
rect 182 10667 210 11298
rect 628 11288 684 11336
rect 1364 11288 1420 11336
rect 67 9912 95 10643
rect 168 10619 224 10667
rect 421 10619 477 10667
rect 789 10619 845 10667
rect 1157 10619 1213 10667
rect 1525 10619 1581 10667
rect 67 9884 210 9912
rect 182 9177 210 9884
rect 628 9874 684 9922
rect 1364 9874 1420 9922
rect 67 8498 95 9153
rect 168 9129 224 9177
rect 421 9129 477 9177
rect 789 9129 845 9177
rect 1157 9129 1213 9177
rect 1525 9129 1581 9177
rect 67 8470 210 8498
rect 182 7839 210 8470
rect 628 8460 684 8508
rect 1364 8460 1420 8508
rect 67 7084 95 7815
rect 168 7791 224 7839
rect 421 7791 477 7839
rect 789 7791 845 7839
rect 1157 7791 1213 7839
rect 1525 7791 1581 7839
rect 67 7056 210 7084
rect 182 6349 210 7056
rect 628 7046 684 7094
rect 1364 7046 1420 7094
rect 67 5670 95 6325
rect 168 6301 224 6349
rect 421 6301 477 6349
rect 789 6301 845 6349
rect 1157 6301 1213 6349
rect 1525 6301 1581 6349
rect 67 5642 210 5670
rect 182 5011 210 5642
rect 628 5632 684 5680
rect 1364 5632 1420 5680
rect 67 4256 95 4987
rect 168 4963 224 5011
rect 421 4963 477 5011
rect 789 4963 845 5011
rect 1157 4963 1213 5011
rect 1525 4963 1581 5011
rect 67 4228 210 4256
rect 182 3521 210 4228
rect 628 4218 684 4266
rect 1364 4218 1420 4266
rect 67 2842 95 3497
rect 168 3473 224 3521
rect 421 3473 477 3521
rect 789 3473 845 3521
rect 1157 3473 1213 3521
rect 1525 3473 1581 3521
rect 67 2814 210 2842
rect 182 2183 210 2814
rect 628 2804 684 2852
rect 1364 2804 1420 2852
rect 67 1428 95 2159
rect 168 2135 224 2183
rect 421 2135 477 2183
rect 789 2135 845 2183
rect 1157 2135 1213 2183
rect 1525 2135 1581 2183
rect 67 1400 210 1428
rect 182 693 210 1400
rect 628 1390 684 1438
rect 1364 1390 1420 1438
rect -57 655 -29 683
rect 168 645 224 693
rect 421 645 477 693
rect 789 645 845 693
rect 1157 645 1213 693
rect 1525 645 1581 693
rect 628 -24 684 24
rect 1364 -24 1420 24
<< metal3 >>
rect 607 12677 705 12775
rect 1343 12677 1441 12775
rect 196 11951 1553 12011
rect 607 11263 705 11361
rect 1343 11263 1441 11361
rect 196 10613 1553 10673
rect 607 9849 705 9947
rect 1343 9849 1441 9947
rect 196 9123 1553 9183
rect 607 8435 705 8533
rect 1343 8435 1441 8533
rect 196 7785 1553 7845
rect 607 7021 705 7119
rect 1343 7021 1441 7119
rect 196 6295 1553 6355
rect 607 5607 705 5705
rect 1343 5607 1441 5705
rect 196 4957 1553 5017
rect 607 4193 705 4291
rect 1343 4193 1441 4291
rect 196 3467 1553 3527
rect 607 2779 705 2877
rect 1343 2779 1441 2877
rect 196 2129 1553 2189
rect 607 1365 705 1463
rect 1343 1365 1441 1463
rect 196 639 1553 699
rect 607 -49 705 49
rect 1343 -49 1441 49
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 -75 0 1 637
box 0 0 64 64
use contact_7  contact_7_1
timestamp 1624494425
transform 1 0 -72 0 1 636
box 0 0 58 66
use contact_9  contact_9_76
timestamp 1624494425
transform 1 0 163 0 1 632
box 0 0 66 74
use contact_8  contact_8_85
timestamp 1624494425
transform 1 0 164 0 1 637
box 0 0 64 64
use contact_7  contact_7_86
timestamp 1624494425
transform 1 0 167 0 1 636
box 0 0 58 66
use contact_8  contact_8_86
timestamp 1624494425
transform 1 0 49 0 1 637
box 0 0 64 64
use contact_7  contact_7_87
timestamp 1624494425
transform 1 0 52 0 1 636
box 0 0 58 66
use pinv_19  pinv_19_44
timestamp 1624494425
transform 1 0 0 0 1 0
box -36 -17 404 1471
use pinv_19  pinv_19_43
timestamp 1624494425
transform 1 0 368 0 1 0
box -36 -17 404 1471
use pinv_19  pinv_19_39
timestamp 1624494425
transform 1 0 0 0 -1 2828
box -36 -17 404 1471
use pinv_19  pinv_19_38
timestamp 1624494425
transform 1 0 368 0 -1 2828
box -36 -17 404 1471
use contact_9  contact_9_33
timestamp 1624494425
transform 1 0 623 0 1 -37
box 0 0 66 74
use contact_8  contact_8_34
timestamp 1624494425
transform 1 0 624 0 1 -32
box 0 0 64 64
use contact_7  contact_7_35
timestamp 1624494425
transform 1 0 627 0 1 -33
box 0 0 58 66
use contact_9  contact_9_79
timestamp 1624494425
transform 1 0 784 0 1 632
box 0 0 66 74
use contact_8  contact_8_89
timestamp 1624494425
transform 1 0 785 0 1 637
box 0 0 64 64
use contact_7  contact_7_90
timestamp 1624494425
transform 1 0 788 0 1 636
box 0 0 58 66
use contact_9  contact_9_80
timestamp 1624494425
transform 1 0 416 0 1 632
box 0 0 66 74
use contact_8  contact_8_90
timestamp 1624494425
transform 1 0 417 0 1 637
box 0 0 64 64
use contact_7  contact_7_91
timestamp 1624494425
transform 1 0 420 0 1 636
box 0 0 58 66
use contact_9  contact_9_31
timestamp 1624494425
transform 1 0 623 0 1 1377
box 0 0 66 74
use contact_8  contact_8_32
timestamp 1624494425
transform 1 0 624 0 1 1382
box 0 0 64 64
use contact_7  contact_7_33
timestamp 1624494425
transform 1 0 627 0 1 1381
box 0 0 58 66
use contact_9  contact_9_35
timestamp 1624494425
transform 1 0 623 0 1 1377
box 0 0 66 74
use contact_8  contact_8_36
timestamp 1624494425
transform 1 0 624 0 1 1382
box 0 0 64 64
use contact_7  contact_7_37
timestamp 1624494425
transform 1 0 627 0 1 1381
box 0 0 58 66
use pinv_19  pinv_19_42
timestamp 1624494425
transform 1 0 736 0 1 0
box -36 -17 404 1471
use pinv_19  pinv_19_37
timestamp 1624494425
transform 1 0 736 0 -1 2828
box -36 -17 404 1471
use contact_7  contact_7_89
timestamp 1624494425
transform 1 0 1156 0 1 636
box 0 0 58 66
use contact_8  contact_8_88
timestamp 1624494425
transform 1 0 1153 0 1 637
box 0 0 64 64
use contact_9  contact_9_78
timestamp 1624494425
transform 1 0 1152 0 1 632
box 0 0 66 74
use pinv_19  pinv_19_36
timestamp 1624494425
transform 1 0 1104 0 -1 2828
box -36 -17 404 1471
use pinv_19  pinv_19_41
timestamp 1624494425
transform 1 0 1104 0 1 0
box -36 -17 404 1471
use contact_9  contact_9_32
timestamp 1624494425
transform 1 0 1359 0 1 -37
box 0 0 66 74
use contact_8  contact_8_33
timestamp 1624494425
transform 1 0 1360 0 1 -32
box 0 0 64 64
use contact_7  contact_7_34
timestamp 1624494425
transform 1 0 1363 0 1 -33
box 0 0 58 66
use contact_9  contact_9_77
timestamp 1624494425
transform 1 0 1520 0 1 632
box 0 0 66 74
use contact_8  contact_8_87
timestamp 1624494425
transform 1 0 1521 0 1 637
box 0 0 64 64
use contact_7  contact_7_88
timestamp 1624494425
transform 1 0 1524 0 1 636
box 0 0 58 66
use contact_9  contact_9_30
timestamp 1624494425
transform 1 0 1359 0 1 1377
box 0 0 66 74
use contact_8  contact_8_31
timestamp 1624494425
transform 1 0 1360 0 1 1382
box 0 0 64 64
use contact_7  contact_7_32
timestamp 1624494425
transform 1 0 1363 0 1 1381
box 0 0 58 66
use contact_9  contact_9_34
timestamp 1624494425
transform 1 0 1359 0 1 1377
box 0 0 66 74
use contact_8  contact_8_35
timestamp 1624494425
transform 1 0 1360 0 1 1382
box 0 0 64 64
use contact_7  contact_7_36
timestamp 1624494425
transform 1 0 1363 0 1 1381
box 0 0 58 66
use pinv_19  pinv_19_40
timestamp 1624494425
transform 1 0 1472 0 1 0
box -36 -17 404 1471
use pinv_19  pinv_19_35
timestamp 1624494425
transform 1 0 1472 0 -1 2828
box -36 -17 404 1471
use contact_7  contact_7_81
timestamp 1624494425
transform 1 0 52 0 1 2126
box 0 0 58 66
use contact_8  contact_8_80
timestamp 1624494425
transform 1 0 49 0 1 2127
box 0 0 64 64
use contact_7  contact_7_80
timestamp 1624494425
transform 1 0 167 0 1 2126
box 0 0 58 66
use contact_8  contact_8_79
timestamp 1624494425
transform 1 0 164 0 1 2127
box 0 0 64 64
use contact_9  contact_9_71
timestamp 1624494425
transform 1 0 163 0 1 2122
box 0 0 66 74
use pinv_19  pinv_19_33
timestamp 1624494425
transform 1 0 368 0 1 2828
box -36 -17 404 1471
use pinv_19  pinv_19_34
timestamp 1624494425
transform 1 0 0 0 1 2828
box -36 -17 404 1471
use contact_9  contact_9_74
timestamp 1624494425
transform 1 0 784 0 1 2122
box 0 0 66 74
use contact_8  contact_8_83
timestamp 1624494425
transform 1 0 785 0 1 2127
box 0 0 64 64
use contact_7  contact_7_84
timestamp 1624494425
transform 1 0 788 0 1 2126
box 0 0 58 66
use contact_9  contact_9_75
timestamp 1624494425
transform 1 0 416 0 1 2122
box 0 0 66 74
use contact_8  contact_8_84
timestamp 1624494425
transform 1 0 417 0 1 2127
box 0 0 64 64
use contact_7  contact_7_85
timestamp 1624494425
transform 1 0 420 0 1 2126
box 0 0 58 66
use contact_9  contact_9_25
timestamp 1624494425
transform 1 0 623 0 1 2791
box 0 0 66 74
use contact_8  contact_8_26
timestamp 1624494425
transform 1 0 624 0 1 2796
box 0 0 64 64
use contact_7  contact_7_27
timestamp 1624494425
transform 1 0 627 0 1 2795
box 0 0 58 66
use contact_9  contact_9_29
timestamp 1624494425
transform 1 0 623 0 1 2791
box 0 0 66 74
use contact_8  contact_8_30
timestamp 1624494425
transform 1 0 624 0 1 2796
box 0 0 64 64
use contact_7  contact_7_31
timestamp 1624494425
transform 1 0 627 0 1 2795
box 0 0 58 66
use pinv_19  pinv_19_32
timestamp 1624494425
transform 1 0 736 0 1 2828
box -36 -17 404 1471
use contact_7  contact_7_83
timestamp 1624494425
transform 1 0 1156 0 1 2126
box 0 0 58 66
use contact_8  contact_8_82
timestamp 1624494425
transform 1 0 1153 0 1 2127
box 0 0 64 64
use contact_9  contact_9_73
timestamp 1624494425
transform 1 0 1152 0 1 2122
box 0 0 66 74
use pinv_19  pinv_19_31
timestamp 1624494425
transform 1 0 1104 0 1 2828
box -36 -17 404 1471
use contact_9  contact_9_72
timestamp 1624494425
transform 1 0 1520 0 1 2122
box 0 0 66 74
use contact_8  contact_8_81
timestamp 1624494425
transform 1 0 1521 0 1 2127
box 0 0 64 64
use contact_7  contact_7_82
timestamp 1624494425
transform 1 0 1524 0 1 2126
box 0 0 58 66
use contact_9  contact_9_24
timestamp 1624494425
transform 1 0 1359 0 1 2791
box 0 0 66 74
use contact_8  contact_8_25
timestamp 1624494425
transform 1 0 1360 0 1 2796
box 0 0 64 64
use contact_7  contact_7_26
timestamp 1624494425
transform 1 0 1363 0 1 2795
box 0 0 58 66
use contact_9  contact_9_28
timestamp 1624494425
transform 1 0 1359 0 1 2791
box 0 0 66 74
use contact_8  contact_8_29
timestamp 1624494425
transform 1 0 1360 0 1 2796
box 0 0 64 64
use contact_7  contact_7_30
timestamp 1624494425
transform 1 0 1363 0 1 2795
box 0 0 58 66
use pinv_19  pinv_19_30
timestamp 1624494425
transform 1 0 1472 0 1 2828
box -36 -17 404 1471
use contact_7  contact_7_75
timestamp 1624494425
transform 1 0 52 0 1 3464
box 0 0 58 66
use contact_8  contact_8_74
timestamp 1624494425
transform 1 0 49 0 1 3465
box 0 0 64 64
use contact_7  contact_7_74
timestamp 1624494425
transform 1 0 167 0 1 3464
box 0 0 58 66
use contact_8  contact_8_73
timestamp 1624494425
transform 1 0 164 0 1 3465
box 0 0 64 64
use contact_9  contact_9_66
timestamp 1624494425
transform 1 0 163 0 1 3460
box 0 0 66 74
use pinv_19  pinv_19_28
timestamp 1624494425
transform 1 0 368 0 -1 5656
box -36 -17 404 1471
use pinv_19  pinv_19_29
timestamp 1624494425
transform 1 0 0 0 -1 5656
box -36 -17 404 1471
use contact_9  contact_9_69
timestamp 1624494425
transform 1 0 784 0 1 3460
box 0 0 66 74
use contact_8  contact_8_77
timestamp 1624494425
transform 1 0 785 0 1 3465
box 0 0 64 64
use contact_7  contact_7_78
timestamp 1624494425
transform 1 0 788 0 1 3464
box 0 0 58 66
use contact_9  contact_9_70
timestamp 1624494425
transform 1 0 416 0 1 3460
box 0 0 66 74
use contact_8  contact_8_78
timestamp 1624494425
transform 1 0 417 0 1 3465
box 0 0 64 64
use contact_7  contact_7_79
timestamp 1624494425
transform 1 0 420 0 1 3464
box 0 0 58 66
use contact_9  contact_9_23
timestamp 1624494425
transform 1 0 623 0 1 4205
box 0 0 66 74
use contact_8  contact_8_24
timestamp 1624494425
transform 1 0 624 0 1 4210
box 0 0 64 64
use contact_7  contact_7_25
timestamp 1624494425
transform 1 0 627 0 1 4209
box 0 0 58 66
use contact_9  contact_9_27
timestamp 1624494425
transform 1 0 623 0 1 4205
box 0 0 66 74
use contact_8  contact_8_28
timestamp 1624494425
transform 1 0 624 0 1 4210
box 0 0 64 64
use contact_7  contact_7_29
timestamp 1624494425
transform 1 0 627 0 1 4209
box 0 0 58 66
use pinv_19  pinv_19_27
timestamp 1624494425
transform 1 0 736 0 -1 5656
box -36 -17 404 1471
use contact_7  contact_7_77
timestamp 1624494425
transform 1 0 1156 0 1 3464
box 0 0 58 66
use contact_8  contact_8_76
timestamp 1624494425
transform 1 0 1153 0 1 3465
box 0 0 64 64
use contact_9  contact_9_68
timestamp 1624494425
transform 1 0 1152 0 1 3460
box 0 0 66 74
use pinv_19  pinv_19_26
timestamp 1624494425
transform 1 0 1104 0 -1 5656
box -36 -17 404 1471
use contact_9  contact_9_67
timestamp 1624494425
transform 1 0 1520 0 1 3460
box 0 0 66 74
use contact_8  contact_8_75
timestamp 1624494425
transform 1 0 1521 0 1 3465
box 0 0 64 64
use contact_7  contact_7_76
timestamp 1624494425
transform 1 0 1524 0 1 3464
box 0 0 58 66
use contact_9  contact_9_22
timestamp 1624494425
transform 1 0 1359 0 1 4205
box 0 0 66 74
use contact_8  contact_8_23
timestamp 1624494425
transform 1 0 1360 0 1 4210
box 0 0 64 64
use contact_7  contact_7_24
timestamp 1624494425
transform 1 0 1363 0 1 4209
box 0 0 58 66
use contact_9  contact_9_26
timestamp 1624494425
transform 1 0 1359 0 1 4205
box 0 0 66 74
use contact_8  contact_8_27
timestamp 1624494425
transform 1 0 1360 0 1 4210
box 0 0 64 64
use contact_7  contact_7_28
timestamp 1624494425
transform 1 0 1363 0 1 4209
box 0 0 58 66
use pinv_19  pinv_19_25
timestamp 1624494425
transform 1 0 1472 0 -1 5656
box -36 -17 404 1471
use contact_7  contact_7_69
timestamp 1624494425
transform 1 0 52 0 1 4954
box 0 0 58 66
use contact_8  contact_8_68
timestamp 1624494425
transform 1 0 49 0 1 4955
box 0 0 64 64
use contact_7  contact_7_68
timestamp 1624494425
transform 1 0 167 0 1 4954
box 0 0 58 66
use contact_8  contact_8_67
timestamp 1624494425
transform 1 0 164 0 1 4955
box 0 0 64 64
use contact_9  contact_9_61
timestamp 1624494425
transform 1 0 163 0 1 4950
box 0 0 66 74
use pinv_19  pinv_19_23
timestamp 1624494425
transform 1 0 368 0 1 5656
box -36 -17 404 1471
use pinv_19  pinv_19_24
timestamp 1624494425
transform 1 0 0 0 1 5656
box -36 -17 404 1471
use contact_9  contact_9_64
timestamp 1624494425
transform 1 0 784 0 1 4950
box 0 0 66 74
use contact_8  contact_8_71
timestamp 1624494425
transform 1 0 785 0 1 4955
box 0 0 64 64
use contact_7  contact_7_72
timestamp 1624494425
transform 1 0 788 0 1 4954
box 0 0 58 66
use contact_9  contact_9_65
timestamp 1624494425
transform 1 0 416 0 1 4950
box 0 0 66 74
use contact_8  contact_8_72
timestamp 1624494425
transform 1 0 417 0 1 4955
box 0 0 64 64
use contact_7  contact_7_73
timestamp 1624494425
transform 1 0 420 0 1 4954
box 0 0 58 66
use contact_9  contact_9_17
timestamp 1624494425
transform 1 0 623 0 1 5619
box 0 0 66 74
use contact_8  contact_8_18
timestamp 1624494425
transform 1 0 624 0 1 5624
box 0 0 64 64
use contact_7  contact_7_19
timestamp 1624494425
transform 1 0 627 0 1 5623
box 0 0 58 66
use contact_9  contact_9_21
timestamp 1624494425
transform 1 0 623 0 1 5619
box 0 0 66 74
use contact_8  contact_8_22
timestamp 1624494425
transform 1 0 624 0 1 5624
box 0 0 64 64
use contact_7  contact_7_23
timestamp 1624494425
transform 1 0 627 0 1 5623
box 0 0 58 66
use pinv_19  pinv_19_22
timestamp 1624494425
transform 1 0 736 0 1 5656
box -36 -17 404 1471
use contact_7  contact_7_71
timestamp 1624494425
transform 1 0 1156 0 1 4954
box 0 0 58 66
use contact_8  contact_8_70
timestamp 1624494425
transform 1 0 1153 0 1 4955
box 0 0 64 64
use contact_9  contact_9_63
timestamp 1624494425
transform 1 0 1152 0 1 4950
box 0 0 66 74
use pinv_19  pinv_19_21
timestamp 1624494425
transform 1 0 1104 0 1 5656
box -36 -17 404 1471
use contact_9  contact_9_62
timestamp 1624494425
transform 1 0 1520 0 1 4950
box 0 0 66 74
use contact_8  contact_8_69
timestamp 1624494425
transform 1 0 1521 0 1 4955
box 0 0 64 64
use contact_7  contact_7_70
timestamp 1624494425
transform 1 0 1524 0 1 4954
box 0 0 58 66
use contact_9  contact_9_16
timestamp 1624494425
transform 1 0 1359 0 1 5619
box 0 0 66 74
use contact_8  contact_8_17
timestamp 1624494425
transform 1 0 1360 0 1 5624
box 0 0 64 64
use contact_7  contact_7_18
timestamp 1624494425
transform 1 0 1363 0 1 5623
box 0 0 58 66
use contact_9  contact_9_20
timestamp 1624494425
transform 1 0 1359 0 1 5619
box 0 0 66 74
use contact_8  contact_8_21
timestamp 1624494425
transform 1 0 1360 0 1 5624
box 0 0 64 64
use contact_7  contact_7_22
timestamp 1624494425
transform 1 0 1363 0 1 5623
box 0 0 58 66
use pinv_19  pinv_19_20
timestamp 1624494425
transform 1 0 1472 0 1 5656
box -36 -17 404 1471
use contact_7  contact_7_63
timestamp 1624494425
transform 1 0 52 0 1 6292
box 0 0 58 66
use contact_8  contact_8_62
timestamp 1624494425
transform 1 0 49 0 1 6293
box 0 0 64 64
use contact_7  contact_7_62
timestamp 1624494425
transform 1 0 167 0 1 6292
box 0 0 58 66
use contact_8  contact_8_61
timestamp 1624494425
transform 1 0 164 0 1 6293
box 0 0 64 64
use contact_9  contact_9_56
timestamp 1624494425
transform 1 0 163 0 1 6288
box 0 0 66 74
use pinv_19  pinv_19_18
timestamp 1624494425
transform 1 0 368 0 -1 8484
box -36 -17 404 1471
use pinv_19  pinv_19_19
timestamp 1624494425
transform 1 0 0 0 -1 8484
box -36 -17 404 1471
use contact_9  contact_9_59
timestamp 1624494425
transform 1 0 784 0 1 6288
box 0 0 66 74
use contact_8  contact_8_65
timestamp 1624494425
transform 1 0 785 0 1 6293
box 0 0 64 64
use contact_7  contact_7_66
timestamp 1624494425
transform 1 0 788 0 1 6292
box 0 0 58 66
use contact_9  contact_9_60
timestamp 1624494425
transform 1 0 416 0 1 6288
box 0 0 66 74
use contact_8  contact_8_66
timestamp 1624494425
transform 1 0 417 0 1 6293
box 0 0 64 64
use contact_7  contact_7_67
timestamp 1624494425
transform 1 0 420 0 1 6292
box 0 0 58 66
use contact_9  contact_9_15
timestamp 1624494425
transform 1 0 623 0 1 7033
box 0 0 66 74
use contact_8  contact_8_16
timestamp 1624494425
transform 1 0 624 0 1 7038
box 0 0 64 64
use contact_7  contact_7_17
timestamp 1624494425
transform 1 0 627 0 1 7037
box 0 0 58 66
use contact_9  contact_9_19
timestamp 1624494425
transform 1 0 623 0 1 7033
box 0 0 66 74
use contact_8  contact_8_20
timestamp 1624494425
transform 1 0 624 0 1 7038
box 0 0 64 64
use contact_7  contact_7_21
timestamp 1624494425
transform 1 0 627 0 1 7037
box 0 0 58 66
use pinv_19  pinv_19_17
timestamp 1624494425
transform 1 0 736 0 -1 8484
box -36 -17 404 1471
use contact_7  contact_7_65
timestamp 1624494425
transform 1 0 1156 0 1 6292
box 0 0 58 66
use contact_8  contact_8_64
timestamp 1624494425
transform 1 0 1153 0 1 6293
box 0 0 64 64
use contact_9  contact_9_58
timestamp 1624494425
transform 1 0 1152 0 1 6288
box 0 0 66 74
use pinv_19  pinv_19_16
timestamp 1624494425
transform 1 0 1104 0 -1 8484
box -36 -17 404 1471
use contact_9  contact_9_57
timestamp 1624494425
transform 1 0 1520 0 1 6288
box 0 0 66 74
use contact_8  contact_8_63
timestamp 1624494425
transform 1 0 1521 0 1 6293
box 0 0 64 64
use contact_7  contact_7_64
timestamp 1624494425
transform 1 0 1524 0 1 6292
box 0 0 58 66
use contact_9  contact_9_14
timestamp 1624494425
transform 1 0 1359 0 1 7033
box 0 0 66 74
use contact_8  contact_8_15
timestamp 1624494425
transform 1 0 1360 0 1 7038
box 0 0 64 64
use contact_7  contact_7_16
timestamp 1624494425
transform 1 0 1363 0 1 7037
box 0 0 58 66
use contact_9  contact_9_18
timestamp 1624494425
transform 1 0 1359 0 1 7033
box 0 0 66 74
use contact_8  contact_8_19
timestamp 1624494425
transform 1 0 1360 0 1 7038
box 0 0 64 64
use contact_7  contact_7_20
timestamp 1624494425
transform 1 0 1363 0 1 7037
box 0 0 58 66
use pinv_19  pinv_19_15
timestamp 1624494425
transform 1 0 1472 0 -1 8484
box -36 -17 404 1471
use contact_7  contact_7_57
timestamp 1624494425
transform 1 0 52 0 1 7782
box 0 0 58 66
use contact_8  contact_8_56
timestamp 1624494425
transform 1 0 49 0 1 7783
box 0 0 64 64
use contact_7  contact_7_56
timestamp 1624494425
transform 1 0 167 0 1 7782
box 0 0 58 66
use contact_8  contact_8_55
timestamp 1624494425
transform 1 0 164 0 1 7783
box 0 0 64 64
use contact_9  contact_9_51
timestamp 1624494425
transform 1 0 163 0 1 7778
box 0 0 66 74
use pinv_19  pinv_19_13
timestamp 1624494425
transform 1 0 368 0 1 8484
box -36 -17 404 1471
use pinv_19  pinv_19_14
timestamp 1624494425
transform 1 0 0 0 1 8484
box -36 -17 404 1471
use contact_9  contact_9_54
timestamp 1624494425
transform 1 0 784 0 1 7778
box 0 0 66 74
use contact_8  contact_8_59
timestamp 1624494425
transform 1 0 785 0 1 7783
box 0 0 64 64
use contact_7  contact_7_60
timestamp 1624494425
transform 1 0 788 0 1 7782
box 0 0 58 66
use contact_9  contact_9_55
timestamp 1624494425
transform 1 0 416 0 1 7778
box 0 0 66 74
use contact_8  contact_8_60
timestamp 1624494425
transform 1 0 417 0 1 7783
box 0 0 64 64
use contact_7  contact_7_61
timestamp 1624494425
transform 1 0 420 0 1 7782
box 0 0 58 66
use contact_9  contact_9_9
timestamp 1624494425
transform 1 0 623 0 1 8447
box 0 0 66 74
use contact_8  contact_8_10
timestamp 1624494425
transform 1 0 624 0 1 8452
box 0 0 64 64
use contact_7  contact_7_11
timestamp 1624494425
transform 1 0 627 0 1 8451
box 0 0 58 66
use contact_9  contact_9_13
timestamp 1624494425
transform 1 0 623 0 1 8447
box 0 0 66 74
use contact_8  contact_8_14
timestamp 1624494425
transform 1 0 624 0 1 8452
box 0 0 64 64
use contact_7  contact_7_15
timestamp 1624494425
transform 1 0 627 0 1 8451
box 0 0 58 66
use pinv_19  pinv_19_12
timestamp 1624494425
transform 1 0 736 0 1 8484
box -36 -17 404 1471
use contact_7  contact_7_59
timestamp 1624494425
transform 1 0 1156 0 1 7782
box 0 0 58 66
use contact_8  contact_8_58
timestamp 1624494425
transform 1 0 1153 0 1 7783
box 0 0 64 64
use contact_9  contact_9_53
timestamp 1624494425
transform 1 0 1152 0 1 7778
box 0 0 66 74
use pinv_19  pinv_19_11
timestamp 1624494425
transform 1 0 1104 0 1 8484
box -36 -17 404 1471
use contact_9  contact_9_52
timestamp 1624494425
transform 1 0 1520 0 1 7778
box 0 0 66 74
use contact_8  contact_8_57
timestamp 1624494425
transform 1 0 1521 0 1 7783
box 0 0 64 64
use contact_7  contact_7_58
timestamp 1624494425
transform 1 0 1524 0 1 7782
box 0 0 58 66
use contact_9  contact_9_8
timestamp 1624494425
transform 1 0 1359 0 1 8447
box 0 0 66 74
use contact_8  contact_8_9
timestamp 1624494425
transform 1 0 1360 0 1 8452
box 0 0 64 64
use contact_7  contact_7_10
timestamp 1624494425
transform 1 0 1363 0 1 8451
box 0 0 58 66
use contact_9  contact_9_12
timestamp 1624494425
transform 1 0 1359 0 1 8447
box 0 0 66 74
use contact_8  contact_8_13
timestamp 1624494425
transform 1 0 1360 0 1 8452
box 0 0 64 64
use contact_7  contact_7_14
timestamp 1624494425
transform 1 0 1363 0 1 8451
box 0 0 58 66
use pinv_19  pinv_19_10
timestamp 1624494425
transform 1 0 1472 0 1 8484
box -36 -17 404 1471
use contact_7  contact_7_51
timestamp 1624494425
transform 1 0 52 0 1 9120
box 0 0 58 66
use contact_8  contact_8_50
timestamp 1624494425
transform 1 0 49 0 1 9121
box 0 0 64 64
use contact_7  contact_7_50
timestamp 1624494425
transform 1 0 167 0 1 9120
box 0 0 58 66
use contact_8  contact_8_49
timestamp 1624494425
transform 1 0 164 0 1 9121
box 0 0 64 64
use contact_9  contact_9_46
timestamp 1624494425
transform 1 0 163 0 1 9116
box 0 0 66 74
use pinv_19  pinv_19_8
timestamp 1624494425
transform 1 0 368 0 -1 11312
box -36 -17 404 1471
use pinv_19  pinv_19_9
timestamp 1624494425
transform 1 0 0 0 -1 11312
box -36 -17 404 1471
use contact_9  contact_9_49
timestamp 1624494425
transform 1 0 784 0 1 9116
box 0 0 66 74
use contact_8  contact_8_53
timestamp 1624494425
transform 1 0 785 0 1 9121
box 0 0 64 64
use contact_7  contact_7_54
timestamp 1624494425
transform 1 0 788 0 1 9120
box 0 0 58 66
use contact_9  contact_9_50
timestamp 1624494425
transform 1 0 416 0 1 9116
box 0 0 66 74
use contact_8  contact_8_54
timestamp 1624494425
transform 1 0 417 0 1 9121
box 0 0 64 64
use contact_7  contact_7_55
timestamp 1624494425
transform 1 0 420 0 1 9120
box 0 0 58 66
use contact_9  contact_9_7
timestamp 1624494425
transform 1 0 623 0 1 9861
box 0 0 66 74
use contact_8  contact_8_8
timestamp 1624494425
transform 1 0 624 0 1 9866
box 0 0 64 64
use contact_7  contact_7_9
timestamp 1624494425
transform 1 0 627 0 1 9865
box 0 0 58 66
use contact_9  contact_9_11
timestamp 1624494425
transform 1 0 623 0 1 9861
box 0 0 66 74
use contact_8  contact_8_12
timestamp 1624494425
transform 1 0 624 0 1 9866
box 0 0 64 64
use contact_7  contact_7_13
timestamp 1624494425
transform 1 0 627 0 1 9865
box 0 0 58 66
use pinv_19  pinv_19_7
timestamp 1624494425
transform 1 0 736 0 -1 11312
box -36 -17 404 1471
use contact_7  contact_7_53
timestamp 1624494425
transform 1 0 1156 0 1 9120
box 0 0 58 66
use contact_8  contact_8_52
timestamp 1624494425
transform 1 0 1153 0 1 9121
box 0 0 64 64
use contact_9  contact_9_48
timestamp 1624494425
transform 1 0 1152 0 1 9116
box 0 0 66 74
use pinv_19  pinv_19_6
timestamp 1624494425
transform 1 0 1104 0 -1 11312
box -36 -17 404 1471
use contact_9  contact_9_47
timestamp 1624494425
transform 1 0 1520 0 1 9116
box 0 0 66 74
use contact_8  contact_8_51
timestamp 1624494425
transform 1 0 1521 0 1 9121
box 0 0 64 64
use contact_7  contact_7_52
timestamp 1624494425
transform 1 0 1524 0 1 9120
box 0 0 58 66
use contact_9  contact_9_6
timestamp 1624494425
transform 1 0 1359 0 1 9861
box 0 0 66 74
use contact_8  contact_8_7
timestamp 1624494425
transform 1 0 1360 0 1 9866
box 0 0 64 64
use contact_7  contact_7_8
timestamp 1624494425
transform 1 0 1363 0 1 9865
box 0 0 58 66
use contact_9  contact_9_10
timestamp 1624494425
transform 1 0 1359 0 1 9861
box 0 0 66 74
use contact_8  contact_8_11
timestamp 1624494425
transform 1 0 1360 0 1 9866
box 0 0 64 64
use contact_7  contact_7_12
timestamp 1624494425
transform 1 0 1363 0 1 9865
box 0 0 58 66
use pinv_19  pinv_19_5
timestamp 1624494425
transform 1 0 1472 0 -1 11312
box -36 -17 404 1471
use contact_7  contact_7_45
timestamp 1624494425
transform 1 0 52 0 1 10610
box 0 0 58 66
use contact_8  contact_8_44
timestamp 1624494425
transform 1 0 49 0 1 10611
box 0 0 64 64
use contact_7  contact_7_44
timestamp 1624494425
transform 1 0 167 0 1 10610
box 0 0 58 66
use contact_8  contact_8_43
timestamp 1624494425
transform 1 0 164 0 1 10611
box 0 0 64 64
use contact_9  contact_9_41
timestamp 1624494425
transform 1 0 163 0 1 10606
box 0 0 66 74
use pinv_19  pinv_19_3
timestamp 1624494425
transform 1 0 368 0 1 11312
box -36 -17 404 1471
use pinv_19  pinv_19_4
timestamp 1624494425
transform 1 0 0 0 1 11312
box -36 -17 404 1471
use contact_9  contact_9_44
timestamp 1624494425
transform 1 0 784 0 1 10606
box 0 0 66 74
use contact_8  contact_8_47
timestamp 1624494425
transform 1 0 785 0 1 10611
box 0 0 64 64
use contact_7  contact_7_48
timestamp 1624494425
transform 1 0 788 0 1 10610
box 0 0 58 66
use contact_9  contact_9_45
timestamp 1624494425
transform 1 0 416 0 1 10606
box 0 0 66 74
use contact_8  contact_8_48
timestamp 1624494425
transform 1 0 417 0 1 10611
box 0 0 64 64
use contact_7  contact_7_49
timestamp 1624494425
transform 1 0 420 0 1 10610
box 0 0 58 66
use contact_9  contact_9_1
timestamp 1624494425
transform 1 0 623 0 1 11275
box 0 0 66 74
use contact_8  contact_8_2
timestamp 1624494425
transform 1 0 624 0 1 11280
box 0 0 64 64
use contact_7  contact_7_3
timestamp 1624494425
transform 1 0 627 0 1 11279
box 0 0 58 66
use contact_9  contact_9_5
timestamp 1624494425
transform 1 0 623 0 1 11275
box 0 0 66 74
use contact_8  contact_8_6
timestamp 1624494425
transform 1 0 624 0 1 11280
box 0 0 64 64
use contact_7  contact_7_7
timestamp 1624494425
transform 1 0 627 0 1 11279
box 0 0 58 66
use pinv_19  pinv_19_2
timestamp 1624494425
transform 1 0 736 0 1 11312
box -36 -17 404 1471
use contact_7  contact_7_47
timestamp 1624494425
transform 1 0 1156 0 1 10610
box 0 0 58 66
use contact_8  contact_8_46
timestamp 1624494425
transform 1 0 1153 0 1 10611
box 0 0 64 64
use contact_9  contact_9_43
timestamp 1624494425
transform 1 0 1152 0 1 10606
box 0 0 66 74
use pinv_19  pinv_19_1
timestamp 1624494425
transform 1 0 1104 0 1 11312
box -36 -17 404 1471
use contact_9  contact_9_42
timestamp 1624494425
transform 1 0 1520 0 1 10606
box 0 0 66 74
use contact_8  contact_8_45
timestamp 1624494425
transform 1 0 1521 0 1 10611
box 0 0 64 64
use contact_7  contact_7_46
timestamp 1624494425
transform 1 0 1524 0 1 10610
box 0 0 58 66
use contact_9  contact_9_0
timestamp 1624494425
transform 1 0 1359 0 1 11275
box 0 0 66 74
use contact_8  contact_8_1
timestamp 1624494425
transform 1 0 1360 0 1 11280
box 0 0 64 64
use contact_7  contact_7_2
timestamp 1624494425
transform 1 0 1363 0 1 11279
box 0 0 58 66
use contact_9  contact_9_4
timestamp 1624494425
transform 1 0 1359 0 1 11275
box 0 0 66 74
use contact_8  contact_8_5
timestamp 1624494425
transform 1 0 1360 0 1 11280
box 0 0 64 64
use contact_7  contact_7_6
timestamp 1624494425
transform 1 0 1363 0 1 11279
box 0 0 58 66
use pinv_19  pinv_19_0
timestamp 1624494425
transform 1 0 1472 0 1 11312
box -36 -17 404 1471
use contact_7  contact_7_39
timestamp 1624494425
transform 1 0 52 0 1 11948
box 0 0 58 66
use contact_8  contact_8_38
timestamp 1624494425
transform 1 0 49 0 1 11949
box 0 0 64 64
use contact_7  contact_7_38
timestamp 1624494425
transform 1 0 167 0 1 11948
box 0 0 58 66
use contact_8  contact_8_37
timestamp 1624494425
transform 1 0 164 0 1 11949
box 0 0 64 64
use contact_9  contact_9_36
timestamp 1624494425
transform 1 0 163 0 1 11944
box 0 0 66 74
use contact_7  contact_7_43
timestamp 1624494425
transform 1 0 420 0 1 11948
box 0 0 58 66
use contact_8  contact_8_42
timestamp 1624494425
transform 1 0 417 0 1 11949
box 0 0 64 64
use contact_9  contact_9_40
timestamp 1624494425
transform 1 0 416 0 1 11944
box 0 0 66 74
use contact_7  contact_7_42
timestamp 1624494425
transform 1 0 788 0 1 11948
box 0 0 58 66
use contact_8  contact_8_41
timestamp 1624494425
transform 1 0 785 0 1 11949
box 0 0 64 64
use contact_9  contact_9_39
timestamp 1624494425
transform 1 0 784 0 1 11944
box 0 0 66 74
use contact_7  contact_7_5
timestamp 1624494425
transform 1 0 627 0 1 12693
box 0 0 58 66
use contact_8  contact_8_4
timestamp 1624494425
transform 1 0 624 0 1 12694
box 0 0 64 64
use contact_9  contact_9_3
timestamp 1624494425
transform 1 0 623 0 1 12689
box 0 0 66 74
use contact_7  contact_7_41
timestamp 1624494425
transform 1 0 1156 0 1 11948
box 0 0 58 66
use contact_8  contact_8_40
timestamp 1624494425
transform 1 0 1153 0 1 11949
box 0 0 64 64
use contact_9  contact_9_38
timestamp 1624494425
transform 1 0 1152 0 1 11944
box 0 0 66 74
use contact_7  contact_7_40
timestamp 1624494425
transform 1 0 1524 0 1 11948
box 0 0 58 66
use contact_8  contact_8_39
timestamp 1624494425
transform 1 0 1521 0 1 11949
box 0 0 64 64
use contact_9  contact_9_37
timestamp 1624494425
transform 1 0 1520 0 1 11944
box 0 0 66 74
use contact_7  contact_7_4
timestamp 1624494425
transform 1 0 1363 0 1 12693
box 0 0 58 66
use contact_8  contact_8_3
timestamp 1624494425
transform 1 0 1360 0 1 12694
box 0 0 64 64
use contact_9  contact_9_2
timestamp 1624494425
transform 1 0 1359 0 1 12689
box 0 0 66 74
use contact_7  contact_7_0
timestamp 1624494425
transform 1 0 1524 0 1 11948
box 0 0 58 66
<< labels >>
rlabel metal3 s 1343 7021 1441 7119 4 vdd
rlabel metal3 s 1343 1365 1441 1463 4 vdd
rlabel metal3 s 607 9849 705 9947 4 vdd
rlabel metal3 s 1343 9849 1441 9947 4 vdd
rlabel metal3 s 607 4193 705 4291 4 vdd
rlabel metal3 s 1343 4193 1441 4291 4 vdd
rlabel metal3 s 607 1365 705 1463 4 vdd
rlabel metal3 s 607 7021 705 7119 4 vdd
rlabel metal3 s 607 12677 705 12775 4 vdd
rlabel metal3 s 1343 12677 1441 12775 4 vdd
rlabel metal3 s 1343 5607 1441 5705 4 gnd
rlabel metal3 s 1343 8435 1441 8533 4 gnd
rlabel metal3 s 607 8435 705 8533 4 gnd
rlabel metal3 s 607 11263 705 11361 4 gnd
rlabel metal3 s 1343 11263 1441 11361 4 gnd
rlabel metal3 s 1343 2779 1441 2877 4 gnd
rlabel metal3 s 607 5607 705 5705 4 gnd
rlabel metal3 s 607 -49 705 49 4 gnd
rlabel metal3 s 1343 -49 1441 49 4 gnd
rlabel metal3 s 607 2779 705 2877 4 gnd
rlabel metal2 s -57 655 -29 683 4 in
rlabel metal1 s 1539 11967 1567 11995 4 out
<< properties >>
string FIXED_BBOX 0 0 1840 12726
<< end >>
