magic
tech sky130A
magscale 1 2
timestamp 1624426885
<< nwell >>
rect 25786 -42362 50302 -27620
rect 52120 -41876 58318 -38944
rect 52120 -43036 55580 -41876
rect 10260 -57542 12494 -56702
rect -27720 -67242 -25324 -64390
rect -23720 -67242 -21324 -64390
rect -19720 -67242 -17324 -64390
rect -15720 -67242 -13324 -64390
rect -11720 -67242 -9324 -64390
rect -7720 -67242 -5324 -64390
rect -3720 -67242 -1324 -64390
rect 280 -67242 2676 -64390
rect 4280 -67242 6676 -64390
rect -28112 -67566 -25324 -67242
rect -24112 -67566 -21324 -67242
rect -20112 -67566 -17324 -67242
rect -16112 -67566 -13324 -67242
rect -12112 -67566 -9324 -67242
rect -8112 -67566 -5324 -67242
rect -4112 -67566 -1324 -67242
rect -112 -67566 2676 -67242
rect 3888 -67566 6676 -67242
rect -28112 -72954 -25324 -72630
rect -24112 -72954 -21324 -72630
rect -20112 -72954 -17324 -72630
rect -16112 -72954 -13324 -72630
rect -12112 -72954 -9324 -72630
rect -8112 -72954 -5324 -72630
rect -4112 -72954 -1324 -72630
rect -112 -72954 2676 -72630
rect 3888 -72954 6676 -72630
rect -27720 -75806 -25324 -72954
rect -23720 -75806 -21324 -72954
rect -19720 -75806 -17324 -72954
rect -15720 -75806 -13324 -72954
rect -11720 -75806 -9324 -72954
rect -7720 -75806 -5324 -72954
rect -3720 -75806 -1324 -72954
rect 280 -75806 2676 -72954
rect 4280 -75806 6676 -72954
<< pwell >>
rect 55864 -41933 56834 -41932
rect 55864 -41942 56931 -41933
rect 56952 -41942 58318 -41932
rect 12118 -57600 12148 -57598
rect 12198 -57599 12410 -57598
rect 12198 -57600 12414 -57599
rect 12118 -57636 12414 -57600
rect 10260 -57785 12414 -57636
rect 10260 -57819 12427 -57785
rect 10260 -58256 12410 -57819
rect 13086 -59236 50402 -43120
rect 55864 -43922 58318 -41942
rect -28030 -67730 -27844 -67623
rect -24030 -67730 -23844 -67623
rect -20030 -67730 -19844 -67623
rect -16030 -67730 -15844 -67623
rect -12030 -67730 -11844 -67623
rect -8030 -67730 -7844 -67623
rect -4030 -67730 -3844 -67623
rect -30 -67730 156 -67623
rect 3970 -67730 4156 -67623
rect -28032 -67809 -25324 -67730
rect -24032 -67809 -21324 -67730
rect -20032 -67809 -17324 -67730
rect -16032 -67809 -13324 -67730
rect -12032 -67809 -9324 -67730
rect -8032 -67809 -5324 -67730
rect -4032 -67809 -1324 -67730
rect -32 -67809 2676 -67730
rect 3968 -67809 6676 -67730
rect -28043 -67843 -25324 -67809
rect -24043 -67843 -21324 -67809
rect -20043 -67843 -17324 -67809
rect -16043 -67843 -13324 -67809
rect -12043 -67843 -9324 -67809
rect -8043 -67843 -5324 -67809
rect -4043 -67843 -1324 -67809
rect -43 -67843 2676 -67809
rect 3957 -67843 6676 -67809
rect -28032 -67874 -25324 -67843
rect -24032 -67874 -21324 -67843
rect -20032 -67874 -17324 -67843
rect -16032 -67874 -13324 -67843
rect -12032 -67874 -9324 -67843
rect -8032 -67874 -5324 -67843
rect -4032 -67874 -1324 -67843
rect -32 -67874 2676 -67843
rect 3968 -67874 6676 -67843
rect -27720 -69846 -25324 -67874
rect -23720 -69846 -21324 -67874
rect -19720 -69846 -17324 -67874
rect -15720 -69846 -13324 -67874
rect -11720 -69846 -9324 -67874
rect -7720 -69846 -5324 -67874
rect -3720 -69846 -1324 -67874
rect 280 -69846 2676 -67874
rect 4280 -69846 6676 -67874
rect -27720 -72322 -25324 -70350
rect -23720 -72322 -21324 -70350
rect -19720 -72322 -17324 -70350
rect -15720 -72322 -13324 -70350
rect -11720 -72322 -9324 -70350
rect -7720 -72322 -5324 -70350
rect -3720 -72322 -1324 -70350
rect 280 -72322 2676 -70350
rect 4280 -72322 6676 -70350
rect -28032 -72353 -25324 -72322
rect -24032 -72353 -21324 -72322
rect -20032 -72353 -17324 -72322
rect -16032 -72353 -13324 -72322
rect -12032 -72353 -9324 -72322
rect -8032 -72353 -5324 -72322
rect -4032 -72353 -1324 -72322
rect -32 -72353 2676 -72322
rect 3968 -72353 6676 -72322
rect -28043 -72387 -25324 -72353
rect -24043 -72387 -21324 -72353
rect -20043 -72387 -17324 -72353
rect -16043 -72387 -13324 -72353
rect -12043 -72387 -9324 -72353
rect -8043 -72387 -5324 -72353
rect -4043 -72387 -1324 -72353
rect -43 -72387 2676 -72353
rect 3957 -72387 6676 -72353
rect -28032 -72466 -25324 -72387
rect -24032 -72466 -21324 -72387
rect -20032 -72466 -17324 -72387
rect -16032 -72466 -13324 -72387
rect -12032 -72466 -9324 -72387
rect -8032 -72466 -5324 -72387
rect -4032 -72466 -1324 -72387
rect -32 -72466 2676 -72387
rect 3968 -72466 6676 -72387
rect -28030 -72573 -27844 -72466
rect -24030 -72573 -23844 -72466
rect -20030 -72573 -19844 -72466
rect -16030 -72573 -15844 -72466
rect -12030 -72573 -11844 -72466
rect -8030 -72573 -7844 -72466
rect -4030 -72573 -3844 -72466
rect -30 -72573 156 -72466
rect 3970 -72573 4156 -72466
<< nmos >>
rect 56062 -42902 56122 -42702
rect 56608 -42816 56668 -42616
rect 56726 -42816 56786 -42616
rect 56844 -42816 56904 -42616
rect 56962 -42816 57022 -42616
rect 57080 -42816 57140 -42616
rect 57198 -42816 57258 -42616
rect 57316 -42816 57376 -42616
rect 57434 -42816 57494 -42616
rect 10456 -58046 10656 -57846
rect 10714 -58046 10914 -57846
rect 10972 -58046 11172 -57846
rect 11230 -58046 11430 -57846
rect 11488 -58046 11688 -57846
rect 11746 -58046 11946 -57846
rect 28072 -44614 29032 -44014
rect 29090 -44614 30050 -44014
rect 30108 -44614 31068 -44014
rect 31126 -44614 32086 -44014
rect 32144 -44614 33104 -44014
rect 33162 -44614 34122 -44014
rect 34180 -44614 35140 -44014
rect 35198 -44614 36158 -44014
rect 36216 -44614 37176 -44014
rect 37234 -44614 38194 -44014
rect 38252 -44614 39212 -44014
rect 39270 -44614 40230 -44014
rect 40288 -44614 41248 -44014
rect 41306 -44614 42266 -44014
rect 42324 -44614 43284 -44014
rect 43342 -44614 44302 -44014
rect 44360 -44614 45320 -44014
rect 45378 -44614 46338 -44014
rect 46396 -44614 47356 -44014
rect 47414 -44614 48374 -44014
rect 28072 -45432 29032 -44832
rect 29090 -45432 30050 -44832
rect 30108 -45432 31068 -44832
rect 31126 -45432 32086 -44832
rect 32144 -45432 33104 -44832
rect 33162 -45432 34122 -44832
rect 34180 -45432 35140 -44832
rect 35198 -45432 36158 -44832
rect 36216 -45432 37176 -44832
rect 37234 -45432 38194 -44832
rect 38252 -45432 39212 -44832
rect 39270 -45432 40230 -44832
rect 40288 -45432 41248 -44832
rect 41306 -45432 42266 -44832
rect 42324 -45432 43284 -44832
rect 43342 -45432 44302 -44832
rect 44360 -45432 45320 -44832
rect 45378 -45432 46338 -44832
rect 46396 -45432 47356 -44832
rect 47414 -45432 48374 -44832
rect 28072 -46810 29032 -46210
rect 29090 -46810 30050 -46210
rect 30108 -46810 31068 -46210
rect 31126 -46810 32086 -46210
rect 32144 -46810 33104 -46210
rect 33162 -46810 34122 -46210
rect 34180 -46810 35140 -46210
rect 35198 -46810 36158 -46210
rect 36216 -46810 37176 -46210
rect 37234 -46810 38194 -46210
rect 38252 -46810 39212 -46210
rect 39270 -46810 40230 -46210
rect 40288 -46810 41248 -46210
rect 41306 -46810 42266 -46210
rect 42324 -46810 43284 -46210
rect 43342 -46810 44302 -46210
rect 44360 -46810 45320 -46210
rect 45378 -46810 46338 -46210
rect 46396 -46810 47356 -46210
rect 47414 -46810 48374 -46210
rect 28072 -48042 29032 -47442
rect 29090 -48042 30050 -47442
rect 30108 -48042 31068 -47442
rect 31126 -48042 32086 -47442
rect 32144 -48042 33104 -47442
rect 33162 -48042 34122 -47442
rect 34180 -48042 35140 -47442
rect 35198 -48042 36158 -47442
rect 36216 -48042 37176 -47442
rect 37234 -48042 38194 -47442
rect 38252 -48042 39212 -47442
rect 39270 -48042 40230 -47442
rect 40288 -48042 41248 -47442
rect 41306 -48042 42266 -47442
rect 42324 -48042 43284 -47442
rect 43342 -48042 44302 -47442
rect 44360 -48042 45320 -47442
rect 45378 -48042 46338 -47442
rect 46396 -48042 47356 -47442
rect 47414 -48042 48374 -47442
rect 28070 -49276 29030 -48676
rect 29088 -49276 30048 -48676
rect 30106 -49276 31066 -48676
rect 31124 -49276 32084 -48676
rect 32142 -49276 33102 -48676
rect 33160 -49276 34120 -48676
rect 34178 -49276 35138 -48676
rect 35196 -49276 36156 -48676
rect 36214 -49276 37174 -48676
rect 37232 -49276 38192 -48676
rect 38250 -49276 39210 -48676
rect 39268 -49276 40228 -48676
rect 40286 -49276 41246 -48676
rect 41304 -49276 42264 -48676
rect 42322 -49276 43282 -48676
rect 43340 -49276 44300 -48676
rect 44358 -49276 45318 -48676
rect 45376 -49276 46336 -48676
rect 46394 -49276 47354 -48676
rect 47412 -49276 48372 -48676
rect 28070 -50510 29030 -49910
rect 29088 -50510 30048 -49910
rect 30106 -50510 31066 -49910
rect 31124 -50510 32084 -49910
rect 32142 -50510 33102 -49910
rect 33160 -50510 34120 -49910
rect 34178 -50510 35138 -49910
rect 35196 -50510 36156 -49910
rect 36214 -50510 37174 -49910
rect 37232 -50510 38192 -49910
rect 38250 -50510 39210 -49910
rect 39268 -50510 40228 -49910
rect 40286 -50510 41246 -49910
rect 41304 -50510 42264 -49910
rect 42322 -50510 43282 -49910
rect 43340 -50510 44300 -49910
rect 44358 -50510 45318 -49910
rect 45376 -50510 46336 -49910
rect 46394 -50510 47354 -49910
rect 47412 -50510 48372 -49910
rect 28070 -51742 29030 -51142
rect 29088 -51742 30048 -51142
rect 30106 -51742 31066 -51142
rect 31124 -51742 32084 -51142
rect 32142 -51742 33102 -51142
rect 33160 -51742 34120 -51142
rect 34178 -51742 35138 -51142
rect 35196 -51742 36156 -51142
rect 36214 -51742 37174 -51142
rect 37232 -51742 38192 -51142
rect 38250 -51742 39210 -51142
rect 39268 -51742 40228 -51142
rect 40286 -51742 41246 -51142
rect 41304 -51742 42264 -51142
rect 42322 -51742 43282 -51142
rect 43340 -51742 44300 -51142
rect 44358 -51742 45318 -51142
rect 45376 -51742 46336 -51142
rect 46394 -51742 47354 -51142
rect 47412 -51742 48372 -51142
rect 28070 -52976 29030 -52376
rect 29088 -52976 30048 -52376
rect 30106 -52976 31066 -52376
rect 31124 -52976 32084 -52376
rect 32142 -52976 33102 -52376
rect 33160 -52976 34120 -52376
rect 34178 -52976 35138 -52376
rect 35196 -52976 36156 -52376
rect 36214 -52976 37174 -52376
rect 37232 -52976 38192 -52376
rect 38250 -52976 39210 -52376
rect 39268 -52976 40228 -52376
rect 40286 -52976 41246 -52376
rect 41304 -52976 42264 -52376
rect 42322 -52976 43282 -52376
rect 43340 -52976 44300 -52376
rect 44358 -52976 45318 -52376
rect 45376 -52976 46336 -52376
rect 46394 -52976 47354 -52376
rect 47412 -52976 48372 -52376
rect 28070 -54210 29030 -53610
rect 29088 -54210 30048 -53610
rect 30106 -54210 31066 -53610
rect 31124 -54210 32084 -53610
rect 32142 -54210 33102 -53610
rect 33160 -54210 34120 -53610
rect 34178 -54210 35138 -53610
rect 35196 -54210 36156 -53610
rect 36214 -54210 37174 -53610
rect 37232 -54210 38192 -53610
rect 38250 -54210 39210 -53610
rect 39268 -54210 40228 -53610
rect 40286 -54210 41246 -53610
rect 41304 -54210 42264 -53610
rect 42322 -54210 43282 -53610
rect 43340 -54210 44300 -53610
rect 44358 -54210 45318 -53610
rect 45376 -54210 46336 -53610
rect 46394 -54210 47354 -53610
rect 47412 -54210 48372 -53610
rect 28070 -55442 29030 -54842
rect 29088 -55442 30048 -54842
rect 30106 -55442 31066 -54842
rect 31124 -55442 32084 -54842
rect 32142 -55442 33102 -54842
rect 33160 -55442 34120 -54842
rect 34178 -55442 35138 -54842
rect 35196 -55442 36156 -54842
rect 36214 -55442 37174 -54842
rect 37232 -55442 38192 -54842
rect 38250 -55442 39210 -54842
rect 39268 -55442 40228 -54842
rect 40286 -55442 41246 -54842
rect 41304 -55442 42264 -54842
rect 42322 -55442 43282 -54842
rect 43340 -55442 44300 -54842
rect 44358 -55442 45318 -54842
rect 45376 -55442 46336 -54842
rect 46394 -55442 47354 -54842
rect 47412 -55442 48372 -54842
rect 28070 -56676 29030 -56076
rect 29088 -56676 30048 -56076
rect 30106 -56676 31066 -56076
rect 31124 -56676 32084 -56076
rect 32142 -56676 33102 -56076
rect 33160 -56676 34120 -56076
rect 34178 -56676 35138 -56076
rect 35196 -56676 36156 -56076
rect 36214 -56676 37174 -56076
rect 37232 -56676 38192 -56076
rect 38250 -56676 39210 -56076
rect 39268 -56676 40228 -56076
rect 40286 -56676 41246 -56076
rect 41304 -56676 42264 -56076
rect 42322 -56676 43282 -56076
rect 43340 -56676 44300 -56076
rect 44358 -56676 45318 -56076
rect 45376 -56676 46336 -56076
rect 46394 -56676 47354 -56076
rect 47412 -56676 48372 -56076
rect 15440 -57718 16400 -57118
rect 16458 -57718 17418 -57118
rect 17476 -57718 18436 -57118
rect 18494 -57718 19454 -57118
rect 19512 -57718 20472 -57118
rect 20530 -57718 21490 -57118
rect 21548 -57718 22508 -57118
rect 22566 -57718 23526 -57118
rect 23584 -57718 24544 -57118
rect 24602 -57718 25562 -57118
rect 28070 -57908 29030 -57308
rect 29088 -57908 30048 -57308
rect 30106 -57908 31066 -57308
rect 31124 -57908 32084 -57308
rect 32142 -57908 33102 -57308
rect 33160 -57908 34120 -57308
rect 34178 -57908 35138 -57308
rect 35196 -57908 36156 -57308
rect 36214 -57908 37174 -57308
rect 37232 -57908 38192 -57308
rect 38250 -57908 39210 -57308
rect 39268 -57908 40228 -57308
rect 40286 -57908 41246 -57308
rect 41304 -57908 42264 -57308
rect 42322 -57908 43282 -57308
rect 43340 -57908 44300 -57308
rect 44358 -57908 45318 -57308
rect 45376 -57908 46336 -57308
rect 46394 -57908 47354 -57308
rect 47412 -57908 48372 -57308
rect 57966 -42902 58026 -42702
rect -27296 -68718 -27096 -68318
rect -27038 -68718 -26838 -68318
rect -26780 -68718 -26580 -68318
rect -26522 -68718 -26322 -68318
rect -26264 -68718 -26064 -68318
rect -26006 -68718 -25806 -68318
rect -23296 -68718 -23096 -68318
rect -23038 -68718 -22838 -68318
rect -22780 -68718 -22580 -68318
rect -22522 -68718 -22322 -68318
rect -22264 -68718 -22064 -68318
rect -22006 -68718 -21806 -68318
rect -19296 -68718 -19096 -68318
rect -19038 -68718 -18838 -68318
rect -18780 -68718 -18580 -68318
rect -18522 -68718 -18322 -68318
rect -18264 -68718 -18064 -68318
rect -18006 -68718 -17806 -68318
rect -15296 -68718 -15096 -68318
rect -15038 -68718 -14838 -68318
rect -14780 -68718 -14580 -68318
rect -14522 -68718 -14322 -68318
rect -14264 -68718 -14064 -68318
rect -14006 -68718 -13806 -68318
rect -11296 -68718 -11096 -68318
rect -11038 -68718 -10838 -68318
rect -10780 -68718 -10580 -68318
rect -10522 -68718 -10322 -68318
rect -10264 -68718 -10064 -68318
rect -10006 -68718 -9806 -68318
rect -7296 -68718 -7096 -68318
rect -7038 -68718 -6838 -68318
rect -6780 -68718 -6580 -68318
rect -6522 -68718 -6322 -68318
rect -6264 -68718 -6064 -68318
rect -6006 -68718 -5806 -68318
rect -3296 -68718 -3096 -68318
rect -3038 -68718 -2838 -68318
rect -2780 -68718 -2580 -68318
rect -2522 -68718 -2322 -68318
rect -2264 -68718 -2064 -68318
rect -2006 -68718 -1806 -68318
rect 704 -68718 904 -68318
rect 962 -68718 1162 -68318
rect 1220 -68718 1420 -68318
rect 1478 -68718 1678 -68318
rect 1736 -68718 1936 -68318
rect 1994 -68718 2194 -68318
rect 4704 -68718 4904 -68318
rect 4962 -68718 5162 -68318
rect 5220 -68718 5420 -68318
rect 5478 -68718 5678 -68318
rect 5736 -68718 5936 -68318
rect 5994 -68718 6194 -68318
rect -27296 -71878 -27096 -71478
rect -27038 -71878 -26838 -71478
rect -26780 -71878 -26580 -71478
rect -26522 -71878 -26322 -71478
rect -26264 -71878 -26064 -71478
rect -26006 -71878 -25806 -71478
rect -23296 -71878 -23096 -71478
rect -23038 -71878 -22838 -71478
rect -22780 -71878 -22580 -71478
rect -22522 -71878 -22322 -71478
rect -22264 -71878 -22064 -71478
rect -22006 -71878 -21806 -71478
rect -19296 -71878 -19096 -71478
rect -19038 -71878 -18838 -71478
rect -18780 -71878 -18580 -71478
rect -18522 -71878 -18322 -71478
rect -18264 -71878 -18064 -71478
rect -18006 -71878 -17806 -71478
rect -15296 -71878 -15096 -71478
rect -15038 -71878 -14838 -71478
rect -14780 -71878 -14580 -71478
rect -14522 -71878 -14322 -71478
rect -14264 -71878 -14064 -71478
rect -14006 -71878 -13806 -71478
rect -11296 -71878 -11096 -71478
rect -11038 -71878 -10838 -71478
rect -10780 -71878 -10580 -71478
rect -10522 -71878 -10322 -71478
rect -10264 -71878 -10064 -71478
rect -10006 -71878 -9806 -71478
rect -7296 -71878 -7096 -71478
rect -7038 -71878 -6838 -71478
rect -6780 -71878 -6580 -71478
rect -6522 -71878 -6322 -71478
rect -6264 -71878 -6064 -71478
rect -6006 -71878 -5806 -71478
rect -3296 -71878 -3096 -71478
rect -3038 -71878 -2838 -71478
rect -2780 -71878 -2580 -71478
rect -2522 -71878 -2322 -71478
rect -2264 -71878 -2064 -71478
rect -2006 -71878 -1806 -71478
rect 704 -71878 904 -71478
rect 962 -71878 1162 -71478
rect 1220 -71878 1420 -71478
rect 1478 -71878 1678 -71478
rect 1736 -71878 1936 -71478
rect 1994 -71878 2194 -71478
rect 4704 -71878 4904 -71478
rect 4962 -71878 5162 -71478
rect 5220 -71878 5420 -71478
rect 5478 -71878 5678 -71478
rect 5736 -71878 5936 -71478
rect 5994 -71878 6194 -71478
<< scnmos >>
rect 56224 -42089 56254 -41959
rect 56500 -42089 56530 -41959
rect 56739 -42089 56769 -41959
rect 56823 -42089 56853 -41959
rect 57197 -42089 57227 -41959
rect 57281 -42089 57311 -41959
rect 57520 -42089 57550 -41959
rect 57796 -42089 57826 -41959
rect 12306 -57755 12336 -57625
rect -27952 -67779 -27922 -67649
rect -23952 -67779 -23922 -67649
rect -19952 -67779 -19922 -67649
rect -15952 -67779 -15922 -67649
rect -11952 -67779 -11922 -67649
rect -7952 -67779 -7922 -67649
rect -3952 -67779 -3922 -67649
rect 48 -67779 78 -67649
rect 4048 -67779 4078 -67649
rect -27952 -72547 -27922 -72417
rect -23952 -72547 -23922 -72417
rect -19952 -72547 -19922 -72417
rect -15952 -72547 -15922 -72417
rect -11952 -72547 -11922 -72417
rect -7952 -72547 -7922 -72417
rect -3952 -72547 -3922 -72417
rect 48 -72547 78 -72417
rect 4048 -72547 4078 -72417
<< pmos >>
rect 32964 -37650 33924 -37050
rect 33982 -37650 34942 -37050
rect 35000 -37650 35960 -37050
rect 36018 -37650 36978 -37050
rect 37036 -37650 37996 -37050
rect 38054 -37650 39014 -37050
rect 39072 -37650 40032 -37050
rect 40090 -37650 41050 -37050
rect 41108 -37650 42068 -37050
rect 42126 -37650 43086 -37050
rect 43144 -37650 44104 -37050
rect 44162 -37650 45122 -37050
rect 45180 -37650 46140 -37050
rect 46198 -37650 47158 -37050
rect 47216 -37650 48176 -37050
rect 32964 -38906 33924 -38306
rect 33982 -38906 34942 -38306
rect 35000 -38906 35960 -38306
rect 36018 -38906 36978 -38306
rect 37036 -38906 37996 -38306
rect 38054 -38906 39014 -38306
rect 39072 -38906 40032 -38306
rect 40090 -38906 41050 -38306
rect 41108 -38906 42068 -38306
rect 42126 -38906 43086 -38306
rect 43144 -38906 44104 -38306
rect 44162 -38906 45122 -38306
rect 45180 -38906 46140 -38306
rect 46198 -38906 47158 -38306
rect 47216 -38906 48176 -38306
rect 32964 -40162 33924 -39562
rect 33982 -40162 34942 -39562
rect 35000 -40162 35960 -39562
rect 36018 -40162 36978 -39562
rect 37036 -40162 37996 -39562
rect 38054 -40162 39014 -39562
rect 39072 -40162 40032 -39562
rect 40090 -40162 41050 -39562
rect 41108 -40162 42068 -39562
rect 42126 -40162 43086 -39562
rect 43144 -40162 44104 -39562
rect 44162 -40162 45122 -39562
rect 45180 -40162 46140 -39562
rect 46198 -40162 47158 -39562
rect 47216 -40162 48176 -39562
rect 32964 -41418 33924 -40818
rect 33982 -41418 34942 -40818
rect 35000 -41418 35960 -40818
rect 36018 -41418 36978 -40818
rect 37036 -41418 37996 -40818
rect 38054 -41418 39014 -40818
rect 39072 -41418 40032 -40818
rect 40090 -41418 41050 -40818
rect 41108 -41418 42068 -40818
rect 42126 -41418 43086 -40818
rect 43144 -41418 44104 -40818
rect 44162 -41418 45122 -40818
rect 45180 -41418 46140 -40818
rect 46198 -41418 47158 -40818
rect 47216 -41418 48176 -40818
rect 52488 -39880 52888 -39680
rect 52946 -39880 53346 -39680
rect 53404 -39880 53804 -39680
rect 53862 -39880 54262 -39680
rect 54320 -39880 54720 -39680
rect 54778 -39880 55178 -39680
rect 56116 -40280 56316 -39880
rect 56374 -40280 56574 -39880
rect 56632 -40280 56832 -39880
rect 56890 -40280 57090 -39880
rect 57148 -40280 57348 -39880
rect 57406 -40280 57606 -39880
rect 57664 -40280 57864 -39880
rect 56116 -41140 56316 -40740
rect 56374 -41140 56574 -40740
rect 56632 -41140 56832 -40740
rect 56890 -41140 57090 -40740
rect 57148 -41140 57348 -40740
rect 57406 -41140 57606 -40740
rect 57664 -41140 57864 -40740
<< scpmoshvt >>
rect 56224 -41839 56254 -41639
rect 56500 -41839 56530 -41639
rect 56739 -41839 56769 -41639
rect 56823 -41839 56853 -41639
rect 57197 -41839 57227 -41639
rect 57281 -41839 57311 -41639
rect 57520 -41839 57550 -41639
rect 57796 -41839 57826 -41639
rect 12306 -57505 12336 -57305
rect -27952 -67529 -27922 -67329
rect -23952 -67529 -23922 -67329
rect -19952 -67529 -19922 -67329
rect -15952 -67529 -15922 -67329
rect -11952 -67529 -11922 -67329
rect -7952 -67529 -7922 -67329
rect -3952 -67529 -3922 -67329
rect 48 -67529 78 -67329
rect 4048 -67529 4078 -67329
rect -27952 -72867 -27922 -72667
rect -23952 -72867 -23922 -72667
rect -19952 -72867 -19922 -72667
rect -15952 -72867 -15922 -72667
rect -11952 -72867 -11922 -72667
rect -7952 -72867 -7922 -72667
rect -3952 -72867 -3922 -72667
rect 48 -72867 78 -72667
rect 4048 -72867 4078 -72667
<< pmoslvt >>
rect 31978 -31104 32938 -30504
rect 32996 -31104 33956 -30504
rect 34014 -31104 34974 -30504
rect 35032 -31104 35992 -30504
rect 36050 -31104 37010 -30504
rect 37068 -31104 38028 -30504
rect 38086 -31104 39046 -30504
rect 39104 -31104 40064 -30504
rect 40122 -31104 41082 -30504
rect 41140 -31104 42100 -30504
rect 42158 -31104 43118 -30504
rect 43176 -31104 44136 -30504
rect 44194 -31104 45154 -30504
rect 45212 -31104 46172 -30504
rect 46230 -31104 47190 -30504
rect 47248 -31104 48208 -30504
rect 31978 -32240 32938 -31640
rect 32996 -32240 33956 -31640
rect 34014 -32240 34974 -31640
rect 35032 -32240 35992 -31640
rect 36050 -32240 37010 -31640
rect 37068 -32240 38028 -31640
rect 38086 -32240 39046 -31640
rect 39104 -32240 40064 -31640
rect 40122 -32240 41082 -31640
rect 41140 -32240 42100 -31640
rect 42158 -32240 43118 -31640
rect 43176 -32240 44136 -31640
rect 44194 -32240 45154 -31640
rect 45212 -32240 46172 -31640
rect 46230 -32240 47190 -31640
rect 47248 -32240 48208 -31640
rect 31978 -33376 32938 -32776
rect 32996 -33376 33956 -32776
rect 34014 -33376 34974 -32776
rect 35032 -33376 35992 -32776
rect 36050 -33376 37010 -32776
rect 37068 -33376 38028 -32776
rect 38086 -33376 39046 -32776
rect 39104 -33376 40064 -32776
rect 40122 -33376 41082 -32776
rect 41140 -33376 42100 -32776
rect 42158 -33376 43118 -32776
rect 43176 -33376 44136 -32776
rect 44194 -33376 45154 -32776
rect 45212 -33376 46172 -32776
rect 46230 -33376 47190 -32776
rect 47248 -33376 48208 -32776
rect 33172 -35014 34132 -34414
rect 34190 -35014 35150 -34414
rect 35208 -35014 36168 -34414
rect 36226 -35014 37186 -34414
rect 37244 -35014 38204 -34414
rect 38262 -35014 39222 -34414
rect 39280 -35014 40240 -34414
rect 40298 -35014 41258 -34414
rect 41316 -35014 42276 -34414
rect 42334 -35014 43294 -34414
rect 43352 -35014 44312 -34414
rect 44370 -35014 45330 -34414
rect 45388 -35014 46348 -34414
rect 46406 -35014 47366 -34414
rect 33172 -36046 34132 -35446
rect 34190 -36046 35150 -35446
rect 35208 -36046 36168 -35446
rect 36226 -36046 37186 -35446
rect 37244 -36046 38204 -35446
rect 38262 -36046 39222 -35446
rect 39280 -36046 40240 -35446
rect 40298 -36046 41258 -35446
rect 41316 -36046 42276 -35446
rect 42334 -36046 43294 -35446
rect 43352 -36046 44312 -35446
rect 44370 -36046 45330 -35446
rect 45388 -36046 46348 -35446
rect 46406 -36046 47366 -35446
rect 27660 -37754 28620 -37154
rect 28678 -37754 29638 -37154
rect 29696 -37754 30656 -37154
rect 30714 -37754 31674 -37154
rect 27660 -38786 28620 -38186
rect 28678 -38786 29638 -38186
rect 29696 -38786 30656 -38186
rect 30714 -38786 31674 -38186
rect 27660 -39818 28620 -39218
rect 28678 -39818 29638 -39218
rect 29696 -39818 30656 -39218
rect 30714 -39818 31674 -39218
rect 27660 -40850 28620 -40250
rect 28678 -40850 29638 -40250
rect 29696 -40850 30656 -40250
rect 30714 -40850 31674 -40250
rect 52547 -40963 52747 -40563
rect 52805 -40963 53005 -40563
rect 53063 -40963 53263 -40563
rect 53321 -40963 53521 -40563
rect 53579 -40963 53779 -40563
rect 53837 -40963 54037 -40563
rect 54095 -40963 54295 -40563
rect 54353 -40963 54553 -40563
rect 54611 -40963 54811 -40563
rect 54869 -40963 55069 -40563
rect 52547 -41823 52747 -41423
rect 52805 -41823 53005 -41423
rect 53063 -41823 53263 -41423
rect 53321 -41823 53521 -41423
rect 53579 -41823 53779 -41423
rect 53837 -41823 54037 -41423
rect 54095 -41823 54295 -41423
rect 54353 -41823 54553 -41423
rect 54611 -41823 54811 -41423
rect 54869 -41823 55069 -41423
rect 54264 -42794 54334 -42594
rect 54392 -42794 54462 -42594
rect 54520 -42794 54590 -42594
rect 54648 -42794 54718 -42594
rect 54776 -42794 54846 -42594
rect 54904 -42794 54974 -42594
rect 55032 -42794 55102 -42594
rect 55160 -42794 55230 -42594
rect 55288 -42794 55358 -42594
<< pmoshvt >>
rect 10456 -57322 10656 -56922
rect 10714 -57322 10914 -56922
rect 10972 -57322 11172 -56922
rect 11230 -57322 11430 -56922
rect 11488 -57322 11688 -56922
rect 11746 -57322 11946 -56922
rect -27291 -66025 -27091 -65625
rect -27033 -66025 -26833 -65625
rect -26775 -66025 -26575 -65625
rect -26517 -66025 -26317 -65625
rect -26259 -66025 -26059 -65625
rect -26001 -66025 -25801 -65625
rect -27291 -66885 -27091 -66485
rect -27033 -66885 -26833 -66485
rect -26775 -66885 -26575 -66485
rect -26517 -66885 -26317 -66485
rect -26259 -66885 -26059 -66485
rect -26001 -66885 -25801 -66485
rect -23291 -66025 -23091 -65625
rect -23033 -66025 -22833 -65625
rect -22775 -66025 -22575 -65625
rect -22517 -66025 -22317 -65625
rect -22259 -66025 -22059 -65625
rect -22001 -66025 -21801 -65625
rect -23291 -66885 -23091 -66485
rect -23033 -66885 -22833 -66485
rect -22775 -66885 -22575 -66485
rect -22517 -66885 -22317 -66485
rect -22259 -66885 -22059 -66485
rect -22001 -66885 -21801 -66485
rect -19291 -66025 -19091 -65625
rect -19033 -66025 -18833 -65625
rect -18775 -66025 -18575 -65625
rect -18517 -66025 -18317 -65625
rect -18259 -66025 -18059 -65625
rect -18001 -66025 -17801 -65625
rect -19291 -66885 -19091 -66485
rect -19033 -66885 -18833 -66485
rect -18775 -66885 -18575 -66485
rect -18517 -66885 -18317 -66485
rect -18259 -66885 -18059 -66485
rect -18001 -66885 -17801 -66485
rect -15291 -66025 -15091 -65625
rect -15033 -66025 -14833 -65625
rect -14775 -66025 -14575 -65625
rect -14517 -66025 -14317 -65625
rect -14259 -66025 -14059 -65625
rect -14001 -66025 -13801 -65625
rect -15291 -66885 -15091 -66485
rect -15033 -66885 -14833 -66485
rect -14775 -66885 -14575 -66485
rect -14517 -66885 -14317 -66485
rect -14259 -66885 -14059 -66485
rect -14001 -66885 -13801 -66485
rect -11291 -66025 -11091 -65625
rect -11033 -66025 -10833 -65625
rect -10775 -66025 -10575 -65625
rect -10517 -66025 -10317 -65625
rect -10259 -66025 -10059 -65625
rect -10001 -66025 -9801 -65625
rect -11291 -66885 -11091 -66485
rect -11033 -66885 -10833 -66485
rect -10775 -66885 -10575 -66485
rect -10517 -66885 -10317 -66485
rect -10259 -66885 -10059 -66485
rect -10001 -66885 -9801 -66485
rect -7291 -66025 -7091 -65625
rect -7033 -66025 -6833 -65625
rect -6775 -66025 -6575 -65625
rect -6517 -66025 -6317 -65625
rect -6259 -66025 -6059 -65625
rect -6001 -66025 -5801 -65625
rect -7291 -66885 -7091 -66485
rect -7033 -66885 -6833 -66485
rect -6775 -66885 -6575 -66485
rect -6517 -66885 -6317 -66485
rect -6259 -66885 -6059 -66485
rect -6001 -66885 -5801 -66485
rect -3291 -66025 -3091 -65625
rect -3033 -66025 -2833 -65625
rect -2775 -66025 -2575 -65625
rect -2517 -66025 -2317 -65625
rect -2259 -66025 -2059 -65625
rect -2001 -66025 -1801 -65625
rect -3291 -66885 -3091 -66485
rect -3033 -66885 -2833 -66485
rect -2775 -66885 -2575 -66485
rect -2517 -66885 -2317 -66485
rect -2259 -66885 -2059 -66485
rect -2001 -66885 -1801 -66485
rect 709 -66025 909 -65625
rect 967 -66025 1167 -65625
rect 1225 -66025 1425 -65625
rect 1483 -66025 1683 -65625
rect 1741 -66025 1941 -65625
rect 1999 -66025 2199 -65625
rect 709 -66885 909 -66485
rect 967 -66885 1167 -66485
rect 1225 -66885 1425 -66485
rect 1483 -66885 1683 -66485
rect 1741 -66885 1941 -66485
rect 1999 -66885 2199 -66485
rect 4709 -66025 4909 -65625
rect 4967 -66025 5167 -65625
rect 5225 -66025 5425 -65625
rect 5483 -66025 5683 -65625
rect 5741 -66025 5941 -65625
rect 5999 -66025 6199 -65625
rect 4709 -66885 4909 -66485
rect 4967 -66885 5167 -66485
rect 5225 -66885 5425 -66485
rect 5483 -66885 5683 -66485
rect 5741 -66885 5941 -66485
rect 5999 -66885 6199 -66485
rect -27291 -73711 -27091 -73311
rect -27033 -73711 -26833 -73311
rect -26775 -73711 -26575 -73311
rect -26517 -73711 -26317 -73311
rect -26259 -73711 -26059 -73311
rect -26001 -73711 -25801 -73311
rect -27291 -74571 -27091 -74171
rect -27033 -74571 -26833 -74171
rect -26775 -74571 -26575 -74171
rect -26517 -74571 -26317 -74171
rect -26259 -74571 -26059 -74171
rect -26001 -74571 -25801 -74171
rect -23291 -73711 -23091 -73311
rect -23033 -73711 -22833 -73311
rect -22775 -73711 -22575 -73311
rect -22517 -73711 -22317 -73311
rect -22259 -73711 -22059 -73311
rect -22001 -73711 -21801 -73311
rect -23291 -74571 -23091 -74171
rect -23033 -74571 -22833 -74171
rect -22775 -74571 -22575 -74171
rect -22517 -74571 -22317 -74171
rect -22259 -74571 -22059 -74171
rect -22001 -74571 -21801 -74171
rect -19291 -73711 -19091 -73311
rect -19033 -73711 -18833 -73311
rect -18775 -73711 -18575 -73311
rect -18517 -73711 -18317 -73311
rect -18259 -73711 -18059 -73311
rect -18001 -73711 -17801 -73311
rect -19291 -74571 -19091 -74171
rect -19033 -74571 -18833 -74171
rect -18775 -74571 -18575 -74171
rect -18517 -74571 -18317 -74171
rect -18259 -74571 -18059 -74171
rect -18001 -74571 -17801 -74171
rect -15291 -73711 -15091 -73311
rect -15033 -73711 -14833 -73311
rect -14775 -73711 -14575 -73311
rect -14517 -73711 -14317 -73311
rect -14259 -73711 -14059 -73311
rect -14001 -73711 -13801 -73311
rect -15291 -74571 -15091 -74171
rect -15033 -74571 -14833 -74171
rect -14775 -74571 -14575 -74171
rect -14517 -74571 -14317 -74171
rect -14259 -74571 -14059 -74171
rect -14001 -74571 -13801 -74171
rect -11291 -73711 -11091 -73311
rect -11033 -73711 -10833 -73311
rect -10775 -73711 -10575 -73311
rect -10517 -73711 -10317 -73311
rect -10259 -73711 -10059 -73311
rect -10001 -73711 -9801 -73311
rect -11291 -74571 -11091 -74171
rect -11033 -74571 -10833 -74171
rect -10775 -74571 -10575 -74171
rect -10517 -74571 -10317 -74171
rect -10259 -74571 -10059 -74171
rect -10001 -74571 -9801 -74171
rect -7291 -73711 -7091 -73311
rect -7033 -73711 -6833 -73311
rect -6775 -73711 -6575 -73311
rect -6517 -73711 -6317 -73311
rect -6259 -73711 -6059 -73311
rect -6001 -73711 -5801 -73311
rect -7291 -74571 -7091 -74171
rect -7033 -74571 -6833 -74171
rect -6775 -74571 -6575 -74171
rect -6517 -74571 -6317 -74171
rect -6259 -74571 -6059 -74171
rect -6001 -74571 -5801 -74171
rect -3291 -73711 -3091 -73311
rect -3033 -73711 -2833 -73311
rect -2775 -73711 -2575 -73311
rect -2517 -73711 -2317 -73311
rect -2259 -73711 -2059 -73311
rect -2001 -73711 -1801 -73311
rect -3291 -74571 -3091 -74171
rect -3033 -74571 -2833 -74171
rect -2775 -74571 -2575 -74171
rect -2517 -74571 -2317 -74171
rect -2259 -74571 -2059 -74171
rect -2001 -74571 -1801 -74171
rect 709 -73711 909 -73311
rect 967 -73711 1167 -73311
rect 1225 -73711 1425 -73311
rect 1483 -73711 1683 -73311
rect 1741 -73711 1941 -73311
rect 1999 -73711 2199 -73311
rect 709 -74571 909 -74171
rect 967 -74571 1167 -74171
rect 1225 -74571 1425 -74171
rect 1483 -74571 1683 -74171
rect 1741 -74571 1941 -74171
rect 1999 -74571 2199 -74171
rect 4709 -73711 4909 -73311
rect 4967 -73711 5167 -73311
rect 5225 -73711 5425 -73311
rect 5483 -73711 5683 -73311
rect 5741 -73711 5941 -73311
rect 5999 -73711 6199 -73311
rect 4709 -74571 4909 -74171
rect 4967 -74571 5167 -74171
rect 5225 -74571 5425 -74171
rect 5483 -74571 5683 -74171
rect 5741 -74571 5941 -74171
rect 5999 -74571 6199 -74171
<< nmoslvt >>
rect 16306 -45090 17266 -44490
rect 17324 -45090 18284 -44490
rect 18342 -45090 19302 -44490
rect 19360 -45090 20320 -44490
rect 20378 -45090 21338 -44490
rect 21396 -45090 22356 -44490
rect 22414 -45090 23374 -44490
rect 23432 -45090 24392 -44490
rect 24450 -45090 25410 -44490
rect 16306 -45908 17266 -45308
rect 17324 -45908 18284 -45308
rect 18342 -45908 19302 -45308
rect 19360 -45908 20320 -45308
rect 20378 -45908 21338 -45308
rect 21396 -45908 22356 -45308
rect 22414 -45908 23374 -45308
rect 23432 -45908 24392 -45308
rect 24450 -45908 25410 -45308
rect 16306 -46726 17266 -46126
rect 17324 -46726 18284 -46126
rect 18342 -46726 19302 -46126
rect 19360 -46726 20320 -46126
rect 20378 -46726 21338 -46126
rect 21396 -46726 22356 -46126
rect 22414 -46726 23374 -46126
rect 23432 -46726 24392 -46126
rect 24450 -46726 25410 -46126
rect 16306 -47544 17266 -46944
rect 17324 -47544 18284 -46944
rect 18342 -47544 19302 -46944
rect 19360 -47544 20320 -46944
rect 20378 -47544 21338 -46944
rect 21396 -47544 22356 -46944
rect 22414 -47544 23374 -46944
rect 23432 -47544 24392 -46944
rect 24450 -47544 25410 -46944
rect 16306 -48362 17266 -47762
rect 17324 -48362 18284 -47762
rect 18342 -48362 19302 -47762
rect 19360 -48362 20320 -47762
rect 20378 -48362 21338 -47762
rect 21396 -48362 22356 -47762
rect 22414 -48362 23374 -47762
rect 23432 -48362 24392 -47762
rect 24450 -48362 25410 -47762
rect 16306 -49180 17266 -48580
rect 17324 -49180 18284 -48580
rect 18342 -49180 19302 -48580
rect 19360 -49180 20320 -48580
rect 20378 -49180 21338 -48580
rect 21396 -49180 22356 -48580
rect 22414 -49180 23374 -48580
rect 23432 -49180 24392 -48580
rect 24450 -49180 25410 -48580
rect 16306 -49998 17266 -49398
rect 17324 -49998 18284 -49398
rect 18342 -49998 19302 -49398
rect 19360 -49998 20320 -49398
rect 20378 -49998 21338 -49398
rect 21396 -49998 22356 -49398
rect 22414 -49998 23374 -49398
rect 23432 -49998 24392 -49398
rect 24450 -49998 25410 -49398
rect 16306 -50816 17266 -50216
rect 17324 -50816 18284 -50216
rect 18342 -50816 19302 -50216
rect 19360 -50816 20320 -50216
rect 20378 -50816 21338 -50216
rect 21396 -50816 22356 -50216
rect 22414 -50816 23374 -50216
rect 23432 -50816 24392 -50216
rect 24450 -50816 25410 -50216
rect 14982 -52840 15942 -52240
rect 16000 -52840 16960 -52240
rect 17018 -52840 17978 -52240
rect 18036 -52840 18996 -52240
rect 19054 -52840 20014 -52240
rect 20072 -52840 21032 -52240
rect 21090 -52840 22050 -52240
rect 22108 -52840 23068 -52240
rect 23126 -52840 24086 -52240
rect 24144 -52840 25104 -52240
rect 25162 -52840 26122 -52240
rect 14982 -53952 15942 -53352
rect 16000 -53952 16960 -53352
rect 17018 -53952 17978 -53352
rect 18036 -53952 18996 -53352
rect 19054 -53952 20014 -53352
rect 20072 -53952 21032 -53352
rect 21090 -53952 22050 -53352
rect 22108 -53952 23068 -53352
rect 23126 -53952 24086 -53352
rect 24144 -53952 25104 -53352
rect 25162 -53952 26122 -53352
rect 14982 -55064 15942 -54464
rect 16000 -55064 16960 -54464
rect 17018 -55064 17978 -54464
rect 18036 -55064 18996 -54464
rect 19054 -55064 20014 -54464
rect 20072 -55064 21032 -54464
rect 21090 -55064 22050 -54464
rect 22108 -55064 23068 -54464
rect 23126 -55064 24086 -54464
rect 24144 -55064 25104 -54464
rect 25162 -55064 26122 -54464
rect 14982 -56176 15942 -55576
rect 16000 -56176 16960 -55576
rect 17018 -56176 17978 -55576
rect 18036 -56176 18996 -55576
rect 19054 -56176 20014 -55576
rect 20072 -56176 21032 -55576
rect 21090 -56176 22050 -55576
rect 22108 -56176 23068 -55576
rect 23126 -56176 24086 -55576
rect 24144 -56176 25104 -55576
rect 25162 -56176 26122 -55576
<< ndiff >>
rect 56172 -41971 56224 -41959
rect 56172 -42005 56180 -41971
rect 56214 -42005 56224 -41971
rect 56172 -42039 56224 -42005
rect 56172 -42073 56180 -42039
rect 56214 -42073 56224 -42039
rect 56172 -42089 56224 -42073
rect 56254 -41971 56306 -41959
rect 56254 -42005 56264 -41971
rect 56298 -42005 56306 -41971
rect 56254 -42039 56306 -42005
rect 56254 -42073 56264 -42039
rect 56298 -42073 56306 -42039
rect 56254 -42089 56306 -42073
rect 56448 -41971 56500 -41959
rect 56448 -42005 56456 -41971
rect 56490 -42005 56500 -41971
rect 56448 -42039 56500 -42005
rect 56448 -42073 56456 -42039
rect 56490 -42073 56500 -42039
rect 56448 -42089 56500 -42073
rect 56530 -41971 56582 -41959
rect 56530 -42005 56540 -41971
rect 56574 -42005 56582 -41971
rect 56530 -42039 56582 -42005
rect 56530 -42073 56540 -42039
rect 56574 -42073 56582 -42039
rect 56530 -42089 56582 -42073
rect 56687 -41975 56739 -41959
rect 56687 -42009 56695 -41975
rect 56729 -42009 56739 -41975
rect 56687 -42043 56739 -42009
rect 56687 -42077 56695 -42043
rect 56729 -42077 56739 -42043
rect 56687 -42089 56739 -42077
rect 56769 -42089 56823 -41959
rect 56853 -41975 56905 -41959
rect 56853 -42009 56863 -41975
rect 56897 -42009 56905 -41975
rect 56853 -42043 56905 -42009
rect 56853 -42077 56863 -42043
rect 56897 -42077 56905 -42043
rect 56853 -42089 56905 -42077
rect 57145 -41975 57197 -41959
rect 57145 -42009 57153 -41975
rect 57187 -42009 57197 -41975
rect 57145 -42043 57197 -42009
rect 57145 -42077 57153 -42043
rect 57187 -42077 57197 -42043
rect 57145 -42089 57197 -42077
rect 57227 -42089 57281 -41959
rect 57311 -41975 57363 -41959
rect 57311 -42009 57321 -41975
rect 57355 -42009 57363 -41975
rect 57311 -42043 57363 -42009
rect 57311 -42077 57321 -42043
rect 57355 -42077 57363 -42043
rect 57311 -42089 57363 -42077
rect 57468 -41971 57520 -41959
rect 57468 -42005 57476 -41971
rect 57510 -42005 57520 -41971
rect 57468 -42039 57520 -42005
rect 57468 -42073 57476 -42039
rect 57510 -42073 57520 -42039
rect 57468 -42089 57520 -42073
rect 57550 -41971 57602 -41959
rect 57550 -42005 57560 -41971
rect 57594 -42005 57602 -41971
rect 57550 -42039 57602 -42005
rect 57550 -42073 57560 -42039
rect 57594 -42073 57602 -42039
rect 57550 -42089 57602 -42073
rect 57744 -41971 57796 -41959
rect 57744 -42005 57752 -41971
rect 57786 -42005 57796 -41971
rect 57744 -42039 57796 -42005
rect 57744 -42073 57752 -42039
rect 57786 -42073 57796 -42039
rect 57744 -42089 57796 -42073
rect 57826 -41971 57878 -41959
rect 57826 -42005 57836 -41971
rect 57870 -42005 57878 -41971
rect 57826 -42039 57878 -42005
rect 57826 -42073 57836 -42039
rect 57870 -42073 57878 -42039
rect 57826 -42089 57878 -42073
rect 56004 -42714 56062 -42702
rect 56004 -42890 56016 -42714
rect 56050 -42890 56062 -42714
rect 56004 -42902 56062 -42890
rect 56122 -42714 56180 -42702
rect 56122 -42890 56134 -42714
rect 56168 -42890 56180 -42714
rect 56122 -42902 56180 -42890
rect 56550 -42628 56608 -42616
rect 56550 -42804 56562 -42628
rect 56596 -42804 56608 -42628
rect 56550 -42816 56608 -42804
rect 56668 -42628 56726 -42616
rect 56668 -42804 56680 -42628
rect 56714 -42804 56726 -42628
rect 56668 -42816 56726 -42804
rect 56786 -42628 56844 -42616
rect 56786 -42804 56798 -42628
rect 56832 -42804 56844 -42628
rect 56786 -42816 56844 -42804
rect 56904 -42628 56962 -42616
rect 56904 -42804 56916 -42628
rect 56950 -42804 56962 -42628
rect 56904 -42816 56962 -42804
rect 57022 -42628 57080 -42616
rect 57022 -42804 57034 -42628
rect 57068 -42804 57080 -42628
rect 57022 -42816 57080 -42804
rect 57140 -42628 57198 -42616
rect 57140 -42804 57152 -42628
rect 57186 -42804 57198 -42628
rect 57140 -42816 57198 -42804
rect 57258 -42628 57316 -42616
rect 57258 -42804 57270 -42628
rect 57304 -42804 57316 -42628
rect 57258 -42816 57316 -42804
rect 57376 -42628 57434 -42616
rect 57376 -42804 57388 -42628
rect 57422 -42804 57434 -42628
rect 57376 -42816 57434 -42804
rect 57494 -42628 57552 -42616
rect 57494 -42804 57506 -42628
rect 57540 -42804 57552 -42628
rect 57494 -42816 57552 -42804
rect 12254 -57637 12306 -57625
rect 12254 -57671 12262 -57637
rect 12296 -57671 12306 -57637
rect 12254 -57705 12306 -57671
rect 12254 -57739 12262 -57705
rect 12296 -57739 12306 -57705
rect 12254 -57755 12306 -57739
rect 12336 -57637 12388 -57625
rect 12336 -57671 12346 -57637
rect 12380 -57671 12388 -57637
rect 12336 -57705 12388 -57671
rect 12336 -57739 12346 -57705
rect 12380 -57739 12388 -57705
rect 12336 -57755 12388 -57739
rect 10398 -57858 10456 -57846
rect 10398 -58034 10410 -57858
rect 10444 -58034 10456 -57858
rect 10398 -58046 10456 -58034
rect 10656 -57858 10714 -57846
rect 10656 -58034 10668 -57858
rect 10702 -58034 10714 -57858
rect 10656 -58046 10714 -58034
rect 10914 -57858 10972 -57846
rect 10914 -58034 10926 -57858
rect 10960 -58034 10972 -57858
rect 10914 -58046 10972 -58034
rect 11172 -57858 11230 -57846
rect 11172 -58034 11184 -57858
rect 11218 -58034 11230 -57858
rect 11172 -58046 11230 -58034
rect 11430 -57858 11488 -57846
rect 11430 -58034 11442 -57858
rect 11476 -58034 11488 -57858
rect 11430 -58046 11488 -58034
rect 11688 -57858 11746 -57846
rect 11688 -58034 11700 -57858
rect 11734 -58034 11746 -57858
rect 11688 -58046 11746 -58034
rect 11946 -57858 12004 -57846
rect 11946 -58034 11958 -57858
rect 11992 -58034 12004 -57858
rect 11946 -58046 12004 -58034
rect 28014 -44026 28072 -44014
rect 16248 -44502 16306 -44490
rect 16248 -45078 16260 -44502
rect 16294 -45078 16306 -44502
rect 16248 -45090 16306 -45078
rect 17266 -44502 17324 -44490
rect 17266 -45078 17278 -44502
rect 17312 -45078 17324 -44502
rect 17266 -45090 17324 -45078
rect 18284 -44502 18342 -44490
rect 18284 -45078 18296 -44502
rect 18330 -45078 18342 -44502
rect 18284 -45090 18342 -45078
rect 19302 -44502 19360 -44490
rect 19302 -45078 19314 -44502
rect 19348 -45078 19360 -44502
rect 19302 -45090 19360 -45078
rect 20320 -44502 20378 -44490
rect 20320 -45078 20332 -44502
rect 20366 -45078 20378 -44502
rect 20320 -45090 20378 -45078
rect 21338 -44502 21396 -44490
rect 21338 -45078 21350 -44502
rect 21384 -45078 21396 -44502
rect 21338 -45090 21396 -45078
rect 22356 -44502 22414 -44490
rect 22356 -45078 22368 -44502
rect 22402 -45078 22414 -44502
rect 22356 -45090 22414 -45078
rect 23374 -44502 23432 -44490
rect 23374 -45078 23386 -44502
rect 23420 -45078 23432 -44502
rect 23374 -45090 23432 -45078
rect 24392 -44502 24450 -44490
rect 24392 -45078 24404 -44502
rect 24438 -45078 24450 -44502
rect 24392 -45090 24450 -45078
rect 25410 -44502 25468 -44490
rect 25410 -45078 25422 -44502
rect 25456 -45078 25468 -44502
rect 28014 -44602 28026 -44026
rect 28060 -44602 28072 -44026
rect 28014 -44614 28072 -44602
rect 29032 -44026 29090 -44014
rect 29032 -44602 29044 -44026
rect 29078 -44602 29090 -44026
rect 29032 -44614 29090 -44602
rect 30050 -44026 30108 -44014
rect 30050 -44602 30062 -44026
rect 30096 -44602 30108 -44026
rect 30050 -44614 30108 -44602
rect 31068 -44026 31126 -44014
rect 31068 -44602 31080 -44026
rect 31114 -44602 31126 -44026
rect 31068 -44614 31126 -44602
rect 32086 -44026 32144 -44014
rect 32086 -44602 32098 -44026
rect 32132 -44602 32144 -44026
rect 32086 -44614 32144 -44602
rect 33104 -44026 33162 -44014
rect 33104 -44602 33116 -44026
rect 33150 -44602 33162 -44026
rect 33104 -44614 33162 -44602
rect 34122 -44026 34180 -44014
rect 34122 -44602 34134 -44026
rect 34168 -44602 34180 -44026
rect 34122 -44614 34180 -44602
rect 35140 -44026 35198 -44014
rect 35140 -44602 35152 -44026
rect 35186 -44602 35198 -44026
rect 35140 -44614 35198 -44602
rect 36158 -44026 36216 -44014
rect 36158 -44602 36170 -44026
rect 36204 -44602 36216 -44026
rect 36158 -44614 36216 -44602
rect 37176 -44026 37234 -44014
rect 37176 -44602 37188 -44026
rect 37222 -44602 37234 -44026
rect 37176 -44614 37234 -44602
rect 38194 -44026 38252 -44014
rect 38194 -44602 38206 -44026
rect 38240 -44602 38252 -44026
rect 38194 -44614 38252 -44602
rect 39212 -44026 39270 -44014
rect 39212 -44602 39224 -44026
rect 39258 -44602 39270 -44026
rect 39212 -44614 39270 -44602
rect 40230 -44026 40288 -44014
rect 40230 -44602 40242 -44026
rect 40276 -44602 40288 -44026
rect 40230 -44614 40288 -44602
rect 41248 -44026 41306 -44014
rect 41248 -44602 41260 -44026
rect 41294 -44602 41306 -44026
rect 41248 -44614 41306 -44602
rect 42266 -44026 42324 -44014
rect 42266 -44602 42278 -44026
rect 42312 -44602 42324 -44026
rect 42266 -44614 42324 -44602
rect 43284 -44026 43342 -44014
rect 43284 -44602 43296 -44026
rect 43330 -44602 43342 -44026
rect 43284 -44614 43342 -44602
rect 44302 -44026 44360 -44014
rect 44302 -44602 44314 -44026
rect 44348 -44602 44360 -44026
rect 44302 -44614 44360 -44602
rect 45320 -44026 45378 -44014
rect 45320 -44602 45332 -44026
rect 45366 -44602 45378 -44026
rect 45320 -44614 45378 -44602
rect 46338 -44026 46396 -44014
rect 46338 -44602 46350 -44026
rect 46384 -44602 46396 -44026
rect 46338 -44614 46396 -44602
rect 47356 -44026 47414 -44014
rect 47356 -44602 47368 -44026
rect 47402 -44602 47414 -44026
rect 47356 -44614 47414 -44602
rect 48374 -44026 48432 -44014
rect 48374 -44602 48386 -44026
rect 48420 -44602 48432 -44026
rect 48374 -44614 48432 -44602
rect 25410 -45090 25468 -45078
rect 28014 -44844 28072 -44832
rect 16248 -45320 16306 -45308
rect 16248 -45896 16260 -45320
rect 16294 -45896 16306 -45320
rect 16248 -45908 16306 -45896
rect 17266 -45320 17324 -45308
rect 17266 -45896 17278 -45320
rect 17312 -45896 17324 -45320
rect 17266 -45908 17324 -45896
rect 18284 -45320 18342 -45308
rect 18284 -45896 18296 -45320
rect 18330 -45896 18342 -45320
rect 18284 -45908 18342 -45896
rect 19302 -45320 19360 -45308
rect 19302 -45896 19314 -45320
rect 19348 -45896 19360 -45320
rect 19302 -45908 19360 -45896
rect 20320 -45320 20378 -45308
rect 20320 -45896 20332 -45320
rect 20366 -45896 20378 -45320
rect 20320 -45908 20378 -45896
rect 21338 -45320 21396 -45308
rect 21338 -45896 21350 -45320
rect 21384 -45896 21396 -45320
rect 21338 -45908 21396 -45896
rect 22356 -45320 22414 -45308
rect 22356 -45896 22368 -45320
rect 22402 -45896 22414 -45320
rect 22356 -45908 22414 -45896
rect 23374 -45320 23432 -45308
rect 23374 -45896 23386 -45320
rect 23420 -45896 23432 -45320
rect 23374 -45908 23432 -45896
rect 24392 -45320 24450 -45308
rect 24392 -45896 24404 -45320
rect 24438 -45896 24450 -45320
rect 24392 -45908 24450 -45896
rect 25410 -45320 25468 -45308
rect 25410 -45896 25422 -45320
rect 25456 -45896 25468 -45320
rect 28014 -45420 28026 -44844
rect 28060 -45420 28072 -44844
rect 28014 -45432 28072 -45420
rect 29032 -44844 29090 -44832
rect 29032 -45420 29044 -44844
rect 29078 -45420 29090 -44844
rect 29032 -45432 29090 -45420
rect 30050 -44844 30108 -44832
rect 30050 -45420 30062 -44844
rect 30096 -45420 30108 -44844
rect 30050 -45432 30108 -45420
rect 31068 -44844 31126 -44832
rect 31068 -45420 31080 -44844
rect 31114 -45420 31126 -44844
rect 31068 -45432 31126 -45420
rect 32086 -44844 32144 -44832
rect 32086 -45420 32098 -44844
rect 32132 -45420 32144 -44844
rect 32086 -45432 32144 -45420
rect 33104 -44844 33162 -44832
rect 33104 -45420 33116 -44844
rect 33150 -45420 33162 -44844
rect 33104 -45432 33162 -45420
rect 34122 -44844 34180 -44832
rect 34122 -45420 34134 -44844
rect 34168 -45420 34180 -44844
rect 34122 -45432 34180 -45420
rect 35140 -44844 35198 -44832
rect 35140 -45420 35152 -44844
rect 35186 -45420 35198 -44844
rect 35140 -45432 35198 -45420
rect 36158 -44844 36216 -44832
rect 36158 -45420 36170 -44844
rect 36204 -45420 36216 -44844
rect 36158 -45432 36216 -45420
rect 37176 -44844 37234 -44832
rect 37176 -45420 37188 -44844
rect 37222 -45420 37234 -44844
rect 37176 -45432 37234 -45420
rect 38194 -44844 38252 -44832
rect 38194 -45420 38206 -44844
rect 38240 -45420 38252 -44844
rect 38194 -45432 38252 -45420
rect 39212 -44844 39270 -44832
rect 39212 -45420 39224 -44844
rect 39258 -45420 39270 -44844
rect 39212 -45432 39270 -45420
rect 40230 -44844 40288 -44832
rect 40230 -45420 40242 -44844
rect 40276 -45420 40288 -44844
rect 40230 -45432 40288 -45420
rect 41248 -44844 41306 -44832
rect 41248 -45420 41260 -44844
rect 41294 -45420 41306 -44844
rect 41248 -45432 41306 -45420
rect 42266 -44844 42324 -44832
rect 42266 -45420 42278 -44844
rect 42312 -45420 42324 -44844
rect 42266 -45432 42324 -45420
rect 43284 -44844 43342 -44832
rect 43284 -45420 43296 -44844
rect 43330 -45420 43342 -44844
rect 43284 -45432 43342 -45420
rect 44302 -44844 44360 -44832
rect 44302 -45420 44314 -44844
rect 44348 -45420 44360 -44844
rect 44302 -45432 44360 -45420
rect 45320 -44844 45378 -44832
rect 45320 -45420 45332 -44844
rect 45366 -45420 45378 -44844
rect 45320 -45432 45378 -45420
rect 46338 -44844 46396 -44832
rect 46338 -45420 46350 -44844
rect 46384 -45420 46396 -44844
rect 46338 -45432 46396 -45420
rect 47356 -44844 47414 -44832
rect 47356 -45420 47368 -44844
rect 47402 -45420 47414 -44844
rect 47356 -45432 47414 -45420
rect 48374 -44844 48432 -44832
rect 48374 -45420 48386 -44844
rect 48420 -45420 48432 -44844
rect 48374 -45432 48432 -45420
rect 25410 -45908 25468 -45896
rect 16248 -46138 16306 -46126
rect 16248 -46714 16260 -46138
rect 16294 -46714 16306 -46138
rect 16248 -46726 16306 -46714
rect 17266 -46138 17324 -46126
rect 17266 -46714 17278 -46138
rect 17312 -46714 17324 -46138
rect 17266 -46726 17324 -46714
rect 18284 -46138 18342 -46126
rect 18284 -46714 18296 -46138
rect 18330 -46714 18342 -46138
rect 18284 -46726 18342 -46714
rect 19302 -46138 19360 -46126
rect 19302 -46714 19314 -46138
rect 19348 -46714 19360 -46138
rect 19302 -46726 19360 -46714
rect 20320 -46138 20378 -46126
rect 20320 -46714 20332 -46138
rect 20366 -46714 20378 -46138
rect 20320 -46726 20378 -46714
rect 21338 -46138 21396 -46126
rect 21338 -46714 21350 -46138
rect 21384 -46714 21396 -46138
rect 21338 -46726 21396 -46714
rect 22356 -46138 22414 -46126
rect 22356 -46714 22368 -46138
rect 22402 -46714 22414 -46138
rect 22356 -46726 22414 -46714
rect 23374 -46138 23432 -46126
rect 23374 -46714 23386 -46138
rect 23420 -46714 23432 -46138
rect 23374 -46726 23432 -46714
rect 24392 -46138 24450 -46126
rect 24392 -46714 24404 -46138
rect 24438 -46714 24450 -46138
rect 24392 -46726 24450 -46714
rect 25410 -46138 25468 -46126
rect 25410 -46714 25422 -46138
rect 25456 -46714 25468 -46138
rect 25410 -46726 25468 -46714
rect 28014 -46222 28072 -46210
rect 28014 -46798 28026 -46222
rect 28060 -46798 28072 -46222
rect 28014 -46810 28072 -46798
rect 29032 -46222 29090 -46210
rect 29032 -46798 29044 -46222
rect 29078 -46798 29090 -46222
rect 29032 -46810 29090 -46798
rect 30050 -46222 30108 -46210
rect 30050 -46798 30062 -46222
rect 30096 -46798 30108 -46222
rect 30050 -46810 30108 -46798
rect 31068 -46222 31126 -46210
rect 31068 -46798 31080 -46222
rect 31114 -46798 31126 -46222
rect 31068 -46810 31126 -46798
rect 32086 -46222 32144 -46210
rect 32086 -46798 32098 -46222
rect 32132 -46798 32144 -46222
rect 32086 -46810 32144 -46798
rect 33104 -46222 33162 -46210
rect 33104 -46798 33116 -46222
rect 33150 -46798 33162 -46222
rect 33104 -46810 33162 -46798
rect 34122 -46222 34180 -46210
rect 34122 -46798 34134 -46222
rect 34168 -46798 34180 -46222
rect 34122 -46810 34180 -46798
rect 35140 -46222 35198 -46210
rect 35140 -46798 35152 -46222
rect 35186 -46798 35198 -46222
rect 35140 -46810 35198 -46798
rect 36158 -46222 36216 -46210
rect 36158 -46798 36170 -46222
rect 36204 -46798 36216 -46222
rect 36158 -46810 36216 -46798
rect 37176 -46222 37234 -46210
rect 37176 -46798 37188 -46222
rect 37222 -46798 37234 -46222
rect 37176 -46810 37234 -46798
rect 38194 -46222 38252 -46210
rect 38194 -46798 38206 -46222
rect 38240 -46798 38252 -46222
rect 38194 -46810 38252 -46798
rect 39212 -46222 39270 -46210
rect 39212 -46798 39224 -46222
rect 39258 -46798 39270 -46222
rect 39212 -46810 39270 -46798
rect 40230 -46222 40288 -46210
rect 40230 -46798 40242 -46222
rect 40276 -46798 40288 -46222
rect 40230 -46810 40288 -46798
rect 41248 -46222 41306 -46210
rect 41248 -46798 41260 -46222
rect 41294 -46798 41306 -46222
rect 41248 -46810 41306 -46798
rect 42266 -46222 42324 -46210
rect 42266 -46798 42278 -46222
rect 42312 -46798 42324 -46222
rect 42266 -46810 42324 -46798
rect 43284 -46222 43342 -46210
rect 43284 -46798 43296 -46222
rect 43330 -46798 43342 -46222
rect 43284 -46810 43342 -46798
rect 44302 -46222 44360 -46210
rect 44302 -46798 44314 -46222
rect 44348 -46798 44360 -46222
rect 44302 -46810 44360 -46798
rect 45320 -46222 45378 -46210
rect 45320 -46798 45332 -46222
rect 45366 -46798 45378 -46222
rect 45320 -46810 45378 -46798
rect 46338 -46222 46396 -46210
rect 46338 -46798 46350 -46222
rect 46384 -46798 46396 -46222
rect 46338 -46810 46396 -46798
rect 47356 -46222 47414 -46210
rect 47356 -46798 47368 -46222
rect 47402 -46798 47414 -46222
rect 47356 -46810 47414 -46798
rect 48374 -46222 48432 -46210
rect 48374 -46798 48386 -46222
rect 48420 -46798 48432 -46222
rect 48374 -46810 48432 -46798
rect 16248 -46956 16306 -46944
rect 16248 -47532 16260 -46956
rect 16294 -47532 16306 -46956
rect 16248 -47544 16306 -47532
rect 17266 -46956 17324 -46944
rect 17266 -47532 17278 -46956
rect 17312 -47532 17324 -46956
rect 17266 -47544 17324 -47532
rect 18284 -46956 18342 -46944
rect 18284 -47532 18296 -46956
rect 18330 -47532 18342 -46956
rect 18284 -47544 18342 -47532
rect 19302 -46956 19360 -46944
rect 19302 -47532 19314 -46956
rect 19348 -47532 19360 -46956
rect 19302 -47544 19360 -47532
rect 20320 -46956 20378 -46944
rect 20320 -47532 20332 -46956
rect 20366 -47532 20378 -46956
rect 20320 -47544 20378 -47532
rect 21338 -46956 21396 -46944
rect 21338 -47532 21350 -46956
rect 21384 -47532 21396 -46956
rect 21338 -47544 21396 -47532
rect 22356 -46956 22414 -46944
rect 22356 -47532 22368 -46956
rect 22402 -47532 22414 -46956
rect 22356 -47544 22414 -47532
rect 23374 -46956 23432 -46944
rect 23374 -47532 23386 -46956
rect 23420 -47532 23432 -46956
rect 23374 -47544 23432 -47532
rect 24392 -46956 24450 -46944
rect 24392 -47532 24404 -46956
rect 24438 -47532 24450 -46956
rect 24392 -47544 24450 -47532
rect 25410 -46956 25468 -46944
rect 25410 -47532 25422 -46956
rect 25456 -47532 25468 -46956
rect 25410 -47544 25468 -47532
rect 28014 -47454 28072 -47442
rect 16248 -47774 16306 -47762
rect 16248 -48350 16260 -47774
rect 16294 -48350 16306 -47774
rect 16248 -48362 16306 -48350
rect 17266 -47774 17324 -47762
rect 17266 -48350 17278 -47774
rect 17312 -48350 17324 -47774
rect 17266 -48362 17324 -48350
rect 18284 -47774 18342 -47762
rect 18284 -48350 18296 -47774
rect 18330 -48350 18342 -47774
rect 18284 -48362 18342 -48350
rect 19302 -47774 19360 -47762
rect 19302 -48350 19314 -47774
rect 19348 -48350 19360 -47774
rect 19302 -48362 19360 -48350
rect 20320 -47774 20378 -47762
rect 20320 -48350 20332 -47774
rect 20366 -48350 20378 -47774
rect 20320 -48362 20378 -48350
rect 21338 -47774 21396 -47762
rect 21338 -48350 21350 -47774
rect 21384 -48350 21396 -47774
rect 21338 -48362 21396 -48350
rect 22356 -47774 22414 -47762
rect 22356 -48350 22368 -47774
rect 22402 -48350 22414 -47774
rect 22356 -48362 22414 -48350
rect 23374 -47774 23432 -47762
rect 23374 -48350 23386 -47774
rect 23420 -48350 23432 -47774
rect 23374 -48362 23432 -48350
rect 24392 -47774 24450 -47762
rect 24392 -48350 24404 -47774
rect 24438 -48350 24450 -47774
rect 24392 -48362 24450 -48350
rect 25410 -47774 25468 -47762
rect 25410 -48350 25422 -47774
rect 25456 -48350 25468 -47774
rect 28014 -48030 28026 -47454
rect 28060 -48030 28072 -47454
rect 28014 -48042 28072 -48030
rect 29032 -47454 29090 -47442
rect 29032 -48030 29044 -47454
rect 29078 -48030 29090 -47454
rect 29032 -48042 29090 -48030
rect 30050 -47454 30108 -47442
rect 30050 -48030 30062 -47454
rect 30096 -48030 30108 -47454
rect 30050 -48042 30108 -48030
rect 31068 -47454 31126 -47442
rect 31068 -48030 31080 -47454
rect 31114 -48030 31126 -47454
rect 31068 -48042 31126 -48030
rect 32086 -47454 32144 -47442
rect 32086 -48030 32098 -47454
rect 32132 -48030 32144 -47454
rect 32086 -48042 32144 -48030
rect 33104 -47454 33162 -47442
rect 33104 -48030 33116 -47454
rect 33150 -48030 33162 -47454
rect 33104 -48042 33162 -48030
rect 34122 -47454 34180 -47442
rect 34122 -48030 34134 -47454
rect 34168 -48030 34180 -47454
rect 34122 -48042 34180 -48030
rect 35140 -47454 35198 -47442
rect 35140 -48030 35152 -47454
rect 35186 -48030 35198 -47454
rect 35140 -48042 35198 -48030
rect 36158 -47454 36216 -47442
rect 36158 -48030 36170 -47454
rect 36204 -48030 36216 -47454
rect 36158 -48042 36216 -48030
rect 37176 -47454 37234 -47442
rect 37176 -48030 37188 -47454
rect 37222 -48030 37234 -47454
rect 37176 -48042 37234 -48030
rect 38194 -47454 38252 -47442
rect 38194 -48030 38206 -47454
rect 38240 -48030 38252 -47454
rect 38194 -48042 38252 -48030
rect 39212 -47454 39270 -47442
rect 39212 -48030 39224 -47454
rect 39258 -48030 39270 -47454
rect 39212 -48042 39270 -48030
rect 40230 -47454 40288 -47442
rect 40230 -48030 40242 -47454
rect 40276 -48030 40288 -47454
rect 40230 -48042 40288 -48030
rect 41248 -47454 41306 -47442
rect 41248 -48030 41260 -47454
rect 41294 -48030 41306 -47454
rect 41248 -48042 41306 -48030
rect 42266 -47454 42324 -47442
rect 42266 -48030 42278 -47454
rect 42312 -48030 42324 -47454
rect 42266 -48042 42324 -48030
rect 43284 -47454 43342 -47442
rect 43284 -48030 43296 -47454
rect 43330 -48030 43342 -47454
rect 43284 -48042 43342 -48030
rect 44302 -47454 44360 -47442
rect 44302 -48030 44314 -47454
rect 44348 -48030 44360 -47454
rect 44302 -48042 44360 -48030
rect 45320 -47454 45378 -47442
rect 45320 -48030 45332 -47454
rect 45366 -48030 45378 -47454
rect 45320 -48042 45378 -48030
rect 46338 -47454 46396 -47442
rect 46338 -48030 46350 -47454
rect 46384 -48030 46396 -47454
rect 46338 -48042 46396 -48030
rect 47356 -47454 47414 -47442
rect 47356 -48030 47368 -47454
rect 47402 -48030 47414 -47454
rect 47356 -48042 47414 -48030
rect 48374 -47454 48432 -47442
rect 48374 -48030 48386 -47454
rect 48420 -48030 48432 -47454
rect 48374 -48042 48432 -48030
rect 25410 -48362 25468 -48350
rect 16248 -48592 16306 -48580
rect 16248 -49168 16260 -48592
rect 16294 -49168 16306 -48592
rect 16248 -49180 16306 -49168
rect 17266 -48592 17324 -48580
rect 17266 -49168 17278 -48592
rect 17312 -49168 17324 -48592
rect 17266 -49180 17324 -49168
rect 18284 -48592 18342 -48580
rect 18284 -49168 18296 -48592
rect 18330 -49168 18342 -48592
rect 18284 -49180 18342 -49168
rect 19302 -48592 19360 -48580
rect 19302 -49168 19314 -48592
rect 19348 -49168 19360 -48592
rect 19302 -49180 19360 -49168
rect 20320 -48592 20378 -48580
rect 20320 -49168 20332 -48592
rect 20366 -49168 20378 -48592
rect 20320 -49180 20378 -49168
rect 21338 -48592 21396 -48580
rect 21338 -49168 21350 -48592
rect 21384 -49168 21396 -48592
rect 21338 -49180 21396 -49168
rect 22356 -48592 22414 -48580
rect 22356 -49168 22368 -48592
rect 22402 -49168 22414 -48592
rect 22356 -49180 22414 -49168
rect 23374 -48592 23432 -48580
rect 23374 -49168 23386 -48592
rect 23420 -49168 23432 -48592
rect 23374 -49180 23432 -49168
rect 24392 -48592 24450 -48580
rect 24392 -49168 24404 -48592
rect 24438 -49168 24450 -48592
rect 24392 -49180 24450 -49168
rect 25410 -48592 25468 -48580
rect 25410 -49168 25422 -48592
rect 25456 -49168 25468 -48592
rect 25410 -49180 25468 -49168
rect 28012 -48688 28070 -48676
rect 28012 -49264 28024 -48688
rect 28058 -49264 28070 -48688
rect 28012 -49276 28070 -49264
rect 29030 -48688 29088 -48676
rect 29030 -49264 29042 -48688
rect 29076 -49264 29088 -48688
rect 29030 -49276 29088 -49264
rect 30048 -48688 30106 -48676
rect 30048 -49264 30060 -48688
rect 30094 -49264 30106 -48688
rect 30048 -49276 30106 -49264
rect 31066 -48688 31124 -48676
rect 31066 -49264 31078 -48688
rect 31112 -49264 31124 -48688
rect 31066 -49276 31124 -49264
rect 32084 -48688 32142 -48676
rect 32084 -49264 32096 -48688
rect 32130 -49264 32142 -48688
rect 32084 -49276 32142 -49264
rect 33102 -48688 33160 -48676
rect 33102 -49264 33114 -48688
rect 33148 -49264 33160 -48688
rect 33102 -49276 33160 -49264
rect 34120 -48688 34178 -48676
rect 34120 -49264 34132 -48688
rect 34166 -49264 34178 -48688
rect 34120 -49276 34178 -49264
rect 35138 -48688 35196 -48676
rect 35138 -49264 35150 -48688
rect 35184 -49264 35196 -48688
rect 35138 -49276 35196 -49264
rect 36156 -48688 36214 -48676
rect 36156 -49264 36168 -48688
rect 36202 -49264 36214 -48688
rect 36156 -49276 36214 -49264
rect 37174 -48688 37232 -48676
rect 37174 -49264 37186 -48688
rect 37220 -49264 37232 -48688
rect 37174 -49276 37232 -49264
rect 38192 -48688 38250 -48676
rect 38192 -49264 38204 -48688
rect 38238 -49264 38250 -48688
rect 38192 -49276 38250 -49264
rect 39210 -48688 39268 -48676
rect 39210 -49264 39222 -48688
rect 39256 -49264 39268 -48688
rect 39210 -49276 39268 -49264
rect 40228 -48688 40286 -48676
rect 40228 -49264 40240 -48688
rect 40274 -49264 40286 -48688
rect 40228 -49276 40286 -49264
rect 41246 -48688 41304 -48676
rect 41246 -49264 41258 -48688
rect 41292 -49264 41304 -48688
rect 41246 -49276 41304 -49264
rect 42264 -48688 42322 -48676
rect 42264 -49264 42276 -48688
rect 42310 -49264 42322 -48688
rect 42264 -49276 42322 -49264
rect 43282 -48688 43340 -48676
rect 43282 -49264 43294 -48688
rect 43328 -49264 43340 -48688
rect 43282 -49276 43340 -49264
rect 44300 -48688 44358 -48676
rect 44300 -49264 44312 -48688
rect 44346 -49264 44358 -48688
rect 44300 -49276 44358 -49264
rect 45318 -48688 45376 -48676
rect 45318 -49264 45330 -48688
rect 45364 -49264 45376 -48688
rect 45318 -49276 45376 -49264
rect 46336 -48688 46394 -48676
rect 46336 -49264 46348 -48688
rect 46382 -49264 46394 -48688
rect 46336 -49276 46394 -49264
rect 47354 -48688 47412 -48676
rect 47354 -49264 47366 -48688
rect 47400 -49264 47412 -48688
rect 47354 -49276 47412 -49264
rect 48372 -48688 48430 -48676
rect 48372 -49264 48384 -48688
rect 48418 -49264 48430 -48688
rect 48372 -49276 48430 -49264
rect 16248 -49410 16306 -49398
rect 16248 -49986 16260 -49410
rect 16294 -49986 16306 -49410
rect 16248 -49998 16306 -49986
rect 17266 -49410 17324 -49398
rect 17266 -49986 17278 -49410
rect 17312 -49986 17324 -49410
rect 17266 -49998 17324 -49986
rect 18284 -49410 18342 -49398
rect 18284 -49986 18296 -49410
rect 18330 -49986 18342 -49410
rect 18284 -49998 18342 -49986
rect 19302 -49410 19360 -49398
rect 19302 -49986 19314 -49410
rect 19348 -49986 19360 -49410
rect 19302 -49998 19360 -49986
rect 20320 -49410 20378 -49398
rect 20320 -49986 20332 -49410
rect 20366 -49986 20378 -49410
rect 20320 -49998 20378 -49986
rect 21338 -49410 21396 -49398
rect 21338 -49986 21350 -49410
rect 21384 -49986 21396 -49410
rect 21338 -49998 21396 -49986
rect 22356 -49410 22414 -49398
rect 22356 -49986 22368 -49410
rect 22402 -49986 22414 -49410
rect 22356 -49998 22414 -49986
rect 23374 -49410 23432 -49398
rect 23374 -49986 23386 -49410
rect 23420 -49986 23432 -49410
rect 23374 -49998 23432 -49986
rect 24392 -49410 24450 -49398
rect 24392 -49986 24404 -49410
rect 24438 -49986 24450 -49410
rect 24392 -49998 24450 -49986
rect 25410 -49410 25468 -49398
rect 25410 -49986 25422 -49410
rect 25456 -49986 25468 -49410
rect 25410 -49998 25468 -49986
rect 28012 -49922 28070 -49910
rect 16248 -50228 16306 -50216
rect 16248 -50804 16260 -50228
rect 16294 -50804 16306 -50228
rect 16248 -50816 16306 -50804
rect 17266 -50228 17324 -50216
rect 17266 -50804 17278 -50228
rect 17312 -50804 17324 -50228
rect 17266 -50816 17324 -50804
rect 18284 -50228 18342 -50216
rect 18284 -50804 18296 -50228
rect 18330 -50804 18342 -50228
rect 18284 -50816 18342 -50804
rect 19302 -50228 19360 -50216
rect 19302 -50804 19314 -50228
rect 19348 -50804 19360 -50228
rect 19302 -50816 19360 -50804
rect 20320 -50228 20378 -50216
rect 20320 -50804 20332 -50228
rect 20366 -50804 20378 -50228
rect 20320 -50816 20378 -50804
rect 21338 -50228 21396 -50216
rect 21338 -50804 21350 -50228
rect 21384 -50804 21396 -50228
rect 21338 -50816 21396 -50804
rect 22356 -50228 22414 -50216
rect 22356 -50804 22368 -50228
rect 22402 -50804 22414 -50228
rect 22356 -50816 22414 -50804
rect 23374 -50228 23432 -50216
rect 23374 -50804 23386 -50228
rect 23420 -50804 23432 -50228
rect 23374 -50816 23432 -50804
rect 24392 -50228 24450 -50216
rect 24392 -50804 24404 -50228
rect 24438 -50804 24450 -50228
rect 24392 -50816 24450 -50804
rect 25410 -50228 25468 -50216
rect 25410 -50804 25422 -50228
rect 25456 -50804 25468 -50228
rect 28012 -50498 28024 -49922
rect 28058 -50498 28070 -49922
rect 28012 -50510 28070 -50498
rect 29030 -49922 29088 -49910
rect 29030 -50498 29042 -49922
rect 29076 -50498 29088 -49922
rect 29030 -50510 29088 -50498
rect 30048 -49922 30106 -49910
rect 30048 -50498 30060 -49922
rect 30094 -50498 30106 -49922
rect 30048 -50510 30106 -50498
rect 31066 -49922 31124 -49910
rect 31066 -50498 31078 -49922
rect 31112 -50498 31124 -49922
rect 31066 -50510 31124 -50498
rect 32084 -49922 32142 -49910
rect 32084 -50498 32096 -49922
rect 32130 -50498 32142 -49922
rect 32084 -50510 32142 -50498
rect 33102 -49922 33160 -49910
rect 33102 -50498 33114 -49922
rect 33148 -50498 33160 -49922
rect 33102 -50510 33160 -50498
rect 34120 -49922 34178 -49910
rect 34120 -50498 34132 -49922
rect 34166 -50498 34178 -49922
rect 34120 -50510 34178 -50498
rect 35138 -49922 35196 -49910
rect 35138 -50498 35150 -49922
rect 35184 -50498 35196 -49922
rect 35138 -50510 35196 -50498
rect 36156 -49922 36214 -49910
rect 36156 -50498 36168 -49922
rect 36202 -50498 36214 -49922
rect 36156 -50510 36214 -50498
rect 37174 -49922 37232 -49910
rect 37174 -50498 37186 -49922
rect 37220 -50498 37232 -49922
rect 37174 -50510 37232 -50498
rect 38192 -49922 38250 -49910
rect 38192 -50498 38204 -49922
rect 38238 -50498 38250 -49922
rect 38192 -50510 38250 -50498
rect 39210 -49922 39268 -49910
rect 39210 -50498 39222 -49922
rect 39256 -50498 39268 -49922
rect 39210 -50510 39268 -50498
rect 40228 -49922 40286 -49910
rect 40228 -50498 40240 -49922
rect 40274 -50498 40286 -49922
rect 40228 -50510 40286 -50498
rect 41246 -49922 41304 -49910
rect 41246 -50498 41258 -49922
rect 41292 -50498 41304 -49922
rect 41246 -50510 41304 -50498
rect 42264 -49922 42322 -49910
rect 42264 -50498 42276 -49922
rect 42310 -50498 42322 -49922
rect 42264 -50510 42322 -50498
rect 43282 -49922 43340 -49910
rect 43282 -50498 43294 -49922
rect 43328 -50498 43340 -49922
rect 43282 -50510 43340 -50498
rect 44300 -49922 44358 -49910
rect 44300 -50498 44312 -49922
rect 44346 -50498 44358 -49922
rect 44300 -50510 44358 -50498
rect 45318 -49922 45376 -49910
rect 45318 -50498 45330 -49922
rect 45364 -50498 45376 -49922
rect 45318 -50510 45376 -50498
rect 46336 -49922 46394 -49910
rect 46336 -50498 46348 -49922
rect 46382 -50498 46394 -49922
rect 46336 -50510 46394 -50498
rect 47354 -49922 47412 -49910
rect 47354 -50498 47366 -49922
rect 47400 -50498 47412 -49922
rect 47354 -50510 47412 -50498
rect 48372 -49922 48430 -49910
rect 48372 -50498 48384 -49922
rect 48418 -50498 48430 -49922
rect 48372 -50510 48430 -50498
rect 25410 -50816 25468 -50804
rect 28012 -51154 28070 -51142
rect 28012 -51730 28024 -51154
rect 28058 -51730 28070 -51154
rect 28012 -51742 28070 -51730
rect 29030 -51154 29088 -51142
rect 29030 -51730 29042 -51154
rect 29076 -51730 29088 -51154
rect 29030 -51742 29088 -51730
rect 30048 -51154 30106 -51142
rect 30048 -51730 30060 -51154
rect 30094 -51730 30106 -51154
rect 30048 -51742 30106 -51730
rect 31066 -51154 31124 -51142
rect 31066 -51730 31078 -51154
rect 31112 -51730 31124 -51154
rect 31066 -51742 31124 -51730
rect 32084 -51154 32142 -51142
rect 32084 -51730 32096 -51154
rect 32130 -51730 32142 -51154
rect 32084 -51742 32142 -51730
rect 33102 -51154 33160 -51142
rect 33102 -51730 33114 -51154
rect 33148 -51730 33160 -51154
rect 33102 -51742 33160 -51730
rect 34120 -51154 34178 -51142
rect 34120 -51730 34132 -51154
rect 34166 -51730 34178 -51154
rect 34120 -51742 34178 -51730
rect 35138 -51154 35196 -51142
rect 35138 -51730 35150 -51154
rect 35184 -51730 35196 -51154
rect 35138 -51742 35196 -51730
rect 36156 -51154 36214 -51142
rect 36156 -51730 36168 -51154
rect 36202 -51730 36214 -51154
rect 36156 -51742 36214 -51730
rect 37174 -51154 37232 -51142
rect 37174 -51730 37186 -51154
rect 37220 -51730 37232 -51154
rect 37174 -51742 37232 -51730
rect 38192 -51154 38250 -51142
rect 38192 -51730 38204 -51154
rect 38238 -51730 38250 -51154
rect 38192 -51742 38250 -51730
rect 39210 -51154 39268 -51142
rect 39210 -51730 39222 -51154
rect 39256 -51730 39268 -51154
rect 39210 -51742 39268 -51730
rect 40228 -51154 40286 -51142
rect 40228 -51730 40240 -51154
rect 40274 -51730 40286 -51154
rect 40228 -51742 40286 -51730
rect 41246 -51154 41304 -51142
rect 41246 -51730 41258 -51154
rect 41292 -51730 41304 -51154
rect 41246 -51742 41304 -51730
rect 42264 -51154 42322 -51142
rect 42264 -51730 42276 -51154
rect 42310 -51730 42322 -51154
rect 42264 -51742 42322 -51730
rect 43282 -51154 43340 -51142
rect 43282 -51730 43294 -51154
rect 43328 -51730 43340 -51154
rect 43282 -51742 43340 -51730
rect 44300 -51154 44358 -51142
rect 44300 -51730 44312 -51154
rect 44346 -51730 44358 -51154
rect 44300 -51742 44358 -51730
rect 45318 -51154 45376 -51142
rect 45318 -51730 45330 -51154
rect 45364 -51730 45376 -51154
rect 45318 -51742 45376 -51730
rect 46336 -51154 46394 -51142
rect 46336 -51730 46348 -51154
rect 46382 -51730 46394 -51154
rect 46336 -51742 46394 -51730
rect 47354 -51154 47412 -51142
rect 47354 -51730 47366 -51154
rect 47400 -51730 47412 -51154
rect 47354 -51742 47412 -51730
rect 48372 -51154 48430 -51142
rect 48372 -51730 48384 -51154
rect 48418 -51730 48430 -51154
rect 48372 -51742 48430 -51730
rect 14924 -52252 14982 -52240
rect 14924 -52828 14936 -52252
rect 14970 -52828 14982 -52252
rect 14924 -52840 14982 -52828
rect 15942 -52252 16000 -52240
rect 15942 -52828 15954 -52252
rect 15988 -52828 16000 -52252
rect 15942 -52840 16000 -52828
rect 16960 -52252 17018 -52240
rect 16960 -52828 16972 -52252
rect 17006 -52828 17018 -52252
rect 16960 -52840 17018 -52828
rect 17978 -52252 18036 -52240
rect 17978 -52828 17990 -52252
rect 18024 -52828 18036 -52252
rect 17978 -52840 18036 -52828
rect 18996 -52252 19054 -52240
rect 18996 -52828 19008 -52252
rect 19042 -52828 19054 -52252
rect 18996 -52840 19054 -52828
rect 20014 -52252 20072 -52240
rect 20014 -52828 20026 -52252
rect 20060 -52828 20072 -52252
rect 20014 -52840 20072 -52828
rect 21032 -52252 21090 -52240
rect 21032 -52828 21044 -52252
rect 21078 -52828 21090 -52252
rect 21032 -52840 21090 -52828
rect 22050 -52252 22108 -52240
rect 22050 -52828 22062 -52252
rect 22096 -52828 22108 -52252
rect 22050 -52840 22108 -52828
rect 23068 -52252 23126 -52240
rect 23068 -52828 23080 -52252
rect 23114 -52828 23126 -52252
rect 23068 -52840 23126 -52828
rect 24086 -52252 24144 -52240
rect 24086 -52828 24098 -52252
rect 24132 -52828 24144 -52252
rect 24086 -52840 24144 -52828
rect 25104 -52252 25162 -52240
rect 25104 -52828 25116 -52252
rect 25150 -52828 25162 -52252
rect 25104 -52840 25162 -52828
rect 26122 -52252 26180 -52240
rect 26122 -52828 26134 -52252
rect 26168 -52828 26180 -52252
rect 26122 -52840 26180 -52828
rect 28012 -52388 28070 -52376
rect 28012 -52964 28024 -52388
rect 28058 -52964 28070 -52388
rect 28012 -52976 28070 -52964
rect 29030 -52388 29088 -52376
rect 29030 -52964 29042 -52388
rect 29076 -52964 29088 -52388
rect 29030 -52976 29088 -52964
rect 30048 -52388 30106 -52376
rect 30048 -52964 30060 -52388
rect 30094 -52964 30106 -52388
rect 30048 -52976 30106 -52964
rect 31066 -52388 31124 -52376
rect 31066 -52964 31078 -52388
rect 31112 -52964 31124 -52388
rect 31066 -52976 31124 -52964
rect 32084 -52388 32142 -52376
rect 32084 -52964 32096 -52388
rect 32130 -52964 32142 -52388
rect 32084 -52976 32142 -52964
rect 33102 -52388 33160 -52376
rect 33102 -52964 33114 -52388
rect 33148 -52964 33160 -52388
rect 33102 -52976 33160 -52964
rect 34120 -52388 34178 -52376
rect 34120 -52964 34132 -52388
rect 34166 -52964 34178 -52388
rect 34120 -52976 34178 -52964
rect 35138 -52388 35196 -52376
rect 35138 -52964 35150 -52388
rect 35184 -52964 35196 -52388
rect 35138 -52976 35196 -52964
rect 36156 -52388 36214 -52376
rect 36156 -52964 36168 -52388
rect 36202 -52964 36214 -52388
rect 36156 -52976 36214 -52964
rect 37174 -52388 37232 -52376
rect 37174 -52964 37186 -52388
rect 37220 -52964 37232 -52388
rect 37174 -52976 37232 -52964
rect 38192 -52388 38250 -52376
rect 38192 -52964 38204 -52388
rect 38238 -52964 38250 -52388
rect 38192 -52976 38250 -52964
rect 39210 -52388 39268 -52376
rect 39210 -52964 39222 -52388
rect 39256 -52964 39268 -52388
rect 39210 -52976 39268 -52964
rect 40228 -52388 40286 -52376
rect 40228 -52964 40240 -52388
rect 40274 -52964 40286 -52388
rect 40228 -52976 40286 -52964
rect 41246 -52388 41304 -52376
rect 41246 -52964 41258 -52388
rect 41292 -52964 41304 -52388
rect 41246 -52976 41304 -52964
rect 42264 -52388 42322 -52376
rect 42264 -52964 42276 -52388
rect 42310 -52964 42322 -52388
rect 42264 -52976 42322 -52964
rect 43282 -52388 43340 -52376
rect 43282 -52964 43294 -52388
rect 43328 -52964 43340 -52388
rect 43282 -52976 43340 -52964
rect 44300 -52388 44358 -52376
rect 44300 -52964 44312 -52388
rect 44346 -52964 44358 -52388
rect 44300 -52976 44358 -52964
rect 45318 -52388 45376 -52376
rect 45318 -52964 45330 -52388
rect 45364 -52964 45376 -52388
rect 45318 -52976 45376 -52964
rect 46336 -52388 46394 -52376
rect 46336 -52964 46348 -52388
rect 46382 -52964 46394 -52388
rect 46336 -52976 46394 -52964
rect 47354 -52388 47412 -52376
rect 47354 -52964 47366 -52388
rect 47400 -52964 47412 -52388
rect 47354 -52976 47412 -52964
rect 48372 -52388 48430 -52376
rect 48372 -52964 48384 -52388
rect 48418 -52964 48430 -52388
rect 48372 -52976 48430 -52964
rect 14924 -53364 14982 -53352
rect 14924 -53940 14936 -53364
rect 14970 -53940 14982 -53364
rect 14924 -53952 14982 -53940
rect 15942 -53364 16000 -53352
rect 15942 -53940 15954 -53364
rect 15988 -53940 16000 -53364
rect 15942 -53952 16000 -53940
rect 16960 -53364 17018 -53352
rect 16960 -53940 16972 -53364
rect 17006 -53940 17018 -53364
rect 16960 -53952 17018 -53940
rect 17978 -53364 18036 -53352
rect 17978 -53940 17990 -53364
rect 18024 -53940 18036 -53364
rect 17978 -53952 18036 -53940
rect 18996 -53364 19054 -53352
rect 18996 -53940 19008 -53364
rect 19042 -53940 19054 -53364
rect 18996 -53952 19054 -53940
rect 20014 -53364 20072 -53352
rect 20014 -53940 20026 -53364
rect 20060 -53940 20072 -53364
rect 20014 -53952 20072 -53940
rect 21032 -53364 21090 -53352
rect 21032 -53940 21044 -53364
rect 21078 -53940 21090 -53364
rect 21032 -53952 21090 -53940
rect 22050 -53364 22108 -53352
rect 22050 -53940 22062 -53364
rect 22096 -53940 22108 -53364
rect 22050 -53952 22108 -53940
rect 23068 -53364 23126 -53352
rect 23068 -53940 23080 -53364
rect 23114 -53940 23126 -53364
rect 23068 -53952 23126 -53940
rect 24086 -53364 24144 -53352
rect 24086 -53940 24098 -53364
rect 24132 -53940 24144 -53364
rect 24086 -53952 24144 -53940
rect 25104 -53364 25162 -53352
rect 25104 -53940 25116 -53364
rect 25150 -53940 25162 -53364
rect 25104 -53952 25162 -53940
rect 26122 -53364 26180 -53352
rect 26122 -53940 26134 -53364
rect 26168 -53940 26180 -53364
rect 26122 -53952 26180 -53940
rect 28012 -53622 28070 -53610
rect 28012 -54198 28024 -53622
rect 28058 -54198 28070 -53622
rect 28012 -54210 28070 -54198
rect 29030 -53622 29088 -53610
rect 29030 -54198 29042 -53622
rect 29076 -54198 29088 -53622
rect 29030 -54210 29088 -54198
rect 30048 -53622 30106 -53610
rect 30048 -54198 30060 -53622
rect 30094 -54198 30106 -53622
rect 30048 -54210 30106 -54198
rect 31066 -53622 31124 -53610
rect 31066 -54198 31078 -53622
rect 31112 -54198 31124 -53622
rect 31066 -54210 31124 -54198
rect 32084 -53622 32142 -53610
rect 32084 -54198 32096 -53622
rect 32130 -54198 32142 -53622
rect 32084 -54210 32142 -54198
rect 33102 -53622 33160 -53610
rect 33102 -54198 33114 -53622
rect 33148 -54198 33160 -53622
rect 33102 -54210 33160 -54198
rect 34120 -53622 34178 -53610
rect 34120 -54198 34132 -53622
rect 34166 -54198 34178 -53622
rect 34120 -54210 34178 -54198
rect 35138 -53622 35196 -53610
rect 35138 -54198 35150 -53622
rect 35184 -54198 35196 -53622
rect 35138 -54210 35196 -54198
rect 36156 -53622 36214 -53610
rect 36156 -54198 36168 -53622
rect 36202 -54198 36214 -53622
rect 36156 -54210 36214 -54198
rect 37174 -53622 37232 -53610
rect 37174 -54198 37186 -53622
rect 37220 -54198 37232 -53622
rect 37174 -54210 37232 -54198
rect 38192 -53622 38250 -53610
rect 38192 -54198 38204 -53622
rect 38238 -54198 38250 -53622
rect 38192 -54210 38250 -54198
rect 39210 -53622 39268 -53610
rect 39210 -54198 39222 -53622
rect 39256 -54198 39268 -53622
rect 39210 -54210 39268 -54198
rect 40228 -53622 40286 -53610
rect 40228 -54198 40240 -53622
rect 40274 -54198 40286 -53622
rect 40228 -54210 40286 -54198
rect 41246 -53622 41304 -53610
rect 41246 -54198 41258 -53622
rect 41292 -54198 41304 -53622
rect 41246 -54210 41304 -54198
rect 42264 -53622 42322 -53610
rect 42264 -54198 42276 -53622
rect 42310 -54198 42322 -53622
rect 42264 -54210 42322 -54198
rect 43282 -53622 43340 -53610
rect 43282 -54198 43294 -53622
rect 43328 -54198 43340 -53622
rect 43282 -54210 43340 -54198
rect 44300 -53622 44358 -53610
rect 44300 -54198 44312 -53622
rect 44346 -54198 44358 -53622
rect 44300 -54210 44358 -54198
rect 45318 -53622 45376 -53610
rect 45318 -54198 45330 -53622
rect 45364 -54198 45376 -53622
rect 45318 -54210 45376 -54198
rect 46336 -53622 46394 -53610
rect 46336 -54198 46348 -53622
rect 46382 -54198 46394 -53622
rect 46336 -54210 46394 -54198
rect 47354 -53622 47412 -53610
rect 47354 -54198 47366 -53622
rect 47400 -54198 47412 -53622
rect 47354 -54210 47412 -54198
rect 48372 -53622 48430 -53610
rect 48372 -54198 48384 -53622
rect 48418 -54198 48430 -53622
rect 48372 -54210 48430 -54198
rect 14924 -54476 14982 -54464
rect 14924 -55052 14936 -54476
rect 14970 -55052 14982 -54476
rect 14924 -55064 14982 -55052
rect 15942 -54476 16000 -54464
rect 15942 -55052 15954 -54476
rect 15988 -55052 16000 -54476
rect 15942 -55064 16000 -55052
rect 16960 -54476 17018 -54464
rect 16960 -55052 16972 -54476
rect 17006 -55052 17018 -54476
rect 16960 -55064 17018 -55052
rect 17978 -54476 18036 -54464
rect 17978 -55052 17990 -54476
rect 18024 -55052 18036 -54476
rect 17978 -55064 18036 -55052
rect 18996 -54476 19054 -54464
rect 18996 -55052 19008 -54476
rect 19042 -55052 19054 -54476
rect 18996 -55064 19054 -55052
rect 20014 -54476 20072 -54464
rect 20014 -55052 20026 -54476
rect 20060 -55052 20072 -54476
rect 20014 -55064 20072 -55052
rect 21032 -54476 21090 -54464
rect 21032 -55052 21044 -54476
rect 21078 -55052 21090 -54476
rect 21032 -55064 21090 -55052
rect 22050 -54476 22108 -54464
rect 22050 -55052 22062 -54476
rect 22096 -55052 22108 -54476
rect 22050 -55064 22108 -55052
rect 23068 -54476 23126 -54464
rect 23068 -55052 23080 -54476
rect 23114 -55052 23126 -54476
rect 23068 -55064 23126 -55052
rect 24086 -54476 24144 -54464
rect 24086 -55052 24098 -54476
rect 24132 -55052 24144 -54476
rect 24086 -55064 24144 -55052
rect 25104 -54476 25162 -54464
rect 25104 -55052 25116 -54476
rect 25150 -55052 25162 -54476
rect 25104 -55064 25162 -55052
rect 26122 -54476 26180 -54464
rect 26122 -55052 26134 -54476
rect 26168 -55052 26180 -54476
rect 26122 -55064 26180 -55052
rect 28012 -54854 28070 -54842
rect 28012 -55430 28024 -54854
rect 28058 -55430 28070 -54854
rect 28012 -55442 28070 -55430
rect 29030 -54854 29088 -54842
rect 29030 -55430 29042 -54854
rect 29076 -55430 29088 -54854
rect 29030 -55442 29088 -55430
rect 30048 -54854 30106 -54842
rect 30048 -55430 30060 -54854
rect 30094 -55430 30106 -54854
rect 30048 -55442 30106 -55430
rect 31066 -54854 31124 -54842
rect 31066 -55430 31078 -54854
rect 31112 -55430 31124 -54854
rect 31066 -55442 31124 -55430
rect 32084 -54854 32142 -54842
rect 32084 -55430 32096 -54854
rect 32130 -55430 32142 -54854
rect 32084 -55442 32142 -55430
rect 33102 -54854 33160 -54842
rect 33102 -55430 33114 -54854
rect 33148 -55430 33160 -54854
rect 33102 -55442 33160 -55430
rect 34120 -54854 34178 -54842
rect 34120 -55430 34132 -54854
rect 34166 -55430 34178 -54854
rect 34120 -55442 34178 -55430
rect 35138 -54854 35196 -54842
rect 35138 -55430 35150 -54854
rect 35184 -55430 35196 -54854
rect 35138 -55442 35196 -55430
rect 36156 -54854 36214 -54842
rect 36156 -55430 36168 -54854
rect 36202 -55430 36214 -54854
rect 36156 -55442 36214 -55430
rect 37174 -54854 37232 -54842
rect 37174 -55430 37186 -54854
rect 37220 -55430 37232 -54854
rect 37174 -55442 37232 -55430
rect 38192 -54854 38250 -54842
rect 38192 -55430 38204 -54854
rect 38238 -55430 38250 -54854
rect 38192 -55442 38250 -55430
rect 39210 -54854 39268 -54842
rect 39210 -55430 39222 -54854
rect 39256 -55430 39268 -54854
rect 39210 -55442 39268 -55430
rect 40228 -54854 40286 -54842
rect 40228 -55430 40240 -54854
rect 40274 -55430 40286 -54854
rect 40228 -55442 40286 -55430
rect 41246 -54854 41304 -54842
rect 41246 -55430 41258 -54854
rect 41292 -55430 41304 -54854
rect 41246 -55442 41304 -55430
rect 42264 -54854 42322 -54842
rect 42264 -55430 42276 -54854
rect 42310 -55430 42322 -54854
rect 42264 -55442 42322 -55430
rect 43282 -54854 43340 -54842
rect 43282 -55430 43294 -54854
rect 43328 -55430 43340 -54854
rect 43282 -55442 43340 -55430
rect 44300 -54854 44358 -54842
rect 44300 -55430 44312 -54854
rect 44346 -55430 44358 -54854
rect 44300 -55442 44358 -55430
rect 45318 -54854 45376 -54842
rect 45318 -55430 45330 -54854
rect 45364 -55430 45376 -54854
rect 45318 -55442 45376 -55430
rect 46336 -54854 46394 -54842
rect 46336 -55430 46348 -54854
rect 46382 -55430 46394 -54854
rect 46336 -55442 46394 -55430
rect 47354 -54854 47412 -54842
rect 47354 -55430 47366 -54854
rect 47400 -55430 47412 -54854
rect 47354 -55442 47412 -55430
rect 48372 -54854 48430 -54842
rect 48372 -55430 48384 -54854
rect 48418 -55430 48430 -54854
rect 48372 -55442 48430 -55430
rect 14924 -55588 14982 -55576
rect 14924 -56164 14936 -55588
rect 14970 -56164 14982 -55588
rect 14924 -56176 14982 -56164
rect 15942 -55588 16000 -55576
rect 15942 -56164 15954 -55588
rect 15988 -56164 16000 -55588
rect 15942 -56176 16000 -56164
rect 16960 -55588 17018 -55576
rect 16960 -56164 16972 -55588
rect 17006 -56164 17018 -55588
rect 16960 -56176 17018 -56164
rect 17978 -55588 18036 -55576
rect 17978 -56164 17990 -55588
rect 18024 -56164 18036 -55588
rect 17978 -56176 18036 -56164
rect 18996 -55588 19054 -55576
rect 18996 -56164 19008 -55588
rect 19042 -56164 19054 -55588
rect 18996 -56176 19054 -56164
rect 20014 -55588 20072 -55576
rect 20014 -56164 20026 -55588
rect 20060 -56164 20072 -55588
rect 20014 -56176 20072 -56164
rect 21032 -55588 21090 -55576
rect 21032 -56164 21044 -55588
rect 21078 -56164 21090 -55588
rect 21032 -56176 21090 -56164
rect 22050 -55588 22108 -55576
rect 22050 -56164 22062 -55588
rect 22096 -56164 22108 -55588
rect 22050 -56176 22108 -56164
rect 23068 -55588 23126 -55576
rect 23068 -56164 23080 -55588
rect 23114 -56164 23126 -55588
rect 23068 -56176 23126 -56164
rect 24086 -55588 24144 -55576
rect 24086 -56164 24098 -55588
rect 24132 -56164 24144 -55588
rect 24086 -56176 24144 -56164
rect 25104 -55588 25162 -55576
rect 25104 -56164 25116 -55588
rect 25150 -56164 25162 -55588
rect 25104 -56176 25162 -56164
rect 26122 -55588 26180 -55576
rect 26122 -56164 26134 -55588
rect 26168 -56164 26180 -55588
rect 26122 -56176 26180 -56164
rect 28012 -56088 28070 -56076
rect 28012 -56664 28024 -56088
rect 28058 -56664 28070 -56088
rect 28012 -56676 28070 -56664
rect 29030 -56088 29088 -56076
rect 29030 -56664 29042 -56088
rect 29076 -56664 29088 -56088
rect 29030 -56676 29088 -56664
rect 30048 -56088 30106 -56076
rect 30048 -56664 30060 -56088
rect 30094 -56664 30106 -56088
rect 30048 -56676 30106 -56664
rect 31066 -56088 31124 -56076
rect 31066 -56664 31078 -56088
rect 31112 -56664 31124 -56088
rect 31066 -56676 31124 -56664
rect 32084 -56088 32142 -56076
rect 32084 -56664 32096 -56088
rect 32130 -56664 32142 -56088
rect 32084 -56676 32142 -56664
rect 33102 -56088 33160 -56076
rect 33102 -56664 33114 -56088
rect 33148 -56664 33160 -56088
rect 33102 -56676 33160 -56664
rect 34120 -56088 34178 -56076
rect 34120 -56664 34132 -56088
rect 34166 -56664 34178 -56088
rect 34120 -56676 34178 -56664
rect 35138 -56088 35196 -56076
rect 35138 -56664 35150 -56088
rect 35184 -56664 35196 -56088
rect 35138 -56676 35196 -56664
rect 36156 -56088 36214 -56076
rect 36156 -56664 36168 -56088
rect 36202 -56664 36214 -56088
rect 36156 -56676 36214 -56664
rect 37174 -56088 37232 -56076
rect 37174 -56664 37186 -56088
rect 37220 -56664 37232 -56088
rect 37174 -56676 37232 -56664
rect 38192 -56088 38250 -56076
rect 38192 -56664 38204 -56088
rect 38238 -56664 38250 -56088
rect 38192 -56676 38250 -56664
rect 39210 -56088 39268 -56076
rect 39210 -56664 39222 -56088
rect 39256 -56664 39268 -56088
rect 39210 -56676 39268 -56664
rect 40228 -56088 40286 -56076
rect 40228 -56664 40240 -56088
rect 40274 -56664 40286 -56088
rect 40228 -56676 40286 -56664
rect 41246 -56088 41304 -56076
rect 41246 -56664 41258 -56088
rect 41292 -56664 41304 -56088
rect 41246 -56676 41304 -56664
rect 42264 -56088 42322 -56076
rect 42264 -56664 42276 -56088
rect 42310 -56664 42322 -56088
rect 42264 -56676 42322 -56664
rect 43282 -56088 43340 -56076
rect 43282 -56664 43294 -56088
rect 43328 -56664 43340 -56088
rect 43282 -56676 43340 -56664
rect 44300 -56088 44358 -56076
rect 44300 -56664 44312 -56088
rect 44346 -56664 44358 -56088
rect 44300 -56676 44358 -56664
rect 45318 -56088 45376 -56076
rect 45318 -56664 45330 -56088
rect 45364 -56664 45376 -56088
rect 45318 -56676 45376 -56664
rect 46336 -56088 46394 -56076
rect 46336 -56664 46348 -56088
rect 46382 -56664 46394 -56088
rect 46336 -56676 46394 -56664
rect 47354 -56088 47412 -56076
rect 47354 -56664 47366 -56088
rect 47400 -56664 47412 -56088
rect 47354 -56676 47412 -56664
rect 48372 -56088 48430 -56076
rect 48372 -56664 48384 -56088
rect 48418 -56664 48430 -56088
rect 48372 -56676 48430 -56664
rect 15382 -57130 15440 -57118
rect 15382 -57706 15394 -57130
rect 15428 -57706 15440 -57130
rect 15382 -57718 15440 -57706
rect 16400 -57130 16458 -57118
rect 16400 -57706 16412 -57130
rect 16446 -57706 16458 -57130
rect 16400 -57718 16458 -57706
rect 17418 -57130 17476 -57118
rect 17418 -57706 17430 -57130
rect 17464 -57706 17476 -57130
rect 17418 -57718 17476 -57706
rect 18436 -57130 18494 -57118
rect 18436 -57706 18448 -57130
rect 18482 -57706 18494 -57130
rect 18436 -57718 18494 -57706
rect 19454 -57130 19512 -57118
rect 19454 -57706 19466 -57130
rect 19500 -57706 19512 -57130
rect 19454 -57718 19512 -57706
rect 20472 -57130 20530 -57118
rect 20472 -57706 20484 -57130
rect 20518 -57706 20530 -57130
rect 20472 -57718 20530 -57706
rect 21490 -57130 21548 -57118
rect 21490 -57706 21502 -57130
rect 21536 -57706 21548 -57130
rect 21490 -57718 21548 -57706
rect 22508 -57130 22566 -57118
rect 22508 -57706 22520 -57130
rect 22554 -57706 22566 -57130
rect 22508 -57718 22566 -57706
rect 23526 -57130 23584 -57118
rect 23526 -57706 23538 -57130
rect 23572 -57706 23584 -57130
rect 23526 -57718 23584 -57706
rect 24544 -57130 24602 -57118
rect 24544 -57706 24556 -57130
rect 24590 -57706 24602 -57130
rect 24544 -57718 24602 -57706
rect 25562 -57130 25620 -57118
rect 25562 -57706 25574 -57130
rect 25608 -57706 25620 -57130
rect 25562 -57718 25620 -57706
rect 28012 -57320 28070 -57308
rect 28012 -57896 28024 -57320
rect 28058 -57896 28070 -57320
rect 28012 -57908 28070 -57896
rect 29030 -57320 29088 -57308
rect 29030 -57896 29042 -57320
rect 29076 -57896 29088 -57320
rect 29030 -57908 29088 -57896
rect 30048 -57320 30106 -57308
rect 30048 -57896 30060 -57320
rect 30094 -57896 30106 -57320
rect 30048 -57908 30106 -57896
rect 31066 -57320 31124 -57308
rect 31066 -57896 31078 -57320
rect 31112 -57896 31124 -57320
rect 31066 -57908 31124 -57896
rect 32084 -57320 32142 -57308
rect 32084 -57896 32096 -57320
rect 32130 -57896 32142 -57320
rect 32084 -57908 32142 -57896
rect 33102 -57320 33160 -57308
rect 33102 -57896 33114 -57320
rect 33148 -57896 33160 -57320
rect 33102 -57908 33160 -57896
rect 34120 -57320 34178 -57308
rect 34120 -57896 34132 -57320
rect 34166 -57896 34178 -57320
rect 34120 -57908 34178 -57896
rect 35138 -57320 35196 -57308
rect 35138 -57896 35150 -57320
rect 35184 -57896 35196 -57320
rect 35138 -57908 35196 -57896
rect 36156 -57320 36214 -57308
rect 36156 -57896 36168 -57320
rect 36202 -57896 36214 -57320
rect 36156 -57908 36214 -57896
rect 37174 -57320 37232 -57308
rect 37174 -57896 37186 -57320
rect 37220 -57896 37232 -57320
rect 37174 -57908 37232 -57896
rect 38192 -57320 38250 -57308
rect 38192 -57896 38204 -57320
rect 38238 -57896 38250 -57320
rect 38192 -57908 38250 -57896
rect 39210 -57320 39268 -57308
rect 39210 -57896 39222 -57320
rect 39256 -57896 39268 -57320
rect 39210 -57908 39268 -57896
rect 40228 -57320 40286 -57308
rect 40228 -57896 40240 -57320
rect 40274 -57896 40286 -57320
rect 40228 -57908 40286 -57896
rect 41246 -57320 41304 -57308
rect 41246 -57896 41258 -57320
rect 41292 -57896 41304 -57320
rect 41246 -57908 41304 -57896
rect 42264 -57320 42322 -57308
rect 42264 -57896 42276 -57320
rect 42310 -57896 42322 -57320
rect 42264 -57908 42322 -57896
rect 43282 -57320 43340 -57308
rect 43282 -57896 43294 -57320
rect 43328 -57896 43340 -57320
rect 43282 -57908 43340 -57896
rect 44300 -57320 44358 -57308
rect 44300 -57896 44312 -57320
rect 44346 -57896 44358 -57320
rect 44300 -57908 44358 -57896
rect 45318 -57320 45376 -57308
rect 45318 -57896 45330 -57320
rect 45364 -57896 45376 -57320
rect 45318 -57908 45376 -57896
rect 46336 -57320 46394 -57308
rect 46336 -57896 46348 -57320
rect 46382 -57896 46394 -57320
rect 46336 -57908 46394 -57896
rect 47354 -57320 47412 -57308
rect 47354 -57896 47366 -57320
rect 47400 -57896 47412 -57320
rect 47354 -57908 47412 -57896
rect 48372 -57320 48430 -57308
rect 48372 -57896 48384 -57320
rect 48418 -57896 48430 -57320
rect 48372 -57908 48430 -57896
rect 57908 -42714 57966 -42702
rect 57908 -42890 57920 -42714
rect 57954 -42890 57966 -42714
rect 57908 -42902 57966 -42890
rect 58026 -42714 58084 -42702
rect 58026 -42890 58038 -42714
rect 58072 -42890 58084 -42714
rect 58026 -42902 58084 -42890
rect -28004 -67661 -27952 -67649
rect -28004 -67695 -27996 -67661
rect -27962 -67695 -27952 -67661
rect -28004 -67729 -27952 -67695
rect -28004 -67763 -27996 -67729
rect -27962 -67763 -27952 -67729
rect -28004 -67779 -27952 -67763
rect -27922 -67661 -27870 -67649
rect -27922 -67695 -27912 -67661
rect -27878 -67695 -27870 -67661
rect -27922 -67729 -27870 -67695
rect -27922 -67763 -27912 -67729
rect -27878 -67763 -27870 -67729
rect -27922 -67779 -27870 -67763
rect -24004 -67661 -23952 -67649
rect -24004 -67695 -23996 -67661
rect -23962 -67695 -23952 -67661
rect -24004 -67729 -23952 -67695
rect -24004 -67763 -23996 -67729
rect -23962 -67763 -23952 -67729
rect -24004 -67779 -23952 -67763
rect -23922 -67661 -23870 -67649
rect -23922 -67695 -23912 -67661
rect -23878 -67695 -23870 -67661
rect -23922 -67729 -23870 -67695
rect -23922 -67763 -23912 -67729
rect -23878 -67763 -23870 -67729
rect -23922 -67779 -23870 -67763
rect -20004 -67661 -19952 -67649
rect -20004 -67695 -19996 -67661
rect -19962 -67695 -19952 -67661
rect -20004 -67729 -19952 -67695
rect -20004 -67763 -19996 -67729
rect -19962 -67763 -19952 -67729
rect -27354 -68330 -27296 -68318
rect -27354 -68706 -27342 -68330
rect -27308 -68706 -27296 -68330
rect -27354 -68718 -27296 -68706
rect -27096 -68330 -27038 -68318
rect -27096 -68706 -27084 -68330
rect -27050 -68706 -27038 -68330
rect -27096 -68718 -27038 -68706
rect -26838 -68330 -26780 -68318
rect -26838 -68706 -26826 -68330
rect -26792 -68706 -26780 -68330
rect -26838 -68718 -26780 -68706
rect -26580 -68330 -26522 -68318
rect -26580 -68706 -26568 -68330
rect -26534 -68706 -26522 -68330
rect -26580 -68718 -26522 -68706
rect -26322 -68330 -26264 -68318
rect -26322 -68706 -26310 -68330
rect -26276 -68706 -26264 -68330
rect -26322 -68718 -26264 -68706
rect -26064 -68330 -26006 -68318
rect -26064 -68706 -26052 -68330
rect -26018 -68706 -26006 -68330
rect -26064 -68718 -26006 -68706
rect -25806 -68330 -25748 -68318
rect -25806 -68706 -25794 -68330
rect -25760 -68706 -25748 -68330
rect -25806 -68718 -25748 -68706
rect -20004 -67779 -19952 -67763
rect -19922 -67661 -19870 -67649
rect -19922 -67695 -19912 -67661
rect -19878 -67695 -19870 -67661
rect -19922 -67729 -19870 -67695
rect -19922 -67763 -19912 -67729
rect -19878 -67763 -19870 -67729
rect -19922 -67779 -19870 -67763
rect -16004 -67661 -15952 -67649
rect -16004 -67695 -15996 -67661
rect -15962 -67695 -15952 -67661
rect -16004 -67729 -15952 -67695
rect -16004 -67763 -15996 -67729
rect -15962 -67763 -15952 -67729
rect -23354 -68330 -23296 -68318
rect -23354 -68706 -23342 -68330
rect -23308 -68706 -23296 -68330
rect -23354 -68718 -23296 -68706
rect -23096 -68330 -23038 -68318
rect -23096 -68706 -23084 -68330
rect -23050 -68706 -23038 -68330
rect -23096 -68718 -23038 -68706
rect -22838 -68330 -22780 -68318
rect -22838 -68706 -22826 -68330
rect -22792 -68706 -22780 -68330
rect -22838 -68718 -22780 -68706
rect -22580 -68330 -22522 -68318
rect -22580 -68706 -22568 -68330
rect -22534 -68706 -22522 -68330
rect -22580 -68718 -22522 -68706
rect -22322 -68330 -22264 -68318
rect -22322 -68706 -22310 -68330
rect -22276 -68706 -22264 -68330
rect -22322 -68718 -22264 -68706
rect -22064 -68330 -22006 -68318
rect -22064 -68706 -22052 -68330
rect -22018 -68706 -22006 -68330
rect -22064 -68718 -22006 -68706
rect -21806 -68330 -21748 -68318
rect -21806 -68706 -21794 -68330
rect -21760 -68706 -21748 -68330
rect -21806 -68718 -21748 -68706
rect -16004 -67779 -15952 -67763
rect -15922 -67661 -15870 -67649
rect -15922 -67695 -15912 -67661
rect -15878 -67695 -15870 -67661
rect -15922 -67729 -15870 -67695
rect -15922 -67763 -15912 -67729
rect -15878 -67763 -15870 -67729
rect -15922 -67779 -15870 -67763
rect -12004 -67661 -11952 -67649
rect -12004 -67695 -11996 -67661
rect -11962 -67695 -11952 -67661
rect -12004 -67729 -11952 -67695
rect -12004 -67763 -11996 -67729
rect -11962 -67763 -11952 -67729
rect -19354 -68330 -19296 -68318
rect -19354 -68706 -19342 -68330
rect -19308 -68706 -19296 -68330
rect -19354 -68718 -19296 -68706
rect -19096 -68330 -19038 -68318
rect -19096 -68706 -19084 -68330
rect -19050 -68706 -19038 -68330
rect -19096 -68718 -19038 -68706
rect -18838 -68330 -18780 -68318
rect -18838 -68706 -18826 -68330
rect -18792 -68706 -18780 -68330
rect -18838 -68718 -18780 -68706
rect -18580 -68330 -18522 -68318
rect -18580 -68706 -18568 -68330
rect -18534 -68706 -18522 -68330
rect -18580 -68718 -18522 -68706
rect -18322 -68330 -18264 -68318
rect -18322 -68706 -18310 -68330
rect -18276 -68706 -18264 -68330
rect -18322 -68718 -18264 -68706
rect -18064 -68330 -18006 -68318
rect -18064 -68706 -18052 -68330
rect -18018 -68706 -18006 -68330
rect -18064 -68718 -18006 -68706
rect -17806 -68330 -17748 -68318
rect -17806 -68706 -17794 -68330
rect -17760 -68706 -17748 -68330
rect -17806 -68718 -17748 -68706
rect -12004 -67779 -11952 -67763
rect -11922 -67661 -11870 -67649
rect -11922 -67695 -11912 -67661
rect -11878 -67695 -11870 -67661
rect -11922 -67729 -11870 -67695
rect -11922 -67763 -11912 -67729
rect -11878 -67763 -11870 -67729
rect -11922 -67779 -11870 -67763
rect -8004 -67661 -7952 -67649
rect -8004 -67695 -7996 -67661
rect -7962 -67695 -7952 -67661
rect -8004 -67729 -7952 -67695
rect -8004 -67763 -7996 -67729
rect -7962 -67763 -7952 -67729
rect -15354 -68330 -15296 -68318
rect -15354 -68706 -15342 -68330
rect -15308 -68706 -15296 -68330
rect -15354 -68718 -15296 -68706
rect -15096 -68330 -15038 -68318
rect -15096 -68706 -15084 -68330
rect -15050 -68706 -15038 -68330
rect -15096 -68718 -15038 -68706
rect -14838 -68330 -14780 -68318
rect -14838 -68706 -14826 -68330
rect -14792 -68706 -14780 -68330
rect -14838 -68718 -14780 -68706
rect -14580 -68330 -14522 -68318
rect -14580 -68706 -14568 -68330
rect -14534 -68706 -14522 -68330
rect -14580 -68718 -14522 -68706
rect -14322 -68330 -14264 -68318
rect -14322 -68706 -14310 -68330
rect -14276 -68706 -14264 -68330
rect -14322 -68718 -14264 -68706
rect -14064 -68330 -14006 -68318
rect -14064 -68706 -14052 -68330
rect -14018 -68706 -14006 -68330
rect -14064 -68718 -14006 -68706
rect -13806 -68330 -13748 -68318
rect -13806 -68706 -13794 -68330
rect -13760 -68706 -13748 -68330
rect -13806 -68718 -13748 -68706
rect -8004 -67779 -7952 -67763
rect -7922 -67661 -7870 -67649
rect -7922 -67695 -7912 -67661
rect -7878 -67695 -7870 -67661
rect -7922 -67729 -7870 -67695
rect -7922 -67763 -7912 -67729
rect -7878 -67763 -7870 -67729
rect -7922 -67779 -7870 -67763
rect -4004 -67661 -3952 -67649
rect -4004 -67695 -3996 -67661
rect -3962 -67695 -3952 -67661
rect -4004 -67729 -3952 -67695
rect -4004 -67763 -3996 -67729
rect -3962 -67763 -3952 -67729
rect -11354 -68330 -11296 -68318
rect -11354 -68706 -11342 -68330
rect -11308 -68706 -11296 -68330
rect -11354 -68718 -11296 -68706
rect -11096 -68330 -11038 -68318
rect -11096 -68706 -11084 -68330
rect -11050 -68706 -11038 -68330
rect -11096 -68718 -11038 -68706
rect -10838 -68330 -10780 -68318
rect -10838 -68706 -10826 -68330
rect -10792 -68706 -10780 -68330
rect -10838 -68718 -10780 -68706
rect -10580 -68330 -10522 -68318
rect -10580 -68706 -10568 -68330
rect -10534 -68706 -10522 -68330
rect -10580 -68718 -10522 -68706
rect -10322 -68330 -10264 -68318
rect -10322 -68706 -10310 -68330
rect -10276 -68706 -10264 -68330
rect -10322 -68718 -10264 -68706
rect -10064 -68330 -10006 -68318
rect -10064 -68706 -10052 -68330
rect -10018 -68706 -10006 -68330
rect -10064 -68718 -10006 -68706
rect -9806 -68330 -9748 -68318
rect -9806 -68706 -9794 -68330
rect -9760 -68706 -9748 -68330
rect -9806 -68718 -9748 -68706
rect -4004 -67779 -3952 -67763
rect -3922 -67661 -3870 -67649
rect -3922 -67695 -3912 -67661
rect -3878 -67695 -3870 -67661
rect -3922 -67729 -3870 -67695
rect -3922 -67763 -3912 -67729
rect -3878 -67763 -3870 -67729
rect -3922 -67779 -3870 -67763
rect -4 -67661 48 -67649
rect -4 -67695 4 -67661
rect 38 -67695 48 -67661
rect -4 -67729 48 -67695
rect -4 -67763 4 -67729
rect 38 -67763 48 -67729
rect -7354 -68330 -7296 -68318
rect -7354 -68706 -7342 -68330
rect -7308 -68706 -7296 -68330
rect -7354 -68718 -7296 -68706
rect -7096 -68330 -7038 -68318
rect -7096 -68706 -7084 -68330
rect -7050 -68706 -7038 -68330
rect -7096 -68718 -7038 -68706
rect -6838 -68330 -6780 -68318
rect -6838 -68706 -6826 -68330
rect -6792 -68706 -6780 -68330
rect -6838 -68718 -6780 -68706
rect -6580 -68330 -6522 -68318
rect -6580 -68706 -6568 -68330
rect -6534 -68706 -6522 -68330
rect -6580 -68718 -6522 -68706
rect -6322 -68330 -6264 -68318
rect -6322 -68706 -6310 -68330
rect -6276 -68706 -6264 -68330
rect -6322 -68718 -6264 -68706
rect -6064 -68330 -6006 -68318
rect -6064 -68706 -6052 -68330
rect -6018 -68706 -6006 -68330
rect -6064 -68718 -6006 -68706
rect -5806 -68330 -5748 -68318
rect -5806 -68706 -5794 -68330
rect -5760 -68706 -5748 -68330
rect -5806 -68718 -5748 -68706
rect -4 -67779 48 -67763
rect 78 -67661 130 -67649
rect 78 -67695 88 -67661
rect 122 -67695 130 -67661
rect 78 -67729 130 -67695
rect 78 -67763 88 -67729
rect 122 -67763 130 -67729
rect 78 -67779 130 -67763
rect 3996 -67661 4048 -67649
rect 3996 -67695 4004 -67661
rect 4038 -67695 4048 -67661
rect 3996 -67729 4048 -67695
rect 3996 -67763 4004 -67729
rect 4038 -67763 4048 -67729
rect -3354 -68330 -3296 -68318
rect -3354 -68706 -3342 -68330
rect -3308 -68706 -3296 -68330
rect -3354 -68718 -3296 -68706
rect -3096 -68330 -3038 -68318
rect -3096 -68706 -3084 -68330
rect -3050 -68706 -3038 -68330
rect -3096 -68718 -3038 -68706
rect -2838 -68330 -2780 -68318
rect -2838 -68706 -2826 -68330
rect -2792 -68706 -2780 -68330
rect -2838 -68718 -2780 -68706
rect -2580 -68330 -2522 -68318
rect -2580 -68706 -2568 -68330
rect -2534 -68706 -2522 -68330
rect -2580 -68718 -2522 -68706
rect -2322 -68330 -2264 -68318
rect -2322 -68706 -2310 -68330
rect -2276 -68706 -2264 -68330
rect -2322 -68718 -2264 -68706
rect -2064 -68330 -2006 -68318
rect -2064 -68706 -2052 -68330
rect -2018 -68706 -2006 -68330
rect -2064 -68718 -2006 -68706
rect -1806 -68330 -1748 -68318
rect -1806 -68706 -1794 -68330
rect -1760 -68706 -1748 -68330
rect -1806 -68718 -1748 -68706
rect 3996 -67779 4048 -67763
rect 4078 -67661 4130 -67649
rect 4078 -67695 4088 -67661
rect 4122 -67695 4130 -67661
rect 4078 -67729 4130 -67695
rect 4078 -67763 4088 -67729
rect 4122 -67763 4130 -67729
rect 4078 -67779 4130 -67763
rect 646 -68330 704 -68318
rect 646 -68706 658 -68330
rect 692 -68706 704 -68330
rect 646 -68718 704 -68706
rect 904 -68330 962 -68318
rect 904 -68706 916 -68330
rect 950 -68706 962 -68330
rect 904 -68718 962 -68706
rect 1162 -68330 1220 -68318
rect 1162 -68706 1174 -68330
rect 1208 -68706 1220 -68330
rect 1162 -68718 1220 -68706
rect 1420 -68330 1478 -68318
rect 1420 -68706 1432 -68330
rect 1466 -68706 1478 -68330
rect 1420 -68718 1478 -68706
rect 1678 -68330 1736 -68318
rect 1678 -68706 1690 -68330
rect 1724 -68706 1736 -68330
rect 1678 -68718 1736 -68706
rect 1936 -68330 1994 -68318
rect 1936 -68706 1948 -68330
rect 1982 -68706 1994 -68330
rect 1936 -68718 1994 -68706
rect 2194 -68330 2252 -68318
rect 2194 -68706 2206 -68330
rect 2240 -68706 2252 -68330
rect 2194 -68718 2252 -68706
rect 4646 -68330 4704 -68318
rect 4646 -68706 4658 -68330
rect 4692 -68706 4704 -68330
rect 4646 -68718 4704 -68706
rect 4904 -68330 4962 -68318
rect 4904 -68706 4916 -68330
rect 4950 -68706 4962 -68330
rect 4904 -68718 4962 -68706
rect 5162 -68330 5220 -68318
rect 5162 -68706 5174 -68330
rect 5208 -68706 5220 -68330
rect 5162 -68718 5220 -68706
rect 5420 -68330 5478 -68318
rect 5420 -68706 5432 -68330
rect 5466 -68706 5478 -68330
rect 5420 -68718 5478 -68706
rect 5678 -68330 5736 -68318
rect 5678 -68706 5690 -68330
rect 5724 -68706 5736 -68330
rect 5678 -68718 5736 -68706
rect 5936 -68330 5994 -68318
rect 5936 -68706 5948 -68330
rect 5982 -68706 5994 -68330
rect 5936 -68718 5994 -68706
rect 6194 -68330 6252 -68318
rect 6194 -68706 6206 -68330
rect 6240 -68706 6252 -68330
rect 6194 -68718 6252 -68706
rect -27354 -71490 -27296 -71478
rect -27354 -71866 -27342 -71490
rect -27308 -71866 -27296 -71490
rect -27354 -71878 -27296 -71866
rect -27096 -71490 -27038 -71478
rect -27096 -71866 -27084 -71490
rect -27050 -71866 -27038 -71490
rect -27096 -71878 -27038 -71866
rect -26838 -71490 -26780 -71478
rect -26838 -71866 -26826 -71490
rect -26792 -71866 -26780 -71490
rect -26838 -71878 -26780 -71866
rect -26580 -71490 -26522 -71478
rect -26580 -71866 -26568 -71490
rect -26534 -71866 -26522 -71490
rect -26580 -71878 -26522 -71866
rect -26322 -71490 -26264 -71478
rect -26322 -71866 -26310 -71490
rect -26276 -71866 -26264 -71490
rect -26322 -71878 -26264 -71866
rect -26064 -71490 -26006 -71478
rect -26064 -71866 -26052 -71490
rect -26018 -71866 -26006 -71490
rect -26064 -71878 -26006 -71866
rect -25806 -71490 -25748 -71478
rect -25806 -71866 -25794 -71490
rect -25760 -71866 -25748 -71490
rect -25806 -71878 -25748 -71866
rect -28004 -72433 -27952 -72417
rect -28004 -72467 -27996 -72433
rect -27962 -72467 -27952 -72433
rect -28004 -72501 -27952 -72467
rect -28004 -72535 -27996 -72501
rect -27962 -72535 -27952 -72501
rect -28004 -72547 -27952 -72535
rect -27922 -72433 -27870 -72417
rect -23354 -71490 -23296 -71478
rect -23354 -71866 -23342 -71490
rect -23308 -71866 -23296 -71490
rect -23354 -71878 -23296 -71866
rect -23096 -71490 -23038 -71478
rect -23096 -71866 -23084 -71490
rect -23050 -71866 -23038 -71490
rect -23096 -71878 -23038 -71866
rect -22838 -71490 -22780 -71478
rect -22838 -71866 -22826 -71490
rect -22792 -71866 -22780 -71490
rect -22838 -71878 -22780 -71866
rect -22580 -71490 -22522 -71478
rect -22580 -71866 -22568 -71490
rect -22534 -71866 -22522 -71490
rect -22580 -71878 -22522 -71866
rect -22322 -71490 -22264 -71478
rect -22322 -71866 -22310 -71490
rect -22276 -71866 -22264 -71490
rect -22322 -71878 -22264 -71866
rect -22064 -71490 -22006 -71478
rect -22064 -71866 -22052 -71490
rect -22018 -71866 -22006 -71490
rect -22064 -71878 -22006 -71866
rect -21806 -71490 -21748 -71478
rect -21806 -71866 -21794 -71490
rect -21760 -71866 -21748 -71490
rect -21806 -71878 -21748 -71866
rect -27922 -72467 -27912 -72433
rect -27878 -72467 -27870 -72433
rect -27922 -72501 -27870 -72467
rect -27922 -72535 -27912 -72501
rect -27878 -72535 -27870 -72501
rect -27922 -72547 -27870 -72535
rect -24004 -72433 -23952 -72417
rect -24004 -72467 -23996 -72433
rect -23962 -72467 -23952 -72433
rect -24004 -72501 -23952 -72467
rect -24004 -72535 -23996 -72501
rect -23962 -72535 -23952 -72501
rect -24004 -72547 -23952 -72535
rect -23922 -72433 -23870 -72417
rect -19354 -71490 -19296 -71478
rect -19354 -71866 -19342 -71490
rect -19308 -71866 -19296 -71490
rect -19354 -71878 -19296 -71866
rect -19096 -71490 -19038 -71478
rect -19096 -71866 -19084 -71490
rect -19050 -71866 -19038 -71490
rect -19096 -71878 -19038 -71866
rect -18838 -71490 -18780 -71478
rect -18838 -71866 -18826 -71490
rect -18792 -71866 -18780 -71490
rect -18838 -71878 -18780 -71866
rect -18580 -71490 -18522 -71478
rect -18580 -71866 -18568 -71490
rect -18534 -71866 -18522 -71490
rect -18580 -71878 -18522 -71866
rect -18322 -71490 -18264 -71478
rect -18322 -71866 -18310 -71490
rect -18276 -71866 -18264 -71490
rect -18322 -71878 -18264 -71866
rect -18064 -71490 -18006 -71478
rect -18064 -71866 -18052 -71490
rect -18018 -71866 -18006 -71490
rect -18064 -71878 -18006 -71866
rect -17806 -71490 -17748 -71478
rect -17806 -71866 -17794 -71490
rect -17760 -71866 -17748 -71490
rect -17806 -71878 -17748 -71866
rect -23922 -72467 -23912 -72433
rect -23878 -72467 -23870 -72433
rect -23922 -72501 -23870 -72467
rect -23922 -72535 -23912 -72501
rect -23878 -72535 -23870 -72501
rect -23922 -72547 -23870 -72535
rect -20004 -72433 -19952 -72417
rect -20004 -72467 -19996 -72433
rect -19962 -72467 -19952 -72433
rect -20004 -72501 -19952 -72467
rect -20004 -72535 -19996 -72501
rect -19962 -72535 -19952 -72501
rect -20004 -72547 -19952 -72535
rect -19922 -72433 -19870 -72417
rect -15354 -71490 -15296 -71478
rect -15354 -71866 -15342 -71490
rect -15308 -71866 -15296 -71490
rect -15354 -71878 -15296 -71866
rect -15096 -71490 -15038 -71478
rect -15096 -71866 -15084 -71490
rect -15050 -71866 -15038 -71490
rect -15096 -71878 -15038 -71866
rect -14838 -71490 -14780 -71478
rect -14838 -71866 -14826 -71490
rect -14792 -71866 -14780 -71490
rect -14838 -71878 -14780 -71866
rect -14580 -71490 -14522 -71478
rect -14580 -71866 -14568 -71490
rect -14534 -71866 -14522 -71490
rect -14580 -71878 -14522 -71866
rect -14322 -71490 -14264 -71478
rect -14322 -71866 -14310 -71490
rect -14276 -71866 -14264 -71490
rect -14322 -71878 -14264 -71866
rect -14064 -71490 -14006 -71478
rect -14064 -71866 -14052 -71490
rect -14018 -71866 -14006 -71490
rect -14064 -71878 -14006 -71866
rect -13806 -71490 -13748 -71478
rect -13806 -71866 -13794 -71490
rect -13760 -71866 -13748 -71490
rect -13806 -71878 -13748 -71866
rect -19922 -72467 -19912 -72433
rect -19878 -72467 -19870 -72433
rect -19922 -72501 -19870 -72467
rect -19922 -72535 -19912 -72501
rect -19878 -72535 -19870 -72501
rect -19922 -72547 -19870 -72535
rect -16004 -72433 -15952 -72417
rect -16004 -72467 -15996 -72433
rect -15962 -72467 -15952 -72433
rect -16004 -72501 -15952 -72467
rect -16004 -72535 -15996 -72501
rect -15962 -72535 -15952 -72501
rect -16004 -72547 -15952 -72535
rect -15922 -72433 -15870 -72417
rect -11354 -71490 -11296 -71478
rect -11354 -71866 -11342 -71490
rect -11308 -71866 -11296 -71490
rect -11354 -71878 -11296 -71866
rect -11096 -71490 -11038 -71478
rect -11096 -71866 -11084 -71490
rect -11050 -71866 -11038 -71490
rect -11096 -71878 -11038 -71866
rect -10838 -71490 -10780 -71478
rect -10838 -71866 -10826 -71490
rect -10792 -71866 -10780 -71490
rect -10838 -71878 -10780 -71866
rect -10580 -71490 -10522 -71478
rect -10580 -71866 -10568 -71490
rect -10534 -71866 -10522 -71490
rect -10580 -71878 -10522 -71866
rect -10322 -71490 -10264 -71478
rect -10322 -71866 -10310 -71490
rect -10276 -71866 -10264 -71490
rect -10322 -71878 -10264 -71866
rect -10064 -71490 -10006 -71478
rect -10064 -71866 -10052 -71490
rect -10018 -71866 -10006 -71490
rect -10064 -71878 -10006 -71866
rect -9806 -71490 -9748 -71478
rect -9806 -71866 -9794 -71490
rect -9760 -71866 -9748 -71490
rect -9806 -71878 -9748 -71866
rect -15922 -72467 -15912 -72433
rect -15878 -72467 -15870 -72433
rect -15922 -72501 -15870 -72467
rect -15922 -72535 -15912 -72501
rect -15878 -72535 -15870 -72501
rect -15922 -72547 -15870 -72535
rect -12004 -72433 -11952 -72417
rect -12004 -72467 -11996 -72433
rect -11962 -72467 -11952 -72433
rect -12004 -72501 -11952 -72467
rect -12004 -72535 -11996 -72501
rect -11962 -72535 -11952 -72501
rect -12004 -72547 -11952 -72535
rect -11922 -72433 -11870 -72417
rect -7354 -71490 -7296 -71478
rect -7354 -71866 -7342 -71490
rect -7308 -71866 -7296 -71490
rect -7354 -71878 -7296 -71866
rect -7096 -71490 -7038 -71478
rect -7096 -71866 -7084 -71490
rect -7050 -71866 -7038 -71490
rect -7096 -71878 -7038 -71866
rect -6838 -71490 -6780 -71478
rect -6838 -71866 -6826 -71490
rect -6792 -71866 -6780 -71490
rect -6838 -71878 -6780 -71866
rect -6580 -71490 -6522 -71478
rect -6580 -71866 -6568 -71490
rect -6534 -71866 -6522 -71490
rect -6580 -71878 -6522 -71866
rect -6322 -71490 -6264 -71478
rect -6322 -71866 -6310 -71490
rect -6276 -71866 -6264 -71490
rect -6322 -71878 -6264 -71866
rect -6064 -71490 -6006 -71478
rect -6064 -71866 -6052 -71490
rect -6018 -71866 -6006 -71490
rect -6064 -71878 -6006 -71866
rect -5806 -71490 -5748 -71478
rect -5806 -71866 -5794 -71490
rect -5760 -71866 -5748 -71490
rect -5806 -71878 -5748 -71866
rect -11922 -72467 -11912 -72433
rect -11878 -72467 -11870 -72433
rect -11922 -72501 -11870 -72467
rect -11922 -72535 -11912 -72501
rect -11878 -72535 -11870 -72501
rect -11922 -72547 -11870 -72535
rect -8004 -72433 -7952 -72417
rect -8004 -72467 -7996 -72433
rect -7962 -72467 -7952 -72433
rect -8004 -72501 -7952 -72467
rect -8004 -72535 -7996 -72501
rect -7962 -72535 -7952 -72501
rect -8004 -72547 -7952 -72535
rect -7922 -72433 -7870 -72417
rect -3354 -71490 -3296 -71478
rect -3354 -71866 -3342 -71490
rect -3308 -71866 -3296 -71490
rect -3354 -71878 -3296 -71866
rect -3096 -71490 -3038 -71478
rect -3096 -71866 -3084 -71490
rect -3050 -71866 -3038 -71490
rect -3096 -71878 -3038 -71866
rect -2838 -71490 -2780 -71478
rect -2838 -71866 -2826 -71490
rect -2792 -71866 -2780 -71490
rect -2838 -71878 -2780 -71866
rect -2580 -71490 -2522 -71478
rect -2580 -71866 -2568 -71490
rect -2534 -71866 -2522 -71490
rect -2580 -71878 -2522 -71866
rect -2322 -71490 -2264 -71478
rect -2322 -71866 -2310 -71490
rect -2276 -71866 -2264 -71490
rect -2322 -71878 -2264 -71866
rect -2064 -71490 -2006 -71478
rect -2064 -71866 -2052 -71490
rect -2018 -71866 -2006 -71490
rect -2064 -71878 -2006 -71866
rect -1806 -71490 -1748 -71478
rect -1806 -71866 -1794 -71490
rect -1760 -71866 -1748 -71490
rect -1806 -71878 -1748 -71866
rect -7922 -72467 -7912 -72433
rect -7878 -72467 -7870 -72433
rect -7922 -72501 -7870 -72467
rect -7922 -72535 -7912 -72501
rect -7878 -72535 -7870 -72501
rect -7922 -72547 -7870 -72535
rect -4004 -72433 -3952 -72417
rect -4004 -72467 -3996 -72433
rect -3962 -72467 -3952 -72433
rect -4004 -72501 -3952 -72467
rect -4004 -72535 -3996 -72501
rect -3962 -72535 -3952 -72501
rect -4004 -72547 -3952 -72535
rect -3922 -72433 -3870 -72417
rect 646 -71490 704 -71478
rect 646 -71866 658 -71490
rect 692 -71866 704 -71490
rect 646 -71878 704 -71866
rect 904 -71490 962 -71478
rect 904 -71866 916 -71490
rect 950 -71866 962 -71490
rect 904 -71878 962 -71866
rect 1162 -71490 1220 -71478
rect 1162 -71866 1174 -71490
rect 1208 -71866 1220 -71490
rect 1162 -71878 1220 -71866
rect 1420 -71490 1478 -71478
rect 1420 -71866 1432 -71490
rect 1466 -71866 1478 -71490
rect 1420 -71878 1478 -71866
rect 1678 -71490 1736 -71478
rect 1678 -71866 1690 -71490
rect 1724 -71866 1736 -71490
rect 1678 -71878 1736 -71866
rect 1936 -71490 1994 -71478
rect 1936 -71866 1948 -71490
rect 1982 -71866 1994 -71490
rect 1936 -71878 1994 -71866
rect 2194 -71490 2252 -71478
rect 2194 -71866 2206 -71490
rect 2240 -71866 2252 -71490
rect 2194 -71878 2252 -71866
rect -3922 -72467 -3912 -72433
rect -3878 -72467 -3870 -72433
rect -3922 -72501 -3870 -72467
rect -3922 -72535 -3912 -72501
rect -3878 -72535 -3870 -72501
rect -3922 -72547 -3870 -72535
rect -4 -72433 48 -72417
rect -4 -72467 4 -72433
rect 38 -72467 48 -72433
rect -4 -72501 48 -72467
rect -4 -72535 4 -72501
rect 38 -72535 48 -72501
rect -4 -72547 48 -72535
rect 78 -72433 130 -72417
rect 4646 -71490 4704 -71478
rect 4646 -71866 4658 -71490
rect 4692 -71866 4704 -71490
rect 4646 -71878 4704 -71866
rect 4904 -71490 4962 -71478
rect 4904 -71866 4916 -71490
rect 4950 -71866 4962 -71490
rect 4904 -71878 4962 -71866
rect 5162 -71490 5220 -71478
rect 5162 -71866 5174 -71490
rect 5208 -71866 5220 -71490
rect 5162 -71878 5220 -71866
rect 5420 -71490 5478 -71478
rect 5420 -71866 5432 -71490
rect 5466 -71866 5478 -71490
rect 5420 -71878 5478 -71866
rect 5678 -71490 5736 -71478
rect 5678 -71866 5690 -71490
rect 5724 -71866 5736 -71490
rect 5678 -71878 5736 -71866
rect 5936 -71490 5994 -71478
rect 5936 -71866 5948 -71490
rect 5982 -71866 5994 -71490
rect 5936 -71878 5994 -71866
rect 6194 -71490 6252 -71478
rect 6194 -71866 6206 -71490
rect 6240 -71866 6252 -71490
rect 6194 -71878 6252 -71866
rect 78 -72467 88 -72433
rect 122 -72467 130 -72433
rect 78 -72501 130 -72467
rect 78 -72535 88 -72501
rect 122 -72535 130 -72501
rect 78 -72547 130 -72535
rect 3996 -72433 4048 -72417
rect 3996 -72467 4004 -72433
rect 4038 -72467 4048 -72433
rect 3996 -72501 4048 -72467
rect 3996 -72535 4004 -72501
rect 4038 -72535 4048 -72501
rect 3996 -72547 4048 -72535
rect 4078 -72433 4130 -72417
rect 4078 -72467 4088 -72433
rect 4122 -72467 4130 -72433
rect 4078 -72501 4130 -72467
rect 4078 -72535 4088 -72501
rect 4122 -72535 4130 -72501
rect 4078 -72547 4130 -72535
<< pdiff >>
rect 31920 -30516 31978 -30504
rect 31920 -31092 31932 -30516
rect 31966 -31092 31978 -30516
rect 31920 -31104 31978 -31092
rect 32938 -30516 32996 -30504
rect 32938 -31092 32950 -30516
rect 32984 -31092 32996 -30516
rect 32938 -31104 32996 -31092
rect 33956 -30516 34014 -30504
rect 33956 -31092 33968 -30516
rect 34002 -31092 34014 -30516
rect 33956 -31104 34014 -31092
rect 34974 -30516 35032 -30504
rect 34974 -31092 34986 -30516
rect 35020 -31092 35032 -30516
rect 34974 -31104 35032 -31092
rect 35992 -30516 36050 -30504
rect 35992 -31092 36004 -30516
rect 36038 -31092 36050 -30516
rect 35992 -31104 36050 -31092
rect 37010 -30516 37068 -30504
rect 37010 -31092 37022 -30516
rect 37056 -31092 37068 -30516
rect 37010 -31104 37068 -31092
rect 38028 -30516 38086 -30504
rect 38028 -31092 38040 -30516
rect 38074 -31092 38086 -30516
rect 38028 -31104 38086 -31092
rect 39046 -30516 39104 -30504
rect 39046 -31092 39058 -30516
rect 39092 -31092 39104 -30516
rect 39046 -31104 39104 -31092
rect 40064 -30516 40122 -30504
rect 40064 -31092 40076 -30516
rect 40110 -31092 40122 -30516
rect 40064 -31104 40122 -31092
rect 41082 -30516 41140 -30504
rect 41082 -31092 41094 -30516
rect 41128 -31092 41140 -30516
rect 41082 -31104 41140 -31092
rect 42100 -30516 42158 -30504
rect 42100 -31092 42112 -30516
rect 42146 -31092 42158 -30516
rect 42100 -31104 42158 -31092
rect 43118 -30516 43176 -30504
rect 43118 -31092 43130 -30516
rect 43164 -31092 43176 -30516
rect 43118 -31104 43176 -31092
rect 44136 -30516 44194 -30504
rect 44136 -31092 44148 -30516
rect 44182 -31092 44194 -30516
rect 44136 -31104 44194 -31092
rect 45154 -30516 45212 -30504
rect 45154 -31092 45166 -30516
rect 45200 -31092 45212 -30516
rect 45154 -31104 45212 -31092
rect 46172 -30516 46230 -30504
rect 46172 -31092 46184 -30516
rect 46218 -31092 46230 -30516
rect 46172 -31104 46230 -31092
rect 47190 -30516 47248 -30504
rect 47190 -31092 47202 -30516
rect 47236 -31092 47248 -30516
rect 47190 -31104 47248 -31092
rect 48208 -30516 48266 -30504
rect 48208 -31092 48220 -30516
rect 48254 -31092 48266 -30516
rect 48208 -31104 48266 -31092
rect 31920 -31652 31978 -31640
rect 31920 -32228 31932 -31652
rect 31966 -32228 31978 -31652
rect 31920 -32240 31978 -32228
rect 32938 -31652 32996 -31640
rect 32938 -32228 32950 -31652
rect 32984 -32228 32996 -31652
rect 32938 -32240 32996 -32228
rect 33956 -31652 34014 -31640
rect 33956 -32228 33968 -31652
rect 34002 -32228 34014 -31652
rect 33956 -32240 34014 -32228
rect 34974 -31652 35032 -31640
rect 34974 -32228 34986 -31652
rect 35020 -32228 35032 -31652
rect 34974 -32240 35032 -32228
rect 35992 -31652 36050 -31640
rect 35992 -32228 36004 -31652
rect 36038 -32228 36050 -31652
rect 35992 -32240 36050 -32228
rect 37010 -31652 37068 -31640
rect 37010 -32228 37022 -31652
rect 37056 -32228 37068 -31652
rect 37010 -32240 37068 -32228
rect 38028 -31652 38086 -31640
rect 38028 -32228 38040 -31652
rect 38074 -32228 38086 -31652
rect 38028 -32240 38086 -32228
rect 39046 -31652 39104 -31640
rect 39046 -32228 39058 -31652
rect 39092 -32228 39104 -31652
rect 39046 -32240 39104 -32228
rect 40064 -31652 40122 -31640
rect 40064 -32228 40076 -31652
rect 40110 -32228 40122 -31652
rect 40064 -32240 40122 -32228
rect 41082 -31652 41140 -31640
rect 41082 -32228 41094 -31652
rect 41128 -32228 41140 -31652
rect 41082 -32240 41140 -32228
rect 42100 -31652 42158 -31640
rect 42100 -32228 42112 -31652
rect 42146 -32228 42158 -31652
rect 42100 -32240 42158 -32228
rect 43118 -31652 43176 -31640
rect 43118 -32228 43130 -31652
rect 43164 -32228 43176 -31652
rect 43118 -32240 43176 -32228
rect 44136 -31652 44194 -31640
rect 44136 -32228 44148 -31652
rect 44182 -32228 44194 -31652
rect 44136 -32240 44194 -32228
rect 45154 -31652 45212 -31640
rect 45154 -32228 45166 -31652
rect 45200 -32228 45212 -31652
rect 45154 -32240 45212 -32228
rect 46172 -31652 46230 -31640
rect 46172 -32228 46184 -31652
rect 46218 -32228 46230 -31652
rect 46172 -32240 46230 -32228
rect 47190 -31652 47248 -31640
rect 47190 -32228 47202 -31652
rect 47236 -32228 47248 -31652
rect 47190 -32240 47248 -32228
rect 48208 -31652 48266 -31640
rect 48208 -32228 48220 -31652
rect 48254 -32228 48266 -31652
rect 48208 -32240 48266 -32228
rect 31920 -32788 31978 -32776
rect 31920 -33364 31932 -32788
rect 31966 -33364 31978 -32788
rect 31920 -33376 31978 -33364
rect 32938 -32788 32996 -32776
rect 32938 -33364 32950 -32788
rect 32984 -33364 32996 -32788
rect 32938 -33376 32996 -33364
rect 33956 -32788 34014 -32776
rect 33956 -33364 33968 -32788
rect 34002 -33364 34014 -32788
rect 33956 -33376 34014 -33364
rect 34974 -32788 35032 -32776
rect 34974 -33364 34986 -32788
rect 35020 -33364 35032 -32788
rect 34974 -33376 35032 -33364
rect 35992 -32788 36050 -32776
rect 35992 -33364 36004 -32788
rect 36038 -33364 36050 -32788
rect 35992 -33376 36050 -33364
rect 37010 -32788 37068 -32776
rect 37010 -33364 37022 -32788
rect 37056 -33364 37068 -32788
rect 37010 -33376 37068 -33364
rect 38028 -32788 38086 -32776
rect 38028 -33364 38040 -32788
rect 38074 -33364 38086 -32788
rect 38028 -33376 38086 -33364
rect 39046 -32788 39104 -32776
rect 39046 -33364 39058 -32788
rect 39092 -33364 39104 -32788
rect 39046 -33376 39104 -33364
rect 40064 -32788 40122 -32776
rect 40064 -33364 40076 -32788
rect 40110 -33364 40122 -32788
rect 40064 -33376 40122 -33364
rect 41082 -32788 41140 -32776
rect 41082 -33364 41094 -32788
rect 41128 -33364 41140 -32788
rect 41082 -33376 41140 -33364
rect 42100 -32788 42158 -32776
rect 42100 -33364 42112 -32788
rect 42146 -33364 42158 -32788
rect 42100 -33376 42158 -33364
rect 43118 -32788 43176 -32776
rect 43118 -33364 43130 -32788
rect 43164 -33364 43176 -32788
rect 43118 -33376 43176 -33364
rect 44136 -32788 44194 -32776
rect 44136 -33364 44148 -32788
rect 44182 -33364 44194 -32788
rect 44136 -33376 44194 -33364
rect 45154 -32788 45212 -32776
rect 45154 -33364 45166 -32788
rect 45200 -33364 45212 -32788
rect 45154 -33376 45212 -33364
rect 46172 -32788 46230 -32776
rect 46172 -33364 46184 -32788
rect 46218 -33364 46230 -32788
rect 46172 -33376 46230 -33364
rect 47190 -32788 47248 -32776
rect 47190 -33364 47202 -32788
rect 47236 -33364 47248 -32788
rect 47190 -33376 47248 -33364
rect 48208 -32788 48266 -32776
rect 48208 -33364 48220 -32788
rect 48254 -33364 48266 -32788
rect 48208 -33376 48266 -33364
rect 33114 -34426 33172 -34414
rect 33114 -35002 33126 -34426
rect 33160 -35002 33172 -34426
rect 33114 -35014 33172 -35002
rect 34132 -34426 34190 -34414
rect 34132 -35002 34144 -34426
rect 34178 -35002 34190 -34426
rect 34132 -35014 34190 -35002
rect 35150 -34426 35208 -34414
rect 35150 -35002 35162 -34426
rect 35196 -35002 35208 -34426
rect 35150 -35014 35208 -35002
rect 36168 -34426 36226 -34414
rect 36168 -35002 36180 -34426
rect 36214 -35002 36226 -34426
rect 36168 -35014 36226 -35002
rect 37186 -34426 37244 -34414
rect 37186 -35002 37198 -34426
rect 37232 -35002 37244 -34426
rect 37186 -35014 37244 -35002
rect 38204 -34426 38262 -34414
rect 38204 -35002 38216 -34426
rect 38250 -35002 38262 -34426
rect 38204 -35014 38262 -35002
rect 39222 -34426 39280 -34414
rect 39222 -35002 39234 -34426
rect 39268 -35002 39280 -34426
rect 39222 -35014 39280 -35002
rect 40240 -34426 40298 -34414
rect 40240 -35002 40252 -34426
rect 40286 -35002 40298 -34426
rect 40240 -35014 40298 -35002
rect 41258 -34426 41316 -34414
rect 41258 -35002 41270 -34426
rect 41304 -35002 41316 -34426
rect 41258 -35014 41316 -35002
rect 42276 -34426 42334 -34414
rect 42276 -35002 42288 -34426
rect 42322 -35002 42334 -34426
rect 42276 -35014 42334 -35002
rect 43294 -34426 43352 -34414
rect 43294 -35002 43306 -34426
rect 43340 -35002 43352 -34426
rect 43294 -35014 43352 -35002
rect 44312 -34426 44370 -34414
rect 44312 -35002 44324 -34426
rect 44358 -35002 44370 -34426
rect 44312 -35014 44370 -35002
rect 45330 -34426 45388 -34414
rect 45330 -35002 45342 -34426
rect 45376 -35002 45388 -34426
rect 45330 -35014 45388 -35002
rect 46348 -34426 46406 -34414
rect 46348 -35002 46360 -34426
rect 46394 -35002 46406 -34426
rect 46348 -35014 46406 -35002
rect 47366 -34426 47424 -34414
rect 47366 -35002 47378 -34426
rect 47412 -35002 47424 -34426
rect 47366 -35014 47424 -35002
rect 33114 -35458 33172 -35446
rect 33114 -36034 33126 -35458
rect 33160 -36034 33172 -35458
rect 33114 -36046 33172 -36034
rect 34132 -35458 34190 -35446
rect 34132 -36034 34144 -35458
rect 34178 -36034 34190 -35458
rect 34132 -36046 34190 -36034
rect 35150 -35458 35208 -35446
rect 35150 -36034 35162 -35458
rect 35196 -36034 35208 -35458
rect 35150 -36046 35208 -36034
rect 36168 -35458 36226 -35446
rect 36168 -36034 36180 -35458
rect 36214 -36034 36226 -35458
rect 36168 -36046 36226 -36034
rect 37186 -35458 37244 -35446
rect 37186 -36034 37198 -35458
rect 37232 -36034 37244 -35458
rect 37186 -36046 37244 -36034
rect 38204 -35458 38262 -35446
rect 38204 -36034 38216 -35458
rect 38250 -36034 38262 -35458
rect 38204 -36046 38262 -36034
rect 39222 -35458 39280 -35446
rect 39222 -36034 39234 -35458
rect 39268 -36034 39280 -35458
rect 39222 -36046 39280 -36034
rect 40240 -35458 40298 -35446
rect 40240 -36034 40252 -35458
rect 40286 -36034 40298 -35458
rect 40240 -36046 40298 -36034
rect 41258 -35458 41316 -35446
rect 41258 -36034 41270 -35458
rect 41304 -36034 41316 -35458
rect 41258 -36046 41316 -36034
rect 42276 -35458 42334 -35446
rect 42276 -36034 42288 -35458
rect 42322 -36034 42334 -35458
rect 42276 -36046 42334 -36034
rect 43294 -35458 43352 -35446
rect 43294 -36034 43306 -35458
rect 43340 -36034 43352 -35458
rect 43294 -36046 43352 -36034
rect 44312 -35458 44370 -35446
rect 44312 -36034 44324 -35458
rect 44358 -36034 44370 -35458
rect 44312 -36046 44370 -36034
rect 45330 -35458 45388 -35446
rect 45330 -36034 45342 -35458
rect 45376 -36034 45388 -35458
rect 45330 -36046 45388 -36034
rect 46348 -35458 46406 -35446
rect 46348 -36034 46360 -35458
rect 46394 -36034 46406 -35458
rect 46348 -36046 46406 -36034
rect 47366 -35458 47424 -35446
rect 47366 -36034 47378 -35458
rect 47412 -36034 47424 -35458
rect 47366 -36046 47424 -36034
rect 32906 -37062 32964 -37050
rect 27602 -37166 27660 -37154
rect 27602 -37742 27614 -37166
rect 27648 -37742 27660 -37166
rect 27602 -37754 27660 -37742
rect 28620 -37166 28678 -37154
rect 28620 -37742 28632 -37166
rect 28666 -37742 28678 -37166
rect 28620 -37754 28678 -37742
rect 29638 -37166 29696 -37154
rect 29638 -37742 29650 -37166
rect 29684 -37742 29696 -37166
rect 29638 -37754 29696 -37742
rect 30656 -37166 30714 -37154
rect 30656 -37742 30668 -37166
rect 30702 -37742 30714 -37166
rect 30656 -37754 30714 -37742
rect 31674 -37166 31732 -37154
rect 31674 -37742 31686 -37166
rect 31720 -37742 31732 -37166
rect 32906 -37638 32918 -37062
rect 32952 -37638 32964 -37062
rect 32906 -37650 32964 -37638
rect 33924 -37062 33982 -37050
rect 33924 -37638 33936 -37062
rect 33970 -37638 33982 -37062
rect 33924 -37650 33982 -37638
rect 34942 -37062 35000 -37050
rect 34942 -37638 34954 -37062
rect 34988 -37638 35000 -37062
rect 34942 -37650 35000 -37638
rect 35960 -37062 36018 -37050
rect 35960 -37638 35972 -37062
rect 36006 -37638 36018 -37062
rect 35960 -37650 36018 -37638
rect 36978 -37062 37036 -37050
rect 36978 -37638 36990 -37062
rect 37024 -37638 37036 -37062
rect 36978 -37650 37036 -37638
rect 37996 -37062 38054 -37050
rect 37996 -37638 38008 -37062
rect 38042 -37638 38054 -37062
rect 37996 -37650 38054 -37638
rect 39014 -37062 39072 -37050
rect 39014 -37638 39026 -37062
rect 39060 -37638 39072 -37062
rect 39014 -37650 39072 -37638
rect 40032 -37062 40090 -37050
rect 40032 -37638 40044 -37062
rect 40078 -37638 40090 -37062
rect 40032 -37650 40090 -37638
rect 41050 -37062 41108 -37050
rect 41050 -37638 41062 -37062
rect 41096 -37638 41108 -37062
rect 41050 -37650 41108 -37638
rect 42068 -37062 42126 -37050
rect 42068 -37638 42080 -37062
rect 42114 -37638 42126 -37062
rect 42068 -37650 42126 -37638
rect 43086 -37062 43144 -37050
rect 43086 -37638 43098 -37062
rect 43132 -37638 43144 -37062
rect 43086 -37650 43144 -37638
rect 44104 -37062 44162 -37050
rect 44104 -37638 44116 -37062
rect 44150 -37638 44162 -37062
rect 44104 -37650 44162 -37638
rect 45122 -37062 45180 -37050
rect 45122 -37638 45134 -37062
rect 45168 -37638 45180 -37062
rect 45122 -37650 45180 -37638
rect 46140 -37062 46198 -37050
rect 46140 -37638 46152 -37062
rect 46186 -37638 46198 -37062
rect 46140 -37650 46198 -37638
rect 47158 -37062 47216 -37050
rect 47158 -37638 47170 -37062
rect 47204 -37638 47216 -37062
rect 47158 -37650 47216 -37638
rect 48176 -37062 48234 -37050
rect 48176 -37638 48188 -37062
rect 48222 -37638 48234 -37062
rect 48176 -37650 48234 -37638
rect 31674 -37754 31732 -37742
rect 27602 -38198 27660 -38186
rect 27602 -38774 27614 -38198
rect 27648 -38774 27660 -38198
rect 27602 -38786 27660 -38774
rect 28620 -38198 28678 -38186
rect 28620 -38774 28632 -38198
rect 28666 -38774 28678 -38198
rect 28620 -38786 28678 -38774
rect 29638 -38198 29696 -38186
rect 29638 -38774 29650 -38198
rect 29684 -38774 29696 -38198
rect 29638 -38786 29696 -38774
rect 30656 -38198 30714 -38186
rect 30656 -38774 30668 -38198
rect 30702 -38774 30714 -38198
rect 30656 -38786 30714 -38774
rect 31674 -38198 31732 -38186
rect 31674 -38774 31686 -38198
rect 31720 -38774 31732 -38198
rect 31674 -38786 31732 -38774
rect 32906 -38318 32964 -38306
rect 32906 -38894 32918 -38318
rect 32952 -38894 32964 -38318
rect 32906 -38906 32964 -38894
rect 33924 -38318 33982 -38306
rect 33924 -38894 33936 -38318
rect 33970 -38894 33982 -38318
rect 33924 -38906 33982 -38894
rect 34942 -38318 35000 -38306
rect 34942 -38894 34954 -38318
rect 34988 -38894 35000 -38318
rect 34942 -38906 35000 -38894
rect 35960 -38318 36018 -38306
rect 35960 -38894 35972 -38318
rect 36006 -38894 36018 -38318
rect 35960 -38906 36018 -38894
rect 36978 -38318 37036 -38306
rect 36978 -38894 36990 -38318
rect 37024 -38894 37036 -38318
rect 36978 -38906 37036 -38894
rect 37996 -38318 38054 -38306
rect 37996 -38894 38008 -38318
rect 38042 -38894 38054 -38318
rect 37996 -38906 38054 -38894
rect 39014 -38318 39072 -38306
rect 39014 -38894 39026 -38318
rect 39060 -38894 39072 -38318
rect 39014 -38906 39072 -38894
rect 40032 -38318 40090 -38306
rect 40032 -38894 40044 -38318
rect 40078 -38894 40090 -38318
rect 40032 -38906 40090 -38894
rect 41050 -38318 41108 -38306
rect 41050 -38894 41062 -38318
rect 41096 -38894 41108 -38318
rect 41050 -38906 41108 -38894
rect 42068 -38318 42126 -38306
rect 42068 -38894 42080 -38318
rect 42114 -38894 42126 -38318
rect 42068 -38906 42126 -38894
rect 43086 -38318 43144 -38306
rect 43086 -38894 43098 -38318
rect 43132 -38894 43144 -38318
rect 43086 -38906 43144 -38894
rect 44104 -38318 44162 -38306
rect 44104 -38894 44116 -38318
rect 44150 -38894 44162 -38318
rect 44104 -38906 44162 -38894
rect 45122 -38318 45180 -38306
rect 45122 -38894 45134 -38318
rect 45168 -38894 45180 -38318
rect 45122 -38906 45180 -38894
rect 46140 -38318 46198 -38306
rect 46140 -38894 46152 -38318
rect 46186 -38894 46198 -38318
rect 46140 -38906 46198 -38894
rect 47158 -38318 47216 -38306
rect 47158 -38894 47170 -38318
rect 47204 -38894 47216 -38318
rect 47158 -38906 47216 -38894
rect 48176 -38318 48234 -38306
rect 48176 -38894 48188 -38318
rect 48222 -38894 48234 -38318
rect 48176 -38906 48234 -38894
rect 27602 -39230 27660 -39218
rect 27602 -39806 27614 -39230
rect 27648 -39806 27660 -39230
rect 27602 -39818 27660 -39806
rect 28620 -39230 28678 -39218
rect 28620 -39806 28632 -39230
rect 28666 -39806 28678 -39230
rect 28620 -39818 28678 -39806
rect 29638 -39230 29696 -39218
rect 29638 -39806 29650 -39230
rect 29684 -39806 29696 -39230
rect 29638 -39818 29696 -39806
rect 30656 -39230 30714 -39218
rect 30656 -39806 30668 -39230
rect 30702 -39806 30714 -39230
rect 30656 -39818 30714 -39806
rect 31674 -39230 31732 -39218
rect 31674 -39806 31686 -39230
rect 31720 -39806 31732 -39230
rect 31674 -39818 31732 -39806
rect 32906 -39574 32964 -39562
rect 32906 -40150 32918 -39574
rect 32952 -40150 32964 -39574
rect 32906 -40162 32964 -40150
rect 33924 -39574 33982 -39562
rect 33924 -40150 33936 -39574
rect 33970 -40150 33982 -39574
rect 33924 -40162 33982 -40150
rect 34942 -39574 35000 -39562
rect 34942 -40150 34954 -39574
rect 34988 -40150 35000 -39574
rect 34942 -40162 35000 -40150
rect 35960 -39574 36018 -39562
rect 35960 -40150 35972 -39574
rect 36006 -40150 36018 -39574
rect 35960 -40162 36018 -40150
rect 36978 -39574 37036 -39562
rect 36978 -40150 36990 -39574
rect 37024 -40150 37036 -39574
rect 36978 -40162 37036 -40150
rect 37996 -39574 38054 -39562
rect 37996 -40150 38008 -39574
rect 38042 -40150 38054 -39574
rect 37996 -40162 38054 -40150
rect 39014 -39574 39072 -39562
rect 39014 -40150 39026 -39574
rect 39060 -40150 39072 -39574
rect 39014 -40162 39072 -40150
rect 40032 -39574 40090 -39562
rect 40032 -40150 40044 -39574
rect 40078 -40150 40090 -39574
rect 40032 -40162 40090 -40150
rect 41050 -39574 41108 -39562
rect 41050 -40150 41062 -39574
rect 41096 -40150 41108 -39574
rect 41050 -40162 41108 -40150
rect 42068 -39574 42126 -39562
rect 42068 -40150 42080 -39574
rect 42114 -40150 42126 -39574
rect 42068 -40162 42126 -40150
rect 43086 -39574 43144 -39562
rect 43086 -40150 43098 -39574
rect 43132 -40150 43144 -39574
rect 43086 -40162 43144 -40150
rect 44104 -39574 44162 -39562
rect 44104 -40150 44116 -39574
rect 44150 -40150 44162 -39574
rect 44104 -40162 44162 -40150
rect 45122 -39574 45180 -39562
rect 45122 -40150 45134 -39574
rect 45168 -40150 45180 -39574
rect 45122 -40162 45180 -40150
rect 46140 -39574 46198 -39562
rect 46140 -40150 46152 -39574
rect 46186 -40150 46198 -39574
rect 46140 -40162 46198 -40150
rect 47158 -39574 47216 -39562
rect 47158 -40150 47170 -39574
rect 47204 -40150 47216 -39574
rect 47158 -40162 47216 -40150
rect 48176 -39574 48234 -39562
rect 48176 -40150 48188 -39574
rect 48222 -40150 48234 -39574
rect 48176 -40162 48234 -40150
rect 27602 -40262 27660 -40250
rect 27602 -40838 27614 -40262
rect 27648 -40838 27660 -40262
rect 27602 -40850 27660 -40838
rect 28620 -40262 28678 -40250
rect 28620 -40838 28632 -40262
rect 28666 -40838 28678 -40262
rect 28620 -40850 28678 -40838
rect 29638 -40262 29696 -40250
rect 29638 -40838 29650 -40262
rect 29684 -40838 29696 -40262
rect 29638 -40850 29696 -40838
rect 30656 -40262 30714 -40250
rect 30656 -40838 30668 -40262
rect 30702 -40838 30714 -40262
rect 30656 -40850 30714 -40838
rect 31674 -40262 31732 -40250
rect 31674 -40838 31686 -40262
rect 31720 -40838 31732 -40262
rect 31674 -40850 31732 -40838
rect 32906 -40830 32964 -40818
rect 32906 -41406 32918 -40830
rect 32952 -41406 32964 -40830
rect 32906 -41418 32964 -41406
rect 33924 -40830 33982 -40818
rect 33924 -41406 33936 -40830
rect 33970 -41406 33982 -40830
rect 33924 -41418 33982 -41406
rect 34942 -40830 35000 -40818
rect 34942 -41406 34954 -40830
rect 34988 -41406 35000 -40830
rect 34942 -41418 35000 -41406
rect 35960 -40830 36018 -40818
rect 35960 -41406 35972 -40830
rect 36006 -41406 36018 -40830
rect 35960 -41418 36018 -41406
rect 36978 -40830 37036 -40818
rect 36978 -41406 36990 -40830
rect 37024 -41406 37036 -40830
rect 36978 -41418 37036 -41406
rect 37996 -40830 38054 -40818
rect 37996 -41406 38008 -40830
rect 38042 -41406 38054 -40830
rect 37996 -41418 38054 -41406
rect 39014 -40830 39072 -40818
rect 39014 -41406 39026 -40830
rect 39060 -41406 39072 -40830
rect 39014 -41418 39072 -41406
rect 40032 -40830 40090 -40818
rect 40032 -41406 40044 -40830
rect 40078 -41406 40090 -40830
rect 40032 -41418 40090 -41406
rect 41050 -40830 41108 -40818
rect 41050 -41406 41062 -40830
rect 41096 -41406 41108 -40830
rect 41050 -41418 41108 -41406
rect 42068 -40830 42126 -40818
rect 42068 -41406 42080 -40830
rect 42114 -41406 42126 -40830
rect 42068 -41418 42126 -41406
rect 43086 -40830 43144 -40818
rect 43086 -41406 43098 -40830
rect 43132 -41406 43144 -40830
rect 43086 -41418 43144 -41406
rect 44104 -40830 44162 -40818
rect 44104 -41406 44116 -40830
rect 44150 -41406 44162 -40830
rect 44104 -41418 44162 -41406
rect 45122 -40830 45180 -40818
rect 45122 -41406 45134 -40830
rect 45168 -41406 45180 -40830
rect 45122 -41418 45180 -41406
rect 46140 -40830 46198 -40818
rect 46140 -41406 46152 -40830
rect 46186 -41406 46198 -40830
rect 46140 -41418 46198 -41406
rect 47158 -40830 47216 -40818
rect 47158 -41406 47170 -40830
rect 47204 -41406 47216 -40830
rect 47158 -41418 47216 -41406
rect 48176 -40830 48234 -40818
rect 48176 -41406 48188 -40830
rect 48222 -41406 48234 -40830
rect 48176 -41418 48234 -41406
rect 52430 -39692 52488 -39680
rect 52430 -39868 52442 -39692
rect 52476 -39868 52488 -39692
rect 52430 -39880 52488 -39868
rect 52888 -39692 52946 -39680
rect 52888 -39868 52900 -39692
rect 52934 -39868 52946 -39692
rect 52888 -39880 52946 -39868
rect 53346 -39692 53404 -39680
rect 53346 -39868 53358 -39692
rect 53392 -39868 53404 -39692
rect 53346 -39880 53404 -39868
rect 53804 -39692 53862 -39680
rect 53804 -39868 53816 -39692
rect 53850 -39868 53862 -39692
rect 53804 -39880 53862 -39868
rect 54262 -39692 54320 -39680
rect 54262 -39868 54274 -39692
rect 54308 -39868 54320 -39692
rect 54262 -39880 54320 -39868
rect 54720 -39692 54778 -39680
rect 54720 -39868 54732 -39692
rect 54766 -39868 54778 -39692
rect 54720 -39880 54778 -39868
rect 55178 -39692 55236 -39680
rect 55178 -39868 55190 -39692
rect 55224 -39868 55236 -39692
rect 55178 -39880 55236 -39868
rect 52489 -40575 52547 -40563
rect 52489 -40951 52501 -40575
rect 52535 -40951 52547 -40575
rect 52489 -40963 52547 -40951
rect 52747 -40575 52805 -40563
rect 52747 -40951 52759 -40575
rect 52793 -40951 52805 -40575
rect 52747 -40963 52805 -40951
rect 53005 -40575 53063 -40563
rect 53005 -40951 53017 -40575
rect 53051 -40951 53063 -40575
rect 53005 -40963 53063 -40951
rect 53263 -40575 53321 -40563
rect 53263 -40951 53275 -40575
rect 53309 -40951 53321 -40575
rect 53263 -40963 53321 -40951
rect 53521 -40575 53579 -40563
rect 53521 -40951 53533 -40575
rect 53567 -40951 53579 -40575
rect 53521 -40963 53579 -40951
rect 53779 -40575 53837 -40563
rect 53779 -40951 53791 -40575
rect 53825 -40951 53837 -40575
rect 53779 -40963 53837 -40951
rect 54037 -40575 54095 -40563
rect 54037 -40951 54049 -40575
rect 54083 -40951 54095 -40575
rect 54037 -40963 54095 -40951
rect 54295 -40575 54353 -40563
rect 54295 -40951 54307 -40575
rect 54341 -40951 54353 -40575
rect 54295 -40963 54353 -40951
rect 54553 -40575 54611 -40563
rect 54553 -40951 54565 -40575
rect 54599 -40951 54611 -40575
rect 54553 -40963 54611 -40951
rect 54811 -40575 54869 -40563
rect 54811 -40951 54823 -40575
rect 54857 -40951 54869 -40575
rect 54811 -40963 54869 -40951
rect 55069 -40575 55127 -40563
rect 55069 -40951 55081 -40575
rect 55115 -40951 55127 -40575
rect 55069 -40963 55127 -40951
rect 52489 -41435 52547 -41423
rect 52489 -41811 52501 -41435
rect 52535 -41811 52547 -41435
rect 52489 -41823 52547 -41811
rect 52747 -41435 52805 -41423
rect 52747 -41811 52759 -41435
rect 52793 -41811 52805 -41435
rect 52747 -41823 52805 -41811
rect 53005 -41435 53063 -41423
rect 53005 -41811 53017 -41435
rect 53051 -41811 53063 -41435
rect 53005 -41823 53063 -41811
rect 53263 -41435 53321 -41423
rect 53263 -41811 53275 -41435
rect 53309 -41811 53321 -41435
rect 53263 -41823 53321 -41811
rect 53521 -41435 53579 -41423
rect 53521 -41811 53533 -41435
rect 53567 -41811 53579 -41435
rect 53521 -41823 53579 -41811
rect 53779 -41435 53837 -41423
rect 53779 -41811 53791 -41435
rect 53825 -41811 53837 -41435
rect 53779 -41823 53837 -41811
rect 54037 -41435 54095 -41423
rect 54037 -41811 54049 -41435
rect 54083 -41811 54095 -41435
rect 54037 -41823 54095 -41811
rect 54295 -41435 54353 -41423
rect 54295 -41811 54307 -41435
rect 54341 -41811 54353 -41435
rect 54295 -41823 54353 -41811
rect 54553 -41435 54611 -41423
rect 54553 -41811 54565 -41435
rect 54599 -41811 54611 -41435
rect 54553 -41823 54611 -41811
rect 54811 -41435 54869 -41423
rect 54811 -41811 54823 -41435
rect 54857 -41811 54869 -41435
rect 54811 -41823 54869 -41811
rect 55069 -41435 55127 -41423
rect 55069 -41811 55081 -41435
rect 55115 -41811 55127 -41435
rect 55069 -41823 55127 -41811
rect 56058 -39892 56116 -39880
rect 56058 -40268 56070 -39892
rect 56104 -40268 56116 -39892
rect 56058 -40280 56116 -40268
rect 56316 -39892 56374 -39880
rect 56316 -40268 56328 -39892
rect 56362 -40268 56374 -39892
rect 56316 -40280 56374 -40268
rect 56574 -39892 56632 -39880
rect 56574 -40268 56586 -39892
rect 56620 -40268 56632 -39892
rect 56574 -40280 56632 -40268
rect 56832 -39892 56890 -39880
rect 56832 -40268 56844 -39892
rect 56878 -40268 56890 -39892
rect 56832 -40280 56890 -40268
rect 57090 -39892 57148 -39880
rect 57090 -40268 57102 -39892
rect 57136 -40268 57148 -39892
rect 57090 -40280 57148 -40268
rect 57348 -39892 57406 -39880
rect 57348 -40268 57360 -39892
rect 57394 -40268 57406 -39892
rect 57348 -40280 57406 -40268
rect 57606 -39892 57664 -39880
rect 57606 -40268 57618 -39892
rect 57652 -40268 57664 -39892
rect 57606 -40280 57664 -40268
rect 57864 -39892 57922 -39880
rect 57864 -40268 57876 -39892
rect 57910 -40268 57922 -39892
rect 57864 -40280 57922 -40268
rect 56058 -40752 56116 -40740
rect 56058 -41128 56070 -40752
rect 56104 -41128 56116 -40752
rect 56058 -41140 56116 -41128
rect 56316 -40752 56374 -40740
rect 56316 -41128 56328 -40752
rect 56362 -41128 56374 -40752
rect 56316 -41140 56374 -41128
rect 56574 -40752 56632 -40740
rect 56574 -41128 56586 -40752
rect 56620 -41128 56632 -40752
rect 56574 -41140 56632 -41128
rect 56832 -40752 56890 -40740
rect 56832 -41128 56844 -40752
rect 56878 -41128 56890 -40752
rect 56832 -41140 56890 -41128
rect 57090 -40752 57148 -40740
rect 57090 -41128 57102 -40752
rect 57136 -41128 57148 -40752
rect 57090 -41140 57148 -41128
rect 57348 -40752 57406 -40740
rect 57348 -41128 57360 -40752
rect 57394 -41128 57406 -40752
rect 57348 -41140 57406 -41128
rect 57606 -40752 57664 -40740
rect 57606 -41128 57618 -40752
rect 57652 -41128 57664 -40752
rect 57606 -41140 57664 -41128
rect 57864 -40752 57922 -40740
rect 57864 -41128 57876 -40752
rect 57910 -41128 57922 -40752
rect 57864 -41140 57922 -41128
rect 56172 -41651 56224 -41639
rect 56172 -41685 56180 -41651
rect 56214 -41685 56224 -41651
rect 56172 -41719 56224 -41685
rect 56172 -41753 56180 -41719
rect 56214 -41753 56224 -41719
rect 56172 -41787 56224 -41753
rect 56172 -41821 56180 -41787
rect 56214 -41821 56224 -41787
rect 56172 -41839 56224 -41821
rect 56254 -41651 56306 -41639
rect 56254 -41685 56264 -41651
rect 56298 -41685 56306 -41651
rect 56254 -41719 56306 -41685
rect 56254 -41753 56264 -41719
rect 56298 -41753 56306 -41719
rect 56254 -41787 56306 -41753
rect 56254 -41821 56264 -41787
rect 56298 -41821 56306 -41787
rect 56254 -41839 56306 -41821
rect 56448 -41651 56500 -41639
rect 56448 -41685 56456 -41651
rect 56490 -41685 56500 -41651
rect 56448 -41719 56500 -41685
rect 56448 -41753 56456 -41719
rect 56490 -41753 56500 -41719
rect 56448 -41787 56500 -41753
rect 56448 -41821 56456 -41787
rect 56490 -41821 56500 -41787
rect 56448 -41839 56500 -41821
rect 56530 -41651 56582 -41639
rect 56530 -41685 56540 -41651
rect 56574 -41685 56582 -41651
rect 56530 -41719 56582 -41685
rect 56530 -41753 56540 -41719
rect 56574 -41753 56582 -41719
rect 56530 -41787 56582 -41753
rect 56530 -41821 56540 -41787
rect 56574 -41821 56582 -41787
rect 56530 -41839 56582 -41821
rect 56687 -41651 56739 -41639
rect 56687 -41685 56695 -41651
rect 56729 -41685 56739 -41651
rect 56687 -41719 56739 -41685
rect 56687 -41753 56695 -41719
rect 56729 -41753 56739 -41719
rect 56687 -41787 56739 -41753
rect 56687 -41821 56695 -41787
rect 56729 -41821 56739 -41787
rect 56687 -41839 56739 -41821
rect 56769 -41651 56823 -41639
rect 56769 -41685 56779 -41651
rect 56813 -41685 56823 -41651
rect 56769 -41719 56823 -41685
rect 56769 -41753 56779 -41719
rect 56813 -41753 56823 -41719
rect 56769 -41787 56823 -41753
rect 56769 -41821 56779 -41787
rect 56813 -41821 56823 -41787
rect 56769 -41839 56823 -41821
rect 56853 -41651 56905 -41639
rect 56853 -41685 56863 -41651
rect 56897 -41685 56905 -41651
rect 56853 -41719 56905 -41685
rect 56853 -41753 56863 -41719
rect 56897 -41753 56905 -41719
rect 56853 -41787 56905 -41753
rect 56853 -41821 56863 -41787
rect 56897 -41821 56905 -41787
rect 56853 -41839 56905 -41821
rect 57145 -41651 57197 -41639
rect 57145 -41685 57153 -41651
rect 57187 -41685 57197 -41651
rect 57145 -41719 57197 -41685
rect 57145 -41753 57153 -41719
rect 57187 -41753 57197 -41719
rect 57145 -41787 57197 -41753
rect 57145 -41821 57153 -41787
rect 57187 -41821 57197 -41787
rect 57145 -41839 57197 -41821
rect 57227 -41651 57281 -41639
rect 57227 -41685 57237 -41651
rect 57271 -41685 57281 -41651
rect 57227 -41719 57281 -41685
rect 57227 -41753 57237 -41719
rect 57271 -41753 57281 -41719
rect 57227 -41787 57281 -41753
rect 57227 -41821 57237 -41787
rect 57271 -41821 57281 -41787
rect 57227 -41839 57281 -41821
rect 57311 -41651 57363 -41639
rect 57311 -41685 57321 -41651
rect 57355 -41685 57363 -41651
rect 57311 -41719 57363 -41685
rect 57311 -41753 57321 -41719
rect 57355 -41753 57363 -41719
rect 57311 -41787 57363 -41753
rect 57311 -41821 57321 -41787
rect 57355 -41821 57363 -41787
rect 57311 -41839 57363 -41821
rect 57468 -41651 57520 -41639
rect 57468 -41685 57476 -41651
rect 57510 -41685 57520 -41651
rect 57468 -41719 57520 -41685
rect 57468 -41753 57476 -41719
rect 57510 -41753 57520 -41719
rect 57468 -41787 57520 -41753
rect 57468 -41821 57476 -41787
rect 57510 -41821 57520 -41787
rect 57468 -41839 57520 -41821
rect 57550 -41651 57602 -41639
rect 57550 -41685 57560 -41651
rect 57594 -41685 57602 -41651
rect 57550 -41719 57602 -41685
rect 57550 -41753 57560 -41719
rect 57594 -41753 57602 -41719
rect 57550 -41787 57602 -41753
rect 57550 -41821 57560 -41787
rect 57594 -41821 57602 -41787
rect 57550 -41839 57602 -41821
rect 57744 -41651 57796 -41639
rect 57744 -41685 57752 -41651
rect 57786 -41685 57796 -41651
rect 57744 -41719 57796 -41685
rect 57744 -41753 57752 -41719
rect 57786 -41753 57796 -41719
rect 57744 -41787 57796 -41753
rect 57744 -41821 57752 -41787
rect 57786 -41821 57796 -41787
rect 57744 -41839 57796 -41821
rect 57826 -41651 57878 -41639
rect 57826 -41685 57836 -41651
rect 57870 -41685 57878 -41651
rect 57826 -41719 57878 -41685
rect 57826 -41753 57836 -41719
rect 57870 -41753 57878 -41719
rect 57826 -41787 57878 -41753
rect 57826 -41821 57836 -41787
rect 57870 -41821 57878 -41787
rect 57826 -41839 57878 -41821
rect 54206 -42606 54264 -42594
rect 54206 -42782 54218 -42606
rect 54252 -42782 54264 -42606
rect 54206 -42794 54264 -42782
rect 54334 -42606 54392 -42594
rect 54334 -42782 54346 -42606
rect 54380 -42782 54392 -42606
rect 54334 -42794 54392 -42782
rect 54462 -42606 54520 -42594
rect 54462 -42782 54474 -42606
rect 54508 -42782 54520 -42606
rect 54462 -42794 54520 -42782
rect 54590 -42606 54648 -42594
rect 54590 -42782 54602 -42606
rect 54636 -42782 54648 -42606
rect 54590 -42794 54648 -42782
rect 54718 -42606 54776 -42594
rect 54718 -42782 54730 -42606
rect 54764 -42782 54776 -42606
rect 54718 -42794 54776 -42782
rect 54846 -42606 54904 -42594
rect 54846 -42782 54858 -42606
rect 54892 -42782 54904 -42606
rect 54846 -42794 54904 -42782
rect 54974 -42606 55032 -42594
rect 54974 -42782 54986 -42606
rect 55020 -42782 55032 -42606
rect 54974 -42794 55032 -42782
rect 55102 -42606 55160 -42594
rect 55102 -42782 55114 -42606
rect 55148 -42782 55160 -42606
rect 55102 -42794 55160 -42782
rect 55230 -42606 55288 -42594
rect 55230 -42782 55242 -42606
rect 55276 -42782 55288 -42606
rect 55230 -42794 55288 -42782
rect 55358 -42606 55416 -42594
rect 55358 -42782 55370 -42606
rect 55404 -42782 55416 -42606
rect 55358 -42794 55416 -42782
rect 10398 -56934 10456 -56922
rect 10398 -57310 10410 -56934
rect 10444 -57310 10456 -56934
rect 10398 -57322 10456 -57310
rect 10656 -56934 10714 -56922
rect 10656 -57310 10668 -56934
rect 10702 -57310 10714 -56934
rect 10656 -57322 10714 -57310
rect 10914 -56934 10972 -56922
rect 10914 -57310 10926 -56934
rect 10960 -57310 10972 -56934
rect 10914 -57322 10972 -57310
rect 11172 -56934 11230 -56922
rect 11172 -57310 11184 -56934
rect 11218 -57310 11230 -56934
rect 11172 -57322 11230 -57310
rect 11430 -56934 11488 -56922
rect 11430 -57310 11442 -56934
rect 11476 -57310 11488 -56934
rect 11430 -57322 11488 -57310
rect 11688 -56934 11746 -56922
rect 11688 -57310 11700 -56934
rect 11734 -57310 11746 -56934
rect 11688 -57322 11746 -57310
rect 11946 -56934 12004 -56922
rect 11946 -57310 11958 -56934
rect 11992 -57310 12004 -56934
rect 11946 -57322 12004 -57310
rect 12254 -57317 12306 -57305
rect 12254 -57351 12262 -57317
rect 12296 -57351 12306 -57317
rect 12254 -57385 12306 -57351
rect 12254 -57419 12262 -57385
rect 12296 -57419 12306 -57385
rect 12254 -57453 12306 -57419
rect 12254 -57487 12262 -57453
rect 12296 -57487 12306 -57453
rect 12254 -57505 12306 -57487
rect 12336 -57317 12388 -57305
rect 12336 -57351 12346 -57317
rect 12380 -57351 12388 -57317
rect 12336 -57385 12388 -57351
rect 12336 -57419 12346 -57385
rect 12380 -57419 12388 -57385
rect 12336 -57453 12388 -57419
rect 12336 -57487 12346 -57453
rect 12380 -57487 12388 -57453
rect 12336 -57505 12388 -57487
rect -28004 -67341 -27952 -67329
rect -28004 -67375 -27996 -67341
rect -27962 -67375 -27952 -67341
rect -28004 -67409 -27952 -67375
rect -28004 -67443 -27996 -67409
rect -27962 -67443 -27952 -67409
rect -28004 -67477 -27952 -67443
rect -28004 -67511 -27996 -67477
rect -27962 -67511 -27952 -67477
rect -28004 -67529 -27952 -67511
rect -27922 -67341 -27870 -67329
rect -27922 -67375 -27912 -67341
rect -27878 -67375 -27870 -67341
rect -27922 -67409 -27870 -67375
rect -27922 -67443 -27912 -67409
rect -27878 -67443 -27870 -67409
rect -27922 -67477 -27870 -67443
rect -27922 -67511 -27912 -67477
rect -27878 -67511 -27870 -67477
rect -27922 -67529 -27870 -67511
rect -27349 -65637 -27291 -65625
rect -27349 -66013 -27337 -65637
rect -27303 -66013 -27291 -65637
rect -27349 -66025 -27291 -66013
rect -27091 -65637 -27033 -65625
rect -27091 -66013 -27079 -65637
rect -27045 -66013 -27033 -65637
rect -27091 -66025 -27033 -66013
rect -26833 -65637 -26775 -65625
rect -26833 -66013 -26821 -65637
rect -26787 -66013 -26775 -65637
rect -26833 -66025 -26775 -66013
rect -26575 -65637 -26517 -65625
rect -26575 -66013 -26563 -65637
rect -26529 -66013 -26517 -65637
rect -26575 -66025 -26517 -66013
rect -26317 -65637 -26259 -65625
rect -26317 -66013 -26305 -65637
rect -26271 -66013 -26259 -65637
rect -26317 -66025 -26259 -66013
rect -26059 -65637 -26001 -65625
rect -26059 -66013 -26047 -65637
rect -26013 -66013 -26001 -65637
rect -26059 -66025 -26001 -66013
rect -25801 -65637 -25743 -65625
rect -25801 -66013 -25789 -65637
rect -25755 -66013 -25743 -65637
rect -25801 -66025 -25743 -66013
rect -27349 -66497 -27291 -66485
rect -27349 -66873 -27337 -66497
rect -27303 -66873 -27291 -66497
rect -27349 -66885 -27291 -66873
rect -27091 -66497 -27033 -66485
rect -27091 -66873 -27079 -66497
rect -27045 -66873 -27033 -66497
rect -27091 -66885 -27033 -66873
rect -26833 -66497 -26775 -66485
rect -26833 -66873 -26821 -66497
rect -26787 -66873 -26775 -66497
rect -26833 -66885 -26775 -66873
rect -26575 -66497 -26517 -66485
rect -26575 -66873 -26563 -66497
rect -26529 -66873 -26517 -66497
rect -26575 -66885 -26517 -66873
rect -26317 -66497 -26259 -66485
rect -26317 -66873 -26305 -66497
rect -26271 -66873 -26259 -66497
rect -26317 -66885 -26259 -66873
rect -26059 -66497 -26001 -66485
rect -26059 -66873 -26047 -66497
rect -26013 -66873 -26001 -66497
rect -26059 -66885 -26001 -66873
rect -25801 -66497 -25743 -66485
rect -25801 -66873 -25789 -66497
rect -25755 -66873 -25743 -66497
rect -25801 -66885 -25743 -66873
rect -24004 -67341 -23952 -67329
rect -24004 -67375 -23996 -67341
rect -23962 -67375 -23952 -67341
rect -24004 -67409 -23952 -67375
rect -24004 -67443 -23996 -67409
rect -23962 -67443 -23952 -67409
rect -24004 -67477 -23952 -67443
rect -24004 -67511 -23996 -67477
rect -23962 -67511 -23952 -67477
rect -24004 -67529 -23952 -67511
rect -23922 -67341 -23870 -67329
rect -23922 -67375 -23912 -67341
rect -23878 -67375 -23870 -67341
rect -23922 -67409 -23870 -67375
rect -23922 -67443 -23912 -67409
rect -23878 -67443 -23870 -67409
rect -23922 -67477 -23870 -67443
rect -23922 -67511 -23912 -67477
rect -23878 -67511 -23870 -67477
rect -23922 -67529 -23870 -67511
rect -23349 -65637 -23291 -65625
rect -23349 -66013 -23337 -65637
rect -23303 -66013 -23291 -65637
rect -23349 -66025 -23291 -66013
rect -23091 -65637 -23033 -65625
rect -23091 -66013 -23079 -65637
rect -23045 -66013 -23033 -65637
rect -23091 -66025 -23033 -66013
rect -22833 -65637 -22775 -65625
rect -22833 -66013 -22821 -65637
rect -22787 -66013 -22775 -65637
rect -22833 -66025 -22775 -66013
rect -22575 -65637 -22517 -65625
rect -22575 -66013 -22563 -65637
rect -22529 -66013 -22517 -65637
rect -22575 -66025 -22517 -66013
rect -22317 -65637 -22259 -65625
rect -22317 -66013 -22305 -65637
rect -22271 -66013 -22259 -65637
rect -22317 -66025 -22259 -66013
rect -22059 -65637 -22001 -65625
rect -22059 -66013 -22047 -65637
rect -22013 -66013 -22001 -65637
rect -22059 -66025 -22001 -66013
rect -21801 -65637 -21743 -65625
rect -21801 -66013 -21789 -65637
rect -21755 -66013 -21743 -65637
rect -21801 -66025 -21743 -66013
rect -23349 -66497 -23291 -66485
rect -23349 -66873 -23337 -66497
rect -23303 -66873 -23291 -66497
rect -23349 -66885 -23291 -66873
rect -23091 -66497 -23033 -66485
rect -23091 -66873 -23079 -66497
rect -23045 -66873 -23033 -66497
rect -23091 -66885 -23033 -66873
rect -22833 -66497 -22775 -66485
rect -22833 -66873 -22821 -66497
rect -22787 -66873 -22775 -66497
rect -22833 -66885 -22775 -66873
rect -22575 -66497 -22517 -66485
rect -22575 -66873 -22563 -66497
rect -22529 -66873 -22517 -66497
rect -22575 -66885 -22517 -66873
rect -22317 -66497 -22259 -66485
rect -22317 -66873 -22305 -66497
rect -22271 -66873 -22259 -66497
rect -22317 -66885 -22259 -66873
rect -22059 -66497 -22001 -66485
rect -22059 -66873 -22047 -66497
rect -22013 -66873 -22001 -66497
rect -22059 -66885 -22001 -66873
rect -21801 -66497 -21743 -66485
rect -21801 -66873 -21789 -66497
rect -21755 -66873 -21743 -66497
rect -21801 -66885 -21743 -66873
rect -20004 -67341 -19952 -67329
rect -20004 -67375 -19996 -67341
rect -19962 -67375 -19952 -67341
rect -20004 -67409 -19952 -67375
rect -20004 -67443 -19996 -67409
rect -19962 -67443 -19952 -67409
rect -20004 -67477 -19952 -67443
rect -20004 -67511 -19996 -67477
rect -19962 -67511 -19952 -67477
rect -20004 -67529 -19952 -67511
rect -19922 -67341 -19870 -67329
rect -19922 -67375 -19912 -67341
rect -19878 -67375 -19870 -67341
rect -19922 -67409 -19870 -67375
rect -19922 -67443 -19912 -67409
rect -19878 -67443 -19870 -67409
rect -19922 -67477 -19870 -67443
rect -19922 -67511 -19912 -67477
rect -19878 -67511 -19870 -67477
rect -19922 -67529 -19870 -67511
rect -19349 -65637 -19291 -65625
rect -19349 -66013 -19337 -65637
rect -19303 -66013 -19291 -65637
rect -19349 -66025 -19291 -66013
rect -19091 -65637 -19033 -65625
rect -19091 -66013 -19079 -65637
rect -19045 -66013 -19033 -65637
rect -19091 -66025 -19033 -66013
rect -18833 -65637 -18775 -65625
rect -18833 -66013 -18821 -65637
rect -18787 -66013 -18775 -65637
rect -18833 -66025 -18775 -66013
rect -18575 -65637 -18517 -65625
rect -18575 -66013 -18563 -65637
rect -18529 -66013 -18517 -65637
rect -18575 -66025 -18517 -66013
rect -18317 -65637 -18259 -65625
rect -18317 -66013 -18305 -65637
rect -18271 -66013 -18259 -65637
rect -18317 -66025 -18259 -66013
rect -18059 -65637 -18001 -65625
rect -18059 -66013 -18047 -65637
rect -18013 -66013 -18001 -65637
rect -18059 -66025 -18001 -66013
rect -17801 -65637 -17743 -65625
rect -17801 -66013 -17789 -65637
rect -17755 -66013 -17743 -65637
rect -17801 -66025 -17743 -66013
rect -19349 -66497 -19291 -66485
rect -19349 -66873 -19337 -66497
rect -19303 -66873 -19291 -66497
rect -19349 -66885 -19291 -66873
rect -19091 -66497 -19033 -66485
rect -19091 -66873 -19079 -66497
rect -19045 -66873 -19033 -66497
rect -19091 -66885 -19033 -66873
rect -18833 -66497 -18775 -66485
rect -18833 -66873 -18821 -66497
rect -18787 -66873 -18775 -66497
rect -18833 -66885 -18775 -66873
rect -18575 -66497 -18517 -66485
rect -18575 -66873 -18563 -66497
rect -18529 -66873 -18517 -66497
rect -18575 -66885 -18517 -66873
rect -18317 -66497 -18259 -66485
rect -18317 -66873 -18305 -66497
rect -18271 -66873 -18259 -66497
rect -18317 -66885 -18259 -66873
rect -18059 -66497 -18001 -66485
rect -18059 -66873 -18047 -66497
rect -18013 -66873 -18001 -66497
rect -18059 -66885 -18001 -66873
rect -17801 -66497 -17743 -66485
rect -17801 -66873 -17789 -66497
rect -17755 -66873 -17743 -66497
rect -17801 -66885 -17743 -66873
rect -16004 -67341 -15952 -67329
rect -16004 -67375 -15996 -67341
rect -15962 -67375 -15952 -67341
rect -16004 -67409 -15952 -67375
rect -16004 -67443 -15996 -67409
rect -15962 -67443 -15952 -67409
rect -16004 -67477 -15952 -67443
rect -16004 -67511 -15996 -67477
rect -15962 -67511 -15952 -67477
rect -16004 -67529 -15952 -67511
rect -15922 -67341 -15870 -67329
rect -15922 -67375 -15912 -67341
rect -15878 -67375 -15870 -67341
rect -15922 -67409 -15870 -67375
rect -15922 -67443 -15912 -67409
rect -15878 -67443 -15870 -67409
rect -15922 -67477 -15870 -67443
rect -15922 -67511 -15912 -67477
rect -15878 -67511 -15870 -67477
rect -15922 -67529 -15870 -67511
rect -15349 -65637 -15291 -65625
rect -15349 -66013 -15337 -65637
rect -15303 -66013 -15291 -65637
rect -15349 -66025 -15291 -66013
rect -15091 -65637 -15033 -65625
rect -15091 -66013 -15079 -65637
rect -15045 -66013 -15033 -65637
rect -15091 -66025 -15033 -66013
rect -14833 -65637 -14775 -65625
rect -14833 -66013 -14821 -65637
rect -14787 -66013 -14775 -65637
rect -14833 -66025 -14775 -66013
rect -14575 -65637 -14517 -65625
rect -14575 -66013 -14563 -65637
rect -14529 -66013 -14517 -65637
rect -14575 -66025 -14517 -66013
rect -14317 -65637 -14259 -65625
rect -14317 -66013 -14305 -65637
rect -14271 -66013 -14259 -65637
rect -14317 -66025 -14259 -66013
rect -14059 -65637 -14001 -65625
rect -14059 -66013 -14047 -65637
rect -14013 -66013 -14001 -65637
rect -14059 -66025 -14001 -66013
rect -13801 -65637 -13743 -65625
rect -13801 -66013 -13789 -65637
rect -13755 -66013 -13743 -65637
rect -13801 -66025 -13743 -66013
rect -15349 -66497 -15291 -66485
rect -15349 -66873 -15337 -66497
rect -15303 -66873 -15291 -66497
rect -15349 -66885 -15291 -66873
rect -15091 -66497 -15033 -66485
rect -15091 -66873 -15079 -66497
rect -15045 -66873 -15033 -66497
rect -15091 -66885 -15033 -66873
rect -14833 -66497 -14775 -66485
rect -14833 -66873 -14821 -66497
rect -14787 -66873 -14775 -66497
rect -14833 -66885 -14775 -66873
rect -14575 -66497 -14517 -66485
rect -14575 -66873 -14563 -66497
rect -14529 -66873 -14517 -66497
rect -14575 -66885 -14517 -66873
rect -14317 -66497 -14259 -66485
rect -14317 -66873 -14305 -66497
rect -14271 -66873 -14259 -66497
rect -14317 -66885 -14259 -66873
rect -14059 -66497 -14001 -66485
rect -14059 -66873 -14047 -66497
rect -14013 -66873 -14001 -66497
rect -14059 -66885 -14001 -66873
rect -13801 -66497 -13743 -66485
rect -13801 -66873 -13789 -66497
rect -13755 -66873 -13743 -66497
rect -13801 -66885 -13743 -66873
rect -12004 -67341 -11952 -67329
rect -12004 -67375 -11996 -67341
rect -11962 -67375 -11952 -67341
rect -12004 -67409 -11952 -67375
rect -12004 -67443 -11996 -67409
rect -11962 -67443 -11952 -67409
rect -12004 -67477 -11952 -67443
rect -12004 -67511 -11996 -67477
rect -11962 -67511 -11952 -67477
rect -12004 -67529 -11952 -67511
rect -11922 -67341 -11870 -67329
rect -11922 -67375 -11912 -67341
rect -11878 -67375 -11870 -67341
rect -11922 -67409 -11870 -67375
rect -11922 -67443 -11912 -67409
rect -11878 -67443 -11870 -67409
rect -11922 -67477 -11870 -67443
rect -11922 -67511 -11912 -67477
rect -11878 -67511 -11870 -67477
rect -11922 -67529 -11870 -67511
rect -11349 -65637 -11291 -65625
rect -11349 -66013 -11337 -65637
rect -11303 -66013 -11291 -65637
rect -11349 -66025 -11291 -66013
rect -11091 -65637 -11033 -65625
rect -11091 -66013 -11079 -65637
rect -11045 -66013 -11033 -65637
rect -11091 -66025 -11033 -66013
rect -10833 -65637 -10775 -65625
rect -10833 -66013 -10821 -65637
rect -10787 -66013 -10775 -65637
rect -10833 -66025 -10775 -66013
rect -10575 -65637 -10517 -65625
rect -10575 -66013 -10563 -65637
rect -10529 -66013 -10517 -65637
rect -10575 -66025 -10517 -66013
rect -10317 -65637 -10259 -65625
rect -10317 -66013 -10305 -65637
rect -10271 -66013 -10259 -65637
rect -10317 -66025 -10259 -66013
rect -10059 -65637 -10001 -65625
rect -10059 -66013 -10047 -65637
rect -10013 -66013 -10001 -65637
rect -10059 -66025 -10001 -66013
rect -9801 -65637 -9743 -65625
rect -9801 -66013 -9789 -65637
rect -9755 -66013 -9743 -65637
rect -9801 -66025 -9743 -66013
rect -11349 -66497 -11291 -66485
rect -11349 -66873 -11337 -66497
rect -11303 -66873 -11291 -66497
rect -11349 -66885 -11291 -66873
rect -11091 -66497 -11033 -66485
rect -11091 -66873 -11079 -66497
rect -11045 -66873 -11033 -66497
rect -11091 -66885 -11033 -66873
rect -10833 -66497 -10775 -66485
rect -10833 -66873 -10821 -66497
rect -10787 -66873 -10775 -66497
rect -10833 -66885 -10775 -66873
rect -10575 -66497 -10517 -66485
rect -10575 -66873 -10563 -66497
rect -10529 -66873 -10517 -66497
rect -10575 -66885 -10517 -66873
rect -10317 -66497 -10259 -66485
rect -10317 -66873 -10305 -66497
rect -10271 -66873 -10259 -66497
rect -10317 -66885 -10259 -66873
rect -10059 -66497 -10001 -66485
rect -10059 -66873 -10047 -66497
rect -10013 -66873 -10001 -66497
rect -10059 -66885 -10001 -66873
rect -9801 -66497 -9743 -66485
rect -9801 -66873 -9789 -66497
rect -9755 -66873 -9743 -66497
rect -9801 -66885 -9743 -66873
rect -8004 -67341 -7952 -67329
rect -8004 -67375 -7996 -67341
rect -7962 -67375 -7952 -67341
rect -8004 -67409 -7952 -67375
rect -8004 -67443 -7996 -67409
rect -7962 -67443 -7952 -67409
rect -8004 -67477 -7952 -67443
rect -8004 -67511 -7996 -67477
rect -7962 -67511 -7952 -67477
rect -8004 -67529 -7952 -67511
rect -7922 -67341 -7870 -67329
rect -7922 -67375 -7912 -67341
rect -7878 -67375 -7870 -67341
rect -7922 -67409 -7870 -67375
rect -7922 -67443 -7912 -67409
rect -7878 -67443 -7870 -67409
rect -7922 -67477 -7870 -67443
rect -7922 -67511 -7912 -67477
rect -7878 -67511 -7870 -67477
rect -7922 -67529 -7870 -67511
rect -7349 -65637 -7291 -65625
rect -7349 -66013 -7337 -65637
rect -7303 -66013 -7291 -65637
rect -7349 -66025 -7291 -66013
rect -7091 -65637 -7033 -65625
rect -7091 -66013 -7079 -65637
rect -7045 -66013 -7033 -65637
rect -7091 -66025 -7033 -66013
rect -6833 -65637 -6775 -65625
rect -6833 -66013 -6821 -65637
rect -6787 -66013 -6775 -65637
rect -6833 -66025 -6775 -66013
rect -6575 -65637 -6517 -65625
rect -6575 -66013 -6563 -65637
rect -6529 -66013 -6517 -65637
rect -6575 -66025 -6517 -66013
rect -6317 -65637 -6259 -65625
rect -6317 -66013 -6305 -65637
rect -6271 -66013 -6259 -65637
rect -6317 -66025 -6259 -66013
rect -6059 -65637 -6001 -65625
rect -6059 -66013 -6047 -65637
rect -6013 -66013 -6001 -65637
rect -6059 -66025 -6001 -66013
rect -5801 -65637 -5743 -65625
rect -5801 -66013 -5789 -65637
rect -5755 -66013 -5743 -65637
rect -5801 -66025 -5743 -66013
rect -7349 -66497 -7291 -66485
rect -7349 -66873 -7337 -66497
rect -7303 -66873 -7291 -66497
rect -7349 -66885 -7291 -66873
rect -7091 -66497 -7033 -66485
rect -7091 -66873 -7079 -66497
rect -7045 -66873 -7033 -66497
rect -7091 -66885 -7033 -66873
rect -6833 -66497 -6775 -66485
rect -6833 -66873 -6821 -66497
rect -6787 -66873 -6775 -66497
rect -6833 -66885 -6775 -66873
rect -6575 -66497 -6517 -66485
rect -6575 -66873 -6563 -66497
rect -6529 -66873 -6517 -66497
rect -6575 -66885 -6517 -66873
rect -6317 -66497 -6259 -66485
rect -6317 -66873 -6305 -66497
rect -6271 -66873 -6259 -66497
rect -6317 -66885 -6259 -66873
rect -6059 -66497 -6001 -66485
rect -6059 -66873 -6047 -66497
rect -6013 -66873 -6001 -66497
rect -6059 -66885 -6001 -66873
rect -5801 -66497 -5743 -66485
rect -5801 -66873 -5789 -66497
rect -5755 -66873 -5743 -66497
rect -5801 -66885 -5743 -66873
rect -4004 -67341 -3952 -67329
rect -4004 -67375 -3996 -67341
rect -3962 -67375 -3952 -67341
rect -4004 -67409 -3952 -67375
rect -4004 -67443 -3996 -67409
rect -3962 -67443 -3952 -67409
rect -4004 -67477 -3952 -67443
rect -4004 -67511 -3996 -67477
rect -3962 -67511 -3952 -67477
rect -4004 -67529 -3952 -67511
rect -3922 -67341 -3870 -67329
rect -3922 -67375 -3912 -67341
rect -3878 -67375 -3870 -67341
rect -3922 -67409 -3870 -67375
rect -3922 -67443 -3912 -67409
rect -3878 -67443 -3870 -67409
rect -3922 -67477 -3870 -67443
rect -3922 -67511 -3912 -67477
rect -3878 -67511 -3870 -67477
rect -3922 -67529 -3870 -67511
rect -3349 -65637 -3291 -65625
rect -3349 -66013 -3337 -65637
rect -3303 -66013 -3291 -65637
rect -3349 -66025 -3291 -66013
rect -3091 -65637 -3033 -65625
rect -3091 -66013 -3079 -65637
rect -3045 -66013 -3033 -65637
rect -3091 -66025 -3033 -66013
rect -2833 -65637 -2775 -65625
rect -2833 -66013 -2821 -65637
rect -2787 -66013 -2775 -65637
rect -2833 -66025 -2775 -66013
rect -2575 -65637 -2517 -65625
rect -2575 -66013 -2563 -65637
rect -2529 -66013 -2517 -65637
rect -2575 -66025 -2517 -66013
rect -2317 -65637 -2259 -65625
rect -2317 -66013 -2305 -65637
rect -2271 -66013 -2259 -65637
rect -2317 -66025 -2259 -66013
rect -2059 -65637 -2001 -65625
rect -2059 -66013 -2047 -65637
rect -2013 -66013 -2001 -65637
rect -2059 -66025 -2001 -66013
rect -1801 -65637 -1743 -65625
rect -1801 -66013 -1789 -65637
rect -1755 -66013 -1743 -65637
rect -1801 -66025 -1743 -66013
rect -3349 -66497 -3291 -66485
rect -3349 -66873 -3337 -66497
rect -3303 -66873 -3291 -66497
rect -3349 -66885 -3291 -66873
rect -3091 -66497 -3033 -66485
rect -3091 -66873 -3079 -66497
rect -3045 -66873 -3033 -66497
rect -3091 -66885 -3033 -66873
rect -2833 -66497 -2775 -66485
rect -2833 -66873 -2821 -66497
rect -2787 -66873 -2775 -66497
rect -2833 -66885 -2775 -66873
rect -2575 -66497 -2517 -66485
rect -2575 -66873 -2563 -66497
rect -2529 -66873 -2517 -66497
rect -2575 -66885 -2517 -66873
rect -2317 -66497 -2259 -66485
rect -2317 -66873 -2305 -66497
rect -2271 -66873 -2259 -66497
rect -2317 -66885 -2259 -66873
rect -2059 -66497 -2001 -66485
rect -2059 -66873 -2047 -66497
rect -2013 -66873 -2001 -66497
rect -2059 -66885 -2001 -66873
rect -1801 -66497 -1743 -66485
rect -1801 -66873 -1789 -66497
rect -1755 -66873 -1743 -66497
rect -1801 -66885 -1743 -66873
rect -4 -67341 48 -67329
rect -4 -67375 4 -67341
rect 38 -67375 48 -67341
rect -4 -67409 48 -67375
rect -4 -67443 4 -67409
rect 38 -67443 48 -67409
rect -4 -67477 48 -67443
rect -4 -67511 4 -67477
rect 38 -67511 48 -67477
rect -4 -67529 48 -67511
rect 78 -67341 130 -67329
rect 78 -67375 88 -67341
rect 122 -67375 130 -67341
rect 78 -67409 130 -67375
rect 78 -67443 88 -67409
rect 122 -67443 130 -67409
rect 78 -67477 130 -67443
rect 78 -67511 88 -67477
rect 122 -67511 130 -67477
rect 78 -67529 130 -67511
rect 651 -65637 709 -65625
rect 651 -66013 663 -65637
rect 697 -66013 709 -65637
rect 651 -66025 709 -66013
rect 909 -65637 967 -65625
rect 909 -66013 921 -65637
rect 955 -66013 967 -65637
rect 909 -66025 967 -66013
rect 1167 -65637 1225 -65625
rect 1167 -66013 1179 -65637
rect 1213 -66013 1225 -65637
rect 1167 -66025 1225 -66013
rect 1425 -65637 1483 -65625
rect 1425 -66013 1437 -65637
rect 1471 -66013 1483 -65637
rect 1425 -66025 1483 -66013
rect 1683 -65637 1741 -65625
rect 1683 -66013 1695 -65637
rect 1729 -66013 1741 -65637
rect 1683 -66025 1741 -66013
rect 1941 -65637 1999 -65625
rect 1941 -66013 1953 -65637
rect 1987 -66013 1999 -65637
rect 1941 -66025 1999 -66013
rect 2199 -65637 2257 -65625
rect 2199 -66013 2211 -65637
rect 2245 -66013 2257 -65637
rect 2199 -66025 2257 -66013
rect 651 -66497 709 -66485
rect 651 -66873 663 -66497
rect 697 -66873 709 -66497
rect 651 -66885 709 -66873
rect 909 -66497 967 -66485
rect 909 -66873 921 -66497
rect 955 -66873 967 -66497
rect 909 -66885 967 -66873
rect 1167 -66497 1225 -66485
rect 1167 -66873 1179 -66497
rect 1213 -66873 1225 -66497
rect 1167 -66885 1225 -66873
rect 1425 -66497 1483 -66485
rect 1425 -66873 1437 -66497
rect 1471 -66873 1483 -66497
rect 1425 -66885 1483 -66873
rect 1683 -66497 1741 -66485
rect 1683 -66873 1695 -66497
rect 1729 -66873 1741 -66497
rect 1683 -66885 1741 -66873
rect 1941 -66497 1999 -66485
rect 1941 -66873 1953 -66497
rect 1987 -66873 1999 -66497
rect 1941 -66885 1999 -66873
rect 2199 -66497 2257 -66485
rect 2199 -66873 2211 -66497
rect 2245 -66873 2257 -66497
rect 2199 -66885 2257 -66873
rect 3996 -67341 4048 -67329
rect 3996 -67375 4004 -67341
rect 4038 -67375 4048 -67341
rect 3996 -67409 4048 -67375
rect 3996 -67443 4004 -67409
rect 4038 -67443 4048 -67409
rect 3996 -67477 4048 -67443
rect 3996 -67511 4004 -67477
rect 4038 -67511 4048 -67477
rect 3996 -67529 4048 -67511
rect 4078 -67341 4130 -67329
rect 4078 -67375 4088 -67341
rect 4122 -67375 4130 -67341
rect 4078 -67409 4130 -67375
rect 4078 -67443 4088 -67409
rect 4122 -67443 4130 -67409
rect 4078 -67477 4130 -67443
rect 4078 -67511 4088 -67477
rect 4122 -67511 4130 -67477
rect 4078 -67529 4130 -67511
rect 4651 -65637 4709 -65625
rect 4651 -66013 4663 -65637
rect 4697 -66013 4709 -65637
rect 4651 -66025 4709 -66013
rect 4909 -65637 4967 -65625
rect 4909 -66013 4921 -65637
rect 4955 -66013 4967 -65637
rect 4909 -66025 4967 -66013
rect 5167 -65637 5225 -65625
rect 5167 -66013 5179 -65637
rect 5213 -66013 5225 -65637
rect 5167 -66025 5225 -66013
rect 5425 -65637 5483 -65625
rect 5425 -66013 5437 -65637
rect 5471 -66013 5483 -65637
rect 5425 -66025 5483 -66013
rect 5683 -65637 5741 -65625
rect 5683 -66013 5695 -65637
rect 5729 -66013 5741 -65637
rect 5683 -66025 5741 -66013
rect 5941 -65637 5999 -65625
rect 5941 -66013 5953 -65637
rect 5987 -66013 5999 -65637
rect 5941 -66025 5999 -66013
rect 6199 -65637 6257 -65625
rect 6199 -66013 6211 -65637
rect 6245 -66013 6257 -65637
rect 6199 -66025 6257 -66013
rect 4651 -66497 4709 -66485
rect 4651 -66873 4663 -66497
rect 4697 -66873 4709 -66497
rect 4651 -66885 4709 -66873
rect 4909 -66497 4967 -66485
rect 4909 -66873 4921 -66497
rect 4955 -66873 4967 -66497
rect 4909 -66885 4967 -66873
rect 5167 -66497 5225 -66485
rect 5167 -66873 5179 -66497
rect 5213 -66873 5225 -66497
rect 5167 -66885 5225 -66873
rect 5425 -66497 5483 -66485
rect 5425 -66873 5437 -66497
rect 5471 -66873 5483 -66497
rect 5425 -66885 5483 -66873
rect 5683 -66497 5741 -66485
rect 5683 -66873 5695 -66497
rect 5729 -66873 5741 -66497
rect 5683 -66885 5741 -66873
rect 5941 -66497 5999 -66485
rect 5941 -66873 5953 -66497
rect 5987 -66873 5999 -66497
rect 5941 -66885 5999 -66873
rect 6199 -66497 6257 -66485
rect 6199 -66873 6211 -66497
rect 6245 -66873 6257 -66497
rect 6199 -66885 6257 -66873
rect -28004 -72685 -27952 -72667
rect -28004 -72719 -27996 -72685
rect -27962 -72719 -27952 -72685
rect -28004 -72753 -27952 -72719
rect -28004 -72787 -27996 -72753
rect -27962 -72787 -27952 -72753
rect -28004 -72821 -27952 -72787
rect -28004 -72855 -27996 -72821
rect -27962 -72855 -27952 -72821
rect -28004 -72867 -27952 -72855
rect -27922 -72685 -27870 -72667
rect -27922 -72719 -27912 -72685
rect -27878 -72719 -27870 -72685
rect -27922 -72753 -27870 -72719
rect -27922 -72787 -27912 -72753
rect -27878 -72787 -27870 -72753
rect -27922 -72821 -27870 -72787
rect -27922 -72855 -27912 -72821
rect -27878 -72855 -27870 -72821
rect -27922 -72867 -27870 -72855
rect -27349 -73323 -27291 -73311
rect -27349 -73699 -27337 -73323
rect -27303 -73699 -27291 -73323
rect -27349 -73711 -27291 -73699
rect -27091 -73323 -27033 -73311
rect -27091 -73699 -27079 -73323
rect -27045 -73699 -27033 -73323
rect -27091 -73711 -27033 -73699
rect -26833 -73323 -26775 -73311
rect -26833 -73699 -26821 -73323
rect -26787 -73699 -26775 -73323
rect -26833 -73711 -26775 -73699
rect -26575 -73323 -26517 -73311
rect -26575 -73699 -26563 -73323
rect -26529 -73699 -26517 -73323
rect -26575 -73711 -26517 -73699
rect -26317 -73323 -26259 -73311
rect -26317 -73699 -26305 -73323
rect -26271 -73699 -26259 -73323
rect -26317 -73711 -26259 -73699
rect -26059 -73323 -26001 -73311
rect -26059 -73699 -26047 -73323
rect -26013 -73699 -26001 -73323
rect -26059 -73711 -26001 -73699
rect -25801 -73323 -25743 -73311
rect -25801 -73699 -25789 -73323
rect -25755 -73699 -25743 -73323
rect -25801 -73711 -25743 -73699
rect -27349 -74183 -27291 -74171
rect -27349 -74559 -27337 -74183
rect -27303 -74559 -27291 -74183
rect -27349 -74571 -27291 -74559
rect -27091 -74183 -27033 -74171
rect -27091 -74559 -27079 -74183
rect -27045 -74559 -27033 -74183
rect -27091 -74571 -27033 -74559
rect -26833 -74183 -26775 -74171
rect -26833 -74559 -26821 -74183
rect -26787 -74559 -26775 -74183
rect -26833 -74571 -26775 -74559
rect -26575 -74183 -26517 -74171
rect -26575 -74559 -26563 -74183
rect -26529 -74559 -26517 -74183
rect -26575 -74571 -26517 -74559
rect -26317 -74183 -26259 -74171
rect -26317 -74559 -26305 -74183
rect -26271 -74559 -26259 -74183
rect -26317 -74571 -26259 -74559
rect -26059 -74183 -26001 -74171
rect -26059 -74559 -26047 -74183
rect -26013 -74559 -26001 -74183
rect -26059 -74571 -26001 -74559
rect -25801 -74183 -25743 -74171
rect -25801 -74559 -25789 -74183
rect -25755 -74559 -25743 -74183
rect -25801 -74571 -25743 -74559
rect -24004 -72685 -23952 -72667
rect -24004 -72719 -23996 -72685
rect -23962 -72719 -23952 -72685
rect -24004 -72753 -23952 -72719
rect -24004 -72787 -23996 -72753
rect -23962 -72787 -23952 -72753
rect -24004 -72821 -23952 -72787
rect -24004 -72855 -23996 -72821
rect -23962 -72855 -23952 -72821
rect -24004 -72867 -23952 -72855
rect -23922 -72685 -23870 -72667
rect -23922 -72719 -23912 -72685
rect -23878 -72719 -23870 -72685
rect -23922 -72753 -23870 -72719
rect -23922 -72787 -23912 -72753
rect -23878 -72787 -23870 -72753
rect -23922 -72821 -23870 -72787
rect -23922 -72855 -23912 -72821
rect -23878 -72855 -23870 -72821
rect -23922 -72867 -23870 -72855
rect -23349 -73323 -23291 -73311
rect -23349 -73699 -23337 -73323
rect -23303 -73699 -23291 -73323
rect -23349 -73711 -23291 -73699
rect -23091 -73323 -23033 -73311
rect -23091 -73699 -23079 -73323
rect -23045 -73699 -23033 -73323
rect -23091 -73711 -23033 -73699
rect -22833 -73323 -22775 -73311
rect -22833 -73699 -22821 -73323
rect -22787 -73699 -22775 -73323
rect -22833 -73711 -22775 -73699
rect -22575 -73323 -22517 -73311
rect -22575 -73699 -22563 -73323
rect -22529 -73699 -22517 -73323
rect -22575 -73711 -22517 -73699
rect -22317 -73323 -22259 -73311
rect -22317 -73699 -22305 -73323
rect -22271 -73699 -22259 -73323
rect -22317 -73711 -22259 -73699
rect -22059 -73323 -22001 -73311
rect -22059 -73699 -22047 -73323
rect -22013 -73699 -22001 -73323
rect -22059 -73711 -22001 -73699
rect -21801 -73323 -21743 -73311
rect -21801 -73699 -21789 -73323
rect -21755 -73699 -21743 -73323
rect -21801 -73711 -21743 -73699
rect -23349 -74183 -23291 -74171
rect -23349 -74559 -23337 -74183
rect -23303 -74559 -23291 -74183
rect -23349 -74571 -23291 -74559
rect -23091 -74183 -23033 -74171
rect -23091 -74559 -23079 -74183
rect -23045 -74559 -23033 -74183
rect -23091 -74571 -23033 -74559
rect -22833 -74183 -22775 -74171
rect -22833 -74559 -22821 -74183
rect -22787 -74559 -22775 -74183
rect -22833 -74571 -22775 -74559
rect -22575 -74183 -22517 -74171
rect -22575 -74559 -22563 -74183
rect -22529 -74559 -22517 -74183
rect -22575 -74571 -22517 -74559
rect -22317 -74183 -22259 -74171
rect -22317 -74559 -22305 -74183
rect -22271 -74559 -22259 -74183
rect -22317 -74571 -22259 -74559
rect -22059 -74183 -22001 -74171
rect -22059 -74559 -22047 -74183
rect -22013 -74559 -22001 -74183
rect -22059 -74571 -22001 -74559
rect -21801 -74183 -21743 -74171
rect -21801 -74559 -21789 -74183
rect -21755 -74559 -21743 -74183
rect -21801 -74571 -21743 -74559
rect -20004 -72685 -19952 -72667
rect -20004 -72719 -19996 -72685
rect -19962 -72719 -19952 -72685
rect -20004 -72753 -19952 -72719
rect -20004 -72787 -19996 -72753
rect -19962 -72787 -19952 -72753
rect -20004 -72821 -19952 -72787
rect -20004 -72855 -19996 -72821
rect -19962 -72855 -19952 -72821
rect -20004 -72867 -19952 -72855
rect -19922 -72685 -19870 -72667
rect -19922 -72719 -19912 -72685
rect -19878 -72719 -19870 -72685
rect -19922 -72753 -19870 -72719
rect -19922 -72787 -19912 -72753
rect -19878 -72787 -19870 -72753
rect -19922 -72821 -19870 -72787
rect -19922 -72855 -19912 -72821
rect -19878 -72855 -19870 -72821
rect -19922 -72867 -19870 -72855
rect -19349 -73323 -19291 -73311
rect -19349 -73699 -19337 -73323
rect -19303 -73699 -19291 -73323
rect -19349 -73711 -19291 -73699
rect -19091 -73323 -19033 -73311
rect -19091 -73699 -19079 -73323
rect -19045 -73699 -19033 -73323
rect -19091 -73711 -19033 -73699
rect -18833 -73323 -18775 -73311
rect -18833 -73699 -18821 -73323
rect -18787 -73699 -18775 -73323
rect -18833 -73711 -18775 -73699
rect -18575 -73323 -18517 -73311
rect -18575 -73699 -18563 -73323
rect -18529 -73699 -18517 -73323
rect -18575 -73711 -18517 -73699
rect -18317 -73323 -18259 -73311
rect -18317 -73699 -18305 -73323
rect -18271 -73699 -18259 -73323
rect -18317 -73711 -18259 -73699
rect -18059 -73323 -18001 -73311
rect -18059 -73699 -18047 -73323
rect -18013 -73699 -18001 -73323
rect -18059 -73711 -18001 -73699
rect -17801 -73323 -17743 -73311
rect -17801 -73699 -17789 -73323
rect -17755 -73699 -17743 -73323
rect -17801 -73711 -17743 -73699
rect -19349 -74183 -19291 -74171
rect -19349 -74559 -19337 -74183
rect -19303 -74559 -19291 -74183
rect -19349 -74571 -19291 -74559
rect -19091 -74183 -19033 -74171
rect -19091 -74559 -19079 -74183
rect -19045 -74559 -19033 -74183
rect -19091 -74571 -19033 -74559
rect -18833 -74183 -18775 -74171
rect -18833 -74559 -18821 -74183
rect -18787 -74559 -18775 -74183
rect -18833 -74571 -18775 -74559
rect -18575 -74183 -18517 -74171
rect -18575 -74559 -18563 -74183
rect -18529 -74559 -18517 -74183
rect -18575 -74571 -18517 -74559
rect -18317 -74183 -18259 -74171
rect -18317 -74559 -18305 -74183
rect -18271 -74559 -18259 -74183
rect -18317 -74571 -18259 -74559
rect -18059 -74183 -18001 -74171
rect -18059 -74559 -18047 -74183
rect -18013 -74559 -18001 -74183
rect -18059 -74571 -18001 -74559
rect -17801 -74183 -17743 -74171
rect -17801 -74559 -17789 -74183
rect -17755 -74559 -17743 -74183
rect -17801 -74571 -17743 -74559
rect -16004 -72685 -15952 -72667
rect -16004 -72719 -15996 -72685
rect -15962 -72719 -15952 -72685
rect -16004 -72753 -15952 -72719
rect -16004 -72787 -15996 -72753
rect -15962 -72787 -15952 -72753
rect -16004 -72821 -15952 -72787
rect -16004 -72855 -15996 -72821
rect -15962 -72855 -15952 -72821
rect -16004 -72867 -15952 -72855
rect -15922 -72685 -15870 -72667
rect -15922 -72719 -15912 -72685
rect -15878 -72719 -15870 -72685
rect -15922 -72753 -15870 -72719
rect -15922 -72787 -15912 -72753
rect -15878 -72787 -15870 -72753
rect -15922 -72821 -15870 -72787
rect -15922 -72855 -15912 -72821
rect -15878 -72855 -15870 -72821
rect -15922 -72867 -15870 -72855
rect -15349 -73323 -15291 -73311
rect -15349 -73699 -15337 -73323
rect -15303 -73699 -15291 -73323
rect -15349 -73711 -15291 -73699
rect -15091 -73323 -15033 -73311
rect -15091 -73699 -15079 -73323
rect -15045 -73699 -15033 -73323
rect -15091 -73711 -15033 -73699
rect -14833 -73323 -14775 -73311
rect -14833 -73699 -14821 -73323
rect -14787 -73699 -14775 -73323
rect -14833 -73711 -14775 -73699
rect -14575 -73323 -14517 -73311
rect -14575 -73699 -14563 -73323
rect -14529 -73699 -14517 -73323
rect -14575 -73711 -14517 -73699
rect -14317 -73323 -14259 -73311
rect -14317 -73699 -14305 -73323
rect -14271 -73699 -14259 -73323
rect -14317 -73711 -14259 -73699
rect -14059 -73323 -14001 -73311
rect -14059 -73699 -14047 -73323
rect -14013 -73699 -14001 -73323
rect -14059 -73711 -14001 -73699
rect -13801 -73323 -13743 -73311
rect -13801 -73699 -13789 -73323
rect -13755 -73699 -13743 -73323
rect -13801 -73711 -13743 -73699
rect -15349 -74183 -15291 -74171
rect -15349 -74559 -15337 -74183
rect -15303 -74559 -15291 -74183
rect -15349 -74571 -15291 -74559
rect -15091 -74183 -15033 -74171
rect -15091 -74559 -15079 -74183
rect -15045 -74559 -15033 -74183
rect -15091 -74571 -15033 -74559
rect -14833 -74183 -14775 -74171
rect -14833 -74559 -14821 -74183
rect -14787 -74559 -14775 -74183
rect -14833 -74571 -14775 -74559
rect -14575 -74183 -14517 -74171
rect -14575 -74559 -14563 -74183
rect -14529 -74559 -14517 -74183
rect -14575 -74571 -14517 -74559
rect -14317 -74183 -14259 -74171
rect -14317 -74559 -14305 -74183
rect -14271 -74559 -14259 -74183
rect -14317 -74571 -14259 -74559
rect -14059 -74183 -14001 -74171
rect -14059 -74559 -14047 -74183
rect -14013 -74559 -14001 -74183
rect -14059 -74571 -14001 -74559
rect -13801 -74183 -13743 -74171
rect -13801 -74559 -13789 -74183
rect -13755 -74559 -13743 -74183
rect -13801 -74571 -13743 -74559
rect -12004 -72685 -11952 -72667
rect -12004 -72719 -11996 -72685
rect -11962 -72719 -11952 -72685
rect -12004 -72753 -11952 -72719
rect -12004 -72787 -11996 -72753
rect -11962 -72787 -11952 -72753
rect -12004 -72821 -11952 -72787
rect -12004 -72855 -11996 -72821
rect -11962 -72855 -11952 -72821
rect -12004 -72867 -11952 -72855
rect -11922 -72685 -11870 -72667
rect -11922 -72719 -11912 -72685
rect -11878 -72719 -11870 -72685
rect -11922 -72753 -11870 -72719
rect -11922 -72787 -11912 -72753
rect -11878 -72787 -11870 -72753
rect -11922 -72821 -11870 -72787
rect -11922 -72855 -11912 -72821
rect -11878 -72855 -11870 -72821
rect -11922 -72867 -11870 -72855
rect -11349 -73323 -11291 -73311
rect -11349 -73699 -11337 -73323
rect -11303 -73699 -11291 -73323
rect -11349 -73711 -11291 -73699
rect -11091 -73323 -11033 -73311
rect -11091 -73699 -11079 -73323
rect -11045 -73699 -11033 -73323
rect -11091 -73711 -11033 -73699
rect -10833 -73323 -10775 -73311
rect -10833 -73699 -10821 -73323
rect -10787 -73699 -10775 -73323
rect -10833 -73711 -10775 -73699
rect -10575 -73323 -10517 -73311
rect -10575 -73699 -10563 -73323
rect -10529 -73699 -10517 -73323
rect -10575 -73711 -10517 -73699
rect -10317 -73323 -10259 -73311
rect -10317 -73699 -10305 -73323
rect -10271 -73699 -10259 -73323
rect -10317 -73711 -10259 -73699
rect -10059 -73323 -10001 -73311
rect -10059 -73699 -10047 -73323
rect -10013 -73699 -10001 -73323
rect -10059 -73711 -10001 -73699
rect -9801 -73323 -9743 -73311
rect -9801 -73699 -9789 -73323
rect -9755 -73699 -9743 -73323
rect -9801 -73711 -9743 -73699
rect -11349 -74183 -11291 -74171
rect -11349 -74559 -11337 -74183
rect -11303 -74559 -11291 -74183
rect -11349 -74571 -11291 -74559
rect -11091 -74183 -11033 -74171
rect -11091 -74559 -11079 -74183
rect -11045 -74559 -11033 -74183
rect -11091 -74571 -11033 -74559
rect -10833 -74183 -10775 -74171
rect -10833 -74559 -10821 -74183
rect -10787 -74559 -10775 -74183
rect -10833 -74571 -10775 -74559
rect -10575 -74183 -10517 -74171
rect -10575 -74559 -10563 -74183
rect -10529 -74559 -10517 -74183
rect -10575 -74571 -10517 -74559
rect -10317 -74183 -10259 -74171
rect -10317 -74559 -10305 -74183
rect -10271 -74559 -10259 -74183
rect -10317 -74571 -10259 -74559
rect -10059 -74183 -10001 -74171
rect -10059 -74559 -10047 -74183
rect -10013 -74559 -10001 -74183
rect -10059 -74571 -10001 -74559
rect -9801 -74183 -9743 -74171
rect -9801 -74559 -9789 -74183
rect -9755 -74559 -9743 -74183
rect -9801 -74571 -9743 -74559
rect -8004 -72685 -7952 -72667
rect -8004 -72719 -7996 -72685
rect -7962 -72719 -7952 -72685
rect -8004 -72753 -7952 -72719
rect -8004 -72787 -7996 -72753
rect -7962 -72787 -7952 -72753
rect -8004 -72821 -7952 -72787
rect -8004 -72855 -7996 -72821
rect -7962 -72855 -7952 -72821
rect -8004 -72867 -7952 -72855
rect -7922 -72685 -7870 -72667
rect -7922 -72719 -7912 -72685
rect -7878 -72719 -7870 -72685
rect -7922 -72753 -7870 -72719
rect -7922 -72787 -7912 -72753
rect -7878 -72787 -7870 -72753
rect -7922 -72821 -7870 -72787
rect -7922 -72855 -7912 -72821
rect -7878 -72855 -7870 -72821
rect -7922 -72867 -7870 -72855
rect -7349 -73323 -7291 -73311
rect -7349 -73699 -7337 -73323
rect -7303 -73699 -7291 -73323
rect -7349 -73711 -7291 -73699
rect -7091 -73323 -7033 -73311
rect -7091 -73699 -7079 -73323
rect -7045 -73699 -7033 -73323
rect -7091 -73711 -7033 -73699
rect -6833 -73323 -6775 -73311
rect -6833 -73699 -6821 -73323
rect -6787 -73699 -6775 -73323
rect -6833 -73711 -6775 -73699
rect -6575 -73323 -6517 -73311
rect -6575 -73699 -6563 -73323
rect -6529 -73699 -6517 -73323
rect -6575 -73711 -6517 -73699
rect -6317 -73323 -6259 -73311
rect -6317 -73699 -6305 -73323
rect -6271 -73699 -6259 -73323
rect -6317 -73711 -6259 -73699
rect -6059 -73323 -6001 -73311
rect -6059 -73699 -6047 -73323
rect -6013 -73699 -6001 -73323
rect -6059 -73711 -6001 -73699
rect -5801 -73323 -5743 -73311
rect -5801 -73699 -5789 -73323
rect -5755 -73699 -5743 -73323
rect -5801 -73711 -5743 -73699
rect -7349 -74183 -7291 -74171
rect -7349 -74559 -7337 -74183
rect -7303 -74559 -7291 -74183
rect -7349 -74571 -7291 -74559
rect -7091 -74183 -7033 -74171
rect -7091 -74559 -7079 -74183
rect -7045 -74559 -7033 -74183
rect -7091 -74571 -7033 -74559
rect -6833 -74183 -6775 -74171
rect -6833 -74559 -6821 -74183
rect -6787 -74559 -6775 -74183
rect -6833 -74571 -6775 -74559
rect -6575 -74183 -6517 -74171
rect -6575 -74559 -6563 -74183
rect -6529 -74559 -6517 -74183
rect -6575 -74571 -6517 -74559
rect -6317 -74183 -6259 -74171
rect -6317 -74559 -6305 -74183
rect -6271 -74559 -6259 -74183
rect -6317 -74571 -6259 -74559
rect -6059 -74183 -6001 -74171
rect -6059 -74559 -6047 -74183
rect -6013 -74559 -6001 -74183
rect -6059 -74571 -6001 -74559
rect -5801 -74183 -5743 -74171
rect -5801 -74559 -5789 -74183
rect -5755 -74559 -5743 -74183
rect -5801 -74571 -5743 -74559
rect -4004 -72685 -3952 -72667
rect -4004 -72719 -3996 -72685
rect -3962 -72719 -3952 -72685
rect -4004 -72753 -3952 -72719
rect -4004 -72787 -3996 -72753
rect -3962 -72787 -3952 -72753
rect -4004 -72821 -3952 -72787
rect -4004 -72855 -3996 -72821
rect -3962 -72855 -3952 -72821
rect -4004 -72867 -3952 -72855
rect -3922 -72685 -3870 -72667
rect -3922 -72719 -3912 -72685
rect -3878 -72719 -3870 -72685
rect -3922 -72753 -3870 -72719
rect -3922 -72787 -3912 -72753
rect -3878 -72787 -3870 -72753
rect -3922 -72821 -3870 -72787
rect -3922 -72855 -3912 -72821
rect -3878 -72855 -3870 -72821
rect -3922 -72867 -3870 -72855
rect -3349 -73323 -3291 -73311
rect -3349 -73699 -3337 -73323
rect -3303 -73699 -3291 -73323
rect -3349 -73711 -3291 -73699
rect -3091 -73323 -3033 -73311
rect -3091 -73699 -3079 -73323
rect -3045 -73699 -3033 -73323
rect -3091 -73711 -3033 -73699
rect -2833 -73323 -2775 -73311
rect -2833 -73699 -2821 -73323
rect -2787 -73699 -2775 -73323
rect -2833 -73711 -2775 -73699
rect -2575 -73323 -2517 -73311
rect -2575 -73699 -2563 -73323
rect -2529 -73699 -2517 -73323
rect -2575 -73711 -2517 -73699
rect -2317 -73323 -2259 -73311
rect -2317 -73699 -2305 -73323
rect -2271 -73699 -2259 -73323
rect -2317 -73711 -2259 -73699
rect -2059 -73323 -2001 -73311
rect -2059 -73699 -2047 -73323
rect -2013 -73699 -2001 -73323
rect -2059 -73711 -2001 -73699
rect -1801 -73323 -1743 -73311
rect -1801 -73699 -1789 -73323
rect -1755 -73699 -1743 -73323
rect -1801 -73711 -1743 -73699
rect -3349 -74183 -3291 -74171
rect -3349 -74559 -3337 -74183
rect -3303 -74559 -3291 -74183
rect -3349 -74571 -3291 -74559
rect -3091 -74183 -3033 -74171
rect -3091 -74559 -3079 -74183
rect -3045 -74559 -3033 -74183
rect -3091 -74571 -3033 -74559
rect -2833 -74183 -2775 -74171
rect -2833 -74559 -2821 -74183
rect -2787 -74559 -2775 -74183
rect -2833 -74571 -2775 -74559
rect -2575 -74183 -2517 -74171
rect -2575 -74559 -2563 -74183
rect -2529 -74559 -2517 -74183
rect -2575 -74571 -2517 -74559
rect -2317 -74183 -2259 -74171
rect -2317 -74559 -2305 -74183
rect -2271 -74559 -2259 -74183
rect -2317 -74571 -2259 -74559
rect -2059 -74183 -2001 -74171
rect -2059 -74559 -2047 -74183
rect -2013 -74559 -2001 -74183
rect -2059 -74571 -2001 -74559
rect -1801 -74183 -1743 -74171
rect -1801 -74559 -1789 -74183
rect -1755 -74559 -1743 -74183
rect -1801 -74571 -1743 -74559
rect -4 -72685 48 -72667
rect -4 -72719 4 -72685
rect 38 -72719 48 -72685
rect -4 -72753 48 -72719
rect -4 -72787 4 -72753
rect 38 -72787 48 -72753
rect -4 -72821 48 -72787
rect -4 -72855 4 -72821
rect 38 -72855 48 -72821
rect -4 -72867 48 -72855
rect 78 -72685 130 -72667
rect 78 -72719 88 -72685
rect 122 -72719 130 -72685
rect 78 -72753 130 -72719
rect 78 -72787 88 -72753
rect 122 -72787 130 -72753
rect 78 -72821 130 -72787
rect 78 -72855 88 -72821
rect 122 -72855 130 -72821
rect 78 -72867 130 -72855
rect 651 -73323 709 -73311
rect 651 -73699 663 -73323
rect 697 -73699 709 -73323
rect 651 -73711 709 -73699
rect 909 -73323 967 -73311
rect 909 -73699 921 -73323
rect 955 -73699 967 -73323
rect 909 -73711 967 -73699
rect 1167 -73323 1225 -73311
rect 1167 -73699 1179 -73323
rect 1213 -73699 1225 -73323
rect 1167 -73711 1225 -73699
rect 1425 -73323 1483 -73311
rect 1425 -73699 1437 -73323
rect 1471 -73699 1483 -73323
rect 1425 -73711 1483 -73699
rect 1683 -73323 1741 -73311
rect 1683 -73699 1695 -73323
rect 1729 -73699 1741 -73323
rect 1683 -73711 1741 -73699
rect 1941 -73323 1999 -73311
rect 1941 -73699 1953 -73323
rect 1987 -73699 1999 -73323
rect 1941 -73711 1999 -73699
rect 2199 -73323 2257 -73311
rect 2199 -73699 2211 -73323
rect 2245 -73699 2257 -73323
rect 2199 -73711 2257 -73699
rect 651 -74183 709 -74171
rect 651 -74559 663 -74183
rect 697 -74559 709 -74183
rect 651 -74571 709 -74559
rect 909 -74183 967 -74171
rect 909 -74559 921 -74183
rect 955 -74559 967 -74183
rect 909 -74571 967 -74559
rect 1167 -74183 1225 -74171
rect 1167 -74559 1179 -74183
rect 1213 -74559 1225 -74183
rect 1167 -74571 1225 -74559
rect 1425 -74183 1483 -74171
rect 1425 -74559 1437 -74183
rect 1471 -74559 1483 -74183
rect 1425 -74571 1483 -74559
rect 1683 -74183 1741 -74171
rect 1683 -74559 1695 -74183
rect 1729 -74559 1741 -74183
rect 1683 -74571 1741 -74559
rect 1941 -74183 1999 -74171
rect 1941 -74559 1953 -74183
rect 1987 -74559 1999 -74183
rect 1941 -74571 1999 -74559
rect 2199 -74183 2257 -74171
rect 2199 -74559 2211 -74183
rect 2245 -74559 2257 -74183
rect 2199 -74571 2257 -74559
rect 3996 -72685 4048 -72667
rect 3996 -72719 4004 -72685
rect 4038 -72719 4048 -72685
rect 3996 -72753 4048 -72719
rect 3996 -72787 4004 -72753
rect 4038 -72787 4048 -72753
rect 3996 -72821 4048 -72787
rect 3996 -72855 4004 -72821
rect 4038 -72855 4048 -72821
rect 3996 -72867 4048 -72855
rect 4078 -72685 4130 -72667
rect 4078 -72719 4088 -72685
rect 4122 -72719 4130 -72685
rect 4078 -72753 4130 -72719
rect 4078 -72787 4088 -72753
rect 4122 -72787 4130 -72753
rect 4078 -72821 4130 -72787
rect 4078 -72855 4088 -72821
rect 4122 -72855 4130 -72821
rect 4078 -72867 4130 -72855
rect 4651 -73323 4709 -73311
rect 4651 -73699 4663 -73323
rect 4697 -73699 4709 -73323
rect 4651 -73711 4709 -73699
rect 4909 -73323 4967 -73311
rect 4909 -73699 4921 -73323
rect 4955 -73699 4967 -73323
rect 4909 -73711 4967 -73699
rect 5167 -73323 5225 -73311
rect 5167 -73699 5179 -73323
rect 5213 -73699 5225 -73323
rect 5167 -73711 5225 -73699
rect 5425 -73323 5483 -73311
rect 5425 -73699 5437 -73323
rect 5471 -73699 5483 -73323
rect 5425 -73711 5483 -73699
rect 5683 -73323 5741 -73311
rect 5683 -73699 5695 -73323
rect 5729 -73699 5741 -73323
rect 5683 -73711 5741 -73699
rect 5941 -73323 5999 -73311
rect 5941 -73699 5953 -73323
rect 5987 -73699 5999 -73323
rect 5941 -73711 5999 -73699
rect 6199 -73323 6257 -73311
rect 6199 -73699 6211 -73323
rect 6245 -73699 6257 -73323
rect 6199 -73711 6257 -73699
rect 4651 -74183 4709 -74171
rect 4651 -74559 4663 -74183
rect 4697 -74559 4709 -74183
rect 4651 -74571 4709 -74559
rect 4909 -74183 4967 -74171
rect 4909 -74559 4921 -74183
rect 4955 -74559 4967 -74183
rect 4909 -74571 4967 -74559
rect 5167 -74183 5225 -74171
rect 5167 -74559 5179 -74183
rect 5213 -74559 5225 -74183
rect 5167 -74571 5225 -74559
rect 5425 -74183 5483 -74171
rect 5425 -74559 5437 -74183
rect 5471 -74559 5483 -74183
rect 5425 -74571 5483 -74559
rect 5683 -74183 5741 -74171
rect 5683 -74559 5695 -74183
rect 5729 -74559 5741 -74183
rect 5683 -74571 5741 -74559
rect 5941 -74183 5999 -74171
rect 5941 -74559 5953 -74183
rect 5987 -74559 5999 -74183
rect 5941 -74571 5999 -74559
rect 6199 -74183 6257 -74171
rect 6199 -74559 6211 -74183
rect 6245 -74559 6257 -74183
rect 6199 -74571 6257 -74559
<< ndiffc >>
rect 56180 -42005 56214 -41971
rect 56180 -42073 56214 -42039
rect 56264 -42005 56298 -41971
rect 56264 -42073 56298 -42039
rect 56456 -42005 56490 -41971
rect 56456 -42073 56490 -42039
rect 56540 -42005 56574 -41971
rect 56540 -42073 56574 -42039
rect 56695 -42009 56729 -41975
rect 56695 -42077 56729 -42043
rect 56863 -42009 56897 -41975
rect 56863 -42077 56897 -42043
rect 57153 -42009 57187 -41975
rect 57153 -42077 57187 -42043
rect 57321 -42009 57355 -41975
rect 57321 -42077 57355 -42043
rect 57476 -42005 57510 -41971
rect 57476 -42073 57510 -42039
rect 57560 -42005 57594 -41971
rect 57560 -42073 57594 -42039
rect 57752 -42005 57786 -41971
rect 57752 -42073 57786 -42039
rect 57836 -42005 57870 -41971
rect 57836 -42073 57870 -42039
rect 56016 -42890 56050 -42714
rect 56134 -42890 56168 -42714
rect 56562 -42804 56596 -42628
rect 56680 -42804 56714 -42628
rect 56798 -42804 56832 -42628
rect 56916 -42804 56950 -42628
rect 57034 -42804 57068 -42628
rect 57152 -42804 57186 -42628
rect 57270 -42804 57304 -42628
rect 57388 -42804 57422 -42628
rect 57506 -42804 57540 -42628
rect 12262 -57671 12296 -57637
rect 12262 -57739 12296 -57705
rect 12346 -57671 12380 -57637
rect 12346 -57739 12380 -57705
rect 10410 -58034 10444 -57858
rect 10668 -58034 10702 -57858
rect 10926 -58034 10960 -57858
rect 11184 -58034 11218 -57858
rect 11442 -58034 11476 -57858
rect 11700 -58034 11734 -57858
rect 11958 -58034 11992 -57858
rect 16260 -45078 16294 -44502
rect 17278 -45078 17312 -44502
rect 18296 -45078 18330 -44502
rect 19314 -45078 19348 -44502
rect 20332 -45078 20366 -44502
rect 21350 -45078 21384 -44502
rect 22368 -45078 22402 -44502
rect 23386 -45078 23420 -44502
rect 24404 -45078 24438 -44502
rect 25422 -45078 25456 -44502
rect 28026 -44602 28060 -44026
rect 29044 -44602 29078 -44026
rect 30062 -44602 30096 -44026
rect 31080 -44602 31114 -44026
rect 32098 -44602 32132 -44026
rect 33116 -44602 33150 -44026
rect 34134 -44602 34168 -44026
rect 35152 -44602 35186 -44026
rect 36170 -44602 36204 -44026
rect 37188 -44602 37222 -44026
rect 38206 -44602 38240 -44026
rect 39224 -44602 39258 -44026
rect 40242 -44602 40276 -44026
rect 41260 -44602 41294 -44026
rect 42278 -44602 42312 -44026
rect 43296 -44602 43330 -44026
rect 44314 -44602 44348 -44026
rect 45332 -44602 45366 -44026
rect 46350 -44602 46384 -44026
rect 47368 -44602 47402 -44026
rect 48386 -44602 48420 -44026
rect 16260 -45896 16294 -45320
rect 17278 -45896 17312 -45320
rect 18296 -45896 18330 -45320
rect 19314 -45896 19348 -45320
rect 20332 -45896 20366 -45320
rect 21350 -45896 21384 -45320
rect 22368 -45896 22402 -45320
rect 23386 -45896 23420 -45320
rect 24404 -45896 24438 -45320
rect 25422 -45896 25456 -45320
rect 28026 -45420 28060 -44844
rect 29044 -45420 29078 -44844
rect 30062 -45420 30096 -44844
rect 31080 -45420 31114 -44844
rect 32098 -45420 32132 -44844
rect 33116 -45420 33150 -44844
rect 34134 -45420 34168 -44844
rect 35152 -45420 35186 -44844
rect 36170 -45420 36204 -44844
rect 37188 -45420 37222 -44844
rect 38206 -45420 38240 -44844
rect 39224 -45420 39258 -44844
rect 40242 -45420 40276 -44844
rect 41260 -45420 41294 -44844
rect 42278 -45420 42312 -44844
rect 43296 -45420 43330 -44844
rect 44314 -45420 44348 -44844
rect 45332 -45420 45366 -44844
rect 46350 -45420 46384 -44844
rect 47368 -45420 47402 -44844
rect 48386 -45420 48420 -44844
rect 16260 -46714 16294 -46138
rect 17278 -46714 17312 -46138
rect 18296 -46714 18330 -46138
rect 19314 -46714 19348 -46138
rect 20332 -46714 20366 -46138
rect 21350 -46714 21384 -46138
rect 22368 -46714 22402 -46138
rect 23386 -46714 23420 -46138
rect 24404 -46714 24438 -46138
rect 25422 -46714 25456 -46138
rect 28026 -46798 28060 -46222
rect 29044 -46798 29078 -46222
rect 30062 -46798 30096 -46222
rect 31080 -46798 31114 -46222
rect 32098 -46798 32132 -46222
rect 33116 -46798 33150 -46222
rect 34134 -46798 34168 -46222
rect 35152 -46798 35186 -46222
rect 36170 -46798 36204 -46222
rect 37188 -46798 37222 -46222
rect 38206 -46798 38240 -46222
rect 39224 -46798 39258 -46222
rect 40242 -46798 40276 -46222
rect 41260 -46798 41294 -46222
rect 42278 -46798 42312 -46222
rect 43296 -46798 43330 -46222
rect 44314 -46798 44348 -46222
rect 45332 -46798 45366 -46222
rect 46350 -46798 46384 -46222
rect 47368 -46798 47402 -46222
rect 48386 -46798 48420 -46222
rect 16260 -47532 16294 -46956
rect 17278 -47532 17312 -46956
rect 18296 -47532 18330 -46956
rect 19314 -47532 19348 -46956
rect 20332 -47532 20366 -46956
rect 21350 -47532 21384 -46956
rect 22368 -47532 22402 -46956
rect 23386 -47532 23420 -46956
rect 24404 -47532 24438 -46956
rect 25422 -47532 25456 -46956
rect 16260 -48350 16294 -47774
rect 17278 -48350 17312 -47774
rect 18296 -48350 18330 -47774
rect 19314 -48350 19348 -47774
rect 20332 -48350 20366 -47774
rect 21350 -48350 21384 -47774
rect 22368 -48350 22402 -47774
rect 23386 -48350 23420 -47774
rect 24404 -48350 24438 -47774
rect 25422 -48350 25456 -47774
rect 28026 -48030 28060 -47454
rect 29044 -48030 29078 -47454
rect 30062 -48030 30096 -47454
rect 31080 -48030 31114 -47454
rect 32098 -48030 32132 -47454
rect 33116 -48030 33150 -47454
rect 34134 -48030 34168 -47454
rect 35152 -48030 35186 -47454
rect 36170 -48030 36204 -47454
rect 37188 -48030 37222 -47454
rect 38206 -48030 38240 -47454
rect 39224 -48030 39258 -47454
rect 40242 -48030 40276 -47454
rect 41260 -48030 41294 -47454
rect 42278 -48030 42312 -47454
rect 43296 -48030 43330 -47454
rect 44314 -48030 44348 -47454
rect 45332 -48030 45366 -47454
rect 46350 -48030 46384 -47454
rect 47368 -48030 47402 -47454
rect 48386 -48030 48420 -47454
rect 16260 -49168 16294 -48592
rect 17278 -49168 17312 -48592
rect 18296 -49168 18330 -48592
rect 19314 -49168 19348 -48592
rect 20332 -49168 20366 -48592
rect 21350 -49168 21384 -48592
rect 22368 -49168 22402 -48592
rect 23386 -49168 23420 -48592
rect 24404 -49168 24438 -48592
rect 25422 -49168 25456 -48592
rect 28024 -49264 28058 -48688
rect 29042 -49264 29076 -48688
rect 30060 -49264 30094 -48688
rect 31078 -49264 31112 -48688
rect 32096 -49264 32130 -48688
rect 33114 -49264 33148 -48688
rect 34132 -49264 34166 -48688
rect 35150 -49264 35184 -48688
rect 36168 -49264 36202 -48688
rect 37186 -49264 37220 -48688
rect 38204 -49264 38238 -48688
rect 39222 -49264 39256 -48688
rect 40240 -49264 40274 -48688
rect 41258 -49264 41292 -48688
rect 42276 -49264 42310 -48688
rect 43294 -49264 43328 -48688
rect 44312 -49264 44346 -48688
rect 45330 -49264 45364 -48688
rect 46348 -49264 46382 -48688
rect 47366 -49264 47400 -48688
rect 48384 -49264 48418 -48688
rect 16260 -49986 16294 -49410
rect 17278 -49986 17312 -49410
rect 18296 -49986 18330 -49410
rect 19314 -49986 19348 -49410
rect 20332 -49986 20366 -49410
rect 21350 -49986 21384 -49410
rect 22368 -49986 22402 -49410
rect 23386 -49986 23420 -49410
rect 24404 -49986 24438 -49410
rect 25422 -49986 25456 -49410
rect 16260 -50804 16294 -50228
rect 17278 -50804 17312 -50228
rect 18296 -50804 18330 -50228
rect 19314 -50804 19348 -50228
rect 20332 -50804 20366 -50228
rect 21350 -50804 21384 -50228
rect 22368 -50804 22402 -50228
rect 23386 -50804 23420 -50228
rect 24404 -50804 24438 -50228
rect 25422 -50804 25456 -50228
rect 28024 -50498 28058 -49922
rect 29042 -50498 29076 -49922
rect 30060 -50498 30094 -49922
rect 31078 -50498 31112 -49922
rect 32096 -50498 32130 -49922
rect 33114 -50498 33148 -49922
rect 34132 -50498 34166 -49922
rect 35150 -50498 35184 -49922
rect 36168 -50498 36202 -49922
rect 37186 -50498 37220 -49922
rect 38204 -50498 38238 -49922
rect 39222 -50498 39256 -49922
rect 40240 -50498 40274 -49922
rect 41258 -50498 41292 -49922
rect 42276 -50498 42310 -49922
rect 43294 -50498 43328 -49922
rect 44312 -50498 44346 -49922
rect 45330 -50498 45364 -49922
rect 46348 -50498 46382 -49922
rect 47366 -50498 47400 -49922
rect 48384 -50498 48418 -49922
rect 28024 -51730 28058 -51154
rect 29042 -51730 29076 -51154
rect 30060 -51730 30094 -51154
rect 31078 -51730 31112 -51154
rect 32096 -51730 32130 -51154
rect 33114 -51730 33148 -51154
rect 34132 -51730 34166 -51154
rect 35150 -51730 35184 -51154
rect 36168 -51730 36202 -51154
rect 37186 -51730 37220 -51154
rect 38204 -51730 38238 -51154
rect 39222 -51730 39256 -51154
rect 40240 -51730 40274 -51154
rect 41258 -51730 41292 -51154
rect 42276 -51730 42310 -51154
rect 43294 -51730 43328 -51154
rect 44312 -51730 44346 -51154
rect 45330 -51730 45364 -51154
rect 46348 -51730 46382 -51154
rect 47366 -51730 47400 -51154
rect 48384 -51730 48418 -51154
rect 14936 -52828 14970 -52252
rect 15954 -52828 15988 -52252
rect 16972 -52828 17006 -52252
rect 17990 -52828 18024 -52252
rect 19008 -52828 19042 -52252
rect 20026 -52828 20060 -52252
rect 21044 -52828 21078 -52252
rect 22062 -52828 22096 -52252
rect 23080 -52828 23114 -52252
rect 24098 -52828 24132 -52252
rect 25116 -52828 25150 -52252
rect 26134 -52828 26168 -52252
rect 28024 -52964 28058 -52388
rect 29042 -52964 29076 -52388
rect 30060 -52964 30094 -52388
rect 31078 -52964 31112 -52388
rect 32096 -52964 32130 -52388
rect 33114 -52964 33148 -52388
rect 34132 -52964 34166 -52388
rect 35150 -52964 35184 -52388
rect 36168 -52964 36202 -52388
rect 37186 -52964 37220 -52388
rect 38204 -52964 38238 -52388
rect 39222 -52964 39256 -52388
rect 40240 -52964 40274 -52388
rect 41258 -52964 41292 -52388
rect 42276 -52964 42310 -52388
rect 43294 -52964 43328 -52388
rect 44312 -52964 44346 -52388
rect 45330 -52964 45364 -52388
rect 46348 -52964 46382 -52388
rect 47366 -52964 47400 -52388
rect 48384 -52964 48418 -52388
rect 14936 -53940 14970 -53364
rect 15954 -53940 15988 -53364
rect 16972 -53940 17006 -53364
rect 17990 -53940 18024 -53364
rect 19008 -53940 19042 -53364
rect 20026 -53940 20060 -53364
rect 21044 -53940 21078 -53364
rect 22062 -53940 22096 -53364
rect 23080 -53940 23114 -53364
rect 24098 -53940 24132 -53364
rect 25116 -53940 25150 -53364
rect 26134 -53940 26168 -53364
rect 28024 -54198 28058 -53622
rect 29042 -54198 29076 -53622
rect 30060 -54198 30094 -53622
rect 31078 -54198 31112 -53622
rect 32096 -54198 32130 -53622
rect 33114 -54198 33148 -53622
rect 34132 -54198 34166 -53622
rect 35150 -54198 35184 -53622
rect 36168 -54198 36202 -53622
rect 37186 -54198 37220 -53622
rect 38204 -54198 38238 -53622
rect 39222 -54198 39256 -53622
rect 40240 -54198 40274 -53622
rect 41258 -54198 41292 -53622
rect 42276 -54198 42310 -53622
rect 43294 -54198 43328 -53622
rect 44312 -54198 44346 -53622
rect 45330 -54198 45364 -53622
rect 46348 -54198 46382 -53622
rect 47366 -54198 47400 -53622
rect 48384 -54198 48418 -53622
rect 14936 -55052 14970 -54476
rect 15954 -55052 15988 -54476
rect 16972 -55052 17006 -54476
rect 17990 -55052 18024 -54476
rect 19008 -55052 19042 -54476
rect 20026 -55052 20060 -54476
rect 21044 -55052 21078 -54476
rect 22062 -55052 22096 -54476
rect 23080 -55052 23114 -54476
rect 24098 -55052 24132 -54476
rect 25116 -55052 25150 -54476
rect 26134 -55052 26168 -54476
rect 28024 -55430 28058 -54854
rect 29042 -55430 29076 -54854
rect 30060 -55430 30094 -54854
rect 31078 -55430 31112 -54854
rect 32096 -55430 32130 -54854
rect 33114 -55430 33148 -54854
rect 34132 -55430 34166 -54854
rect 35150 -55430 35184 -54854
rect 36168 -55430 36202 -54854
rect 37186 -55430 37220 -54854
rect 38204 -55430 38238 -54854
rect 39222 -55430 39256 -54854
rect 40240 -55430 40274 -54854
rect 41258 -55430 41292 -54854
rect 42276 -55430 42310 -54854
rect 43294 -55430 43328 -54854
rect 44312 -55430 44346 -54854
rect 45330 -55430 45364 -54854
rect 46348 -55430 46382 -54854
rect 47366 -55430 47400 -54854
rect 48384 -55430 48418 -54854
rect 14936 -56164 14970 -55588
rect 15954 -56164 15988 -55588
rect 16972 -56164 17006 -55588
rect 17990 -56164 18024 -55588
rect 19008 -56164 19042 -55588
rect 20026 -56164 20060 -55588
rect 21044 -56164 21078 -55588
rect 22062 -56164 22096 -55588
rect 23080 -56164 23114 -55588
rect 24098 -56164 24132 -55588
rect 25116 -56164 25150 -55588
rect 26134 -56164 26168 -55588
rect 28024 -56664 28058 -56088
rect 29042 -56664 29076 -56088
rect 30060 -56664 30094 -56088
rect 31078 -56664 31112 -56088
rect 32096 -56664 32130 -56088
rect 33114 -56664 33148 -56088
rect 34132 -56664 34166 -56088
rect 35150 -56664 35184 -56088
rect 36168 -56664 36202 -56088
rect 37186 -56664 37220 -56088
rect 38204 -56664 38238 -56088
rect 39222 -56664 39256 -56088
rect 40240 -56664 40274 -56088
rect 41258 -56664 41292 -56088
rect 42276 -56664 42310 -56088
rect 43294 -56664 43328 -56088
rect 44312 -56664 44346 -56088
rect 45330 -56664 45364 -56088
rect 46348 -56664 46382 -56088
rect 47366 -56664 47400 -56088
rect 48384 -56664 48418 -56088
rect 15394 -57706 15428 -57130
rect 16412 -57706 16446 -57130
rect 17430 -57706 17464 -57130
rect 18448 -57706 18482 -57130
rect 19466 -57706 19500 -57130
rect 20484 -57706 20518 -57130
rect 21502 -57706 21536 -57130
rect 22520 -57706 22554 -57130
rect 23538 -57706 23572 -57130
rect 24556 -57706 24590 -57130
rect 25574 -57706 25608 -57130
rect 28024 -57896 28058 -57320
rect 29042 -57896 29076 -57320
rect 30060 -57896 30094 -57320
rect 31078 -57896 31112 -57320
rect 32096 -57896 32130 -57320
rect 33114 -57896 33148 -57320
rect 34132 -57896 34166 -57320
rect 35150 -57896 35184 -57320
rect 36168 -57896 36202 -57320
rect 37186 -57896 37220 -57320
rect 38204 -57896 38238 -57320
rect 39222 -57896 39256 -57320
rect 40240 -57896 40274 -57320
rect 41258 -57896 41292 -57320
rect 42276 -57896 42310 -57320
rect 43294 -57896 43328 -57320
rect 44312 -57896 44346 -57320
rect 45330 -57896 45364 -57320
rect 46348 -57896 46382 -57320
rect 47366 -57896 47400 -57320
rect 48384 -57896 48418 -57320
rect 57920 -42890 57954 -42714
rect 58038 -42890 58072 -42714
rect -27996 -67695 -27962 -67661
rect -27996 -67763 -27962 -67729
rect -27912 -67695 -27878 -67661
rect -27912 -67763 -27878 -67729
rect -23996 -67695 -23962 -67661
rect -23996 -67763 -23962 -67729
rect -23912 -67695 -23878 -67661
rect -23912 -67763 -23878 -67729
rect -19996 -67695 -19962 -67661
rect -19996 -67763 -19962 -67729
rect -27342 -68706 -27308 -68330
rect -27084 -68706 -27050 -68330
rect -26826 -68706 -26792 -68330
rect -26568 -68706 -26534 -68330
rect -26310 -68706 -26276 -68330
rect -26052 -68706 -26018 -68330
rect -25794 -68706 -25760 -68330
rect -19912 -67695 -19878 -67661
rect -19912 -67763 -19878 -67729
rect -15996 -67695 -15962 -67661
rect -15996 -67763 -15962 -67729
rect -23342 -68706 -23308 -68330
rect -23084 -68706 -23050 -68330
rect -22826 -68706 -22792 -68330
rect -22568 -68706 -22534 -68330
rect -22310 -68706 -22276 -68330
rect -22052 -68706 -22018 -68330
rect -21794 -68706 -21760 -68330
rect -15912 -67695 -15878 -67661
rect -15912 -67763 -15878 -67729
rect -11996 -67695 -11962 -67661
rect -11996 -67763 -11962 -67729
rect -19342 -68706 -19308 -68330
rect -19084 -68706 -19050 -68330
rect -18826 -68706 -18792 -68330
rect -18568 -68706 -18534 -68330
rect -18310 -68706 -18276 -68330
rect -18052 -68706 -18018 -68330
rect -17794 -68706 -17760 -68330
rect -11912 -67695 -11878 -67661
rect -11912 -67763 -11878 -67729
rect -7996 -67695 -7962 -67661
rect -7996 -67763 -7962 -67729
rect -15342 -68706 -15308 -68330
rect -15084 -68706 -15050 -68330
rect -14826 -68706 -14792 -68330
rect -14568 -68706 -14534 -68330
rect -14310 -68706 -14276 -68330
rect -14052 -68706 -14018 -68330
rect -13794 -68706 -13760 -68330
rect -7912 -67695 -7878 -67661
rect -7912 -67763 -7878 -67729
rect -3996 -67695 -3962 -67661
rect -3996 -67763 -3962 -67729
rect -11342 -68706 -11308 -68330
rect -11084 -68706 -11050 -68330
rect -10826 -68706 -10792 -68330
rect -10568 -68706 -10534 -68330
rect -10310 -68706 -10276 -68330
rect -10052 -68706 -10018 -68330
rect -9794 -68706 -9760 -68330
rect -3912 -67695 -3878 -67661
rect -3912 -67763 -3878 -67729
rect 4 -67695 38 -67661
rect 4 -67763 38 -67729
rect -7342 -68706 -7308 -68330
rect -7084 -68706 -7050 -68330
rect -6826 -68706 -6792 -68330
rect -6568 -68706 -6534 -68330
rect -6310 -68706 -6276 -68330
rect -6052 -68706 -6018 -68330
rect -5794 -68706 -5760 -68330
rect 88 -67695 122 -67661
rect 88 -67763 122 -67729
rect 4004 -67695 4038 -67661
rect 4004 -67763 4038 -67729
rect -3342 -68706 -3308 -68330
rect -3084 -68706 -3050 -68330
rect -2826 -68706 -2792 -68330
rect -2568 -68706 -2534 -68330
rect -2310 -68706 -2276 -68330
rect -2052 -68706 -2018 -68330
rect -1794 -68706 -1760 -68330
rect 4088 -67695 4122 -67661
rect 4088 -67763 4122 -67729
rect 658 -68706 692 -68330
rect 916 -68706 950 -68330
rect 1174 -68706 1208 -68330
rect 1432 -68706 1466 -68330
rect 1690 -68706 1724 -68330
rect 1948 -68706 1982 -68330
rect 2206 -68706 2240 -68330
rect 4658 -68706 4692 -68330
rect 4916 -68706 4950 -68330
rect 5174 -68706 5208 -68330
rect 5432 -68706 5466 -68330
rect 5690 -68706 5724 -68330
rect 5948 -68706 5982 -68330
rect 6206 -68706 6240 -68330
rect -27342 -71866 -27308 -71490
rect -27084 -71866 -27050 -71490
rect -26826 -71866 -26792 -71490
rect -26568 -71866 -26534 -71490
rect -26310 -71866 -26276 -71490
rect -26052 -71866 -26018 -71490
rect -25794 -71866 -25760 -71490
rect -27996 -72467 -27962 -72433
rect -27996 -72535 -27962 -72501
rect -23342 -71866 -23308 -71490
rect -23084 -71866 -23050 -71490
rect -22826 -71866 -22792 -71490
rect -22568 -71866 -22534 -71490
rect -22310 -71866 -22276 -71490
rect -22052 -71866 -22018 -71490
rect -21794 -71866 -21760 -71490
rect -27912 -72467 -27878 -72433
rect -27912 -72535 -27878 -72501
rect -23996 -72467 -23962 -72433
rect -23996 -72535 -23962 -72501
rect -19342 -71866 -19308 -71490
rect -19084 -71866 -19050 -71490
rect -18826 -71866 -18792 -71490
rect -18568 -71866 -18534 -71490
rect -18310 -71866 -18276 -71490
rect -18052 -71866 -18018 -71490
rect -17794 -71866 -17760 -71490
rect -23912 -72467 -23878 -72433
rect -23912 -72535 -23878 -72501
rect -19996 -72467 -19962 -72433
rect -19996 -72535 -19962 -72501
rect -15342 -71866 -15308 -71490
rect -15084 -71866 -15050 -71490
rect -14826 -71866 -14792 -71490
rect -14568 -71866 -14534 -71490
rect -14310 -71866 -14276 -71490
rect -14052 -71866 -14018 -71490
rect -13794 -71866 -13760 -71490
rect -19912 -72467 -19878 -72433
rect -19912 -72535 -19878 -72501
rect -15996 -72467 -15962 -72433
rect -15996 -72535 -15962 -72501
rect -11342 -71866 -11308 -71490
rect -11084 -71866 -11050 -71490
rect -10826 -71866 -10792 -71490
rect -10568 -71866 -10534 -71490
rect -10310 -71866 -10276 -71490
rect -10052 -71866 -10018 -71490
rect -9794 -71866 -9760 -71490
rect -15912 -72467 -15878 -72433
rect -15912 -72535 -15878 -72501
rect -11996 -72467 -11962 -72433
rect -11996 -72535 -11962 -72501
rect -7342 -71866 -7308 -71490
rect -7084 -71866 -7050 -71490
rect -6826 -71866 -6792 -71490
rect -6568 -71866 -6534 -71490
rect -6310 -71866 -6276 -71490
rect -6052 -71866 -6018 -71490
rect -5794 -71866 -5760 -71490
rect -11912 -72467 -11878 -72433
rect -11912 -72535 -11878 -72501
rect -7996 -72467 -7962 -72433
rect -7996 -72535 -7962 -72501
rect -3342 -71866 -3308 -71490
rect -3084 -71866 -3050 -71490
rect -2826 -71866 -2792 -71490
rect -2568 -71866 -2534 -71490
rect -2310 -71866 -2276 -71490
rect -2052 -71866 -2018 -71490
rect -1794 -71866 -1760 -71490
rect -7912 -72467 -7878 -72433
rect -7912 -72535 -7878 -72501
rect -3996 -72467 -3962 -72433
rect -3996 -72535 -3962 -72501
rect 658 -71866 692 -71490
rect 916 -71866 950 -71490
rect 1174 -71866 1208 -71490
rect 1432 -71866 1466 -71490
rect 1690 -71866 1724 -71490
rect 1948 -71866 1982 -71490
rect 2206 -71866 2240 -71490
rect -3912 -72467 -3878 -72433
rect -3912 -72535 -3878 -72501
rect 4 -72467 38 -72433
rect 4 -72535 38 -72501
rect 4658 -71866 4692 -71490
rect 4916 -71866 4950 -71490
rect 5174 -71866 5208 -71490
rect 5432 -71866 5466 -71490
rect 5690 -71866 5724 -71490
rect 5948 -71866 5982 -71490
rect 6206 -71866 6240 -71490
rect 88 -72467 122 -72433
rect 88 -72535 122 -72501
rect 4004 -72467 4038 -72433
rect 4004 -72535 4038 -72501
rect 4088 -72467 4122 -72433
rect 4088 -72535 4122 -72501
<< pdiffc >>
rect 31932 -31092 31966 -30516
rect 32950 -31092 32984 -30516
rect 33968 -31092 34002 -30516
rect 34986 -31092 35020 -30516
rect 36004 -31092 36038 -30516
rect 37022 -31092 37056 -30516
rect 38040 -31092 38074 -30516
rect 39058 -31092 39092 -30516
rect 40076 -31092 40110 -30516
rect 41094 -31092 41128 -30516
rect 42112 -31092 42146 -30516
rect 43130 -31092 43164 -30516
rect 44148 -31092 44182 -30516
rect 45166 -31092 45200 -30516
rect 46184 -31092 46218 -30516
rect 47202 -31092 47236 -30516
rect 48220 -31092 48254 -30516
rect 31932 -32228 31966 -31652
rect 32950 -32228 32984 -31652
rect 33968 -32228 34002 -31652
rect 34986 -32228 35020 -31652
rect 36004 -32228 36038 -31652
rect 37022 -32228 37056 -31652
rect 38040 -32228 38074 -31652
rect 39058 -32228 39092 -31652
rect 40076 -32228 40110 -31652
rect 41094 -32228 41128 -31652
rect 42112 -32228 42146 -31652
rect 43130 -32228 43164 -31652
rect 44148 -32228 44182 -31652
rect 45166 -32228 45200 -31652
rect 46184 -32228 46218 -31652
rect 47202 -32228 47236 -31652
rect 48220 -32228 48254 -31652
rect 31932 -33364 31966 -32788
rect 32950 -33364 32984 -32788
rect 33968 -33364 34002 -32788
rect 34986 -33364 35020 -32788
rect 36004 -33364 36038 -32788
rect 37022 -33364 37056 -32788
rect 38040 -33364 38074 -32788
rect 39058 -33364 39092 -32788
rect 40076 -33364 40110 -32788
rect 41094 -33364 41128 -32788
rect 42112 -33364 42146 -32788
rect 43130 -33364 43164 -32788
rect 44148 -33364 44182 -32788
rect 45166 -33364 45200 -32788
rect 46184 -33364 46218 -32788
rect 47202 -33364 47236 -32788
rect 48220 -33364 48254 -32788
rect 33126 -35002 33160 -34426
rect 34144 -35002 34178 -34426
rect 35162 -35002 35196 -34426
rect 36180 -35002 36214 -34426
rect 37198 -35002 37232 -34426
rect 38216 -35002 38250 -34426
rect 39234 -35002 39268 -34426
rect 40252 -35002 40286 -34426
rect 41270 -35002 41304 -34426
rect 42288 -35002 42322 -34426
rect 43306 -35002 43340 -34426
rect 44324 -35002 44358 -34426
rect 45342 -35002 45376 -34426
rect 46360 -35002 46394 -34426
rect 47378 -35002 47412 -34426
rect 33126 -36034 33160 -35458
rect 34144 -36034 34178 -35458
rect 35162 -36034 35196 -35458
rect 36180 -36034 36214 -35458
rect 37198 -36034 37232 -35458
rect 38216 -36034 38250 -35458
rect 39234 -36034 39268 -35458
rect 40252 -36034 40286 -35458
rect 41270 -36034 41304 -35458
rect 42288 -36034 42322 -35458
rect 43306 -36034 43340 -35458
rect 44324 -36034 44358 -35458
rect 45342 -36034 45376 -35458
rect 46360 -36034 46394 -35458
rect 47378 -36034 47412 -35458
rect 27614 -37742 27648 -37166
rect 28632 -37742 28666 -37166
rect 29650 -37742 29684 -37166
rect 30668 -37742 30702 -37166
rect 31686 -37742 31720 -37166
rect 32918 -37638 32952 -37062
rect 33936 -37638 33970 -37062
rect 34954 -37638 34988 -37062
rect 35972 -37638 36006 -37062
rect 36990 -37638 37024 -37062
rect 38008 -37638 38042 -37062
rect 39026 -37638 39060 -37062
rect 40044 -37638 40078 -37062
rect 41062 -37638 41096 -37062
rect 42080 -37638 42114 -37062
rect 43098 -37638 43132 -37062
rect 44116 -37638 44150 -37062
rect 45134 -37638 45168 -37062
rect 46152 -37638 46186 -37062
rect 47170 -37638 47204 -37062
rect 48188 -37638 48222 -37062
rect 27614 -38774 27648 -38198
rect 28632 -38774 28666 -38198
rect 29650 -38774 29684 -38198
rect 30668 -38774 30702 -38198
rect 31686 -38774 31720 -38198
rect 32918 -38894 32952 -38318
rect 33936 -38894 33970 -38318
rect 34954 -38894 34988 -38318
rect 35972 -38894 36006 -38318
rect 36990 -38894 37024 -38318
rect 38008 -38894 38042 -38318
rect 39026 -38894 39060 -38318
rect 40044 -38894 40078 -38318
rect 41062 -38894 41096 -38318
rect 42080 -38894 42114 -38318
rect 43098 -38894 43132 -38318
rect 44116 -38894 44150 -38318
rect 45134 -38894 45168 -38318
rect 46152 -38894 46186 -38318
rect 47170 -38894 47204 -38318
rect 48188 -38894 48222 -38318
rect 27614 -39806 27648 -39230
rect 28632 -39806 28666 -39230
rect 29650 -39806 29684 -39230
rect 30668 -39806 30702 -39230
rect 31686 -39806 31720 -39230
rect 32918 -40150 32952 -39574
rect 33936 -40150 33970 -39574
rect 34954 -40150 34988 -39574
rect 35972 -40150 36006 -39574
rect 36990 -40150 37024 -39574
rect 38008 -40150 38042 -39574
rect 39026 -40150 39060 -39574
rect 40044 -40150 40078 -39574
rect 41062 -40150 41096 -39574
rect 42080 -40150 42114 -39574
rect 43098 -40150 43132 -39574
rect 44116 -40150 44150 -39574
rect 45134 -40150 45168 -39574
rect 46152 -40150 46186 -39574
rect 47170 -40150 47204 -39574
rect 48188 -40150 48222 -39574
rect 27614 -40838 27648 -40262
rect 28632 -40838 28666 -40262
rect 29650 -40838 29684 -40262
rect 30668 -40838 30702 -40262
rect 31686 -40838 31720 -40262
rect 32918 -41406 32952 -40830
rect 33936 -41406 33970 -40830
rect 34954 -41406 34988 -40830
rect 35972 -41406 36006 -40830
rect 36990 -41406 37024 -40830
rect 38008 -41406 38042 -40830
rect 39026 -41406 39060 -40830
rect 40044 -41406 40078 -40830
rect 41062 -41406 41096 -40830
rect 42080 -41406 42114 -40830
rect 43098 -41406 43132 -40830
rect 44116 -41406 44150 -40830
rect 45134 -41406 45168 -40830
rect 46152 -41406 46186 -40830
rect 47170 -41406 47204 -40830
rect 48188 -41406 48222 -40830
rect 52442 -39868 52476 -39692
rect 52900 -39868 52934 -39692
rect 53358 -39868 53392 -39692
rect 53816 -39868 53850 -39692
rect 54274 -39868 54308 -39692
rect 54732 -39868 54766 -39692
rect 55190 -39868 55224 -39692
rect 52501 -40951 52535 -40575
rect 52759 -40951 52793 -40575
rect 53017 -40951 53051 -40575
rect 53275 -40951 53309 -40575
rect 53533 -40951 53567 -40575
rect 53791 -40951 53825 -40575
rect 54049 -40951 54083 -40575
rect 54307 -40951 54341 -40575
rect 54565 -40951 54599 -40575
rect 54823 -40951 54857 -40575
rect 55081 -40951 55115 -40575
rect 52501 -41811 52535 -41435
rect 52759 -41811 52793 -41435
rect 53017 -41811 53051 -41435
rect 53275 -41811 53309 -41435
rect 53533 -41811 53567 -41435
rect 53791 -41811 53825 -41435
rect 54049 -41811 54083 -41435
rect 54307 -41811 54341 -41435
rect 54565 -41811 54599 -41435
rect 54823 -41811 54857 -41435
rect 55081 -41811 55115 -41435
rect 56070 -40268 56104 -39892
rect 56328 -40268 56362 -39892
rect 56586 -40268 56620 -39892
rect 56844 -40268 56878 -39892
rect 57102 -40268 57136 -39892
rect 57360 -40268 57394 -39892
rect 57618 -40268 57652 -39892
rect 57876 -40268 57910 -39892
rect 56070 -41128 56104 -40752
rect 56328 -41128 56362 -40752
rect 56586 -41128 56620 -40752
rect 56844 -41128 56878 -40752
rect 57102 -41128 57136 -40752
rect 57360 -41128 57394 -40752
rect 57618 -41128 57652 -40752
rect 57876 -41128 57910 -40752
rect 56180 -41685 56214 -41651
rect 56180 -41753 56214 -41719
rect 56180 -41821 56214 -41787
rect 56264 -41685 56298 -41651
rect 56264 -41753 56298 -41719
rect 56264 -41821 56298 -41787
rect 56456 -41685 56490 -41651
rect 56456 -41753 56490 -41719
rect 56456 -41821 56490 -41787
rect 56540 -41685 56574 -41651
rect 56540 -41753 56574 -41719
rect 56540 -41821 56574 -41787
rect 56695 -41685 56729 -41651
rect 56695 -41753 56729 -41719
rect 56695 -41821 56729 -41787
rect 56779 -41685 56813 -41651
rect 56779 -41753 56813 -41719
rect 56779 -41821 56813 -41787
rect 56863 -41685 56897 -41651
rect 56863 -41753 56897 -41719
rect 56863 -41821 56897 -41787
rect 57153 -41685 57187 -41651
rect 57153 -41753 57187 -41719
rect 57153 -41821 57187 -41787
rect 57237 -41685 57271 -41651
rect 57237 -41753 57271 -41719
rect 57237 -41821 57271 -41787
rect 57321 -41685 57355 -41651
rect 57321 -41753 57355 -41719
rect 57321 -41821 57355 -41787
rect 57476 -41685 57510 -41651
rect 57476 -41753 57510 -41719
rect 57476 -41821 57510 -41787
rect 57560 -41685 57594 -41651
rect 57560 -41753 57594 -41719
rect 57560 -41821 57594 -41787
rect 57752 -41685 57786 -41651
rect 57752 -41753 57786 -41719
rect 57752 -41821 57786 -41787
rect 57836 -41685 57870 -41651
rect 57836 -41753 57870 -41719
rect 57836 -41821 57870 -41787
rect 54218 -42782 54252 -42606
rect 54346 -42782 54380 -42606
rect 54474 -42782 54508 -42606
rect 54602 -42782 54636 -42606
rect 54730 -42782 54764 -42606
rect 54858 -42782 54892 -42606
rect 54986 -42782 55020 -42606
rect 55114 -42782 55148 -42606
rect 55242 -42782 55276 -42606
rect 55370 -42782 55404 -42606
rect 10410 -57310 10444 -56934
rect 10668 -57310 10702 -56934
rect 10926 -57310 10960 -56934
rect 11184 -57310 11218 -56934
rect 11442 -57310 11476 -56934
rect 11700 -57310 11734 -56934
rect 11958 -57310 11992 -56934
rect 12262 -57351 12296 -57317
rect 12262 -57419 12296 -57385
rect 12262 -57487 12296 -57453
rect 12346 -57351 12380 -57317
rect 12346 -57419 12380 -57385
rect 12346 -57487 12380 -57453
rect -27996 -67375 -27962 -67341
rect -27996 -67443 -27962 -67409
rect -27996 -67511 -27962 -67477
rect -27912 -67375 -27878 -67341
rect -27912 -67443 -27878 -67409
rect -27912 -67511 -27878 -67477
rect -27337 -66013 -27303 -65637
rect -27079 -66013 -27045 -65637
rect -26821 -66013 -26787 -65637
rect -26563 -66013 -26529 -65637
rect -26305 -66013 -26271 -65637
rect -26047 -66013 -26013 -65637
rect -25789 -66013 -25755 -65637
rect -27337 -66873 -27303 -66497
rect -27079 -66873 -27045 -66497
rect -26821 -66873 -26787 -66497
rect -26563 -66873 -26529 -66497
rect -26305 -66873 -26271 -66497
rect -26047 -66873 -26013 -66497
rect -25789 -66873 -25755 -66497
rect -23996 -67375 -23962 -67341
rect -23996 -67443 -23962 -67409
rect -23996 -67511 -23962 -67477
rect -23912 -67375 -23878 -67341
rect -23912 -67443 -23878 -67409
rect -23912 -67511 -23878 -67477
rect -23337 -66013 -23303 -65637
rect -23079 -66013 -23045 -65637
rect -22821 -66013 -22787 -65637
rect -22563 -66013 -22529 -65637
rect -22305 -66013 -22271 -65637
rect -22047 -66013 -22013 -65637
rect -21789 -66013 -21755 -65637
rect -23337 -66873 -23303 -66497
rect -23079 -66873 -23045 -66497
rect -22821 -66873 -22787 -66497
rect -22563 -66873 -22529 -66497
rect -22305 -66873 -22271 -66497
rect -22047 -66873 -22013 -66497
rect -21789 -66873 -21755 -66497
rect -19996 -67375 -19962 -67341
rect -19996 -67443 -19962 -67409
rect -19996 -67511 -19962 -67477
rect -19912 -67375 -19878 -67341
rect -19912 -67443 -19878 -67409
rect -19912 -67511 -19878 -67477
rect -19337 -66013 -19303 -65637
rect -19079 -66013 -19045 -65637
rect -18821 -66013 -18787 -65637
rect -18563 -66013 -18529 -65637
rect -18305 -66013 -18271 -65637
rect -18047 -66013 -18013 -65637
rect -17789 -66013 -17755 -65637
rect -19337 -66873 -19303 -66497
rect -19079 -66873 -19045 -66497
rect -18821 -66873 -18787 -66497
rect -18563 -66873 -18529 -66497
rect -18305 -66873 -18271 -66497
rect -18047 -66873 -18013 -66497
rect -17789 -66873 -17755 -66497
rect -15996 -67375 -15962 -67341
rect -15996 -67443 -15962 -67409
rect -15996 -67511 -15962 -67477
rect -15912 -67375 -15878 -67341
rect -15912 -67443 -15878 -67409
rect -15912 -67511 -15878 -67477
rect -15337 -66013 -15303 -65637
rect -15079 -66013 -15045 -65637
rect -14821 -66013 -14787 -65637
rect -14563 -66013 -14529 -65637
rect -14305 -66013 -14271 -65637
rect -14047 -66013 -14013 -65637
rect -13789 -66013 -13755 -65637
rect -15337 -66873 -15303 -66497
rect -15079 -66873 -15045 -66497
rect -14821 -66873 -14787 -66497
rect -14563 -66873 -14529 -66497
rect -14305 -66873 -14271 -66497
rect -14047 -66873 -14013 -66497
rect -13789 -66873 -13755 -66497
rect -11996 -67375 -11962 -67341
rect -11996 -67443 -11962 -67409
rect -11996 -67511 -11962 -67477
rect -11912 -67375 -11878 -67341
rect -11912 -67443 -11878 -67409
rect -11912 -67511 -11878 -67477
rect -11337 -66013 -11303 -65637
rect -11079 -66013 -11045 -65637
rect -10821 -66013 -10787 -65637
rect -10563 -66013 -10529 -65637
rect -10305 -66013 -10271 -65637
rect -10047 -66013 -10013 -65637
rect -9789 -66013 -9755 -65637
rect -11337 -66873 -11303 -66497
rect -11079 -66873 -11045 -66497
rect -10821 -66873 -10787 -66497
rect -10563 -66873 -10529 -66497
rect -10305 -66873 -10271 -66497
rect -10047 -66873 -10013 -66497
rect -9789 -66873 -9755 -66497
rect -7996 -67375 -7962 -67341
rect -7996 -67443 -7962 -67409
rect -7996 -67511 -7962 -67477
rect -7912 -67375 -7878 -67341
rect -7912 -67443 -7878 -67409
rect -7912 -67511 -7878 -67477
rect -7337 -66013 -7303 -65637
rect -7079 -66013 -7045 -65637
rect -6821 -66013 -6787 -65637
rect -6563 -66013 -6529 -65637
rect -6305 -66013 -6271 -65637
rect -6047 -66013 -6013 -65637
rect -5789 -66013 -5755 -65637
rect -7337 -66873 -7303 -66497
rect -7079 -66873 -7045 -66497
rect -6821 -66873 -6787 -66497
rect -6563 -66873 -6529 -66497
rect -6305 -66873 -6271 -66497
rect -6047 -66873 -6013 -66497
rect -5789 -66873 -5755 -66497
rect -3996 -67375 -3962 -67341
rect -3996 -67443 -3962 -67409
rect -3996 -67511 -3962 -67477
rect -3912 -67375 -3878 -67341
rect -3912 -67443 -3878 -67409
rect -3912 -67511 -3878 -67477
rect -3337 -66013 -3303 -65637
rect -3079 -66013 -3045 -65637
rect -2821 -66013 -2787 -65637
rect -2563 -66013 -2529 -65637
rect -2305 -66013 -2271 -65637
rect -2047 -66013 -2013 -65637
rect -1789 -66013 -1755 -65637
rect -3337 -66873 -3303 -66497
rect -3079 -66873 -3045 -66497
rect -2821 -66873 -2787 -66497
rect -2563 -66873 -2529 -66497
rect -2305 -66873 -2271 -66497
rect -2047 -66873 -2013 -66497
rect -1789 -66873 -1755 -66497
rect 4 -67375 38 -67341
rect 4 -67443 38 -67409
rect 4 -67511 38 -67477
rect 88 -67375 122 -67341
rect 88 -67443 122 -67409
rect 88 -67511 122 -67477
rect 663 -66013 697 -65637
rect 921 -66013 955 -65637
rect 1179 -66013 1213 -65637
rect 1437 -66013 1471 -65637
rect 1695 -66013 1729 -65637
rect 1953 -66013 1987 -65637
rect 2211 -66013 2245 -65637
rect 663 -66873 697 -66497
rect 921 -66873 955 -66497
rect 1179 -66873 1213 -66497
rect 1437 -66873 1471 -66497
rect 1695 -66873 1729 -66497
rect 1953 -66873 1987 -66497
rect 2211 -66873 2245 -66497
rect 4004 -67375 4038 -67341
rect 4004 -67443 4038 -67409
rect 4004 -67511 4038 -67477
rect 4088 -67375 4122 -67341
rect 4088 -67443 4122 -67409
rect 4088 -67511 4122 -67477
rect 4663 -66013 4697 -65637
rect 4921 -66013 4955 -65637
rect 5179 -66013 5213 -65637
rect 5437 -66013 5471 -65637
rect 5695 -66013 5729 -65637
rect 5953 -66013 5987 -65637
rect 6211 -66013 6245 -65637
rect 4663 -66873 4697 -66497
rect 4921 -66873 4955 -66497
rect 5179 -66873 5213 -66497
rect 5437 -66873 5471 -66497
rect 5695 -66873 5729 -66497
rect 5953 -66873 5987 -66497
rect 6211 -66873 6245 -66497
rect -27996 -72719 -27962 -72685
rect -27996 -72787 -27962 -72753
rect -27996 -72855 -27962 -72821
rect -27912 -72719 -27878 -72685
rect -27912 -72787 -27878 -72753
rect -27912 -72855 -27878 -72821
rect -27337 -73699 -27303 -73323
rect -27079 -73699 -27045 -73323
rect -26821 -73699 -26787 -73323
rect -26563 -73699 -26529 -73323
rect -26305 -73699 -26271 -73323
rect -26047 -73699 -26013 -73323
rect -25789 -73699 -25755 -73323
rect -27337 -74559 -27303 -74183
rect -27079 -74559 -27045 -74183
rect -26821 -74559 -26787 -74183
rect -26563 -74559 -26529 -74183
rect -26305 -74559 -26271 -74183
rect -26047 -74559 -26013 -74183
rect -25789 -74559 -25755 -74183
rect -23996 -72719 -23962 -72685
rect -23996 -72787 -23962 -72753
rect -23996 -72855 -23962 -72821
rect -23912 -72719 -23878 -72685
rect -23912 -72787 -23878 -72753
rect -23912 -72855 -23878 -72821
rect -23337 -73699 -23303 -73323
rect -23079 -73699 -23045 -73323
rect -22821 -73699 -22787 -73323
rect -22563 -73699 -22529 -73323
rect -22305 -73699 -22271 -73323
rect -22047 -73699 -22013 -73323
rect -21789 -73699 -21755 -73323
rect -23337 -74559 -23303 -74183
rect -23079 -74559 -23045 -74183
rect -22821 -74559 -22787 -74183
rect -22563 -74559 -22529 -74183
rect -22305 -74559 -22271 -74183
rect -22047 -74559 -22013 -74183
rect -21789 -74559 -21755 -74183
rect -19996 -72719 -19962 -72685
rect -19996 -72787 -19962 -72753
rect -19996 -72855 -19962 -72821
rect -19912 -72719 -19878 -72685
rect -19912 -72787 -19878 -72753
rect -19912 -72855 -19878 -72821
rect -19337 -73699 -19303 -73323
rect -19079 -73699 -19045 -73323
rect -18821 -73699 -18787 -73323
rect -18563 -73699 -18529 -73323
rect -18305 -73699 -18271 -73323
rect -18047 -73699 -18013 -73323
rect -17789 -73699 -17755 -73323
rect -19337 -74559 -19303 -74183
rect -19079 -74559 -19045 -74183
rect -18821 -74559 -18787 -74183
rect -18563 -74559 -18529 -74183
rect -18305 -74559 -18271 -74183
rect -18047 -74559 -18013 -74183
rect -17789 -74559 -17755 -74183
rect -15996 -72719 -15962 -72685
rect -15996 -72787 -15962 -72753
rect -15996 -72855 -15962 -72821
rect -15912 -72719 -15878 -72685
rect -15912 -72787 -15878 -72753
rect -15912 -72855 -15878 -72821
rect -15337 -73699 -15303 -73323
rect -15079 -73699 -15045 -73323
rect -14821 -73699 -14787 -73323
rect -14563 -73699 -14529 -73323
rect -14305 -73699 -14271 -73323
rect -14047 -73699 -14013 -73323
rect -13789 -73699 -13755 -73323
rect -15337 -74559 -15303 -74183
rect -15079 -74559 -15045 -74183
rect -14821 -74559 -14787 -74183
rect -14563 -74559 -14529 -74183
rect -14305 -74559 -14271 -74183
rect -14047 -74559 -14013 -74183
rect -13789 -74559 -13755 -74183
rect -11996 -72719 -11962 -72685
rect -11996 -72787 -11962 -72753
rect -11996 -72855 -11962 -72821
rect -11912 -72719 -11878 -72685
rect -11912 -72787 -11878 -72753
rect -11912 -72855 -11878 -72821
rect -11337 -73699 -11303 -73323
rect -11079 -73699 -11045 -73323
rect -10821 -73699 -10787 -73323
rect -10563 -73699 -10529 -73323
rect -10305 -73699 -10271 -73323
rect -10047 -73699 -10013 -73323
rect -9789 -73699 -9755 -73323
rect -11337 -74559 -11303 -74183
rect -11079 -74559 -11045 -74183
rect -10821 -74559 -10787 -74183
rect -10563 -74559 -10529 -74183
rect -10305 -74559 -10271 -74183
rect -10047 -74559 -10013 -74183
rect -9789 -74559 -9755 -74183
rect -7996 -72719 -7962 -72685
rect -7996 -72787 -7962 -72753
rect -7996 -72855 -7962 -72821
rect -7912 -72719 -7878 -72685
rect -7912 -72787 -7878 -72753
rect -7912 -72855 -7878 -72821
rect -7337 -73699 -7303 -73323
rect -7079 -73699 -7045 -73323
rect -6821 -73699 -6787 -73323
rect -6563 -73699 -6529 -73323
rect -6305 -73699 -6271 -73323
rect -6047 -73699 -6013 -73323
rect -5789 -73699 -5755 -73323
rect -7337 -74559 -7303 -74183
rect -7079 -74559 -7045 -74183
rect -6821 -74559 -6787 -74183
rect -6563 -74559 -6529 -74183
rect -6305 -74559 -6271 -74183
rect -6047 -74559 -6013 -74183
rect -5789 -74559 -5755 -74183
rect -3996 -72719 -3962 -72685
rect -3996 -72787 -3962 -72753
rect -3996 -72855 -3962 -72821
rect -3912 -72719 -3878 -72685
rect -3912 -72787 -3878 -72753
rect -3912 -72855 -3878 -72821
rect -3337 -73699 -3303 -73323
rect -3079 -73699 -3045 -73323
rect -2821 -73699 -2787 -73323
rect -2563 -73699 -2529 -73323
rect -2305 -73699 -2271 -73323
rect -2047 -73699 -2013 -73323
rect -1789 -73699 -1755 -73323
rect -3337 -74559 -3303 -74183
rect -3079 -74559 -3045 -74183
rect -2821 -74559 -2787 -74183
rect -2563 -74559 -2529 -74183
rect -2305 -74559 -2271 -74183
rect -2047 -74559 -2013 -74183
rect -1789 -74559 -1755 -74183
rect 4 -72719 38 -72685
rect 4 -72787 38 -72753
rect 4 -72855 38 -72821
rect 88 -72719 122 -72685
rect 88 -72787 122 -72753
rect 88 -72855 122 -72821
rect 663 -73699 697 -73323
rect 921 -73699 955 -73323
rect 1179 -73699 1213 -73323
rect 1437 -73699 1471 -73323
rect 1695 -73699 1729 -73323
rect 1953 -73699 1987 -73323
rect 2211 -73699 2245 -73323
rect 663 -74559 697 -74183
rect 921 -74559 955 -74183
rect 1179 -74559 1213 -74183
rect 1437 -74559 1471 -74183
rect 1695 -74559 1729 -74183
rect 1953 -74559 1987 -74183
rect 2211 -74559 2245 -74183
rect 4004 -72719 4038 -72685
rect 4004 -72787 4038 -72753
rect 4004 -72855 4038 -72821
rect 4088 -72719 4122 -72685
rect 4088 -72787 4122 -72753
rect 4088 -72855 4122 -72821
rect 4663 -73699 4697 -73323
rect 4921 -73699 4955 -73323
rect 5179 -73699 5213 -73323
rect 5437 -73699 5471 -73323
rect 5695 -73699 5729 -73323
rect 5953 -73699 5987 -73323
rect 6211 -73699 6245 -73323
rect 4663 -74559 4697 -74183
rect 4921 -74559 4955 -74183
rect 5179 -74559 5213 -74183
rect 5437 -74559 5471 -74183
rect 5695 -74559 5729 -74183
rect 5953 -74559 5987 -74183
rect 6211 -74559 6245 -74183
<< psubdiff >>
rect 56370 -42446 56532 -42346
rect 57516 -42446 57728 -42346
rect 56370 -42508 56470 -42446
rect 55902 -42562 55998 -42528
rect 56186 -42562 56282 -42528
rect 55902 -42624 55936 -42562
rect 56248 -42624 56282 -42562
rect 55902 -42980 55936 -42918
rect 56248 -42980 56282 -42918
rect 55902 -43014 55998 -42980
rect 56186 -43014 56282 -42980
rect 57628 -42510 57728 -42446
rect 13122 -43256 13284 -43156
rect 50204 -43256 50366 -43156
rect 13122 -43318 13222 -43256
rect 10296 -57706 10392 -57672
rect 12010 -57706 12106 -57672
rect 10296 -57768 10330 -57706
rect 12072 -57768 12106 -57706
rect 10296 -58186 10330 -58124
rect 12072 -58186 12106 -58124
rect 10296 -58220 10392 -58186
rect 12010 -58220 12106 -58186
rect 50266 -43318 50366 -43256
rect 28530 -43762 28612 -43738
rect 28530 -43796 28554 -43762
rect 28588 -43796 28612 -43762
rect 28530 -43820 28612 -43796
rect 29548 -43762 29630 -43738
rect 29548 -43796 29572 -43762
rect 29606 -43796 29630 -43762
rect 29548 -43820 29630 -43796
rect 30566 -43762 30648 -43738
rect 30566 -43796 30590 -43762
rect 30624 -43796 30648 -43762
rect 30566 -43820 30648 -43796
rect 31584 -43762 31666 -43738
rect 31584 -43796 31608 -43762
rect 31642 -43796 31666 -43762
rect 31584 -43820 31666 -43796
rect 32602 -43762 32684 -43738
rect 32602 -43796 32626 -43762
rect 32660 -43796 32684 -43762
rect 32602 -43820 32684 -43796
rect 33620 -43762 33702 -43738
rect 33620 -43796 33644 -43762
rect 33678 -43796 33702 -43762
rect 33620 -43820 33702 -43796
rect 34638 -43762 34720 -43738
rect 34638 -43796 34662 -43762
rect 34696 -43796 34720 -43762
rect 34638 -43820 34720 -43796
rect 35656 -43762 35738 -43738
rect 35656 -43796 35680 -43762
rect 35714 -43796 35738 -43762
rect 35656 -43820 35738 -43796
rect 36674 -43762 36756 -43738
rect 36674 -43796 36698 -43762
rect 36732 -43796 36756 -43762
rect 36674 -43820 36756 -43796
rect 37692 -43762 37774 -43738
rect 37692 -43796 37716 -43762
rect 37750 -43796 37774 -43762
rect 37692 -43820 37774 -43796
rect 38710 -43762 38792 -43738
rect 38710 -43796 38734 -43762
rect 38768 -43796 38792 -43762
rect 38710 -43820 38792 -43796
rect 39728 -43762 39810 -43738
rect 39728 -43796 39752 -43762
rect 39786 -43796 39810 -43762
rect 39728 -43820 39810 -43796
rect 40746 -43762 40828 -43738
rect 40746 -43796 40770 -43762
rect 40804 -43796 40828 -43762
rect 40746 -43820 40828 -43796
rect 41764 -43762 41846 -43738
rect 41764 -43796 41788 -43762
rect 41822 -43796 41846 -43762
rect 41764 -43820 41846 -43796
rect 42782 -43762 42864 -43738
rect 42782 -43796 42806 -43762
rect 42840 -43796 42864 -43762
rect 42782 -43820 42864 -43796
rect 43800 -43762 43882 -43738
rect 43800 -43796 43824 -43762
rect 43858 -43796 43882 -43762
rect 43800 -43820 43882 -43796
rect 44818 -43762 44900 -43738
rect 44818 -43796 44842 -43762
rect 44876 -43796 44900 -43762
rect 44818 -43820 44900 -43796
rect 45836 -43762 45918 -43738
rect 45836 -43796 45860 -43762
rect 45894 -43796 45918 -43762
rect 45836 -43820 45918 -43796
rect 46854 -43762 46936 -43738
rect 46854 -43796 46878 -43762
rect 46912 -43796 46936 -43762
rect 46854 -43820 46936 -43796
rect 47872 -43762 47954 -43738
rect 47872 -43796 47896 -43762
rect 47930 -43796 47954 -43762
rect 47872 -43820 47954 -43796
rect 16236 -44364 16318 -44340
rect 16236 -44398 16260 -44364
rect 16294 -44398 16318 -44364
rect 16236 -44422 16318 -44398
rect 17254 -44364 17336 -44340
rect 17254 -44398 17278 -44364
rect 17312 -44398 17336 -44364
rect 17254 -44422 17336 -44398
rect 18272 -44364 18354 -44340
rect 18272 -44398 18296 -44364
rect 18330 -44398 18354 -44364
rect 18272 -44422 18354 -44398
rect 19290 -44364 19372 -44340
rect 19290 -44398 19314 -44364
rect 19348 -44398 19372 -44364
rect 19290 -44422 19372 -44398
rect 20308 -44364 20390 -44340
rect 20308 -44398 20332 -44364
rect 20366 -44398 20390 -44364
rect 20308 -44422 20390 -44398
rect 21326 -44364 21408 -44340
rect 21326 -44398 21350 -44364
rect 21384 -44398 21408 -44364
rect 21326 -44422 21408 -44398
rect 22344 -44364 22426 -44340
rect 22344 -44398 22368 -44364
rect 22402 -44398 22426 -44364
rect 22344 -44422 22426 -44398
rect 23362 -44364 23444 -44340
rect 23362 -44398 23386 -44364
rect 23420 -44398 23444 -44364
rect 23362 -44422 23444 -44398
rect 24380 -44364 24462 -44340
rect 24380 -44398 24404 -44364
rect 24438 -44398 24462 -44364
rect 24380 -44422 24462 -44398
rect 25408 -44364 25490 -44340
rect 25408 -44398 25432 -44364
rect 25466 -44398 25490 -44364
rect 25408 -44422 25490 -44398
rect 16236 -45182 16318 -45158
rect 16236 -45216 16260 -45182
rect 16294 -45216 16318 -45182
rect 16236 -45240 16318 -45216
rect 17254 -45182 17336 -45158
rect 17254 -45216 17278 -45182
rect 17312 -45216 17336 -45182
rect 17254 -45240 17336 -45216
rect 18272 -45182 18354 -45158
rect 18272 -45216 18296 -45182
rect 18330 -45216 18354 -45182
rect 18272 -45240 18354 -45216
rect 19290 -45182 19372 -45158
rect 19290 -45216 19314 -45182
rect 19348 -45216 19372 -45182
rect 19290 -45240 19372 -45216
rect 20308 -45182 20390 -45158
rect 20308 -45216 20332 -45182
rect 20366 -45216 20390 -45182
rect 20308 -45240 20390 -45216
rect 21326 -45182 21408 -45158
rect 21326 -45216 21350 -45182
rect 21384 -45216 21408 -45182
rect 21326 -45240 21408 -45216
rect 22344 -45182 22426 -45158
rect 22344 -45216 22368 -45182
rect 22402 -45216 22426 -45182
rect 22344 -45240 22426 -45216
rect 23362 -45182 23444 -45158
rect 23362 -45216 23386 -45182
rect 23420 -45216 23444 -45182
rect 23362 -45240 23444 -45216
rect 24380 -45182 24462 -45158
rect 24380 -45216 24404 -45182
rect 24438 -45216 24462 -45182
rect 24380 -45240 24462 -45216
rect 25408 -45182 25490 -45158
rect 25408 -45216 25432 -45182
rect 25466 -45216 25490 -45182
rect 25408 -45240 25490 -45216
rect 28542 -45788 28624 -45764
rect 28542 -45822 28566 -45788
rect 28600 -45822 28624 -45788
rect 28542 -45846 28624 -45822
rect 29560 -45788 29642 -45764
rect 29560 -45822 29584 -45788
rect 29618 -45822 29642 -45788
rect 29560 -45846 29642 -45822
rect 30578 -45788 30660 -45764
rect 30578 -45822 30602 -45788
rect 30636 -45822 30660 -45788
rect 30578 -45846 30660 -45822
rect 31596 -45788 31678 -45764
rect 31596 -45822 31620 -45788
rect 31654 -45822 31678 -45788
rect 31596 -45846 31678 -45822
rect 32614 -45788 32696 -45764
rect 32614 -45822 32638 -45788
rect 32672 -45822 32696 -45788
rect 32614 -45846 32696 -45822
rect 33632 -45788 33714 -45764
rect 33632 -45822 33656 -45788
rect 33690 -45822 33714 -45788
rect 33632 -45846 33714 -45822
rect 34650 -45788 34732 -45764
rect 34650 -45822 34674 -45788
rect 34708 -45822 34732 -45788
rect 34650 -45846 34732 -45822
rect 35668 -45788 35750 -45764
rect 35668 -45822 35692 -45788
rect 35726 -45822 35750 -45788
rect 35668 -45846 35750 -45822
rect 36686 -45788 36768 -45764
rect 36686 -45822 36710 -45788
rect 36744 -45822 36768 -45788
rect 36686 -45846 36768 -45822
rect 37704 -45788 37786 -45764
rect 37704 -45822 37728 -45788
rect 37762 -45822 37786 -45788
rect 37704 -45846 37786 -45822
rect 38722 -45788 38804 -45764
rect 38722 -45822 38746 -45788
rect 38780 -45822 38804 -45788
rect 38722 -45846 38804 -45822
rect 39740 -45788 39822 -45764
rect 39740 -45822 39764 -45788
rect 39798 -45822 39822 -45788
rect 39740 -45846 39822 -45822
rect 40758 -45788 40840 -45764
rect 40758 -45822 40782 -45788
rect 40816 -45822 40840 -45788
rect 40758 -45846 40840 -45822
rect 41776 -45788 41858 -45764
rect 41776 -45822 41800 -45788
rect 41834 -45822 41858 -45788
rect 41776 -45846 41858 -45822
rect 42794 -45788 42876 -45764
rect 42794 -45822 42818 -45788
rect 42852 -45822 42876 -45788
rect 42794 -45846 42876 -45822
rect 43812 -45788 43894 -45764
rect 43812 -45822 43836 -45788
rect 43870 -45822 43894 -45788
rect 43812 -45846 43894 -45822
rect 44830 -45788 44912 -45764
rect 44830 -45822 44854 -45788
rect 44888 -45822 44912 -45788
rect 44830 -45846 44912 -45822
rect 45848 -45788 45930 -45764
rect 45848 -45822 45872 -45788
rect 45906 -45822 45930 -45788
rect 45848 -45846 45930 -45822
rect 46866 -45788 46948 -45764
rect 46866 -45822 46890 -45788
rect 46924 -45822 46948 -45788
rect 46866 -45846 46948 -45822
rect 47884 -45788 47966 -45764
rect 47884 -45822 47908 -45788
rect 47942 -45822 47966 -45788
rect 47884 -45846 47966 -45822
rect 16236 -46000 16318 -45976
rect 16236 -46034 16260 -46000
rect 16294 -46034 16318 -46000
rect 16236 -46058 16318 -46034
rect 17254 -46000 17336 -45976
rect 17254 -46034 17278 -46000
rect 17312 -46034 17336 -46000
rect 17254 -46058 17336 -46034
rect 18272 -46000 18354 -45976
rect 18272 -46034 18296 -46000
rect 18330 -46034 18354 -46000
rect 18272 -46058 18354 -46034
rect 19290 -46000 19372 -45976
rect 19290 -46034 19314 -46000
rect 19348 -46034 19372 -46000
rect 19290 -46058 19372 -46034
rect 20308 -46000 20390 -45976
rect 20308 -46034 20332 -46000
rect 20366 -46034 20390 -46000
rect 20308 -46058 20390 -46034
rect 21326 -46000 21408 -45976
rect 21326 -46034 21350 -46000
rect 21384 -46034 21408 -46000
rect 21326 -46058 21408 -46034
rect 22344 -46000 22426 -45976
rect 22344 -46034 22368 -46000
rect 22402 -46034 22426 -46000
rect 22344 -46058 22426 -46034
rect 23362 -46000 23444 -45976
rect 23362 -46034 23386 -46000
rect 23420 -46034 23444 -46000
rect 23362 -46058 23444 -46034
rect 24380 -46000 24462 -45976
rect 24380 -46034 24404 -46000
rect 24438 -46034 24462 -46000
rect 24380 -46058 24462 -46034
rect 25408 -46000 25490 -45976
rect 25408 -46034 25432 -46000
rect 25466 -46034 25490 -46000
rect 25408 -46058 25490 -46034
rect 16236 -46818 16318 -46794
rect 16236 -46852 16260 -46818
rect 16294 -46852 16318 -46818
rect 16236 -46876 16318 -46852
rect 17254 -46818 17336 -46794
rect 17254 -46852 17278 -46818
rect 17312 -46852 17336 -46818
rect 17254 -46876 17336 -46852
rect 18272 -46818 18354 -46794
rect 18272 -46852 18296 -46818
rect 18330 -46852 18354 -46818
rect 18272 -46876 18354 -46852
rect 19290 -46818 19372 -46794
rect 19290 -46852 19314 -46818
rect 19348 -46852 19372 -46818
rect 19290 -46876 19372 -46852
rect 20308 -46818 20390 -46794
rect 20308 -46852 20332 -46818
rect 20366 -46852 20390 -46818
rect 20308 -46876 20390 -46852
rect 21326 -46818 21408 -46794
rect 21326 -46852 21350 -46818
rect 21384 -46852 21408 -46818
rect 21326 -46876 21408 -46852
rect 22344 -46818 22426 -46794
rect 22344 -46852 22368 -46818
rect 22402 -46852 22426 -46818
rect 22344 -46876 22426 -46852
rect 23362 -46818 23444 -46794
rect 23362 -46852 23386 -46818
rect 23420 -46852 23444 -46818
rect 23362 -46876 23444 -46852
rect 24380 -46818 24462 -46794
rect 24380 -46852 24404 -46818
rect 24438 -46852 24462 -46818
rect 24380 -46876 24462 -46852
rect 25408 -46818 25490 -46794
rect 25408 -46852 25432 -46818
rect 25466 -46852 25490 -46818
rect 25408 -46876 25490 -46852
rect 28530 -47094 28612 -47070
rect 28530 -47128 28554 -47094
rect 28588 -47128 28612 -47094
rect 28530 -47152 28612 -47128
rect 29548 -47094 29630 -47070
rect 29548 -47128 29572 -47094
rect 29606 -47128 29630 -47094
rect 29548 -47152 29630 -47128
rect 30566 -47094 30648 -47070
rect 30566 -47128 30590 -47094
rect 30624 -47128 30648 -47094
rect 30566 -47152 30648 -47128
rect 31584 -47094 31666 -47070
rect 31584 -47128 31608 -47094
rect 31642 -47128 31666 -47094
rect 31584 -47152 31666 -47128
rect 32602 -47094 32684 -47070
rect 32602 -47128 32626 -47094
rect 32660 -47128 32684 -47094
rect 32602 -47152 32684 -47128
rect 33620 -47094 33702 -47070
rect 33620 -47128 33644 -47094
rect 33678 -47128 33702 -47094
rect 33620 -47152 33702 -47128
rect 34638 -47094 34720 -47070
rect 34638 -47128 34662 -47094
rect 34696 -47128 34720 -47094
rect 34638 -47152 34720 -47128
rect 35656 -47094 35738 -47070
rect 35656 -47128 35680 -47094
rect 35714 -47128 35738 -47094
rect 35656 -47152 35738 -47128
rect 36674 -47094 36756 -47070
rect 36674 -47128 36698 -47094
rect 36732 -47128 36756 -47094
rect 36674 -47152 36756 -47128
rect 37692 -47094 37774 -47070
rect 37692 -47128 37716 -47094
rect 37750 -47128 37774 -47094
rect 37692 -47152 37774 -47128
rect 38710 -47094 38792 -47070
rect 38710 -47128 38734 -47094
rect 38768 -47128 38792 -47094
rect 38710 -47152 38792 -47128
rect 39728 -47094 39810 -47070
rect 39728 -47128 39752 -47094
rect 39786 -47128 39810 -47094
rect 39728 -47152 39810 -47128
rect 40746 -47094 40828 -47070
rect 40746 -47128 40770 -47094
rect 40804 -47128 40828 -47094
rect 40746 -47152 40828 -47128
rect 41764 -47094 41846 -47070
rect 41764 -47128 41788 -47094
rect 41822 -47128 41846 -47094
rect 41764 -47152 41846 -47128
rect 42782 -47094 42864 -47070
rect 42782 -47128 42806 -47094
rect 42840 -47128 42864 -47094
rect 42782 -47152 42864 -47128
rect 43800 -47094 43882 -47070
rect 43800 -47128 43824 -47094
rect 43858 -47128 43882 -47094
rect 43800 -47152 43882 -47128
rect 44818 -47094 44900 -47070
rect 44818 -47128 44842 -47094
rect 44876 -47128 44900 -47094
rect 44818 -47152 44900 -47128
rect 45836 -47094 45918 -47070
rect 45836 -47128 45860 -47094
rect 45894 -47128 45918 -47094
rect 45836 -47152 45918 -47128
rect 46854 -47094 46936 -47070
rect 46854 -47128 46878 -47094
rect 46912 -47128 46936 -47094
rect 46854 -47152 46936 -47128
rect 47872 -47094 47954 -47070
rect 47872 -47128 47896 -47094
rect 47930 -47128 47954 -47094
rect 47872 -47152 47954 -47128
rect 16236 -47636 16318 -47612
rect 16236 -47670 16260 -47636
rect 16294 -47670 16318 -47636
rect 16236 -47694 16318 -47670
rect 17254 -47636 17336 -47612
rect 17254 -47670 17278 -47636
rect 17312 -47670 17336 -47636
rect 17254 -47694 17336 -47670
rect 18272 -47636 18354 -47612
rect 18272 -47670 18296 -47636
rect 18330 -47670 18354 -47636
rect 18272 -47694 18354 -47670
rect 19290 -47636 19372 -47612
rect 19290 -47670 19314 -47636
rect 19348 -47670 19372 -47636
rect 19290 -47694 19372 -47670
rect 20308 -47636 20390 -47612
rect 20308 -47670 20332 -47636
rect 20366 -47670 20390 -47636
rect 20308 -47694 20390 -47670
rect 21326 -47636 21408 -47612
rect 21326 -47670 21350 -47636
rect 21384 -47670 21408 -47636
rect 21326 -47694 21408 -47670
rect 22344 -47636 22426 -47612
rect 22344 -47670 22368 -47636
rect 22402 -47670 22426 -47636
rect 22344 -47694 22426 -47670
rect 23362 -47636 23444 -47612
rect 23362 -47670 23386 -47636
rect 23420 -47670 23444 -47636
rect 23362 -47694 23444 -47670
rect 24380 -47636 24462 -47612
rect 24380 -47670 24404 -47636
rect 24438 -47670 24462 -47636
rect 24380 -47694 24462 -47670
rect 25408 -47636 25490 -47612
rect 25408 -47670 25432 -47636
rect 25466 -47670 25490 -47636
rect 25408 -47694 25490 -47670
rect 28518 -48330 28600 -48306
rect 16236 -48454 16318 -48430
rect 16236 -48488 16260 -48454
rect 16294 -48488 16318 -48454
rect 16236 -48512 16318 -48488
rect 17254 -48454 17336 -48430
rect 17254 -48488 17278 -48454
rect 17312 -48488 17336 -48454
rect 17254 -48512 17336 -48488
rect 18272 -48454 18354 -48430
rect 18272 -48488 18296 -48454
rect 18330 -48488 18354 -48454
rect 18272 -48512 18354 -48488
rect 19290 -48454 19372 -48430
rect 19290 -48488 19314 -48454
rect 19348 -48488 19372 -48454
rect 19290 -48512 19372 -48488
rect 20308 -48454 20390 -48430
rect 20308 -48488 20332 -48454
rect 20366 -48488 20390 -48454
rect 20308 -48512 20390 -48488
rect 21326 -48454 21408 -48430
rect 21326 -48488 21350 -48454
rect 21384 -48488 21408 -48454
rect 21326 -48512 21408 -48488
rect 22344 -48454 22426 -48430
rect 22344 -48488 22368 -48454
rect 22402 -48488 22426 -48454
rect 22344 -48512 22426 -48488
rect 23362 -48454 23444 -48430
rect 28518 -48364 28542 -48330
rect 28576 -48364 28600 -48330
rect 28518 -48388 28600 -48364
rect 29536 -48330 29618 -48306
rect 29536 -48364 29560 -48330
rect 29594 -48364 29618 -48330
rect 29536 -48388 29618 -48364
rect 30554 -48330 30636 -48306
rect 30554 -48364 30578 -48330
rect 30612 -48364 30636 -48330
rect 30554 -48388 30636 -48364
rect 31572 -48330 31654 -48306
rect 31572 -48364 31596 -48330
rect 31630 -48364 31654 -48330
rect 31572 -48388 31654 -48364
rect 32590 -48330 32672 -48306
rect 32590 -48364 32614 -48330
rect 32648 -48364 32672 -48330
rect 32590 -48388 32672 -48364
rect 33608 -48330 33690 -48306
rect 33608 -48364 33632 -48330
rect 33666 -48364 33690 -48330
rect 33608 -48388 33690 -48364
rect 34626 -48330 34708 -48306
rect 34626 -48364 34650 -48330
rect 34684 -48364 34708 -48330
rect 34626 -48388 34708 -48364
rect 35644 -48330 35726 -48306
rect 35644 -48364 35668 -48330
rect 35702 -48364 35726 -48330
rect 35644 -48388 35726 -48364
rect 36662 -48330 36744 -48306
rect 36662 -48364 36686 -48330
rect 36720 -48364 36744 -48330
rect 36662 -48388 36744 -48364
rect 37680 -48330 37762 -48306
rect 37680 -48364 37704 -48330
rect 37738 -48364 37762 -48330
rect 37680 -48388 37762 -48364
rect 38698 -48330 38780 -48306
rect 38698 -48364 38722 -48330
rect 38756 -48364 38780 -48330
rect 38698 -48388 38780 -48364
rect 39716 -48330 39798 -48306
rect 39716 -48364 39740 -48330
rect 39774 -48364 39798 -48330
rect 39716 -48388 39798 -48364
rect 40734 -48330 40816 -48306
rect 40734 -48364 40758 -48330
rect 40792 -48364 40816 -48330
rect 40734 -48388 40816 -48364
rect 41752 -48330 41834 -48306
rect 41752 -48364 41776 -48330
rect 41810 -48364 41834 -48330
rect 41752 -48388 41834 -48364
rect 42770 -48330 42852 -48306
rect 42770 -48364 42794 -48330
rect 42828 -48364 42852 -48330
rect 42770 -48388 42852 -48364
rect 43788 -48330 43870 -48306
rect 43788 -48364 43812 -48330
rect 43846 -48364 43870 -48330
rect 43788 -48388 43870 -48364
rect 44806 -48330 44888 -48306
rect 44806 -48364 44830 -48330
rect 44864 -48364 44888 -48330
rect 44806 -48388 44888 -48364
rect 45824 -48330 45906 -48306
rect 45824 -48364 45848 -48330
rect 45882 -48364 45906 -48330
rect 45824 -48388 45906 -48364
rect 46842 -48330 46924 -48306
rect 46842 -48364 46866 -48330
rect 46900 -48364 46924 -48330
rect 46842 -48388 46924 -48364
rect 47860 -48330 47942 -48306
rect 47860 -48364 47884 -48330
rect 47918 -48364 47942 -48330
rect 47860 -48388 47942 -48364
rect 23362 -48488 23386 -48454
rect 23420 -48488 23444 -48454
rect 23362 -48512 23444 -48488
rect 24380 -48454 24462 -48430
rect 24380 -48488 24404 -48454
rect 24438 -48488 24462 -48454
rect 24380 -48512 24462 -48488
rect 25408 -48454 25490 -48430
rect 25408 -48488 25432 -48454
rect 25466 -48488 25490 -48454
rect 25408 -48512 25490 -48488
rect 16236 -49272 16318 -49248
rect 16236 -49306 16260 -49272
rect 16294 -49306 16318 -49272
rect 16236 -49330 16318 -49306
rect 17254 -49272 17336 -49248
rect 17254 -49306 17278 -49272
rect 17312 -49306 17336 -49272
rect 17254 -49330 17336 -49306
rect 18272 -49272 18354 -49248
rect 18272 -49306 18296 -49272
rect 18330 -49306 18354 -49272
rect 18272 -49330 18354 -49306
rect 19290 -49272 19372 -49248
rect 19290 -49306 19314 -49272
rect 19348 -49306 19372 -49272
rect 19290 -49330 19372 -49306
rect 20308 -49272 20390 -49248
rect 20308 -49306 20332 -49272
rect 20366 -49306 20390 -49272
rect 20308 -49330 20390 -49306
rect 21326 -49272 21408 -49248
rect 21326 -49306 21350 -49272
rect 21384 -49306 21408 -49272
rect 21326 -49330 21408 -49306
rect 22344 -49272 22426 -49248
rect 22344 -49306 22368 -49272
rect 22402 -49306 22426 -49272
rect 22344 -49330 22426 -49306
rect 23362 -49272 23444 -49248
rect 23362 -49306 23386 -49272
rect 23420 -49306 23444 -49272
rect 23362 -49330 23444 -49306
rect 24380 -49272 24462 -49248
rect 24380 -49306 24404 -49272
rect 24438 -49306 24462 -49272
rect 24380 -49330 24462 -49306
rect 25408 -49272 25490 -49248
rect 25408 -49306 25432 -49272
rect 25466 -49306 25490 -49272
rect 25408 -49330 25490 -49306
rect 28518 -49554 28600 -49530
rect 28518 -49588 28542 -49554
rect 28576 -49588 28600 -49554
rect 28518 -49612 28600 -49588
rect 29536 -49554 29618 -49530
rect 29536 -49588 29560 -49554
rect 29594 -49588 29618 -49554
rect 29536 -49612 29618 -49588
rect 30554 -49554 30636 -49530
rect 30554 -49588 30578 -49554
rect 30612 -49588 30636 -49554
rect 30554 -49612 30636 -49588
rect 31572 -49554 31654 -49530
rect 31572 -49588 31596 -49554
rect 31630 -49588 31654 -49554
rect 31572 -49612 31654 -49588
rect 32590 -49554 32672 -49530
rect 32590 -49588 32614 -49554
rect 32648 -49588 32672 -49554
rect 32590 -49612 32672 -49588
rect 33608 -49554 33690 -49530
rect 33608 -49588 33632 -49554
rect 33666 -49588 33690 -49554
rect 33608 -49612 33690 -49588
rect 34626 -49554 34708 -49530
rect 34626 -49588 34650 -49554
rect 34684 -49588 34708 -49554
rect 34626 -49612 34708 -49588
rect 35644 -49554 35726 -49530
rect 35644 -49588 35668 -49554
rect 35702 -49588 35726 -49554
rect 35644 -49612 35726 -49588
rect 36662 -49554 36744 -49530
rect 36662 -49588 36686 -49554
rect 36720 -49588 36744 -49554
rect 36662 -49612 36744 -49588
rect 37680 -49554 37762 -49530
rect 37680 -49588 37704 -49554
rect 37738 -49588 37762 -49554
rect 37680 -49612 37762 -49588
rect 38698 -49554 38780 -49530
rect 38698 -49588 38722 -49554
rect 38756 -49588 38780 -49554
rect 38698 -49612 38780 -49588
rect 39716 -49554 39798 -49530
rect 39716 -49588 39740 -49554
rect 39774 -49588 39798 -49554
rect 39716 -49612 39798 -49588
rect 40734 -49554 40816 -49530
rect 40734 -49588 40758 -49554
rect 40792 -49588 40816 -49554
rect 40734 -49612 40816 -49588
rect 41752 -49554 41834 -49530
rect 41752 -49588 41776 -49554
rect 41810 -49588 41834 -49554
rect 41752 -49612 41834 -49588
rect 42770 -49554 42852 -49530
rect 42770 -49588 42794 -49554
rect 42828 -49588 42852 -49554
rect 42770 -49612 42852 -49588
rect 43788 -49554 43870 -49530
rect 43788 -49588 43812 -49554
rect 43846 -49588 43870 -49554
rect 43788 -49612 43870 -49588
rect 44806 -49554 44888 -49530
rect 44806 -49588 44830 -49554
rect 44864 -49588 44888 -49554
rect 44806 -49612 44888 -49588
rect 45824 -49554 45906 -49530
rect 45824 -49588 45848 -49554
rect 45882 -49588 45906 -49554
rect 45824 -49612 45906 -49588
rect 46842 -49554 46924 -49530
rect 46842 -49588 46866 -49554
rect 46900 -49588 46924 -49554
rect 46842 -49612 46924 -49588
rect 47860 -49554 47942 -49530
rect 47860 -49588 47884 -49554
rect 47918 -49588 47942 -49554
rect 47860 -49612 47942 -49588
rect 16236 -50090 16318 -50066
rect 16236 -50124 16260 -50090
rect 16294 -50124 16318 -50090
rect 16236 -50148 16318 -50124
rect 17254 -50090 17336 -50066
rect 17254 -50124 17278 -50090
rect 17312 -50124 17336 -50090
rect 17254 -50148 17336 -50124
rect 18272 -50090 18354 -50066
rect 18272 -50124 18296 -50090
rect 18330 -50124 18354 -50090
rect 18272 -50148 18354 -50124
rect 19290 -50090 19372 -50066
rect 19290 -50124 19314 -50090
rect 19348 -50124 19372 -50090
rect 19290 -50148 19372 -50124
rect 20308 -50090 20390 -50066
rect 20308 -50124 20332 -50090
rect 20366 -50124 20390 -50090
rect 20308 -50148 20390 -50124
rect 21326 -50090 21408 -50066
rect 21326 -50124 21350 -50090
rect 21384 -50124 21408 -50090
rect 21326 -50148 21408 -50124
rect 22344 -50090 22426 -50066
rect 22344 -50124 22368 -50090
rect 22402 -50124 22426 -50090
rect 22344 -50148 22426 -50124
rect 23362 -50090 23444 -50066
rect 23362 -50124 23386 -50090
rect 23420 -50124 23444 -50090
rect 23362 -50148 23444 -50124
rect 24380 -50090 24462 -50066
rect 24380 -50124 24404 -50090
rect 24438 -50124 24462 -50090
rect 24380 -50148 24462 -50124
rect 25408 -50090 25490 -50066
rect 25408 -50124 25432 -50090
rect 25466 -50124 25490 -50090
rect 25408 -50148 25490 -50124
rect 28530 -50790 28612 -50766
rect 28530 -50824 28554 -50790
rect 28588 -50824 28612 -50790
rect 28530 -50848 28612 -50824
rect 29548 -50790 29630 -50766
rect 29548 -50824 29572 -50790
rect 29606 -50824 29630 -50790
rect 29548 -50848 29630 -50824
rect 30566 -50790 30648 -50766
rect 30566 -50824 30590 -50790
rect 30624 -50824 30648 -50790
rect 30566 -50848 30648 -50824
rect 31584 -50790 31666 -50766
rect 31584 -50824 31608 -50790
rect 31642 -50824 31666 -50790
rect 31584 -50848 31666 -50824
rect 32602 -50790 32684 -50766
rect 32602 -50824 32626 -50790
rect 32660 -50824 32684 -50790
rect 32602 -50848 32684 -50824
rect 33620 -50790 33702 -50766
rect 33620 -50824 33644 -50790
rect 33678 -50824 33702 -50790
rect 33620 -50848 33702 -50824
rect 34638 -50790 34720 -50766
rect 34638 -50824 34662 -50790
rect 34696 -50824 34720 -50790
rect 34638 -50848 34720 -50824
rect 35656 -50790 35738 -50766
rect 35656 -50824 35680 -50790
rect 35714 -50824 35738 -50790
rect 35656 -50848 35738 -50824
rect 36674 -50790 36756 -50766
rect 36674 -50824 36698 -50790
rect 36732 -50824 36756 -50790
rect 36674 -50848 36756 -50824
rect 37692 -50790 37774 -50766
rect 37692 -50824 37716 -50790
rect 37750 -50824 37774 -50790
rect 37692 -50848 37774 -50824
rect 38710 -50790 38792 -50766
rect 38710 -50824 38734 -50790
rect 38768 -50824 38792 -50790
rect 38710 -50848 38792 -50824
rect 39728 -50790 39810 -50766
rect 39728 -50824 39752 -50790
rect 39786 -50824 39810 -50790
rect 39728 -50848 39810 -50824
rect 40746 -50790 40828 -50766
rect 40746 -50824 40770 -50790
rect 40804 -50824 40828 -50790
rect 40746 -50848 40828 -50824
rect 41764 -50790 41846 -50766
rect 41764 -50824 41788 -50790
rect 41822 -50824 41846 -50790
rect 41764 -50848 41846 -50824
rect 42782 -50790 42864 -50766
rect 42782 -50824 42806 -50790
rect 42840 -50824 42864 -50790
rect 42782 -50848 42864 -50824
rect 43800 -50790 43882 -50766
rect 43800 -50824 43824 -50790
rect 43858 -50824 43882 -50790
rect 43800 -50848 43882 -50824
rect 44818 -50790 44900 -50766
rect 44818 -50824 44842 -50790
rect 44876 -50824 44900 -50790
rect 44818 -50848 44900 -50824
rect 45836 -50790 45918 -50766
rect 45836 -50824 45860 -50790
rect 45894 -50824 45918 -50790
rect 45836 -50848 45918 -50824
rect 46854 -50790 46936 -50766
rect 46854 -50824 46878 -50790
rect 46912 -50824 46936 -50790
rect 46854 -50848 46936 -50824
rect 47872 -50790 47954 -50766
rect 47872 -50824 47896 -50790
rect 47930 -50824 47954 -50790
rect 47872 -50848 47954 -50824
rect 16224 -50984 16306 -50960
rect 16224 -51018 16248 -50984
rect 16282 -51018 16306 -50984
rect 16224 -51042 16306 -51018
rect 17242 -50984 17324 -50960
rect 17242 -51018 17266 -50984
rect 17300 -51018 17324 -50984
rect 17242 -51042 17324 -51018
rect 18260 -50984 18342 -50960
rect 18260 -51018 18284 -50984
rect 18318 -51018 18342 -50984
rect 18260 -51042 18342 -51018
rect 19278 -50984 19360 -50960
rect 19278 -51018 19302 -50984
rect 19336 -51018 19360 -50984
rect 19278 -51042 19360 -51018
rect 20296 -50984 20378 -50960
rect 20296 -51018 20320 -50984
rect 20354 -51018 20378 -50984
rect 20296 -51042 20378 -51018
rect 21314 -50984 21396 -50960
rect 21314 -51018 21338 -50984
rect 21372 -51018 21396 -50984
rect 21314 -51042 21396 -51018
rect 22332 -50984 22414 -50960
rect 22332 -51018 22356 -50984
rect 22390 -51018 22414 -50984
rect 22332 -51042 22414 -51018
rect 23350 -50984 23432 -50960
rect 23350 -51018 23374 -50984
rect 23408 -51018 23432 -50984
rect 23350 -51042 23432 -51018
rect 24368 -50984 24450 -50960
rect 24368 -51018 24392 -50984
rect 24426 -51018 24450 -50984
rect 24368 -51042 24450 -51018
rect 25396 -50984 25478 -50960
rect 25396 -51018 25420 -50984
rect 25454 -51018 25478 -50984
rect 25396 -51042 25478 -51018
rect 15428 -51932 15510 -51908
rect 15428 -51966 15452 -51932
rect 15486 -51966 15510 -51932
rect 15428 -51990 15510 -51966
rect 16446 -51932 16528 -51908
rect 16446 -51966 16470 -51932
rect 16504 -51966 16528 -51932
rect 16446 -51990 16528 -51966
rect 17464 -51932 17546 -51908
rect 17464 -51966 17488 -51932
rect 17522 -51966 17546 -51932
rect 17464 -51990 17546 -51966
rect 18482 -51932 18564 -51908
rect 18482 -51966 18506 -51932
rect 18540 -51966 18564 -51932
rect 18482 -51990 18564 -51966
rect 19500 -51932 19582 -51908
rect 19500 -51966 19524 -51932
rect 19558 -51966 19582 -51932
rect 19500 -51990 19582 -51966
rect 20518 -51932 20600 -51908
rect 20518 -51966 20542 -51932
rect 20576 -51966 20600 -51932
rect 20518 -51990 20600 -51966
rect 21536 -51932 21618 -51908
rect 21536 -51966 21560 -51932
rect 21594 -51966 21618 -51932
rect 21536 -51990 21618 -51966
rect 22554 -51932 22636 -51908
rect 22554 -51966 22578 -51932
rect 22612 -51966 22636 -51932
rect 22554 -51990 22636 -51966
rect 23572 -51932 23654 -51908
rect 23572 -51966 23596 -51932
rect 23630 -51966 23654 -51932
rect 23572 -51990 23654 -51966
rect 24590 -51932 24672 -51908
rect 24590 -51966 24614 -51932
rect 24648 -51966 24672 -51932
rect 24590 -51990 24672 -51966
rect 25608 -51932 25690 -51908
rect 25608 -51966 25632 -51932
rect 25666 -51966 25690 -51932
rect 25608 -51990 25690 -51966
rect 28530 -52038 28612 -52014
rect 28530 -52072 28554 -52038
rect 28588 -52072 28612 -52038
rect 28530 -52096 28612 -52072
rect 29548 -52038 29630 -52014
rect 29548 -52072 29572 -52038
rect 29606 -52072 29630 -52038
rect 29548 -52096 29630 -52072
rect 30566 -52038 30648 -52014
rect 30566 -52072 30590 -52038
rect 30624 -52072 30648 -52038
rect 30566 -52096 30648 -52072
rect 31584 -52038 31666 -52014
rect 31584 -52072 31608 -52038
rect 31642 -52072 31666 -52038
rect 31584 -52096 31666 -52072
rect 32602 -52038 32684 -52014
rect 32602 -52072 32626 -52038
rect 32660 -52072 32684 -52038
rect 32602 -52096 32684 -52072
rect 33620 -52038 33702 -52014
rect 33620 -52072 33644 -52038
rect 33678 -52072 33702 -52038
rect 33620 -52096 33702 -52072
rect 34638 -52038 34720 -52014
rect 34638 -52072 34662 -52038
rect 34696 -52072 34720 -52038
rect 34638 -52096 34720 -52072
rect 35656 -52038 35738 -52014
rect 35656 -52072 35680 -52038
rect 35714 -52072 35738 -52038
rect 35656 -52096 35738 -52072
rect 36674 -52038 36756 -52014
rect 36674 -52072 36698 -52038
rect 36732 -52072 36756 -52038
rect 36674 -52096 36756 -52072
rect 37692 -52038 37774 -52014
rect 37692 -52072 37716 -52038
rect 37750 -52072 37774 -52038
rect 37692 -52096 37774 -52072
rect 38710 -52038 38792 -52014
rect 38710 -52072 38734 -52038
rect 38768 -52072 38792 -52038
rect 38710 -52096 38792 -52072
rect 39728 -52038 39810 -52014
rect 39728 -52072 39752 -52038
rect 39786 -52072 39810 -52038
rect 39728 -52096 39810 -52072
rect 40746 -52038 40828 -52014
rect 40746 -52072 40770 -52038
rect 40804 -52072 40828 -52038
rect 40746 -52096 40828 -52072
rect 41764 -52038 41846 -52014
rect 41764 -52072 41788 -52038
rect 41822 -52072 41846 -52038
rect 41764 -52096 41846 -52072
rect 42782 -52038 42864 -52014
rect 42782 -52072 42806 -52038
rect 42840 -52072 42864 -52038
rect 42782 -52096 42864 -52072
rect 43800 -52038 43882 -52014
rect 43800 -52072 43824 -52038
rect 43858 -52072 43882 -52038
rect 43800 -52096 43882 -52072
rect 44818 -52038 44900 -52014
rect 44818 -52072 44842 -52038
rect 44876 -52072 44900 -52038
rect 44818 -52096 44900 -52072
rect 45836 -52038 45918 -52014
rect 45836 -52072 45860 -52038
rect 45894 -52072 45918 -52038
rect 45836 -52096 45918 -52072
rect 46854 -52038 46936 -52014
rect 46854 -52072 46878 -52038
rect 46912 -52072 46936 -52038
rect 46854 -52096 46936 -52072
rect 47872 -52038 47954 -52014
rect 47872 -52072 47896 -52038
rect 47930 -52072 47954 -52038
rect 47872 -52096 47954 -52072
rect 15440 -53074 15522 -53050
rect 15440 -53108 15464 -53074
rect 15498 -53108 15522 -53074
rect 15440 -53132 15522 -53108
rect 16458 -53074 16540 -53050
rect 16458 -53108 16482 -53074
rect 16516 -53108 16540 -53074
rect 16458 -53132 16540 -53108
rect 17476 -53074 17558 -53050
rect 17476 -53108 17500 -53074
rect 17534 -53108 17558 -53074
rect 17476 -53132 17558 -53108
rect 18494 -53074 18576 -53050
rect 18494 -53108 18518 -53074
rect 18552 -53108 18576 -53074
rect 18494 -53132 18576 -53108
rect 19512 -53074 19594 -53050
rect 19512 -53108 19536 -53074
rect 19570 -53108 19594 -53074
rect 19512 -53132 19594 -53108
rect 20530 -53074 20612 -53050
rect 20530 -53108 20554 -53074
rect 20588 -53108 20612 -53074
rect 20530 -53132 20612 -53108
rect 21548 -53074 21630 -53050
rect 21548 -53108 21572 -53074
rect 21606 -53108 21630 -53074
rect 21548 -53132 21630 -53108
rect 22566 -53074 22648 -53050
rect 22566 -53108 22590 -53074
rect 22624 -53108 22648 -53074
rect 22566 -53132 22648 -53108
rect 23584 -53074 23666 -53050
rect 23584 -53108 23608 -53074
rect 23642 -53108 23666 -53074
rect 23584 -53132 23666 -53108
rect 24602 -53074 24684 -53050
rect 24602 -53108 24626 -53074
rect 24660 -53108 24684 -53074
rect 24602 -53132 24684 -53108
rect 25620 -53074 25702 -53050
rect 25620 -53108 25644 -53074
rect 25678 -53108 25702 -53074
rect 25620 -53132 25702 -53108
rect 28506 -53274 28588 -53250
rect 28506 -53308 28530 -53274
rect 28564 -53308 28588 -53274
rect 28506 -53332 28588 -53308
rect 29524 -53274 29606 -53250
rect 29524 -53308 29548 -53274
rect 29582 -53308 29606 -53274
rect 29524 -53332 29606 -53308
rect 30542 -53274 30624 -53250
rect 30542 -53308 30566 -53274
rect 30600 -53308 30624 -53274
rect 30542 -53332 30624 -53308
rect 31560 -53274 31642 -53250
rect 31560 -53308 31584 -53274
rect 31618 -53308 31642 -53274
rect 31560 -53332 31642 -53308
rect 32578 -53274 32660 -53250
rect 32578 -53308 32602 -53274
rect 32636 -53308 32660 -53274
rect 32578 -53332 32660 -53308
rect 33596 -53274 33678 -53250
rect 33596 -53308 33620 -53274
rect 33654 -53308 33678 -53274
rect 33596 -53332 33678 -53308
rect 34614 -53274 34696 -53250
rect 34614 -53308 34638 -53274
rect 34672 -53308 34696 -53274
rect 34614 -53332 34696 -53308
rect 35632 -53274 35714 -53250
rect 35632 -53308 35656 -53274
rect 35690 -53308 35714 -53274
rect 35632 -53332 35714 -53308
rect 36650 -53274 36732 -53250
rect 36650 -53308 36674 -53274
rect 36708 -53308 36732 -53274
rect 36650 -53332 36732 -53308
rect 37668 -53274 37750 -53250
rect 37668 -53308 37692 -53274
rect 37726 -53308 37750 -53274
rect 37668 -53332 37750 -53308
rect 38686 -53274 38768 -53250
rect 38686 -53308 38710 -53274
rect 38744 -53308 38768 -53274
rect 38686 -53332 38768 -53308
rect 39704 -53274 39786 -53250
rect 39704 -53308 39728 -53274
rect 39762 -53308 39786 -53274
rect 39704 -53332 39786 -53308
rect 40722 -53274 40804 -53250
rect 40722 -53308 40746 -53274
rect 40780 -53308 40804 -53274
rect 40722 -53332 40804 -53308
rect 41740 -53274 41822 -53250
rect 41740 -53308 41764 -53274
rect 41798 -53308 41822 -53274
rect 41740 -53332 41822 -53308
rect 42758 -53274 42840 -53250
rect 42758 -53308 42782 -53274
rect 42816 -53308 42840 -53274
rect 42758 -53332 42840 -53308
rect 43776 -53274 43858 -53250
rect 43776 -53308 43800 -53274
rect 43834 -53308 43858 -53274
rect 43776 -53332 43858 -53308
rect 44794 -53274 44876 -53250
rect 44794 -53308 44818 -53274
rect 44852 -53308 44876 -53274
rect 44794 -53332 44876 -53308
rect 45812 -53274 45894 -53250
rect 45812 -53308 45836 -53274
rect 45870 -53308 45894 -53274
rect 45812 -53332 45894 -53308
rect 46830 -53274 46912 -53250
rect 46830 -53308 46854 -53274
rect 46888 -53308 46912 -53274
rect 46830 -53332 46912 -53308
rect 47848 -53274 47930 -53250
rect 47848 -53308 47872 -53274
rect 47906 -53308 47930 -53274
rect 47848 -53332 47930 -53308
rect 15418 -54182 15500 -54158
rect 15418 -54216 15442 -54182
rect 15476 -54216 15500 -54182
rect 15418 -54240 15500 -54216
rect 16436 -54182 16518 -54158
rect 16436 -54216 16460 -54182
rect 16494 -54216 16518 -54182
rect 16436 -54240 16518 -54216
rect 17454 -54182 17536 -54158
rect 17454 -54216 17478 -54182
rect 17512 -54216 17536 -54182
rect 17454 -54240 17536 -54216
rect 18472 -54182 18554 -54158
rect 18472 -54216 18496 -54182
rect 18530 -54216 18554 -54182
rect 18472 -54240 18554 -54216
rect 19490 -54182 19572 -54158
rect 19490 -54216 19514 -54182
rect 19548 -54216 19572 -54182
rect 19490 -54240 19572 -54216
rect 20508 -54182 20590 -54158
rect 20508 -54216 20532 -54182
rect 20566 -54216 20590 -54182
rect 20508 -54240 20590 -54216
rect 21526 -54182 21608 -54158
rect 21526 -54216 21550 -54182
rect 21584 -54216 21608 -54182
rect 21526 -54240 21608 -54216
rect 22544 -54182 22626 -54158
rect 22544 -54216 22568 -54182
rect 22602 -54216 22626 -54182
rect 22544 -54240 22626 -54216
rect 23562 -54182 23644 -54158
rect 23562 -54216 23586 -54182
rect 23620 -54216 23644 -54182
rect 23562 -54240 23644 -54216
rect 24580 -54182 24662 -54158
rect 24580 -54216 24604 -54182
rect 24638 -54216 24662 -54182
rect 24580 -54240 24662 -54216
rect 25598 -54182 25680 -54158
rect 25598 -54216 25622 -54182
rect 25656 -54216 25680 -54182
rect 25598 -54240 25680 -54216
rect 28518 -54498 28600 -54474
rect 28518 -54532 28542 -54498
rect 28576 -54532 28600 -54498
rect 28518 -54556 28600 -54532
rect 29536 -54498 29618 -54474
rect 29536 -54532 29560 -54498
rect 29594 -54532 29618 -54498
rect 29536 -54556 29618 -54532
rect 30554 -54498 30636 -54474
rect 30554 -54532 30578 -54498
rect 30612 -54532 30636 -54498
rect 30554 -54556 30636 -54532
rect 31572 -54498 31654 -54474
rect 31572 -54532 31596 -54498
rect 31630 -54532 31654 -54498
rect 31572 -54556 31654 -54532
rect 32590 -54498 32672 -54474
rect 32590 -54532 32614 -54498
rect 32648 -54532 32672 -54498
rect 32590 -54556 32672 -54532
rect 33608 -54498 33690 -54474
rect 33608 -54532 33632 -54498
rect 33666 -54532 33690 -54498
rect 33608 -54556 33690 -54532
rect 34626 -54498 34708 -54474
rect 34626 -54532 34650 -54498
rect 34684 -54532 34708 -54498
rect 34626 -54556 34708 -54532
rect 35644 -54498 35726 -54474
rect 35644 -54532 35668 -54498
rect 35702 -54532 35726 -54498
rect 35644 -54556 35726 -54532
rect 36662 -54498 36744 -54474
rect 36662 -54532 36686 -54498
rect 36720 -54532 36744 -54498
rect 36662 -54556 36744 -54532
rect 37680 -54498 37762 -54474
rect 37680 -54532 37704 -54498
rect 37738 -54532 37762 -54498
rect 37680 -54556 37762 -54532
rect 38698 -54498 38780 -54474
rect 38698 -54532 38722 -54498
rect 38756 -54532 38780 -54498
rect 38698 -54556 38780 -54532
rect 39716 -54498 39798 -54474
rect 39716 -54532 39740 -54498
rect 39774 -54532 39798 -54498
rect 39716 -54556 39798 -54532
rect 40734 -54498 40816 -54474
rect 40734 -54532 40758 -54498
rect 40792 -54532 40816 -54498
rect 40734 -54556 40816 -54532
rect 41752 -54498 41834 -54474
rect 41752 -54532 41776 -54498
rect 41810 -54532 41834 -54498
rect 41752 -54556 41834 -54532
rect 42770 -54498 42852 -54474
rect 42770 -54532 42794 -54498
rect 42828 -54532 42852 -54498
rect 42770 -54556 42852 -54532
rect 43788 -54498 43870 -54474
rect 43788 -54532 43812 -54498
rect 43846 -54532 43870 -54498
rect 43788 -54556 43870 -54532
rect 44806 -54498 44888 -54474
rect 44806 -54532 44830 -54498
rect 44864 -54532 44888 -54498
rect 44806 -54556 44888 -54532
rect 45824 -54498 45906 -54474
rect 45824 -54532 45848 -54498
rect 45882 -54532 45906 -54498
rect 45824 -54556 45906 -54532
rect 46842 -54498 46924 -54474
rect 46842 -54532 46866 -54498
rect 46900 -54532 46924 -54498
rect 46842 -54556 46924 -54532
rect 47860 -54498 47942 -54474
rect 47860 -54532 47884 -54498
rect 47918 -54532 47942 -54498
rect 47860 -54556 47942 -54532
rect 15418 -55288 15500 -55264
rect 15418 -55322 15442 -55288
rect 15476 -55322 15500 -55288
rect 15418 -55346 15500 -55322
rect 16436 -55288 16518 -55264
rect 16436 -55322 16460 -55288
rect 16494 -55322 16518 -55288
rect 16436 -55346 16518 -55322
rect 17454 -55288 17536 -55264
rect 17454 -55322 17478 -55288
rect 17512 -55322 17536 -55288
rect 17454 -55346 17536 -55322
rect 18472 -55288 18554 -55264
rect 18472 -55322 18496 -55288
rect 18530 -55322 18554 -55288
rect 18472 -55346 18554 -55322
rect 19490 -55288 19572 -55264
rect 19490 -55322 19514 -55288
rect 19548 -55322 19572 -55288
rect 19490 -55346 19572 -55322
rect 20508 -55288 20590 -55264
rect 20508 -55322 20532 -55288
rect 20566 -55322 20590 -55288
rect 20508 -55346 20590 -55322
rect 21526 -55288 21608 -55264
rect 21526 -55322 21550 -55288
rect 21584 -55322 21608 -55288
rect 21526 -55346 21608 -55322
rect 22544 -55288 22626 -55264
rect 22544 -55322 22568 -55288
rect 22602 -55322 22626 -55288
rect 22544 -55346 22626 -55322
rect 23562 -55288 23644 -55264
rect 23562 -55322 23586 -55288
rect 23620 -55322 23644 -55288
rect 23562 -55346 23644 -55322
rect 24580 -55288 24662 -55264
rect 24580 -55322 24604 -55288
rect 24638 -55322 24662 -55288
rect 24580 -55346 24662 -55322
rect 25598 -55288 25680 -55264
rect 25598 -55322 25622 -55288
rect 25656 -55322 25680 -55288
rect 25598 -55346 25680 -55322
rect 28518 -55734 28600 -55710
rect 28518 -55768 28542 -55734
rect 28576 -55768 28600 -55734
rect 28518 -55792 28600 -55768
rect 29536 -55734 29618 -55710
rect 29536 -55768 29560 -55734
rect 29594 -55768 29618 -55734
rect 29536 -55792 29618 -55768
rect 30554 -55734 30636 -55710
rect 30554 -55768 30578 -55734
rect 30612 -55768 30636 -55734
rect 30554 -55792 30636 -55768
rect 31572 -55734 31654 -55710
rect 31572 -55768 31596 -55734
rect 31630 -55768 31654 -55734
rect 31572 -55792 31654 -55768
rect 32590 -55734 32672 -55710
rect 32590 -55768 32614 -55734
rect 32648 -55768 32672 -55734
rect 32590 -55792 32672 -55768
rect 33608 -55734 33690 -55710
rect 33608 -55768 33632 -55734
rect 33666 -55768 33690 -55734
rect 33608 -55792 33690 -55768
rect 34626 -55734 34708 -55710
rect 34626 -55768 34650 -55734
rect 34684 -55768 34708 -55734
rect 34626 -55792 34708 -55768
rect 35644 -55734 35726 -55710
rect 35644 -55768 35668 -55734
rect 35702 -55768 35726 -55734
rect 35644 -55792 35726 -55768
rect 36662 -55734 36744 -55710
rect 36662 -55768 36686 -55734
rect 36720 -55768 36744 -55734
rect 36662 -55792 36744 -55768
rect 37680 -55734 37762 -55710
rect 37680 -55768 37704 -55734
rect 37738 -55768 37762 -55734
rect 37680 -55792 37762 -55768
rect 38698 -55734 38780 -55710
rect 38698 -55768 38722 -55734
rect 38756 -55768 38780 -55734
rect 38698 -55792 38780 -55768
rect 39716 -55734 39798 -55710
rect 39716 -55768 39740 -55734
rect 39774 -55768 39798 -55734
rect 39716 -55792 39798 -55768
rect 40734 -55734 40816 -55710
rect 40734 -55768 40758 -55734
rect 40792 -55768 40816 -55734
rect 40734 -55792 40816 -55768
rect 41752 -55734 41834 -55710
rect 41752 -55768 41776 -55734
rect 41810 -55768 41834 -55734
rect 41752 -55792 41834 -55768
rect 42770 -55734 42852 -55710
rect 42770 -55768 42794 -55734
rect 42828 -55768 42852 -55734
rect 42770 -55792 42852 -55768
rect 43788 -55734 43870 -55710
rect 43788 -55768 43812 -55734
rect 43846 -55768 43870 -55734
rect 43788 -55792 43870 -55768
rect 44806 -55734 44888 -55710
rect 44806 -55768 44830 -55734
rect 44864 -55768 44888 -55734
rect 44806 -55792 44888 -55768
rect 45824 -55734 45906 -55710
rect 45824 -55768 45848 -55734
rect 45882 -55768 45906 -55734
rect 45824 -55792 45906 -55768
rect 46842 -55734 46924 -55710
rect 46842 -55768 46866 -55734
rect 46900 -55768 46924 -55734
rect 46842 -55792 46924 -55768
rect 47860 -55734 47942 -55710
rect 47860 -55768 47884 -55734
rect 47918 -55768 47942 -55734
rect 47860 -55792 47942 -55768
rect 15418 -56630 15500 -56606
rect 15418 -56664 15442 -56630
rect 15476 -56664 15500 -56630
rect 15418 -56688 15500 -56664
rect 16436 -56630 16518 -56606
rect 16436 -56664 16460 -56630
rect 16494 -56664 16518 -56630
rect 16436 -56688 16518 -56664
rect 17454 -56630 17536 -56606
rect 17454 -56664 17478 -56630
rect 17512 -56664 17536 -56630
rect 17454 -56688 17536 -56664
rect 18472 -56630 18554 -56606
rect 18472 -56664 18496 -56630
rect 18530 -56664 18554 -56630
rect 18472 -56688 18554 -56664
rect 19490 -56630 19572 -56606
rect 19490 -56664 19514 -56630
rect 19548 -56664 19572 -56630
rect 19490 -56688 19572 -56664
rect 20508 -56630 20590 -56606
rect 20508 -56664 20532 -56630
rect 20566 -56664 20590 -56630
rect 20508 -56688 20590 -56664
rect 21526 -56630 21608 -56606
rect 21526 -56664 21550 -56630
rect 21584 -56664 21608 -56630
rect 21526 -56688 21608 -56664
rect 22544 -56630 22626 -56606
rect 22544 -56664 22568 -56630
rect 22602 -56664 22626 -56630
rect 22544 -56688 22626 -56664
rect 23562 -56630 23644 -56606
rect 23562 -56664 23586 -56630
rect 23620 -56664 23644 -56630
rect 23562 -56688 23644 -56664
rect 24580 -56630 24662 -56606
rect 24580 -56664 24604 -56630
rect 24638 -56664 24662 -56630
rect 24580 -56688 24662 -56664
rect 25598 -56630 25680 -56606
rect 25598 -56664 25622 -56630
rect 25656 -56664 25680 -56630
rect 25598 -56688 25680 -56664
rect 28530 -56980 28612 -56956
rect 28530 -57014 28554 -56980
rect 28588 -57014 28612 -56980
rect 28530 -57038 28612 -57014
rect 29548 -56980 29630 -56956
rect 29548 -57014 29572 -56980
rect 29606 -57014 29630 -56980
rect 29548 -57038 29630 -57014
rect 30566 -56980 30648 -56956
rect 30566 -57014 30590 -56980
rect 30624 -57014 30648 -56980
rect 30566 -57038 30648 -57014
rect 31584 -56980 31666 -56956
rect 31584 -57014 31608 -56980
rect 31642 -57014 31666 -56980
rect 31584 -57038 31666 -57014
rect 32602 -56980 32684 -56956
rect 32602 -57014 32626 -56980
rect 32660 -57014 32684 -56980
rect 32602 -57038 32684 -57014
rect 33620 -56980 33702 -56956
rect 33620 -57014 33644 -56980
rect 33678 -57014 33702 -56980
rect 33620 -57038 33702 -57014
rect 34638 -56980 34720 -56956
rect 34638 -57014 34662 -56980
rect 34696 -57014 34720 -56980
rect 34638 -57038 34720 -57014
rect 35656 -56980 35738 -56956
rect 35656 -57014 35680 -56980
rect 35714 -57014 35738 -56980
rect 35656 -57038 35738 -57014
rect 36674 -56980 36756 -56956
rect 36674 -57014 36698 -56980
rect 36732 -57014 36756 -56980
rect 36674 -57038 36756 -57014
rect 37692 -56980 37774 -56956
rect 37692 -57014 37716 -56980
rect 37750 -57014 37774 -56980
rect 37692 -57038 37774 -57014
rect 38710 -56980 38792 -56956
rect 38710 -57014 38734 -56980
rect 38768 -57014 38792 -56980
rect 38710 -57038 38792 -57014
rect 39728 -56980 39810 -56956
rect 39728 -57014 39752 -56980
rect 39786 -57014 39810 -56980
rect 39728 -57038 39810 -57014
rect 40746 -56980 40828 -56956
rect 40746 -57014 40770 -56980
rect 40804 -57014 40828 -56980
rect 40746 -57038 40828 -57014
rect 41764 -56980 41846 -56956
rect 41764 -57014 41788 -56980
rect 41822 -57014 41846 -56980
rect 41764 -57038 41846 -57014
rect 42782 -56980 42864 -56956
rect 42782 -57014 42806 -56980
rect 42840 -57014 42864 -56980
rect 42782 -57038 42864 -57014
rect 43800 -56980 43882 -56956
rect 43800 -57014 43824 -56980
rect 43858 -57014 43882 -56980
rect 43800 -57038 43882 -57014
rect 44818 -56980 44900 -56956
rect 44818 -57014 44842 -56980
rect 44876 -57014 44900 -56980
rect 44818 -57038 44900 -57014
rect 45836 -56980 45918 -56956
rect 45836 -57014 45860 -56980
rect 45894 -57014 45918 -56980
rect 45836 -57038 45918 -57014
rect 46854 -56980 46936 -56956
rect 46854 -57014 46878 -56980
rect 46912 -57014 46936 -56980
rect 46854 -57038 46936 -57014
rect 47872 -56980 47954 -56956
rect 47872 -57014 47896 -56980
rect 47930 -57014 47954 -56980
rect 47872 -57038 47954 -57014
rect 15228 -58076 15310 -58052
rect 15228 -58110 15252 -58076
rect 15286 -58110 15310 -58076
rect 15228 -58134 15310 -58110
rect 16246 -58076 16328 -58052
rect 16246 -58110 16270 -58076
rect 16304 -58110 16328 -58076
rect 16246 -58134 16328 -58110
rect 17264 -58076 17346 -58052
rect 17264 -58110 17288 -58076
rect 17322 -58110 17346 -58076
rect 17264 -58134 17346 -58110
rect 18282 -58076 18364 -58052
rect 18282 -58110 18306 -58076
rect 18340 -58110 18364 -58076
rect 18282 -58134 18364 -58110
rect 19300 -58076 19382 -58052
rect 19300 -58110 19324 -58076
rect 19358 -58110 19382 -58076
rect 19300 -58134 19382 -58110
rect 20318 -58076 20400 -58052
rect 20318 -58110 20342 -58076
rect 20376 -58110 20400 -58076
rect 20318 -58134 20400 -58110
rect 21336 -58076 21418 -58052
rect 21336 -58110 21360 -58076
rect 21394 -58110 21418 -58076
rect 21336 -58134 21418 -58110
rect 22354 -58076 22436 -58052
rect 22354 -58110 22378 -58076
rect 22412 -58110 22436 -58076
rect 22354 -58134 22436 -58110
rect 23372 -58076 23454 -58052
rect 23372 -58110 23396 -58076
rect 23430 -58110 23454 -58076
rect 23372 -58134 23454 -58110
rect 24390 -58076 24472 -58052
rect 24390 -58110 24414 -58076
rect 24448 -58110 24472 -58076
rect 24390 -58134 24472 -58110
rect 25408 -58076 25490 -58052
rect 25408 -58110 25432 -58076
rect 25466 -58110 25490 -58076
rect 25408 -58134 25490 -58110
rect 28518 -58158 28600 -58134
rect 28518 -58192 28542 -58158
rect 28576 -58192 28600 -58158
rect 28518 -58216 28600 -58192
rect 29536 -58158 29618 -58134
rect 29536 -58192 29560 -58158
rect 29594 -58192 29618 -58158
rect 29536 -58216 29618 -58192
rect 30554 -58158 30636 -58134
rect 30554 -58192 30578 -58158
rect 30612 -58192 30636 -58158
rect 30554 -58216 30636 -58192
rect 31572 -58158 31654 -58134
rect 31572 -58192 31596 -58158
rect 31630 -58192 31654 -58158
rect 31572 -58216 31654 -58192
rect 32590 -58158 32672 -58134
rect 32590 -58192 32614 -58158
rect 32648 -58192 32672 -58158
rect 32590 -58216 32672 -58192
rect 33608 -58158 33690 -58134
rect 33608 -58192 33632 -58158
rect 33666 -58192 33690 -58158
rect 33608 -58216 33690 -58192
rect 34626 -58158 34708 -58134
rect 34626 -58192 34650 -58158
rect 34684 -58192 34708 -58158
rect 34626 -58216 34708 -58192
rect 35644 -58158 35726 -58134
rect 35644 -58192 35668 -58158
rect 35702 -58192 35726 -58158
rect 35644 -58216 35726 -58192
rect 36662 -58158 36744 -58134
rect 36662 -58192 36686 -58158
rect 36720 -58192 36744 -58158
rect 36662 -58216 36744 -58192
rect 37680 -58158 37762 -58134
rect 37680 -58192 37704 -58158
rect 37738 -58192 37762 -58158
rect 37680 -58216 37762 -58192
rect 38698 -58158 38780 -58134
rect 38698 -58192 38722 -58158
rect 38756 -58192 38780 -58158
rect 38698 -58216 38780 -58192
rect 39716 -58158 39798 -58134
rect 39716 -58192 39740 -58158
rect 39774 -58192 39798 -58158
rect 39716 -58216 39798 -58192
rect 40734 -58158 40816 -58134
rect 40734 -58192 40758 -58158
rect 40792 -58192 40816 -58158
rect 40734 -58216 40816 -58192
rect 41752 -58158 41834 -58134
rect 41752 -58192 41776 -58158
rect 41810 -58192 41834 -58158
rect 41752 -58216 41834 -58192
rect 42770 -58158 42852 -58134
rect 42770 -58192 42794 -58158
rect 42828 -58192 42852 -58158
rect 42770 -58216 42852 -58192
rect 43788 -58158 43870 -58134
rect 43788 -58192 43812 -58158
rect 43846 -58192 43870 -58158
rect 43788 -58216 43870 -58192
rect 44806 -58158 44888 -58134
rect 44806 -58192 44830 -58158
rect 44864 -58192 44888 -58158
rect 44806 -58216 44888 -58192
rect 45824 -58158 45906 -58134
rect 45824 -58192 45848 -58158
rect 45882 -58192 45906 -58158
rect 45824 -58216 45906 -58192
rect 46842 -58158 46924 -58134
rect 46842 -58192 46866 -58158
rect 46900 -58192 46924 -58158
rect 46842 -58216 46924 -58192
rect 47860 -58158 47942 -58134
rect 47860 -58192 47884 -58158
rect 47918 -58192 47942 -58158
rect 47860 -58216 47942 -58192
rect 13122 -59100 13222 -59038
rect 56370 -43604 56470 -43070
rect 57806 -42562 57902 -42528
rect 58090 -42562 58186 -42528
rect 57806 -42624 57840 -42562
rect 58152 -42624 58186 -42562
rect 57806 -42980 57840 -42918
rect 58152 -42980 58186 -42918
rect 57806 -43014 57902 -42980
rect 58090 -43014 58186 -42980
rect 57628 -43604 57728 -43144
rect 56370 -43704 56526 -43604
rect 57510 -43704 57728 -43604
rect 50266 -59100 50366 -59038
rect 13122 -59200 13284 -59100
rect 50204 -59200 50366 -59100
rect -27684 -67866 -27522 -67766
rect -25522 -67866 -25360 -67766
rect -27684 -67928 -27584 -67866
rect -25460 -67928 -25360 -67866
rect -27684 -69710 -27584 -69648
rect -25460 -69710 -25360 -69648
rect -27684 -69810 -27522 -69710
rect -25522 -69810 -25360 -69710
rect -23684 -67866 -23522 -67766
rect -21522 -67866 -21360 -67766
rect -23684 -67928 -23584 -67866
rect -21460 -67928 -21360 -67866
rect -23684 -69710 -23584 -69648
rect -21460 -69710 -21360 -69648
rect -23684 -69810 -23522 -69710
rect -21522 -69810 -21360 -69710
rect -19684 -67866 -19522 -67766
rect -17522 -67866 -17360 -67766
rect -19684 -67928 -19584 -67866
rect -17460 -67928 -17360 -67866
rect -19684 -69710 -19584 -69648
rect -17460 -69710 -17360 -69648
rect -19684 -69810 -19522 -69710
rect -17522 -69810 -17360 -69710
rect -15684 -67866 -15522 -67766
rect -13522 -67866 -13360 -67766
rect -15684 -67928 -15584 -67866
rect -13460 -67928 -13360 -67866
rect -15684 -69710 -15584 -69648
rect -13460 -69710 -13360 -69648
rect -15684 -69810 -15522 -69710
rect -13522 -69810 -13360 -69710
rect -11684 -67866 -11522 -67766
rect -9522 -67866 -9360 -67766
rect -11684 -67928 -11584 -67866
rect -9460 -67928 -9360 -67866
rect -11684 -69710 -11584 -69648
rect -9460 -69710 -9360 -69648
rect -11684 -69810 -11522 -69710
rect -9522 -69810 -9360 -69710
rect -7684 -67866 -7522 -67766
rect -5522 -67866 -5360 -67766
rect -7684 -67928 -7584 -67866
rect -5460 -67928 -5360 -67866
rect -7684 -69710 -7584 -69648
rect -5460 -69710 -5360 -69648
rect -7684 -69810 -7522 -69710
rect -5522 -69810 -5360 -69710
rect -3684 -67866 -3522 -67766
rect -1522 -67866 -1360 -67766
rect -3684 -67928 -3584 -67866
rect -1460 -67928 -1360 -67866
rect -3684 -69710 -3584 -69648
rect -1460 -69710 -1360 -69648
rect -3684 -69810 -3522 -69710
rect -1522 -69810 -1360 -69710
rect 316 -67866 478 -67766
rect 2478 -67866 2640 -67766
rect 316 -67928 416 -67866
rect 2540 -67928 2640 -67866
rect 316 -69710 416 -69648
rect 2540 -69710 2640 -69648
rect 316 -69810 478 -69710
rect 2478 -69810 2640 -69710
rect 4316 -67866 4478 -67766
rect 6478 -67866 6640 -67766
rect 4316 -67928 4416 -67866
rect 6540 -67928 6640 -67866
rect 4316 -69710 4416 -69648
rect 6540 -69710 6640 -69648
rect 4316 -69810 4478 -69710
rect 6478 -69810 6640 -69710
rect -27684 -70486 -27522 -70386
rect -25522 -70486 -25360 -70386
rect -27684 -70548 -27584 -70486
rect -25460 -70548 -25360 -70486
rect -27684 -72330 -27584 -72268
rect -25460 -72330 -25360 -72268
rect -27684 -72430 -27522 -72330
rect -25522 -72430 -25360 -72330
rect -23684 -70486 -23522 -70386
rect -21522 -70486 -21360 -70386
rect -23684 -70548 -23584 -70486
rect -21460 -70548 -21360 -70486
rect -23684 -72330 -23584 -72268
rect -21460 -72330 -21360 -72268
rect -23684 -72430 -23522 -72330
rect -21522 -72430 -21360 -72330
rect -19684 -70486 -19522 -70386
rect -17522 -70486 -17360 -70386
rect -19684 -70548 -19584 -70486
rect -17460 -70548 -17360 -70486
rect -19684 -72330 -19584 -72268
rect -17460 -72330 -17360 -72268
rect -19684 -72430 -19522 -72330
rect -17522 -72430 -17360 -72330
rect -15684 -70486 -15522 -70386
rect -13522 -70486 -13360 -70386
rect -15684 -70548 -15584 -70486
rect -13460 -70548 -13360 -70486
rect -15684 -72330 -15584 -72268
rect -13460 -72330 -13360 -72268
rect -15684 -72430 -15522 -72330
rect -13522 -72430 -13360 -72330
rect -11684 -70486 -11522 -70386
rect -9522 -70486 -9360 -70386
rect -11684 -70548 -11584 -70486
rect -9460 -70548 -9360 -70486
rect -11684 -72330 -11584 -72268
rect -9460 -72330 -9360 -72268
rect -11684 -72430 -11522 -72330
rect -9522 -72430 -9360 -72330
rect -7684 -70486 -7522 -70386
rect -5522 -70486 -5360 -70386
rect -7684 -70548 -7584 -70486
rect -5460 -70548 -5360 -70486
rect -7684 -72330 -7584 -72268
rect -5460 -72330 -5360 -72268
rect -7684 -72430 -7522 -72330
rect -5522 -72430 -5360 -72330
rect -3684 -70486 -3522 -70386
rect -1522 -70486 -1360 -70386
rect -3684 -70548 -3584 -70486
rect -1460 -70548 -1360 -70486
rect -3684 -72330 -3584 -72268
rect -1460 -72330 -1360 -72268
rect -3684 -72430 -3522 -72330
rect -1522 -72430 -1360 -72330
rect 316 -70486 478 -70386
rect 2478 -70486 2640 -70386
rect 316 -70548 416 -70486
rect 2540 -70548 2640 -70486
rect 316 -72330 416 -72268
rect 2540 -72330 2640 -72268
rect 316 -72430 478 -72330
rect 2478 -72430 2640 -72330
rect 4316 -70486 4478 -70386
rect 6478 -70486 6640 -70386
rect 4316 -70548 4416 -70486
rect 6540 -70548 6640 -70486
rect 4316 -72330 4416 -72268
rect 6540 -72330 6640 -72268
rect 4316 -72430 4478 -72330
rect 6478 -72430 6640 -72330
<< nsubdiff >>
rect 25822 -27756 25984 -27656
rect 50104 -27756 50266 -27656
rect 25822 -27818 25922 -27756
rect 50166 -27818 50266 -27756
rect 32416 -30200 32498 -30174
rect 32416 -30234 32440 -30200
rect 32474 -30234 32498 -30200
rect 32416 -30258 32498 -30234
rect 33434 -30200 33516 -30174
rect 33434 -30234 33458 -30200
rect 33492 -30234 33516 -30200
rect 33434 -30258 33516 -30234
rect 34452 -30200 34534 -30174
rect 34452 -30234 34476 -30200
rect 34510 -30234 34534 -30200
rect 34452 -30258 34534 -30234
rect 35470 -30200 35552 -30174
rect 35470 -30234 35494 -30200
rect 35528 -30234 35552 -30200
rect 35470 -30258 35552 -30234
rect 36488 -30200 36570 -30174
rect 36488 -30234 36512 -30200
rect 36546 -30234 36570 -30200
rect 36488 -30258 36570 -30234
rect 37506 -30200 37588 -30174
rect 37506 -30234 37530 -30200
rect 37564 -30234 37588 -30200
rect 37506 -30258 37588 -30234
rect 38524 -30200 38606 -30174
rect 38524 -30234 38548 -30200
rect 38582 -30234 38606 -30200
rect 38524 -30258 38606 -30234
rect 39542 -30200 39624 -30174
rect 39542 -30234 39566 -30200
rect 39600 -30234 39624 -30200
rect 39542 -30258 39624 -30234
rect 40560 -30200 40642 -30174
rect 40560 -30234 40584 -30200
rect 40618 -30234 40642 -30200
rect 40560 -30258 40642 -30234
rect 41578 -30200 41660 -30174
rect 41578 -30234 41602 -30200
rect 41636 -30234 41660 -30200
rect 41578 -30258 41660 -30234
rect 42596 -30200 42678 -30174
rect 42596 -30234 42620 -30200
rect 42654 -30234 42678 -30200
rect 42596 -30258 42678 -30234
rect 43614 -30200 43696 -30174
rect 43614 -30234 43638 -30200
rect 43672 -30234 43696 -30200
rect 43614 -30258 43696 -30234
rect 44632 -30200 44714 -30174
rect 44632 -30234 44656 -30200
rect 44690 -30234 44714 -30200
rect 44632 -30258 44714 -30234
rect 45650 -30200 45732 -30174
rect 45650 -30234 45674 -30200
rect 45708 -30234 45732 -30200
rect 45650 -30258 45732 -30234
rect 46668 -30200 46750 -30174
rect 46668 -30234 46692 -30200
rect 46726 -30234 46750 -30200
rect 46668 -30258 46750 -30234
rect 47686 -30200 47768 -30174
rect 47686 -30234 47710 -30200
rect 47744 -30234 47768 -30200
rect 47686 -30258 47768 -30234
rect 32438 -31354 32520 -31328
rect 32438 -31388 32462 -31354
rect 32496 -31388 32520 -31354
rect 32438 -31412 32520 -31388
rect 33456 -31354 33538 -31328
rect 33456 -31388 33480 -31354
rect 33514 -31388 33538 -31354
rect 33456 -31412 33538 -31388
rect 34474 -31354 34556 -31328
rect 34474 -31388 34498 -31354
rect 34532 -31388 34556 -31354
rect 34474 -31412 34556 -31388
rect 35492 -31354 35574 -31328
rect 35492 -31388 35516 -31354
rect 35550 -31388 35574 -31354
rect 35492 -31412 35574 -31388
rect 36510 -31354 36592 -31328
rect 36510 -31388 36534 -31354
rect 36568 -31388 36592 -31354
rect 36510 -31412 36592 -31388
rect 37528 -31354 37610 -31328
rect 37528 -31388 37552 -31354
rect 37586 -31388 37610 -31354
rect 37528 -31412 37610 -31388
rect 38546 -31354 38628 -31328
rect 38546 -31388 38570 -31354
rect 38604 -31388 38628 -31354
rect 38546 -31412 38628 -31388
rect 39564 -31354 39646 -31328
rect 39564 -31388 39588 -31354
rect 39622 -31388 39646 -31354
rect 39564 -31412 39646 -31388
rect 40582 -31354 40664 -31328
rect 40582 -31388 40606 -31354
rect 40640 -31388 40664 -31354
rect 40582 -31412 40664 -31388
rect 41600 -31354 41682 -31328
rect 41600 -31388 41624 -31354
rect 41658 -31388 41682 -31354
rect 41600 -31412 41682 -31388
rect 42618 -31354 42700 -31328
rect 42618 -31388 42642 -31354
rect 42676 -31388 42700 -31354
rect 42618 -31412 42700 -31388
rect 43636 -31354 43718 -31328
rect 43636 -31388 43660 -31354
rect 43694 -31388 43718 -31354
rect 43636 -31412 43718 -31388
rect 44654 -31354 44736 -31328
rect 44654 -31388 44678 -31354
rect 44712 -31388 44736 -31354
rect 44654 -31412 44736 -31388
rect 45672 -31354 45754 -31328
rect 45672 -31388 45696 -31354
rect 45730 -31388 45754 -31354
rect 45672 -31412 45754 -31388
rect 46690 -31354 46772 -31328
rect 46690 -31388 46714 -31354
rect 46748 -31388 46772 -31354
rect 46690 -31412 46772 -31388
rect 47708 -31354 47790 -31328
rect 47708 -31388 47732 -31354
rect 47766 -31388 47790 -31354
rect 47708 -31412 47790 -31388
rect 32416 -32486 32498 -32460
rect 32416 -32520 32440 -32486
rect 32474 -32520 32498 -32486
rect 32416 -32544 32498 -32520
rect 33434 -32486 33516 -32460
rect 33434 -32520 33458 -32486
rect 33492 -32520 33516 -32486
rect 33434 -32544 33516 -32520
rect 34452 -32486 34534 -32460
rect 34452 -32520 34476 -32486
rect 34510 -32520 34534 -32486
rect 34452 -32544 34534 -32520
rect 35470 -32486 35552 -32460
rect 35470 -32520 35494 -32486
rect 35528 -32520 35552 -32486
rect 35470 -32544 35552 -32520
rect 36488 -32486 36570 -32460
rect 36488 -32520 36512 -32486
rect 36546 -32520 36570 -32486
rect 36488 -32544 36570 -32520
rect 37506 -32486 37588 -32460
rect 37506 -32520 37530 -32486
rect 37564 -32520 37588 -32486
rect 37506 -32544 37588 -32520
rect 38524 -32486 38606 -32460
rect 38524 -32520 38548 -32486
rect 38582 -32520 38606 -32486
rect 38524 -32544 38606 -32520
rect 39542 -32486 39624 -32460
rect 39542 -32520 39566 -32486
rect 39600 -32520 39624 -32486
rect 39542 -32544 39624 -32520
rect 40560 -32486 40642 -32460
rect 40560 -32520 40584 -32486
rect 40618 -32520 40642 -32486
rect 40560 -32544 40642 -32520
rect 41578 -32486 41660 -32460
rect 41578 -32520 41602 -32486
rect 41636 -32520 41660 -32486
rect 41578 -32544 41660 -32520
rect 42596 -32486 42678 -32460
rect 42596 -32520 42620 -32486
rect 42654 -32520 42678 -32486
rect 42596 -32544 42678 -32520
rect 43614 -32486 43696 -32460
rect 43614 -32520 43638 -32486
rect 43672 -32520 43696 -32486
rect 43614 -32544 43696 -32520
rect 44632 -32486 44714 -32460
rect 44632 -32520 44656 -32486
rect 44690 -32520 44714 -32486
rect 44632 -32544 44714 -32520
rect 45650 -32486 45732 -32460
rect 45650 -32520 45674 -32486
rect 45708 -32520 45732 -32486
rect 45650 -32544 45732 -32520
rect 46668 -32486 46750 -32460
rect 46668 -32520 46692 -32486
rect 46726 -32520 46750 -32486
rect 46668 -32544 46750 -32520
rect 47686 -32486 47768 -32460
rect 47686 -32520 47710 -32486
rect 47744 -32520 47768 -32486
rect 47686 -32544 47768 -32520
rect 32416 -33868 32498 -33842
rect 32416 -33902 32440 -33868
rect 32474 -33902 32498 -33868
rect 32416 -33926 32498 -33902
rect 33434 -33868 33516 -33842
rect 33434 -33902 33458 -33868
rect 33492 -33902 33516 -33868
rect 33434 -33926 33516 -33902
rect 34452 -33868 34534 -33842
rect 34452 -33902 34476 -33868
rect 34510 -33902 34534 -33868
rect 34452 -33926 34534 -33902
rect 35470 -33868 35552 -33842
rect 35470 -33902 35494 -33868
rect 35528 -33902 35552 -33868
rect 35470 -33926 35552 -33902
rect 36488 -33868 36570 -33842
rect 36488 -33902 36512 -33868
rect 36546 -33902 36570 -33868
rect 36488 -33926 36570 -33902
rect 37506 -33868 37588 -33842
rect 37506 -33902 37530 -33868
rect 37564 -33902 37588 -33868
rect 37506 -33926 37588 -33902
rect 38524 -33868 38606 -33842
rect 38524 -33902 38548 -33868
rect 38582 -33902 38606 -33868
rect 38524 -33926 38606 -33902
rect 39542 -33868 39624 -33842
rect 39542 -33902 39566 -33868
rect 39600 -33902 39624 -33868
rect 39542 -33926 39624 -33902
rect 40560 -33868 40642 -33842
rect 40560 -33902 40584 -33868
rect 40618 -33902 40642 -33868
rect 40560 -33926 40642 -33902
rect 41578 -33868 41660 -33842
rect 41578 -33902 41602 -33868
rect 41636 -33902 41660 -33868
rect 41578 -33926 41660 -33902
rect 42596 -33868 42678 -33842
rect 42596 -33902 42620 -33868
rect 42654 -33902 42678 -33868
rect 42596 -33926 42678 -33902
rect 43614 -33868 43696 -33842
rect 43614 -33902 43638 -33868
rect 43672 -33902 43696 -33868
rect 43614 -33926 43696 -33902
rect 44632 -33868 44714 -33842
rect 44632 -33902 44656 -33868
rect 44690 -33902 44714 -33868
rect 44632 -33926 44714 -33902
rect 45650 -33868 45732 -33842
rect 45650 -33902 45674 -33868
rect 45708 -33902 45732 -33868
rect 45650 -33926 45732 -33902
rect 46668 -33868 46750 -33842
rect 46668 -33902 46692 -33868
rect 46726 -33902 46750 -33868
rect 46668 -33926 46750 -33902
rect 47686 -33868 47768 -33842
rect 47686 -33902 47710 -33868
rect 47744 -33902 47768 -33868
rect 47686 -33926 47768 -33902
rect 33104 -35216 33186 -35190
rect 33104 -35250 33128 -35216
rect 33162 -35250 33186 -35216
rect 33104 -35274 33186 -35250
rect 34122 -35216 34204 -35190
rect 34122 -35250 34146 -35216
rect 34180 -35250 34204 -35216
rect 34122 -35274 34204 -35250
rect 35140 -35216 35222 -35190
rect 35140 -35250 35164 -35216
rect 35198 -35250 35222 -35216
rect 35140 -35274 35222 -35250
rect 36158 -35216 36240 -35190
rect 36158 -35250 36182 -35216
rect 36216 -35250 36240 -35216
rect 36158 -35274 36240 -35250
rect 37176 -35216 37258 -35190
rect 37176 -35250 37200 -35216
rect 37234 -35250 37258 -35216
rect 37176 -35274 37258 -35250
rect 38194 -35216 38276 -35190
rect 38194 -35250 38218 -35216
rect 38252 -35250 38276 -35216
rect 38194 -35274 38276 -35250
rect 39212 -35216 39294 -35190
rect 39212 -35250 39236 -35216
rect 39270 -35250 39294 -35216
rect 39212 -35274 39294 -35250
rect 40230 -35216 40312 -35190
rect 40230 -35250 40254 -35216
rect 40288 -35250 40312 -35216
rect 40230 -35274 40312 -35250
rect 41248 -35216 41330 -35190
rect 41248 -35250 41272 -35216
rect 41306 -35250 41330 -35216
rect 41248 -35274 41330 -35250
rect 42266 -35216 42348 -35190
rect 42266 -35250 42290 -35216
rect 42324 -35250 42348 -35216
rect 42266 -35274 42348 -35250
rect 43284 -35216 43366 -35190
rect 43284 -35250 43308 -35216
rect 43342 -35250 43366 -35216
rect 43284 -35274 43366 -35250
rect 44302 -35216 44384 -35190
rect 44302 -35250 44326 -35216
rect 44360 -35250 44384 -35216
rect 44302 -35274 44384 -35250
rect 45320 -35216 45402 -35190
rect 45320 -35250 45344 -35216
rect 45378 -35250 45402 -35216
rect 45320 -35274 45402 -35250
rect 46338 -35216 46420 -35190
rect 46338 -35250 46362 -35216
rect 46396 -35250 46420 -35216
rect 46338 -35274 46420 -35250
rect 47356 -35216 47438 -35190
rect 47356 -35250 47380 -35216
rect 47414 -35250 47438 -35216
rect 47356 -35274 47438 -35250
rect 32710 -36494 32792 -36468
rect 32710 -36528 32734 -36494
rect 32768 -36528 32792 -36494
rect 32710 -36552 32792 -36528
rect 33728 -36494 33810 -36468
rect 33728 -36528 33752 -36494
rect 33786 -36528 33810 -36494
rect 33728 -36552 33810 -36528
rect 34746 -36494 34828 -36468
rect 34746 -36528 34770 -36494
rect 34804 -36528 34828 -36494
rect 34746 -36552 34828 -36528
rect 35764 -36494 35846 -36468
rect 35764 -36528 35788 -36494
rect 35822 -36528 35846 -36494
rect 35764 -36552 35846 -36528
rect 36782 -36494 36864 -36468
rect 36782 -36528 36806 -36494
rect 36840 -36528 36864 -36494
rect 36782 -36552 36864 -36528
rect 37800 -36494 37882 -36468
rect 37800 -36528 37824 -36494
rect 37858 -36528 37882 -36494
rect 37800 -36552 37882 -36528
rect 38818 -36494 38900 -36468
rect 38818 -36528 38842 -36494
rect 38876 -36528 38900 -36494
rect 38818 -36552 38900 -36528
rect 39836 -36494 39918 -36468
rect 39836 -36528 39860 -36494
rect 39894 -36528 39918 -36494
rect 39836 -36552 39918 -36528
rect 40854 -36494 40936 -36468
rect 40854 -36528 40878 -36494
rect 40912 -36528 40936 -36494
rect 40854 -36552 40936 -36528
rect 41872 -36494 41954 -36468
rect 41872 -36528 41896 -36494
rect 41930 -36528 41954 -36494
rect 41872 -36552 41954 -36528
rect 42890 -36494 42972 -36468
rect 42890 -36528 42914 -36494
rect 42948 -36528 42972 -36494
rect 42890 -36552 42972 -36528
rect 43908 -36494 43990 -36468
rect 43908 -36528 43932 -36494
rect 43966 -36528 43990 -36494
rect 43908 -36552 43990 -36528
rect 44926 -36494 45008 -36468
rect 44926 -36528 44950 -36494
rect 44984 -36528 45008 -36494
rect 44926 -36552 45008 -36528
rect 45944 -36494 46026 -36468
rect 45944 -36528 45968 -36494
rect 46002 -36528 46026 -36494
rect 45944 -36552 46026 -36528
rect 46962 -36494 47044 -36468
rect 46962 -36528 46986 -36494
rect 47020 -36528 47044 -36494
rect 46962 -36552 47044 -36528
rect 47980 -36494 48062 -36468
rect 47980 -36528 48004 -36494
rect 48038 -36528 48062 -36494
rect 47980 -36552 48062 -36528
rect 28112 -36804 28194 -36778
rect 28112 -36838 28136 -36804
rect 28170 -36838 28194 -36804
rect 28112 -36862 28194 -36838
rect 29130 -36804 29212 -36778
rect 29130 -36838 29154 -36804
rect 29188 -36838 29212 -36804
rect 29130 -36862 29212 -36838
rect 30148 -36804 30230 -36778
rect 30148 -36838 30172 -36804
rect 30206 -36838 30230 -36804
rect 30148 -36862 30230 -36838
rect 31166 -36804 31248 -36778
rect 31166 -36838 31190 -36804
rect 31224 -36838 31248 -36804
rect 31166 -36862 31248 -36838
rect 27588 -37958 27670 -37932
rect 27588 -37992 27612 -37958
rect 27646 -37992 27670 -37958
rect 27588 -38016 27670 -37992
rect 28606 -37958 28688 -37932
rect 28606 -37992 28630 -37958
rect 28664 -37992 28688 -37958
rect 28606 -38016 28688 -37992
rect 29624 -37958 29706 -37932
rect 29624 -37992 29648 -37958
rect 29682 -37992 29706 -37958
rect 29624 -38016 29706 -37992
rect 30642 -37958 30724 -37932
rect 30642 -37992 30666 -37958
rect 30700 -37992 30724 -37958
rect 30642 -38016 30724 -37992
rect 32800 -37942 32882 -37916
rect 32800 -37976 32824 -37942
rect 32858 -37976 32882 -37942
rect 32800 -38000 32882 -37976
rect 33818 -37942 33900 -37916
rect 33818 -37976 33842 -37942
rect 33876 -37976 33900 -37942
rect 33818 -38000 33900 -37976
rect 34836 -37942 34918 -37916
rect 34836 -37976 34860 -37942
rect 34894 -37976 34918 -37942
rect 34836 -38000 34918 -37976
rect 35854 -37942 35936 -37916
rect 35854 -37976 35878 -37942
rect 35912 -37976 35936 -37942
rect 35854 -38000 35936 -37976
rect 36872 -37942 36954 -37916
rect 36872 -37976 36896 -37942
rect 36930 -37976 36954 -37942
rect 36872 -38000 36954 -37976
rect 37890 -37942 37972 -37916
rect 37890 -37976 37914 -37942
rect 37948 -37976 37972 -37942
rect 37890 -38000 37972 -37976
rect 38908 -37942 38990 -37916
rect 38908 -37976 38932 -37942
rect 38966 -37976 38990 -37942
rect 38908 -38000 38990 -37976
rect 39926 -37942 40008 -37916
rect 39926 -37976 39950 -37942
rect 39984 -37976 40008 -37942
rect 39926 -38000 40008 -37976
rect 40944 -37942 41026 -37916
rect 40944 -37976 40968 -37942
rect 41002 -37976 41026 -37942
rect 40944 -38000 41026 -37976
rect 41962 -37942 42044 -37916
rect 41962 -37976 41986 -37942
rect 42020 -37976 42044 -37942
rect 41962 -38000 42044 -37976
rect 42980 -37942 43062 -37916
rect 42980 -37976 43004 -37942
rect 43038 -37976 43062 -37942
rect 42980 -38000 43062 -37976
rect 43998 -37942 44080 -37916
rect 43998 -37976 44022 -37942
rect 44056 -37976 44080 -37942
rect 43998 -38000 44080 -37976
rect 45016 -37942 45098 -37916
rect 45016 -37976 45040 -37942
rect 45074 -37976 45098 -37942
rect 45016 -38000 45098 -37976
rect 46034 -37942 46116 -37916
rect 46034 -37976 46058 -37942
rect 46092 -37976 46116 -37942
rect 46034 -38000 46116 -37976
rect 47052 -37942 47134 -37916
rect 47052 -37976 47076 -37942
rect 47110 -37976 47134 -37942
rect 47052 -38000 47134 -37976
rect 48070 -37942 48152 -37916
rect 48070 -37976 48094 -37942
rect 48128 -37976 48152 -37942
rect 48070 -38000 48152 -37976
rect 27598 -38986 27680 -38960
rect 27598 -39020 27622 -38986
rect 27656 -39020 27680 -38986
rect 27598 -39044 27680 -39020
rect 28616 -38986 28698 -38960
rect 28616 -39020 28640 -38986
rect 28674 -39020 28698 -38986
rect 28616 -39044 28698 -39020
rect 29634 -38986 29716 -38960
rect 29634 -39020 29658 -38986
rect 29692 -39020 29716 -38986
rect 29634 -39044 29716 -39020
rect 30652 -38986 30734 -38960
rect 30652 -39020 30676 -38986
rect 30710 -39020 30734 -38986
rect 30652 -39044 30734 -39020
rect 32824 -39210 32906 -39184
rect 32824 -39244 32848 -39210
rect 32882 -39244 32906 -39210
rect 32824 -39268 32906 -39244
rect 33842 -39210 33924 -39184
rect 33842 -39244 33866 -39210
rect 33900 -39244 33924 -39210
rect 33842 -39268 33924 -39244
rect 34860 -39210 34942 -39184
rect 34860 -39244 34884 -39210
rect 34918 -39244 34942 -39210
rect 34860 -39268 34942 -39244
rect 35878 -39210 35960 -39184
rect 35878 -39244 35902 -39210
rect 35936 -39244 35960 -39210
rect 35878 -39268 35960 -39244
rect 36896 -39210 36978 -39184
rect 36896 -39244 36920 -39210
rect 36954 -39244 36978 -39210
rect 36896 -39268 36978 -39244
rect 37914 -39210 37996 -39184
rect 37914 -39244 37938 -39210
rect 37972 -39244 37996 -39210
rect 37914 -39268 37996 -39244
rect 38932 -39210 39014 -39184
rect 38932 -39244 38956 -39210
rect 38990 -39244 39014 -39210
rect 38932 -39268 39014 -39244
rect 39950 -39210 40032 -39184
rect 39950 -39244 39974 -39210
rect 40008 -39244 40032 -39210
rect 39950 -39268 40032 -39244
rect 40968 -39210 41050 -39184
rect 40968 -39244 40992 -39210
rect 41026 -39244 41050 -39210
rect 40968 -39268 41050 -39244
rect 41986 -39210 42068 -39184
rect 41986 -39244 42010 -39210
rect 42044 -39244 42068 -39210
rect 41986 -39268 42068 -39244
rect 43004 -39210 43086 -39184
rect 43004 -39244 43028 -39210
rect 43062 -39244 43086 -39210
rect 43004 -39268 43086 -39244
rect 44022 -39210 44104 -39184
rect 44022 -39244 44046 -39210
rect 44080 -39244 44104 -39210
rect 44022 -39268 44104 -39244
rect 45040 -39210 45122 -39184
rect 45040 -39244 45064 -39210
rect 45098 -39244 45122 -39210
rect 45040 -39268 45122 -39244
rect 46058 -39210 46140 -39184
rect 46058 -39244 46082 -39210
rect 46116 -39244 46140 -39210
rect 46058 -39268 46140 -39244
rect 47076 -39210 47158 -39184
rect 47076 -39244 47100 -39210
rect 47134 -39244 47158 -39210
rect 47076 -39268 47158 -39244
rect 48094 -39210 48176 -39184
rect 48094 -39244 48118 -39210
rect 48152 -39244 48176 -39210
rect 48094 -39268 48176 -39244
rect 27588 -40014 27670 -39988
rect 27588 -40048 27612 -40014
rect 27646 -40048 27670 -40014
rect 27588 -40072 27670 -40048
rect 28606 -40014 28688 -39988
rect 28606 -40048 28630 -40014
rect 28664 -40048 28688 -40014
rect 28606 -40072 28688 -40048
rect 29624 -40014 29706 -39988
rect 29624 -40048 29648 -40014
rect 29682 -40048 29706 -40014
rect 29624 -40072 29706 -40048
rect 30642 -40014 30724 -39988
rect 30642 -40048 30666 -40014
rect 30700 -40048 30724 -40014
rect 30642 -40072 30724 -40048
rect 32688 -40454 32770 -40428
rect 32688 -40488 32712 -40454
rect 32746 -40488 32770 -40454
rect 32688 -40512 32770 -40488
rect 33706 -40454 33788 -40428
rect 33706 -40488 33730 -40454
rect 33764 -40488 33788 -40454
rect 33706 -40512 33788 -40488
rect 34724 -40454 34806 -40428
rect 34724 -40488 34748 -40454
rect 34782 -40488 34806 -40454
rect 34724 -40512 34806 -40488
rect 35742 -40454 35824 -40428
rect 35742 -40488 35766 -40454
rect 35800 -40488 35824 -40454
rect 35742 -40512 35824 -40488
rect 36760 -40454 36842 -40428
rect 36760 -40488 36784 -40454
rect 36818 -40488 36842 -40454
rect 36760 -40512 36842 -40488
rect 37778 -40454 37860 -40428
rect 37778 -40488 37802 -40454
rect 37836 -40488 37860 -40454
rect 37778 -40512 37860 -40488
rect 38796 -40454 38878 -40428
rect 38796 -40488 38820 -40454
rect 38854 -40488 38878 -40454
rect 38796 -40512 38878 -40488
rect 39814 -40454 39896 -40428
rect 39814 -40488 39838 -40454
rect 39872 -40488 39896 -40454
rect 39814 -40512 39896 -40488
rect 40832 -40454 40914 -40428
rect 40832 -40488 40856 -40454
rect 40890 -40488 40914 -40454
rect 40832 -40512 40914 -40488
rect 41850 -40454 41932 -40428
rect 41850 -40488 41874 -40454
rect 41908 -40488 41932 -40454
rect 41850 -40512 41932 -40488
rect 42868 -40454 42950 -40428
rect 42868 -40488 42892 -40454
rect 42926 -40488 42950 -40454
rect 42868 -40512 42950 -40488
rect 43886 -40454 43968 -40428
rect 43886 -40488 43910 -40454
rect 43944 -40488 43968 -40454
rect 43886 -40512 43968 -40488
rect 44904 -40454 44986 -40428
rect 44904 -40488 44928 -40454
rect 44962 -40488 44986 -40454
rect 44904 -40512 44986 -40488
rect 45922 -40454 46004 -40428
rect 45922 -40488 45946 -40454
rect 45980 -40488 46004 -40454
rect 45922 -40512 46004 -40488
rect 46940 -40454 47022 -40428
rect 46940 -40488 46964 -40454
rect 46998 -40488 47022 -40454
rect 46940 -40512 47022 -40488
rect 47958 -40454 48040 -40428
rect 47958 -40488 47982 -40454
rect 48016 -40488 48040 -40454
rect 47958 -40512 48040 -40488
rect 28112 -41166 28194 -41140
rect 28112 -41200 28136 -41166
rect 28170 -41200 28194 -41166
rect 28112 -41224 28194 -41200
rect 29130 -41166 29212 -41140
rect 29130 -41200 29154 -41166
rect 29188 -41200 29212 -41166
rect 29130 -41224 29212 -41200
rect 30148 -41166 30230 -41140
rect 30148 -41200 30172 -41166
rect 30206 -41200 30230 -41166
rect 30148 -41224 30230 -41200
rect 31166 -41166 31248 -41140
rect 31166 -41200 31190 -41166
rect 31224 -41200 31248 -41166
rect 31166 -41224 31248 -41200
rect 25822 -42226 25922 -42164
rect 50166 -42226 50266 -42164
rect 25822 -42326 25984 -42226
rect 50104 -42326 50266 -42226
rect 52156 -39080 52318 -38980
rect 55358 -39080 55520 -38980
rect 52156 -39142 52256 -39080
rect 55420 -39142 55520 -39080
rect 52156 -42224 52256 -42162
rect 55858 -39080 56020 -38980
rect 58100 -39080 58262 -38980
rect 55858 -39142 55958 -39080
rect 58162 -39142 58262 -39080
rect 55858 -41430 55958 -41368
rect 58162 -41430 58262 -41368
rect 55858 -41530 56020 -41430
rect 58100 -41530 58262 -41430
rect 55420 -42224 55520 -42162
rect 52156 -42324 52318 -42224
rect 55358 -42324 55520 -42224
rect 54104 -42418 54200 -42384
rect 55422 -42418 55518 -42384
rect 54104 -42578 54138 -42418
rect 55484 -42578 55518 -42418
rect 54104 -42966 54138 -42810
rect 55484 -42966 55518 -42810
rect 54104 -43000 54200 -42966
rect 55422 -43000 55518 -42966
rect 10296 -56773 10392 -56739
rect 12010 -56773 12106 -56739
rect 10296 -56835 10330 -56773
rect 12072 -56835 12106 -56773
rect 10296 -57471 10330 -57409
rect 12072 -57471 12106 -57409
rect 10296 -57505 10392 -57471
rect 12010 -57505 12106 -57471
rect -27684 -64526 -27522 -64426
rect -25522 -64526 -25360 -64426
rect -27684 -64588 -27584 -64526
rect -25460 -64588 -25360 -64526
rect -27684 -67430 -27584 -67368
rect -23684 -64526 -23522 -64426
rect -21522 -64526 -21360 -64426
rect -23684 -64588 -23584 -64526
rect -25460 -67430 -25360 -67368
rect -27684 -67530 -27522 -67430
rect -25522 -67530 -25360 -67430
rect -21460 -64588 -21360 -64526
rect -23684 -67430 -23584 -67368
rect -19684 -64526 -19522 -64426
rect -17522 -64526 -17360 -64426
rect -19684 -64588 -19584 -64526
rect -21460 -67430 -21360 -67368
rect -23684 -67530 -23522 -67430
rect -21522 -67530 -21360 -67430
rect -17460 -64588 -17360 -64526
rect -19684 -67430 -19584 -67368
rect -15684 -64526 -15522 -64426
rect -13522 -64526 -13360 -64426
rect -15684 -64588 -15584 -64526
rect -17460 -67430 -17360 -67368
rect -19684 -67530 -19522 -67430
rect -17522 -67530 -17360 -67430
rect -13460 -64588 -13360 -64526
rect -15684 -67430 -15584 -67368
rect -11684 -64526 -11522 -64426
rect -9522 -64526 -9360 -64426
rect -11684 -64588 -11584 -64526
rect -13460 -67430 -13360 -67368
rect -15684 -67530 -15522 -67430
rect -13522 -67530 -13360 -67430
rect -9460 -64588 -9360 -64526
rect -11684 -67430 -11584 -67368
rect -7684 -64526 -7522 -64426
rect -5522 -64526 -5360 -64426
rect -7684 -64588 -7584 -64526
rect -9460 -67430 -9360 -67368
rect -11684 -67530 -11522 -67430
rect -9522 -67530 -9360 -67430
rect -5460 -64588 -5360 -64526
rect -7684 -67430 -7584 -67368
rect -3684 -64526 -3522 -64426
rect -1522 -64526 -1360 -64426
rect -3684 -64588 -3584 -64526
rect -5460 -67430 -5360 -67368
rect -7684 -67530 -7522 -67430
rect -5522 -67530 -5360 -67430
rect -1460 -64588 -1360 -64526
rect -3684 -67430 -3584 -67368
rect 316 -64526 478 -64426
rect 2478 -64526 2640 -64426
rect 316 -64588 416 -64526
rect -1460 -67430 -1360 -67368
rect -3684 -67530 -3522 -67430
rect -1522 -67530 -1360 -67430
rect 2540 -64588 2640 -64526
rect 316 -67430 416 -67368
rect 4316 -64526 4478 -64426
rect 6478 -64526 6640 -64426
rect 4316 -64588 4416 -64526
rect 2540 -67430 2640 -67368
rect 316 -67530 478 -67430
rect 2478 -67530 2640 -67430
rect 6540 -64588 6640 -64526
rect 4316 -67430 4416 -67368
rect 6540 -67430 6640 -67368
rect 4316 -67530 4478 -67430
rect 6478 -67530 6640 -67430
rect -27684 -72766 -27522 -72666
rect -25522 -72766 -25360 -72666
rect -27684 -72828 -27584 -72766
rect -25460 -72828 -25360 -72766
rect -27684 -75670 -27584 -75608
rect -23684 -72766 -23522 -72666
rect -21522 -72766 -21360 -72666
rect -23684 -72828 -23584 -72766
rect -25460 -75670 -25360 -75608
rect -27684 -75770 -27522 -75670
rect -25522 -75770 -25360 -75670
rect -21460 -72828 -21360 -72766
rect -23684 -75670 -23584 -75608
rect -19684 -72766 -19522 -72666
rect -17522 -72766 -17360 -72666
rect -19684 -72828 -19584 -72766
rect -21460 -75670 -21360 -75608
rect -23684 -75770 -23522 -75670
rect -21522 -75770 -21360 -75670
rect -17460 -72828 -17360 -72766
rect -19684 -75670 -19584 -75608
rect -15684 -72766 -15522 -72666
rect -13522 -72766 -13360 -72666
rect -15684 -72828 -15584 -72766
rect -17460 -75670 -17360 -75608
rect -19684 -75770 -19522 -75670
rect -17522 -75770 -17360 -75670
rect -13460 -72828 -13360 -72766
rect -15684 -75670 -15584 -75608
rect -11684 -72766 -11522 -72666
rect -9522 -72766 -9360 -72666
rect -11684 -72828 -11584 -72766
rect -13460 -75670 -13360 -75608
rect -15684 -75770 -15522 -75670
rect -13522 -75770 -13360 -75670
rect -9460 -72828 -9360 -72766
rect -11684 -75670 -11584 -75608
rect -7684 -72766 -7522 -72666
rect -5522 -72766 -5360 -72666
rect -7684 -72828 -7584 -72766
rect -9460 -75670 -9360 -75608
rect -11684 -75770 -11522 -75670
rect -9522 -75770 -9360 -75670
rect -5460 -72828 -5360 -72766
rect -7684 -75670 -7584 -75608
rect -3684 -72766 -3522 -72666
rect -1522 -72766 -1360 -72666
rect -3684 -72828 -3584 -72766
rect -5460 -75670 -5360 -75608
rect -7684 -75770 -7522 -75670
rect -5522 -75770 -5360 -75670
rect -1460 -72828 -1360 -72766
rect -3684 -75670 -3584 -75608
rect 316 -72766 478 -72666
rect 2478 -72766 2640 -72666
rect 316 -72828 416 -72766
rect -1460 -75670 -1360 -75608
rect -3684 -75770 -3522 -75670
rect -1522 -75770 -1360 -75670
rect 2540 -72828 2640 -72766
rect 316 -75670 416 -75608
rect 4316 -72766 4478 -72666
rect 6478 -72766 6640 -72666
rect 4316 -72828 4416 -72766
rect 2540 -75670 2640 -75608
rect 316 -75770 478 -75670
rect 2478 -75770 2640 -75670
rect 6540 -72828 6640 -72766
rect 4316 -75670 4416 -75608
rect 6540 -75670 6640 -75608
rect 4316 -75770 4478 -75670
rect 6478 -75770 6640 -75670
<< psubdiffcont >>
rect 56532 -42446 57516 -42346
rect 55998 -42562 56186 -42528
rect 55902 -42918 55936 -42624
rect 56248 -42918 56282 -42624
rect 55998 -43014 56186 -42980
rect 56370 -43070 56470 -42508
rect 13284 -43256 50204 -43156
rect 10392 -57706 12010 -57672
rect 10296 -58124 10330 -57768
rect 12072 -58124 12106 -57768
rect 10392 -58220 12010 -58186
rect 13122 -59038 13222 -43318
rect 28554 -43796 28588 -43762
rect 29572 -43796 29606 -43762
rect 30590 -43796 30624 -43762
rect 31608 -43796 31642 -43762
rect 32626 -43796 32660 -43762
rect 33644 -43796 33678 -43762
rect 34662 -43796 34696 -43762
rect 35680 -43796 35714 -43762
rect 36698 -43796 36732 -43762
rect 37716 -43796 37750 -43762
rect 38734 -43796 38768 -43762
rect 39752 -43796 39786 -43762
rect 40770 -43796 40804 -43762
rect 41788 -43796 41822 -43762
rect 42806 -43796 42840 -43762
rect 43824 -43796 43858 -43762
rect 44842 -43796 44876 -43762
rect 45860 -43796 45894 -43762
rect 46878 -43796 46912 -43762
rect 47896 -43796 47930 -43762
rect 16260 -44398 16294 -44364
rect 17278 -44398 17312 -44364
rect 18296 -44398 18330 -44364
rect 19314 -44398 19348 -44364
rect 20332 -44398 20366 -44364
rect 21350 -44398 21384 -44364
rect 22368 -44398 22402 -44364
rect 23386 -44398 23420 -44364
rect 24404 -44398 24438 -44364
rect 25432 -44398 25466 -44364
rect 16260 -45216 16294 -45182
rect 17278 -45216 17312 -45182
rect 18296 -45216 18330 -45182
rect 19314 -45216 19348 -45182
rect 20332 -45216 20366 -45182
rect 21350 -45216 21384 -45182
rect 22368 -45216 22402 -45182
rect 23386 -45216 23420 -45182
rect 24404 -45216 24438 -45182
rect 25432 -45216 25466 -45182
rect 28566 -45822 28600 -45788
rect 29584 -45822 29618 -45788
rect 30602 -45822 30636 -45788
rect 31620 -45822 31654 -45788
rect 32638 -45822 32672 -45788
rect 33656 -45822 33690 -45788
rect 34674 -45822 34708 -45788
rect 35692 -45822 35726 -45788
rect 36710 -45822 36744 -45788
rect 37728 -45822 37762 -45788
rect 38746 -45822 38780 -45788
rect 39764 -45822 39798 -45788
rect 40782 -45822 40816 -45788
rect 41800 -45822 41834 -45788
rect 42818 -45822 42852 -45788
rect 43836 -45822 43870 -45788
rect 44854 -45822 44888 -45788
rect 45872 -45822 45906 -45788
rect 46890 -45822 46924 -45788
rect 47908 -45822 47942 -45788
rect 16260 -46034 16294 -46000
rect 17278 -46034 17312 -46000
rect 18296 -46034 18330 -46000
rect 19314 -46034 19348 -46000
rect 20332 -46034 20366 -46000
rect 21350 -46034 21384 -46000
rect 22368 -46034 22402 -46000
rect 23386 -46034 23420 -46000
rect 24404 -46034 24438 -46000
rect 25432 -46034 25466 -46000
rect 16260 -46852 16294 -46818
rect 17278 -46852 17312 -46818
rect 18296 -46852 18330 -46818
rect 19314 -46852 19348 -46818
rect 20332 -46852 20366 -46818
rect 21350 -46852 21384 -46818
rect 22368 -46852 22402 -46818
rect 23386 -46852 23420 -46818
rect 24404 -46852 24438 -46818
rect 25432 -46852 25466 -46818
rect 28554 -47128 28588 -47094
rect 29572 -47128 29606 -47094
rect 30590 -47128 30624 -47094
rect 31608 -47128 31642 -47094
rect 32626 -47128 32660 -47094
rect 33644 -47128 33678 -47094
rect 34662 -47128 34696 -47094
rect 35680 -47128 35714 -47094
rect 36698 -47128 36732 -47094
rect 37716 -47128 37750 -47094
rect 38734 -47128 38768 -47094
rect 39752 -47128 39786 -47094
rect 40770 -47128 40804 -47094
rect 41788 -47128 41822 -47094
rect 42806 -47128 42840 -47094
rect 43824 -47128 43858 -47094
rect 44842 -47128 44876 -47094
rect 45860 -47128 45894 -47094
rect 46878 -47128 46912 -47094
rect 47896 -47128 47930 -47094
rect 16260 -47670 16294 -47636
rect 17278 -47670 17312 -47636
rect 18296 -47670 18330 -47636
rect 19314 -47670 19348 -47636
rect 20332 -47670 20366 -47636
rect 21350 -47670 21384 -47636
rect 22368 -47670 22402 -47636
rect 23386 -47670 23420 -47636
rect 24404 -47670 24438 -47636
rect 25432 -47670 25466 -47636
rect 16260 -48488 16294 -48454
rect 17278 -48488 17312 -48454
rect 18296 -48488 18330 -48454
rect 19314 -48488 19348 -48454
rect 20332 -48488 20366 -48454
rect 21350 -48488 21384 -48454
rect 22368 -48488 22402 -48454
rect 28542 -48364 28576 -48330
rect 29560 -48364 29594 -48330
rect 30578 -48364 30612 -48330
rect 31596 -48364 31630 -48330
rect 32614 -48364 32648 -48330
rect 33632 -48364 33666 -48330
rect 34650 -48364 34684 -48330
rect 35668 -48364 35702 -48330
rect 36686 -48364 36720 -48330
rect 37704 -48364 37738 -48330
rect 38722 -48364 38756 -48330
rect 39740 -48364 39774 -48330
rect 40758 -48364 40792 -48330
rect 41776 -48364 41810 -48330
rect 42794 -48364 42828 -48330
rect 43812 -48364 43846 -48330
rect 44830 -48364 44864 -48330
rect 45848 -48364 45882 -48330
rect 46866 -48364 46900 -48330
rect 47884 -48364 47918 -48330
rect 23386 -48488 23420 -48454
rect 24404 -48488 24438 -48454
rect 25432 -48488 25466 -48454
rect 16260 -49306 16294 -49272
rect 17278 -49306 17312 -49272
rect 18296 -49306 18330 -49272
rect 19314 -49306 19348 -49272
rect 20332 -49306 20366 -49272
rect 21350 -49306 21384 -49272
rect 22368 -49306 22402 -49272
rect 23386 -49306 23420 -49272
rect 24404 -49306 24438 -49272
rect 25432 -49306 25466 -49272
rect 28542 -49588 28576 -49554
rect 29560 -49588 29594 -49554
rect 30578 -49588 30612 -49554
rect 31596 -49588 31630 -49554
rect 32614 -49588 32648 -49554
rect 33632 -49588 33666 -49554
rect 34650 -49588 34684 -49554
rect 35668 -49588 35702 -49554
rect 36686 -49588 36720 -49554
rect 37704 -49588 37738 -49554
rect 38722 -49588 38756 -49554
rect 39740 -49588 39774 -49554
rect 40758 -49588 40792 -49554
rect 41776 -49588 41810 -49554
rect 42794 -49588 42828 -49554
rect 43812 -49588 43846 -49554
rect 44830 -49588 44864 -49554
rect 45848 -49588 45882 -49554
rect 46866 -49588 46900 -49554
rect 47884 -49588 47918 -49554
rect 16260 -50124 16294 -50090
rect 17278 -50124 17312 -50090
rect 18296 -50124 18330 -50090
rect 19314 -50124 19348 -50090
rect 20332 -50124 20366 -50090
rect 21350 -50124 21384 -50090
rect 22368 -50124 22402 -50090
rect 23386 -50124 23420 -50090
rect 24404 -50124 24438 -50090
rect 25432 -50124 25466 -50090
rect 28554 -50824 28588 -50790
rect 29572 -50824 29606 -50790
rect 30590 -50824 30624 -50790
rect 31608 -50824 31642 -50790
rect 32626 -50824 32660 -50790
rect 33644 -50824 33678 -50790
rect 34662 -50824 34696 -50790
rect 35680 -50824 35714 -50790
rect 36698 -50824 36732 -50790
rect 37716 -50824 37750 -50790
rect 38734 -50824 38768 -50790
rect 39752 -50824 39786 -50790
rect 40770 -50824 40804 -50790
rect 41788 -50824 41822 -50790
rect 42806 -50824 42840 -50790
rect 43824 -50824 43858 -50790
rect 44842 -50824 44876 -50790
rect 45860 -50824 45894 -50790
rect 46878 -50824 46912 -50790
rect 47896 -50824 47930 -50790
rect 16248 -51018 16282 -50984
rect 17266 -51018 17300 -50984
rect 18284 -51018 18318 -50984
rect 19302 -51018 19336 -50984
rect 20320 -51018 20354 -50984
rect 21338 -51018 21372 -50984
rect 22356 -51018 22390 -50984
rect 23374 -51018 23408 -50984
rect 24392 -51018 24426 -50984
rect 25420 -51018 25454 -50984
rect 15452 -51966 15486 -51932
rect 16470 -51966 16504 -51932
rect 17488 -51966 17522 -51932
rect 18506 -51966 18540 -51932
rect 19524 -51966 19558 -51932
rect 20542 -51966 20576 -51932
rect 21560 -51966 21594 -51932
rect 22578 -51966 22612 -51932
rect 23596 -51966 23630 -51932
rect 24614 -51966 24648 -51932
rect 25632 -51966 25666 -51932
rect 28554 -52072 28588 -52038
rect 29572 -52072 29606 -52038
rect 30590 -52072 30624 -52038
rect 31608 -52072 31642 -52038
rect 32626 -52072 32660 -52038
rect 33644 -52072 33678 -52038
rect 34662 -52072 34696 -52038
rect 35680 -52072 35714 -52038
rect 36698 -52072 36732 -52038
rect 37716 -52072 37750 -52038
rect 38734 -52072 38768 -52038
rect 39752 -52072 39786 -52038
rect 40770 -52072 40804 -52038
rect 41788 -52072 41822 -52038
rect 42806 -52072 42840 -52038
rect 43824 -52072 43858 -52038
rect 44842 -52072 44876 -52038
rect 45860 -52072 45894 -52038
rect 46878 -52072 46912 -52038
rect 47896 -52072 47930 -52038
rect 15464 -53108 15498 -53074
rect 16482 -53108 16516 -53074
rect 17500 -53108 17534 -53074
rect 18518 -53108 18552 -53074
rect 19536 -53108 19570 -53074
rect 20554 -53108 20588 -53074
rect 21572 -53108 21606 -53074
rect 22590 -53108 22624 -53074
rect 23608 -53108 23642 -53074
rect 24626 -53108 24660 -53074
rect 25644 -53108 25678 -53074
rect 28530 -53308 28564 -53274
rect 29548 -53308 29582 -53274
rect 30566 -53308 30600 -53274
rect 31584 -53308 31618 -53274
rect 32602 -53308 32636 -53274
rect 33620 -53308 33654 -53274
rect 34638 -53308 34672 -53274
rect 35656 -53308 35690 -53274
rect 36674 -53308 36708 -53274
rect 37692 -53308 37726 -53274
rect 38710 -53308 38744 -53274
rect 39728 -53308 39762 -53274
rect 40746 -53308 40780 -53274
rect 41764 -53308 41798 -53274
rect 42782 -53308 42816 -53274
rect 43800 -53308 43834 -53274
rect 44818 -53308 44852 -53274
rect 45836 -53308 45870 -53274
rect 46854 -53308 46888 -53274
rect 47872 -53308 47906 -53274
rect 15442 -54216 15476 -54182
rect 16460 -54216 16494 -54182
rect 17478 -54216 17512 -54182
rect 18496 -54216 18530 -54182
rect 19514 -54216 19548 -54182
rect 20532 -54216 20566 -54182
rect 21550 -54216 21584 -54182
rect 22568 -54216 22602 -54182
rect 23586 -54216 23620 -54182
rect 24604 -54216 24638 -54182
rect 25622 -54216 25656 -54182
rect 28542 -54532 28576 -54498
rect 29560 -54532 29594 -54498
rect 30578 -54532 30612 -54498
rect 31596 -54532 31630 -54498
rect 32614 -54532 32648 -54498
rect 33632 -54532 33666 -54498
rect 34650 -54532 34684 -54498
rect 35668 -54532 35702 -54498
rect 36686 -54532 36720 -54498
rect 37704 -54532 37738 -54498
rect 38722 -54532 38756 -54498
rect 39740 -54532 39774 -54498
rect 40758 -54532 40792 -54498
rect 41776 -54532 41810 -54498
rect 42794 -54532 42828 -54498
rect 43812 -54532 43846 -54498
rect 44830 -54532 44864 -54498
rect 45848 -54532 45882 -54498
rect 46866 -54532 46900 -54498
rect 47884 -54532 47918 -54498
rect 15442 -55322 15476 -55288
rect 16460 -55322 16494 -55288
rect 17478 -55322 17512 -55288
rect 18496 -55322 18530 -55288
rect 19514 -55322 19548 -55288
rect 20532 -55322 20566 -55288
rect 21550 -55322 21584 -55288
rect 22568 -55322 22602 -55288
rect 23586 -55322 23620 -55288
rect 24604 -55322 24638 -55288
rect 25622 -55322 25656 -55288
rect 28542 -55768 28576 -55734
rect 29560 -55768 29594 -55734
rect 30578 -55768 30612 -55734
rect 31596 -55768 31630 -55734
rect 32614 -55768 32648 -55734
rect 33632 -55768 33666 -55734
rect 34650 -55768 34684 -55734
rect 35668 -55768 35702 -55734
rect 36686 -55768 36720 -55734
rect 37704 -55768 37738 -55734
rect 38722 -55768 38756 -55734
rect 39740 -55768 39774 -55734
rect 40758 -55768 40792 -55734
rect 41776 -55768 41810 -55734
rect 42794 -55768 42828 -55734
rect 43812 -55768 43846 -55734
rect 44830 -55768 44864 -55734
rect 45848 -55768 45882 -55734
rect 46866 -55768 46900 -55734
rect 47884 -55768 47918 -55734
rect 15442 -56664 15476 -56630
rect 16460 -56664 16494 -56630
rect 17478 -56664 17512 -56630
rect 18496 -56664 18530 -56630
rect 19514 -56664 19548 -56630
rect 20532 -56664 20566 -56630
rect 21550 -56664 21584 -56630
rect 22568 -56664 22602 -56630
rect 23586 -56664 23620 -56630
rect 24604 -56664 24638 -56630
rect 25622 -56664 25656 -56630
rect 28554 -57014 28588 -56980
rect 29572 -57014 29606 -56980
rect 30590 -57014 30624 -56980
rect 31608 -57014 31642 -56980
rect 32626 -57014 32660 -56980
rect 33644 -57014 33678 -56980
rect 34662 -57014 34696 -56980
rect 35680 -57014 35714 -56980
rect 36698 -57014 36732 -56980
rect 37716 -57014 37750 -56980
rect 38734 -57014 38768 -56980
rect 39752 -57014 39786 -56980
rect 40770 -57014 40804 -56980
rect 41788 -57014 41822 -56980
rect 42806 -57014 42840 -56980
rect 43824 -57014 43858 -56980
rect 44842 -57014 44876 -56980
rect 45860 -57014 45894 -56980
rect 46878 -57014 46912 -56980
rect 47896 -57014 47930 -56980
rect 15252 -58110 15286 -58076
rect 16270 -58110 16304 -58076
rect 17288 -58110 17322 -58076
rect 18306 -58110 18340 -58076
rect 19324 -58110 19358 -58076
rect 20342 -58110 20376 -58076
rect 21360 -58110 21394 -58076
rect 22378 -58110 22412 -58076
rect 23396 -58110 23430 -58076
rect 24414 -58110 24448 -58076
rect 25432 -58110 25466 -58076
rect 28542 -58192 28576 -58158
rect 29560 -58192 29594 -58158
rect 30578 -58192 30612 -58158
rect 31596 -58192 31630 -58158
rect 32614 -58192 32648 -58158
rect 33632 -58192 33666 -58158
rect 34650 -58192 34684 -58158
rect 35668 -58192 35702 -58158
rect 36686 -58192 36720 -58158
rect 37704 -58192 37738 -58158
rect 38722 -58192 38756 -58158
rect 39740 -58192 39774 -58158
rect 40758 -58192 40792 -58158
rect 41776 -58192 41810 -58158
rect 42794 -58192 42828 -58158
rect 43812 -58192 43846 -58158
rect 44830 -58192 44864 -58158
rect 45848 -58192 45882 -58158
rect 46866 -58192 46900 -58158
rect 47884 -58192 47918 -58158
rect 50266 -59038 50366 -43318
rect 57628 -43144 57728 -42510
rect 57902 -42562 58090 -42528
rect 57806 -42918 57840 -42624
rect 58152 -42918 58186 -42624
rect 57902 -43014 58090 -42980
rect 56526 -43704 57510 -43604
rect 13284 -59200 50204 -59100
rect -27522 -67866 -25522 -67766
rect -27684 -69648 -27584 -67928
rect -25460 -69648 -25360 -67928
rect -27522 -69810 -25522 -69710
rect -23522 -67866 -21522 -67766
rect -23684 -69648 -23584 -67928
rect -21460 -69648 -21360 -67928
rect -23522 -69810 -21522 -69710
rect -19522 -67866 -17522 -67766
rect -19684 -69648 -19584 -67928
rect -17460 -69648 -17360 -67928
rect -19522 -69810 -17522 -69710
rect -15522 -67866 -13522 -67766
rect -15684 -69648 -15584 -67928
rect -13460 -69648 -13360 -67928
rect -15522 -69810 -13522 -69710
rect -11522 -67866 -9522 -67766
rect -11684 -69648 -11584 -67928
rect -9460 -69648 -9360 -67928
rect -11522 -69810 -9522 -69710
rect -7522 -67866 -5522 -67766
rect -7684 -69648 -7584 -67928
rect -5460 -69648 -5360 -67928
rect -7522 -69810 -5522 -69710
rect -3522 -67866 -1522 -67766
rect -3684 -69648 -3584 -67928
rect -1460 -69648 -1360 -67928
rect -3522 -69810 -1522 -69710
rect 478 -67866 2478 -67766
rect 316 -69648 416 -67928
rect 2540 -69648 2640 -67928
rect 478 -69810 2478 -69710
rect 4478 -67866 6478 -67766
rect 4316 -69648 4416 -67928
rect 6540 -69648 6640 -67928
rect 4478 -69810 6478 -69710
rect -27522 -70486 -25522 -70386
rect -27684 -72268 -27584 -70548
rect -25460 -72268 -25360 -70548
rect -27522 -72430 -25522 -72330
rect -23522 -70486 -21522 -70386
rect -23684 -72268 -23584 -70548
rect -21460 -72268 -21360 -70548
rect -23522 -72430 -21522 -72330
rect -19522 -70486 -17522 -70386
rect -19684 -72268 -19584 -70548
rect -17460 -72268 -17360 -70548
rect -19522 -72430 -17522 -72330
rect -15522 -70486 -13522 -70386
rect -15684 -72268 -15584 -70548
rect -13460 -72268 -13360 -70548
rect -15522 -72430 -13522 -72330
rect -11522 -70486 -9522 -70386
rect -11684 -72268 -11584 -70548
rect -9460 -72268 -9360 -70548
rect -11522 -72430 -9522 -72330
rect -7522 -70486 -5522 -70386
rect -7684 -72268 -7584 -70548
rect -5460 -72268 -5360 -70548
rect -7522 -72430 -5522 -72330
rect -3522 -70486 -1522 -70386
rect -3684 -72268 -3584 -70548
rect -1460 -72268 -1360 -70548
rect -3522 -72430 -1522 -72330
rect 478 -70486 2478 -70386
rect 316 -72268 416 -70548
rect 2540 -72268 2640 -70548
rect 478 -72430 2478 -72330
rect 4478 -70486 6478 -70386
rect 4316 -72268 4416 -70548
rect 6540 -72268 6640 -70548
rect 4478 -72430 6478 -72330
<< nsubdiffcont >>
rect 25984 -27756 50104 -27656
rect 25822 -42164 25922 -27818
rect 32440 -30234 32474 -30200
rect 33458 -30234 33492 -30200
rect 34476 -30234 34510 -30200
rect 35494 -30234 35528 -30200
rect 36512 -30234 36546 -30200
rect 37530 -30234 37564 -30200
rect 38548 -30234 38582 -30200
rect 39566 -30234 39600 -30200
rect 40584 -30234 40618 -30200
rect 41602 -30234 41636 -30200
rect 42620 -30234 42654 -30200
rect 43638 -30234 43672 -30200
rect 44656 -30234 44690 -30200
rect 45674 -30234 45708 -30200
rect 46692 -30234 46726 -30200
rect 47710 -30234 47744 -30200
rect 32462 -31388 32496 -31354
rect 33480 -31388 33514 -31354
rect 34498 -31388 34532 -31354
rect 35516 -31388 35550 -31354
rect 36534 -31388 36568 -31354
rect 37552 -31388 37586 -31354
rect 38570 -31388 38604 -31354
rect 39588 -31388 39622 -31354
rect 40606 -31388 40640 -31354
rect 41624 -31388 41658 -31354
rect 42642 -31388 42676 -31354
rect 43660 -31388 43694 -31354
rect 44678 -31388 44712 -31354
rect 45696 -31388 45730 -31354
rect 46714 -31388 46748 -31354
rect 47732 -31388 47766 -31354
rect 32440 -32520 32474 -32486
rect 33458 -32520 33492 -32486
rect 34476 -32520 34510 -32486
rect 35494 -32520 35528 -32486
rect 36512 -32520 36546 -32486
rect 37530 -32520 37564 -32486
rect 38548 -32520 38582 -32486
rect 39566 -32520 39600 -32486
rect 40584 -32520 40618 -32486
rect 41602 -32520 41636 -32486
rect 42620 -32520 42654 -32486
rect 43638 -32520 43672 -32486
rect 44656 -32520 44690 -32486
rect 45674 -32520 45708 -32486
rect 46692 -32520 46726 -32486
rect 47710 -32520 47744 -32486
rect 32440 -33902 32474 -33868
rect 33458 -33902 33492 -33868
rect 34476 -33902 34510 -33868
rect 35494 -33902 35528 -33868
rect 36512 -33902 36546 -33868
rect 37530 -33902 37564 -33868
rect 38548 -33902 38582 -33868
rect 39566 -33902 39600 -33868
rect 40584 -33902 40618 -33868
rect 41602 -33902 41636 -33868
rect 42620 -33902 42654 -33868
rect 43638 -33902 43672 -33868
rect 44656 -33902 44690 -33868
rect 45674 -33902 45708 -33868
rect 46692 -33902 46726 -33868
rect 47710 -33902 47744 -33868
rect 33128 -35250 33162 -35216
rect 34146 -35250 34180 -35216
rect 35164 -35250 35198 -35216
rect 36182 -35250 36216 -35216
rect 37200 -35250 37234 -35216
rect 38218 -35250 38252 -35216
rect 39236 -35250 39270 -35216
rect 40254 -35250 40288 -35216
rect 41272 -35250 41306 -35216
rect 42290 -35250 42324 -35216
rect 43308 -35250 43342 -35216
rect 44326 -35250 44360 -35216
rect 45344 -35250 45378 -35216
rect 46362 -35250 46396 -35216
rect 47380 -35250 47414 -35216
rect 32734 -36528 32768 -36494
rect 33752 -36528 33786 -36494
rect 34770 -36528 34804 -36494
rect 35788 -36528 35822 -36494
rect 36806 -36528 36840 -36494
rect 37824 -36528 37858 -36494
rect 38842 -36528 38876 -36494
rect 39860 -36528 39894 -36494
rect 40878 -36528 40912 -36494
rect 41896 -36528 41930 -36494
rect 42914 -36528 42948 -36494
rect 43932 -36528 43966 -36494
rect 44950 -36528 44984 -36494
rect 45968 -36528 46002 -36494
rect 46986 -36528 47020 -36494
rect 48004 -36528 48038 -36494
rect 28136 -36838 28170 -36804
rect 29154 -36838 29188 -36804
rect 30172 -36838 30206 -36804
rect 31190 -36838 31224 -36804
rect 27612 -37992 27646 -37958
rect 28630 -37992 28664 -37958
rect 29648 -37992 29682 -37958
rect 30666 -37992 30700 -37958
rect 32824 -37976 32858 -37942
rect 33842 -37976 33876 -37942
rect 34860 -37976 34894 -37942
rect 35878 -37976 35912 -37942
rect 36896 -37976 36930 -37942
rect 37914 -37976 37948 -37942
rect 38932 -37976 38966 -37942
rect 39950 -37976 39984 -37942
rect 40968 -37976 41002 -37942
rect 41986 -37976 42020 -37942
rect 43004 -37976 43038 -37942
rect 44022 -37976 44056 -37942
rect 45040 -37976 45074 -37942
rect 46058 -37976 46092 -37942
rect 47076 -37976 47110 -37942
rect 48094 -37976 48128 -37942
rect 27622 -39020 27656 -38986
rect 28640 -39020 28674 -38986
rect 29658 -39020 29692 -38986
rect 30676 -39020 30710 -38986
rect 32848 -39244 32882 -39210
rect 33866 -39244 33900 -39210
rect 34884 -39244 34918 -39210
rect 35902 -39244 35936 -39210
rect 36920 -39244 36954 -39210
rect 37938 -39244 37972 -39210
rect 38956 -39244 38990 -39210
rect 39974 -39244 40008 -39210
rect 40992 -39244 41026 -39210
rect 42010 -39244 42044 -39210
rect 43028 -39244 43062 -39210
rect 44046 -39244 44080 -39210
rect 45064 -39244 45098 -39210
rect 46082 -39244 46116 -39210
rect 47100 -39244 47134 -39210
rect 48118 -39244 48152 -39210
rect 27612 -40048 27646 -40014
rect 28630 -40048 28664 -40014
rect 29648 -40048 29682 -40014
rect 30666 -40048 30700 -40014
rect 32712 -40488 32746 -40454
rect 33730 -40488 33764 -40454
rect 34748 -40488 34782 -40454
rect 35766 -40488 35800 -40454
rect 36784 -40488 36818 -40454
rect 37802 -40488 37836 -40454
rect 38820 -40488 38854 -40454
rect 39838 -40488 39872 -40454
rect 40856 -40488 40890 -40454
rect 41874 -40488 41908 -40454
rect 42892 -40488 42926 -40454
rect 43910 -40488 43944 -40454
rect 44928 -40488 44962 -40454
rect 45946 -40488 45980 -40454
rect 46964 -40488 46998 -40454
rect 47982 -40488 48016 -40454
rect 28136 -41200 28170 -41166
rect 29154 -41200 29188 -41166
rect 30172 -41200 30206 -41166
rect 31190 -41200 31224 -41166
rect 50166 -42164 50266 -27818
rect 25984 -42326 50104 -42226
rect 52318 -39080 55358 -38980
rect 52156 -42162 52256 -39142
rect 55420 -42162 55520 -39142
rect 56020 -39080 58100 -38980
rect 55858 -41368 55958 -39142
rect 58162 -41368 58262 -39142
rect 56020 -41530 58100 -41430
rect 52318 -42324 55358 -42224
rect 54200 -42418 55422 -42384
rect 54104 -42810 54138 -42578
rect 55484 -42810 55518 -42578
rect 54200 -43000 55422 -42966
rect 10392 -56773 12010 -56739
rect 10296 -57409 10330 -56835
rect 12072 -57409 12106 -56835
rect 10392 -57505 12010 -57471
rect -27522 -64526 -25522 -64426
rect -27684 -67368 -27584 -64588
rect -25460 -67368 -25360 -64588
rect -23522 -64526 -21522 -64426
rect -27522 -67530 -25522 -67430
rect -23684 -67368 -23584 -64588
rect -21460 -67368 -21360 -64588
rect -19522 -64526 -17522 -64426
rect -23522 -67530 -21522 -67430
rect -19684 -67368 -19584 -64588
rect -17460 -67368 -17360 -64588
rect -15522 -64526 -13522 -64426
rect -19522 -67530 -17522 -67430
rect -15684 -67368 -15584 -64588
rect -13460 -67368 -13360 -64588
rect -11522 -64526 -9522 -64426
rect -15522 -67530 -13522 -67430
rect -11684 -67368 -11584 -64588
rect -9460 -67368 -9360 -64588
rect -7522 -64526 -5522 -64426
rect -11522 -67530 -9522 -67430
rect -7684 -67368 -7584 -64588
rect -5460 -67368 -5360 -64588
rect -3522 -64526 -1522 -64426
rect -7522 -67530 -5522 -67430
rect -3684 -67368 -3584 -64588
rect -1460 -67368 -1360 -64588
rect 478 -64526 2478 -64426
rect -3522 -67530 -1522 -67430
rect 316 -67368 416 -64588
rect 2540 -67368 2640 -64588
rect 4478 -64526 6478 -64426
rect 478 -67530 2478 -67430
rect 4316 -67368 4416 -64588
rect 6540 -67368 6640 -64588
rect 4478 -67530 6478 -67430
rect -27522 -72766 -25522 -72666
rect -27684 -75608 -27584 -72828
rect -25460 -75608 -25360 -72828
rect -23522 -72766 -21522 -72666
rect -27522 -75770 -25522 -75670
rect -23684 -75608 -23584 -72828
rect -21460 -75608 -21360 -72828
rect -19522 -72766 -17522 -72666
rect -23522 -75770 -21522 -75670
rect -19684 -75608 -19584 -72828
rect -17460 -75608 -17360 -72828
rect -15522 -72766 -13522 -72666
rect -19522 -75770 -17522 -75670
rect -15684 -75608 -15584 -72828
rect -13460 -75608 -13360 -72828
rect -11522 -72766 -9522 -72666
rect -15522 -75770 -13522 -75670
rect -11684 -75608 -11584 -72828
rect -9460 -75608 -9360 -72828
rect -7522 -72766 -5522 -72666
rect -11522 -75770 -9522 -75670
rect -7684 -75608 -7584 -72828
rect -5460 -75608 -5360 -72828
rect -3522 -72766 -1522 -72666
rect -7522 -75770 -5522 -75670
rect -3684 -75608 -3584 -72828
rect -1460 -75608 -1360 -72828
rect 478 -72766 2478 -72666
rect -3522 -75770 -1522 -75670
rect 316 -75608 416 -72828
rect 2540 -75608 2640 -72828
rect 4478 -72766 6478 -72666
rect 478 -75770 2478 -75670
rect 4316 -75608 4416 -72828
rect 6540 -75608 6640 -72828
rect 4478 -75770 6478 -75670
<< poly >>
rect 32164 -30423 32752 -30407
rect 32164 -30440 32180 -30423
rect 31978 -30457 32180 -30440
rect 32736 -30440 32752 -30423
rect 33182 -30423 33770 -30407
rect 33182 -30440 33198 -30423
rect 32736 -30457 32938 -30440
rect 31978 -30504 32938 -30457
rect 32996 -30457 33198 -30440
rect 33754 -30440 33770 -30423
rect 34200 -30423 34788 -30407
rect 34200 -30440 34216 -30423
rect 33754 -30457 33956 -30440
rect 32996 -30504 33956 -30457
rect 34014 -30457 34216 -30440
rect 34772 -30440 34788 -30423
rect 35218 -30423 35806 -30407
rect 35218 -30440 35234 -30423
rect 34772 -30457 34974 -30440
rect 34014 -30504 34974 -30457
rect 35032 -30457 35234 -30440
rect 35790 -30440 35806 -30423
rect 36236 -30423 36824 -30407
rect 36236 -30440 36252 -30423
rect 35790 -30457 35992 -30440
rect 35032 -30504 35992 -30457
rect 36050 -30457 36252 -30440
rect 36808 -30440 36824 -30423
rect 37254 -30423 37842 -30407
rect 37254 -30440 37270 -30423
rect 36808 -30457 37010 -30440
rect 36050 -30504 37010 -30457
rect 37068 -30457 37270 -30440
rect 37826 -30440 37842 -30423
rect 38272 -30423 38860 -30407
rect 38272 -30440 38288 -30423
rect 37826 -30457 38028 -30440
rect 37068 -30504 38028 -30457
rect 38086 -30457 38288 -30440
rect 38844 -30440 38860 -30423
rect 39290 -30423 39878 -30407
rect 39290 -30440 39306 -30423
rect 38844 -30457 39046 -30440
rect 38086 -30504 39046 -30457
rect 39104 -30457 39306 -30440
rect 39862 -30440 39878 -30423
rect 40308 -30423 40896 -30407
rect 40308 -30440 40324 -30423
rect 39862 -30457 40064 -30440
rect 39104 -30504 40064 -30457
rect 40122 -30457 40324 -30440
rect 40880 -30440 40896 -30423
rect 41326 -30423 41914 -30407
rect 41326 -30440 41342 -30423
rect 40880 -30457 41082 -30440
rect 40122 -30504 41082 -30457
rect 41140 -30457 41342 -30440
rect 41898 -30440 41914 -30423
rect 42344 -30423 42932 -30407
rect 42344 -30440 42360 -30423
rect 41898 -30457 42100 -30440
rect 41140 -30504 42100 -30457
rect 42158 -30457 42360 -30440
rect 42916 -30440 42932 -30423
rect 43362 -30423 43950 -30407
rect 43362 -30440 43378 -30423
rect 42916 -30457 43118 -30440
rect 42158 -30504 43118 -30457
rect 43176 -30457 43378 -30440
rect 43934 -30440 43950 -30423
rect 44380 -30423 44968 -30407
rect 44380 -30440 44396 -30423
rect 43934 -30457 44136 -30440
rect 43176 -30504 44136 -30457
rect 44194 -30457 44396 -30440
rect 44952 -30440 44968 -30423
rect 45398 -30423 45986 -30407
rect 45398 -30440 45414 -30423
rect 44952 -30457 45154 -30440
rect 44194 -30504 45154 -30457
rect 45212 -30457 45414 -30440
rect 45970 -30440 45986 -30423
rect 46416 -30423 47004 -30407
rect 46416 -30440 46432 -30423
rect 45970 -30457 46172 -30440
rect 45212 -30504 46172 -30457
rect 46230 -30457 46432 -30440
rect 46988 -30440 47004 -30423
rect 47434 -30423 48022 -30407
rect 47434 -30440 47450 -30423
rect 46988 -30457 47190 -30440
rect 46230 -30504 47190 -30457
rect 47248 -30457 47450 -30440
rect 48006 -30440 48022 -30423
rect 48006 -30457 48208 -30440
rect 47248 -30504 48208 -30457
rect 31978 -31151 32938 -31104
rect 31978 -31168 32180 -31151
rect 32164 -31185 32180 -31168
rect 32736 -31168 32938 -31151
rect 32996 -31151 33956 -31104
rect 32996 -31168 33198 -31151
rect 32736 -31185 32752 -31168
rect 32164 -31201 32752 -31185
rect 33182 -31185 33198 -31168
rect 33754 -31168 33956 -31151
rect 34014 -31151 34974 -31104
rect 34014 -31168 34216 -31151
rect 33754 -31185 33770 -31168
rect 33182 -31201 33770 -31185
rect 34200 -31185 34216 -31168
rect 34772 -31168 34974 -31151
rect 35032 -31151 35992 -31104
rect 35032 -31168 35234 -31151
rect 34772 -31185 34788 -31168
rect 34200 -31201 34788 -31185
rect 35218 -31185 35234 -31168
rect 35790 -31168 35992 -31151
rect 36050 -31151 37010 -31104
rect 36050 -31168 36252 -31151
rect 35790 -31185 35806 -31168
rect 35218 -31201 35806 -31185
rect 36236 -31185 36252 -31168
rect 36808 -31168 37010 -31151
rect 37068 -31151 38028 -31104
rect 37068 -31168 37270 -31151
rect 36808 -31185 36824 -31168
rect 36236 -31201 36824 -31185
rect 37254 -31185 37270 -31168
rect 37826 -31168 38028 -31151
rect 38086 -31151 39046 -31104
rect 38086 -31168 38288 -31151
rect 37826 -31185 37842 -31168
rect 37254 -31201 37842 -31185
rect 38272 -31185 38288 -31168
rect 38844 -31168 39046 -31151
rect 39104 -31151 40064 -31104
rect 39104 -31168 39306 -31151
rect 38844 -31185 38860 -31168
rect 38272 -31201 38860 -31185
rect 39290 -31185 39306 -31168
rect 39862 -31168 40064 -31151
rect 40122 -31151 41082 -31104
rect 40122 -31168 40324 -31151
rect 39862 -31185 39878 -31168
rect 39290 -31201 39878 -31185
rect 40308 -31185 40324 -31168
rect 40880 -31168 41082 -31151
rect 41140 -31151 42100 -31104
rect 41140 -31168 41342 -31151
rect 40880 -31185 40896 -31168
rect 40308 -31201 40896 -31185
rect 41326 -31185 41342 -31168
rect 41898 -31168 42100 -31151
rect 42158 -31151 43118 -31104
rect 42158 -31168 42360 -31151
rect 41898 -31185 41914 -31168
rect 41326 -31201 41914 -31185
rect 42344 -31185 42360 -31168
rect 42916 -31168 43118 -31151
rect 43176 -31151 44136 -31104
rect 43176 -31168 43378 -31151
rect 42916 -31185 42932 -31168
rect 42344 -31201 42932 -31185
rect 43362 -31185 43378 -31168
rect 43934 -31168 44136 -31151
rect 44194 -31151 45154 -31104
rect 44194 -31168 44396 -31151
rect 43934 -31185 43950 -31168
rect 43362 -31201 43950 -31185
rect 44380 -31185 44396 -31168
rect 44952 -31168 45154 -31151
rect 45212 -31151 46172 -31104
rect 45212 -31168 45414 -31151
rect 44952 -31185 44968 -31168
rect 44380 -31201 44968 -31185
rect 45398 -31185 45414 -31168
rect 45970 -31168 46172 -31151
rect 46230 -31151 47190 -31104
rect 46230 -31168 46432 -31151
rect 45970 -31185 45986 -31168
rect 45398 -31201 45986 -31185
rect 46416 -31185 46432 -31168
rect 46988 -31168 47190 -31151
rect 47248 -31151 48208 -31104
rect 47248 -31168 47450 -31151
rect 46988 -31185 47004 -31168
rect 46416 -31201 47004 -31185
rect 47434 -31185 47450 -31168
rect 48006 -31168 48208 -31151
rect 48006 -31185 48022 -31168
rect 47434 -31201 48022 -31185
rect 32164 -31559 32752 -31543
rect 32164 -31576 32180 -31559
rect 31978 -31593 32180 -31576
rect 32736 -31576 32752 -31559
rect 33182 -31559 33770 -31543
rect 33182 -31576 33198 -31559
rect 32736 -31593 32938 -31576
rect 31978 -31640 32938 -31593
rect 32996 -31593 33198 -31576
rect 33754 -31576 33770 -31559
rect 34200 -31559 34788 -31543
rect 34200 -31576 34216 -31559
rect 33754 -31593 33956 -31576
rect 32996 -31640 33956 -31593
rect 34014 -31593 34216 -31576
rect 34772 -31576 34788 -31559
rect 35218 -31559 35806 -31543
rect 35218 -31576 35234 -31559
rect 34772 -31593 34974 -31576
rect 34014 -31640 34974 -31593
rect 35032 -31593 35234 -31576
rect 35790 -31576 35806 -31559
rect 36236 -31559 36824 -31543
rect 36236 -31576 36252 -31559
rect 35790 -31593 35992 -31576
rect 35032 -31640 35992 -31593
rect 36050 -31593 36252 -31576
rect 36808 -31576 36824 -31559
rect 37254 -31559 37842 -31543
rect 37254 -31576 37270 -31559
rect 36808 -31593 37010 -31576
rect 36050 -31640 37010 -31593
rect 37068 -31593 37270 -31576
rect 37826 -31576 37842 -31559
rect 38272 -31559 38860 -31543
rect 38272 -31576 38288 -31559
rect 37826 -31593 38028 -31576
rect 37068 -31640 38028 -31593
rect 38086 -31593 38288 -31576
rect 38844 -31576 38860 -31559
rect 39290 -31559 39878 -31543
rect 39290 -31576 39306 -31559
rect 38844 -31593 39046 -31576
rect 38086 -31640 39046 -31593
rect 39104 -31593 39306 -31576
rect 39862 -31576 39878 -31559
rect 40308 -31559 40896 -31543
rect 40308 -31576 40324 -31559
rect 39862 -31593 40064 -31576
rect 39104 -31640 40064 -31593
rect 40122 -31593 40324 -31576
rect 40880 -31576 40896 -31559
rect 41326 -31559 41914 -31543
rect 41326 -31576 41342 -31559
rect 40880 -31593 41082 -31576
rect 40122 -31640 41082 -31593
rect 41140 -31593 41342 -31576
rect 41898 -31576 41914 -31559
rect 42344 -31559 42932 -31543
rect 42344 -31576 42360 -31559
rect 41898 -31593 42100 -31576
rect 41140 -31640 42100 -31593
rect 42158 -31593 42360 -31576
rect 42916 -31576 42932 -31559
rect 43362 -31559 43950 -31543
rect 43362 -31576 43378 -31559
rect 42916 -31593 43118 -31576
rect 42158 -31640 43118 -31593
rect 43176 -31593 43378 -31576
rect 43934 -31576 43950 -31559
rect 44380 -31559 44968 -31543
rect 44380 -31576 44396 -31559
rect 43934 -31593 44136 -31576
rect 43176 -31640 44136 -31593
rect 44194 -31593 44396 -31576
rect 44952 -31576 44968 -31559
rect 45398 -31559 45986 -31543
rect 45398 -31576 45414 -31559
rect 44952 -31593 45154 -31576
rect 44194 -31640 45154 -31593
rect 45212 -31593 45414 -31576
rect 45970 -31576 45986 -31559
rect 46416 -31559 47004 -31543
rect 46416 -31576 46432 -31559
rect 45970 -31593 46172 -31576
rect 45212 -31640 46172 -31593
rect 46230 -31593 46432 -31576
rect 46988 -31576 47004 -31559
rect 47434 -31559 48022 -31543
rect 47434 -31576 47450 -31559
rect 46988 -31593 47190 -31576
rect 46230 -31640 47190 -31593
rect 47248 -31593 47450 -31576
rect 48006 -31576 48022 -31559
rect 48006 -31593 48208 -31576
rect 47248 -31640 48208 -31593
rect 31978 -32287 32938 -32240
rect 31978 -32304 32180 -32287
rect 32164 -32321 32180 -32304
rect 32736 -32304 32938 -32287
rect 32996 -32287 33956 -32240
rect 32996 -32304 33198 -32287
rect 32736 -32321 32752 -32304
rect 32164 -32337 32752 -32321
rect 33182 -32321 33198 -32304
rect 33754 -32304 33956 -32287
rect 34014 -32287 34974 -32240
rect 34014 -32304 34216 -32287
rect 33754 -32321 33770 -32304
rect 33182 -32337 33770 -32321
rect 34200 -32321 34216 -32304
rect 34772 -32304 34974 -32287
rect 35032 -32287 35992 -32240
rect 35032 -32304 35234 -32287
rect 34772 -32321 34788 -32304
rect 34200 -32337 34788 -32321
rect 35218 -32321 35234 -32304
rect 35790 -32304 35992 -32287
rect 36050 -32287 37010 -32240
rect 36050 -32304 36252 -32287
rect 35790 -32321 35806 -32304
rect 35218 -32337 35806 -32321
rect 36236 -32321 36252 -32304
rect 36808 -32304 37010 -32287
rect 37068 -32287 38028 -32240
rect 37068 -32304 37270 -32287
rect 36808 -32321 36824 -32304
rect 36236 -32337 36824 -32321
rect 37254 -32321 37270 -32304
rect 37826 -32304 38028 -32287
rect 38086 -32287 39046 -32240
rect 38086 -32304 38288 -32287
rect 37826 -32321 37842 -32304
rect 37254 -32337 37842 -32321
rect 38272 -32321 38288 -32304
rect 38844 -32304 39046 -32287
rect 39104 -32287 40064 -32240
rect 39104 -32304 39306 -32287
rect 38844 -32321 38860 -32304
rect 38272 -32337 38860 -32321
rect 39290 -32321 39306 -32304
rect 39862 -32304 40064 -32287
rect 40122 -32287 41082 -32240
rect 40122 -32304 40324 -32287
rect 39862 -32321 39878 -32304
rect 39290 -32337 39878 -32321
rect 40308 -32321 40324 -32304
rect 40880 -32304 41082 -32287
rect 41140 -32287 42100 -32240
rect 41140 -32304 41342 -32287
rect 40880 -32321 40896 -32304
rect 40308 -32337 40896 -32321
rect 41326 -32321 41342 -32304
rect 41898 -32304 42100 -32287
rect 42158 -32287 43118 -32240
rect 42158 -32304 42360 -32287
rect 41898 -32321 41914 -32304
rect 41326 -32337 41914 -32321
rect 42344 -32321 42360 -32304
rect 42916 -32304 43118 -32287
rect 43176 -32287 44136 -32240
rect 43176 -32304 43378 -32287
rect 42916 -32321 42932 -32304
rect 42344 -32337 42932 -32321
rect 43362 -32321 43378 -32304
rect 43934 -32304 44136 -32287
rect 44194 -32287 45154 -32240
rect 44194 -32304 44396 -32287
rect 43934 -32321 43950 -32304
rect 43362 -32337 43950 -32321
rect 44380 -32321 44396 -32304
rect 44952 -32304 45154 -32287
rect 45212 -32287 46172 -32240
rect 45212 -32304 45414 -32287
rect 44952 -32321 44968 -32304
rect 44380 -32337 44968 -32321
rect 45398 -32321 45414 -32304
rect 45970 -32304 46172 -32287
rect 46230 -32287 47190 -32240
rect 46230 -32304 46432 -32287
rect 45970 -32321 45986 -32304
rect 45398 -32337 45986 -32321
rect 46416 -32321 46432 -32304
rect 46988 -32304 47190 -32287
rect 47248 -32287 48208 -32240
rect 47248 -32304 47450 -32287
rect 46988 -32321 47004 -32304
rect 46416 -32337 47004 -32321
rect 47434 -32321 47450 -32304
rect 48006 -32304 48208 -32287
rect 48006 -32321 48022 -32304
rect 47434 -32337 48022 -32321
rect 32164 -32695 32752 -32679
rect 32164 -32712 32180 -32695
rect 31978 -32729 32180 -32712
rect 32736 -32712 32752 -32695
rect 33182 -32695 33770 -32679
rect 33182 -32712 33198 -32695
rect 32736 -32729 32938 -32712
rect 31978 -32776 32938 -32729
rect 32996 -32729 33198 -32712
rect 33754 -32712 33770 -32695
rect 34200 -32695 34788 -32679
rect 34200 -32712 34216 -32695
rect 33754 -32729 33956 -32712
rect 32996 -32776 33956 -32729
rect 34014 -32729 34216 -32712
rect 34772 -32712 34788 -32695
rect 35218 -32695 35806 -32679
rect 35218 -32712 35234 -32695
rect 34772 -32729 34974 -32712
rect 34014 -32776 34974 -32729
rect 35032 -32729 35234 -32712
rect 35790 -32712 35806 -32695
rect 36236 -32695 36824 -32679
rect 36236 -32712 36252 -32695
rect 35790 -32729 35992 -32712
rect 35032 -32776 35992 -32729
rect 36050 -32729 36252 -32712
rect 36808 -32712 36824 -32695
rect 37254 -32695 37842 -32679
rect 37254 -32712 37270 -32695
rect 36808 -32729 37010 -32712
rect 36050 -32776 37010 -32729
rect 37068 -32729 37270 -32712
rect 37826 -32712 37842 -32695
rect 38272 -32695 38860 -32679
rect 38272 -32712 38288 -32695
rect 37826 -32729 38028 -32712
rect 37068 -32776 38028 -32729
rect 38086 -32729 38288 -32712
rect 38844 -32712 38860 -32695
rect 39290 -32695 39878 -32679
rect 39290 -32712 39306 -32695
rect 38844 -32729 39046 -32712
rect 38086 -32776 39046 -32729
rect 39104 -32729 39306 -32712
rect 39862 -32712 39878 -32695
rect 40308 -32695 40896 -32679
rect 40308 -32712 40324 -32695
rect 39862 -32729 40064 -32712
rect 39104 -32776 40064 -32729
rect 40122 -32729 40324 -32712
rect 40880 -32712 40896 -32695
rect 41326 -32695 41914 -32679
rect 41326 -32712 41342 -32695
rect 40880 -32729 41082 -32712
rect 40122 -32776 41082 -32729
rect 41140 -32729 41342 -32712
rect 41898 -32712 41914 -32695
rect 42344 -32695 42932 -32679
rect 42344 -32712 42360 -32695
rect 41898 -32729 42100 -32712
rect 41140 -32776 42100 -32729
rect 42158 -32729 42360 -32712
rect 42916 -32712 42932 -32695
rect 43362 -32695 43950 -32679
rect 43362 -32712 43378 -32695
rect 42916 -32729 43118 -32712
rect 42158 -32776 43118 -32729
rect 43176 -32729 43378 -32712
rect 43934 -32712 43950 -32695
rect 44380 -32695 44968 -32679
rect 44380 -32712 44396 -32695
rect 43934 -32729 44136 -32712
rect 43176 -32776 44136 -32729
rect 44194 -32729 44396 -32712
rect 44952 -32712 44968 -32695
rect 45398 -32695 45986 -32679
rect 45398 -32712 45414 -32695
rect 44952 -32729 45154 -32712
rect 44194 -32776 45154 -32729
rect 45212 -32729 45414 -32712
rect 45970 -32712 45986 -32695
rect 46416 -32695 47004 -32679
rect 46416 -32712 46432 -32695
rect 45970 -32729 46172 -32712
rect 45212 -32776 46172 -32729
rect 46230 -32729 46432 -32712
rect 46988 -32712 47004 -32695
rect 47434 -32695 48022 -32679
rect 47434 -32712 47450 -32695
rect 46988 -32729 47190 -32712
rect 46230 -32776 47190 -32729
rect 47248 -32729 47450 -32712
rect 48006 -32712 48022 -32695
rect 48006 -32729 48208 -32712
rect 47248 -32776 48208 -32729
rect 31978 -33423 32938 -33376
rect 31978 -33440 32180 -33423
rect 32164 -33457 32180 -33440
rect 32736 -33440 32938 -33423
rect 32996 -33423 33956 -33376
rect 32996 -33440 33198 -33423
rect 32736 -33457 32752 -33440
rect 32164 -33473 32752 -33457
rect 33182 -33457 33198 -33440
rect 33754 -33440 33956 -33423
rect 34014 -33423 34974 -33376
rect 34014 -33440 34216 -33423
rect 33754 -33457 33770 -33440
rect 33182 -33473 33770 -33457
rect 34200 -33457 34216 -33440
rect 34772 -33440 34974 -33423
rect 35032 -33423 35992 -33376
rect 35032 -33440 35234 -33423
rect 34772 -33457 34788 -33440
rect 34200 -33473 34788 -33457
rect 35218 -33457 35234 -33440
rect 35790 -33440 35992 -33423
rect 36050 -33423 37010 -33376
rect 36050 -33440 36252 -33423
rect 35790 -33457 35806 -33440
rect 35218 -33473 35806 -33457
rect 36236 -33457 36252 -33440
rect 36808 -33440 37010 -33423
rect 37068 -33423 38028 -33376
rect 37068 -33440 37270 -33423
rect 36808 -33457 36824 -33440
rect 36236 -33473 36824 -33457
rect 37254 -33457 37270 -33440
rect 37826 -33440 38028 -33423
rect 38086 -33423 39046 -33376
rect 38086 -33440 38288 -33423
rect 37826 -33457 37842 -33440
rect 37254 -33473 37842 -33457
rect 38272 -33457 38288 -33440
rect 38844 -33440 39046 -33423
rect 39104 -33423 40064 -33376
rect 39104 -33440 39306 -33423
rect 38844 -33457 38860 -33440
rect 38272 -33473 38860 -33457
rect 39290 -33457 39306 -33440
rect 39862 -33440 40064 -33423
rect 40122 -33423 41082 -33376
rect 40122 -33440 40324 -33423
rect 39862 -33457 39878 -33440
rect 39290 -33473 39878 -33457
rect 40308 -33457 40324 -33440
rect 40880 -33440 41082 -33423
rect 41140 -33423 42100 -33376
rect 41140 -33440 41342 -33423
rect 40880 -33457 40896 -33440
rect 40308 -33473 40896 -33457
rect 41326 -33457 41342 -33440
rect 41898 -33440 42100 -33423
rect 42158 -33423 43118 -33376
rect 42158 -33440 42360 -33423
rect 41898 -33457 41914 -33440
rect 41326 -33473 41914 -33457
rect 42344 -33457 42360 -33440
rect 42916 -33440 43118 -33423
rect 43176 -33423 44136 -33376
rect 43176 -33440 43378 -33423
rect 42916 -33457 42932 -33440
rect 42344 -33473 42932 -33457
rect 43362 -33457 43378 -33440
rect 43934 -33440 44136 -33423
rect 44194 -33423 45154 -33376
rect 44194 -33440 44396 -33423
rect 43934 -33457 43950 -33440
rect 43362 -33473 43950 -33457
rect 44380 -33457 44396 -33440
rect 44952 -33440 45154 -33423
rect 45212 -33423 46172 -33376
rect 45212 -33440 45414 -33423
rect 44952 -33457 44968 -33440
rect 44380 -33473 44968 -33457
rect 45398 -33457 45414 -33440
rect 45970 -33440 46172 -33423
rect 46230 -33423 47190 -33376
rect 46230 -33440 46432 -33423
rect 45970 -33457 45986 -33440
rect 45398 -33473 45986 -33457
rect 46416 -33457 46432 -33440
rect 46988 -33440 47190 -33423
rect 47248 -33423 48208 -33376
rect 47248 -33440 47450 -33423
rect 46988 -33457 47004 -33440
rect 46416 -33473 47004 -33457
rect 47434 -33457 47450 -33440
rect 48006 -33440 48208 -33423
rect 48006 -33457 48022 -33440
rect 47434 -33473 48022 -33457
rect 33358 -34333 33946 -34317
rect 33358 -34350 33374 -34333
rect 33172 -34367 33374 -34350
rect 33930 -34350 33946 -34333
rect 34376 -34333 34964 -34317
rect 34376 -34350 34392 -34333
rect 33930 -34367 34132 -34350
rect 33172 -34414 34132 -34367
rect 34190 -34367 34392 -34350
rect 34948 -34350 34964 -34333
rect 35394 -34333 35982 -34317
rect 35394 -34350 35410 -34333
rect 34948 -34367 35150 -34350
rect 34190 -34414 35150 -34367
rect 35208 -34367 35410 -34350
rect 35966 -34350 35982 -34333
rect 36412 -34333 37000 -34317
rect 36412 -34350 36428 -34333
rect 35966 -34367 36168 -34350
rect 35208 -34414 36168 -34367
rect 36226 -34367 36428 -34350
rect 36984 -34350 37000 -34333
rect 37430 -34333 38018 -34317
rect 37430 -34350 37446 -34333
rect 36984 -34367 37186 -34350
rect 36226 -34414 37186 -34367
rect 37244 -34367 37446 -34350
rect 38002 -34350 38018 -34333
rect 38448 -34333 39036 -34317
rect 38448 -34350 38464 -34333
rect 38002 -34367 38204 -34350
rect 37244 -34414 38204 -34367
rect 38262 -34367 38464 -34350
rect 39020 -34350 39036 -34333
rect 39466 -34333 40054 -34317
rect 39466 -34350 39482 -34333
rect 39020 -34367 39222 -34350
rect 38262 -34414 39222 -34367
rect 39280 -34367 39482 -34350
rect 40038 -34350 40054 -34333
rect 40484 -34333 41072 -34317
rect 40484 -34350 40500 -34333
rect 40038 -34367 40240 -34350
rect 39280 -34414 40240 -34367
rect 40298 -34367 40500 -34350
rect 41056 -34350 41072 -34333
rect 41502 -34333 42090 -34317
rect 41502 -34350 41518 -34333
rect 41056 -34367 41258 -34350
rect 40298 -34414 41258 -34367
rect 41316 -34367 41518 -34350
rect 42074 -34350 42090 -34333
rect 42520 -34333 43108 -34317
rect 42520 -34350 42536 -34333
rect 42074 -34367 42276 -34350
rect 41316 -34414 42276 -34367
rect 42334 -34367 42536 -34350
rect 43092 -34350 43108 -34333
rect 43538 -34333 44126 -34317
rect 43538 -34350 43554 -34333
rect 43092 -34367 43294 -34350
rect 42334 -34414 43294 -34367
rect 43352 -34367 43554 -34350
rect 44110 -34350 44126 -34333
rect 44556 -34333 45144 -34317
rect 44556 -34350 44572 -34333
rect 44110 -34367 44312 -34350
rect 43352 -34414 44312 -34367
rect 44370 -34367 44572 -34350
rect 45128 -34350 45144 -34333
rect 45574 -34333 46162 -34317
rect 45574 -34350 45590 -34333
rect 45128 -34367 45330 -34350
rect 44370 -34414 45330 -34367
rect 45388 -34367 45590 -34350
rect 46146 -34350 46162 -34333
rect 46592 -34333 47180 -34317
rect 46592 -34350 46608 -34333
rect 46146 -34367 46348 -34350
rect 45388 -34414 46348 -34367
rect 46406 -34367 46608 -34350
rect 47164 -34350 47180 -34333
rect 47164 -34367 47366 -34350
rect 46406 -34414 47366 -34367
rect 33172 -35061 34132 -35014
rect 33172 -35078 33374 -35061
rect 33358 -35095 33374 -35078
rect 33930 -35078 34132 -35061
rect 34190 -35061 35150 -35014
rect 34190 -35078 34392 -35061
rect 33930 -35095 33946 -35078
rect 33358 -35111 33946 -35095
rect 34376 -35095 34392 -35078
rect 34948 -35078 35150 -35061
rect 35208 -35061 36168 -35014
rect 35208 -35078 35410 -35061
rect 34948 -35095 34964 -35078
rect 34376 -35111 34964 -35095
rect 35394 -35095 35410 -35078
rect 35966 -35078 36168 -35061
rect 36226 -35061 37186 -35014
rect 36226 -35078 36428 -35061
rect 35966 -35095 35982 -35078
rect 35394 -35111 35982 -35095
rect 36412 -35095 36428 -35078
rect 36984 -35078 37186 -35061
rect 37244 -35061 38204 -35014
rect 37244 -35078 37446 -35061
rect 36984 -35095 37000 -35078
rect 36412 -35111 37000 -35095
rect 37430 -35095 37446 -35078
rect 38002 -35078 38204 -35061
rect 38262 -35061 39222 -35014
rect 38262 -35078 38464 -35061
rect 38002 -35095 38018 -35078
rect 37430 -35111 38018 -35095
rect 38448 -35095 38464 -35078
rect 39020 -35078 39222 -35061
rect 39280 -35061 40240 -35014
rect 39280 -35078 39482 -35061
rect 39020 -35095 39036 -35078
rect 38448 -35111 39036 -35095
rect 39466 -35095 39482 -35078
rect 40038 -35078 40240 -35061
rect 40298 -35061 41258 -35014
rect 40298 -35078 40500 -35061
rect 40038 -35095 40054 -35078
rect 39466 -35111 40054 -35095
rect 40484 -35095 40500 -35078
rect 41056 -35078 41258 -35061
rect 41316 -35061 42276 -35014
rect 41316 -35078 41518 -35061
rect 41056 -35095 41072 -35078
rect 40484 -35111 41072 -35095
rect 41502 -35095 41518 -35078
rect 42074 -35078 42276 -35061
rect 42334 -35061 43294 -35014
rect 42334 -35078 42536 -35061
rect 42074 -35095 42090 -35078
rect 41502 -35111 42090 -35095
rect 42520 -35095 42536 -35078
rect 43092 -35078 43294 -35061
rect 43352 -35061 44312 -35014
rect 43352 -35078 43554 -35061
rect 43092 -35095 43108 -35078
rect 42520 -35111 43108 -35095
rect 43538 -35095 43554 -35078
rect 44110 -35078 44312 -35061
rect 44370 -35061 45330 -35014
rect 44370 -35078 44572 -35061
rect 44110 -35095 44126 -35078
rect 43538 -35111 44126 -35095
rect 44556 -35095 44572 -35078
rect 45128 -35078 45330 -35061
rect 45388 -35061 46348 -35014
rect 45388 -35078 45590 -35061
rect 45128 -35095 45144 -35078
rect 44556 -35111 45144 -35095
rect 45574 -35095 45590 -35078
rect 46146 -35078 46348 -35061
rect 46406 -35061 47366 -35014
rect 46406 -35078 46608 -35061
rect 46146 -35095 46162 -35078
rect 45574 -35111 46162 -35095
rect 46592 -35095 46608 -35078
rect 47164 -35078 47366 -35061
rect 47164 -35095 47180 -35078
rect 46592 -35111 47180 -35095
rect 33358 -35365 33946 -35349
rect 33358 -35382 33374 -35365
rect 33172 -35399 33374 -35382
rect 33930 -35382 33946 -35365
rect 34376 -35365 34964 -35349
rect 34376 -35382 34392 -35365
rect 33930 -35399 34132 -35382
rect 33172 -35446 34132 -35399
rect 34190 -35399 34392 -35382
rect 34948 -35382 34964 -35365
rect 35394 -35365 35982 -35349
rect 35394 -35382 35410 -35365
rect 34948 -35399 35150 -35382
rect 34190 -35446 35150 -35399
rect 35208 -35399 35410 -35382
rect 35966 -35382 35982 -35365
rect 36412 -35365 37000 -35349
rect 36412 -35382 36428 -35365
rect 35966 -35399 36168 -35382
rect 35208 -35446 36168 -35399
rect 36226 -35399 36428 -35382
rect 36984 -35382 37000 -35365
rect 37430 -35365 38018 -35349
rect 37430 -35382 37446 -35365
rect 36984 -35399 37186 -35382
rect 36226 -35446 37186 -35399
rect 37244 -35399 37446 -35382
rect 38002 -35382 38018 -35365
rect 38448 -35365 39036 -35349
rect 38448 -35382 38464 -35365
rect 38002 -35399 38204 -35382
rect 37244 -35446 38204 -35399
rect 38262 -35399 38464 -35382
rect 39020 -35382 39036 -35365
rect 39466 -35365 40054 -35349
rect 39466 -35382 39482 -35365
rect 39020 -35399 39222 -35382
rect 38262 -35446 39222 -35399
rect 39280 -35399 39482 -35382
rect 40038 -35382 40054 -35365
rect 40484 -35365 41072 -35349
rect 40484 -35382 40500 -35365
rect 40038 -35399 40240 -35382
rect 39280 -35446 40240 -35399
rect 40298 -35399 40500 -35382
rect 41056 -35382 41072 -35365
rect 41502 -35365 42090 -35349
rect 41502 -35382 41518 -35365
rect 41056 -35399 41258 -35382
rect 40298 -35446 41258 -35399
rect 41316 -35399 41518 -35382
rect 42074 -35382 42090 -35365
rect 42520 -35365 43108 -35349
rect 42520 -35382 42536 -35365
rect 42074 -35399 42276 -35382
rect 41316 -35446 42276 -35399
rect 42334 -35399 42536 -35382
rect 43092 -35382 43108 -35365
rect 43538 -35365 44126 -35349
rect 43538 -35382 43554 -35365
rect 43092 -35399 43294 -35382
rect 42334 -35446 43294 -35399
rect 43352 -35399 43554 -35382
rect 44110 -35382 44126 -35365
rect 44556 -35365 45144 -35349
rect 44556 -35382 44572 -35365
rect 44110 -35399 44312 -35382
rect 43352 -35446 44312 -35399
rect 44370 -35399 44572 -35382
rect 45128 -35382 45144 -35365
rect 45574 -35365 46162 -35349
rect 45574 -35382 45590 -35365
rect 45128 -35399 45330 -35382
rect 44370 -35446 45330 -35399
rect 45388 -35399 45590 -35382
rect 46146 -35382 46162 -35365
rect 46592 -35365 47180 -35349
rect 46592 -35382 46608 -35365
rect 46146 -35399 46348 -35382
rect 45388 -35446 46348 -35399
rect 46406 -35399 46608 -35382
rect 47164 -35382 47180 -35365
rect 47164 -35399 47366 -35382
rect 46406 -35446 47366 -35399
rect 33172 -36093 34132 -36046
rect 33172 -36110 33374 -36093
rect 33358 -36127 33374 -36110
rect 33930 -36110 34132 -36093
rect 34190 -36093 35150 -36046
rect 34190 -36110 34392 -36093
rect 33930 -36127 33946 -36110
rect 33358 -36143 33946 -36127
rect 34376 -36127 34392 -36110
rect 34948 -36110 35150 -36093
rect 35208 -36093 36168 -36046
rect 35208 -36110 35410 -36093
rect 34948 -36127 34964 -36110
rect 34376 -36143 34964 -36127
rect 35394 -36127 35410 -36110
rect 35966 -36110 36168 -36093
rect 36226 -36093 37186 -36046
rect 36226 -36110 36428 -36093
rect 35966 -36127 35982 -36110
rect 35394 -36143 35982 -36127
rect 36412 -36127 36428 -36110
rect 36984 -36110 37186 -36093
rect 37244 -36093 38204 -36046
rect 37244 -36110 37446 -36093
rect 36984 -36127 37000 -36110
rect 36412 -36143 37000 -36127
rect 37430 -36127 37446 -36110
rect 38002 -36110 38204 -36093
rect 38262 -36093 39222 -36046
rect 38262 -36110 38464 -36093
rect 38002 -36127 38018 -36110
rect 37430 -36143 38018 -36127
rect 38448 -36127 38464 -36110
rect 39020 -36110 39222 -36093
rect 39280 -36093 40240 -36046
rect 39280 -36110 39482 -36093
rect 39020 -36127 39036 -36110
rect 38448 -36143 39036 -36127
rect 39466 -36127 39482 -36110
rect 40038 -36110 40240 -36093
rect 40298 -36093 41258 -36046
rect 40298 -36110 40500 -36093
rect 40038 -36127 40054 -36110
rect 39466 -36143 40054 -36127
rect 40484 -36127 40500 -36110
rect 41056 -36110 41258 -36093
rect 41316 -36093 42276 -36046
rect 41316 -36110 41518 -36093
rect 41056 -36127 41072 -36110
rect 40484 -36143 41072 -36127
rect 41502 -36127 41518 -36110
rect 42074 -36110 42276 -36093
rect 42334 -36093 43294 -36046
rect 42334 -36110 42536 -36093
rect 42074 -36127 42090 -36110
rect 41502 -36143 42090 -36127
rect 42520 -36127 42536 -36110
rect 43092 -36110 43294 -36093
rect 43352 -36093 44312 -36046
rect 43352 -36110 43554 -36093
rect 43092 -36127 43108 -36110
rect 42520 -36143 43108 -36127
rect 43538 -36127 43554 -36110
rect 44110 -36110 44312 -36093
rect 44370 -36093 45330 -36046
rect 44370 -36110 44572 -36093
rect 44110 -36127 44126 -36110
rect 43538 -36143 44126 -36127
rect 44556 -36127 44572 -36110
rect 45128 -36110 45330 -36093
rect 45388 -36093 46348 -36046
rect 45388 -36110 45590 -36093
rect 45128 -36127 45144 -36110
rect 44556 -36143 45144 -36127
rect 45574 -36127 45590 -36110
rect 46146 -36110 46348 -36093
rect 46406 -36093 47366 -36046
rect 46406 -36110 46608 -36093
rect 46146 -36127 46162 -36110
rect 45574 -36143 46162 -36127
rect 46592 -36127 46608 -36110
rect 47164 -36110 47366 -36093
rect 47164 -36127 47180 -36110
rect 46592 -36143 47180 -36127
rect 33150 -36969 33738 -36953
rect 33150 -36986 33166 -36969
rect 32964 -37003 33166 -36986
rect 33722 -36986 33738 -36969
rect 34168 -36969 34756 -36953
rect 34168 -36986 34184 -36969
rect 33722 -37003 33924 -36986
rect 32964 -37050 33924 -37003
rect 33982 -37003 34184 -36986
rect 34740 -36986 34756 -36969
rect 35186 -36969 35774 -36953
rect 35186 -36986 35202 -36969
rect 34740 -37003 34942 -36986
rect 33982 -37050 34942 -37003
rect 35000 -37003 35202 -36986
rect 35758 -36986 35774 -36969
rect 36204 -36969 36792 -36953
rect 36204 -36986 36220 -36969
rect 35758 -37003 35960 -36986
rect 35000 -37050 35960 -37003
rect 36018 -37003 36220 -36986
rect 36776 -36986 36792 -36969
rect 37222 -36969 37810 -36953
rect 37222 -36986 37238 -36969
rect 36776 -37003 36978 -36986
rect 36018 -37050 36978 -37003
rect 37036 -37003 37238 -36986
rect 37794 -36986 37810 -36969
rect 38240 -36969 38828 -36953
rect 38240 -36986 38256 -36969
rect 37794 -37003 37996 -36986
rect 37036 -37050 37996 -37003
rect 38054 -37003 38256 -36986
rect 38812 -36986 38828 -36969
rect 39258 -36969 39846 -36953
rect 39258 -36986 39274 -36969
rect 38812 -37003 39014 -36986
rect 38054 -37050 39014 -37003
rect 39072 -37003 39274 -36986
rect 39830 -36986 39846 -36969
rect 40276 -36969 40864 -36953
rect 40276 -36986 40292 -36969
rect 39830 -37003 40032 -36986
rect 39072 -37050 40032 -37003
rect 40090 -37003 40292 -36986
rect 40848 -36986 40864 -36969
rect 41294 -36969 41882 -36953
rect 41294 -36986 41310 -36969
rect 40848 -37003 41050 -36986
rect 40090 -37050 41050 -37003
rect 41108 -37003 41310 -36986
rect 41866 -36986 41882 -36969
rect 42312 -36969 42900 -36953
rect 42312 -36986 42328 -36969
rect 41866 -37003 42068 -36986
rect 41108 -37050 42068 -37003
rect 42126 -37003 42328 -36986
rect 42884 -36986 42900 -36969
rect 43330 -36969 43918 -36953
rect 43330 -36986 43346 -36969
rect 42884 -37003 43086 -36986
rect 42126 -37050 43086 -37003
rect 43144 -37003 43346 -36986
rect 43902 -36986 43918 -36969
rect 44348 -36969 44936 -36953
rect 44348 -36986 44364 -36969
rect 43902 -37003 44104 -36986
rect 43144 -37050 44104 -37003
rect 44162 -37003 44364 -36986
rect 44920 -36986 44936 -36969
rect 45366 -36969 45954 -36953
rect 45366 -36986 45382 -36969
rect 44920 -37003 45122 -36986
rect 44162 -37050 45122 -37003
rect 45180 -37003 45382 -36986
rect 45938 -36986 45954 -36969
rect 46384 -36969 46972 -36953
rect 46384 -36986 46400 -36969
rect 45938 -37003 46140 -36986
rect 45180 -37050 46140 -37003
rect 46198 -37003 46400 -36986
rect 46956 -36986 46972 -36969
rect 47402 -36969 47990 -36953
rect 47402 -36986 47418 -36969
rect 46956 -37003 47158 -36986
rect 46198 -37050 47158 -37003
rect 47216 -37003 47418 -36986
rect 47974 -36986 47990 -36969
rect 47974 -37003 48176 -36986
rect 47216 -37050 48176 -37003
rect 27846 -37073 28434 -37057
rect 27846 -37090 27862 -37073
rect 27660 -37107 27862 -37090
rect 28418 -37090 28434 -37073
rect 28864 -37073 29452 -37057
rect 28864 -37090 28880 -37073
rect 28418 -37107 28620 -37090
rect 27660 -37154 28620 -37107
rect 28678 -37107 28880 -37090
rect 29436 -37090 29452 -37073
rect 29882 -37073 30470 -37057
rect 29882 -37090 29898 -37073
rect 29436 -37107 29638 -37090
rect 28678 -37154 29638 -37107
rect 29696 -37107 29898 -37090
rect 30454 -37090 30470 -37073
rect 30900 -37073 31488 -37057
rect 30900 -37090 30916 -37073
rect 30454 -37107 30656 -37090
rect 29696 -37154 30656 -37107
rect 30714 -37107 30916 -37090
rect 31472 -37090 31488 -37073
rect 31472 -37107 31674 -37090
rect 30714 -37154 31674 -37107
rect 32964 -37697 33924 -37650
rect 32964 -37714 33166 -37697
rect 33150 -37731 33166 -37714
rect 33722 -37714 33924 -37697
rect 33982 -37697 34942 -37650
rect 33982 -37714 34184 -37697
rect 33722 -37731 33738 -37714
rect 33150 -37747 33738 -37731
rect 34168 -37731 34184 -37714
rect 34740 -37714 34942 -37697
rect 35000 -37697 35960 -37650
rect 35000 -37714 35202 -37697
rect 34740 -37731 34756 -37714
rect 34168 -37747 34756 -37731
rect 35186 -37731 35202 -37714
rect 35758 -37714 35960 -37697
rect 36018 -37697 36978 -37650
rect 36018 -37714 36220 -37697
rect 35758 -37731 35774 -37714
rect 35186 -37747 35774 -37731
rect 36204 -37731 36220 -37714
rect 36776 -37714 36978 -37697
rect 37036 -37697 37996 -37650
rect 37036 -37714 37238 -37697
rect 36776 -37731 36792 -37714
rect 36204 -37747 36792 -37731
rect 37222 -37731 37238 -37714
rect 37794 -37714 37996 -37697
rect 38054 -37697 39014 -37650
rect 38054 -37714 38256 -37697
rect 37794 -37731 37810 -37714
rect 37222 -37747 37810 -37731
rect 38240 -37731 38256 -37714
rect 38812 -37714 39014 -37697
rect 39072 -37697 40032 -37650
rect 39072 -37714 39274 -37697
rect 38812 -37731 38828 -37714
rect 38240 -37747 38828 -37731
rect 39258 -37731 39274 -37714
rect 39830 -37714 40032 -37697
rect 40090 -37697 41050 -37650
rect 40090 -37714 40292 -37697
rect 39830 -37731 39846 -37714
rect 39258 -37747 39846 -37731
rect 40276 -37731 40292 -37714
rect 40848 -37714 41050 -37697
rect 41108 -37697 42068 -37650
rect 41108 -37714 41310 -37697
rect 40848 -37731 40864 -37714
rect 40276 -37747 40864 -37731
rect 41294 -37731 41310 -37714
rect 41866 -37714 42068 -37697
rect 42126 -37697 43086 -37650
rect 42126 -37714 42328 -37697
rect 41866 -37731 41882 -37714
rect 41294 -37747 41882 -37731
rect 42312 -37731 42328 -37714
rect 42884 -37714 43086 -37697
rect 43144 -37697 44104 -37650
rect 43144 -37714 43346 -37697
rect 42884 -37731 42900 -37714
rect 42312 -37747 42900 -37731
rect 43330 -37731 43346 -37714
rect 43902 -37714 44104 -37697
rect 44162 -37697 45122 -37650
rect 44162 -37714 44364 -37697
rect 43902 -37731 43918 -37714
rect 43330 -37747 43918 -37731
rect 44348 -37731 44364 -37714
rect 44920 -37714 45122 -37697
rect 45180 -37697 46140 -37650
rect 45180 -37714 45382 -37697
rect 44920 -37731 44936 -37714
rect 44348 -37747 44936 -37731
rect 45366 -37731 45382 -37714
rect 45938 -37714 46140 -37697
rect 46198 -37697 47158 -37650
rect 46198 -37714 46400 -37697
rect 45938 -37731 45954 -37714
rect 45366 -37747 45954 -37731
rect 46384 -37731 46400 -37714
rect 46956 -37714 47158 -37697
rect 47216 -37697 48176 -37650
rect 47216 -37714 47418 -37697
rect 46956 -37731 46972 -37714
rect 46384 -37747 46972 -37731
rect 47402 -37731 47418 -37714
rect 47974 -37714 48176 -37697
rect 47974 -37731 47990 -37714
rect 47402 -37747 47990 -37731
rect 27660 -37801 28620 -37754
rect 27660 -37818 27862 -37801
rect 27846 -37835 27862 -37818
rect 28418 -37818 28620 -37801
rect 28678 -37801 29638 -37754
rect 28678 -37818 28880 -37801
rect 28418 -37835 28434 -37818
rect 27846 -37851 28434 -37835
rect 28864 -37835 28880 -37818
rect 29436 -37818 29638 -37801
rect 29696 -37801 30656 -37754
rect 29696 -37818 29898 -37801
rect 29436 -37835 29452 -37818
rect 28864 -37851 29452 -37835
rect 29882 -37835 29898 -37818
rect 30454 -37818 30656 -37801
rect 30714 -37801 31674 -37754
rect 30714 -37818 30916 -37801
rect 30454 -37835 30470 -37818
rect 29882 -37851 30470 -37835
rect 30900 -37835 30916 -37818
rect 31472 -37818 31674 -37801
rect 31472 -37835 31488 -37818
rect 30900 -37851 31488 -37835
rect 27846 -38105 28434 -38089
rect 27846 -38122 27862 -38105
rect 27660 -38139 27862 -38122
rect 28418 -38122 28434 -38105
rect 28864 -38105 29452 -38089
rect 28864 -38122 28880 -38105
rect 28418 -38139 28620 -38122
rect 27660 -38186 28620 -38139
rect 28678 -38139 28880 -38122
rect 29436 -38122 29452 -38105
rect 29882 -38105 30470 -38089
rect 29882 -38122 29898 -38105
rect 29436 -38139 29638 -38122
rect 28678 -38186 29638 -38139
rect 29696 -38139 29898 -38122
rect 30454 -38122 30470 -38105
rect 30900 -38105 31488 -38089
rect 30900 -38122 30916 -38105
rect 30454 -38139 30656 -38122
rect 29696 -38186 30656 -38139
rect 30714 -38139 30916 -38122
rect 31472 -38122 31488 -38105
rect 31472 -38139 31674 -38122
rect 30714 -38186 31674 -38139
rect 33150 -38225 33738 -38209
rect 33150 -38242 33166 -38225
rect 32964 -38259 33166 -38242
rect 33722 -38242 33738 -38225
rect 34168 -38225 34756 -38209
rect 34168 -38242 34184 -38225
rect 33722 -38259 33924 -38242
rect 32964 -38306 33924 -38259
rect 33982 -38259 34184 -38242
rect 34740 -38242 34756 -38225
rect 35186 -38225 35774 -38209
rect 35186 -38242 35202 -38225
rect 34740 -38259 34942 -38242
rect 33982 -38306 34942 -38259
rect 35000 -38259 35202 -38242
rect 35758 -38242 35774 -38225
rect 36204 -38225 36792 -38209
rect 36204 -38242 36220 -38225
rect 35758 -38259 35960 -38242
rect 35000 -38306 35960 -38259
rect 36018 -38259 36220 -38242
rect 36776 -38242 36792 -38225
rect 37222 -38225 37810 -38209
rect 37222 -38242 37238 -38225
rect 36776 -38259 36978 -38242
rect 36018 -38306 36978 -38259
rect 37036 -38259 37238 -38242
rect 37794 -38242 37810 -38225
rect 38240 -38225 38828 -38209
rect 38240 -38242 38256 -38225
rect 37794 -38259 37996 -38242
rect 37036 -38306 37996 -38259
rect 38054 -38259 38256 -38242
rect 38812 -38242 38828 -38225
rect 39258 -38225 39846 -38209
rect 39258 -38242 39274 -38225
rect 38812 -38259 39014 -38242
rect 38054 -38306 39014 -38259
rect 39072 -38259 39274 -38242
rect 39830 -38242 39846 -38225
rect 40276 -38225 40864 -38209
rect 40276 -38242 40292 -38225
rect 39830 -38259 40032 -38242
rect 39072 -38306 40032 -38259
rect 40090 -38259 40292 -38242
rect 40848 -38242 40864 -38225
rect 41294 -38225 41882 -38209
rect 41294 -38242 41310 -38225
rect 40848 -38259 41050 -38242
rect 40090 -38306 41050 -38259
rect 41108 -38259 41310 -38242
rect 41866 -38242 41882 -38225
rect 42312 -38225 42900 -38209
rect 42312 -38242 42328 -38225
rect 41866 -38259 42068 -38242
rect 41108 -38306 42068 -38259
rect 42126 -38259 42328 -38242
rect 42884 -38242 42900 -38225
rect 43330 -38225 43918 -38209
rect 43330 -38242 43346 -38225
rect 42884 -38259 43086 -38242
rect 42126 -38306 43086 -38259
rect 43144 -38259 43346 -38242
rect 43902 -38242 43918 -38225
rect 44348 -38225 44936 -38209
rect 44348 -38242 44364 -38225
rect 43902 -38259 44104 -38242
rect 43144 -38306 44104 -38259
rect 44162 -38259 44364 -38242
rect 44920 -38242 44936 -38225
rect 45366 -38225 45954 -38209
rect 45366 -38242 45382 -38225
rect 44920 -38259 45122 -38242
rect 44162 -38306 45122 -38259
rect 45180 -38259 45382 -38242
rect 45938 -38242 45954 -38225
rect 46384 -38225 46972 -38209
rect 46384 -38242 46400 -38225
rect 45938 -38259 46140 -38242
rect 45180 -38306 46140 -38259
rect 46198 -38259 46400 -38242
rect 46956 -38242 46972 -38225
rect 47402 -38225 47990 -38209
rect 47402 -38242 47418 -38225
rect 46956 -38259 47158 -38242
rect 46198 -38306 47158 -38259
rect 47216 -38259 47418 -38242
rect 47974 -38242 47990 -38225
rect 47974 -38259 48176 -38242
rect 47216 -38306 48176 -38259
rect 27660 -38833 28620 -38786
rect 27660 -38850 27862 -38833
rect 27846 -38867 27862 -38850
rect 28418 -38850 28620 -38833
rect 28678 -38833 29638 -38786
rect 28678 -38850 28880 -38833
rect 28418 -38867 28434 -38850
rect 27846 -38883 28434 -38867
rect 28864 -38867 28880 -38850
rect 29436 -38850 29638 -38833
rect 29696 -38833 30656 -38786
rect 29696 -38850 29898 -38833
rect 29436 -38867 29452 -38850
rect 28864 -38883 29452 -38867
rect 29882 -38867 29898 -38850
rect 30454 -38850 30656 -38833
rect 30714 -38833 31674 -38786
rect 30714 -38850 30916 -38833
rect 30454 -38867 30470 -38850
rect 29882 -38883 30470 -38867
rect 30900 -38867 30916 -38850
rect 31472 -38850 31674 -38833
rect 31472 -38867 31488 -38850
rect 30900 -38883 31488 -38867
rect 32964 -38953 33924 -38906
rect 32964 -38970 33166 -38953
rect 33150 -38987 33166 -38970
rect 33722 -38970 33924 -38953
rect 33982 -38953 34942 -38906
rect 33982 -38970 34184 -38953
rect 33722 -38987 33738 -38970
rect 33150 -39003 33738 -38987
rect 34168 -38987 34184 -38970
rect 34740 -38970 34942 -38953
rect 35000 -38953 35960 -38906
rect 35000 -38970 35202 -38953
rect 34740 -38987 34756 -38970
rect 34168 -39003 34756 -38987
rect 35186 -38987 35202 -38970
rect 35758 -38970 35960 -38953
rect 36018 -38953 36978 -38906
rect 36018 -38970 36220 -38953
rect 35758 -38987 35774 -38970
rect 35186 -39003 35774 -38987
rect 36204 -38987 36220 -38970
rect 36776 -38970 36978 -38953
rect 37036 -38953 37996 -38906
rect 37036 -38970 37238 -38953
rect 36776 -38987 36792 -38970
rect 36204 -39003 36792 -38987
rect 37222 -38987 37238 -38970
rect 37794 -38970 37996 -38953
rect 38054 -38953 39014 -38906
rect 38054 -38970 38256 -38953
rect 37794 -38987 37810 -38970
rect 37222 -39003 37810 -38987
rect 38240 -38987 38256 -38970
rect 38812 -38970 39014 -38953
rect 39072 -38953 40032 -38906
rect 39072 -38970 39274 -38953
rect 38812 -38987 38828 -38970
rect 38240 -39003 38828 -38987
rect 39258 -38987 39274 -38970
rect 39830 -38970 40032 -38953
rect 40090 -38953 41050 -38906
rect 40090 -38970 40292 -38953
rect 39830 -38987 39846 -38970
rect 39258 -39003 39846 -38987
rect 40276 -38987 40292 -38970
rect 40848 -38970 41050 -38953
rect 41108 -38953 42068 -38906
rect 41108 -38970 41310 -38953
rect 40848 -38987 40864 -38970
rect 40276 -39003 40864 -38987
rect 41294 -38987 41310 -38970
rect 41866 -38970 42068 -38953
rect 42126 -38953 43086 -38906
rect 42126 -38970 42328 -38953
rect 41866 -38987 41882 -38970
rect 41294 -39003 41882 -38987
rect 42312 -38987 42328 -38970
rect 42884 -38970 43086 -38953
rect 43144 -38953 44104 -38906
rect 43144 -38970 43346 -38953
rect 42884 -38987 42900 -38970
rect 42312 -39003 42900 -38987
rect 43330 -38987 43346 -38970
rect 43902 -38970 44104 -38953
rect 44162 -38953 45122 -38906
rect 44162 -38970 44364 -38953
rect 43902 -38987 43918 -38970
rect 43330 -39003 43918 -38987
rect 44348 -38987 44364 -38970
rect 44920 -38970 45122 -38953
rect 45180 -38953 46140 -38906
rect 45180 -38970 45382 -38953
rect 44920 -38987 44936 -38970
rect 44348 -39003 44936 -38987
rect 45366 -38987 45382 -38970
rect 45938 -38970 46140 -38953
rect 46198 -38953 47158 -38906
rect 46198 -38970 46400 -38953
rect 45938 -38987 45954 -38970
rect 45366 -39003 45954 -38987
rect 46384 -38987 46400 -38970
rect 46956 -38970 47158 -38953
rect 47216 -38953 48176 -38906
rect 47216 -38970 47418 -38953
rect 46956 -38987 46972 -38970
rect 46384 -39003 46972 -38987
rect 47402 -38987 47418 -38970
rect 47974 -38970 48176 -38953
rect 47974 -38987 47990 -38970
rect 47402 -39003 47990 -38987
rect 27846 -39137 28434 -39121
rect 27846 -39154 27862 -39137
rect 27660 -39171 27862 -39154
rect 28418 -39154 28434 -39137
rect 28864 -39137 29452 -39121
rect 28864 -39154 28880 -39137
rect 28418 -39171 28620 -39154
rect 27660 -39218 28620 -39171
rect 28678 -39171 28880 -39154
rect 29436 -39154 29452 -39137
rect 29882 -39137 30470 -39121
rect 29882 -39154 29898 -39137
rect 29436 -39171 29638 -39154
rect 28678 -39218 29638 -39171
rect 29696 -39171 29898 -39154
rect 30454 -39154 30470 -39137
rect 30900 -39137 31488 -39121
rect 30900 -39154 30916 -39137
rect 30454 -39171 30656 -39154
rect 29696 -39218 30656 -39171
rect 30714 -39171 30916 -39154
rect 31472 -39154 31488 -39137
rect 31472 -39171 31674 -39154
rect 30714 -39218 31674 -39171
rect 33150 -39481 33738 -39465
rect 33150 -39498 33166 -39481
rect 32964 -39515 33166 -39498
rect 33722 -39498 33738 -39481
rect 34168 -39481 34756 -39465
rect 34168 -39498 34184 -39481
rect 33722 -39515 33924 -39498
rect 32964 -39562 33924 -39515
rect 33982 -39515 34184 -39498
rect 34740 -39498 34756 -39481
rect 35186 -39481 35774 -39465
rect 35186 -39498 35202 -39481
rect 34740 -39515 34942 -39498
rect 33982 -39562 34942 -39515
rect 35000 -39515 35202 -39498
rect 35758 -39498 35774 -39481
rect 36204 -39481 36792 -39465
rect 36204 -39498 36220 -39481
rect 35758 -39515 35960 -39498
rect 35000 -39562 35960 -39515
rect 36018 -39515 36220 -39498
rect 36776 -39498 36792 -39481
rect 37222 -39481 37810 -39465
rect 37222 -39498 37238 -39481
rect 36776 -39515 36978 -39498
rect 36018 -39562 36978 -39515
rect 37036 -39515 37238 -39498
rect 37794 -39498 37810 -39481
rect 38240 -39481 38828 -39465
rect 38240 -39498 38256 -39481
rect 37794 -39515 37996 -39498
rect 37036 -39562 37996 -39515
rect 38054 -39515 38256 -39498
rect 38812 -39498 38828 -39481
rect 39258 -39481 39846 -39465
rect 39258 -39498 39274 -39481
rect 38812 -39515 39014 -39498
rect 38054 -39562 39014 -39515
rect 39072 -39515 39274 -39498
rect 39830 -39498 39846 -39481
rect 40276 -39481 40864 -39465
rect 40276 -39498 40292 -39481
rect 39830 -39515 40032 -39498
rect 39072 -39562 40032 -39515
rect 40090 -39515 40292 -39498
rect 40848 -39498 40864 -39481
rect 41294 -39481 41882 -39465
rect 41294 -39498 41310 -39481
rect 40848 -39515 41050 -39498
rect 40090 -39562 41050 -39515
rect 41108 -39515 41310 -39498
rect 41866 -39498 41882 -39481
rect 42312 -39481 42900 -39465
rect 42312 -39498 42328 -39481
rect 41866 -39515 42068 -39498
rect 41108 -39562 42068 -39515
rect 42126 -39515 42328 -39498
rect 42884 -39498 42900 -39481
rect 43330 -39481 43918 -39465
rect 43330 -39498 43346 -39481
rect 42884 -39515 43086 -39498
rect 42126 -39562 43086 -39515
rect 43144 -39515 43346 -39498
rect 43902 -39498 43918 -39481
rect 44348 -39481 44936 -39465
rect 44348 -39498 44364 -39481
rect 43902 -39515 44104 -39498
rect 43144 -39562 44104 -39515
rect 44162 -39515 44364 -39498
rect 44920 -39498 44936 -39481
rect 45366 -39481 45954 -39465
rect 45366 -39498 45382 -39481
rect 44920 -39515 45122 -39498
rect 44162 -39562 45122 -39515
rect 45180 -39515 45382 -39498
rect 45938 -39498 45954 -39481
rect 46384 -39481 46972 -39465
rect 46384 -39498 46400 -39481
rect 45938 -39515 46140 -39498
rect 45180 -39562 46140 -39515
rect 46198 -39515 46400 -39498
rect 46956 -39498 46972 -39481
rect 47402 -39481 47990 -39465
rect 47402 -39498 47418 -39481
rect 46956 -39515 47158 -39498
rect 46198 -39562 47158 -39515
rect 47216 -39515 47418 -39498
rect 47974 -39498 47990 -39481
rect 47974 -39515 48176 -39498
rect 47216 -39562 48176 -39515
rect 27660 -39865 28620 -39818
rect 27660 -39882 27862 -39865
rect 27846 -39899 27862 -39882
rect 28418 -39882 28620 -39865
rect 28678 -39865 29638 -39818
rect 28678 -39882 28880 -39865
rect 28418 -39899 28434 -39882
rect 27846 -39915 28434 -39899
rect 28864 -39899 28880 -39882
rect 29436 -39882 29638 -39865
rect 29696 -39865 30656 -39818
rect 29696 -39882 29898 -39865
rect 29436 -39899 29452 -39882
rect 28864 -39915 29452 -39899
rect 29882 -39899 29898 -39882
rect 30454 -39882 30656 -39865
rect 30714 -39865 31674 -39818
rect 30714 -39882 30916 -39865
rect 30454 -39899 30470 -39882
rect 29882 -39915 30470 -39899
rect 30900 -39899 30916 -39882
rect 31472 -39882 31674 -39865
rect 31472 -39899 31488 -39882
rect 30900 -39915 31488 -39899
rect 27846 -40169 28434 -40153
rect 27846 -40186 27862 -40169
rect 27660 -40203 27862 -40186
rect 28418 -40186 28434 -40169
rect 28864 -40169 29452 -40153
rect 28864 -40186 28880 -40169
rect 28418 -40203 28620 -40186
rect 27660 -40250 28620 -40203
rect 28678 -40203 28880 -40186
rect 29436 -40186 29452 -40169
rect 29882 -40169 30470 -40153
rect 29882 -40186 29898 -40169
rect 29436 -40203 29638 -40186
rect 28678 -40250 29638 -40203
rect 29696 -40203 29898 -40186
rect 30454 -40186 30470 -40169
rect 30900 -40169 31488 -40153
rect 30900 -40186 30916 -40169
rect 30454 -40203 30656 -40186
rect 29696 -40250 30656 -40203
rect 30714 -40203 30916 -40186
rect 31472 -40186 31488 -40169
rect 31472 -40203 31674 -40186
rect 30714 -40250 31674 -40203
rect 32964 -40209 33924 -40162
rect 32964 -40226 33166 -40209
rect 33150 -40243 33166 -40226
rect 33722 -40226 33924 -40209
rect 33982 -40209 34942 -40162
rect 33982 -40226 34184 -40209
rect 33722 -40243 33738 -40226
rect 33150 -40259 33738 -40243
rect 34168 -40243 34184 -40226
rect 34740 -40226 34942 -40209
rect 35000 -40209 35960 -40162
rect 35000 -40226 35202 -40209
rect 34740 -40243 34756 -40226
rect 34168 -40259 34756 -40243
rect 35186 -40243 35202 -40226
rect 35758 -40226 35960 -40209
rect 36018 -40209 36978 -40162
rect 36018 -40226 36220 -40209
rect 35758 -40243 35774 -40226
rect 35186 -40259 35774 -40243
rect 36204 -40243 36220 -40226
rect 36776 -40226 36978 -40209
rect 37036 -40209 37996 -40162
rect 37036 -40226 37238 -40209
rect 36776 -40243 36792 -40226
rect 36204 -40259 36792 -40243
rect 37222 -40243 37238 -40226
rect 37794 -40226 37996 -40209
rect 38054 -40209 39014 -40162
rect 38054 -40226 38256 -40209
rect 37794 -40243 37810 -40226
rect 37222 -40259 37810 -40243
rect 38240 -40243 38256 -40226
rect 38812 -40226 39014 -40209
rect 39072 -40209 40032 -40162
rect 39072 -40226 39274 -40209
rect 38812 -40243 38828 -40226
rect 38240 -40259 38828 -40243
rect 39258 -40243 39274 -40226
rect 39830 -40226 40032 -40209
rect 40090 -40209 41050 -40162
rect 40090 -40226 40292 -40209
rect 39830 -40243 39846 -40226
rect 39258 -40259 39846 -40243
rect 40276 -40243 40292 -40226
rect 40848 -40226 41050 -40209
rect 41108 -40209 42068 -40162
rect 41108 -40226 41310 -40209
rect 40848 -40243 40864 -40226
rect 40276 -40259 40864 -40243
rect 41294 -40243 41310 -40226
rect 41866 -40226 42068 -40209
rect 42126 -40209 43086 -40162
rect 42126 -40226 42328 -40209
rect 41866 -40243 41882 -40226
rect 41294 -40259 41882 -40243
rect 42312 -40243 42328 -40226
rect 42884 -40226 43086 -40209
rect 43144 -40209 44104 -40162
rect 43144 -40226 43346 -40209
rect 42884 -40243 42900 -40226
rect 42312 -40259 42900 -40243
rect 43330 -40243 43346 -40226
rect 43902 -40226 44104 -40209
rect 44162 -40209 45122 -40162
rect 44162 -40226 44364 -40209
rect 43902 -40243 43918 -40226
rect 43330 -40259 43918 -40243
rect 44348 -40243 44364 -40226
rect 44920 -40226 45122 -40209
rect 45180 -40209 46140 -40162
rect 45180 -40226 45382 -40209
rect 44920 -40243 44936 -40226
rect 44348 -40259 44936 -40243
rect 45366 -40243 45382 -40226
rect 45938 -40226 46140 -40209
rect 46198 -40209 47158 -40162
rect 46198 -40226 46400 -40209
rect 45938 -40243 45954 -40226
rect 45366 -40259 45954 -40243
rect 46384 -40243 46400 -40226
rect 46956 -40226 47158 -40209
rect 47216 -40209 48176 -40162
rect 47216 -40226 47418 -40209
rect 46956 -40243 46972 -40226
rect 46384 -40259 46972 -40243
rect 47402 -40243 47418 -40226
rect 47974 -40226 48176 -40209
rect 47974 -40243 47990 -40226
rect 47402 -40259 47990 -40243
rect 33150 -40737 33738 -40721
rect 33150 -40754 33166 -40737
rect 32964 -40771 33166 -40754
rect 33722 -40754 33738 -40737
rect 34168 -40737 34756 -40721
rect 34168 -40754 34184 -40737
rect 33722 -40771 33924 -40754
rect 32964 -40818 33924 -40771
rect 33982 -40771 34184 -40754
rect 34740 -40754 34756 -40737
rect 35186 -40737 35774 -40721
rect 35186 -40754 35202 -40737
rect 34740 -40771 34942 -40754
rect 33982 -40818 34942 -40771
rect 35000 -40771 35202 -40754
rect 35758 -40754 35774 -40737
rect 36204 -40737 36792 -40721
rect 36204 -40754 36220 -40737
rect 35758 -40771 35960 -40754
rect 35000 -40818 35960 -40771
rect 36018 -40771 36220 -40754
rect 36776 -40754 36792 -40737
rect 37222 -40737 37810 -40721
rect 37222 -40754 37238 -40737
rect 36776 -40771 36978 -40754
rect 36018 -40818 36978 -40771
rect 37036 -40771 37238 -40754
rect 37794 -40754 37810 -40737
rect 38240 -40737 38828 -40721
rect 38240 -40754 38256 -40737
rect 37794 -40771 37996 -40754
rect 37036 -40818 37996 -40771
rect 38054 -40771 38256 -40754
rect 38812 -40754 38828 -40737
rect 39258 -40737 39846 -40721
rect 39258 -40754 39274 -40737
rect 38812 -40771 39014 -40754
rect 38054 -40818 39014 -40771
rect 39072 -40771 39274 -40754
rect 39830 -40754 39846 -40737
rect 40276 -40737 40864 -40721
rect 40276 -40754 40292 -40737
rect 39830 -40771 40032 -40754
rect 39072 -40818 40032 -40771
rect 40090 -40771 40292 -40754
rect 40848 -40754 40864 -40737
rect 41294 -40737 41882 -40721
rect 41294 -40754 41310 -40737
rect 40848 -40771 41050 -40754
rect 40090 -40818 41050 -40771
rect 41108 -40771 41310 -40754
rect 41866 -40754 41882 -40737
rect 42312 -40737 42900 -40721
rect 42312 -40754 42328 -40737
rect 41866 -40771 42068 -40754
rect 41108 -40818 42068 -40771
rect 42126 -40771 42328 -40754
rect 42884 -40754 42900 -40737
rect 43330 -40737 43918 -40721
rect 43330 -40754 43346 -40737
rect 42884 -40771 43086 -40754
rect 42126 -40818 43086 -40771
rect 43144 -40771 43346 -40754
rect 43902 -40754 43918 -40737
rect 44348 -40737 44936 -40721
rect 44348 -40754 44364 -40737
rect 43902 -40771 44104 -40754
rect 43144 -40818 44104 -40771
rect 44162 -40771 44364 -40754
rect 44920 -40754 44936 -40737
rect 45366 -40737 45954 -40721
rect 45366 -40754 45382 -40737
rect 44920 -40771 45122 -40754
rect 44162 -40818 45122 -40771
rect 45180 -40771 45382 -40754
rect 45938 -40754 45954 -40737
rect 46384 -40737 46972 -40721
rect 46384 -40754 46400 -40737
rect 45938 -40771 46140 -40754
rect 45180 -40818 46140 -40771
rect 46198 -40771 46400 -40754
rect 46956 -40754 46972 -40737
rect 47402 -40737 47990 -40721
rect 47402 -40754 47418 -40737
rect 46956 -40771 47158 -40754
rect 46198 -40818 47158 -40771
rect 47216 -40771 47418 -40754
rect 47974 -40754 47990 -40737
rect 47974 -40771 48176 -40754
rect 47216 -40818 48176 -40771
rect 27660 -40897 28620 -40850
rect 27660 -40914 27862 -40897
rect 27846 -40931 27862 -40914
rect 28418 -40914 28620 -40897
rect 28678 -40897 29638 -40850
rect 28678 -40914 28880 -40897
rect 28418 -40931 28434 -40914
rect 27846 -40947 28434 -40931
rect 28864 -40931 28880 -40914
rect 29436 -40914 29638 -40897
rect 29696 -40897 30656 -40850
rect 29696 -40914 29898 -40897
rect 29436 -40931 29452 -40914
rect 28864 -40947 29452 -40931
rect 29882 -40931 29898 -40914
rect 30454 -40914 30656 -40897
rect 30714 -40897 31674 -40850
rect 30714 -40914 30916 -40897
rect 30454 -40931 30470 -40914
rect 29882 -40947 30470 -40931
rect 30900 -40931 30916 -40914
rect 31472 -40914 31674 -40897
rect 31472 -40931 31488 -40914
rect 30900 -40947 31488 -40931
rect 32964 -41465 33924 -41418
rect 32964 -41482 33166 -41465
rect 33150 -41499 33166 -41482
rect 33722 -41482 33924 -41465
rect 33982 -41465 34942 -41418
rect 33982 -41482 34184 -41465
rect 33722 -41499 33738 -41482
rect 33150 -41515 33738 -41499
rect 34168 -41499 34184 -41482
rect 34740 -41482 34942 -41465
rect 35000 -41465 35960 -41418
rect 35000 -41482 35202 -41465
rect 34740 -41499 34756 -41482
rect 34168 -41515 34756 -41499
rect 35186 -41499 35202 -41482
rect 35758 -41482 35960 -41465
rect 36018 -41465 36978 -41418
rect 36018 -41482 36220 -41465
rect 35758 -41499 35774 -41482
rect 35186 -41515 35774 -41499
rect 36204 -41499 36220 -41482
rect 36776 -41482 36978 -41465
rect 37036 -41465 37996 -41418
rect 37036 -41482 37238 -41465
rect 36776 -41499 36792 -41482
rect 36204 -41515 36792 -41499
rect 37222 -41499 37238 -41482
rect 37794 -41482 37996 -41465
rect 38054 -41465 39014 -41418
rect 38054 -41482 38256 -41465
rect 37794 -41499 37810 -41482
rect 37222 -41515 37810 -41499
rect 38240 -41499 38256 -41482
rect 38812 -41482 39014 -41465
rect 39072 -41465 40032 -41418
rect 39072 -41482 39274 -41465
rect 38812 -41499 38828 -41482
rect 38240 -41515 38828 -41499
rect 39258 -41499 39274 -41482
rect 39830 -41482 40032 -41465
rect 40090 -41465 41050 -41418
rect 40090 -41482 40292 -41465
rect 39830 -41499 39846 -41482
rect 39258 -41515 39846 -41499
rect 40276 -41499 40292 -41482
rect 40848 -41482 41050 -41465
rect 41108 -41465 42068 -41418
rect 41108 -41482 41310 -41465
rect 40848 -41499 40864 -41482
rect 40276 -41515 40864 -41499
rect 41294 -41499 41310 -41482
rect 41866 -41482 42068 -41465
rect 42126 -41465 43086 -41418
rect 42126 -41482 42328 -41465
rect 41866 -41499 41882 -41482
rect 41294 -41515 41882 -41499
rect 42312 -41499 42328 -41482
rect 42884 -41482 43086 -41465
rect 43144 -41465 44104 -41418
rect 43144 -41482 43346 -41465
rect 42884 -41499 42900 -41482
rect 42312 -41515 42900 -41499
rect 43330 -41499 43346 -41482
rect 43902 -41482 44104 -41465
rect 44162 -41465 45122 -41418
rect 44162 -41482 44364 -41465
rect 43902 -41499 43918 -41482
rect 43330 -41515 43918 -41499
rect 44348 -41499 44364 -41482
rect 44920 -41482 45122 -41465
rect 45180 -41465 46140 -41418
rect 45180 -41482 45382 -41465
rect 44920 -41499 44936 -41482
rect 44348 -41515 44936 -41499
rect 45366 -41499 45382 -41482
rect 45938 -41482 46140 -41465
rect 46198 -41465 47158 -41418
rect 46198 -41482 46400 -41465
rect 45938 -41499 45954 -41482
rect 45366 -41515 45954 -41499
rect 46384 -41499 46400 -41482
rect 46956 -41482 47158 -41465
rect 47216 -41465 48176 -41418
rect 47216 -41482 47418 -41465
rect 46956 -41499 46972 -41482
rect 46384 -41515 46972 -41499
rect 47402 -41499 47418 -41482
rect 47974 -41482 48176 -41465
rect 47974 -41499 47990 -41482
rect 47402 -41515 47990 -41499
rect 52562 -39599 52814 -39583
rect 52562 -39616 52578 -39599
rect 52488 -39633 52578 -39616
rect 52798 -39616 52814 -39599
rect 53020 -39599 53272 -39583
rect 53020 -39616 53036 -39599
rect 52798 -39633 52888 -39616
rect 52488 -39680 52888 -39633
rect 52946 -39633 53036 -39616
rect 53256 -39616 53272 -39599
rect 53478 -39599 53730 -39583
rect 53478 -39616 53494 -39599
rect 53256 -39633 53346 -39616
rect 52946 -39680 53346 -39633
rect 53404 -39633 53494 -39616
rect 53714 -39616 53730 -39599
rect 53936 -39599 54188 -39583
rect 53936 -39616 53952 -39599
rect 53714 -39633 53804 -39616
rect 53404 -39680 53804 -39633
rect 53862 -39633 53952 -39616
rect 54172 -39616 54188 -39599
rect 54394 -39599 54646 -39583
rect 54394 -39616 54410 -39599
rect 54172 -39633 54262 -39616
rect 53862 -39680 54262 -39633
rect 54320 -39633 54410 -39616
rect 54630 -39616 54646 -39599
rect 54852 -39599 55104 -39583
rect 54852 -39616 54868 -39599
rect 54630 -39633 54720 -39616
rect 54320 -39680 54720 -39633
rect 54778 -39633 54868 -39616
rect 55088 -39616 55104 -39599
rect 55088 -39633 55178 -39616
rect 54778 -39680 55178 -39633
rect 52488 -39927 52888 -39880
rect 52488 -39944 52578 -39927
rect 52562 -39961 52578 -39944
rect 52798 -39944 52888 -39927
rect 52946 -39927 53346 -39880
rect 52946 -39944 53036 -39927
rect 52798 -39961 52814 -39944
rect 52562 -39977 52814 -39961
rect 53020 -39961 53036 -39944
rect 53256 -39944 53346 -39927
rect 53404 -39927 53804 -39880
rect 53404 -39944 53494 -39927
rect 53256 -39961 53272 -39944
rect 53020 -39977 53272 -39961
rect 53478 -39961 53494 -39944
rect 53714 -39944 53804 -39927
rect 53862 -39927 54262 -39880
rect 53862 -39944 53952 -39927
rect 53714 -39961 53730 -39944
rect 53478 -39977 53730 -39961
rect 53936 -39961 53952 -39944
rect 54172 -39944 54262 -39927
rect 54320 -39927 54720 -39880
rect 54320 -39944 54410 -39927
rect 54172 -39961 54188 -39944
rect 53936 -39977 54188 -39961
rect 54394 -39961 54410 -39944
rect 54630 -39944 54720 -39927
rect 54778 -39927 55178 -39880
rect 54778 -39944 54868 -39927
rect 54630 -39961 54646 -39944
rect 54394 -39977 54646 -39961
rect 54852 -39961 54868 -39944
rect 55088 -39944 55178 -39927
rect 55088 -39961 55104 -39944
rect 54852 -39977 55104 -39961
rect 52581 -40482 52713 -40466
rect 52581 -40499 52597 -40482
rect 52547 -40516 52597 -40499
rect 52697 -40499 52713 -40482
rect 52839 -40482 52971 -40466
rect 52839 -40499 52855 -40482
rect 52697 -40516 52747 -40499
rect 52547 -40563 52747 -40516
rect 52805 -40516 52855 -40499
rect 52955 -40499 52971 -40482
rect 53097 -40482 53229 -40466
rect 53097 -40499 53113 -40482
rect 52955 -40516 53005 -40499
rect 52805 -40563 53005 -40516
rect 53063 -40516 53113 -40499
rect 53213 -40499 53229 -40482
rect 53355 -40482 53487 -40466
rect 53355 -40499 53371 -40482
rect 53213 -40516 53263 -40499
rect 53063 -40563 53263 -40516
rect 53321 -40516 53371 -40499
rect 53471 -40499 53487 -40482
rect 53613 -40482 53745 -40466
rect 53613 -40499 53629 -40482
rect 53471 -40516 53521 -40499
rect 53321 -40563 53521 -40516
rect 53579 -40516 53629 -40499
rect 53729 -40499 53745 -40482
rect 53871 -40482 54003 -40466
rect 53871 -40499 53887 -40482
rect 53729 -40516 53779 -40499
rect 53579 -40563 53779 -40516
rect 53837 -40516 53887 -40499
rect 53987 -40499 54003 -40482
rect 54129 -40482 54261 -40466
rect 54129 -40499 54145 -40482
rect 53987 -40516 54037 -40499
rect 53837 -40563 54037 -40516
rect 54095 -40516 54145 -40499
rect 54245 -40499 54261 -40482
rect 54387 -40482 54519 -40466
rect 54387 -40499 54403 -40482
rect 54245 -40516 54295 -40499
rect 54095 -40563 54295 -40516
rect 54353 -40516 54403 -40499
rect 54503 -40499 54519 -40482
rect 54645 -40482 54777 -40466
rect 54645 -40499 54661 -40482
rect 54503 -40516 54553 -40499
rect 54353 -40563 54553 -40516
rect 54611 -40516 54661 -40499
rect 54761 -40499 54777 -40482
rect 54903 -40482 55035 -40466
rect 54903 -40499 54919 -40482
rect 54761 -40516 54811 -40499
rect 54611 -40563 54811 -40516
rect 54869 -40516 54919 -40499
rect 55019 -40499 55035 -40482
rect 55019 -40516 55069 -40499
rect 54869 -40563 55069 -40516
rect 52547 -41010 52747 -40963
rect 52547 -41027 52597 -41010
rect 52581 -41044 52597 -41027
rect 52697 -41027 52747 -41010
rect 52805 -41010 53005 -40963
rect 52805 -41027 52855 -41010
rect 52697 -41044 52713 -41027
rect 52581 -41060 52713 -41044
rect 52839 -41044 52855 -41027
rect 52955 -41027 53005 -41010
rect 53063 -41010 53263 -40963
rect 53063 -41027 53113 -41010
rect 52955 -41044 52971 -41027
rect 52839 -41060 52971 -41044
rect 53097 -41044 53113 -41027
rect 53213 -41027 53263 -41010
rect 53321 -41010 53521 -40963
rect 53321 -41027 53371 -41010
rect 53213 -41044 53229 -41027
rect 53097 -41060 53229 -41044
rect 53355 -41044 53371 -41027
rect 53471 -41027 53521 -41010
rect 53579 -41010 53779 -40963
rect 53579 -41027 53629 -41010
rect 53471 -41044 53487 -41027
rect 53355 -41060 53487 -41044
rect 53613 -41044 53629 -41027
rect 53729 -41027 53779 -41010
rect 53837 -41010 54037 -40963
rect 53837 -41027 53887 -41010
rect 53729 -41044 53745 -41027
rect 53613 -41060 53745 -41044
rect 53871 -41044 53887 -41027
rect 53987 -41027 54037 -41010
rect 54095 -41010 54295 -40963
rect 54095 -41027 54145 -41010
rect 53987 -41044 54003 -41027
rect 53871 -41060 54003 -41044
rect 54129 -41044 54145 -41027
rect 54245 -41027 54295 -41010
rect 54353 -41010 54553 -40963
rect 54353 -41027 54403 -41010
rect 54245 -41044 54261 -41027
rect 54129 -41060 54261 -41044
rect 54387 -41044 54403 -41027
rect 54503 -41027 54553 -41010
rect 54611 -41010 54811 -40963
rect 54611 -41027 54661 -41010
rect 54503 -41044 54519 -41027
rect 54387 -41060 54519 -41044
rect 54645 -41044 54661 -41027
rect 54761 -41027 54811 -41010
rect 54869 -41010 55069 -40963
rect 54869 -41027 54919 -41010
rect 54761 -41044 54777 -41027
rect 54645 -41060 54777 -41044
rect 54903 -41044 54919 -41027
rect 55019 -41027 55069 -41010
rect 55019 -41044 55035 -41027
rect 54903 -41060 55035 -41044
rect 52581 -41342 52713 -41326
rect 52581 -41359 52597 -41342
rect 52547 -41376 52597 -41359
rect 52697 -41359 52713 -41342
rect 52839 -41342 52971 -41326
rect 52839 -41359 52855 -41342
rect 52697 -41376 52747 -41359
rect 52547 -41423 52747 -41376
rect 52805 -41376 52855 -41359
rect 52955 -41359 52971 -41342
rect 53097 -41342 53229 -41326
rect 53097 -41359 53113 -41342
rect 52955 -41376 53005 -41359
rect 52805 -41423 53005 -41376
rect 53063 -41376 53113 -41359
rect 53213 -41359 53229 -41342
rect 53355 -41342 53487 -41326
rect 53355 -41359 53371 -41342
rect 53213 -41376 53263 -41359
rect 53063 -41423 53263 -41376
rect 53321 -41376 53371 -41359
rect 53471 -41359 53487 -41342
rect 53613 -41342 53745 -41326
rect 53613 -41359 53629 -41342
rect 53471 -41376 53521 -41359
rect 53321 -41423 53521 -41376
rect 53579 -41376 53629 -41359
rect 53729 -41359 53745 -41342
rect 53871 -41342 54003 -41326
rect 53871 -41359 53887 -41342
rect 53729 -41376 53779 -41359
rect 53579 -41423 53779 -41376
rect 53837 -41376 53887 -41359
rect 53987 -41359 54003 -41342
rect 54129 -41342 54261 -41326
rect 54129 -41359 54145 -41342
rect 53987 -41376 54037 -41359
rect 53837 -41423 54037 -41376
rect 54095 -41376 54145 -41359
rect 54245 -41359 54261 -41342
rect 54387 -41342 54519 -41326
rect 54387 -41359 54403 -41342
rect 54245 -41376 54295 -41359
rect 54095 -41423 54295 -41376
rect 54353 -41376 54403 -41359
rect 54503 -41359 54519 -41342
rect 54645 -41342 54777 -41326
rect 54645 -41359 54661 -41342
rect 54503 -41376 54553 -41359
rect 54353 -41423 54553 -41376
rect 54611 -41376 54661 -41359
rect 54761 -41359 54777 -41342
rect 54903 -41342 55035 -41326
rect 54903 -41359 54919 -41342
rect 54761 -41376 54811 -41359
rect 54611 -41423 54811 -41376
rect 54869 -41376 54919 -41359
rect 55019 -41359 55035 -41342
rect 55019 -41376 55069 -41359
rect 54869 -41423 55069 -41376
rect 52547 -41870 52747 -41823
rect 52547 -41887 52597 -41870
rect 52581 -41904 52597 -41887
rect 52697 -41887 52747 -41870
rect 52805 -41870 53005 -41823
rect 52805 -41887 52855 -41870
rect 52697 -41904 52713 -41887
rect 52581 -41920 52713 -41904
rect 52839 -41904 52855 -41887
rect 52955 -41887 53005 -41870
rect 53063 -41870 53263 -41823
rect 53063 -41887 53113 -41870
rect 52955 -41904 52971 -41887
rect 52839 -41920 52971 -41904
rect 53097 -41904 53113 -41887
rect 53213 -41887 53263 -41870
rect 53321 -41870 53521 -41823
rect 53321 -41887 53371 -41870
rect 53213 -41904 53229 -41887
rect 53097 -41920 53229 -41904
rect 53355 -41904 53371 -41887
rect 53471 -41887 53521 -41870
rect 53579 -41870 53779 -41823
rect 53579 -41887 53629 -41870
rect 53471 -41904 53487 -41887
rect 53355 -41920 53487 -41904
rect 53613 -41904 53629 -41887
rect 53729 -41887 53779 -41870
rect 53837 -41870 54037 -41823
rect 53837 -41887 53887 -41870
rect 53729 -41904 53745 -41887
rect 53613 -41920 53745 -41904
rect 53871 -41904 53887 -41887
rect 53987 -41887 54037 -41870
rect 54095 -41870 54295 -41823
rect 54095 -41887 54145 -41870
rect 53987 -41904 54003 -41887
rect 53871 -41920 54003 -41904
rect 54129 -41904 54145 -41887
rect 54245 -41887 54295 -41870
rect 54353 -41870 54553 -41823
rect 54353 -41887 54403 -41870
rect 54245 -41904 54261 -41887
rect 54129 -41920 54261 -41904
rect 54387 -41904 54403 -41887
rect 54503 -41887 54553 -41870
rect 54611 -41870 54811 -41823
rect 54611 -41887 54661 -41870
rect 54503 -41904 54519 -41887
rect 54387 -41920 54519 -41904
rect 54645 -41904 54661 -41887
rect 54761 -41887 54811 -41870
rect 54869 -41870 55069 -41823
rect 54869 -41887 54919 -41870
rect 54761 -41904 54777 -41887
rect 54645 -41920 54777 -41904
rect 54903 -41904 54919 -41887
rect 55019 -41887 55069 -41870
rect 55019 -41904 55035 -41887
rect 54903 -41920 55035 -41904
rect 56150 -39799 56282 -39783
rect 56150 -39816 56166 -39799
rect 56116 -39833 56166 -39816
rect 56266 -39816 56282 -39799
rect 56408 -39799 56540 -39783
rect 56408 -39816 56424 -39799
rect 56266 -39833 56316 -39816
rect 56116 -39880 56316 -39833
rect 56374 -39833 56424 -39816
rect 56524 -39816 56540 -39799
rect 56666 -39799 56798 -39783
rect 56666 -39816 56682 -39799
rect 56524 -39833 56574 -39816
rect 56374 -39880 56574 -39833
rect 56632 -39833 56682 -39816
rect 56782 -39816 56798 -39799
rect 56924 -39799 57056 -39783
rect 56924 -39816 56940 -39799
rect 56782 -39833 56832 -39816
rect 56632 -39880 56832 -39833
rect 56890 -39833 56940 -39816
rect 57040 -39816 57056 -39799
rect 57182 -39799 57314 -39783
rect 57182 -39816 57198 -39799
rect 57040 -39833 57090 -39816
rect 56890 -39880 57090 -39833
rect 57148 -39833 57198 -39816
rect 57298 -39816 57314 -39799
rect 57440 -39799 57572 -39783
rect 57440 -39816 57456 -39799
rect 57298 -39833 57348 -39816
rect 57148 -39880 57348 -39833
rect 57406 -39833 57456 -39816
rect 57556 -39816 57572 -39799
rect 57698 -39799 57830 -39783
rect 57698 -39816 57714 -39799
rect 57556 -39833 57606 -39816
rect 57406 -39880 57606 -39833
rect 57664 -39833 57714 -39816
rect 57814 -39816 57830 -39799
rect 57814 -39833 57864 -39816
rect 57664 -39880 57864 -39833
rect 56116 -40327 56316 -40280
rect 56116 -40344 56166 -40327
rect 56150 -40361 56166 -40344
rect 56266 -40344 56316 -40327
rect 56374 -40327 56574 -40280
rect 56374 -40344 56424 -40327
rect 56266 -40361 56282 -40344
rect 56150 -40377 56282 -40361
rect 56408 -40361 56424 -40344
rect 56524 -40344 56574 -40327
rect 56632 -40327 56832 -40280
rect 56632 -40344 56682 -40327
rect 56524 -40361 56540 -40344
rect 56408 -40377 56540 -40361
rect 56666 -40361 56682 -40344
rect 56782 -40344 56832 -40327
rect 56890 -40327 57090 -40280
rect 56890 -40344 56940 -40327
rect 56782 -40361 56798 -40344
rect 56666 -40377 56798 -40361
rect 56924 -40361 56940 -40344
rect 57040 -40344 57090 -40327
rect 57148 -40327 57348 -40280
rect 57148 -40344 57198 -40327
rect 57040 -40361 57056 -40344
rect 56924 -40377 57056 -40361
rect 57182 -40361 57198 -40344
rect 57298 -40344 57348 -40327
rect 57406 -40327 57606 -40280
rect 57406 -40344 57456 -40327
rect 57298 -40361 57314 -40344
rect 57182 -40377 57314 -40361
rect 57440 -40361 57456 -40344
rect 57556 -40344 57606 -40327
rect 57664 -40327 57864 -40280
rect 57664 -40344 57714 -40327
rect 57556 -40361 57572 -40344
rect 57440 -40377 57572 -40361
rect 57698 -40361 57714 -40344
rect 57814 -40344 57864 -40327
rect 57814 -40361 57830 -40344
rect 57698 -40377 57830 -40361
rect 56150 -40659 56282 -40643
rect 56150 -40676 56166 -40659
rect 56116 -40693 56166 -40676
rect 56266 -40676 56282 -40659
rect 56408 -40659 56540 -40643
rect 56408 -40676 56424 -40659
rect 56266 -40693 56316 -40676
rect 56116 -40740 56316 -40693
rect 56374 -40693 56424 -40676
rect 56524 -40676 56540 -40659
rect 56666 -40659 56798 -40643
rect 56666 -40676 56682 -40659
rect 56524 -40693 56574 -40676
rect 56374 -40740 56574 -40693
rect 56632 -40693 56682 -40676
rect 56782 -40676 56798 -40659
rect 56924 -40659 57056 -40643
rect 56924 -40676 56940 -40659
rect 56782 -40693 56832 -40676
rect 56632 -40740 56832 -40693
rect 56890 -40693 56940 -40676
rect 57040 -40676 57056 -40659
rect 57182 -40659 57314 -40643
rect 57182 -40676 57198 -40659
rect 57040 -40693 57090 -40676
rect 56890 -40740 57090 -40693
rect 57148 -40693 57198 -40676
rect 57298 -40676 57314 -40659
rect 57440 -40659 57572 -40643
rect 57440 -40676 57456 -40659
rect 57298 -40693 57348 -40676
rect 57148 -40740 57348 -40693
rect 57406 -40693 57456 -40676
rect 57556 -40676 57572 -40659
rect 57698 -40659 57830 -40643
rect 57698 -40676 57714 -40659
rect 57556 -40693 57606 -40676
rect 57406 -40740 57606 -40693
rect 57664 -40693 57714 -40676
rect 57814 -40676 57830 -40659
rect 57814 -40693 57864 -40676
rect 57664 -40740 57864 -40693
rect 56116 -41187 56316 -41140
rect 56116 -41204 56166 -41187
rect 56150 -41221 56166 -41204
rect 56266 -41204 56316 -41187
rect 56374 -41187 56574 -41140
rect 56374 -41204 56424 -41187
rect 56266 -41221 56282 -41204
rect 56150 -41237 56282 -41221
rect 56408 -41221 56424 -41204
rect 56524 -41204 56574 -41187
rect 56632 -41187 56832 -41140
rect 56632 -41204 56682 -41187
rect 56524 -41221 56540 -41204
rect 56408 -41237 56540 -41221
rect 56666 -41221 56682 -41204
rect 56782 -41204 56832 -41187
rect 56890 -41187 57090 -41140
rect 56890 -41204 56940 -41187
rect 56782 -41221 56798 -41204
rect 56666 -41237 56798 -41221
rect 56924 -41221 56940 -41204
rect 57040 -41204 57090 -41187
rect 57148 -41187 57348 -41140
rect 57148 -41204 57198 -41187
rect 57040 -41221 57056 -41204
rect 56924 -41237 57056 -41221
rect 57182 -41221 57198 -41204
rect 57298 -41204 57348 -41187
rect 57406 -41187 57606 -41140
rect 57406 -41204 57456 -41187
rect 57298 -41221 57314 -41204
rect 57182 -41237 57314 -41221
rect 57440 -41221 57456 -41204
rect 57556 -41204 57606 -41187
rect 57664 -41187 57864 -41140
rect 57664 -41204 57714 -41187
rect 57556 -41221 57572 -41204
rect 57440 -41237 57572 -41221
rect 57698 -41221 57714 -41204
rect 57814 -41204 57864 -41187
rect 57814 -41221 57830 -41204
rect 57698 -41237 57830 -41221
rect 56224 -41639 56254 -41613
rect 56500 -41639 56530 -41613
rect 56739 -41639 56769 -41613
rect 56823 -41639 56853 -41613
rect 57197 -41639 57227 -41613
rect 57281 -41639 57311 -41613
rect 57520 -41639 57550 -41613
rect 57796 -41639 57826 -41613
rect 56224 -41871 56254 -41839
rect 56500 -41871 56530 -41839
rect 56739 -41871 56769 -41839
rect 56168 -41887 56254 -41871
rect 56168 -41921 56184 -41887
rect 56218 -41921 56254 -41887
rect 56168 -41937 56254 -41921
rect 56444 -41887 56530 -41871
rect 56444 -41921 56460 -41887
rect 56494 -41921 56530 -41887
rect 56444 -41937 56530 -41921
rect 56677 -41887 56769 -41871
rect 56677 -41921 56692 -41887
rect 56726 -41921 56769 -41887
rect 56677 -41937 56769 -41921
rect 56224 -41959 56254 -41937
rect 56500 -41959 56530 -41937
rect 56739 -41959 56769 -41937
rect 56823 -41871 56853 -41839
rect 57197 -41871 57227 -41839
rect 56823 -41887 56911 -41871
rect 56823 -41921 56860 -41887
rect 56894 -41921 56911 -41887
rect 56823 -41937 56911 -41921
rect 57139 -41887 57227 -41871
rect 57139 -41921 57156 -41887
rect 57190 -41921 57227 -41887
rect 57139 -41937 57227 -41921
rect 56823 -41959 56853 -41937
rect 57197 -41959 57227 -41937
rect 57281 -41871 57311 -41839
rect 57520 -41871 57550 -41839
rect 57796 -41871 57826 -41839
rect 57281 -41887 57373 -41871
rect 57281 -41921 57324 -41887
rect 57358 -41921 57373 -41887
rect 57281 -41937 57373 -41921
rect 57520 -41887 57606 -41871
rect 57520 -41921 57556 -41887
rect 57590 -41921 57606 -41887
rect 57520 -41937 57606 -41921
rect 57796 -41887 57882 -41871
rect 57796 -41921 57832 -41887
rect 57866 -41921 57882 -41887
rect 57796 -41937 57882 -41921
rect 57281 -41959 57311 -41937
rect 57520 -41959 57550 -41937
rect 57796 -41959 57826 -41937
rect 56224 -42115 56254 -42089
rect 56500 -42115 56530 -42089
rect 56739 -42115 56769 -42089
rect 56823 -42115 56853 -42089
rect 57197 -42115 57227 -42089
rect 57281 -42115 57311 -42089
rect 57520 -42115 57550 -42089
rect 57796 -42115 57826 -42089
rect 54386 -42487 54468 -42477
rect 54386 -42537 54402 -42487
rect 54452 -42537 54468 -42487
rect 54386 -42547 54468 -42537
rect 54514 -42487 54596 -42477
rect 54514 -42537 54530 -42487
rect 54580 -42537 54596 -42487
rect 54514 -42547 54596 -42537
rect 54642 -42487 54724 -42477
rect 54642 -42537 54658 -42487
rect 54708 -42537 54724 -42487
rect 54642 -42547 54724 -42537
rect 54770 -42487 54852 -42477
rect 54770 -42537 54786 -42487
rect 54836 -42537 54852 -42487
rect 54770 -42547 54852 -42537
rect 54898 -42487 54980 -42477
rect 54898 -42537 54914 -42487
rect 54964 -42537 54980 -42487
rect 54898 -42547 54980 -42537
rect 55026 -42487 55108 -42477
rect 55026 -42537 55042 -42487
rect 55092 -42537 55108 -42487
rect 55026 -42547 55108 -42537
rect 55154 -42487 55236 -42477
rect 55154 -42537 55170 -42487
rect 55220 -42537 55236 -42487
rect 55154 -42547 55236 -42537
rect 54264 -42594 54334 -42568
rect 54392 -42594 54462 -42547
rect 54520 -42594 54590 -42547
rect 54648 -42594 54718 -42547
rect 54776 -42594 54846 -42547
rect 54904 -42594 54974 -42547
rect 55032 -42594 55102 -42547
rect 55160 -42594 55230 -42547
rect 55288 -42594 55358 -42568
rect 54264 -42839 54334 -42794
rect 54392 -42820 54462 -42794
rect 54520 -42820 54590 -42794
rect 54648 -42820 54718 -42794
rect 54776 -42820 54846 -42794
rect 54904 -42820 54974 -42794
rect 55032 -42820 55102 -42794
rect 55160 -42820 55230 -42794
rect 55288 -42839 55358 -42794
rect 54258 -42849 54340 -42839
rect 54258 -42899 54274 -42849
rect 54324 -42899 54340 -42849
rect 54258 -42909 54340 -42899
rect 55282 -42849 55364 -42839
rect 55282 -42899 55298 -42849
rect 55348 -42899 55364 -42849
rect 55282 -42909 55364 -42899
rect 56059 -42630 56125 -42614
rect 56059 -42664 56075 -42630
rect 56109 -42664 56125 -42630
rect 56059 -42680 56125 -42664
rect 56062 -42702 56122 -42680
rect 56062 -42928 56122 -42902
rect 56726 -42512 56786 -42496
rect 56726 -42552 56736 -42512
rect 56776 -42552 56786 -42512
rect 56608 -42616 56668 -42590
rect 56726 -42616 56786 -42552
rect 56956 -42512 57028 -42502
rect 56956 -42552 56972 -42512
rect 57012 -42552 57028 -42512
rect 56956 -42562 57028 -42552
rect 57074 -42512 57146 -42502
rect 57074 -42552 57090 -42512
rect 57130 -42552 57146 -42512
rect 57074 -42562 57146 -42552
rect 57310 -42512 57382 -42502
rect 57310 -42552 57326 -42512
rect 57366 -42552 57382 -42512
rect 57310 -42562 57382 -42552
rect 56844 -42616 56904 -42590
rect 56962 -42616 57022 -42562
rect 57080 -42616 57140 -42562
rect 57198 -42616 57258 -42590
rect 57316 -42616 57376 -42562
rect 57434 -42616 57494 -42590
rect 56608 -42866 56668 -42816
rect 56726 -42842 56786 -42816
rect 56542 -42876 56668 -42866
rect 56844 -42868 56904 -42816
rect 56962 -42842 57022 -42816
rect 57080 -42842 57140 -42816
rect 57198 -42868 57258 -42816
rect 57316 -42842 57376 -42816
rect 57434 -42866 57494 -42816
rect 56542 -42916 56558 -42876
rect 56598 -42916 56668 -42876
rect 56542 -42926 56668 -42916
rect 56838 -42878 56910 -42868
rect 56838 -42918 56854 -42878
rect 56894 -42918 56910 -42878
rect 56838 -42928 56910 -42918
rect 57192 -42878 57264 -42868
rect 57192 -42918 57208 -42878
rect 57248 -42918 57264 -42878
rect 57192 -42928 57264 -42918
rect 57434 -42876 57562 -42866
rect 57434 -42916 57506 -42876
rect 57546 -42916 57562 -42876
rect 57434 -42926 57562 -42916
rect 10490 -56841 10622 -56825
rect 10490 -56858 10506 -56841
rect 10456 -56875 10506 -56858
rect 10606 -56858 10622 -56841
rect 10748 -56841 10880 -56825
rect 10748 -56858 10764 -56841
rect 10606 -56875 10656 -56858
rect 10456 -56922 10656 -56875
rect 10714 -56875 10764 -56858
rect 10864 -56858 10880 -56841
rect 11006 -56841 11138 -56825
rect 11006 -56858 11022 -56841
rect 10864 -56875 10914 -56858
rect 10714 -56922 10914 -56875
rect 10972 -56875 11022 -56858
rect 11122 -56858 11138 -56841
rect 11264 -56841 11396 -56825
rect 11264 -56858 11280 -56841
rect 11122 -56875 11172 -56858
rect 10972 -56922 11172 -56875
rect 11230 -56875 11280 -56858
rect 11380 -56858 11396 -56841
rect 11522 -56841 11654 -56825
rect 11522 -56858 11538 -56841
rect 11380 -56875 11430 -56858
rect 11230 -56922 11430 -56875
rect 11488 -56875 11538 -56858
rect 11638 -56858 11654 -56841
rect 11780 -56841 11912 -56825
rect 11780 -56858 11796 -56841
rect 11638 -56875 11688 -56858
rect 11488 -56922 11688 -56875
rect 11746 -56875 11796 -56858
rect 11896 -56858 11912 -56841
rect 11896 -56875 11946 -56858
rect 11746 -56922 11946 -56875
rect 10456 -57369 10656 -57322
rect 10456 -57386 10506 -57369
rect 10490 -57403 10506 -57386
rect 10606 -57386 10656 -57369
rect 10714 -57369 10914 -57322
rect 10714 -57386 10764 -57369
rect 10606 -57403 10622 -57386
rect 10490 -57419 10622 -57403
rect 10748 -57403 10764 -57386
rect 10864 -57386 10914 -57369
rect 10972 -57369 11172 -57322
rect 10972 -57386 11022 -57369
rect 10864 -57403 10880 -57386
rect 10748 -57419 10880 -57403
rect 11006 -57403 11022 -57386
rect 11122 -57386 11172 -57369
rect 11230 -57369 11430 -57322
rect 11230 -57386 11280 -57369
rect 11122 -57403 11138 -57386
rect 11006 -57419 11138 -57403
rect 11264 -57403 11280 -57386
rect 11380 -57386 11430 -57369
rect 11488 -57369 11688 -57322
rect 11488 -57386 11538 -57369
rect 11380 -57403 11396 -57386
rect 11264 -57419 11396 -57403
rect 11522 -57403 11538 -57386
rect 11638 -57386 11688 -57369
rect 11746 -57369 11946 -57322
rect 11746 -57386 11796 -57369
rect 11638 -57403 11654 -57386
rect 11522 -57419 11654 -57403
rect 11780 -57403 11796 -57386
rect 11896 -57386 11946 -57369
rect 11896 -57403 11912 -57386
rect 11780 -57419 11912 -57403
rect 12306 -57305 12336 -57279
rect 12306 -57537 12336 -57505
rect 12306 -57553 12392 -57537
rect 12306 -57587 12342 -57553
rect 12376 -57587 12392 -57553
rect 12306 -57603 12392 -57587
rect 12306 -57625 12336 -57603
rect 10490 -57774 10622 -57758
rect 10490 -57791 10506 -57774
rect 10456 -57808 10506 -57791
rect 10606 -57791 10622 -57774
rect 10748 -57774 10880 -57758
rect 10748 -57791 10764 -57774
rect 10606 -57808 10656 -57791
rect 10456 -57846 10656 -57808
rect 10714 -57808 10764 -57791
rect 10864 -57791 10880 -57774
rect 11006 -57774 11138 -57758
rect 11006 -57791 11022 -57774
rect 10864 -57808 10914 -57791
rect 10714 -57846 10914 -57808
rect 10972 -57808 11022 -57791
rect 11122 -57791 11138 -57774
rect 11264 -57774 11396 -57758
rect 11264 -57791 11280 -57774
rect 11122 -57808 11172 -57791
rect 10972 -57846 11172 -57808
rect 11230 -57808 11280 -57791
rect 11380 -57791 11396 -57774
rect 11522 -57774 11654 -57758
rect 11522 -57791 11538 -57774
rect 11380 -57808 11430 -57791
rect 11230 -57846 11430 -57808
rect 11488 -57808 11538 -57791
rect 11638 -57791 11654 -57774
rect 11780 -57774 11912 -57758
rect 11780 -57791 11796 -57774
rect 11638 -57808 11688 -57791
rect 11488 -57846 11688 -57808
rect 11746 -57808 11796 -57791
rect 11896 -57791 11912 -57774
rect 11896 -57808 11946 -57791
rect 11746 -57846 11946 -57808
rect 10456 -58084 10656 -58046
rect 10456 -58101 10506 -58084
rect 10490 -58118 10506 -58101
rect 10606 -58101 10656 -58084
rect 10714 -58084 10914 -58046
rect 10714 -58101 10764 -58084
rect 10606 -58118 10622 -58101
rect 10490 -58134 10622 -58118
rect 10748 -58118 10764 -58101
rect 10864 -58101 10914 -58084
rect 10972 -58084 11172 -58046
rect 10972 -58101 11022 -58084
rect 10864 -58118 10880 -58101
rect 10748 -58134 10880 -58118
rect 11006 -58118 11022 -58101
rect 11122 -58101 11172 -58084
rect 11230 -58084 11430 -58046
rect 11230 -58101 11280 -58084
rect 11122 -58118 11138 -58101
rect 11006 -58134 11138 -58118
rect 11264 -58118 11280 -58101
rect 11380 -58101 11430 -58084
rect 11488 -58084 11688 -58046
rect 11488 -58101 11538 -58084
rect 11380 -58118 11396 -58101
rect 11264 -58134 11396 -58118
rect 11522 -58118 11538 -58101
rect 11638 -58101 11688 -58084
rect 11746 -58084 11946 -58046
rect 11746 -58101 11796 -58084
rect 11638 -58118 11654 -58101
rect 11522 -58134 11654 -58118
rect 11780 -58118 11796 -58101
rect 11896 -58101 11946 -58084
rect 11896 -58118 11912 -58101
rect 11780 -58134 11912 -58118
rect 12306 -57781 12336 -57755
rect 28258 -43942 28846 -43926
rect 28258 -43959 28274 -43942
rect 28072 -43976 28274 -43959
rect 28830 -43959 28846 -43942
rect 29276 -43942 29864 -43926
rect 29276 -43959 29292 -43942
rect 28830 -43976 29032 -43959
rect 28072 -44014 29032 -43976
rect 29090 -43976 29292 -43959
rect 29848 -43959 29864 -43942
rect 30294 -43942 30882 -43926
rect 30294 -43959 30310 -43942
rect 29848 -43976 30050 -43959
rect 29090 -44014 30050 -43976
rect 30108 -43976 30310 -43959
rect 30866 -43959 30882 -43942
rect 31312 -43942 31900 -43926
rect 31312 -43959 31328 -43942
rect 30866 -43976 31068 -43959
rect 30108 -44014 31068 -43976
rect 31126 -43976 31328 -43959
rect 31884 -43959 31900 -43942
rect 32330 -43942 32918 -43926
rect 32330 -43959 32346 -43942
rect 31884 -43976 32086 -43959
rect 31126 -44014 32086 -43976
rect 32144 -43976 32346 -43959
rect 32902 -43959 32918 -43942
rect 33348 -43942 33936 -43926
rect 33348 -43959 33364 -43942
rect 32902 -43976 33104 -43959
rect 32144 -44014 33104 -43976
rect 33162 -43976 33364 -43959
rect 33920 -43959 33936 -43942
rect 34366 -43942 34954 -43926
rect 34366 -43959 34382 -43942
rect 33920 -43976 34122 -43959
rect 33162 -44014 34122 -43976
rect 34180 -43976 34382 -43959
rect 34938 -43959 34954 -43942
rect 35384 -43942 35972 -43926
rect 35384 -43959 35400 -43942
rect 34938 -43976 35140 -43959
rect 34180 -44014 35140 -43976
rect 35198 -43976 35400 -43959
rect 35956 -43959 35972 -43942
rect 36402 -43942 36990 -43926
rect 36402 -43959 36418 -43942
rect 35956 -43976 36158 -43959
rect 35198 -44014 36158 -43976
rect 36216 -43976 36418 -43959
rect 36974 -43959 36990 -43942
rect 37420 -43942 38008 -43926
rect 37420 -43959 37436 -43942
rect 36974 -43976 37176 -43959
rect 36216 -44014 37176 -43976
rect 37234 -43976 37436 -43959
rect 37992 -43959 38008 -43942
rect 38438 -43942 39026 -43926
rect 38438 -43959 38454 -43942
rect 37992 -43976 38194 -43959
rect 37234 -44014 38194 -43976
rect 38252 -43976 38454 -43959
rect 39010 -43959 39026 -43942
rect 39456 -43942 40044 -43926
rect 39456 -43959 39472 -43942
rect 39010 -43976 39212 -43959
rect 38252 -44014 39212 -43976
rect 39270 -43976 39472 -43959
rect 40028 -43959 40044 -43942
rect 40474 -43942 41062 -43926
rect 40474 -43959 40490 -43942
rect 40028 -43976 40230 -43959
rect 39270 -44014 40230 -43976
rect 40288 -43976 40490 -43959
rect 41046 -43959 41062 -43942
rect 41492 -43942 42080 -43926
rect 41492 -43959 41508 -43942
rect 41046 -43976 41248 -43959
rect 40288 -44014 41248 -43976
rect 41306 -43976 41508 -43959
rect 42064 -43959 42080 -43942
rect 42510 -43942 43098 -43926
rect 42510 -43959 42526 -43942
rect 42064 -43976 42266 -43959
rect 41306 -44014 42266 -43976
rect 42324 -43976 42526 -43959
rect 43082 -43959 43098 -43942
rect 43528 -43942 44116 -43926
rect 43528 -43959 43544 -43942
rect 43082 -43976 43284 -43959
rect 42324 -44014 43284 -43976
rect 43342 -43976 43544 -43959
rect 44100 -43959 44116 -43942
rect 44546 -43942 45134 -43926
rect 44546 -43959 44562 -43942
rect 44100 -43976 44302 -43959
rect 43342 -44014 44302 -43976
rect 44360 -43976 44562 -43959
rect 45118 -43959 45134 -43942
rect 45564 -43942 46152 -43926
rect 45564 -43959 45580 -43942
rect 45118 -43976 45320 -43959
rect 44360 -44014 45320 -43976
rect 45378 -43976 45580 -43959
rect 46136 -43959 46152 -43942
rect 46582 -43942 47170 -43926
rect 46582 -43959 46598 -43942
rect 46136 -43976 46338 -43959
rect 45378 -44014 46338 -43976
rect 46396 -43976 46598 -43959
rect 47154 -43959 47170 -43942
rect 47600 -43942 48188 -43926
rect 47600 -43959 47616 -43942
rect 47154 -43976 47356 -43959
rect 46396 -44014 47356 -43976
rect 47414 -43976 47616 -43959
rect 48172 -43959 48188 -43942
rect 48172 -43976 48374 -43959
rect 47414 -44014 48374 -43976
rect 16492 -44418 17080 -44402
rect 16492 -44435 16508 -44418
rect 16306 -44452 16508 -44435
rect 17064 -44435 17080 -44418
rect 17510 -44418 18098 -44402
rect 17510 -44435 17526 -44418
rect 17064 -44452 17266 -44435
rect 16306 -44490 17266 -44452
rect 17324 -44452 17526 -44435
rect 18082 -44435 18098 -44418
rect 18528 -44418 19116 -44402
rect 18528 -44435 18544 -44418
rect 18082 -44452 18284 -44435
rect 17324 -44490 18284 -44452
rect 18342 -44452 18544 -44435
rect 19100 -44435 19116 -44418
rect 19546 -44418 20134 -44402
rect 19546 -44435 19562 -44418
rect 19100 -44452 19302 -44435
rect 18342 -44490 19302 -44452
rect 19360 -44452 19562 -44435
rect 20118 -44435 20134 -44418
rect 20564 -44418 21152 -44402
rect 20564 -44435 20580 -44418
rect 20118 -44452 20320 -44435
rect 19360 -44490 20320 -44452
rect 20378 -44452 20580 -44435
rect 21136 -44435 21152 -44418
rect 21582 -44418 22170 -44402
rect 21582 -44435 21598 -44418
rect 21136 -44452 21338 -44435
rect 20378 -44490 21338 -44452
rect 21396 -44452 21598 -44435
rect 22154 -44435 22170 -44418
rect 22600 -44418 23188 -44402
rect 22600 -44435 22616 -44418
rect 22154 -44452 22356 -44435
rect 21396 -44490 22356 -44452
rect 22414 -44452 22616 -44435
rect 23172 -44435 23188 -44418
rect 23618 -44418 24206 -44402
rect 23618 -44435 23634 -44418
rect 23172 -44452 23374 -44435
rect 22414 -44490 23374 -44452
rect 23432 -44452 23634 -44435
rect 24190 -44435 24206 -44418
rect 24636 -44418 25224 -44402
rect 24636 -44435 24652 -44418
rect 24190 -44452 24392 -44435
rect 23432 -44490 24392 -44452
rect 24450 -44452 24652 -44435
rect 25208 -44435 25224 -44418
rect 25208 -44452 25410 -44435
rect 24450 -44490 25410 -44452
rect 28072 -44652 29032 -44614
rect 28072 -44669 28274 -44652
rect 28258 -44686 28274 -44669
rect 28830 -44669 29032 -44652
rect 29090 -44652 30050 -44614
rect 29090 -44669 29292 -44652
rect 28830 -44686 28846 -44669
rect 28258 -44702 28846 -44686
rect 29276 -44686 29292 -44669
rect 29848 -44669 30050 -44652
rect 30108 -44652 31068 -44614
rect 30108 -44669 30310 -44652
rect 29848 -44686 29864 -44669
rect 29276 -44702 29864 -44686
rect 30294 -44686 30310 -44669
rect 30866 -44669 31068 -44652
rect 31126 -44652 32086 -44614
rect 31126 -44669 31328 -44652
rect 30866 -44686 30882 -44669
rect 30294 -44702 30882 -44686
rect 31312 -44686 31328 -44669
rect 31884 -44669 32086 -44652
rect 32144 -44652 33104 -44614
rect 32144 -44669 32346 -44652
rect 31884 -44686 31900 -44669
rect 31312 -44702 31900 -44686
rect 32330 -44686 32346 -44669
rect 32902 -44669 33104 -44652
rect 33162 -44652 34122 -44614
rect 33162 -44669 33364 -44652
rect 32902 -44686 32918 -44669
rect 32330 -44702 32918 -44686
rect 33348 -44686 33364 -44669
rect 33920 -44669 34122 -44652
rect 34180 -44652 35140 -44614
rect 34180 -44669 34382 -44652
rect 33920 -44686 33936 -44669
rect 33348 -44702 33936 -44686
rect 34366 -44686 34382 -44669
rect 34938 -44669 35140 -44652
rect 35198 -44652 36158 -44614
rect 35198 -44669 35400 -44652
rect 34938 -44686 34954 -44669
rect 34366 -44702 34954 -44686
rect 35384 -44686 35400 -44669
rect 35956 -44669 36158 -44652
rect 36216 -44652 37176 -44614
rect 36216 -44669 36418 -44652
rect 35956 -44686 35972 -44669
rect 35384 -44702 35972 -44686
rect 36402 -44686 36418 -44669
rect 36974 -44669 37176 -44652
rect 37234 -44652 38194 -44614
rect 37234 -44669 37436 -44652
rect 36974 -44686 36990 -44669
rect 36402 -44702 36990 -44686
rect 37420 -44686 37436 -44669
rect 37992 -44669 38194 -44652
rect 38252 -44652 39212 -44614
rect 38252 -44669 38454 -44652
rect 37992 -44686 38008 -44669
rect 37420 -44702 38008 -44686
rect 38438 -44686 38454 -44669
rect 39010 -44669 39212 -44652
rect 39270 -44652 40230 -44614
rect 39270 -44669 39472 -44652
rect 39010 -44686 39026 -44669
rect 38438 -44702 39026 -44686
rect 39456 -44686 39472 -44669
rect 40028 -44669 40230 -44652
rect 40288 -44652 41248 -44614
rect 40288 -44669 40490 -44652
rect 40028 -44686 40044 -44669
rect 39456 -44702 40044 -44686
rect 40474 -44686 40490 -44669
rect 41046 -44669 41248 -44652
rect 41306 -44652 42266 -44614
rect 41306 -44669 41508 -44652
rect 41046 -44686 41062 -44669
rect 40474 -44702 41062 -44686
rect 41492 -44686 41508 -44669
rect 42064 -44669 42266 -44652
rect 42324 -44652 43284 -44614
rect 42324 -44669 42526 -44652
rect 42064 -44686 42080 -44669
rect 41492 -44702 42080 -44686
rect 42510 -44686 42526 -44669
rect 43082 -44669 43284 -44652
rect 43342 -44652 44302 -44614
rect 43342 -44669 43544 -44652
rect 43082 -44686 43098 -44669
rect 42510 -44702 43098 -44686
rect 43528 -44686 43544 -44669
rect 44100 -44669 44302 -44652
rect 44360 -44652 45320 -44614
rect 44360 -44669 44562 -44652
rect 44100 -44686 44116 -44669
rect 43528 -44702 44116 -44686
rect 44546 -44686 44562 -44669
rect 45118 -44669 45320 -44652
rect 45378 -44652 46338 -44614
rect 45378 -44669 45580 -44652
rect 45118 -44686 45134 -44669
rect 44546 -44702 45134 -44686
rect 45564 -44686 45580 -44669
rect 46136 -44669 46338 -44652
rect 46396 -44652 47356 -44614
rect 46396 -44669 46598 -44652
rect 46136 -44686 46152 -44669
rect 45564 -44702 46152 -44686
rect 46582 -44686 46598 -44669
rect 47154 -44669 47356 -44652
rect 47414 -44652 48374 -44614
rect 47414 -44669 47616 -44652
rect 47154 -44686 47170 -44669
rect 46582 -44702 47170 -44686
rect 47600 -44686 47616 -44669
rect 48172 -44669 48374 -44652
rect 48172 -44686 48188 -44669
rect 47600 -44702 48188 -44686
rect 28258 -44760 28846 -44744
rect 28258 -44777 28274 -44760
rect 28072 -44794 28274 -44777
rect 28830 -44777 28846 -44760
rect 29276 -44760 29864 -44744
rect 29276 -44777 29292 -44760
rect 28830 -44794 29032 -44777
rect 28072 -44832 29032 -44794
rect 29090 -44794 29292 -44777
rect 29848 -44777 29864 -44760
rect 30294 -44760 30882 -44744
rect 30294 -44777 30310 -44760
rect 29848 -44794 30050 -44777
rect 29090 -44832 30050 -44794
rect 30108 -44794 30310 -44777
rect 30866 -44777 30882 -44760
rect 31312 -44760 31900 -44744
rect 31312 -44777 31328 -44760
rect 30866 -44794 31068 -44777
rect 30108 -44832 31068 -44794
rect 31126 -44794 31328 -44777
rect 31884 -44777 31900 -44760
rect 32330 -44760 32918 -44744
rect 32330 -44777 32346 -44760
rect 31884 -44794 32086 -44777
rect 31126 -44832 32086 -44794
rect 32144 -44794 32346 -44777
rect 32902 -44777 32918 -44760
rect 33348 -44760 33936 -44744
rect 33348 -44777 33364 -44760
rect 32902 -44794 33104 -44777
rect 32144 -44832 33104 -44794
rect 33162 -44794 33364 -44777
rect 33920 -44777 33936 -44760
rect 34366 -44760 34954 -44744
rect 34366 -44777 34382 -44760
rect 33920 -44794 34122 -44777
rect 33162 -44832 34122 -44794
rect 34180 -44794 34382 -44777
rect 34938 -44777 34954 -44760
rect 35384 -44760 35972 -44744
rect 35384 -44777 35400 -44760
rect 34938 -44794 35140 -44777
rect 34180 -44832 35140 -44794
rect 35198 -44794 35400 -44777
rect 35956 -44777 35972 -44760
rect 36402 -44760 36990 -44744
rect 36402 -44777 36418 -44760
rect 35956 -44794 36158 -44777
rect 35198 -44832 36158 -44794
rect 36216 -44794 36418 -44777
rect 36974 -44777 36990 -44760
rect 37420 -44760 38008 -44744
rect 37420 -44777 37436 -44760
rect 36974 -44794 37176 -44777
rect 36216 -44832 37176 -44794
rect 37234 -44794 37436 -44777
rect 37992 -44777 38008 -44760
rect 38438 -44760 39026 -44744
rect 38438 -44777 38454 -44760
rect 37992 -44794 38194 -44777
rect 37234 -44832 38194 -44794
rect 38252 -44794 38454 -44777
rect 39010 -44777 39026 -44760
rect 39456 -44760 40044 -44744
rect 39456 -44777 39472 -44760
rect 39010 -44794 39212 -44777
rect 38252 -44832 39212 -44794
rect 39270 -44794 39472 -44777
rect 40028 -44777 40044 -44760
rect 40474 -44760 41062 -44744
rect 40474 -44777 40490 -44760
rect 40028 -44794 40230 -44777
rect 39270 -44832 40230 -44794
rect 40288 -44794 40490 -44777
rect 41046 -44777 41062 -44760
rect 41492 -44760 42080 -44744
rect 41492 -44777 41508 -44760
rect 41046 -44794 41248 -44777
rect 40288 -44832 41248 -44794
rect 41306 -44794 41508 -44777
rect 42064 -44777 42080 -44760
rect 42510 -44760 43098 -44744
rect 42510 -44777 42526 -44760
rect 42064 -44794 42266 -44777
rect 41306 -44832 42266 -44794
rect 42324 -44794 42526 -44777
rect 43082 -44777 43098 -44760
rect 43528 -44760 44116 -44744
rect 43528 -44777 43544 -44760
rect 43082 -44794 43284 -44777
rect 42324 -44832 43284 -44794
rect 43342 -44794 43544 -44777
rect 44100 -44777 44116 -44760
rect 44546 -44760 45134 -44744
rect 44546 -44777 44562 -44760
rect 44100 -44794 44302 -44777
rect 43342 -44832 44302 -44794
rect 44360 -44794 44562 -44777
rect 45118 -44777 45134 -44760
rect 45564 -44760 46152 -44744
rect 45564 -44777 45580 -44760
rect 45118 -44794 45320 -44777
rect 44360 -44832 45320 -44794
rect 45378 -44794 45580 -44777
rect 46136 -44777 46152 -44760
rect 46582 -44760 47170 -44744
rect 46582 -44777 46598 -44760
rect 46136 -44794 46338 -44777
rect 45378 -44832 46338 -44794
rect 46396 -44794 46598 -44777
rect 47154 -44777 47170 -44760
rect 47600 -44760 48188 -44744
rect 47600 -44777 47616 -44760
rect 47154 -44794 47356 -44777
rect 46396 -44832 47356 -44794
rect 47414 -44794 47616 -44777
rect 48172 -44777 48188 -44760
rect 48172 -44794 48374 -44777
rect 47414 -44832 48374 -44794
rect 16306 -45128 17266 -45090
rect 16306 -45145 16508 -45128
rect 16492 -45162 16508 -45145
rect 17064 -45145 17266 -45128
rect 17324 -45128 18284 -45090
rect 17324 -45145 17526 -45128
rect 17064 -45162 17080 -45145
rect 16492 -45178 17080 -45162
rect 17510 -45162 17526 -45145
rect 18082 -45145 18284 -45128
rect 18342 -45128 19302 -45090
rect 18342 -45145 18544 -45128
rect 18082 -45162 18098 -45145
rect 17510 -45178 18098 -45162
rect 16492 -45236 17080 -45220
rect 16492 -45253 16508 -45236
rect 16306 -45270 16508 -45253
rect 17064 -45253 17080 -45236
rect 18528 -45162 18544 -45145
rect 19100 -45145 19302 -45128
rect 19360 -45128 20320 -45090
rect 19360 -45145 19562 -45128
rect 19100 -45162 19116 -45145
rect 18528 -45178 19116 -45162
rect 17510 -45236 18098 -45220
rect 17510 -45253 17526 -45236
rect 17064 -45270 17266 -45253
rect 16306 -45308 17266 -45270
rect 17324 -45270 17526 -45253
rect 18082 -45253 18098 -45236
rect 19546 -45162 19562 -45145
rect 20118 -45145 20320 -45128
rect 20378 -45128 21338 -45090
rect 20378 -45145 20580 -45128
rect 20118 -45162 20134 -45145
rect 19546 -45178 20134 -45162
rect 18528 -45236 19116 -45220
rect 18528 -45253 18544 -45236
rect 18082 -45270 18284 -45253
rect 17324 -45308 18284 -45270
rect 18342 -45270 18544 -45253
rect 19100 -45253 19116 -45236
rect 20564 -45162 20580 -45145
rect 21136 -45145 21338 -45128
rect 21396 -45128 22356 -45090
rect 21396 -45145 21598 -45128
rect 21136 -45162 21152 -45145
rect 20564 -45178 21152 -45162
rect 19546 -45236 20134 -45220
rect 19546 -45253 19562 -45236
rect 19100 -45270 19302 -45253
rect 18342 -45308 19302 -45270
rect 19360 -45270 19562 -45253
rect 20118 -45253 20134 -45236
rect 21582 -45162 21598 -45145
rect 22154 -45145 22356 -45128
rect 22414 -45128 23374 -45090
rect 22414 -45145 22616 -45128
rect 22154 -45162 22170 -45145
rect 21582 -45178 22170 -45162
rect 20564 -45236 21152 -45220
rect 20564 -45253 20580 -45236
rect 20118 -45270 20320 -45253
rect 19360 -45308 20320 -45270
rect 20378 -45270 20580 -45253
rect 21136 -45253 21152 -45236
rect 22600 -45162 22616 -45145
rect 23172 -45145 23374 -45128
rect 23432 -45128 24392 -45090
rect 23432 -45145 23634 -45128
rect 23172 -45162 23188 -45145
rect 22600 -45178 23188 -45162
rect 21582 -45236 22170 -45220
rect 21582 -45253 21598 -45236
rect 21136 -45270 21338 -45253
rect 20378 -45308 21338 -45270
rect 21396 -45270 21598 -45253
rect 22154 -45253 22170 -45236
rect 23618 -45162 23634 -45145
rect 24190 -45145 24392 -45128
rect 24450 -45128 25410 -45090
rect 24450 -45145 24652 -45128
rect 24190 -45162 24206 -45145
rect 23618 -45178 24206 -45162
rect 22600 -45236 23188 -45220
rect 22600 -45253 22616 -45236
rect 22154 -45270 22356 -45253
rect 21396 -45308 22356 -45270
rect 22414 -45270 22616 -45253
rect 23172 -45253 23188 -45236
rect 24636 -45162 24652 -45145
rect 25208 -45145 25410 -45128
rect 25208 -45162 25224 -45145
rect 24636 -45178 25224 -45162
rect 23618 -45236 24206 -45220
rect 23618 -45253 23634 -45236
rect 23172 -45270 23374 -45253
rect 22414 -45308 23374 -45270
rect 23432 -45270 23634 -45253
rect 24190 -45253 24206 -45236
rect 24636 -45236 25224 -45220
rect 24636 -45253 24652 -45236
rect 24190 -45270 24392 -45253
rect 23432 -45308 24392 -45270
rect 24450 -45270 24652 -45253
rect 25208 -45253 25224 -45236
rect 25208 -45270 25410 -45253
rect 24450 -45308 25410 -45270
rect 28072 -45470 29032 -45432
rect 28072 -45487 28274 -45470
rect 28258 -45504 28274 -45487
rect 28830 -45487 29032 -45470
rect 29090 -45470 30050 -45432
rect 29090 -45487 29292 -45470
rect 28830 -45504 28846 -45487
rect 28258 -45520 28846 -45504
rect 29276 -45504 29292 -45487
rect 29848 -45487 30050 -45470
rect 30108 -45470 31068 -45432
rect 30108 -45487 30310 -45470
rect 29848 -45504 29864 -45487
rect 29276 -45520 29864 -45504
rect 30294 -45504 30310 -45487
rect 30866 -45487 31068 -45470
rect 31126 -45470 32086 -45432
rect 31126 -45487 31328 -45470
rect 30866 -45504 30882 -45487
rect 30294 -45520 30882 -45504
rect 31312 -45504 31328 -45487
rect 31884 -45487 32086 -45470
rect 32144 -45470 33104 -45432
rect 32144 -45487 32346 -45470
rect 31884 -45504 31900 -45487
rect 31312 -45520 31900 -45504
rect 32330 -45504 32346 -45487
rect 32902 -45487 33104 -45470
rect 33162 -45470 34122 -45432
rect 33162 -45487 33364 -45470
rect 32902 -45504 32918 -45487
rect 32330 -45520 32918 -45504
rect 33348 -45504 33364 -45487
rect 33920 -45487 34122 -45470
rect 34180 -45470 35140 -45432
rect 34180 -45487 34382 -45470
rect 33920 -45504 33936 -45487
rect 33348 -45520 33936 -45504
rect 34366 -45504 34382 -45487
rect 34938 -45487 35140 -45470
rect 35198 -45470 36158 -45432
rect 35198 -45487 35400 -45470
rect 34938 -45504 34954 -45487
rect 34366 -45520 34954 -45504
rect 35384 -45504 35400 -45487
rect 35956 -45487 36158 -45470
rect 36216 -45470 37176 -45432
rect 36216 -45487 36418 -45470
rect 35956 -45504 35972 -45487
rect 35384 -45520 35972 -45504
rect 36402 -45504 36418 -45487
rect 36974 -45487 37176 -45470
rect 37234 -45470 38194 -45432
rect 37234 -45487 37436 -45470
rect 36974 -45504 36990 -45487
rect 36402 -45520 36990 -45504
rect 37420 -45504 37436 -45487
rect 37992 -45487 38194 -45470
rect 38252 -45470 39212 -45432
rect 38252 -45487 38454 -45470
rect 37992 -45504 38008 -45487
rect 37420 -45520 38008 -45504
rect 38438 -45504 38454 -45487
rect 39010 -45487 39212 -45470
rect 39270 -45470 40230 -45432
rect 39270 -45487 39472 -45470
rect 39010 -45504 39026 -45487
rect 38438 -45520 39026 -45504
rect 39456 -45504 39472 -45487
rect 40028 -45487 40230 -45470
rect 40288 -45470 41248 -45432
rect 40288 -45487 40490 -45470
rect 40028 -45504 40044 -45487
rect 39456 -45520 40044 -45504
rect 40474 -45504 40490 -45487
rect 41046 -45487 41248 -45470
rect 41306 -45470 42266 -45432
rect 41306 -45487 41508 -45470
rect 41046 -45504 41062 -45487
rect 40474 -45520 41062 -45504
rect 41492 -45504 41508 -45487
rect 42064 -45487 42266 -45470
rect 42324 -45470 43284 -45432
rect 42324 -45487 42526 -45470
rect 42064 -45504 42080 -45487
rect 41492 -45520 42080 -45504
rect 42510 -45504 42526 -45487
rect 43082 -45487 43284 -45470
rect 43342 -45470 44302 -45432
rect 43342 -45487 43544 -45470
rect 43082 -45504 43098 -45487
rect 42510 -45520 43098 -45504
rect 43528 -45504 43544 -45487
rect 44100 -45487 44302 -45470
rect 44360 -45470 45320 -45432
rect 44360 -45487 44562 -45470
rect 44100 -45504 44116 -45487
rect 43528 -45520 44116 -45504
rect 44546 -45504 44562 -45487
rect 45118 -45487 45320 -45470
rect 45378 -45470 46338 -45432
rect 45378 -45487 45580 -45470
rect 45118 -45504 45134 -45487
rect 44546 -45520 45134 -45504
rect 45564 -45504 45580 -45487
rect 46136 -45487 46338 -45470
rect 46396 -45470 47356 -45432
rect 46396 -45487 46598 -45470
rect 46136 -45504 46152 -45487
rect 45564 -45520 46152 -45504
rect 46582 -45504 46598 -45487
rect 47154 -45487 47356 -45470
rect 47414 -45470 48374 -45432
rect 47414 -45487 47616 -45470
rect 47154 -45504 47170 -45487
rect 46582 -45520 47170 -45504
rect 47600 -45504 47616 -45487
rect 48172 -45487 48374 -45470
rect 48172 -45504 48188 -45487
rect 47600 -45520 48188 -45504
rect 16306 -45946 17266 -45908
rect 16306 -45963 16508 -45946
rect 16492 -45980 16508 -45963
rect 17064 -45963 17266 -45946
rect 17324 -45946 18284 -45908
rect 17324 -45963 17526 -45946
rect 17064 -45980 17080 -45963
rect 16492 -45996 17080 -45980
rect 17510 -45980 17526 -45963
rect 18082 -45963 18284 -45946
rect 18342 -45946 19302 -45908
rect 18342 -45963 18544 -45946
rect 18082 -45980 18098 -45963
rect 17510 -45996 18098 -45980
rect 16492 -46054 17080 -46038
rect 16492 -46071 16508 -46054
rect 16306 -46088 16508 -46071
rect 17064 -46071 17080 -46054
rect 18528 -45980 18544 -45963
rect 19100 -45963 19302 -45946
rect 19360 -45946 20320 -45908
rect 19360 -45963 19562 -45946
rect 19100 -45980 19116 -45963
rect 18528 -45996 19116 -45980
rect 17510 -46054 18098 -46038
rect 17510 -46071 17526 -46054
rect 17064 -46088 17266 -46071
rect 16306 -46126 17266 -46088
rect 17324 -46088 17526 -46071
rect 18082 -46071 18098 -46054
rect 19546 -45980 19562 -45963
rect 20118 -45963 20320 -45946
rect 20378 -45946 21338 -45908
rect 20378 -45963 20580 -45946
rect 20118 -45980 20134 -45963
rect 19546 -45996 20134 -45980
rect 18528 -46054 19116 -46038
rect 18528 -46071 18544 -46054
rect 18082 -46088 18284 -46071
rect 17324 -46126 18284 -46088
rect 18342 -46088 18544 -46071
rect 19100 -46071 19116 -46054
rect 20564 -45980 20580 -45963
rect 21136 -45963 21338 -45946
rect 21396 -45946 22356 -45908
rect 21396 -45963 21598 -45946
rect 21136 -45980 21152 -45963
rect 20564 -45996 21152 -45980
rect 19546 -46054 20134 -46038
rect 19546 -46071 19562 -46054
rect 19100 -46088 19302 -46071
rect 18342 -46126 19302 -46088
rect 19360 -46088 19562 -46071
rect 20118 -46071 20134 -46054
rect 21582 -45980 21598 -45963
rect 22154 -45963 22356 -45946
rect 22414 -45946 23374 -45908
rect 22414 -45963 22616 -45946
rect 22154 -45980 22170 -45963
rect 21582 -45996 22170 -45980
rect 20564 -46054 21152 -46038
rect 20564 -46071 20580 -46054
rect 20118 -46088 20320 -46071
rect 19360 -46126 20320 -46088
rect 20378 -46088 20580 -46071
rect 21136 -46071 21152 -46054
rect 22600 -45980 22616 -45963
rect 23172 -45963 23374 -45946
rect 23432 -45946 24392 -45908
rect 23432 -45963 23634 -45946
rect 23172 -45980 23188 -45963
rect 22600 -45996 23188 -45980
rect 21582 -46054 22170 -46038
rect 21582 -46071 21598 -46054
rect 21136 -46088 21338 -46071
rect 20378 -46126 21338 -46088
rect 21396 -46088 21598 -46071
rect 22154 -46071 22170 -46054
rect 23618 -45980 23634 -45963
rect 24190 -45963 24392 -45946
rect 24450 -45946 25410 -45908
rect 24450 -45963 24652 -45946
rect 24190 -45980 24206 -45963
rect 23618 -45996 24206 -45980
rect 22600 -46054 23188 -46038
rect 22600 -46071 22616 -46054
rect 22154 -46088 22356 -46071
rect 21396 -46126 22356 -46088
rect 22414 -46088 22616 -46071
rect 23172 -46071 23188 -46054
rect 24636 -45980 24652 -45963
rect 25208 -45963 25410 -45946
rect 25208 -45980 25224 -45963
rect 24636 -45996 25224 -45980
rect 23618 -46054 24206 -46038
rect 23618 -46071 23634 -46054
rect 23172 -46088 23374 -46071
rect 22414 -46126 23374 -46088
rect 23432 -46088 23634 -46071
rect 24190 -46071 24206 -46054
rect 24636 -46054 25224 -46038
rect 24636 -46071 24652 -46054
rect 24190 -46088 24392 -46071
rect 23432 -46126 24392 -46088
rect 24450 -46088 24652 -46071
rect 25208 -46071 25224 -46054
rect 25208 -46088 25410 -46071
rect 24450 -46126 25410 -46088
rect 28258 -46138 28846 -46122
rect 28258 -46155 28274 -46138
rect 28072 -46172 28274 -46155
rect 28830 -46155 28846 -46138
rect 29276 -46138 29864 -46122
rect 29276 -46155 29292 -46138
rect 28830 -46172 29032 -46155
rect 28072 -46210 29032 -46172
rect 29090 -46172 29292 -46155
rect 29848 -46155 29864 -46138
rect 30294 -46138 30882 -46122
rect 30294 -46155 30310 -46138
rect 29848 -46172 30050 -46155
rect 29090 -46210 30050 -46172
rect 30108 -46172 30310 -46155
rect 30866 -46155 30882 -46138
rect 31312 -46138 31900 -46122
rect 31312 -46155 31328 -46138
rect 30866 -46172 31068 -46155
rect 30108 -46210 31068 -46172
rect 31126 -46172 31328 -46155
rect 31884 -46155 31900 -46138
rect 32330 -46138 32918 -46122
rect 32330 -46155 32346 -46138
rect 31884 -46172 32086 -46155
rect 31126 -46210 32086 -46172
rect 32144 -46172 32346 -46155
rect 32902 -46155 32918 -46138
rect 33348 -46138 33936 -46122
rect 33348 -46155 33364 -46138
rect 32902 -46172 33104 -46155
rect 32144 -46210 33104 -46172
rect 33162 -46172 33364 -46155
rect 33920 -46155 33936 -46138
rect 34366 -46138 34954 -46122
rect 34366 -46155 34382 -46138
rect 33920 -46172 34122 -46155
rect 33162 -46210 34122 -46172
rect 34180 -46172 34382 -46155
rect 34938 -46155 34954 -46138
rect 35384 -46138 35972 -46122
rect 35384 -46155 35400 -46138
rect 34938 -46172 35140 -46155
rect 34180 -46210 35140 -46172
rect 35198 -46172 35400 -46155
rect 35956 -46155 35972 -46138
rect 36402 -46138 36990 -46122
rect 36402 -46155 36418 -46138
rect 35956 -46172 36158 -46155
rect 35198 -46210 36158 -46172
rect 36216 -46172 36418 -46155
rect 36974 -46155 36990 -46138
rect 37420 -46138 38008 -46122
rect 37420 -46155 37436 -46138
rect 36974 -46172 37176 -46155
rect 36216 -46210 37176 -46172
rect 37234 -46172 37436 -46155
rect 37992 -46155 38008 -46138
rect 38438 -46138 39026 -46122
rect 38438 -46155 38454 -46138
rect 37992 -46172 38194 -46155
rect 37234 -46210 38194 -46172
rect 38252 -46172 38454 -46155
rect 39010 -46155 39026 -46138
rect 39456 -46138 40044 -46122
rect 39456 -46155 39472 -46138
rect 39010 -46172 39212 -46155
rect 38252 -46210 39212 -46172
rect 39270 -46172 39472 -46155
rect 40028 -46155 40044 -46138
rect 40474 -46138 41062 -46122
rect 40474 -46155 40490 -46138
rect 40028 -46172 40230 -46155
rect 39270 -46210 40230 -46172
rect 40288 -46172 40490 -46155
rect 41046 -46155 41062 -46138
rect 41492 -46138 42080 -46122
rect 41492 -46155 41508 -46138
rect 41046 -46172 41248 -46155
rect 40288 -46210 41248 -46172
rect 41306 -46172 41508 -46155
rect 42064 -46155 42080 -46138
rect 42510 -46138 43098 -46122
rect 42510 -46155 42526 -46138
rect 42064 -46172 42266 -46155
rect 41306 -46210 42266 -46172
rect 42324 -46172 42526 -46155
rect 43082 -46155 43098 -46138
rect 43528 -46138 44116 -46122
rect 43528 -46155 43544 -46138
rect 43082 -46172 43284 -46155
rect 42324 -46210 43284 -46172
rect 43342 -46172 43544 -46155
rect 44100 -46155 44116 -46138
rect 44546 -46138 45134 -46122
rect 44546 -46155 44562 -46138
rect 44100 -46172 44302 -46155
rect 43342 -46210 44302 -46172
rect 44360 -46172 44562 -46155
rect 45118 -46155 45134 -46138
rect 45564 -46138 46152 -46122
rect 45564 -46155 45580 -46138
rect 45118 -46172 45320 -46155
rect 44360 -46210 45320 -46172
rect 45378 -46172 45580 -46155
rect 46136 -46155 46152 -46138
rect 46582 -46138 47170 -46122
rect 46582 -46155 46598 -46138
rect 46136 -46172 46338 -46155
rect 45378 -46210 46338 -46172
rect 46396 -46172 46598 -46155
rect 47154 -46155 47170 -46138
rect 47600 -46138 48188 -46122
rect 47600 -46155 47616 -46138
rect 47154 -46172 47356 -46155
rect 46396 -46210 47356 -46172
rect 47414 -46172 47616 -46155
rect 48172 -46155 48188 -46138
rect 48172 -46172 48374 -46155
rect 47414 -46210 48374 -46172
rect 16306 -46764 17266 -46726
rect 16306 -46781 16508 -46764
rect 16492 -46798 16508 -46781
rect 17064 -46781 17266 -46764
rect 17324 -46764 18284 -46726
rect 17324 -46781 17526 -46764
rect 17064 -46798 17080 -46781
rect 16492 -46814 17080 -46798
rect 17510 -46798 17526 -46781
rect 18082 -46781 18284 -46764
rect 18342 -46764 19302 -46726
rect 18342 -46781 18544 -46764
rect 18082 -46798 18098 -46781
rect 17510 -46814 18098 -46798
rect 16492 -46872 17080 -46856
rect 16492 -46889 16508 -46872
rect 16306 -46906 16508 -46889
rect 17064 -46889 17080 -46872
rect 18528 -46798 18544 -46781
rect 19100 -46781 19302 -46764
rect 19360 -46764 20320 -46726
rect 19360 -46781 19562 -46764
rect 19100 -46798 19116 -46781
rect 18528 -46814 19116 -46798
rect 17510 -46872 18098 -46856
rect 17510 -46889 17526 -46872
rect 17064 -46906 17266 -46889
rect 16306 -46944 17266 -46906
rect 17324 -46906 17526 -46889
rect 18082 -46889 18098 -46872
rect 19546 -46798 19562 -46781
rect 20118 -46781 20320 -46764
rect 20378 -46764 21338 -46726
rect 20378 -46781 20580 -46764
rect 20118 -46798 20134 -46781
rect 19546 -46814 20134 -46798
rect 18528 -46872 19116 -46856
rect 18528 -46889 18544 -46872
rect 18082 -46906 18284 -46889
rect 17324 -46944 18284 -46906
rect 18342 -46906 18544 -46889
rect 19100 -46889 19116 -46872
rect 20564 -46798 20580 -46781
rect 21136 -46781 21338 -46764
rect 21396 -46764 22356 -46726
rect 21396 -46781 21598 -46764
rect 21136 -46798 21152 -46781
rect 20564 -46814 21152 -46798
rect 19546 -46872 20134 -46856
rect 19546 -46889 19562 -46872
rect 19100 -46906 19302 -46889
rect 18342 -46944 19302 -46906
rect 19360 -46906 19562 -46889
rect 20118 -46889 20134 -46872
rect 21582 -46798 21598 -46781
rect 22154 -46781 22356 -46764
rect 22414 -46764 23374 -46726
rect 22414 -46781 22616 -46764
rect 22154 -46798 22170 -46781
rect 21582 -46814 22170 -46798
rect 20564 -46872 21152 -46856
rect 20564 -46889 20580 -46872
rect 20118 -46906 20320 -46889
rect 19360 -46944 20320 -46906
rect 20378 -46906 20580 -46889
rect 21136 -46889 21152 -46872
rect 22600 -46798 22616 -46781
rect 23172 -46781 23374 -46764
rect 23432 -46764 24392 -46726
rect 23432 -46781 23634 -46764
rect 23172 -46798 23188 -46781
rect 22600 -46814 23188 -46798
rect 21582 -46872 22170 -46856
rect 21582 -46889 21598 -46872
rect 21136 -46906 21338 -46889
rect 20378 -46944 21338 -46906
rect 21396 -46906 21598 -46889
rect 22154 -46889 22170 -46872
rect 23618 -46798 23634 -46781
rect 24190 -46781 24392 -46764
rect 24450 -46764 25410 -46726
rect 24450 -46781 24652 -46764
rect 24190 -46798 24206 -46781
rect 23618 -46814 24206 -46798
rect 22600 -46872 23188 -46856
rect 22600 -46889 22616 -46872
rect 22154 -46906 22356 -46889
rect 21396 -46944 22356 -46906
rect 22414 -46906 22616 -46889
rect 23172 -46889 23188 -46872
rect 24636 -46798 24652 -46781
rect 25208 -46781 25410 -46764
rect 25208 -46798 25224 -46781
rect 24636 -46814 25224 -46798
rect 23618 -46872 24206 -46856
rect 23618 -46889 23634 -46872
rect 23172 -46906 23374 -46889
rect 22414 -46944 23374 -46906
rect 23432 -46906 23634 -46889
rect 24190 -46889 24206 -46872
rect 24636 -46872 25224 -46856
rect 24636 -46889 24652 -46872
rect 24190 -46906 24392 -46889
rect 23432 -46944 24392 -46906
rect 24450 -46906 24652 -46889
rect 25208 -46889 25224 -46872
rect 28072 -46848 29032 -46810
rect 28072 -46865 28274 -46848
rect 28258 -46882 28274 -46865
rect 28830 -46865 29032 -46848
rect 29090 -46848 30050 -46810
rect 29090 -46865 29292 -46848
rect 28830 -46882 28846 -46865
rect 25208 -46906 25410 -46889
rect 28258 -46898 28846 -46882
rect 29276 -46882 29292 -46865
rect 29848 -46865 30050 -46848
rect 30108 -46848 31068 -46810
rect 30108 -46865 30310 -46848
rect 29848 -46882 29864 -46865
rect 29276 -46898 29864 -46882
rect 30294 -46882 30310 -46865
rect 30866 -46865 31068 -46848
rect 31126 -46848 32086 -46810
rect 31126 -46865 31328 -46848
rect 30866 -46882 30882 -46865
rect 30294 -46898 30882 -46882
rect 31312 -46882 31328 -46865
rect 31884 -46865 32086 -46848
rect 32144 -46848 33104 -46810
rect 32144 -46865 32346 -46848
rect 31884 -46882 31900 -46865
rect 31312 -46898 31900 -46882
rect 32330 -46882 32346 -46865
rect 32902 -46865 33104 -46848
rect 33162 -46848 34122 -46810
rect 33162 -46865 33364 -46848
rect 32902 -46882 32918 -46865
rect 32330 -46898 32918 -46882
rect 33348 -46882 33364 -46865
rect 33920 -46865 34122 -46848
rect 34180 -46848 35140 -46810
rect 34180 -46865 34382 -46848
rect 33920 -46882 33936 -46865
rect 33348 -46898 33936 -46882
rect 34366 -46882 34382 -46865
rect 34938 -46865 35140 -46848
rect 35198 -46848 36158 -46810
rect 35198 -46865 35400 -46848
rect 34938 -46882 34954 -46865
rect 34366 -46898 34954 -46882
rect 35384 -46882 35400 -46865
rect 35956 -46865 36158 -46848
rect 36216 -46848 37176 -46810
rect 36216 -46865 36418 -46848
rect 35956 -46882 35972 -46865
rect 35384 -46898 35972 -46882
rect 36402 -46882 36418 -46865
rect 36974 -46865 37176 -46848
rect 37234 -46848 38194 -46810
rect 37234 -46865 37436 -46848
rect 36974 -46882 36990 -46865
rect 36402 -46898 36990 -46882
rect 37420 -46882 37436 -46865
rect 37992 -46865 38194 -46848
rect 38252 -46848 39212 -46810
rect 38252 -46865 38454 -46848
rect 37992 -46882 38008 -46865
rect 37420 -46898 38008 -46882
rect 38438 -46882 38454 -46865
rect 39010 -46865 39212 -46848
rect 39270 -46848 40230 -46810
rect 39270 -46865 39472 -46848
rect 39010 -46882 39026 -46865
rect 38438 -46898 39026 -46882
rect 39456 -46882 39472 -46865
rect 40028 -46865 40230 -46848
rect 40288 -46848 41248 -46810
rect 40288 -46865 40490 -46848
rect 40028 -46882 40044 -46865
rect 39456 -46898 40044 -46882
rect 40474 -46882 40490 -46865
rect 41046 -46865 41248 -46848
rect 41306 -46848 42266 -46810
rect 41306 -46865 41508 -46848
rect 41046 -46882 41062 -46865
rect 40474 -46898 41062 -46882
rect 41492 -46882 41508 -46865
rect 42064 -46865 42266 -46848
rect 42324 -46848 43284 -46810
rect 42324 -46865 42526 -46848
rect 42064 -46882 42080 -46865
rect 41492 -46898 42080 -46882
rect 42510 -46882 42526 -46865
rect 43082 -46865 43284 -46848
rect 43342 -46848 44302 -46810
rect 43342 -46865 43544 -46848
rect 43082 -46882 43098 -46865
rect 42510 -46898 43098 -46882
rect 43528 -46882 43544 -46865
rect 44100 -46865 44302 -46848
rect 44360 -46848 45320 -46810
rect 44360 -46865 44562 -46848
rect 44100 -46882 44116 -46865
rect 43528 -46898 44116 -46882
rect 44546 -46882 44562 -46865
rect 45118 -46865 45320 -46848
rect 45378 -46848 46338 -46810
rect 45378 -46865 45580 -46848
rect 45118 -46882 45134 -46865
rect 44546 -46898 45134 -46882
rect 45564 -46882 45580 -46865
rect 46136 -46865 46338 -46848
rect 46396 -46848 47356 -46810
rect 46396 -46865 46598 -46848
rect 46136 -46882 46152 -46865
rect 45564 -46898 46152 -46882
rect 46582 -46882 46598 -46865
rect 47154 -46865 47356 -46848
rect 47414 -46848 48374 -46810
rect 47414 -46865 47616 -46848
rect 47154 -46882 47170 -46865
rect 46582 -46898 47170 -46882
rect 47600 -46882 47616 -46865
rect 48172 -46865 48374 -46848
rect 48172 -46882 48188 -46865
rect 47600 -46898 48188 -46882
rect 24450 -46944 25410 -46906
rect 28258 -47370 28846 -47354
rect 28258 -47387 28274 -47370
rect 28072 -47404 28274 -47387
rect 28830 -47387 28846 -47370
rect 29276 -47370 29864 -47354
rect 29276 -47387 29292 -47370
rect 28830 -47404 29032 -47387
rect 28072 -47442 29032 -47404
rect 29090 -47404 29292 -47387
rect 29848 -47387 29864 -47370
rect 30294 -47370 30882 -47354
rect 30294 -47387 30310 -47370
rect 29848 -47404 30050 -47387
rect 29090 -47442 30050 -47404
rect 30108 -47404 30310 -47387
rect 30866 -47387 30882 -47370
rect 31312 -47370 31900 -47354
rect 31312 -47387 31328 -47370
rect 30866 -47404 31068 -47387
rect 30108 -47442 31068 -47404
rect 31126 -47404 31328 -47387
rect 31884 -47387 31900 -47370
rect 32330 -47370 32918 -47354
rect 32330 -47387 32346 -47370
rect 31884 -47404 32086 -47387
rect 31126 -47442 32086 -47404
rect 32144 -47404 32346 -47387
rect 32902 -47387 32918 -47370
rect 33348 -47370 33936 -47354
rect 33348 -47387 33364 -47370
rect 32902 -47404 33104 -47387
rect 32144 -47442 33104 -47404
rect 33162 -47404 33364 -47387
rect 33920 -47387 33936 -47370
rect 34366 -47370 34954 -47354
rect 34366 -47387 34382 -47370
rect 33920 -47404 34122 -47387
rect 33162 -47442 34122 -47404
rect 34180 -47404 34382 -47387
rect 34938 -47387 34954 -47370
rect 35384 -47370 35972 -47354
rect 35384 -47387 35400 -47370
rect 34938 -47404 35140 -47387
rect 34180 -47442 35140 -47404
rect 35198 -47404 35400 -47387
rect 35956 -47387 35972 -47370
rect 36402 -47370 36990 -47354
rect 36402 -47387 36418 -47370
rect 35956 -47404 36158 -47387
rect 35198 -47442 36158 -47404
rect 36216 -47404 36418 -47387
rect 36974 -47387 36990 -47370
rect 37420 -47370 38008 -47354
rect 37420 -47387 37436 -47370
rect 36974 -47404 37176 -47387
rect 36216 -47442 37176 -47404
rect 37234 -47404 37436 -47387
rect 37992 -47387 38008 -47370
rect 38438 -47370 39026 -47354
rect 38438 -47387 38454 -47370
rect 37992 -47404 38194 -47387
rect 37234 -47442 38194 -47404
rect 38252 -47404 38454 -47387
rect 39010 -47387 39026 -47370
rect 39456 -47370 40044 -47354
rect 39456 -47387 39472 -47370
rect 39010 -47404 39212 -47387
rect 38252 -47442 39212 -47404
rect 39270 -47404 39472 -47387
rect 40028 -47387 40044 -47370
rect 40474 -47370 41062 -47354
rect 40474 -47387 40490 -47370
rect 40028 -47404 40230 -47387
rect 39270 -47442 40230 -47404
rect 40288 -47404 40490 -47387
rect 41046 -47387 41062 -47370
rect 41492 -47370 42080 -47354
rect 41492 -47387 41508 -47370
rect 41046 -47404 41248 -47387
rect 40288 -47442 41248 -47404
rect 41306 -47404 41508 -47387
rect 42064 -47387 42080 -47370
rect 42510 -47370 43098 -47354
rect 42510 -47387 42526 -47370
rect 42064 -47404 42266 -47387
rect 41306 -47442 42266 -47404
rect 42324 -47404 42526 -47387
rect 43082 -47387 43098 -47370
rect 43528 -47370 44116 -47354
rect 43528 -47387 43544 -47370
rect 43082 -47404 43284 -47387
rect 42324 -47442 43284 -47404
rect 43342 -47404 43544 -47387
rect 44100 -47387 44116 -47370
rect 44546 -47370 45134 -47354
rect 44546 -47387 44562 -47370
rect 44100 -47404 44302 -47387
rect 43342 -47442 44302 -47404
rect 44360 -47404 44562 -47387
rect 45118 -47387 45134 -47370
rect 45564 -47370 46152 -47354
rect 45564 -47387 45580 -47370
rect 45118 -47404 45320 -47387
rect 44360 -47442 45320 -47404
rect 45378 -47404 45580 -47387
rect 46136 -47387 46152 -47370
rect 46582 -47370 47170 -47354
rect 46582 -47387 46598 -47370
rect 46136 -47404 46338 -47387
rect 45378 -47442 46338 -47404
rect 46396 -47404 46598 -47387
rect 47154 -47387 47170 -47370
rect 47600 -47370 48188 -47354
rect 47600 -47387 47616 -47370
rect 47154 -47404 47356 -47387
rect 46396 -47442 47356 -47404
rect 47414 -47404 47616 -47387
rect 48172 -47387 48188 -47370
rect 48172 -47404 48374 -47387
rect 47414 -47442 48374 -47404
rect 16306 -47582 17266 -47544
rect 16306 -47599 16508 -47582
rect 16492 -47616 16508 -47599
rect 17064 -47599 17266 -47582
rect 17324 -47582 18284 -47544
rect 17324 -47599 17526 -47582
rect 17064 -47616 17080 -47599
rect 16492 -47632 17080 -47616
rect 17510 -47616 17526 -47599
rect 18082 -47599 18284 -47582
rect 18342 -47582 19302 -47544
rect 18342 -47599 18544 -47582
rect 18082 -47616 18098 -47599
rect 17510 -47632 18098 -47616
rect 16492 -47690 17080 -47674
rect 16492 -47707 16508 -47690
rect 16306 -47724 16508 -47707
rect 17064 -47707 17080 -47690
rect 18528 -47616 18544 -47599
rect 19100 -47599 19302 -47582
rect 19360 -47582 20320 -47544
rect 19360 -47599 19562 -47582
rect 19100 -47616 19116 -47599
rect 18528 -47632 19116 -47616
rect 17510 -47690 18098 -47674
rect 17510 -47707 17526 -47690
rect 17064 -47724 17266 -47707
rect 16306 -47762 17266 -47724
rect 17324 -47724 17526 -47707
rect 18082 -47707 18098 -47690
rect 19546 -47616 19562 -47599
rect 20118 -47599 20320 -47582
rect 20378 -47582 21338 -47544
rect 20378 -47599 20580 -47582
rect 20118 -47616 20134 -47599
rect 19546 -47632 20134 -47616
rect 18528 -47690 19116 -47674
rect 18528 -47707 18544 -47690
rect 18082 -47724 18284 -47707
rect 17324 -47762 18284 -47724
rect 18342 -47724 18544 -47707
rect 19100 -47707 19116 -47690
rect 20564 -47616 20580 -47599
rect 21136 -47599 21338 -47582
rect 21396 -47582 22356 -47544
rect 21396 -47599 21598 -47582
rect 21136 -47616 21152 -47599
rect 20564 -47632 21152 -47616
rect 19546 -47690 20134 -47674
rect 19546 -47707 19562 -47690
rect 19100 -47724 19302 -47707
rect 18342 -47762 19302 -47724
rect 19360 -47724 19562 -47707
rect 20118 -47707 20134 -47690
rect 21582 -47616 21598 -47599
rect 22154 -47599 22356 -47582
rect 22414 -47582 23374 -47544
rect 22414 -47599 22616 -47582
rect 22154 -47616 22170 -47599
rect 21582 -47632 22170 -47616
rect 20564 -47690 21152 -47674
rect 20564 -47707 20580 -47690
rect 20118 -47724 20320 -47707
rect 19360 -47762 20320 -47724
rect 20378 -47724 20580 -47707
rect 21136 -47707 21152 -47690
rect 22600 -47616 22616 -47599
rect 23172 -47599 23374 -47582
rect 23432 -47582 24392 -47544
rect 23432 -47599 23634 -47582
rect 23172 -47616 23188 -47599
rect 22600 -47632 23188 -47616
rect 21582 -47690 22170 -47674
rect 21582 -47707 21598 -47690
rect 21136 -47724 21338 -47707
rect 20378 -47762 21338 -47724
rect 21396 -47724 21598 -47707
rect 22154 -47707 22170 -47690
rect 23618 -47616 23634 -47599
rect 24190 -47599 24392 -47582
rect 24450 -47582 25410 -47544
rect 24450 -47599 24652 -47582
rect 24190 -47616 24206 -47599
rect 23618 -47632 24206 -47616
rect 22600 -47690 23188 -47674
rect 22600 -47707 22616 -47690
rect 22154 -47724 22356 -47707
rect 21396 -47762 22356 -47724
rect 22414 -47724 22616 -47707
rect 23172 -47707 23188 -47690
rect 24636 -47616 24652 -47599
rect 25208 -47599 25410 -47582
rect 25208 -47616 25224 -47599
rect 24636 -47632 25224 -47616
rect 23618 -47690 24206 -47674
rect 23618 -47707 23634 -47690
rect 23172 -47724 23374 -47707
rect 22414 -47762 23374 -47724
rect 23432 -47724 23634 -47707
rect 24190 -47707 24206 -47690
rect 24636 -47690 25224 -47674
rect 24636 -47707 24652 -47690
rect 24190 -47724 24392 -47707
rect 23432 -47762 24392 -47724
rect 24450 -47724 24652 -47707
rect 25208 -47707 25224 -47690
rect 25208 -47724 25410 -47707
rect 24450 -47762 25410 -47724
rect 28072 -48080 29032 -48042
rect 28072 -48097 28274 -48080
rect 28258 -48114 28274 -48097
rect 28830 -48097 29032 -48080
rect 29090 -48080 30050 -48042
rect 29090 -48097 29292 -48080
rect 28830 -48114 28846 -48097
rect 28258 -48130 28846 -48114
rect 29276 -48114 29292 -48097
rect 29848 -48097 30050 -48080
rect 30108 -48080 31068 -48042
rect 30108 -48097 30310 -48080
rect 29848 -48114 29864 -48097
rect 29276 -48130 29864 -48114
rect 30294 -48114 30310 -48097
rect 30866 -48097 31068 -48080
rect 31126 -48080 32086 -48042
rect 31126 -48097 31328 -48080
rect 30866 -48114 30882 -48097
rect 30294 -48130 30882 -48114
rect 31312 -48114 31328 -48097
rect 31884 -48097 32086 -48080
rect 32144 -48080 33104 -48042
rect 32144 -48097 32346 -48080
rect 31884 -48114 31900 -48097
rect 31312 -48130 31900 -48114
rect 32330 -48114 32346 -48097
rect 32902 -48097 33104 -48080
rect 33162 -48080 34122 -48042
rect 33162 -48097 33364 -48080
rect 32902 -48114 32918 -48097
rect 32330 -48130 32918 -48114
rect 33348 -48114 33364 -48097
rect 33920 -48097 34122 -48080
rect 34180 -48080 35140 -48042
rect 34180 -48097 34382 -48080
rect 33920 -48114 33936 -48097
rect 33348 -48130 33936 -48114
rect 34366 -48114 34382 -48097
rect 34938 -48097 35140 -48080
rect 35198 -48080 36158 -48042
rect 35198 -48097 35400 -48080
rect 34938 -48114 34954 -48097
rect 34366 -48130 34954 -48114
rect 35384 -48114 35400 -48097
rect 35956 -48097 36158 -48080
rect 36216 -48080 37176 -48042
rect 36216 -48097 36418 -48080
rect 35956 -48114 35972 -48097
rect 35384 -48130 35972 -48114
rect 36402 -48114 36418 -48097
rect 36974 -48097 37176 -48080
rect 37234 -48080 38194 -48042
rect 37234 -48097 37436 -48080
rect 36974 -48114 36990 -48097
rect 36402 -48130 36990 -48114
rect 37420 -48114 37436 -48097
rect 37992 -48097 38194 -48080
rect 38252 -48080 39212 -48042
rect 38252 -48097 38454 -48080
rect 37992 -48114 38008 -48097
rect 37420 -48130 38008 -48114
rect 38438 -48114 38454 -48097
rect 39010 -48097 39212 -48080
rect 39270 -48080 40230 -48042
rect 39270 -48097 39472 -48080
rect 39010 -48114 39026 -48097
rect 38438 -48130 39026 -48114
rect 39456 -48114 39472 -48097
rect 40028 -48097 40230 -48080
rect 40288 -48080 41248 -48042
rect 40288 -48097 40490 -48080
rect 40028 -48114 40044 -48097
rect 39456 -48130 40044 -48114
rect 40474 -48114 40490 -48097
rect 41046 -48097 41248 -48080
rect 41306 -48080 42266 -48042
rect 41306 -48097 41508 -48080
rect 41046 -48114 41062 -48097
rect 40474 -48130 41062 -48114
rect 41492 -48114 41508 -48097
rect 42064 -48097 42266 -48080
rect 42324 -48080 43284 -48042
rect 42324 -48097 42526 -48080
rect 42064 -48114 42080 -48097
rect 41492 -48130 42080 -48114
rect 42510 -48114 42526 -48097
rect 43082 -48097 43284 -48080
rect 43342 -48080 44302 -48042
rect 43342 -48097 43544 -48080
rect 43082 -48114 43098 -48097
rect 42510 -48130 43098 -48114
rect 43528 -48114 43544 -48097
rect 44100 -48097 44302 -48080
rect 44360 -48080 45320 -48042
rect 44360 -48097 44562 -48080
rect 44100 -48114 44116 -48097
rect 43528 -48130 44116 -48114
rect 44546 -48114 44562 -48097
rect 45118 -48097 45320 -48080
rect 45378 -48080 46338 -48042
rect 45378 -48097 45580 -48080
rect 45118 -48114 45134 -48097
rect 44546 -48130 45134 -48114
rect 45564 -48114 45580 -48097
rect 46136 -48097 46338 -48080
rect 46396 -48080 47356 -48042
rect 46396 -48097 46598 -48080
rect 46136 -48114 46152 -48097
rect 45564 -48130 46152 -48114
rect 46582 -48114 46598 -48097
rect 47154 -48097 47356 -48080
rect 47414 -48080 48374 -48042
rect 47414 -48097 47616 -48080
rect 47154 -48114 47170 -48097
rect 46582 -48130 47170 -48114
rect 47600 -48114 47616 -48097
rect 48172 -48097 48374 -48080
rect 48172 -48114 48188 -48097
rect 47600 -48130 48188 -48114
rect 16306 -48400 17266 -48362
rect 16306 -48417 16508 -48400
rect 16492 -48434 16508 -48417
rect 17064 -48417 17266 -48400
rect 17324 -48400 18284 -48362
rect 17324 -48417 17526 -48400
rect 17064 -48434 17080 -48417
rect 16492 -48450 17080 -48434
rect 17510 -48434 17526 -48417
rect 18082 -48417 18284 -48400
rect 18342 -48400 19302 -48362
rect 18342 -48417 18544 -48400
rect 18082 -48434 18098 -48417
rect 17510 -48450 18098 -48434
rect 16492 -48508 17080 -48492
rect 16492 -48525 16508 -48508
rect 16306 -48542 16508 -48525
rect 17064 -48525 17080 -48508
rect 18528 -48434 18544 -48417
rect 19100 -48417 19302 -48400
rect 19360 -48400 20320 -48362
rect 19360 -48417 19562 -48400
rect 19100 -48434 19116 -48417
rect 18528 -48450 19116 -48434
rect 17510 -48508 18098 -48492
rect 17510 -48525 17526 -48508
rect 17064 -48542 17266 -48525
rect 16306 -48580 17266 -48542
rect 17324 -48542 17526 -48525
rect 18082 -48525 18098 -48508
rect 19546 -48434 19562 -48417
rect 20118 -48417 20320 -48400
rect 20378 -48400 21338 -48362
rect 20378 -48417 20580 -48400
rect 20118 -48434 20134 -48417
rect 19546 -48450 20134 -48434
rect 18528 -48508 19116 -48492
rect 18528 -48525 18544 -48508
rect 18082 -48542 18284 -48525
rect 17324 -48580 18284 -48542
rect 18342 -48542 18544 -48525
rect 19100 -48525 19116 -48508
rect 20564 -48434 20580 -48417
rect 21136 -48417 21338 -48400
rect 21396 -48400 22356 -48362
rect 21396 -48417 21598 -48400
rect 21136 -48434 21152 -48417
rect 20564 -48450 21152 -48434
rect 19546 -48508 20134 -48492
rect 19546 -48525 19562 -48508
rect 19100 -48542 19302 -48525
rect 18342 -48580 19302 -48542
rect 19360 -48542 19562 -48525
rect 20118 -48525 20134 -48508
rect 21582 -48434 21598 -48417
rect 22154 -48417 22356 -48400
rect 22414 -48400 23374 -48362
rect 22414 -48417 22616 -48400
rect 22154 -48434 22170 -48417
rect 21582 -48450 22170 -48434
rect 20564 -48508 21152 -48492
rect 20564 -48525 20580 -48508
rect 20118 -48542 20320 -48525
rect 19360 -48580 20320 -48542
rect 20378 -48542 20580 -48525
rect 21136 -48525 21152 -48508
rect 22600 -48434 22616 -48417
rect 23172 -48417 23374 -48400
rect 23432 -48400 24392 -48362
rect 23432 -48417 23634 -48400
rect 23172 -48434 23188 -48417
rect 22600 -48450 23188 -48434
rect 21582 -48508 22170 -48492
rect 21582 -48525 21598 -48508
rect 21136 -48542 21338 -48525
rect 20378 -48580 21338 -48542
rect 21396 -48542 21598 -48525
rect 22154 -48525 22170 -48508
rect 23618 -48434 23634 -48417
rect 24190 -48417 24392 -48400
rect 24450 -48400 25410 -48362
rect 24450 -48417 24652 -48400
rect 24190 -48434 24206 -48417
rect 23618 -48450 24206 -48434
rect 22600 -48508 23188 -48492
rect 22600 -48525 22616 -48508
rect 22154 -48542 22356 -48525
rect 21396 -48580 22356 -48542
rect 22414 -48542 22616 -48525
rect 23172 -48525 23188 -48508
rect 24636 -48434 24652 -48417
rect 25208 -48417 25410 -48400
rect 25208 -48434 25224 -48417
rect 24636 -48450 25224 -48434
rect 23618 -48508 24206 -48492
rect 23618 -48525 23634 -48508
rect 23172 -48542 23374 -48525
rect 22414 -48580 23374 -48542
rect 23432 -48542 23634 -48525
rect 24190 -48525 24206 -48508
rect 24636 -48508 25224 -48492
rect 24636 -48525 24652 -48508
rect 24190 -48542 24392 -48525
rect 23432 -48580 24392 -48542
rect 24450 -48542 24652 -48525
rect 25208 -48525 25224 -48508
rect 25208 -48542 25410 -48525
rect 24450 -48580 25410 -48542
rect 28256 -48604 28844 -48588
rect 28256 -48621 28272 -48604
rect 28070 -48638 28272 -48621
rect 28828 -48621 28844 -48604
rect 29274 -48604 29862 -48588
rect 29274 -48621 29290 -48604
rect 28828 -48638 29030 -48621
rect 28070 -48676 29030 -48638
rect 29088 -48638 29290 -48621
rect 29846 -48621 29862 -48604
rect 30292 -48604 30880 -48588
rect 30292 -48621 30308 -48604
rect 29846 -48638 30048 -48621
rect 29088 -48676 30048 -48638
rect 30106 -48638 30308 -48621
rect 30864 -48621 30880 -48604
rect 31310 -48604 31898 -48588
rect 31310 -48621 31326 -48604
rect 30864 -48638 31066 -48621
rect 30106 -48676 31066 -48638
rect 31124 -48638 31326 -48621
rect 31882 -48621 31898 -48604
rect 32328 -48604 32916 -48588
rect 32328 -48621 32344 -48604
rect 31882 -48638 32084 -48621
rect 31124 -48676 32084 -48638
rect 32142 -48638 32344 -48621
rect 32900 -48621 32916 -48604
rect 33346 -48604 33934 -48588
rect 33346 -48621 33362 -48604
rect 32900 -48638 33102 -48621
rect 32142 -48676 33102 -48638
rect 33160 -48638 33362 -48621
rect 33918 -48621 33934 -48604
rect 34364 -48604 34952 -48588
rect 34364 -48621 34380 -48604
rect 33918 -48638 34120 -48621
rect 33160 -48676 34120 -48638
rect 34178 -48638 34380 -48621
rect 34936 -48621 34952 -48604
rect 35382 -48604 35970 -48588
rect 35382 -48621 35398 -48604
rect 34936 -48638 35138 -48621
rect 34178 -48676 35138 -48638
rect 35196 -48638 35398 -48621
rect 35954 -48621 35970 -48604
rect 36400 -48604 36988 -48588
rect 36400 -48621 36416 -48604
rect 35954 -48638 36156 -48621
rect 35196 -48676 36156 -48638
rect 36214 -48638 36416 -48621
rect 36972 -48621 36988 -48604
rect 37418 -48604 38006 -48588
rect 37418 -48621 37434 -48604
rect 36972 -48638 37174 -48621
rect 36214 -48676 37174 -48638
rect 37232 -48638 37434 -48621
rect 37990 -48621 38006 -48604
rect 38436 -48604 39024 -48588
rect 38436 -48621 38452 -48604
rect 37990 -48638 38192 -48621
rect 37232 -48676 38192 -48638
rect 38250 -48638 38452 -48621
rect 39008 -48621 39024 -48604
rect 39454 -48604 40042 -48588
rect 39454 -48621 39470 -48604
rect 39008 -48638 39210 -48621
rect 38250 -48676 39210 -48638
rect 39268 -48638 39470 -48621
rect 40026 -48621 40042 -48604
rect 40472 -48604 41060 -48588
rect 40472 -48621 40488 -48604
rect 40026 -48638 40228 -48621
rect 39268 -48676 40228 -48638
rect 40286 -48638 40488 -48621
rect 41044 -48621 41060 -48604
rect 41490 -48604 42078 -48588
rect 41490 -48621 41506 -48604
rect 41044 -48638 41246 -48621
rect 40286 -48676 41246 -48638
rect 41304 -48638 41506 -48621
rect 42062 -48621 42078 -48604
rect 42508 -48604 43096 -48588
rect 42508 -48621 42524 -48604
rect 42062 -48638 42264 -48621
rect 41304 -48676 42264 -48638
rect 42322 -48638 42524 -48621
rect 43080 -48621 43096 -48604
rect 43526 -48604 44114 -48588
rect 43526 -48621 43542 -48604
rect 43080 -48638 43282 -48621
rect 42322 -48676 43282 -48638
rect 43340 -48638 43542 -48621
rect 44098 -48621 44114 -48604
rect 44544 -48604 45132 -48588
rect 44544 -48621 44560 -48604
rect 44098 -48638 44300 -48621
rect 43340 -48676 44300 -48638
rect 44358 -48638 44560 -48621
rect 45116 -48621 45132 -48604
rect 45562 -48604 46150 -48588
rect 45562 -48621 45578 -48604
rect 45116 -48638 45318 -48621
rect 44358 -48676 45318 -48638
rect 45376 -48638 45578 -48621
rect 46134 -48621 46150 -48604
rect 46580 -48604 47168 -48588
rect 46580 -48621 46596 -48604
rect 46134 -48638 46336 -48621
rect 45376 -48676 46336 -48638
rect 46394 -48638 46596 -48621
rect 47152 -48621 47168 -48604
rect 47598 -48604 48186 -48588
rect 47598 -48621 47614 -48604
rect 47152 -48638 47354 -48621
rect 46394 -48676 47354 -48638
rect 47412 -48638 47614 -48621
rect 48170 -48621 48186 -48604
rect 48170 -48638 48372 -48621
rect 47412 -48676 48372 -48638
rect 16306 -49218 17266 -49180
rect 16306 -49235 16508 -49218
rect 16492 -49252 16508 -49235
rect 17064 -49235 17266 -49218
rect 17324 -49218 18284 -49180
rect 17324 -49235 17526 -49218
rect 17064 -49252 17080 -49235
rect 16492 -49268 17080 -49252
rect 17510 -49252 17526 -49235
rect 18082 -49235 18284 -49218
rect 18342 -49218 19302 -49180
rect 18342 -49235 18544 -49218
rect 18082 -49252 18098 -49235
rect 17510 -49268 18098 -49252
rect 16492 -49326 17080 -49310
rect 16492 -49343 16508 -49326
rect 16306 -49360 16508 -49343
rect 17064 -49343 17080 -49326
rect 18528 -49252 18544 -49235
rect 19100 -49235 19302 -49218
rect 19360 -49218 20320 -49180
rect 19360 -49235 19562 -49218
rect 19100 -49252 19116 -49235
rect 18528 -49268 19116 -49252
rect 17510 -49326 18098 -49310
rect 17510 -49343 17526 -49326
rect 17064 -49360 17266 -49343
rect 16306 -49398 17266 -49360
rect 17324 -49360 17526 -49343
rect 18082 -49343 18098 -49326
rect 19546 -49252 19562 -49235
rect 20118 -49235 20320 -49218
rect 20378 -49218 21338 -49180
rect 20378 -49235 20580 -49218
rect 20118 -49252 20134 -49235
rect 19546 -49268 20134 -49252
rect 18528 -49326 19116 -49310
rect 18528 -49343 18544 -49326
rect 18082 -49360 18284 -49343
rect 17324 -49398 18284 -49360
rect 18342 -49360 18544 -49343
rect 19100 -49343 19116 -49326
rect 20564 -49252 20580 -49235
rect 21136 -49235 21338 -49218
rect 21396 -49218 22356 -49180
rect 21396 -49235 21598 -49218
rect 21136 -49252 21152 -49235
rect 20564 -49268 21152 -49252
rect 19546 -49326 20134 -49310
rect 19546 -49343 19562 -49326
rect 19100 -49360 19302 -49343
rect 18342 -49398 19302 -49360
rect 19360 -49360 19562 -49343
rect 20118 -49343 20134 -49326
rect 21582 -49252 21598 -49235
rect 22154 -49235 22356 -49218
rect 22414 -49218 23374 -49180
rect 22414 -49235 22616 -49218
rect 22154 -49252 22170 -49235
rect 21582 -49268 22170 -49252
rect 20564 -49326 21152 -49310
rect 20564 -49343 20580 -49326
rect 20118 -49360 20320 -49343
rect 19360 -49398 20320 -49360
rect 20378 -49360 20580 -49343
rect 21136 -49343 21152 -49326
rect 22600 -49252 22616 -49235
rect 23172 -49235 23374 -49218
rect 23432 -49218 24392 -49180
rect 23432 -49235 23634 -49218
rect 23172 -49252 23188 -49235
rect 22600 -49268 23188 -49252
rect 21582 -49326 22170 -49310
rect 21582 -49343 21598 -49326
rect 21136 -49360 21338 -49343
rect 20378 -49398 21338 -49360
rect 21396 -49360 21598 -49343
rect 22154 -49343 22170 -49326
rect 23618 -49252 23634 -49235
rect 24190 -49235 24392 -49218
rect 24450 -49218 25410 -49180
rect 24450 -49235 24652 -49218
rect 24190 -49252 24206 -49235
rect 23618 -49268 24206 -49252
rect 22600 -49326 23188 -49310
rect 22600 -49343 22616 -49326
rect 22154 -49360 22356 -49343
rect 21396 -49398 22356 -49360
rect 22414 -49360 22616 -49343
rect 23172 -49343 23188 -49326
rect 24636 -49252 24652 -49235
rect 25208 -49235 25410 -49218
rect 25208 -49252 25224 -49235
rect 24636 -49268 25224 -49252
rect 23618 -49326 24206 -49310
rect 23618 -49343 23634 -49326
rect 23172 -49360 23374 -49343
rect 22414 -49398 23374 -49360
rect 23432 -49360 23634 -49343
rect 24190 -49343 24206 -49326
rect 24636 -49326 25224 -49310
rect 24636 -49343 24652 -49326
rect 24190 -49360 24392 -49343
rect 23432 -49398 24392 -49360
rect 24450 -49360 24652 -49343
rect 25208 -49343 25224 -49326
rect 28070 -49314 29030 -49276
rect 28070 -49331 28272 -49314
rect 25208 -49360 25410 -49343
rect 24450 -49398 25410 -49360
rect 28256 -49348 28272 -49331
rect 28828 -49331 29030 -49314
rect 29088 -49314 30048 -49276
rect 29088 -49331 29290 -49314
rect 28828 -49348 28844 -49331
rect 28256 -49364 28844 -49348
rect 29274 -49348 29290 -49331
rect 29846 -49331 30048 -49314
rect 30106 -49314 31066 -49276
rect 30106 -49331 30308 -49314
rect 29846 -49348 29862 -49331
rect 29274 -49364 29862 -49348
rect 30292 -49348 30308 -49331
rect 30864 -49331 31066 -49314
rect 31124 -49314 32084 -49276
rect 31124 -49331 31326 -49314
rect 30864 -49348 30880 -49331
rect 30292 -49364 30880 -49348
rect 31310 -49348 31326 -49331
rect 31882 -49331 32084 -49314
rect 32142 -49314 33102 -49276
rect 32142 -49331 32344 -49314
rect 31882 -49348 31898 -49331
rect 31310 -49364 31898 -49348
rect 32328 -49348 32344 -49331
rect 32900 -49331 33102 -49314
rect 33160 -49314 34120 -49276
rect 33160 -49331 33362 -49314
rect 32900 -49348 32916 -49331
rect 32328 -49364 32916 -49348
rect 33346 -49348 33362 -49331
rect 33918 -49331 34120 -49314
rect 34178 -49314 35138 -49276
rect 34178 -49331 34380 -49314
rect 33918 -49348 33934 -49331
rect 33346 -49364 33934 -49348
rect 34364 -49348 34380 -49331
rect 34936 -49331 35138 -49314
rect 35196 -49314 36156 -49276
rect 35196 -49331 35398 -49314
rect 34936 -49348 34952 -49331
rect 34364 -49364 34952 -49348
rect 35382 -49348 35398 -49331
rect 35954 -49331 36156 -49314
rect 36214 -49314 37174 -49276
rect 36214 -49331 36416 -49314
rect 35954 -49348 35970 -49331
rect 35382 -49364 35970 -49348
rect 36400 -49348 36416 -49331
rect 36972 -49331 37174 -49314
rect 37232 -49314 38192 -49276
rect 37232 -49331 37434 -49314
rect 36972 -49348 36988 -49331
rect 36400 -49364 36988 -49348
rect 37418 -49348 37434 -49331
rect 37990 -49331 38192 -49314
rect 38250 -49314 39210 -49276
rect 38250 -49331 38452 -49314
rect 37990 -49348 38006 -49331
rect 37418 -49364 38006 -49348
rect 38436 -49348 38452 -49331
rect 39008 -49331 39210 -49314
rect 39268 -49314 40228 -49276
rect 39268 -49331 39470 -49314
rect 39008 -49348 39024 -49331
rect 38436 -49364 39024 -49348
rect 39454 -49348 39470 -49331
rect 40026 -49331 40228 -49314
rect 40286 -49314 41246 -49276
rect 40286 -49331 40488 -49314
rect 40026 -49348 40042 -49331
rect 39454 -49364 40042 -49348
rect 40472 -49348 40488 -49331
rect 41044 -49331 41246 -49314
rect 41304 -49314 42264 -49276
rect 41304 -49331 41506 -49314
rect 41044 -49348 41060 -49331
rect 40472 -49364 41060 -49348
rect 41490 -49348 41506 -49331
rect 42062 -49331 42264 -49314
rect 42322 -49314 43282 -49276
rect 42322 -49331 42524 -49314
rect 42062 -49348 42078 -49331
rect 41490 -49364 42078 -49348
rect 42508 -49348 42524 -49331
rect 43080 -49331 43282 -49314
rect 43340 -49314 44300 -49276
rect 43340 -49331 43542 -49314
rect 43080 -49348 43096 -49331
rect 42508 -49364 43096 -49348
rect 43526 -49348 43542 -49331
rect 44098 -49331 44300 -49314
rect 44358 -49314 45318 -49276
rect 44358 -49331 44560 -49314
rect 44098 -49348 44114 -49331
rect 43526 -49364 44114 -49348
rect 44544 -49348 44560 -49331
rect 45116 -49331 45318 -49314
rect 45376 -49314 46336 -49276
rect 45376 -49331 45578 -49314
rect 45116 -49348 45132 -49331
rect 44544 -49364 45132 -49348
rect 45562 -49348 45578 -49331
rect 46134 -49331 46336 -49314
rect 46394 -49314 47354 -49276
rect 46394 -49331 46596 -49314
rect 46134 -49348 46150 -49331
rect 45562 -49364 46150 -49348
rect 46580 -49348 46596 -49331
rect 47152 -49331 47354 -49314
rect 47412 -49314 48372 -49276
rect 47412 -49331 47614 -49314
rect 47152 -49348 47168 -49331
rect 46580 -49364 47168 -49348
rect 47598 -49348 47614 -49331
rect 48170 -49331 48372 -49314
rect 48170 -49348 48186 -49331
rect 47598 -49364 48186 -49348
rect 28256 -49838 28844 -49822
rect 28256 -49855 28272 -49838
rect 28070 -49872 28272 -49855
rect 28828 -49855 28844 -49838
rect 29274 -49838 29862 -49822
rect 29274 -49855 29290 -49838
rect 28828 -49872 29030 -49855
rect 28070 -49910 29030 -49872
rect 29088 -49872 29290 -49855
rect 29846 -49855 29862 -49838
rect 30292 -49838 30880 -49822
rect 30292 -49855 30308 -49838
rect 29846 -49872 30048 -49855
rect 29088 -49910 30048 -49872
rect 30106 -49872 30308 -49855
rect 30864 -49855 30880 -49838
rect 31310 -49838 31898 -49822
rect 31310 -49855 31326 -49838
rect 30864 -49872 31066 -49855
rect 30106 -49910 31066 -49872
rect 31124 -49872 31326 -49855
rect 31882 -49855 31898 -49838
rect 32328 -49838 32916 -49822
rect 32328 -49855 32344 -49838
rect 31882 -49872 32084 -49855
rect 31124 -49910 32084 -49872
rect 32142 -49872 32344 -49855
rect 32900 -49855 32916 -49838
rect 33346 -49838 33934 -49822
rect 33346 -49855 33362 -49838
rect 32900 -49872 33102 -49855
rect 32142 -49910 33102 -49872
rect 33160 -49872 33362 -49855
rect 33918 -49855 33934 -49838
rect 34364 -49838 34952 -49822
rect 34364 -49855 34380 -49838
rect 33918 -49872 34120 -49855
rect 33160 -49910 34120 -49872
rect 34178 -49872 34380 -49855
rect 34936 -49855 34952 -49838
rect 35382 -49838 35970 -49822
rect 35382 -49855 35398 -49838
rect 34936 -49872 35138 -49855
rect 34178 -49910 35138 -49872
rect 35196 -49872 35398 -49855
rect 35954 -49855 35970 -49838
rect 36400 -49838 36988 -49822
rect 36400 -49855 36416 -49838
rect 35954 -49872 36156 -49855
rect 35196 -49910 36156 -49872
rect 36214 -49872 36416 -49855
rect 36972 -49855 36988 -49838
rect 37418 -49838 38006 -49822
rect 37418 -49855 37434 -49838
rect 36972 -49872 37174 -49855
rect 36214 -49910 37174 -49872
rect 37232 -49872 37434 -49855
rect 37990 -49855 38006 -49838
rect 38436 -49838 39024 -49822
rect 38436 -49855 38452 -49838
rect 37990 -49872 38192 -49855
rect 37232 -49910 38192 -49872
rect 38250 -49872 38452 -49855
rect 39008 -49855 39024 -49838
rect 39454 -49838 40042 -49822
rect 39454 -49855 39470 -49838
rect 39008 -49872 39210 -49855
rect 38250 -49910 39210 -49872
rect 39268 -49872 39470 -49855
rect 40026 -49855 40042 -49838
rect 40472 -49838 41060 -49822
rect 40472 -49855 40488 -49838
rect 40026 -49872 40228 -49855
rect 39268 -49910 40228 -49872
rect 40286 -49872 40488 -49855
rect 41044 -49855 41060 -49838
rect 41490 -49838 42078 -49822
rect 41490 -49855 41506 -49838
rect 41044 -49872 41246 -49855
rect 40286 -49910 41246 -49872
rect 41304 -49872 41506 -49855
rect 42062 -49855 42078 -49838
rect 42508 -49838 43096 -49822
rect 42508 -49855 42524 -49838
rect 42062 -49872 42264 -49855
rect 41304 -49910 42264 -49872
rect 42322 -49872 42524 -49855
rect 43080 -49855 43096 -49838
rect 43526 -49838 44114 -49822
rect 43526 -49855 43542 -49838
rect 43080 -49872 43282 -49855
rect 42322 -49910 43282 -49872
rect 43340 -49872 43542 -49855
rect 44098 -49855 44114 -49838
rect 44544 -49838 45132 -49822
rect 44544 -49855 44560 -49838
rect 44098 -49872 44300 -49855
rect 43340 -49910 44300 -49872
rect 44358 -49872 44560 -49855
rect 45116 -49855 45132 -49838
rect 45562 -49838 46150 -49822
rect 45562 -49855 45578 -49838
rect 45116 -49872 45318 -49855
rect 44358 -49910 45318 -49872
rect 45376 -49872 45578 -49855
rect 46134 -49855 46150 -49838
rect 46580 -49838 47168 -49822
rect 46580 -49855 46596 -49838
rect 46134 -49872 46336 -49855
rect 45376 -49910 46336 -49872
rect 46394 -49872 46596 -49855
rect 47152 -49855 47168 -49838
rect 47598 -49838 48186 -49822
rect 47598 -49855 47614 -49838
rect 47152 -49872 47354 -49855
rect 46394 -49910 47354 -49872
rect 47412 -49872 47614 -49855
rect 48170 -49855 48186 -49838
rect 48170 -49872 48372 -49855
rect 47412 -49910 48372 -49872
rect 16306 -50036 17266 -49998
rect 16306 -50053 16508 -50036
rect 16492 -50070 16508 -50053
rect 17064 -50053 17266 -50036
rect 17324 -50036 18284 -49998
rect 17324 -50053 17526 -50036
rect 17064 -50070 17080 -50053
rect 16492 -50086 17080 -50070
rect 17510 -50070 17526 -50053
rect 18082 -50053 18284 -50036
rect 18342 -50036 19302 -49998
rect 18342 -50053 18544 -50036
rect 18082 -50070 18098 -50053
rect 17510 -50086 18098 -50070
rect 16492 -50144 17080 -50128
rect 16492 -50161 16508 -50144
rect 16306 -50178 16508 -50161
rect 17064 -50161 17080 -50144
rect 18528 -50070 18544 -50053
rect 19100 -50053 19302 -50036
rect 19360 -50036 20320 -49998
rect 19360 -50053 19562 -50036
rect 19100 -50070 19116 -50053
rect 18528 -50086 19116 -50070
rect 17510 -50144 18098 -50128
rect 17510 -50161 17526 -50144
rect 17064 -50178 17266 -50161
rect 16306 -50216 17266 -50178
rect 17324 -50178 17526 -50161
rect 18082 -50161 18098 -50144
rect 19546 -50070 19562 -50053
rect 20118 -50053 20320 -50036
rect 20378 -50036 21338 -49998
rect 20378 -50053 20580 -50036
rect 20118 -50070 20134 -50053
rect 19546 -50086 20134 -50070
rect 18528 -50144 19116 -50128
rect 18528 -50161 18544 -50144
rect 18082 -50178 18284 -50161
rect 17324 -50216 18284 -50178
rect 18342 -50178 18544 -50161
rect 19100 -50161 19116 -50144
rect 20564 -50070 20580 -50053
rect 21136 -50053 21338 -50036
rect 21396 -50036 22356 -49998
rect 21396 -50053 21598 -50036
rect 21136 -50070 21152 -50053
rect 20564 -50086 21152 -50070
rect 19546 -50144 20134 -50128
rect 19546 -50161 19562 -50144
rect 19100 -50178 19302 -50161
rect 18342 -50216 19302 -50178
rect 19360 -50178 19562 -50161
rect 20118 -50161 20134 -50144
rect 21582 -50070 21598 -50053
rect 22154 -50053 22356 -50036
rect 22414 -50036 23374 -49998
rect 22414 -50053 22616 -50036
rect 22154 -50070 22170 -50053
rect 21582 -50086 22170 -50070
rect 20564 -50144 21152 -50128
rect 20564 -50161 20580 -50144
rect 20118 -50178 20320 -50161
rect 19360 -50216 20320 -50178
rect 20378 -50178 20580 -50161
rect 21136 -50161 21152 -50144
rect 22600 -50070 22616 -50053
rect 23172 -50053 23374 -50036
rect 23432 -50036 24392 -49998
rect 23432 -50053 23634 -50036
rect 23172 -50070 23188 -50053
rect 22600 -50086 23188 -50070
rect 21582 -50144 22170 -50128
rect 21582 -50161 21598 -50144
rect 21136 -50178 21338 -50161
rect 20378 -50216 21338 -50178
rect 21396 -50178 21598 -50161
rect 22154 -50161 22170 -50144
rect 23618 -50070 23634 -50053
rect 24190 -50053 24392 -50036
rect 24450 -50036 25410 -49998
rect 24450 -50053 24652 -50036
rect 24190 -50070 24206 -50053
rect 23618 -50086 24206 -50070
rect 22600 -50144 23188 -50128
rect 22600 -50161 22616 -50144
rect 22154 -50178 22356 -50161
rect 21396 -50216 22356 -50178
rect 22414 -50178 22616 -50161
rect 23172 -50161 23188 -50144
rect 24636 -50070 24652 -50053
rect 25208 -50053 25410 -50036
rect 25208 -50070 25224 -50053
rect 24636 -50086 25224 -50070
rect 23618 -50144 24206 -50128
rect 23618 -50161 23634 -50144
rect 23172 -50178 23374 -50161
rect 22414 -50216 23374 -50178
rect 23432 -50178 23634 -50161
rect 24190 -50161 24206 -50144
rect 24636 -50144 25224 -50128
rect 24636 -50161 24652 -50144
rect 24190 -50178 24392 -50161
rect 23432 -50216 24392 -50178
rect 24450 -50178 24652 -50161
rect 25208 -50161 25224 -50144
rect 25208 -50178 25410 -50161
rect 24450 -50216 25410 -50178
rect 28070 -50548 29030 -50510
rect 28070 -50565 28272 -50548
rect 28256 -50582 28272 -50565
rect 28828 -50565 29030 -50548
rect 29088 -50548 30048 -50510
rect 29088 -50565 29290 -50548
rect 28828 -50582 28844 -50565
rect 28256 -50598 28844 -50582
rect 29274 -50582 29290 -50565
rect 29846 -50565 30048 -50548
rect 30106 -50548 31066 -50510
rect 30106 -50565 30308 -50548
rect 29846 -50582 29862 -50565
rect 29274 -50598 29862 -50582
rect 30292 -50582 30308 -50565
rect 30864 -50565 31066 -50548
rect 31124 -50548 32084 -50510
rect 31124 -50565 31326 -50548
rect 30864 -50582 30880 -50565
rect 30292 -50598 30880 -50582
rect 31310 -50582 31326 -50565
rect 31882 -50565 32084 -50548
rect 32142 -50548 33102 -50510
rect 32142 -50565 32344 -50548
rect 31882 -50582 31898 -50565
rect 31310 -50598 31898 -50582
rect 32328 -50582 32344 -50565
rect 32900 -50565 33102 -50548
rect 33160 -50548 34120 -50510
rect 33160 -50565 33362 -50548
rect 32900 -50582 32916 -50565
rect 32328 -50598 32916 -50582
rect 33346 -50582 33362 -50565
rect 33918 -50565 34120 -50548
rect 34178 -50548 35138 -50510
rect 34178 -50565 34380 -50548
rect 33918 -50582 33934 -50565
rect 33346 -50598 33934 -50582
rect 34364 -50582 34380 -50565
rect 34936 -50565 35138 -50548
rect 35196 -50548 36156 -50510
rect 35196 -50565 35398 -50548
rect 34936 -50582 34952 -50565
rect 34364 -50598 34952 -50582
rect 35382 -50582 35398 -50565
rect 35954 -50565 36156 -50548
rect 36214 -50548 37174 -50510
rect 36214 -50565 36416 -50548
rect 35954 -50582 35970 -50565
rect 35382 -50598 35970 -50582
rect 36400 -50582 36416 -50565
rect 36972 -50565 37174 -50548
rect 37232 -50548 38192 -50510
rect 37232 -50565 37434 -50548
rect 36972 -50582 36988 -50565
rect 36400 -50598 36988 -50582
rect 37418 -50582 37434 -50565
rect 37990 -50565 38192 -50548
rect 38250 -50548 39210 -50510
rect 38250 -50565 38452 -50548
rect 37990 -50582 38006 -50565
rect 37418 -50598 38006 -50582
rect 38436 -50582 38452 -50565
rect 39008 -50565 39210 -50548
rect 39268 -50548 40228 -50510
rect 39268 -50565 39470 -50548
rect 39008 -50582 39024 -50565
rect 38436 -50598 39024 -50582
rect 39454 -50582 39470 -50565
rect 40026 -50565 40228 -50548
rect 40286 -50548 41246 -50510
rect 40286 -50565 40488 -50548
rect 40026 -50582 40042 -50565
rect 39454 -50598 40042 -50582
rect 40472 -50582 40488 -50565
rect 41044 -50565 41246 -50548
rect 41304 -50548 42264 -50510
rect 41304 -50565 41506 -50548
rect 41044 -50582 41060 -50565
rect 40472 -50598 41060 -50582
rect 41490 -50582 41506 -50565
rect 42062 -50565 42264 -50548
rect 42322 -50548 43282 -50510
rect 42322 -50565 42524 -50548
rect 42062 -50582 42078 -50565
rect 41490 -50598 42078 -50582
rect 42508 -50582 42524 -50565
rect 43080 -50565 43282 -50548
rect 43340 -50548 44300 -50510
rect 43340 -50565 43542 -50548
rect 43080 -50582 43096 -50565
rect 42508 -50598 43096 -50582
rect 43526 -50582 43542 -50565
rect 44098 -50565 44300 -50548
rect 44358 -50548 45318 -50510
rect 44358 -50565 44560 -50548
rect 44098 -50582 44114 -50565
rect 43526 -50598 44114 -50582
rect 44544 -50582 44560 -50565
rect 45116 -50565 45318 -50548
rect 45376 -50548 46336 -50510
rect 45376 -50565 45578 -50548
rect 45116 -50582 45132 -50565
rect 44544 -50598 45132 -50582
rect 45562 -50582 45578 -50565
rect 46134 -50565 46336 -50548
rect 46394 -50548 47354 -50510
rect 46394 -50565 46596 -50548
rect 46134 -50582 46150 -50565
rect 45562 -50598 46150 -50582
rect 46580 -50582 46596 -50565
rect 47152 -50565 47354 -50548
rect 47412 -50548 48372 -50510
rect 47412 -50565 47614 -50548
rect 47152 -50582 47168 -50565
rect 46580 -50598 47168 -50582
rect 47598 -50582 47614 -50565
rect 48170 -50565 48372 -50548
rect 48170 -50582 48186 -50565
rect 47598 -50598 48186 -50582
rect 16306 -50854 17266 -50816
rect 16306 -50871 16508 -50854
rect 16492 -50888 16508 -50871
rect 17064 -50871 17266 -50854
rect 17324 -50854 18284 -50816
rect 17324 -50871 17526 -50854
rect 17064 -50888 17080 -50871
rect 16492 -50904 17080 -50888
rect 17510 -50888 17526 -50871
rect 18082 -50871 18284 -50854
rect 18342 -50854 19302 -50816
rect 18342 -50871 18544 -50854
rect 18082 -50888 18098 -50871
rect 17510 -50904 18098 -50888
rect 18528 -50888 18544 -50871
rect 19100 -50871 19302 -50854
rect 19360 -50854 20320 -50816
rect 19360 -50871 19562 -50854
rect 19100 -50888 19116 -50871
rect 18528 -50904 19116 -50888
rect 19546 -50888 19562 -50871
rect 20118 -50871 20320 -50854
rect 20378 -50854 21338 -50816
rect 20378 -50871 20580 -50854
rect 20118 -50888 20134 -50871
rect 19546 -50904 20134 -50888
rect 20564 -50888 20580 -50871
rect 21136 -50871 21338 -50854
rect 21396 -50854 22356 -50816
rect 21396 -50871 21598 -50854
rect 21136 -50888 21152 -50871
rect 20564 -50904 21152 -50888
rect 21582 -50888 21598 -50871
rect 22154 -50871 22356 -50854
rect 22414 -50854 23374 -50816
rect 22414 -50871 22616 -50854
rect 22154 -50888 22170 -50871
rect 21582 -50904 22170 -50888
rect 22600 -50888 22616 -50871
rect 23172 -50871 23374 -50854
rect 23432 -50854 24392 -50816
rect 23432 -50871 23634 -50854
rect 23172 -50888 23188 -50871
rect 22600 -50904 23188 -50888
rect 23618 -50888 23634 -50871
rect 24190 -50871 24392 -50854
rect 24450 -50854 25410 -50816
rect 24450 -50871 24652 -50854
rect 24190 -50888 24206 -50871
rect 23618 -50904 24206 -50888
rect 24636 -50888 24652 -50871
rect 25208 -50871 25410 -50854
rect 25208 -50888 25224 -50871
rect 24636 -50904 25224 -50888
rect 28256 -51070 28844 -51054
rect 28256 -51087 28272 -51070
rect 28070 -51104 28272 -51087
rect 28828 -51087 28844 -51070
rect 29274 -51070 29862 -51054
rect 29274 -51087 29290 -51070
rect 28828 -51104 29030 -51087
rect 28070 -51142 29030 -51104
rect 29088 -51104 29290 -51087
rect 29846 -51087 29862 -51070
rect 30292 -51070 30880 -51054
rect 30292 -51087 30308 -51070
rect 29846 -51104 30048 -51087
rect 29088 -51142 30048 -51104
rect 30106 -51104 30308 -51087
rect 30864 -51087 30880 -51070
rect 31310 -51070 31898 -51054
rect 31310 -51087 31326 -51070
rect 30864 -51104 31066 -51087
rect 30106 -51142 31066 -51104
rect 31124 -51104 31326 -51087
rect 31882 -51087 31898 -51070
rect 32328 -51070 32916 -51054
rect 32328 -51087 32344 -51070
rect 31882 -51104 32084 -51087
rect 31124 -51142 32084 -51104
rect 32142 -51104 32344 -51087
rect 32900 -51087 32916 -51070
rect 33346 -51070 33934 -51054
rect 33346 -51087 33362 -51070
rect 32900 -51104 33102 -51087
rect 32142 -51142 33102 -51104
rect 33160 -51104 33362 -51087
rect 33918 -51087 33934 -51070
rect 34364 -51070 34952 -51054
rect 34364 -51087 34380 -51070
rect 33918 -51104 34120 -51087
rect 33160 -51142 34120 -51104
rect 34178 -51104 34380 -51087
rect 34936 -51087 34952 -51070
rect 35382 -51070 35970 -51054
rect 35382 -51087 35398 -51070
rect 34936 -51104 35138 -51087
rect 34178 -51142 35138 -51104
rect 35196 -51104 35398 -51087
rect 35954 -51087 35970 -51070
rect 36400 -51070 36988 -51054
rect 36400 -51087 36416 -51070
rect 35954 -51104 36156 -51087
rect 35196 -51142 36156 -51104
rect 36214 -51104 36416 -51087
rect 36972 -51087 36988 -51070
rect 37418 -51070 38006 -51054
rect 37418 -51087 37434 -51070
rect 36972 -51104 37174 -51087
rect 36214 -51142 37174 -51104
rect 37232 -51104 37434 -51087
rect 37990 -51087 38006 -51070
rect 38436 -51070 39024 -51054
rect 38436 -51087 38452 -51070
rect 37990 -51104 38192 -51087
rect 37232 -51142 38192 -51104
rect 38250 -51104 38452 -51087
rect 39008 -51087 39024 -51070
rect 39454 -51070 40042 -51054
rect 39454 -51087 39470 -51070
rect 39008 -51104 39210 -51087
rect 38250 -51142 39210 -51104
rect 39268 -51104 39470 -51087
rect 40026 -51087 40042 -51070
rect 40472 -51070 41060 -51054
rect 40472 -51087 40488 -51070
rect 40026 -51104 40228 -51087
rect 39268 -51142 40228 -51104
rect 40286 -51104 40488 -51087
rect 41044 -51087 41060 -51070
rect 41490 -51070 42078 -51054
rect 41490 -51087 41506 -51070
rect 41044 -51104 41246 -51087
rect 40286 -51142 41246 -51104
rect 41304 -51104 41506 -51087
rect 42062 -51087 42078 -51070
rect 42508 -51070 43096 -51054
rect 42508 -51087 42524 -51070
rect 42062 -51104 42264 -51087
rect 41304 -51142 42264 -51104
rect 42322 -51104 42524 -51087
rect 43080 -51087 43096 -51070
rect 43526 -51070 44114 -51054
rect 43526 -51087 43542 -51070
rect 43080 -51104 43282 -51087
rect 42322 -51142 43282 -51104
rect 43340 -51104 43542 -51087
rect 44098 -51087 44114 -51070
rect 44544 -51070 45132 -51054
rect 44544 -51087 44560 -51070
rect 44098 -51104 44300 -51087
rect 43340 -51142 44300 -51104
rect 44358 -51104 44560 -51087
rect 45116 -51087 45132 -51070
rect 45562 -51070 46150 -51054
rect 45562 -51087 45578 -51070
rect 45116 -51104 45318 -51087
rect 44358 -51142 45318 -51104
rect 45376 -51104 45578 -51087
rect 46134 -51087 46150 -51070
rect 46580 -51070 47168 -51054
rect 46580 -51087 46596 -51070
rect 46134 -51104 46336 -51087
rect 45376 -51142 46336 -51104
rect 46394 -51104 46596 -51087
rect 47152 -51087 47168 -51070
rect 47598 -51070 48186 -51054
rect 47598 -51087 47614 -51070
rect 47152 -51104 47354 -51087
rect 46394 -51142 47354 -51104
rect 47412 -51104 47614 -51087
rect 48170 -51087 48186 -51070
rect 48170 -51104 48372 -51087
rect 47412 -51142 48372 -51104
rect 28070 -51780 29030 -51742
rect 28070 -51797 28272 -51780
rect 28256 -51814 28272 -51797
rect 28828 -51797 29030 -51780
rect 29088 -51780 30048 -51742
rect 29088 -51797 29290 -51780
rect 28828 -51814 28844 -51797
rect 28256 -51830 28844 -51814
rect 29274 -51814 29290 -51797
rect 29846 -51797 30048 -51780
rect 30106 -51780 31066 -51742
rect 30106 -51797 30308 -51780
rect 29846 -51814 29862 -51797
rect 29274 -51830 29862 -51814
rect 30292 -51814 30308 -51797
rect 30864 -51797 31066 -51780
rect 31124 -51780 32084 -51742
rect 31124 -51797 31326 -51780
rect 30864 -51814 30880 -51797
rect 30292 -51830 30880 -51814
rect 31310 -51814 31326 -51797
rect 31882 -51797 32084 -51780
rect 32142 -51780 33102 -51742
rect 32142 -51797 32344 -51780
rect 31882 -51814 31898 -51797
rect 31310 -51830 31898 -51814
rect 32328 -51814 32344 -51797
rect 32900 -51797 33102 -51780
rect 33160 -51780 34120 -51742
rect 33160 -51797 33362 -51780
rect 32900 -51814 32916 -51797
rect 32328 -51830 32916 -51814
rect 33346 -51814 33362 -51797
rect 33918 -51797 34120 -51780
rect 34178 -51780 35138 -51742
rect 34178 -51797 34380 -51780
rect 33918 -51814 33934 -51797
rect 33346 -51830 33934 -51814
rect 34364 -51814 34380 -51797
rect 34936 -51797 35138 -51780
rect 35196 -51780 36156 -51742
rect 35196 -51797 35398 -51780
rect 34936 -51814 34952 -51797
rect 34364 -51830 34952 -51814
rect 35382 -51814 35398 -51797
rect 35954 -51797 36156 -51780
rect 36214 -51780 37174 -51742
rect 36214 -51797 36416 -51780
rect 35954 -51814 35970 -51797
rect 35382 -51830 35970 -51814
rect 36400 -51814 36416 -51797
rect 36972 -51797 37174 -51780
rect 37232 -51780 38192 -51742
rect 37232 -51797 37434 -51780
rect 36972 -51814 36988 -51797
rect 36400 -51830 36988 -51814
rect 37418 -51814 37434 -51797
rect 37990 -51797 38192 -51780
rect 38250 -51780 39210 -51742
rect 38250 -51797 38452 -51780
rect 37990 -51814 38006 -51797
rect 37418 -51830 38006 -51814
rect 38436 -51814 38452 -51797
rect 39008 -51797 39210 -51780
rect 39268 -51780 40228 -51742
rect 39268 -51797 39470 -51780
rect 39008 -51814 39024 -51797
rect 38436 -51830 39024 -51814
rect 39454 -51814 39470 -51797
rect 40026 -51797 40228 -51780
rect 40286 -51780 41246 -51742
rect 40286 -51797 40488 -51780
rect 40026 -51814 40042 -51797
rect 39454 -51830 40042 -51814
rect 40472 -51814 40488 -51797
rect 41044 -51797 41246 -51780
rect 41304 -51780 42264 -51742
rect 41304 -51797 41506 -51780
rect 41044 -51814 41060 -51797
rect 40472 -51830 41060 -51814
rect 41490 -51814 41506 -51797
rect 42062 -51797 42264 -51780
rect 42322 -51780 43282 -51742
rect 42322 -51797 42524 -51780
rect 42062 -51814 42078 -51797
rect 41490 -51830 42078 -51814
rect 42508 -51814 42524 -51797
rect 43080 -51797 43282 -51780
rect 43340 -51780 44300 -51742
rect 43340 -51797 43542 -51780
rect 43080 -51814 43096 -51797
rect 42508 -51830 43096 -51814
rect 43526 -51814 43542 -51797
rect 44098 -51797 44300 -51780
rect 44358 -51780 45318 -51742
rect 44358 -51797 44560 -51780
rect 44098 -51814 44114 -51797
rect 43526 -51830 44114 -51814
rect 44544 -51814 44560 -51797
rect 45116 -51797 45318 -51780
rect 45376 -51780 46336 -51742
rect 45376 -51797 45578 -51780
rect 45116 -51814 45132 -51797
rect 44544 -51830 45132 -51814
rect 45562 -51814 45578 -51797
rect 46134 -51797 46336 -51780
rect 46394 -51780 47354 -51742
rect 46394 -51797 46596 -51780
rect 46134 -51814 46150 -51797
rect 45562 -51830 46150 -51814
rect 46580 -51814 46596 -51797
rect 47152 -51797 47354 -51780
rect 47412 -51780 48372 -51742
rect 47412 -51797 47614 -51780
rect 47152 -51814 47168 -51797
rect 46580 -51830 47168 -51814
rect 47598 -51814 47614 -51797
rect 48170 -51797 48372 -51780
rect 48170 -51814 48186 -51797
rect 47598 -51830 48186 -51814
rect 15168 -52168 15756 -52152
rect 15168 -52185 15184 -52168
rect 14982 -52202 15184 -52185
rect 15740 -52185 15756 -52168
rect 16186 -52168 16774 -52152
rect 16186 -52185 16202 -52168
rect 15740 -52202 15942 -52185
rect 14982 -52240 15942 -52202
rect 16000 -52202 16202 -52185
rect 16758 -52185 16774 -52168
rect 17204 -52168 17792 -52152
rect 17204 -52185 17220 -52168
rect 16758 -52202 16960 -52185
rect 16000 -52240 16960 -52202
rect 17018 -52202 17220 -52185
rect 17776 -52185 17792 -52168
rect 18222 -52168 18810 -52152
rect 18222 -52185 18238 -52168
rect 17776 -52202 17978 -52185
rect 17018 -52240 17978 -52202
rect 18036 -52202 18238 -52185
rect 18794 -52185 18810 -52168
rect 19240 -52168 19828 -52152
rect 19240 -52185 19256 -52168
rect 18794 -52202 18996 -52185
rect 18036 -52240 18996 -52202
rect 19054 -52202 19256 -52185
rect 19812 -52185 19828 -52168
rect 20258 -52168 20846 -52152
rect 20258 -52185 20274 -52168
rect 19812 -52202 20014 -52185
rect 19054 -52240 20014 -52202
rect 20072 -52202 20274 -52185
rect 20830 -52185 20846 -52168
rect 21276 -52168 21864 -52152
rect 21276 -52185 21292 -52168
rect 20830 -52202 21032 -52185
rect 20072 -52240 21032 -52202
rect 21090 -52202 21292 -52185
rect 21848 -52185 21864 -52168
rect 22294 -52168 22882 -52152
rect 22294 -52185 22310 -52168
rect 21848 -52202 22050 -52185
rect 21090 -52240 22050 -52202
rect 22108 -52202 22310 -52185
rect 22866 -52185 22882 -52168
rect 23312 -52168 23900 -52152
rect 23312 -52185 23328 -52168
rect 22866 -52202 23068 -52185
rect 22108 -52240 23068 -52202
rect 23126 -52202 23328 -52185
rect 23884 -52185 23900 -52168
rect 24330 -52168 24918 -52152
rect 24330 -52185 24346 -52168
rect 23884 -52202 24086 -52185
rect 23126 -52240 24086 -52202
rect 24144 -52202 24346 -52185
rect 24902 -52185 24918 -52168
rect 25348 -52168 25936 -52152
rect 25348 -52185 25364 -52168
rect 24902 -52202 25104 -52185
rect 24144 -52240 25104 -52202
rect 25162 -52202 25364 -52185
rect 25920 -52185 25936 -52168
rect 25920 -52202 26122 -52185
rect 25162 -52240 26122 -52202
rect 28256 -52304 28844 -52288
rect 28256 -52321 28272 -52304
rect 28070 -52338 28272 -52321
rect 28828 -52321 28844 -52304
rect 29274 -52304 29862 -52288
rect 29274 -52321 29290 -52304
rect 28828 -52338 29030 -52321
rect 28070 -52376 29030 -52338
rect 29088 -52338 29290 -52321
rect 29846 -52321 29862 -52304
rect 30292 -52304 30880 -52288
rect 30292 -52321 30308 -52304
rect 29846 -52338 30048 -52321
rect 29088 -52376 30048 -52338
rect 30106 -52338 30308 -52321
rect 30864 -52321 30880 -52304
rect 31310 -52304 31898 -52288
rect 31310 -52321 31326 -52304
rect 30864 -52338 31066 -52321
rect 30106 -52376 31066 -52338
rect 31124 -52338 31326 -52321
rect 31882 -52321 31898 -52304
rect 32328 -52304 32916 -52288
rect 32328 -52321 32344 -52304
rect 31882 -52338 32084 -52321
rect 31124 -52376 32084 -52338
rect 32142 -52338 32344 -52321
rect 32900 -52321 32916 -52304
rect 33346 -52304 33934 -52288
rect 33346 -52321 33362 -52304
rect 32900 -52338 33102 -52321
rect 32142 -52376 33102 -52338
rect 33160 -52338 33362 -52321
rect 33918 -52321 33934 -52304
rect 34364 -52304 34952 -52288
rect 34364 -52321 34380 -52304
rect 33918 -52338 34120 -52321
rect 33160 -52376 34120 -52338
rect 34178 -52338 34380 -52321
rect 34936 -52321 34952 -52304
rect 35382 -52304 35970 -52288
rect 35382 -52321 35398 -52304
rect 34936 -52338 35138 -52321
rect 34178 -52376 35138 -52338
rect 35196 -52338 35398 -52321
rect 35954 -52321 35970 -52304
rect 36400 -52304 36988 -52288
rect 36400 -52321 36416 -52304
rect 35954 -52338 36156 -52321
rect 35196 -52376 36156 -52338
rect 36214 -52338 36416 -52321
rect 36972 -52321 36988 -52304
rect 37418 -52304 38006 -52288
rect 37418 -52321 37434 -52304
rect 36972 -52338 37174 -52321
rect 36214 -52376 37174 -52338
rect 37232 -52338 37434 -52321
rect 37990 -52321 38006 -52304
rect 38436 -52304 39024 -52288
rect 38436 -52321 38452 -52304
rect 37990 -52338 38192 -52321
rect 37232 -52376 38192 -52338
rect 38250 -52338 38452 -52321
rect 39008 -52321 39024 -52304
rect 39454 -52304 40042 -52288
rect 39454 -52321 39470 -52304
rect 39008 -52338 39210 -52321
rect 38250 -52376 39210 -52338
rect 39268 -52338 39470 -52321
rect 40026 -52321 40042 -52304
rect 40472 -52304 41060 -52288
rect 40472 -52321 40488 -52304
rect 40026 -52338 40228 -52321
rect 39268 -52376 40228 -52338
rect 40286 -52338 40488 -52321
rect 41044 -52321 41060 -52304
rect 41490 -52304 42078 -52288
rect 41490 -52321 41506 -52304
rect 41044 -52338 41246 -52321
rect 40286 -52376 41246 -52338
rect 41304 -52338 41506 -52321
rect 42062 -52321 42078 -52304
rect 42508 -52304 43096 -52288
rect 42508 -52321 42524 -52304
rect 42062 -52338 42264 -52321
rect 41304 -52376 42264 -52338
rect 42322 -52338 42524 -52321
rect 43080 -52321 43096 -52304
rect 43526 -52304 44114 -52288
rect 43526 -52321 43542 -52304
rect 43080 -52338 43282 -52321
rect 42322 -52376 43282 -52338
rect 43340 -52338 43542 -52321
rect 44098 -52321 44114 -52304
rect 44544 -52304 45132 -52288
rect 44544 -52321 44560 -52304
rect 44098 -52338 44300 -52321
rect 43340 -52376 44300 -52338
rect 44358 -52338 44560 -52321
rect 45116 -52321 45132 -52304
rect 45562 -52304 46150 -52288
rect 45562 -52321 45578 -52304
rect 45116 -52338 45318 -52321
rect 44358 -52376 45318 -52338
rect 45376 -52338 45578 -52321
rect 46134 -52321 46150 -52304
rect 46580 -52304 47168 -52288
rect 46580 -52321 46596 -52304
rect 46134 -52338 46336 -52321
rect 45376 -52376 46336 -52338
rect 46394 -52338 46596 -52321
rect 47152 -52321 47168 -52304
rect 47598 -52304 48186 -52288
rect 47598 -52321 47614 -52304
rect 47152 -52338 47354 -52321
rect 46394 -52376 47354 -52338
rect 47412 -52338 47614 -52321
rect 48170 -52321 48186 -52304
rect 48170 -52338 48372 -52321
rect 47412 -52376 48372 -52338
rect 14982 -52878 15942 -52840
rect 14982 -52895 15184 -52878
rect 15168 -52912 15184 -52895
rect 15740 -52895 15942 -52878
rect 16000 -52878 16960 -52840
rect 16000 -52895 16202 -52878
rect 15740 -52912 15756 -52895
rect 15168 -52928 15756 -52912
rect 16186 -52912 16202 -52895
rect 16758 -52895 16960 -52878
rect 17018 -52878 17978 -52840
rect 17018 -52895 17220 -52878
rect 16758 -52912 16774 -52895
rect 16186 -52928 16774 -52912
rect 17204 -52912 17220 -52895
rect 17776 -52895 17978 -52878
rect 18036 -52878 18996 -52840
rect 18036 -52895 18238 -52878
rect 17776 -52912 17792 -52895
rect 17204 -52928 17792 -52912
rect 18222 -52912 18238 -52895
rect 18794 -52895 18996 -52878
rect 19054 -52878 20014 -52840
rect 19054 -52895 19256 -52878
rect 18794 -52912 18810 -52895
rect 18222 -52928 18810 -52912
rect 19240 -52912 19256 -52895
rect 19812 -52895 20014 -52878
rect 20072 -52878 21032 -52840
rect 20072 -52895 20274 -52878
rect 19812 -52912 19828 -52895
rect 19240 -52928 19828 -52912
rect 20258 -52912 20274 -52895
rect 20830 -52895 21032 -52878
rect 21090 -52878 22050 -52840
rect 21090 -52895 21292 -52878
rect 20830 -52912 20846 -52895
rect 20258 -52928 20846 -52912
rect 21276 -52912 21292 -52895
rect 21848 -52895 22050 -52878
rect 22108 -52878 23068 -52840
rect 22108 -52895 22310 -52878
rect 21848 -52912 21864 -52895
rect 21276 -52928 21864 -52912
rect 22294 -52912 22310 -52895
rect 22866 -52895 23068 -52878
rect 23126 -52878 24086 -52840
rect 23126 -52895 23328 -52878
rect 22866 -52912 22882 -52895
rect 22294 -52928 22882 -52912
rect 23312 -52912 23328 -52895
rect 23884 -52895 24086 -52878
rect 24144 -52878 25104 -52840
rect 24144 -52895 24346 -52878
rect 23884 -52912 23900 -52895
rect 23312 -52928 23900 -52912
rect 24330 -52912 24346 -52895
rect 24902 -52895 25104 -52878
rect 25162 -52878 26122 -52840
rect 25162 -52895 25364 -52878
rect 24902 -52912 24918 -52895
rect 24330 -52928 24918 -52912
rect 25348 -52912 25364 -52895
rect 25920 -52895 26122 -52878
rect 25920 -52912 25936 -52895
rect 25348 -52928 25936 -52912
rect 28070 -53014 29030 -52976
rect 28070 -53031 28272 -53014
rect 28256 -53048 28272 -53031
rect 28828 -53031 29030 -53014
rect 29088 -53014 30048 -52976
rect 29088 -53031 29290 -53014
rect 28828 -53048 28844 -53031
rect 28256 -53064 28844 -53048
rect 29274 -53048 29290 -53031
rect 29846 -53031 30048 -53014
rect 30106 -53014 31066 -52976
rect 30106 -53031 30308 -53014
rect 29846 -53048 29862 -53031
rect 29274 -53064 29862 -53048
rect 30292 -53048 30308 -53031
rect 30864 -53031 31066 -53014
rect 31124 -53014 32084 -52976
rect 31124 -53031 31326 -53014
rect 30864 -53048 30880 -53031
rect 30292 -53064 30880 -53048
rect 31310 -53048 31326 -53031
rect 31882 -53031 32084 -53014
rect 32142 -53014 33102 -52976
rect 32142 -53031 32344 -53014
rect 31882 -53048 31898 -53031
rect 31310 -53064 31898 -53048
rect 32328 -53048 32344 -53031
rect 32900 -53031 33102 -53014
rect 33160 -53014 34120 -52976
rect 33160 -53031 33362 -53014
rect 32900 -53048 32916 -53031
rect 32328 -53064 32916 -53048
rect 33346 -53048 33362 -53031
rect 33918 -53031 34120 -53014
rect 34178 -53014 35138 -52976
rect 34178 -53031 34380 -53014
rect 33918 -53048 33934 -53031
rect 33346 -53064 33934 -53048
rect 34364 -53048 34380 -53031
rect 34936 -53031 35138 -53014
rect 35196 -53014 36156 -52976
rect 35196 -53031 35398 -53014
rect 34936 -53048 34952 -53031
rect 34364 -53064 34952 -53048
rect 35382 -53048 35398 -53031
rect 35954 -53031 36156 -53014
rect 36214 -53014 37174 -52976
rect 36214 -53031 36416 -53014
rect 35954 -53048 35970 -53031
rect 35382 -53064 35970 -53048
rect 36400 -53048 36416 -53031
rect 36972 -53031 37174 -53014
rect 37232 -53014 38192 -52976
rect 37232 -53031 37434 -53014
rect 36972 -53048 36988 -53031
rect 36400 -53064 36988 -53048
rect 37418 -53048 37434 -53031
rect 37990 -53031 38192 -53014
rect 38250 -53014 39210 -52976
rect 38250 -53031 38452 -53014
rect 37990 -53048 38006 -53031
rect 37418 -53064 38006 -53048
rect 38436 -53048 38452 -53031
rect 39008 -53031 39210 -53014
rect 39268 -53014 40228 -52976
rect 39268 -53031 39470 -53014
rect 39008 -53048 39024 -53031
rect 38436 -53064 39024 -53048
rect 39454 -53048 39470 -53031
rect 40026 -53031 40228 -53014
rect 40286 -53014 41246 -52976
rect 40286 -53031 40488 -53014
rect 40026 -53048 40042 -53031
rect 39454 -53064 40042 -53048
rect 40472 -53048 40488 -53031
rect 41044 -53031 41246 -53014
rect 41304 -53014 42264 -52976
rect 41304 -53031 41506 -53014
rect 41044 -53048 41060 -53031
rect 40472 -53064 41060 -53048
rect 41490 -53048 41506 -53031
rect 42062 -53031 42264 -53014
rect 42322 -53014 43282 -52976
rect 42322 -53031 42524 -53014
rect 42062 -53048 42078 -53031
rect 41490 -53064 42078 -53048
rect 42508 -53048 42524 -53031
rect 43080 -53031 43282 -53014
rect 43340 -53014 44300 -52976
rect 43340 -53031 43542 -53014
rect 43080 -53048 43096 -53031
rect 42508 -53064 43096 -53048
rect 43526 -53048 43542 -53031
rect 44098 -53031 44300 -53014
rect 44358 -53014 45318 -52976
rect 44358 -53031 44560 -53014
rect 44098 -53048 44114 -53031
rect 43526 -53064 44114 -53048
rect 44544 -53048 44560 -53031
rect 45116 -53031 45318 -53014
rect 45376 -53014 46336 -52976
rect 45376 -53031 45578 -53014
rect 45116 -53048 45132 -53031
rect 44544 -53064 45132 -53048
rect 45562 -53048 45578 -53031
rect 46134 -53031 46336 -53014
rect 46394 -53014 47354 -52976
rect 46394 -53031 46596 -53014
rect 46134 -53048 46150 -53031
rect 45562 -53064 46150 -53048
rect 46580 -53048 46596 -53031
rect 47152 -53031 47354 -53014
rect 47412 -53014 48372 -52976
rect 47412 -53031 47614 -53014
rect 47152 -53048 47168 -53031
rect 46580 -53064 47168 -53048
rect 47598 -53048 47614 -53031
rect 48170 -53031 48372 -53014
rect 48170 -53048 48186 -53031
rect 47598 -53064 48186 -53048
rect 15168 -53280 15756 -53264
rect 15168 -53297 15184 -53280
rect 14982 -53314 15184 -53297
rect 15740 -53297 15756 -53280
rect 16186 -53280 16774 -53264
rect 16186 -53297 16202 -53280
rect 15740 -53314 15942 -53297
rect 14982 -53352 15942 -53314
rect 16000 -53314 16202 -53297
rect 16758 -53297 16774 -53280
rect 17204 -53280 17792 -53264
rect 17204 -53297 17220 -53280
rect 16758 -53314 16960 -53297
rect 16000 -53352 16960 -53314
rect 17018 -53314 17220 -53297
rect 17776 -53297 17792 -53280
rect 18222 -53280 18810 -53264
rect 18222 -53297 18238 -53280
rect 17776 -53314 17978 -53297
rect 17018 -53352 17978 -53314
rect 18036 -53314 18238 -53297
rect 18794 -53297 18810 -53280
rect 19240 -53280 19828 -53264
rect 19240 -53297 19256 -53280
rect 18794 -53314 18996 -53297
rect 18036 -53352 18996 -53314
rect 19054 -53314 19256 -53297
rect 19812 -53297 19828 -53280
rect 20258 -53280 20846 -53264
rect 20258 -53297 20274 -53280
rect 19812 -53314 20014 -53297
rect 19054 -53352 20014 -53314
rect 20072 -53314 20274 -53297
rect 20830 -53297 20846 -53280
rect 21276 -53280 21864 -53264
rect 21276 -53297 21292 -53280
rect 20830 -53314 21032 -53297
rect 20072 -53352 21032 -53314
rect 21090 -53314 21292 -53297
rect 21848 -53297 21864 -53280
rect 22294 -53280 22882 -53264
rect 22294 -53297 22310 -53280
rect 21848 -53314 22050 -53297
rect 21090 -53352 22050 -53314
rect 22108 -53314 22310 -53297
rect 22866 -53297 22882 -53280
rect 23312 -53280 23900 -53264
rect 23312 -53297 23328 -53280
rect 22866 -53314 23068 -53297
rect 22108 -53352 23068 -53314
rect 23126 -53314 23328 -53297
rect 23884 -53297 23900 -53280
rect 24330 -53280 24918 -53264
rect 24330 -53297 24346 -53280
rect 23884 -53314 24086 -53297
rect 23126 -53352 24086 -53314
rect 24144 -53314 24346 -53297
rect 24902 -53297 24918 -53280
rect 25348 -53280 25936 -53264
rect 25348 -53297 25364 -53280
rect 24902 -53314 25104 -53297
rect 24144 -53352 25104 -53314
rect 25162 -53314 25364 -53297
rect 25920 -53297 25936 -53280
rect 25920 -53314 26122 -53297
rect 25162 -53352 26122 -53314
rect 28256 -53538 28844 -53522
rect 28256 -53555 28272 -53538
rect 28070 -53572 28272 -53555
rect 28828 -53555 28844 -53538
rect 29274 -53538 29862 -53522
rect 29274 -53555 29290 -53538
rect 28828 -53572 29030 -53555
rect 28070 -53610 29030 -53572
rect 29088 -53572 29290 -53555
rect 29846 -53555 29862 -53538
rect 30292 -53538 30880 -53522
rect 30292 -53555 30308 -53538
rect 29846 -53572 30048 -53555
rect 29088 -53610 30048 -53572
rect 30106 -53572 30308 -53555
rect 30864 -53555 30880 -53538
rect 31310 -53538 31898 -53522
rect 31310 -53555 31326 -53538
rect 30864 -53572 31066 -53555
rect 30106 -53610 31066 -53572
rect 31124 -53572 31326 -53555
rect 31882 -53555 31898 -53538
rect 32328 -53538 32916 -53522
rect 32328 -53555 32344 -53538
rect 31882 -53572 32084 -53555
rect 31124 -53610 32084 -53572
rect 32142 -53572 32344 -53555
rect 32900 -53555 32916 -53538
rect 33346 -53538 33934 -53522
rect 33346 -53555 33362 -53538
rect 32900 -53572 33102 -53555
rect 32142 -53610 33102 -53572
rect 33160 -53572 33362 -53555
rect 33918 -53555 33934 -53538
rect 34364 -53538 34952 -53522
rect 34364 -53555 34380 -53538
rect 33918 -53572 34120 -53555
rect 33160 -53610 34120 -53572
rect 34178 -53572 34380 -53555
rect 34936 -53555 34952 -53538
rect 35382 -53538 35970 -53522
rect 35382 -53555 35398 -53538
rect 34936 -53572 35138 -53555
rect 34178 -53610 35138 -53572
rect 35196 -53572 35398 -53555
rect 35954 -53555 35970 -53538
rect 36400 -53538 36988 -53522
rect 36400 -53555 36416 -53538
rect 35954 -53572 36156 -53555
rect 35196 -53610 36156 -53572
rect 36214 -53572 36416 -53555
rect 36972 -53555 36988 -53538
rect 37418 -53538 38006 -53522
rect 37418 -53555 37434 -53538
rect 36972 -53572 37174 -53555
rect 36214 -53610 37174 -53572
rect 37232 -53572 37434 -53555
rect 37990 -53555 38006 -53538
rect 38436 -53538 39024 -53522
rect 38436 -53555 38452 -53538
rect 37990 -53572 38192 -53555
rect 37232 -53610 38192 -53572
rect 38250 -53572 38452 -53555
rect 39008 -53555 39024 -53538
rect 39454 -53538 40042 -53522
rect 39454 -53555 39470 -53538
rect 39008 -53572 39210 -53555
rect 38250 -53610 39210 -53572
rect 39268 -53572 39470 -53555
rect 40026 -53555 40042 -53538
rect 40472 -53538 41060 -53522
rect 40472 -53555 40488 -53538
rect 40026 -53572 40228 -53555
rect 39268 -53610 40228 -53572
rect 40286 -53572 40488 -53555
rect 41044 -53555 41060 -53538
rect 41490 -53538 42078 -53522
rect 41490 -53555 41506 -53538
rect 41044 -53572 41246 -53555
rect 40286 -53610 41246 -53572
rect 41304 -53572 41506 -53555
rect 42062 -53555 42078 -53538
rect 42508 -53538 43096 -53522
rect 42508 -53555 42524 -53538
rect 42062 -53572 42264 -53555
rect 41304 -53610 42264 -53572
rect 42322 -53572 42524 -53555
rect 43080 -53555 43096 -53538
rect 43526 -53538 44114 -53522
rect 43526 -53555 43542 -53538
rect 43080 -53572 43282 -53555
rect 42322 -53610 43282 -53572
rect 43340 -53572 43542 -53555
rect 44098 -53555 44114 -53538
rect 44544 -53538 45132 -53522
rect 44544 -53555 44560 -53538
rect 44098 -53572 44300 -53555
rect 43340 -53610 44300 -53572
rect 44358 -53572 44560 -53555
rect 45116 -53555 45132 -53538
rect 45562 -53538 46150 -53522
rect 45562 -53555 45578 -53538
rect 45116 -53572 45318 -53555
rect 44358 -53610 45318 -53572
rect 45376 -53572 45578 -53555
rect 46134 -53555 46150 -53538
rect 46580 -53538 47168 -53522
rect 46580 -53555 46596 -53538
rect 46134 -53572 46336 -53555
rect 45376 -53610 46336 -53572
rect 46394 -53572 46596 -53555
rect 47152 -53555 47168 -53538
rect 47598 -53538 48186 -53522
rect 47598 -53555 47614 -53538
rect 47152 -53572 47354 -53555
rect 46394 -53610 47354 -53572
rect 47412 -53572 47614 -53555
rect 48170 -53555 48186 -53538
rect 48170 -53572 48372 -53555
rect 47412 -53610 48372 -53572
rect 14982 -53990 15942 -53952
rect 14982 -54007 15184 -53990
rect 15168 -54024 15184 -54007
rect 15740 -54007 15942 -53990
rect 16000 -53990 16960 -53952
rect 16000 -54007 16202 -53990
rect 15740 -54024 15756 -54007
rect 15168 -54040 15756 -54024
rect 16186 -54024 16202 -54007
rect 16758 -54007 16960 -53990
rect 17018 -53990 17978 -53952
rect 17018 -54007 17220 -53990
rect 16758 -54024 16774 -54007
rect 16186 -54040 16774 -54024
rect 17204 -54024 17220 -54007
rect 17776 -54007 17978 -53990
rect 18036 -53990 18996 -53952
rect 18036 -54007 18238 -53990
rect 17776 -54024 17792 -54007
rect 17204 -54040 17792 -54024
rect 18222 -54024 18238 -54007
rect 18794 -54007 18996 -53990
rect 19054 -53990 20014 -53952
rect 19054 -54007 19256 -53990
rect 18794 -54024 18810 -54007
rect 18222 -54040 18810 -54024
rect 19240 -54024 19256 -54007
rect 19812 -54007 20014 -53990
rect 20072 -53990 21032 -53952
rect 20072 -54007 20274 -53990
rect 19812 -54024 19828 -54007
rect 19240 -54040 19828 -54024
rect 20258 -54024 20274 -54007
rect 20830 -54007 21032 -53990
rect 21090 -53990 22050 -53952
rect 21090 -54007 21292 -53990
rect 20830 -54024 20846 -54007
rect 20258 -54040 20846 -54024
rect 21276 -54024 21292 -54007
rect 21848 -54007 22050 -53990
rect 22108 -53990 23068 -53952
rect 22108 -54007 22310 -53990
rect 21848 -54024 21864 -54007
rect 21276 -54040 21864 -54024
rect 22294 -54024 22310 -54007
rect 22866 -54007 23068 -53990
rect 23126 -53990 24086 -53952
rect 23126 -54007 23328 -53990
rect 22866 -54024 22882 -54007
rect 22294 -54040 22882 -54024
rect 23312 -54024 23328 -54007
rect 23884 -54007 24086 -53990
rect 24144 -53990 25104 -53952
rect 24144 -54007 24346 -53990
rect 23884 -54024 23900 -54007
rect 23312 -54040 23900 -54024
rect 24330 -54024 24346 -54007
rect 24902 -54007 25104 -53990
rect 25162 -53990 26122 -53952
rect 25162 -54007 25364 -53990
rect 24902 -54024 24918 -54007
rect 24330 -54040 24918 -54024
rect 25348 -54024 25364 -54007
rect 25920 -54007 26122 -53990
rect 25920 -54024 25936 -54007
rect 25348 -54040 25936 -54024
rect 28070 -54248 29030 -54210
rect 28070 -54265 28272 -54248
rect 28256 -54282 28272 -54265
rect 28828 -54265 29030 -54248
rect 29088 -54248 30048 -54210
rect 29088 -54265 29290 -54248
rect 28828 -54282 28844 -54265
rect 28256 -54298 28844 -54282
rect 29274 -54282 29290 -54265
rect 29846 -54265 30048 -54248
rect 30106 -54248 31066 -54210
rect 30106 -54265 30308 -54248
rect 29846 -54282 29862 -54265
rect 29274 -54298 29862 -54282
rect 30292 -54282 30308 -54265
rect 30864 -54265 31066 -54248
rect 31124 -54248 32084 -54210
rect 31124 -54265 31326 -54248
rect 30864 -54282 30880 -54265
rect 30292 -54298 30880 -54282
rect 31310 -54282 31326 -54265
rect 31882 -54265 32084 -54248
rect 32142 -54248 33102 -54210
rect 32142 -54265 32344 -54248
rect 31882 -54282 31898 -54265
rect 31310 -54298 31898 -54282
rect 32328 -54282 32344 -54265
rect 32900 -54265 33102 -54248
rect 33160 -54248 34120 -54210
rect 33160 -54265 33362 -54248
rect 32900 -54282 32916 -54265
rect 32328 -54298 32916 -54282
rect 33346 -54282 33362 -54265
rect 33918 -54265 34120 -54248
rect 34178 -54248 35138 -54210
rect 34178 -54265 34380 -54248
rect 33918 -54282 33934 -54265
rect 33346 -54298 33934 -54282
rect 34364 -54282 34380 -54265
rect 34936 -54265 35138 -54248
rect 35196 -54248 36156 -54210
rect 35196 -54265 35398 -54248
rect 34936 -54282 34952 -54265
rect 34364 -54298 34952 -54282
rect 35382 -54282 35398 -54265
rect 35954 -54265 36156 -54248
rect 36214 -54248 37174 -54210
rect 36214 -54265 36416 -54248
rect 35954 -54282 35970 -54265
rect 35382 -54298 35970 -54282
rect 36400 -54282 36416 -54265
rect 36972 -54265 37174 -54248
rect 37232 -54248 38192 -54210
rect 37232 -54265 37434 -54248
rect 36972 -54282 36988 -54265
rect 36400 -54298 36988 -54282
rect 37418 -54282 37434 -54265
rect 37990 -54265 38192 -54248
rect 38250 -54248 39210 -54210
rect 38250 -54265 38452 -54248
rect 37990 -54282 38006 -54265
rect 37418 -54298 38006 -54282
rect 38436 -54282 38452 -54265
rect 39008 -54265 39210 -54248
rect 39268 -54248 40228 -54210
rect 39268 -54265 39470 -54248
rect 39008 -54282 39024 -54265
rect 38436 -54298 39024 -54282
rect 39454 -54282 39470 -54265
rect 40026 -54265 40228 -54248
rect 40286 -54248 41246 -54210
rect 40286 -54265 40488 -54248
rect 40026 -54282 40042 -54265
rect 39454 -54298 40042 -54282
rect 40472 -54282 40488 -54265
rect 41044 -54265 41246 -54248
rect 41304 -54248 42264 -54210
rect 41304 -54265 41506 -54248
rect 41044 -54282 41060 -54265
rect 40472 -54298 41060 -54282
rect 41490 -54282 41506 -54265
rect 42062 -54265 42264 -54248
rect 42322 -54248 43282 -54210
rect 42322 -54265 42524 -54248
rect 42062 -54282 42078 -54265
rect 41490 -54298 42078 -54282
rect 42508 -54282 42524 -54265
rect 43080 -54265 43282 -54248
rect 43340 -54248 44300 -54210
rect 43340 -54265 43542 -54248
rect 43080 -54282 43096 -54265
rect 42508 -54298 43096 -54282
rect 43526 -54282 43542 -54265
rect 44098 -54265 44300 -54248
rect 44358 -54248 45318 -54210
rect 44358 -54265 44560 -54248
rect 44098 -54282 44114 -54265
rect 43526 -54298 44114 -54282
rect 44544 -54282 44560 -54265
rect 45116 -54265 45318 -54248
rect 45376 -54248 46336 -54210
rect 45376 -54265 45578 -54248
rect 45116 -54282 45132 -54265
rect 44544 -54298 45132 -54282
rect 45562 -54282 45578 -54265
rect 46134 -54265 46336 -54248
rect 46394 -54248 47354 -54210
rect 46394 -54265 46596 -54248
rect 46134 -54282 46150 -54265
rect 45562 -54298 46150 -54282
rect 46580 -54282 46596 -54265
rect 47152 -54265 47354 -54248
rect 47412 -54248 48372 -54210
rect 47412 -54265 47614 -54248
rect 47152 -54282 47168 -54265
rect 46580 -54298 47168 -54282
rect 47598 -54282 47614 -54265
rect 48170 -54265 48372 -54248
rect 48170 -54282 48186 -54265
rect 47598 -54298 48186 -54282
rect 15168 -54392 15756 -54376
rect 15168 -54409 15184 -54392
rect 14982 -54426 15184 -54409
rect 15740 -54409 15756 -54392
rect 16186 -54392 16774 -54376
rect 16186 -54409 16202 -54392
rect 15740 -54426 15942 -54409
rect 14982 -54464 15942 -54426
rect 16000 -54426 16202 -54409
rect 16758 -54409 16774 -54392
rect 17204 -54392 17792 -54376
rect 17204 -54409 17220 -54392
rect 16758 -54426 16960 -54409
rect 16000 -54464 16960 -54426
rect 17018 -54426 17220 -54409
rect 17776 -54409 17792 -54392
rect 18222 -54392 18810 -54376
rect 18222 -54409 18238 -54392
rect 17776 -54426 17978 -54409
rect 17018 -54464 17978 -54426
rect 18036 -54426 18238 -54409
rect 18794 -54409 18810 -54392
rect 19240 -54392 19828 -54376
rect 19240 -54409 19256 -54392
rect 18794 -54426 18996 -54409
rect 18036 -54464 18996 -54426
rect 19054 -54426 19256 -54409
rect 19812 -54409 19828 -54392
rect 20258 -54392 20846 -54376
rect 20258 -54409 20274 -54392
rect 19812 -54426 20014 -54409
rect 19054 -54464 20014 -54426
rect 20072 -54426 20274 -54409
rect 20830 -54409 20846 -54392
rect 21276 -54392 21864 -54376
rect 21276 -54409 21292 -54392
rect 20830 -54426 21032 -54409
rect 20072 -54464 21032 -54426
rect 21090 -54426 21292 -54409
rect 21848 -54409 21864 -54392
rect 22294 -54392 22882 -54376
rect 22294 -54409 22310 -54392
rect 21848 -54426 22050 -54409
rect 21090 -54464 22050 -54426
rect 22108 -54426 22310 -54409
rect 22866 -54409 22882 -54392
rect 23312 -54392 23900 -54376
rect 23312 -54409 23328 -54392
rect 22866 -54426 23068 -54409
rect 22108 -54464 23068 -54426
rect 23126 -54426 23328 -54409
rect 23884 -54409 23900 -54392
rect 24330 -54392 24918 -54376
rect 24330 -54409 24346 -54392
rect 23884 -54426 24086 -54409
rect 23126 -54464 24086 -54426
rect 24144 -54426 24346 -54409
rect 24902 -54409 24918 -54392
rect 25348 -54392 25936 -54376
rect 25348 -54409 25364 -54392
rect 24902 -54426 25104 -54409
rect 24144 -54464 25104 -54426
rect 25162 -54426 25364 -54409
rect 25920 -54409 25936 -54392
rect 25920 -54426 26122 -54409
rect 25162 -54464 26122 -54426
rect 28256 -54770 28844 -54754
rect 28256 -54787 28272 -54770
rect 28070 -54804 28272 -54787
rect 28828 -54787 28844 -54770
rect 29274 -54770 29862 -54754
rect 29274 -54787 29290 -54770
rect 28828 -54804 29030 -54787
rect 28070 -54842 29030 -54804
rect 29088 -54804 29290 -54787
rect 29846 -54787 29862 -54770
rect 30292 -54770 30880 -54754
rect 30292 -54787 30308 -54770
rect 29846 -54804 30048 -54787
rect 29088 -54842 30048 -54804
rect 30106 -54804 30308 -54787
rect 30864 -54787 30880 -54770
rect 31310 -54770 31898 -54754
rect 31310 -54787 31326 -54770
rect 30864 -54804 31066 -54787
rect 30106 -54842 31066 -54804
rect 31124 -54804 31326 -54787
rect 31882 -54787 31898 -54770
rect 32328 -54770 32916 -54754
rect 32328 -54787 32344 -54770
rect 31882 -54804 32084 -54787
rect 31124 -54842 32084 -54804
rect 32142 -54804 32344 -54787
rect 32900 -54787 32916 -54770
rect 33346 -54770 33934 -54754
rect 33346 -54787 33362 -54770
rect 32900 -54804 33102 -54787
rect 32142 -54842 33102 -54804
rect 33160 -54804 33362 -54787
rect 33918 -54787 33934 -54770
rect 34364 -54770 34952 -54754
rect 34364 -54787 34380 -54770
rect 33918 -54804 34120 -54787
rect 33160 -54842 34120 -54804
rect 34178 -54804 34380 -54787
rect 34936 -54787 34952 -54770
rect 35382 -54770 35970 -54754
rect 35382 -54787 35398 -54770
rect 34936 -54804 35138 -54787
rect 34178 -54842 35138 -54804
rect 35196 -54804 35398 -54787
rect 35954 -54787 35970 -54770
rect 36400 -54770 36988 -54754
rect 36400 -54787 36416 -54770
rect 35954 -54804 36156 -54787
rect 35196 -54842 36156 -54804
rect 36214 -54804 36416 -54787
rect 36972 -54787 36988 -54770
rect 37418 -54770 38006 -54754
rect 37418 -54787 37434 -54770
rect 36972 -54804 37174 -54787
rect 36214 -54842 37174 -54804
rect 37232 -54804 37434 -54787
rect 37990 -54787 38006 -54770
rect 38436 -54770 39024 -54754
rect 38436 -54787 38452 -54770
rect 37990 -54804 38192 -54787
rect 37232 -54842 38192 -54804
rect 38250 -54804 38452 -54787
rect 39008 -54787 39024 -54770
rect 39454 -54770 40042 -54754
rect 39454 -54787 39470 -54770
rect 39008 -54804 39210 -54787
rect 38250 -54842 39210 -54804
rect 39268 -54804 39470 -54787
rect 40026 -54787 40042 -54770
rect 40472 -54770 41060 -54754
rect 40472 -54787 40488 -54770
rect 40026 -54804 40228 -54787
rect 39268 -54842 40228 -54804
rect 40286 -54804 40488 -54787
rect 41044 -54787 41060 -54770
rect 41490 -54770 42078 -54754
rect 41490 -54787 41506 -54770
rect 41044 -54804 41246 -54787
rect 40286 -54842 41246 -54804
rect 41304 -54804 41506 -54787
rect 42062 -54787 42078 -54770
rect 42508 -54770 43096 -54754
rect 42508 -54787 42524 -54770
rect 42062 -54804 42264 -54787
rect 41304 -54842 42264 -54804
rect 42322 -54804 42524 -54787
rect 43080 -54787 43096 -54770
rect 43526 -54770 44114 -54754
rect 43526 -54787 43542 -54770
rect 43080 -54804 43282 -54787
rect 42322 -54842 43282 -54804
rect 43340 -54804 43542 -54787
rect 44098 -54787 44114 -54770
rect 44544 -54770 45132 -54754
rect 44544 -54787 44560 -54770
rect 44098 -54804 44300 -54787
rect 43340 -54842 44300 -54804
rect 44358 -54804 44560 -54787
rect 45116 -54787 45132 -54770
rect 45562 -54770 46150 -54754
rect 45562 -54787 45578 -54770
rect 45116 -54804 45318 -54787
rect 44358 -54842 45318 -54804
rect 45376 -54804 45578 -54787
rect 46134 -54787 46150 -54770
rect 46580 -54770 47168 -54754
rect 46580 -54787 46596 -54770
rect 46134 -54804 46336 -54787
rect 45376 -54842 46336 -54804
rect 46394 -54804 46596 -54787
rect 47152 -54787 47168 -54770
rect 47598 -54770 48186 -54754
rect 47598 -54787 47614 -54770
rect 47152 -54804 47354 -54787
rect 46394 -54842 47354 -54804
rect 47412 -54804 47614 -54787
rect 48170 -54787 48186 -54770
rect 48170 -54804 48372 -54787
rect 47412 -54842 48372 -54804
rect 14982 -55102 15942 -55064
rect 14982 -55119 15184 -55102
rect 15168 -55136 15184 -55119
rect 15740 -55119 15942 -55102
rect 16000 -55102 16960 -55064
rect 16000 -55119 16202 -55102
rect 15740 -55136 15756 -55119
rect 15168 -55152 15756 -55136
rect 16186 -55136 16202 -55119
rect 16758 -55119 16960 -55102
rect 17018 -55102 17978 -55064
rect 17018 -55119 17220 -55102
rect 16758 -55136 16774 -55119
rect 16186 -55152 16774 -55136
rect 17204 -55136 17220 -55119
rect 17776 -55119 17978 -55102
rect 18036 -55102 18996 -55064
rect 18036 -55119 18238 -55102
rect 17776 -55136 17792 -55119
rect 17204 -55152 17792 -55136
rect 18222 -55136 18238 -55119
rect 18794 -55119 18996 -55102
rect 19054 -55102 20014 -55064
rect 19054 -55119 19256 -55102
rect 18794 -55136 18810 -55119
rect 18222 -55152 18810 -55136
rect 19240 -55136 19256 -55119
rect 19812 -55119 20014 -55102
rect 20072 -55102 21032 -55064
rect 20072 -55119 20274 -55102
rect 19812 -55136 19828 -55119
rect 19240 -55152 19828 -55136
rect 20258 -55136 20274 -55119
rect 20830 -55119 21032 -55102
rect 21090 -55102 22050 -55064
rect 21090 -55119 21292 -55102
rect 20830 -55136 20846 -55119
rect 20258 -55152 20846 -55136
rect 21276 -55136 21292 -55119
rect 21848 -55119 22050 -55102
rect 22108 -55102 23068 -55064
rect 22108 -55119 22310 -55102
rect 21848 -55136 21864 -55119
rect 21276 -55152 21864 -55136
rect 22294 -55136 22310 -55119
rect 22866 -55119 23068 -55102
rect 23126 -55102 24086 -55064
rect 23126 -55119 23328 -55102
rect 22866 -55136 22882 -55119
rect 22294 -55152 22882 -55136
rect 23312 -55136 23328 -55119
rect 23884 -55119 24086 -55102
rect 24144 -55102 25104 -55064
rect 24144 -55119 24346 -55102
rect 23884 -55136 23900 -55119
rect 23312 -55152 23900 -55136
rect 24330 -55136 24346 -55119
rect 24902 -55119 25104 -55102
rect 25162 -55102 26122 -55064
rect 25162 -55119 25364 -55102
rect 24902 -55136 24918 -55119
rect 24330 -55152 24918 -55136
rect 25348 -55136 25364 -55119
rect 25920 -55119 26122 -55102
rect 25920 -55136 25936 -55119
rect 25348 -55152 25936 -55136
rect 28070 -55480 29030 -55442
rect 15168 -55504 15756 -55488
rect 15168 -55521 15184 -55504
rect 14982 -55538 15184 -55521
rect 15740 -55521 15756 -55504
rect 16186 -55504 16774 -55488
rect 16186 -55521 16202 -55504
rect 15740 -55538 15942 -55521
rect 14982 -55576 15942 -55538
rect 16000 -55538 16202 -55521
rect 16758 -55521 16774 -55504
rect 17204 -55504 17792 -55488
rect 17204 -55521 17220 -55504
rect 16758 -55538 16960 -55521
rect 16000 -55576 16960 -55538
rect 17018 -55538 17220 -55521
rect 17776 -55521 17792 -55504
rect 18222 -55504 18810 -55488
rect 18222 -55521 18238 -55504
rect 17776 -55538 17978 -55521
rect 17018 -55576 17978 -55538
rect 18036 -55538 18238 -55521
rect 18794 -55521 18810 -55504
rect 19240 -55504 19828 -55488
rect 19240 -55521 19256 -55504
rect 18794 -55538 18996 -55521
rect 18036 -55576 18996 -55538
rect 19054 -55538 19256 -55521
rect 19812 -55521 19828 -55504
rect 20258 -55504 20846 -55488
rect 20258 -55521 20274 -55504
rect 19812 -55538 20014 -55521
rect 19054 -55576 20014 -55538
rect 20072 -55538 20274 -55521
rect 20830 -55521 20846 -55504
rect 21276 -55504 21864 -55488
rect 21276 -55521 21292 -55504
rect 20830 -55538 21032 -55521
rect 20072 -55576 21032 -55538
rect 21090 -55538 21292 -55521
rect 21848 -55521 21864 -55504
rect 22294 -55504 22882 -55488
rect 22294 -55521 22310 -55504
rect 21848 -55538 22050 -55521
rect 21090 -55576 22050 -55538
rect 22108 -55538 22310 -55521
rect 22866 -55521 22882 -55504
rect 23312 -55504 23900 -55488
rect 23312 -55521 23328 -55504
rect 22866 -55538 23068 -55521
rect 22108 -55576 23068 -55538
rect 23126 -55538 23328 -55521
rect 23884 -55521 23900 -55504
rect 24330 -55504 24918 -55488
rect 24330 -55521 24346 -55504
rect 23884 -55538 24086 -55521
rect 23126 -55576 24086 -55538
rect 24144 -55538 24346 -55521
rect 24902 -55521 24918 -55504
rect 25348 -55504 25936 -55488
rect 28070 -55497 28272 -55480
rect 25348 -55521 25364 -55504
rect 24902 -55538 25104 -55521
rect 24144 -55576 25104 -55538
rect 25162 -55538 25364 -55521
rect 25920 -55521 25936 -55504
rect 28256 -55514 28272 -55497
rect 28828 -55497 29030 -55480
rect 29088 -55480 30048 -55442
rect 29088 -55497 29290 -55480
rect 28828 -55514 28844 -55497
rect 25920 -55538 26122 -55521
rect 28256 -55530 28844 -55514
rect 29274 -55514 29290 -55497
rect 29846 -55497 30048 -55480
rect 30106 -55480 31066 -55442
rect 30106 -55497 30308 -55480
rect 29846 -55514 29862 -55497
rect 29274 -55530 29862 -55514
rect 30292 -55514 30308 -55497
rect 30864 -55497 31066 -55480
rect 31124 -55480 32084 -55442
rect 31124 -55497 31326 -55480
rect 30864 -55514 30880 -55497
rect 30292 -55530 30880 -55514
rect 31310 -55514 31326 -55497
rect 31882 -55497 32084 -55480
rect 32142 -55480 33102 -55442
rect 32142 -55497 32344 -55480
rect 31882 -55514 31898 -55497
rect 31310 -55530 31898 -55514
rect 32328 -55514 32344 -55497
rect 32900 -55497 33102 -55480
rect 33160 -55480 34120 -55442
rect 33160 -55497 33362 -55480
rect 32900 -55514 32916 -55497
rect 32328 -55530 32916 -55514
rect 33346 -55514 33362 -55497
rect 33918 -55497 34120 -55480
rect 34178 -55480 35138 -55442
rect 34178 -55497 34380 -55480
rect 33918 -55514 33934 -55497
rect 33346 -55530 33934 -55514
rect 34364 -55514 34380 -55497
rect 34936 -55497 35138 -55480
rect 35196 -55480 36156 -55442
rect 35196 -55497 35398 -55480
rect 34936 -55514 34952 -55497
rect 34364 -55530 34952 -55514
rect 35382 -55514 35398 -55497
rect 35954 -55497 36156 -55480
rect 36214 -55480 37174 -55442
rect 36214 -55497 36416 -55480
rect 35954 -55514 35970 -55497
rect 35382 -55530 35970 -55514
rect 36400 -55514 36416 -55497
rect 36972 -55497 37174 -55480
rect 37232 -55480 38192 -55442
rect 37232 -55497 37434 -55480
rect 36972 -55514 36988 -55497
rect 36400 -55530 36988 -55514
rect 37418 -55514 37434 -55497
rect 37990 -55497 38192 -55480
rect 38250 -55480 39210 -55442
rect 38250 -55497 38452 -55480
rect 37990 -55514 38006 -55497
rect 37418 -55530 38006 -55514
rect 38436 -55514 38452 -55497
rect 39008 -55497 39210 -55480
rect 39268 -55480 40228 -55442
rect 39268 -55497 39470 -55480
rect 39008 -55514 39024 -55497
rect 38436 -55530 39024 -55514
rect 39454 -55514 39470 -55497
rect 40026 -55497 40228 -55480
rect 40286 -55480 41246 -55442
rect 40286 -55497 40488 -55480
rect 40026 -55514 40042 -55497
rect 39454 -55530 40042 -55514
rect 40472 -55514 40488 -55497
rect 41044 -55497 41246 -55480
rect 41304 -55480 42264 -55442
rect 41304 -55497 41506 -55480
rect 41044 -55514 41060 -55497
rect 40472 -55530 41060 -55514
rect 41490 -55514 41506 -55497
rect 42062 -55497 42264 -55480
rect 42322 -55480 43282 -55442
rect 42322 -55497 42524 -55480
rect 42062 -55514 42078 -55497
rect 41490 -55530 42078 -55514
rect 42508 -55514 42524 -55497
rect 43080 -55497 43282 -55480
rect 43340 -55480 44300 -55442
rect 43340 -55497 43542 -55480
rect 43080 -55514 43096 -55497
rect 42508 -55530 43096 -55514
rect 43526 -55514 43542 -55497
rect 44098 -55497 44300 -55480
rect 44358 -55480 45318 -55442
rect 44358 -55497 44560 -55480
rect 44098 -55514 44114 -55497
rect 43526 -55530 44114 -55514
rect 44544 -55514 44560 -55497
rect 45116 -55497 45318 -55480
rect 45376 -55480 46336 -55442
rect 45376 -55497 45578 -55480
rect 45116 -55514 45132 -55497
rect 44544 -55530 45132 -55514
rect 45562 -55514 45578 -55497
rect 46134 -55497 46336 -55480
rect 46394 -55480 47354 -55442
rect 46394 -55497 46596 -55480
rect 46134 -55514 46150 -55497
rect 45562 -55530 46150 -55514
rect 46580 -55514 46596 -55497
rect 47152 -55497 47354 -55480
rect 47412 -55480 48372 -55442
rect 47412 -55497 47614 -55480
rect 47152 -55514 47168 -55497
rect 46580 -55530 47168 -55514
rect 47598 -55514 47614 -55497
rect 48170 -55497 48372 -55480
rect 48170 -55514 48186 -55497
rect 47598 -55530 48186 -55514
rect 25162 -55576 26122 -55538
rect 28256 -56004 28844 -55988
rect 28256 -56021 28272 -56004
rect 28070 -56038 28272 -56021
rect 28828 -56021 28844 -56004
rect 29274 -56004 29862 -55988
rect 29274 -56021 29290 -56004
rect 28828 -56038 29030 -56021
rect 28070 -56076 29030 -56038
rect 29088 -56038 29290 -56021
rect 29846 -56021 29862 -56004
rect 30292 -56004 30880 -55988
rect 30292 -56021 30308 -56004
rect 29846 -56038 30048 -56021
rect 29088 -56076 30048 -56038
rect 30106 -56038 30308 -56021
rect 30864 -56021 30880 -56004
rect 31310 -56004 31898 -55988
rect 31310 -56021 31326 -56004
rect 30864 -56038 31066 -56021
rect 30106 -56076 31066 -56038
rect 31124 -56038 31326 -56021
rect 31882 -56021 31898 -56004
rect 32328 -56004 32916 -55988
rect 32328 -56021 32344 -56004
rect 31882 -56038 32084 -56021
rect 31124 -56076 32084 -56038
rect 32142 -56038 32344 -56021
rect 32900 -56021 32916 -56004
rect 33346 -56004 33934 -55988
rect 33346 -56021 33362 -56004
rect 32900 -56038 33102 -56021
rect 32142 -56076 33102 -56038
rect 33160 -56038 33362 -56021
rect 33918 -56021 33934 -56004
rect 34364 -56004 34952 -55988
rect 34364 -56021 34380 -56004
rect 33918 -56038 34120 -56021
rect 33160 -56076 34120 -56038
rect 34178 -56038 34380 -56021
rect 34936 -56021 34952 -56004
rect 35382 -56004 35970 -55988
rect 35382 -56021 35398 -56004
rect 34936 -56038 35138 -56021
rect 34178 -56076 35138 -56038
rect 35196 -56038 35398 -56021
rect 35954 -56021 35970 -56004
rect 36400 -56004 36988 -55988
rect 36400 -56021 36416 -56004
rect 35954 -56038 36156 -56021
rect 35196 -56076 36156 -56038
rect 36214 -56038 36416 -56021
rect 36972 -56021 36988 -56004
rect 37418 -56004 38006 -55988
rect 37418 -56021 37434 -56004
rect 36972 -56038 37174 -56021
rect 36214 -56076 37174 -56038
rect 37232 -56038 37434 -56021
rect 37990 -56021 38006 -56004
rect 38436 -56004 39024 -55988
rect 38436 -56021 38452 -56004
rect 37990 -56038 38192 -56021
rect 37232 -56076 38192 -56038
rect 38250 -56038 38452 -56021
rect 39008 -56021 39024 -56004
rect 39454 -56004 40042 -55988
rect 39454 -56021 39470 -56004
rect 39008 -56038 39210 -56021
rect 38250 -56076 39210 -56038
rect 39268 -56038 39470 -56021
rect 40026 -56021 40042 -56004
rect 40472 -56004 41060 -55988
rect 40472 -56021 40488 -56004
rect 40026 -56038 40228 -56021
rect 39268 -56076 40228 -56038
rect 40286 -56038 40488 -56021
rect 41044 -56021 41060 -56004
rect 41490 -56004 42078 -55988
rect 41490 -56021 41506 -56004
rect 41044 -56038 41246 -56021
rect 40286 -56076 41246 -56038
rect 41304 -56038 41506 -56021
rect 42062 -56021 42078 -56004
rect 42508 -56004 43096 -55988
rect 42508 -56021 42524 -56004
rect 42062 -56038 42264 -56021
rect 41304 -56076 42264 -56038
rect 42322 -56038 42524 -56021
rect 43080 -56021 43096 -56004
rect 43526 -56004 44114 -55988
rect 43526 -56021 43542 -56004
rect 43080 -56038 43282 -56021
rect 42322 -56076 43282 -56038
rect 43340 -56038 43542 -56021
rect 44098 -56021 44114 -56004
rect 44544 -56004 45132 -55988
rect 44544 -56021 44560 -56004
rect 44098 -56038 44300 -56021
rect 43340 -56076 44300 -56038
rect 44358 -56038 44560 -56021
rect 45116 -56021 45132 -56004
rect 45562 -56004 46150 -55988
rect 45562 -56021 45578 -56004
rect 45116 -56038 45318 -56021
rect 44358 -56076 45318 -56038
rect 45376 -56038 45578 -56021
rect 46134 -56021 46150 -56004
rect 46580 -56004 47168 -55988
rect 46580 -56021 46596 -56004
rect 46134 -56038 46336 -56021
rect 45376 -56076 46336 -56038
rect 46394 -56038 46596 -56021
rect 47152 -56021 47168 -56004
rect 47598 -56004 48186 -55988
rect 47598 -56021 47614 -56004
rect 47152 -56038 47354 -56021
rect 46394 -56076 47354 -56038
rect 47412 -56038 47614 -56021
rect 48170 -56021 48186 -56004
rect 48170 -56038 48372 -56021
rect 47412 -56076 48372 -56038
rect 14982 -56214 15942 -56176
rect 14982 -56231 15184 -56214
rect 15168 -56248 15184 -56231
rect 15740 -56231 15942 -56214
rect 16000 -56214 16960 -56176
rect 16000 -56231 16202 -56214
rect 15740 -56248 15756 -56231
rect 15168 -56264 15756 -56248
rect 16186 -56248 16202 -56231
rect 16758 -56231 16960 -56214
rect 17018 -56214 17978 -56176
rect 17018 -56231 17220 -56214
rect 16758 -56248 16774 -56231
rect 16186 -56264 16774 -56248
rect 17204 -56248 17220 -56231
rect 17776 -56231 17978 -56214
rect 18036 -56214 18996 -56176
rect 18036 -56231 18238 -56214
rect 17776 -56248 17792 -56231
rect 17204 -56264 17792 -56248
rect 18222 -56248 18238 -56231
rect 18794 -56231 18996 -56214
rect 19054 -56214 20014 -56176
rect 19054 -56231 19256 -56214
rect 18794 -56248 18810 -56231
rect 18222 -56264 18810 -56248
rect 19240 -56248 19256 -56231
rect 19812 -56231 20014 -56214
rect 20072 -56214 21032 -56176
rect 20072 -56231 20274 -56214
rect 19812 -56248 19828 -56231
rect 19240 -56264 19828 -56248
rect 20258 -56248 20274 -56231
rect 20830 -56231 21032 -56214
rect 21090 -56214 22050 -56176
rect 21090 -56231 21292 -56214
rect 20830 -56248 20846 -56231
rect 20258 -56264 20846 -56248
rect 21276 -56248 21292 -56231
rect 21848 -56231 22050 -56214
rect 22108 -56214 23068 -56176
rect 22108 -56231 22310 -56214
rect 21848 -56248 21864 -56231
rect 21276 -56264 21864 -56248
rect 22294 -56248 22310 -56231
rect 22866 -56231 23068 -56214
rect 23126 -56214 24086 -56176
rect 23126 -56231 23328 -56214
rect 22866 -56248 22882 -56231
rect 22294 -56264 22882 -56248
rect 23312 -56248 23328 -56231
rect 23884 -56231 24086 -56214
rect 24144 -56214 25104 -56176
rect 24144 -56231 24346 -56214
rect 23884 -56248 23900 -56231
rect 23312 -56264 23900 -56248
rect 24330 -56248 24346 -56231
rect 24902 -56231 25104 -56214
rect 25162 -56214 26122 -56176
rect 25162 -56231 25364 -56214
rect 24902 -56248 24918 -56231
rect 24330 -56264 24918 -56248
rect 25348 -56248 25364 -56231
rect 25920 -56231 26122 -56214
rect 25920 -56248 25936 -56231
rect 25348 -56264 25936 -56248
rect 28070 -56714 29030 -56676
rect 28070 -56731 28272 -56714
rect 28256 -56748 28272 -56731
rect 28828 -56731 29030 -56714
rect 29088 -56714 30048 -56676
rect 29088 -56731 29290 -56714
rect 28828 -56748 28844 -56731
rect 28256 -56764 28844 -56748
rect 29274 -56748 29290 -56731
rect 29846 -56731 30048 -56714
rect 30106 -56714 31066 -56676
rect 30106 -56731 30308 -56714
rect 29846 -56748 29862 -56731
rect 29274 -56764 29862 -56748
rect 30292 -56748 30308 -56731
rect 30864 -56731 31066 -56714
rect 31124 -56714 32084 -56676
rect 31124 -56731 31326 -56714
rect 30864 -56748 30880 -56731
rect 30292 -56764 30880 -56748
rect 31310 -56748 31326 -56731
rect 31882 -56731 32084 -56714
rect 32142 -56714 33102 -56676
rect 32142 -56731 32344 -56714
rect 31882 -56748 31898 -56731
rect 31310 -56764 31898 -56748
rect 32328 -56748 32344 -56731
rect 32900 -56731 33102 -56714
rect 33160 -56714 34120 -56676
rect 33160 -56731 33362 -56714
rect 32900 -56748 32916 -56731
rect 32328 -56764 32916 -56748
rect 33346 -56748 33362 -56731
rect 33918 -56731 34120 -56714
rect 34178 -56714 35138 -56676
rect 34178 -56731 34380 -56714
rect 33918 -56748 33934 -56731
rect 33346 -56764 33934 -56748
rect 34364 -56748 34380 -56731
rect 34936 -56731 35138 -56714
rect 35196 -56714 36156 -56676
rect 35196 -56731 35398 -56714
rect 34936 -56748 34952 -56731
rect 34364 -56764 34952 -56748
rect 35382 -56748 35398 -56731
rect 35954 -56731 36156 -56714
rect 36214 -56714 37174 -56676
rect 36214 -56731 36416 -56714
rect 35954 -56748 35970 -56731
rect 35382 -56764 35970 -56748
rect 36400 -56748 36416 -56731
rect 36972 -56731 37174 -56714
rect 37232 -56714 38192 -56676
rect 37232 -56731 37434 -56714
rect 36972 -56748 36988 -56731
rect 36400 -56764 36988 -56748
rect 37418 -56748 37434 -56731
rect 37990 -56731 38192 -56714
rect 38250 -56714 39210 -56676
rect 38250 -56731 38452 -56714
rect 37990 -56748 38006 -56731
rect 37418 -56764 38006 -56748
rect 38436 -56748 38452 -56731
rect 39008 -56731 39210 -56714
rect 39268 -56714 40228 -56676
rect 39268 -56731 39470 -56714
rect 39008 -56748 39024 -56731
rect 38436 -56764 39024 -56748
rect 39454 -56748 39470 -56731
rect 40026 -56731 40228 -56714
rect 40286 -56714 41246 -56676
rect 40286 -56731 40488 -56714
rect 40026 -56748 40042 -56731
rect 39454 -56764 40042 -56748
rect 40472 -56748 40488 -56731
rect 41044 -56731 41246 -56714
rect 41304 -56714 42264 -56676
rect 41304 -56731 41506 -56714
rect 41044 -56748 41060 -56731
rect 40472 -56764 41060 -56748
rect 41490 -56748 41506 -56731
rect 42062 -56731 42264 -56714
rect 42322 -56714 43282 -56676
rect 42322 -56731 42524 -56714
rect 42062 -56748 42078 -56731
rect 41490 -56764 42078 -56748
rect 42508 -56748 42524 -56731
rect 43080 -56731 43282 -56714
rect 43340 -56714 44300 -56676
rect 43340 -56731 43542 -56714
rect 43080 -56748 43096 -56731
rect 42508 -56764 43096 -56748
rect 43526 -56748 43542 -56731
rect 44098 -56731 44300 -56714
rect 44358 -56714 45318 -56676
rect 44358 -56731 44560 -56714
rect 44098 -56748 44114 -56731
rect 43526 -56764 44114 -56748
rect 44544 -56748 44560 -56731
rect 45116 -56731 45318 -56714
rect 45376 -56714 46336 -56676
rect 45376 -56731 45578 -56714
rect 45116 -56748 45132 -56731
rect 44544 -56764 45132 -56748
rect 45562 -56748 45578 -56731
rect 46134 -56731 46336 -56714
rect 46394 -56714 47354 -56676
rect 46394 -56731 46596 -56714
rect 46134 -56748 46150 -56731
rect 45562 -56764 46150 -56748
rect 46580 -56748 46596 -56731
rect 47152 -56731 47354 -56714
rect 47412 -56714 48372 -56676
rect 47412 -56731 47614 -56714
rect 47152 -56748 47168 -56731
rect 46580 -56764 47168 -56748
rect 47598 -56748 47614 -56731
rect 48170 -56731 48372 -56714
rect 48170 -56748 48186 -56731
rect 47598 -56764 48186 -56748
rect 15626 -57046 16214 -57030
rect 15626 -57063 15642 -57046
rect 15440 -57080 15642 -57063
rect 16198 -57063 16214 -57046
rect 16644 -57046 17232 -57030
rect 16644 -57063 16660 -57046
rect 16198 -57080 16400 -57063
rect 15440 -57118 16400 -57080
rect 16458 -57080 16660 -57063
rect 17216 -57063 17232 -57046
rect 17662 -57046 18250 -57030
rect 17662 -57063 17678 -57046
rect 17216 -57080 17418 -57063
rect 16458 -57118 17418 -57080
rect 17476 -57080 17678 -57063
rect 18234 -57063 18250 -57046
rect 18680 -57046 19268 -57030
rect 18680 -57063 18696 -57046
rect 18234 -57080 18436 -57063
rect 17476 -57118 18436 -57080
rect 18494 -57080 18696 -57063
rect 19252 -57063 19268 -57046
rect 19698 -57046 20286 -57030
rect 19698 -57063 19714 -57046
rect 19252 -57080 19454 -57063
rect 18494 -57118 19454 -57080
rect 19512 -57080 19714 -57063
rect 20270 -57063 20286 -57046
rect 20716 -57046 21304 -57030
rect 20716 -57063 20732 -57046
rect 20270 -57080 20472 -57063
rect 19512 -57118 20472 -57080
rect 20530 -57080 20732 -57063
rect 21288 -57063 21304 -57046
rect 21734 -57046 22322 -57030
rect 21734 -57063 21750 -57046
rect 21288 -57080 21490 -57063
rect 20530 -57118 21490 -57080
rect 21548 -57080 21750 -57063
rect 22306 -57063 22322 -57046
rect 22752 -57046 23340 -57030
rect 22752 -57063 22768 -57046
rect 22306 -57080 22508 -57063
rect 21548 -57118 22508 -57080
rect 22566 -57080 22768 -57063
rect 23324 -57063 23340 -57046
rect 23770 -57046 24358 -57030
rect 23770 -57063 23786 -57046
rect 23324 -57080 23526 -57063
rect 22566 -57118 23526 -57080
rect 23584 -57080 23786 -57063
rect 24342 -57063 24358 -57046
rect 24788 -57046 25376 -57030
rect 24788 -57063 24804 -57046
rect 24342 -57080 24544 -57063
rect 23584 -57118 24544 -57080
rect 24602 -57080 24804 -57063
rect 25360 -57063 25376 -57046
rect 25360 -57080 25562 -57063
rect 24602 -57118 25562 -57080
rect 28256 -57236 28844 -57220
rect 28256 -57253 28272 -57236
rect 28070 -57270 28272 -57253
rect 28828 -57253 28844 -57236
rect 29274 -57236 29862 -57220
rect 29274 -57253 29290 -57236
rect 28828 -57270 29030 -57253
rect 28070 -57308 29030 -57270
rect 29088 -57270 29290 -57253
rect 29846 -57253 29862 -57236
rect 30292 -57236 30880 -57220
rect 30292 -57253 30308 -57236
rect 29846 -57270 30048 -57253
rect 29088 -57308 30048 -57270
rect 30106 -57270 30308 -57253
rect 30864 -57253 30880 -57236
rect 31310 -57236 31898 -57220
rect 31310 -57253 31326 -57236
rect 30864 -57270 31066 -57253
rect 30106 -57308 31066 -57270
rect 31124 -57270 31326 -57253
rect 31882 -57253 31898 -57236
rect 32328 -57236 32916 -57220
rect 32328 -57253 32344 -57236
rect 31882 -57270 32084 -57253
rect 31124 -57308 32084 -57270
rect 32142 -57270 32344 -57253
rect 32900 -57253 32916 -57236
rect 33346 -57236 33934 -57220
rect 33346 -57253 33362 -57236
rect 32900 -57270 33102 -57253
rect 32142 -57308 33102 -57270
rect 33160 -57270 33362 -57253
rect 33918 -57253 33934 -57236
rect 34364 -57236 34952 -57220
rect 34364 -57253 34380 -57236
rect 33918 -57270 34120 -57253
rect 33160 -57308 34120 -57270
rect 34178 -57270 34380 -57253
rect 34936 -57253 34952 -57236
rect 35382 -57236 35970 -57220
rect 35382 -57253 35398 -57236
rect 34936 -57270 35138 -57253
rect 34178 -57308 35138 -57270
rect 35196 -57270 35398 -57253
rect 35954 -57253 35970 -57236
rect 36400 -57236 36988 -57220
rect 36400 -57253 36416 -57236
rect 35954 -57270 36156 -57253
rect 35196 -57308 36156 -57270
rect 36214 -57270 36416 -57253
rect 36972 -57253 36988 -57236
rect 37418 -57236 38006 -57220
rect 37418 -57253 37434 -57236
rect 36972 -57270 37174 -57253
rect 36214 -57308 37174 -57270
rect 37232 -57270 37434 -57253
rect 37990 -57253 38006 -57236
rect 38436 -57236 39024 -57220
rect 38436 -57253 38452 -57236
rect 37990 -57270 38192 -57253
rect 37232 -57308 38192 -57270
rect 38250 -57270 38452 -57253
rect 39008 -57253 39024 -57236
rect 39454 -57236 40042 -57220
rect 39454 -57253 39470 -57236
rect 39008 -57270 39210 -57253
rect 38250 -57308 39210 -57270
rect 39268 -57270 39470 -57253
rect 40026 -57253 40042 -57236
rect 40472 -57236 41060 -57220
rect 40472 -57253 40488 -57236
rect 40026 -57270 40228 -57253
rect 39268 -57308 40228 -57270
rect 40286 -57270 40488 -57253
rect 41044 -57253 41060 -57236
rect 41490 -57236 42078 -57220
rect 41490 -57253 41506 -57236
rect 41044 -57270 41246 -57253
rect 40286 -57308 41246 -57270
rect 41304 -57270 41506 -57253
rect 42062 -57253 42078 -57236
rect 42508 -57236 43096 -57220
rect 42508 -57253 42524 -57236
rect 42062 -57270 42264 -57253
rect 41304 -57308 42264 -57270
rect 42322 -57270 42524 -57253
rect 43080 -57253 43096 -57236
rect 43526 -57236 44114 -57220
rect 43526 -57253 43542 -57236
rect 43080 -57270 43282 -57253
rect 42322 -57308 43282 -57270
rect 43340 -57270 43542 -57253
rect 44098 -57253 44114 -57236
rect 44544 -57236 45132 -57220
rect 44544 -57253 44560 -57236
rect 44098 -57270 44300 -57253
rect 43340 -57308 44300 -57270
rect 44358 -57270 44560 -57253
rect 45116 -57253 45132 -57236
rect 45562 -57236 46150 -57220
rect 45562 -57253 45578 -57236
rect 45116 -57270 45318 -57253
rect 44358 -57308 45318 -57270
rect 45376 -57270 45578 -57253
rect 46134 -57253 46150 -57236
rect 46580 -57236 47168 -57220
rect 46580 -57253 46596 -57236
rect 46134 -57270 46336 -57253
rect 45376 -57308 46336 -57270
rect 46394 -57270 46596 -57253
rect 47152 -57253 47168 -57236
rect 47598 -57236 48186 -57220
rect 47598 -57253 47614 -57236
rect 47152 -57270 47354 -57253
rect 46394 -57308 47354 -57270
rect 47412 -57270 47614 -57253
rect 48170 -57253 48186 -57236
rect 48170 -57270 48372 -57253
rect 47412 -57308 48372 -57270
rect 15440 -57756 16400 -57718
rect 15440 -57773 15642 -57756
rect 15626 -57790 15642 -57773
rect 16198 -57773 16400 -57756
rect 16458 -57756 17418 -57718
rect 16458 -57773 16660 -57756
rect 16198 -57790 16214 -57773
rect 15626 -57806 16214 -57790
rect 16644 -57790 16660 -57773
rect 17216 -57773 17418 -57756
rect 17476 -57756 18436 -57718
rect 17476 -57773 17678 -57756
rect 17216 -57790 17232 -57773
rect 16644 -57806 17232 -57790
rect 17662 -57790 17678 -57773
rect 18234 -57773 18436 -57756
rect 18494 -57756 19454 -57718
rect 18494 -57773 18696 -57756
rect 18234 -57790 18250 -57773
rect 17662 -57806 18250 -57790
rect 18680 -57790 18696 -57773
rect 19252 -57773 19454 -57756
rect 19512 -57756 20472 -57718
rect 19512 -57773 19714 -57756
rect 19252 -57790 19268 -57773
rect 18680 -57806 19268 -57790
rect 19698 -57790 19714 -57773
rect 20270 -57773 20472 -57756
rect 20530 -57756 21490 -57718
rect 20530 -57773 20732 -57756
rect 20270 -57790 20286 -57773
rect 19698 -57806 20286 -57790
rect 20716 -57790 20732 -57773
rect 21288 -57773 21490 -57756
rect 21548 -57756 22508 -57718
rect 21548 -57773 21750 -57756
rect 21288 -57790 21304 -57773
rect 20716 -57806 21304 -57790
rect 21734 -57790 21750 -57773
rect 22306 -57773 22508 -57756
rect 22566 -57756 23526 -57718
rect 22566 -57773 22768 -57756
rect 22306 -57790 22322 -57773
rect 21734 -57806 22322 -57790
rect 22752 -57790 22768 -57773
rect 23324 -57773 23526 -57756
rect 23584 -57756 24544 -57718
rect 23584 -57773 23786 -57756
rect 23324 -57790 23340 -57773
rect 22752 -57806 23340 -57790
rect 23770 -57790 23786 -57773
rect 24342 -57773 24544 -57756
rect 24602 -57756 25562 -57718
rect 24602 -57773 24804 -57756
rect 24342 -57790 24358 -57773
rect 23770 -57806 24358 -57790
rect 24788 -57790 24804 -57773
rect 25360 -57773 25562 -57756
rect 25360 -57790 25376 -57773
rect 24788 -57806 25376 -57790
rect 28070 -57946 29030 -57908
rect 28070 -57963 28272 -57946
rect 28256 -57980 28272 -57963
rect 28828 -57963 29030 -57946
rect 29088 -57946 30048 -57908
rect 29088 -57963 29290 -57946
rect 28828 -57980 28844 -57963
rect 28256 -57996 28844 -57980
rect 29274 -57980 29290 -57963
rect 29846 -57963 30048 -57946
rect 30106 -57946 31066 -57908
rect 30106 -57963 30308 -57946
rect 29846 -57980 29862 -57963
rect 29274 -57996 29862 -57980
rect 30292 -57980 30308 -57963
rect 30864 -57963 31066 -57946
rect 31124 -57946 32084 -57908
rect 31124 -57963 31326 -57946
rect 30864 -57980 30880 -57963
rect 30292 -57996 30880 -57980
rect 31310 -57980 31326 -57963
rect 31882 -57963 32084 -57946
rect 32142 -57946 33102 -57908
rect 32142 -57963 32344 -57946
rect 31882 -57980 31898 -57963
rect 31310 -57996 31898 -57980
rect 32328 -57980 32344 -57963
rect 32900 -57963 33102 -57946
rect 33160 -57946 34120 -57908
rect 33160 -57963 33362 -57946
rect 32900 -57980 32916 -57963
rect 32328 -57996 32916 -57980
rect 33346 -57980 33362 -57963
rect 33918 -57963 34120 -57946
rect 34178 -57946 35138 -57908
rect 34178 -57963 34380 -57946
rect 33918 -57980 33934 -57963
rect 33346 -57996 33934 -57980
rect 34364 -57980 34380 -57963
rect 34936 -57963 35138 -57946
rect 35196 -57946 36156 -57908
rect 35196 -57963 35398 -57946
rect 34936 -57980 34952 -57963
rect 34364 -57996 34952 -57980
rect 35382 -57980 35398 -57963
rect 35954 -57963 36156 -57946
rect 36214 -57946 37174 -57908
rect 36214 -57963 36416 -57946
rect 35954 -57980 35970 -57963
rect 35382 -57996 35970 -57980
rect 36400 -57980 36416 -57963
rect 36972 -57963 37174 -57946
rect 37232 -57946 38192 -57908
rect 37232 -57963 37434 -57946
rect 36972 -57980 36988 -57963
rect 36400 -57996 36988 -57980
rect 37418 -57980 37434 -57963
rect 37990 -57963 38192 -57946
rect 38250 -57946 39210 -57908
rect 38250 -57963 38452 -57946
rect 37990 -57980 38006 -57963
rect 37418 -57996 38006 -57980
rect 38436 -57980 38452 -57963
rect 39008 -57963 39210 -57946
rect 39268 -57946 40228 -57908
rect 39268 -57963 39470 -57946
rect 39008 -57980 39024 -57963
rect 38436 -57996 39024 -57980
rect 39454 -57980 39470 -57963
rect 40026 -57963 40228 -57946
rect 40286 -57946 41246 -57908
rect 40286 -57963 40488 -57946
rect 40026 -57980 40042 -57963
rect 39454 -57996 40042 -57980
rect 40472 -57980 40488 -57963
rect 41044 -57963 41246 -57946
rect 41304 -57946 42264 -57908
rect 41304 -57963 41506 -57946
rect 41044 -57980 41060 -57963
rect 40472 -57996 41060 -57980
rect 41490 -57980 41506 -57963
rect 42062 -57963 42264 -57946
rect 42322 -57946 43282 -57908
rect 42322 -57963 42524 -57946
rect 42062 -57980 42078 -57963
rect 41490 -57996 42078 -57980
rect 42508 -57980 42524 -57963
rect 43080 -57963 43282 -57946
rect 43340 -57946 44300 -57908
rect 43340 -57963 43542 -57946
rect 43080 -57980 43096 -57963
rect 42508 -57996 43096 -57980
rect 43526 -57980 43542 -57963
rect 44098 -57963 44300 -57946
rect 44358 -57946 45318 -57908
rect 44358 -57963 44560 -57946
rect 44098 -57980 44114 -57963
rect 43526 -57996 44114 -57980
rect 44544 -57980 44560 -57963
rect 45116 -57963 45318 -57946
rect 45376 -57946 46336 -57908
rect 45376 -57963 45578 -57946
rect 45116 -57980 45132 -57963
rect 44544 -57996 45132 -57980
rect 45562 -57980 45578 -57963
rect 46134 -57963 46336 -57946
rect 46394 -57946 47354 -57908
rect 46394 -57963 46596 -57946
rect 46134 -57980 46150 -57963
rect 45562 -57996 46150 -57980
rect 46580 -57980 46596 -57963
rect 47152 -57963 47354 -57946
rect 47412 -57946 48372 -57908
rect 47412 -57963 47614 -57946
rect 47152 -57980 47168 -57963
rect 46580 -57996 47168 -57980
rect 47598 -57980 47614 -57963
rect 48170 -57963 48372 -57946
rect 48170 -57980 48186 -57963
rect 47598 -57996 48186 -57980
rect 57963 -42630 58029 -42614
rect 57963 -42664 57979 -42630
rect 58013 -42664 58029 -42630
rect 57963 -42680 58029 -42664
rect 57966 -42702 58026 -42680
rect 57966 -42928 58026 -42902
rect -27952 -67329 -27922 -67303
rect -27257 -65544 -27125 -65528
rect -27257 -65561 -27241 -65544
rect -27291 -65578 -27241 -65561
rect -27141 -65561 -27125 -65544
rect -26999 -65544 -26867 -65528
rect -26999 -65561 -26983 -65544
rect -27141 -65578 -27091 -65561
rect -27291 -65625 -27091 -65578
rect -27033 -65578 -26983 -65561
rect -26883 -65561 -26867 -65544
rect -26741 -65544 -26609 -65528
rect -26741 -65561 -26725 -65544
rect -26883 -65578 -26833 -65561
rect -27033 -65625 -26833 -65578
rect -26775 -65578 -26725 -65561
rect -26625 -65561 -26609 -65544
rect -26483 -65544 -26351 -65528
rect -26483 -65561 -26467 -65544
rect -26625 -65578 -26575 -65561
rect -26775 -65625 -26575 -65578
rect -26517 -65578 -26467 -65561
rect -26367 -65561 -26351 -65544
rect -26225 -65544 -26093 -65528
rect -26225 -65561 -26209 -65544
rect -26367 -65578 -26317 -65561
rect -26517 -65625 -26317 -65578
rect -26259 -65578 -26209 -65561
rect -26109 -65561 -26093 -65544
rect -25967 -65544 -25835 -65528
rect -25967 -65561 -25951 -65544
rect -26109 -65578 -26059 -65561
rect -26259 -65625 -26059 -65578
rect -26001 -65578 -25951 -65561
rect -25851 -65561 -25835 -65544
rect -25851 -65578 -25801 -65561
rect -26001 -65625 -25801 -65578
rect -27291 -66072 -27091 -66025
rect -27291 -66089 -27241 -66072
rect -27257 -66106 -27241 -66089
rect -27141 -66089 -27091 -66072
rect -27033 -66072 -26833 -66025
rect -27033 -66089 -26983 -66072
rect -27141 -66106 -27125 -66089
rect -27257 -66122 -27125 -66106
rect -26999 -66106 -26983 -66089
rect -26883 -66089 -26833 -66072
rect -26775 -66072 -26575 -66025
rect -26775 -66089 -26725 -66072
rect -26883 -66106 -26867 -66089
rect -26999 -66122 -26867 -66106
rect -26741 -66106 -26725 -66089
rect -26625 -66089 -26575 -66072
rect -26517 -66072 -26317 -66025
rect -26517 -66089 -26467 -66072
rect -26625 -66106 -26609 -66089
rect -26741 -66122 -26609 -66106
rect -26483 -66106 -26467 -66089
rect -26367 -66089 -26317 -66072
rect -26259 -66072 -26059 -66025
rect -26259 -66089 -26209 -66072
rect -26367 -66106 -26351 -66089
rect -26483 -66122 -26351 -66106
rect -26225 -66106 -26209 -66089
rect -26109 -66089 -26059 -66072
rect -26001 -66072 -25801 -66025
rect -26001 -66089 -25951 -66072
rect -26109 -66106 -26093 -66089
rect -26225 -66122 -26093 -66106
rect -25967 -66106 -25951 -66089
rect -25851 -66089 -25801 -66072
rect -25851 -66106 -25835 -66089
rect -25967 -66122 -25835 -66106
rect -27257 -66404 -27125 -66388
rect -27257 -66421 -27241 -66404
rect -27291 -66438 -27241 -66421
rect -27141 -66421 -27125 -66404
rect -26999 -66404 -26867 -66388
rect -26999 -66421 -26983 -66404
rect -27141 -66438 -27091 -66421
rect -27291 -66485 -27091 -66438
rect -27033 -66438 -26983 -66421
rect -26883 -66421 -26867 -66404
rect -26741 -66404 -26609 -66388
rect -26741 -66421 -26725 -66404
rect -26883 -66438 -26833 -66421
rect -27033 -66485 -26833 -66438
rect -26775 -66438 -26725 -66421
rect -26625 -66421 -26609 -66404
rect -26483 -66404 -26351 -66388
rect -26483 -66421 -26467 -66404
rect -26625 -66438 -26575 -66421
rect -26775 -66485 -26575 -66438
rect -26517 -66438 -26467 -66421
rect -26367 -66421 -26351 -66404
rect -26225 -66404 -26093 -66388
rect -26225 -66421 -26209 -66404
rect -26367 -66438 -26317 -66421
rect -26517 -66485 -26317 -66438
rect -26259 -66438 -26209 -66421
rect -26109 -66421 -26093 -66404
rect -25967 -66404 -25835 -66388
rect -25967 -66421 -25951 -66404
rect -26109 -66438 -26059 -66421
rect -26259 -66485 -26059 -66438
rect -26001 -66438 -25951 -66421
rect -25851 -66421 -25835 -66404
rect -25851 -66438 -25801 -66421
rect -26001 -66485 -25801 -66438
rect -27291 -66932 -27091 -66885
rect -27291 -66949 -27241 -66932
rect -27257 -66966 -27241 -66949
rect -27141 -66949 -27091 -66932
rect -27033 -66932 -26833 -66885
rect -27033 -66949 -26983 -66932
rect -27141 -66966 -27125 -66949
rect -27257 -66982 -27125 -66966
rect -26999 -66966 -26983 -66949
rect -26883 -66949 -26833 -66932
rect -26775 -66932 -26575 -66885
rect -26775 -66949 -26725 -66932
rect -26883 -66966 -26867 -66949
rect -26999 -66982 -26867 -66966
rect -26741 -66966 -26725 -66949
rect -26625 -66949 -26575 -66932
rect -26517 -66932 -26317 -66885
rect -26517 -66949 -26467 -66932
rect -26625 -66966 -26609 -66949
rect -26741 -66982 -26609 -66966
rect -26483 -66966 -26467 -66949
rect -26367 -66949 -26317 -66932
rect -26259 -66932 -26059 -66885
rect -26259 -66949 -26209 -66932
rect -26367 -66966 -26351 -66949
rect -26483 -66982 -26351 -66966
rect -26225 -66966 -26209 -66949
rect -26109 -66949 -26059 -66932
rect -26001 -66932 -25801 -66885
rect -26001 -66949 -25951 -66932
rect -26109 -66966 -26093 -66949
rect -26225 -66982 -26093 -66966
rect -25967 -66966 -25951 -66949
rect -25851 -66949 -25801 -66932
rect -25851 -66966 -25835 -66949
rect -25967 -66982 -25835 -66966
rect -23952 -67329 -23922 -67303
rect -27952 -67561 -27922 -67529
rect -23257 -65544 -23125 -65528
rect -23257 -65561 -23241 -65544
rect -23291 -65578 -23241 -65561
rect -23141 -65561 -23125 -65544
rect -22999 -65544 -22867 -65528
rect -22999 -65561 -22983 -65544
rect -23141 -65578 -23091 -65561
rect -23291 -65625 -23091 -65578
rect -23033 -65578 -22983 -65561
rect -22883 -65561 -22867 -65544
rect -22741 -65544 -22609 -65528
rect -22741 -65561 -22725 -65544
rect -22883 -65578 -22833 -65561
rect -23033 -65625 -22833 -65578
rect -22775 -65578 -22725 -65561
rect -22625 -65561 -22609 -65544
rect -22483 -65544 -22351 -65528
rect -22483 -65561 -22467 -65544
rect -22625 -65578 -22575 -65561
rect -22775 -65625 -22575 -65578
rect -22517 -65578 -22467 -65561
rect -22367 -65561 -22351 -65544
rect -22225 -65544 -22093 -65528
rect -22225 -65561 -22209 -65544
rect -22367 -65578 -22317 -65561
rect -22517 -65625 -22317 -65578
rect -22259 -65578 -22209 -65561
rect -22109 -65561 -22093 -65544
rect -21967 -65544 -21835 -65528
rect -21967 -65561 -21951 -65544
rect -22109 -65578 -22059 -65561
rect -22259 -65625 -22059 -65578
rect -22001 -65578 -21951 -65561
rect -21851 -65561 -21835 -65544
rect -21851 -65578 -21801 -65561
rect -22001 -65625 -21801 -65578
rect -23291 -66072 -23091 -66025
rect -23291 -66089 -23241 -66072
rect -23257 -66106 -23241 -66089
rect -23141 -66089 -23091 -66072
rect -23033 -66072 -22833 -66025
rect -23033 -66089 -22983 -66072
rect -23141 -66106 -23125 -66089
rect -23257 -66122 -23125 -66106
rect -22999 -66106 -22983 -66089
rect -22883 -66089 -22833 -66072
rect -22775 -66072 -22575 -66025
rect -22775 -66089 -22725 -66072
rect -22883 -66106 -22867 -66089
rect -22999 -66122 -22867 -66106
rect -22741 -66106 -22725 -66089
rect -22625 -66089 -22575 -66072
rect -22517 -66072 -22317 -66025
rect -22517 -66089 -22467 -66072
rect -22625 -66106 -22609 -66089
rect -22741 -66122 -22609 -66106
rect -22483 -66106 -22467 -66089
rect -22367 -66089 -22317 -66072
rect -22259 -66072 -22059 -66025
rect -22259 -66089 -22209 -66072
rect -22367 -66106 -22351 -66089
rect -22483 -66122 -22351 -66106
rect -22225 -66106 -22209 -66089
rect -22109 -66089 -22059 -66072
rect -22001 -66072 -21801 -66025
rect -22001 -66089 -21951 -66072
rect -22109 -66106 -22093 -66089
rect -22225 -66122 -22093 -66106
rect -21967 -66106 -21951 -66089
rect -21851 -66089 -21801 -66072
rect -21851 -66106 -21835 -66089
rect -21967 -66122 -21835 -66106
rect -23257 -66404 -23125 -66388
rect -23257 -66421 -23241 -66404
rect -23291 -66438 -23241 -66421
rect -23141 -66421 -23125 -66404
rect -22999 -66404 -22867 -66388
rect -22999 -66421 -22983 -66404
rect -23141 -66438 -23091 -66421
rect -23291 -66485 -23091 -66438
rect -23033 -66438 -22983 -66421
rect -22883 -66421 -22867 -66404
rect -22741 -66404 -22609 -66388
rect -22741 -66421 -22725 -66404
rect -22883 -66438 -22833 -66421
rect -23033 -66485 -22833 -66438
rect -22775 -66438 -22725 -66421
rect -22625 -66421 -22609 -66404
rect -22483 -66404 -22351 -66388
rect -22483 -66421 -22467 -66404
rect -22625 -66438 -22575 -66421
rect -22775 -66485 -22575 -66438
rect -22517 -66438 -22467 -66421
rect -22367 -66421 -22351 -66404
rect -22225 -66404 -22093 -66388
rect -22225 -66421 -22209 -66404
rect -22367 -66438 -22317 -66421
rect -22517 -66485 -22317 -66438
rect -22259 -66438 -22209 -66421
rect -22109 -66421 -22093 -66404
rect -21967 -66404 -21835 -66388
rect -21967 -66421 -21951 -66404
rect -22109 -66438 -22059 -66421
rect -22259 -66485 -22059 -66438
rect -22001 -66438 -21951 -66421
rect -21851 -66421 -21835 -66404
rect -21851 -66438 -21801 -66421
rect -22001 -66485 -21801 -66438
rect -23291 -66932 -23091 -66885
rect -23291 -66949 -23241 -66932
rect -23257 -66966 -23241 -66949
rect -23141 -66949 -23091 -66932
rect -23033 -66932 -22833 -66885
rect -23033 -66949 -22983 -66932
rect -23141 -66966 -23125 -66949
rect -23257 -66982 -23125 -66966
rect -22999 -66966 -22983 -66949
rect -22883 -66949 -22833 -66932
rect -22775 -66932 -22575 -66885
rect -22775 -66949 -22725 -66932
rect -22883 -66966 -22867 -66949
rect -22999 -66982 -22867 -66966
rect -22741 -66966 -22725 -66949
rect -22625 -66949 -22575 -66932
rect -22517 -66932 -22317 -66885
rect -22517 -66949 -22467 -66932
rect -22625 -66966 -22609 -66949
rect -22741 -66982 -22609 -66966
rect -22483 -66966 -22467 -66949
rect -22367 -66949 -22317 -66932
rect -22259 -66932 -22059 -66885
rect -22259 -66949 -22209 -66932
rect -22367 -66966 -22351 -66949
rect -22483 -66982 -22351 -66966
rect -22225 -66966 -22209 -66949
rect -22109 -66949 -22059 -66932
rect -22001 -66932 -21801 -66885
rect -22001 -66949 -21951 -66932
rect -22109 -66966 -22093 -66949
rect -22225 -66982 -22093 -66966
rect -21967 -66966 -21951 -66949
rect -21851 -66949 -21801 -66932
rect -21851 -66966 -21835 -66949
rect -21967 -66982 -21835 -66966
rect -19952 -67329 -19922 -67303
rect -23952 -67561 -23922 -67529
rect -19257 -65544 -19125 -65528
rect -19257 -65561 -19241 -65544
rect -19291 -65578 -19241 -65561
rect -19141 -65561 -19125 -65544
rect -18999 -65544 -18867 -65528
rect -18999 -65561 -18983 -65544
rect -19141 -65578 -19091 -65561
rect -19291 -65625 -19091 -65578
rect -19033 -65578 -18983 -65561
rect -18883 -65561 -18867 -65544
rect -18741 -65544 -18609 -65528
rect -18741 -65561 -18725 -65544
rect -18883 -65578 -18833 -65561
rect -19033 -65625 -18833 -65578
rect -18775 -65578 -18725 -65561
rect -18625 -65561 -18609 -65544
rect -18483 -65544 -18351 -65528
rect -18483 -65561 -18467 -65544
rect -18625 -65578 -18575 -65561
rect -18775 -65625 -18575 -65578
rect -18517 -65578 -18467 -65561
rect -18367 -65561 -18351 -65544
rect -18225 -65544 -18093 -65528
rect -18225 -65561 -18209 -65544
rect -18367 -65578 -18317 -65561
rect -18517 -65625 -18317 -65578
rect -18259 -65578 -18209 -65561
rect -18109 -65561 -18093 -65544
rect -17967 -65544 -17835 -65528
rect -17967 -65561 -17951 -65544
rect -18109 -65578 -18059 -65561
rect -18259 -65625 -18059 -65578
rect -18001 -65578 -17951 -65561
rect -17851 -65561 -17835 -65544
rect -17851 -65578 -17801 -65561
rect -18001 -65625 -17801 -65578
rect -19291 -66072 -19091 -66025
rect -19291 -66089 -19241 -66072
rect -19257 -66106 -19241 -66089
rect -19141 -66089 -19091 -66072
rect -19033 -66072 -18833 -66025
rect -19033 -66089 -18983 -66072
rect -19141 -66106 -19125 -66089
rect -19257 -66122 -19125 -66106
rect -18999 -66106 -18983 -66089
rect -18883 -66089 -18833 -66072
rect -18775 -66072 -18575 -66025
rect -18775 -66089 -18725 -66072
rect -18883 -66106 -18867 -66089
rect -18999 -66122 -18867 -66106
rect -18741 -66106 -18725 -66089
rect -18625 -66089 -18575 -66072
rect -18517 -66072 -18317 -66025
rect -18517 -66089 -18467 -66072
rect -18625 -66106 -18609 -66089
rect -18741 -66122 -18609 -66106
rect -18483 -66106 -18467 -66089
rect -18367 -66089 -18317 -66072
rect -18259 -66072 -18059 -66025
rect -18259 -66089 -18209 -66072
rect -18367 -66106 -18351 -66089
rect -18483 -66122 -18351 -66106
rect -18225 -66106 -18209 -66089
rect -18109 -66089 -18059 -66072
rect -18001 -66072 -17801 -66025
rect -18001 -66089 -17951 -66072
rect -18109 -66106 -18093 -66089
rect -18225 -66122 -18093 -66106
rect -17967 -66106 -17951 -66089
rect -17851 -66089 -17801 -66072
rect -17851 -66106 -17835 -66089
rect -17967 -66122 -17835 -66106
rect -19257 -66404 -19125 -66388
rect -19257 -66421 -19241 -66404
rect -19291 -66438 -19241 -66421
rect -19141 -66421 -19125 -66404
rect -18999 -66404 -18867 -66388
rect -18999 -66421 -18983 -66404
rect -19141 -66438 -19091 -66421
rect -19291 -66485 -19091 -66438
rect -19033 -66438 -18983 -66421
rect -18883 -66421 -18867 -66404
rect -18741 -66404 -18609 -66388
rect -18741 -66421 -18725 -66404
rect -18883 -66438 -18833 -66421
rect -19033 -66485 -18833 -66438
rect -18775 -66438 -18725 -66421
rect -18625 -66421 -18609 -66404
rect -18483 -66404 -18351 -66388
rect -18483 -66421 -18467 -66404
rect -18625 -66438 -18575 -66421
rect -18775 -66485 -18575 -66438
rect -18517 -66438 -18467 -66421
rect -18367 -66421 -18351 -66404
rect -18225 -66404 -18093 -66388
rect -18225 -66421 -18209 -66404
rect -18367 -66438 -18317 -66421
rect -18517 -66485 -18317 -66438
rect -18259 -66438 -18209 -66421
rect -18109 -66421 -18093 -66404
rect -17967 -66404 -17835 -66388
rect -17967 -66421 -17951 -66404
rect -18109 -66438 -18059 -66421
rect -18259 -66485 -18059 -66438
rect -18001 -66438 -17951 -66421
rect -17851 -66421 -17835 -66404
rect -17851 -66438 -17801 -66421
rect -18001 -66485 -17801 -66438
rect -19291 -66932 -19091 -66885
rect -19291 -66949 -19241 -66932
rect -19257 -66966 -19241 -66949
rect -19141 -66949 -19091 -66932
rect -19033 -66932 -18833 -66885
rect -19033 -66949 -18983 -66932
rect -19141 -66966 -19125 -66949
rect -19257 -66982 -19125 -66966
rect -18999 -66966 -18983 -66949
rect -18883 -66949 -18833 -66932
rect -18775 -66932 -18575 -66885
rect -18775 -66949 -18725 -66932
rect -18883 -66966 -18867 -66949
rect -18999 -66982 -18867 -66966
rect -18741 -66966 -18725 -66949
rect -18625 -66949 -18575 -66932
rect -18517 -66932 -18317 -66885
rect -18517 -66949 -18467 -66932
rect -18625 -66966 -18609 -66949
rect -18741 -66982 -18609 -66966
rect -18483 -66966 -18467 -66949
rect -18367 -66949 -18317 -66932
rect -18259 -66932 -18059 -66885
rect -18259 -66949 -18209 -66932
rect -18367 -66966 -18351 -66949
rect -18483 -66982 -18351 -66966
rect -18225 -66966 -18209 -66949
rect -18109 -66949 -18059 -66932
rect -18001 -66932 -17801 -66885
rect -18001 -66949 -17951 -66932
rect -18109 -66966 -18093 -66949
rect -18225 -66982 -18093 -66966
rect -17967 -66966 -17951 -66949
rect -17851 -66949 -17801 -66932
rect -17851 -66966 -17835 -66949
rect -17967 -66982 -17835 -66966
rect -15952 -67329 -15922 -67303
rect -19952 -67561 -19922 -67529
rect -15257 -65544 -15125 -65528
rect -15257 -65561 -15241 -65544
rect -15291 -65578 -15241 -65561
rect -15141 -65561 -15125 -65544
rect -14999 -65544 -14867 -65528
rect -14999 -65561 -14983 -65544
rect -15141 -65578 -15091 -65561
rect -15291 -65625 -15091 -65578
rect -15033 -65578 -14983 -65561
rect -14883 -65561 -14867 -65544
rect -14741 -65544 -14609 -65528
rect -14741 -65561 -14725 -65544
rect -14883 -65578 -14833 -65561
rect -15033 -65625 -14833 -65578
rect -14775 -65578 -14725 -65561
rect -14625 -65561 -14609 -65544
rect -14483 -65544 -14351 -65528
rect -14483 -65561 -14467 -65544
rect -14625 -65578 -14575 -65561
rect -14775 -65625 -14575 -65578
rect -14517 -65578 -14467 -65561
rect -14367 -65561 -14351 -65544
rect -14225 -65544 -14093 -65528
rect -14225 -65561 -14209 -65544
rect -14367 -65578 -14317 -65561
rect -14517 -65625 -14317 -65578
rect -14259 -65578 -14209 -65561
rect -14109 -65561 -14093 -65544
rect -13967 -65544 -13835 -65528
rect -13967 -65561 -13951 -65544
rect -14109 -65578 -14059 -65561
rect -14259 -65625 -14059 -65578
rect -14001 -65578 -13951 -65561
rect -13851 -65561 -13835 -65544
rect -13851 -65578 -13801 -65561
rect -14001 -65625 -13801 -65578
rect -15291 -66072 -15091 -66025
rect -15291 -66089 -15241 -66072
rect -15257 -66106 -15241 -66089
rect -15141 -66089 -15091 -66072
rect -15033 -66072 -14833 -66025
rect -15033 -66089 -14983 -66072
rect -15141 -66106 -15125 -66089
rect -15257 -66122 -15125 -66106
rect -14999 -66106 -14983 -66089
rect -14883 -66089 -14833 -66072
rect -14775 -66072 -14575 -66025
rect -14775 -66089 -14725 -66072
rect -14883 -66106 -14867 -66089
rect -14999 -66122 -14867 -66106
rect -14741 -66106 -14725 -66089
rect -14625 -66089 -14575 -66072
rect -14517 -66072 -14317 -66025
rect -14517 -66089 -14467 -66072
rect -14625 -66106 -14609 -66089
rect -14741 -66122 -14609 -66106
rect -14483 -66106 -14467 -66089
rect -14367 -66089 -14317 -66072
rect -14259 -66072 -14059 -66025
rect -14259 -66089 -14209 -66072
rect -14367 -66106 -14351 -66089
rect -14483 -66122 -14351 -66106
rect -14225 -66106 -14209 -66089
rect -14109 -66089 -14059 -66072
rect -14001 -66072 -13801 -66025
rect -14001 -66089 -13951 -66072
rect -14109 -66106 -14093 -66089
rect -14225 -66122 -14093 -66106
rect -13967 -66106 -13951 -66089
rect -13851 -66089 -13801 -66072
rect -13851 -66106 -13835 -66089
rect -13967 -66122 -13835 -66106
rect -15257 -66404 -15125 -66388
rect -15257 -66421 -15241 -66404
rect -15291 -66438 -15241 -66421
rect -15141 -66421 -15125 -66404
rect -14999 -66404 -14867 -66388
rect -14999 -66421 -14983 -66404
rect -15141 -66438 -15091 -66421
rect -15291 -66485 -15091 -66438
rect -15033 -66438 -14983 -66421
rect -14883 -66421 -14867 -66404
rect -14741 -66404 -14609 -66388
rect -14741 -66421 -14725 -66404
rect -14883 -66438 -14833 -66421
rect -15033 -66485 -14833 -66438
rect -14775 -66438 -14725 -66421
rect -14625 -66421 -14609 -66404
rect -14483 -66404 -14351 -66388
rect -14483 -66421 -14467 -66404
rect -14625 -66438 -14575 -66421
rect -14775 -66485 -14575 -66438
rect -14517 -66438 -14467 -66421
rect -14367 -66421 -14351 -66404
rect -14225 -66404 -14093 -66388
rect -14225 -66421 -14209 -66404
rect -14367 -66438 -14317 -66421
rect -14517 -66485 -14317 -66438
rect -14259 -66438 -14209 -66421
rect -14109 -66421 -14093 -66404
rect -13967 -66404 -13835 -66388
rect -13967 -66421 -13951 -66404
rect -14109 -66438 -14059 -66421
rect -14259 -66485 -14059 -66438
rect -14001 -66438 -13951 -66421
rect -13851 -66421 -13835 -66404
rect -13851 -66438 -13801 -66421
rect -14001 -66485 -13801 -66438
rect -15291 -66932 -15091 -66885
rect -15291 -66949 -15241 -66932
rect -15257 -66966 -15241 -66949
rect -15141 -66949 -15091 -66932
rect -15033 -66932 -14833 -66885
rect -15033 -66949 -14983 -66932
rect -15141 -66966 -15125 -66949
rect -15257 -66982 -15125 -66966
rect -14999 -66966 -14983 -66949
rect -14883 -66949 -14833 -66932
rect -14775 -66932 -14575 -66885
rect -14775 -66949 -14725 -66932
rect -14883 -66966 -14867 -66949
rect -14999 -66982 -14867 -66966
rect -14741 -66966 -14725 -66949
rect -14625 -66949 -14575 -66932
rect -14517 -66932 -14317 -66885
rect -14517 -66949 -14467 -66932
rect -14625 -66966 -14609 -66949
rect -14741 -66982 -14609 -66966
rect -14483 -66966 -14467 -66949
rect -14367 -66949 -14317 -66932
rect -14259 -66932 -14059 -66885
rect -14259 -66949 -14209 -66932
rect -14367 -66966 -14351 -66949
rect -14483 -66982 -14351 -66966
rect -14225 -66966 -14209 -66949
rect -14109 -66949 -14059 -66932
rect -14001 -66932 -13801 -66885
rect -14001 -66949 -13951 -66932
rect -14109 -66966 -14093 -66949
rect -14225 -66982 -14093 -66966
rect -13967 -66966 -13951 -66949
rect -13851 -66949 -13801 -66932
rect -13851 -66966 -13835 -66949
rect -13967 -66982 -13835 -66966
rect -11952 -67329 -11922 -67303
rect -15952 -67561 -15922 -67529
rect -11257 -65544 -11125 -65528
rect -11257 -65561 -11241 -65544
rect -11291 -65578 -11241 -65561
rect -11141 -65561 -11125 -65544
rect -10999 -65544 -10867 -65528
rect -10999 -65561 -10983 -65544
rect -11141 -65578 -11091 -65561
rect -11291 -65625 -11091 -65578
rect -11033 -65578 -10983 -65561
rect -10883 -65561 -10867 -65544
rect -10741 -65544 -10609 -65528
rect -10741 -65561 -10725 -65544
rect -10883 -65578 -10833 -65561
rect -11033 -65625 -10833 -65578
rect -10775 -65578 -10725 -65561
rect -10625 -65561 -10609 -65544
rect -10483 -65544 -10351 -65528
rect -10483 -65561 -10467 -65544
rect -10625 -65578 -10575 -65561
rect -10775 -65625 -10575 -65578
rect -10517 -65578 -10467 -65561
rect -10367 -65561 -10351 -65544
rect -10225 -65544 -10093 -65528
rect -10225 -65561 -10209 -65544
rect -10367 -65578 -10317 -65561
rect -10517 -65625 -10317 -65578
rect -10259 -65578 -10209 -65561
rect -10109 -65561 -10093 -65544
rect -9967 -65544 -9835 -65528
rect -9967 -65561 -9951 -65544
rect -10109 -65578 -10059 -65561
rect -10259 -65625 -10059 -65578
rect -10001 -65578 -9951 -65561
rect -9851 -65561 -9835 -65544
rect -9851 -65578 -9801 -65561
rect -10001 -65625 -9801 -65578
rect -11291 -66072 -11091 -66025
rect -11291 -66089 -11241 -66072
rect -11257 -66106 -11241 -66089
rect -11141 -66089 -11091 -66072
rect -11033 -66072 -10833 -66025
rect -11033 -66089 -10983 -66072
rect -11141 -66106 -11125 -66089
rect -11257 -66122 -11125 -66106
rect -10999 -66106 -10983 -66089
rect -10883 -66089 -10833 -66072
rect -10775 -66072 -10575 -66025
rect -10775 -66089 -10725 -66072
rect -10883 -66106 -10867 -66089
rect -10999 -66122 -10867 -66106
rect -10741 -66106 -10725 -66089
rect -10625 -66089 -10575 -66072
rect -10517 -66072 -10317 -66025
rect -10517 -66089 -10467 -66072
rect -10625 -66106 -10609 -66089
rect -10741 -66122 -10609 -66106
rect -10483 -66106 -10467 -66089
rect -10367 -66089 -10317 -66072
rect -10259 -66072 -10059 -66025
rect -10259 -66089 -10209 -66072
rect -10367 -66106 -10351 -66089
rect -10483 -66122 -10351 -66106
rect -10225 -66106 -10209 -66089
rect -10109 -66089 -10059 -66072
rect -10001 -66072 -9801 -66025
rect -10001 -66089 -9951 -66072
rect -10109 -66106 -10093 -66089
rect -10225 -66122 -10093 -66106
rect -9967 -66106 -9951 -66089
rect -9851 -66089 -9801 -66072
rect -9851 -66106 -9835 -66089
rect -9967 -66122 -9835 -66106
rect -11257 -66404 -11125 -66388
rect -11257 -66421 -11241 -66404
rect -11291 -66438 -11241 -66421
rect -11141 -66421 -11125 -66404
rect -10999 -66404 -10867 -66388
rect -10999 -66421 -10983 -66404
rect -11141 -66438 -11091 -66421
rect -11291 -66485 -11091 -66438
rect -11033 -66438 -10983 -66421
rect -10883 -66421 -10867 -66404
rect -10741 -66404 -10609 -66388
rect -10741 -66421 -10725 -66404
rect -10883 -66438 -10833 -66421
rect -11033 -66485 -10833 -66438
rect -10775 -66438 -10725 -66421
rect -10625 -66421 -10609 -66404
rect -10483 -66404 -10351 -66388
rect -10483 -66421 -10467 -66404
rect -10625 -66438 -10575 -66421
rect -10775 -66485 -10575 -66438
rect -10517 -66438 -10467 -66421
rect -10367 -66421 -10351 -66404
rect -10225 -66404 -10093 -66388
rect -10225 -66421 -10209 -66404
rect -10367 -66438 -10317 -66421
rect -10517 -66485 -10317 -66438
rect -10259 -66438 -10209 -66421
rect -10109 -66421 -10093 -66404
rect -9967 -66404 -9835 -66388
rect -9967 -66421 -9951 -66404
rect -10109 -66438 -10059 -66421
rect -10259 -66485 -10059 -66438
rect -10001 -66438 -9951 -66421
rect -9851 -66421 -9835 -66404
rect -9851 -66438 -9801 -66421
rect -10001 -66485 -9801 -66438
rect -11291 -66932 -11091 -66885
rect -11291 -66949 -11241 -66932
rect -11257 -66966 -11241 -66949
rect -11141 -66949 -11091 -66932
rect -11033 -66932 -10833 -66885
rect -11033 -66949 -10983 -66932
rect -11141 -66966 -11125 -66949
rect -11257 -66982 -11125 -66966
rect -10999 -66966 -10983 -66949
rect -10883 -66949 -10833 -66932
rect -10775 -66932 -10575 -66885
rect -10775 -66949 -10725 -66932
rect -10883 -66966 -10867 -66949
rect -10999 -66982 -10867 -66966
rect -10741 -66966 -10725 -66949
rect -10625 -66949 -10575 -66932
rect -10517 -66932 -10317 -66885
rect -10517 -66949 -10467 -66932
rect -10625 -66966 -10609 -66949
rect -10741 -66982 -10609 -66966
rect -10483 -66966 -10467 -66949
rect -10367 -66949 -10317 -66932
rect -10259 -66932 -10059 -66885
rect -10259 -66949 -10209 -66932
rect -10367 -66966 -10351 -66949
rect -10483 -66982 -10351 -66966
rect -10225 -66966 -10209 -66949
rect -10109 -66949 -10059 -66932
rect -10001 -66932 -9801 -66885
rect -10001 -66949 -9951 -66932
rect -10109 -66966 -10093 -66949
rect -10225 -66982 -10093 -66966
rect -9967 -66966 -9951 -66949
rect -9851 -66949 -9801 -66932
rect -9851 -66966 -9835 -66949
rect -9967 -66982 -9835 -66966
rect -7952 -67329 -7922 -67303
rect -11952 -67561 -11922 -67529
rect -7257 -65544 -7125 -65528
rect -7257 -65561 -7241 -65544
rect -7291 -65578 -7241 -65561
rect -7141 -65561 -7125 -65544
rect -6999 -65544 -6867 -65528
rect -6999 -65561 -6983 -65544
rect -7141 -65578 -7091 -65561
rect -7291 -65625 -7091 -65578
rect -7033 -65578 -6983 -65561
rect -6883 -65561 -6867 -65544
rect -6741 -65544 -6609 -65528
rect -6741 -65561 -6725 -65544
rect -6883 -65578 -6833 -65561
rect -7033 -65625 -6833 -65578
rect -6775 -65578 -6725 -65561
rect -6625 -65561 -6609 -65544
rect -6483 -65544 -6351 -65528
rect -6483 -65561 -6467 -65544
rect -6625 -65578 -6575 -65561
rect -6775 -65625 -6575 -65578
rect -6517 -65578 -6467 -65561
rect -6367 -65561 -6351 -65544
rect -6225 -65544 -6093 -65528
rect -6225 -65561 -6209 -65544
rect -6367 -65578 -6317 -65561
rect -6517 -65625 -6317 -65578
rect -6259 -65578 -6209 -65561
rect -6109 -65561 -6093 -65544
rect -5967 -65544 -5835 -65528
rect -5967 -65561 -5951 -65544
rect -6109 -65578 -6059 -65561
rect -6259 -65625 -6059 -65578
rect -6001 -65578 -5951 -65561
rect -5851 -65561 -5835 -65544
rect -5851 -65578 -5801 -65561
rect -6001 -65625 -5801 -65578
rect -7291 -66072 -7091 -66025
rect -7291 -66089 -7241 -66072
rect -7257 -66106 -7241 -66089
rect -7141 -66089 -7091 -66072
rect -7033 -66072 -6833 -66025
rect -7033 -66089 -6983 -66072
rect -7141 -66106 -7125 -66089
rect -7257 -66122 -7125 -66106
rect -6999 -66106 -6983 -66089
rect -6883 -66089 -6833 -66072
rect -6775 -66072 -6575 -66025
rect -6775 -66089 -6725 -66072
rect -6883 -66106 -6867 -66089
rect -6999 -66122 -6867 -66106
rect -6741 -66106 -6725 -66089
rect -6625 -66089 -6575 -66072
rect -6517 -66072 -6317 -66025
rect -6517 -66089 -6467 -66072
rect -6625 -66106 -6609 -66089
rect -6741 -66122 -6609 -66106
rect -6483 -66106 -6467 -66089
rect -6367 -66089 -6317 -66072
rect -6259 -66072 -6059 -66025
rect -6259 -66089 -6209 -66072
rect -6367 -66106 -6351 -66089
rect -6483 -66122 -6351 -66106
rect -6225 -66106 -6209 -66089
rect -6109 -66089 -6059 -66072
rect -6001 -66072 -5801 -66025
rect -6001 -66089 -5951 -66072
rect -6109 -66106 -6093 -66089
rect -6225 -66122 -6093 -66106
rect -5967 -66106 -5951 -66089
rect -5851 -66089 -5801 -66072
rect -5851 -66106 -5835 -66089
rect -5967 -66122 -5835 -66106
rect -7257 -66404 -7125 -66388
rect -7257 -66421 -7241 -66404
rect -7291 -66438 -7241 -66421
rect -7141 -66421 -7125 -66404
rect -6999 -66404 -6867 -66388
rect -6999 -66421 -6983 -66404
rect -7141 -66438 -7091 -66421
rect -7291 -66485 -7091 -66438
rect -7033 -66438 -6983 -66421
rect -6883 -66421 -6867 -66404
rect -6741 -66404 -6609 -66388
rect -6741 -66421 -6725 -66404
rect -6883 -66438 -6833 -66421
rect -7033 -66485 -6833 -66438
rect -6775 -66438 -6725 -66421
rect -6625 -66421 -6609 -66404
rect -6483 -66404 -6351 -66388
rect -6483 -66421 -6467 -66404
rect -6625 -66438 -6575 -66421
rect -6775 -66485 -6575 -66438
rect -6517 -66438 -6467 -66421
rect -6367 -66421 -6351 -66404
rect -6225 -66404 -6093 -66388
rect -6225 -66421 -6209 -66404
rect -6367 -66438 -6317 -66421
rect -6517 -66485 -6317 -66438
rect -6259 -66438 -6209 -66421
rect -6109 -66421 -6093 -66404
rect -5967 -66404 -5835 -66388
rect -5967 -66421 -5951 -66404
rect -6109 -66438 -6059 -66421
rect -6259 -66485 -6059 -66438
rect -6001 -66438 -5951 -66421
rect -5851 -66421 -5835 -66404
rect -5851 -66438 -5801 -66421
rect -6001 -66485 -5801 -66438
rect -7291 -66932 -7091 -66885
rect -7291 -66949 -7241 -66932
rect -7257 -66966 -7241 -66949
rect -7141 -66949 -7091 -66932
rect -7033 -66932 -6833 -66885
rect -7033 -66949 -6983 -66932
rect -7141 -66966 -7125 -66949
rect -7257 -66982 -7125 -66966
rect -6999 -66966 -6983 -66949
rect -6883 -66949 -6833 -66932
rect -6775 -66932 -6575 -66885
rect -6775 -66949 -6725 -66932
rect -6883 -66966 -6867 -66949
rect -6999 -66982 -6867 -66966
rect -6741 -66966 -6725 -66949
rect -6625 -66949 -6575 -66932
rect -6517 -66932 -6317 -66885
rect -6517 -66949 -6467 -66932
rect -6625 -66966 -6609 -66949
rect -6741 -66982 -6609 -66966
rect -6483 -66966 -6467 -66949
rect -6367 -66949 -6317 -66932
rect -6259 -66932 -6059 -66885
rect -6259 -66949 -6209 -66932
rect -6367 -66966 -6351 -66949
rect -6483 -66982 -6351 -66966
rect -6225 -66966 -6209 -66949
rect -6109 -66949 -6059 -66932
rect -6001 -66932 -5801 -66885
rect -6001 -66949 -5951 -66932
rect -6109 -66966 -6093 -66949
rect -6225 -66982 -6093 -66966
rect -5967 -66966 -5951 -66949
rect -5851 -66949 -5801 -66932
rect -5851 -66966 -5835 -66949
rect -5967 -66982 -5835 -66966
rect -3952 -67329 -3922 -67303
rect -7952 -67561 -7922 -67529
rect -3257 -65544 -3125 -65528
rect -3257 -65561 -3241 -65544
rect -3291 -65578 -3241 -65561
rect -3141 -65561 -3125 -65544
rect -2999 -65544 -2867 -65528
rect -2999 -65561 -2983 -65544
rect -3141 -65578 -3091 -65561
rect -3291 -65625 -3091 -65578
rect -3033 -65578 -2983 -65561
rect -2883 -65561 -2867 -65544
rect -2741 -65544 -2609 -65528
rect -2741 -65561 -2725 -65544
rect -2883 -65578 -2833 -65561
rect -3033 -65625 -2833 -65578
rect -2775 -65578 -2725 -65561
rect -2625 -65561 -2609 -65544
rect -2483 -65544 -2351 -65528
rect -2483 -65561 -2467 -65544
rect -2625 -65578 -2575 -65561
rect -2775 -65625 -2575 -65578
rect -2517 -65578 -2467 -65561
rect -2367 -65561 -2351 -65544
rect -2225 -65544 -2093 -65528
rect -2225 -65561 -2209 -65544
rect -2367 -65578 -2317 -65561
rect -2517 -65625 -2317 -65578
rect -2259 -65578 -2209 -65561
rect -2109 -65561 -2093 -65544
rect -1967 -65544 -1835 -65528
rect -1967 -65561 -1951 -65544
rect -2109 -65578 -2059 -65561
rect -2259 -65625 -2059 -65578
rect -2001 -65578 -1951 -65561
rect -1851 -65561 -1835 -65544
rect -1851 -65578 -1801 -65561
rect -2001 -65625 -1801 -65578
rect -3291 -66072 -3091 -66025
rect -3291 -66089 -3241 -66072
rect -3257 -66106 -3241 -66089
rect -3141 -66089 -3091 -66072
rect -3033 -66072 -2833 -66025
rect -3033 -66089 -2983 -66072
rect -3141 -66106 -3125 -66089
rect -3257 -66122 -3125 -66106
rect -2999 -66106 -2983 -66089
rect -2883 -66089 -2833 -66072
rect -2775 -66072 -2575 -66025
rect -2775 -66089 -2725 -66072
rect -2883 -66106 -2867 -66089
rect -2999 -66122 -2867 -66106
rect -2741 -66106 -2725 -66089
rect -2625 -66089 -2575 -66072
rect -2517 -66072 -2317 -66025
rect -2517 -66089 -2467 -66072
rect -2625 -66106 -2609 -66089
rect -2741 -66122 -2609 -66106
rect -2483 -66106 -2467 -66089
rect -2367 -66089 -2317 -66072
rect -2259 -66072 -2059 -66025
rect -2259 -66089 -2209 -66072
rect -2367 -66106 -2351 -66089
rect -2483 -66122 -2351 -66106
rect -2225 -66106 -2209 -66089
rect -2109 -66089 -2059 -66072
rect -2001 -66072 -1801 -66025
rect -2001 -66089 -1951 -66072
rect -2109 -66106 -2093 -66089
rect -2225 -66122 -2093 -66106
rect -1967 -66106 -1951 -66089
rect -1851 -66089 -1801 -66072
rect -1851 -66106 -1835 -66089
rect -1967 -66122 -1835 -66106
rect -3257 -66404 -3125 -66388
rect -3257 -66421 -3241 -66404
rect -3291 -66438 -3241 -66421
rect -3141 -66421 -3125 -66404
rect -2999 -66404 -2867 -66388
rect -2999 -66421 -2983 -66404
rect -3141 -66438 -3091 -66421
rect -3291 -66485 -3091 -66438
rect -3033 -66438 -2983 -66421
rect -2883 -66421 -2867 -66404
rect -2741 -66404 -2609 -66388
rect -2741 -66421 -2725 -66404
rect -2883 -66438 -2833 -66421
rect -3033 -66485 -2833 -66438
rect -2775 -66438 -2725 -66421
rect -2625 -66421 -2609 -66404
rect -2483 -66404 -2351 -66388
rect -2483 -66421 -2467 -66404
rect -2625 -66438 -2575 -66421
rect -2775 -66485 -2575 -66438
rect -2517 -66438 -2467 -66421
rect -2367 -66421 -2351 -66404
rect -2225 -66404 -2093 -66388
rect -2225 -66421 -2209 -66404
rect -2367 -66438 -2317 -66421
rect -2517 -66485 -2317 -66438
rect -2259 -66438 -2209 -66421
rect -2109 -66421 -2093 -66404
rect -1967 -66404 -1835 -66388
rect -1967 -66421 -1951 -66404
rect -2109 -66438 -2059 -66421
rect -2259 -66485 -2059 -66438
rect -2001 -66438 -1951 -66421
rect -1851 -66421 -1835 -66404
rect -1851 -66438 -1801 -66421
rect -2001 -66485 -1801 -66438
rect -3291 -66932 -3091 -66885
rect -3291 -66949 -3241 -66932
rect -3257 -66966 -3241 -66949
rect -3141 -66949 -3091 -66932
rect -3033 -66932 -2833 -66885
rect -3033 -66949 -2983 -66932
rect -3141 -66966 -3125 -66949
rect -3257 -66982 -3125 -66966
rect -2999 -66966 -2983 -66949
rect -2883 -66949 -2833 -66932
rect -2775 -66932 -2575 -66885
rect -2775 -66949 -2725 -66932
rect -2883 -66966 -2867 -66949
rect -2999 -66982 -2867 -66966
rect -2741 -66966 -2725 -66949
rect -2625 -66949 -2575 -66932
rect -2517 -66932 -2317 -66885
rect -2517 -66949 -2467 -66932
rect -2625 -66966 -2609 -66949
rect -2741 -66982 -2609 -66966
rect -2483 -66966 -2467 -66949
rect -2367 -66949 -2317 -66932
rect -2259 -66932 -2059 -66885
rect -2259 -66949 -2209 -66932
rect -2367 -66966 -2351 -66949
rect -2483 -66982 -2351 -66966
rect -2225 -66966 -2209 -66949
rect -2109 -66949 -2059 -66932
rect -2001 -66932 -1801 -66885
rect -2001 -66949 -1951 -66932
rect -2109 -66966 -2093 -66949
rect -2225 -66982 -2093 -66966
rect -1967 -66966 -1951 -66949
rect -1851 -66949 -1801 -66932
rect -1851 -66966 -1835 -66949
rect -1967 -66982 -1835 -66966
rect 48 -67329 78 -67303
rect -3952 -67561 -3922 -67529
rect 743 -65544 875 -65528
rect 743 -65561 759 -65544
rect 709 -65578 759 -65561
rect 859 -65561 875 -65544
rect 1001 -65544 1133 -65528
rect 1001 -65561 1017 -65544
rect 859 -65578 909 -65561
rect 709 -65625 909 -65578
rect 967 -65578 1017 -65561
rect 1117 -65561 1133 -65544
rect 1259 -65544 1391 -65528
rect 1259 -65561 1275 -65544
rect 1117 -65578 1167 -65561
rect 967 -65625 1167 -65578
rect 1225 -65578 1275 -65561
rect 1375 -65561 1391 -65544
rect 1517 -65544 1649 -65528
rect 1517 -65561 1533 -65544
rect 1375 -65578 1425 -65561
rect 1225 -65625 1425 -65578
rect 1483 -65578 1533 -65561
rect 1633 -65561 1649 -65544
rect 1775 -65544 1907 -65528
rect 1775 -65561 1791 -65544
rect 1633 -65578 1683 -65561
rect 1483 -65625 1683 -65578
rect 1741 -65578 1791 -65561
rect 1891 -65561 1907 -65544
rect 2033 -65544 2165 -65528
rect 2033 -65561 2049 -65544
rect 1891 -65578 1941 -65561
rect 1741 -65625 1941 -65578
rect 1999 -65578 2049 -65561
rect 2149 -65561 2165 -65544
rect 2149 -65578 2199 -65561
rect 1999 -65625 2199 -65578
rect 709 -66072 909 -66025
rect 709 -66089 759 -66072
rect 743 -66106 759 -66089
rect 859 -66089 909 -66072
rect 967 -66072 1167 -66025
rect 967 -66089 1017 -66072
rect 859 -66106 875 -66089
rect 743 -66122 875 -66106
rect 1001 -66106 1017 -66089
rect 1117 -66089 1167 -66072
rect 1225 -66072 1425 -66025
rect 1225 -66089 1275 -66072
rect 1117 -66106 1133 -66089
rect 1001 -66122 1133 -66106
rect 1259 -66106 1275 -66089
rect 1375 -66089 1425 -66072
rect 1483 -66072 1683 -66025
rect 1483 -66089 1533 -66072
rect 1375 -66106 1391 -66089
rect 1259 -66122 1391 -66106
rect 1517 -66106 1533 -66089
rect 1633 -66089 1683 -66072
rect 1741 -66072 1941 -66025
rect 1741 -66089 1791 -66072
rect 1633 -66106 1649 -66089
rect 1517 -66122 1649 -66106
rect 1775 -66106 1791 -66089
rect 1891 -66089 1941 -66072
rect 1999 -66072 2199 -66025
rect 1999 -66089 2049 -66072
rect 1891 -66106 1907 -66089
rect 1775 -66122 1907 -66106
rect 2033 -66106 2049 -66089
rect 2149 -66089 2199 -66072
rect 2149 -66106 2165 -66089
rect 2033 -66122 2165 -66106
rect 743 -66404 875 -66388
rect 743 -66421 759 -66404
rect 709 -66438 759 -66421
rect 859 -66421 875 -66404
rect 1001 -66404 1133 -66388
rect 1001 -66421 1017 -66404
rect 859 -66438 909 -66421
rect 709 -66485 909 -66438
rect 967 -66438 1017 -66421
rect 1117 -66421 1133 -66404
rect 1259 -66404 1391 -66388
rect 1259 -66421 1275 -66404
rect 1117 -66438 1167 -66421
rect 967 -66485 1167 -66438
rect 1225 -66438 1275 -66421
rect 1375 -66421 1391 -66404
rect 1517 -66404 1649 -66388
rect 1517 -66421 1533 -66404
rect 1375 -66438 1425 -66421
rect 1225 -66485 1425 -66438
rect 1483 -66438 1533 -66421
rect 1633 -66421 1649 -66404
rect 1775 -66404 1907 -66388
rect 1775 -66421 1791 -66404
rect 1633 -66438 1683 -66421
rect 1483 -66485 1683 -66438
rect 1741 -66438 1791 -66421
rect 1891 -66421 1907 -66404
rect 2033 -66404 2165 -66388
rect 2033 -66421 2049 -66404
rect 1891 -66438 1941 -66421
rect 1741 -66485 1941 -66438
rect 1999 -66438 2049 -66421
rect 2149 -66421 2165 -66404
rect 2149 -66438 2199 -66421
rect 1999 -66485 2199 -66438
rect 709 -66932 909 -66885
rect 709 -66949 759 -66932
rect 743 -66966 759 -66949
rect 859 -66949 909 -66932
rect 967 -66932 1167 -66885
rect 967 -66949 1017 -66932
rect 859 -66966 875 -66949
rect 743 -66982 875 -66966
rect 1001 -66966 1017 -66949
rect 1117 -66949 1167 -66932
rect 1225 -66932 1425 -66885
rect 1225 -66949 1275 -66932
rect 1117 -66966 1133 -66949
rect 1001 -66982 1133 -66966
rect 1259 -66966 1275 -66949
rect 1375 -66949 1425 -66932
rect 1483 -66932 1683 -66885
rect 1483 -66949 1533 -66932
rect 1375 -66966 1391 -66949
rect 1259 -66982 1391 -66966
rect 1517 -66966 1533 -66949
rect 1633 -66949 1683 -66932
rect 1741 -66932 1941 -66885
rect 1741 -66949 1791 -66932
rect 1633 -66966 1649 -66949
rect 1517 -66982 1649 -66966
rect 1775 -66966 1791 -66949
rect 1891 -66949 1941 -66932
rect 1999 -66932 2199 -66885
rect 1999 -66949 2049 -66932
rect 1891 -66966 1907 -66949
rect 1775 -66982 1907 -66966
rect 2033 -66966 2049 -66949
rect 2149 -66949 2199 -66932
rect 2149 -66966 2165 -66949
rect 2033 -66982 2165 -66966
rect 4048 -67329 4078 -67303
rect 48 -67561 78 -67529
rect 4743 -65544 4875 -65528
rect 4743 -65561 4759 -65544
rect 4709 -65578 4759 -65561
rect 4859 -65561 4875 -65544
rect 5001 -65544 5133 -65528
rect 5001 -65561 5017 -65544
rect 4859 -65578 4909 -65561
rect 4709 -65625 4909 -65578
rect 4967 -65578 5017 -65561
rect 5117 -65561 5133 -65544
rect 5259 -65544 5391 -65528
rect 5259 -65561 5275 -65544
rect 5117 -65578 5167 -65561
rect 4967 -65625 5167 -65578
rect 5225 -65578 5275 -65561
rect 5375 -65561 5391 -65544
rect 5517 -65544 5649 -65528
rect 5517 -65561 5533 -65544
rect 5375 -65578 5425 -65561
rect 5225 -65625 5425 -65578
rect 5483 -65578 5533 -65561
rect 5633 -65561 5649 -65544
rect 5775 -65544 5907 -65528
rect 5775 -65561 5791 -65544
rect 5633 -65578 5683 -65561
rect 5483 -65625 5683 -65578
rect 5741 -65578 5791 -65561
rect 5891 -65561 5907 -65544
rect 6033 -65544 6165 -65528
rect 6033 -65561 6049 -65544
rect 5891 -65578 5941 -65561
rect 5741 -65625 5941 -65578
rect 5999 -65578 6049 -65561
rect 6149 -65561 6165 -65544
rect 6149 -65578 6199 -65561
rect 5999 -65625 6199 -65578
rect 4709 -66072 4909 -66025
rect 4709 -66089 4759 -66072
rect 4743 -66106 4759 -66089
rect 4859 -66089 4909 -66072
rect 4967 -66072 5167 -66025
rect 4967 -66089 5017 -66072
rect 4859 -66106 4875 -66089
rect 4743 -66122 4875 -66106
rect 5001 -66106 5017 -66089
rect 5117 -66089 5167 -66072
rect 5225 -66072 5425 -66025
rect 5225 -66089 5275 -66072
rect 5117 -66106 5133 -66089
rect 5001 -66122 5133 -66106
rect 5259 -66106 5275 -66089
rect 5375 -66089 5425 -66072
rect 5483 -66072 5683 -66025
rect 5483 -66089 5533 -66072
rect 5375 -66106 5391 -66089
rect 5259 -66122 5391 -66106
rect 5517 -66106 5533 -66089
rect 5633 -66089 5683 -66072
rect 5741 -66072 5941 -66025
rect 5741 -66089 5791 -66072
rect 5633 -66106 5649 -66089
rect 5517 -66122 5649 -66106
rect 5775 -66106 5791 -66089
rect 5891 -66089 5941 -66072
rect 5999 -66072 6199 -66025
rect 5999 -66089 6049 -66072
rect 5891 -66106 5907 -66089
rect 5775 -66122 5907 -66106
rect 6033 -66106 6049 -66089
rect 6149 -66089 6199 -66072
rect 6149 -66106 6165 -66089
rect 6033 -66122 6165 -66106
rect 4743 -66404 4875 -66388
rect 4743 -66421 4759 -66404
rect 4709 -66438 4759 -66421
rect 4859 -66421 4875 -66404
rect 5001 -66404 5133 -66388
rect 5001 -66421 5017 -66404
rect 4859 -66438 4909 -66421
rect 4709 -66485 4909 -66438
rect 4967 -66438 5017 -66421
rect 5117 -66421 5133 -66404
rect 5259 -66404 5391 -66388
rect 5259 -66421 5275 -66404
rect 5117 -66438 5167 -66421
rect 4967 -66485 5167 -66438
rect 5225 -66438 5275 -66421
rect 5375 -66421 5391 -66404
rect 5517 -66404 5649 -66388
rect 5517 -66421 5533 -66404
rect 5375 -66438 5425 -66421
rect 5225 -66485 5425 -66438
rect 5483 -66438 5533 -66421
rect 5633 -66421 5649 -66404
rect 5775 -66404 5907 -66388
rect 5775 -66421 5791 -66404
rect 5633 -66438 5683 -66421
rect 5483 -66485 5683 -66438
rect 5741 -66438 5791 -66421
rect 5891 -66421 5907 -66404
rect 6033 -66404 6165 -66388
rect 6033 -66421 6049 -66404
rect 5891 -66438 5941 -66421
rect 5741 -66485 5941 -66438
rect 5999 -66438 6049 -66421
rect 6149 -66421 6165 -66404
rect 6149 -66438 6199 -66421
rect 5999 -66485 6199 -66438
rect 4709 -66932 4909 -66885
rect 4709 -66949 4759 -66932
rect 4743 -66966 4759 -66949
rect 4859 -66949 4909 -66932
rect 4967 -66932 5167 -66885
rect 4967 -66949 5017 -66932
rect 4859 -66966 4875 -66949
rect 4743 -66982 4875 -66966
rect 5001 -66966 5017 -66949
rect 5117 -66949 5167 -66932
rect 5225 -66932 5425 -66885
rect 5225 -66949 5275 -66932
rect 5117 -66966 5133 -66949
rect 5001 -66982 5133 -66966
rect 5259 -66966 5275 -66949
rect 5375 -66949 5425 -66932
rect 5483 -66932 5683 -66885
rect 5483 -66949 5533 -66932
rect 5375 -66966 5391 -66949
rect 5259 -66982 5391 -66966
rect 5517 -66966 5533 -66949
rect 5633 -66949 5683 -66932
rect 5741 -66932 5941 -66885
rect 5741 -66949 5791 -66932
rect 5633 -66966 5649 -66949
rect 5517 -66982 5649 -66966
rect 5775 -66966 5791 -66949
rect 5891 -66949 5941 -66932
rect 5999 -66932 6199 -66885
rect 5999 -66949 6049 -66932
rect 5891 -66966 5907 -66949
rect 5775 -66982 5907 -66966
rect 6033 -66966 6049 -66949
rect 6149 -66949 6199 -66932
rect 6149 -66966 6165 -66949
rect 6033 -66982 6165 -66966
rect 4048 -67561 4078 -67529
rect -28008 -67577 -27922 -67561
rect -28008 -67611 -27992 -67577
rect -27958 -67611 -27922 -67577
rect -28008 -67627 -27922 -67611
rect -24008 -67577 -23922 -67561
rect -24008 -67611 -23992 -67577
rect -23958 -67611 -23922 -67577
rect -24008 -67627 -23922 -67611
rect -20008 -67577 -19922 -67561
rect -20008 -67611 -19992 -67577
rect -19958 -67611 -19922 -67577
rect -20008 -67627 -19922 -67611
rect -16008 -67577 -15922 -67561
rect -16008 -67611 -15992 -67577
rect -15958 -67611 -15922 -67577
rect -16008 -67627 -15922 -67611
rect -12008 -67577 -11922 -67561
rect -12008 -67611 -11992 -67577
rect -11958 -67611 -11922 -67577
rect -12008 -67627 -11922 -67611
rect -8008 -67577 -7922 -67561
rect -8008 -67611 -7992 -67577
rect -7958 -67611 -7922 -67577
rect -8008 -67627 -7922 -67611
rect -4008 -67577 -3922 -67561
rect -4008 -67611 -3992 -67577
rect -3958 -67611 -3922 -67577
rect -4008 -67627 -3922 -67611
rect -8 -67577 78 -67561
rect -8 -67611 8 -67577
rect 42 -67611 78 -67577
rect -8 -67627 78 -67611
rect 3992 -67577 4078 -67561
rect 3992 -67611 4008 -67577
rect 4042 -67611 4078 -67577
rect 3992 -67627 4078 -67611
rect -27952 -67649 -27922 -67627
rect -23952 -67649 -23922 -67627
rect -19952 -67649 -19922 -67627
rect -15952 -67649 -15922 -67627
rect -11952 -67649 -11922 -67627
rect -7952 -67649 -7922 -67627
rect -3952 -67649 -3922 -67627
rect 48 -67649 78 -67627
rect 4048 -67649 4078 -67627
rect -27952 -67805 -27922 -67779
rect -23952 -67805 -23922 -67779
rect -27262 -68246 -27130 -68230
rect -27262 -68263 -27246 -68246
rect -27296 -68280 -27246 -68263
rect -27146 -68263 -27130 -68246
rect -27004 -68246 -26872 -68230
rect -27004 -68263 -26988 -68246
rect -27146 -68280 -27096 -68263
rect -27296 -68318 -27096 -68280
rect -27038 -68280 -26988 -68263
rect -26888 -68263 -26872 -68246
rect -26746 -68246 -26614 -68230
rect -26746 -68263 -26730 -68246
rect -26888 -68280 -26838 -68263
rect -27038 -68318 -26838 -68280
rect -26780 -68280 -26730 -68263
rect -26630 -68263 -26614 -68246
rect -26488 -68246 -26356 -68230
rect -26488 -68263 -26472 -68246
rect -26630 -68280 -26580 -68263
rect -26780 -68318 -26580 -68280
rect -26522 -68280 -26472 -68263
rect -26372 -68263 -26356 -68246
rect -26230 -68246 -26098 -68230
rect -26230 -68263 -26214 -68246
rect -26372 -68280 -26322 -68263
rect -26522 -68318 -26322 -68280
rect -26264 -68280 -26214 -68263
rect -26114 -68263 -26098 -68246
rect -25972 -68246 -25840 -68230
rect -25972 -68263 -25956 -68246
rect -26114 -68280 -26064 -68263
rect -26264 -68318 -26064 -68280
rect -26006 -68280 -25956 -68263
rect -25856 -68263 -25840 -68246
rect -25856 -68280 -25806 -68263
rect -26006 -68318 -25806 -68280
rect -27296 -68756 -27096 -68718
rect -27296 -68773 -27246 -68756
rect -27262 -68790 -27246 -68773
rect -27146 -68773 -27096 -68756
rect -27038 -68756 -26838 -68718
rect -27038 -68773 -26988 -68756
rect -27146 -68790 -27130 -68773
rect -27262 -68806 -27130 -68790
rect -27004 -68790 -26988 -68773
rect -26888 -68773 -26838 -68756
rect -26780 -68756 -26580 -68718
rect -26780 -68773 -26730 -68756
rect -26888 -68790 -26872 -68773
rect -27004 -68806 -26872 -68790
rect -26746 -68790 -26730 -68773
rect -26630 -68773 -26580 -68756
rect -26522 -68756 -26322 -68718
rect -26522 -68773 -26472 -68756
rect -26630 -68790 -26614 -68773
rect -26746 -68806 -26614 -68790
rect -26488 -68790 -26472 -68773
rect -26372 -68773 -26322 -68756
rect -26264 -68756 -26064 -68718
rect -26264 -68773 -26214 -68756
rect -26372 -68790 -26356 -68773
rect -26488 -68806 -26356 -68790
rect -26230 -68790 -26214 -68773
rect -26114 -68773 -26064 -68756
rect -26006 -68756 -25806 -68718
rect -26006 -68773 -25956 -68756
rect -26114 -68790 -26098 -68773
rect -26230 -68806 -26098 -68790
rect -25972 -68790 -25956 -68773
rect -25856 -68773 -25806 -68756
rect -25856 -68790 -25840 -68773
rect -25972 -68806 -25840 -68790
rect -19952 -67805 -19922 -67779
rect -23262 -68246 -23130 -68230
rect -23262 -68263 -23246 -68246
rect -23296 -68280 -23246 -68263
rect -23146 -68263 -23130 -68246
rect -23004 -68246 -22872 -68230
rect -23004 -68263 -22988 -68246
rect -23146 -68280 -23096 -68263
rect -23296 -68318 -23096 -68280
rect -23038 -68280 -22988 -68263
rect -22888 -68263 -22872 -68246
rect -22746 -68246 -22614 -68230
rect -22746 -68263 -22730 -68246
rect -22888 -68280 -22838 -68263
rect -23038 -68318 -22838 -68280
rect -22780 -68280 -22730 -68263
rect -22630 -68263 -22614 -68246
rect -22488 -68246 -22356 -68230
rect -22488 -68263 -22472 -68246
rect -22630 -68280 -22580 -68263
rect -22780 -68318 -22580 -68280
rect -22522 -68280 -22472 -68263
rect -22372 -68263 -22356 -68246
rect -22230 -68246 -22098 -68230
rect -22230 -68263 -22214 -68246
rect -22372 -68280 -22322 -68263
rect -22522 -68318 -22322 -68280
rect -22264 -68280 -22214 -68263
rect -22114 -68263 -22098 -68246
rect -21972 -68246 -21840 -68230
rect -21972 -68263 -21956 -68246
rect -22114 -68280 -22064 -68263
rect -22264 -68318 -22064 -68280
rect -22006 -68280 -21956 -68263
rect -21856 -68263 -21840 -68246
rect -21856 -68280 -21806 -68263
rect -22006 -68318 -21806 -68280
rect -23296 -68756 -23096 -68718
rect -23296 -68773 -23246 -68756
rect -23262 -68790 -23246 -68773
rect -23146 -68773 -23096 -68756
rect -23038 -68756 -22838 -68718
rect -23038 -68773 -22988 -68756
rect -23146 -68790 -23130 -68773
rect -23262 -68806 -23130 -68790
rect -23004 -68790 -22988 -68773
rect -22888 -68773 -22838 -68756
rect -22780 -68756 -22580 -68718
rect -22780 -68773 -22730 -68756
rect -22888 -68790 -22872 -68773
rect -23004 -68806 -22872 -68790
rect -22746 -68790 -22730 -68773
rect -22630 -68773 -22580 -68756
rect -22522 -68756 -22322 -68718
rect -22522 -68773 -22472 -68756
rect -22630 -68790 -22614 -68773
rect -22746 -68806 -22614 -68790
rect -22488 -68790 -22472 -68773
rect -22372 -68773 -22322 -68756
rect -22264 -68756 -22064 -68718
rect -22264 -68773 -22214 -68756
rect -22372 -68790 -22356 -68773
rect -22488 -68806 -22356 -68790
rect -22230 -68790 -22214 -68773
rect -22114 -68773 -22064 -68756
rect -22006 -68756 -21806 -68718
rect -22006 -68773 -21956 -68756
rect -22114 -68790 -22098 -68773
rect -22230 -68806 -22098 -68790
rect -21972 -68790 -21956 -68773
rect -21856 -68773 -21806 -68756
rect -21856 -68790 -21840 -68773
rect -21972 -68806 -21840 -68790
rect -15952 -67805 -15922 -67779
rect -19262 -68246 -19130 -68230
rect -19262 -68263 -19246 -68246
rect -19296 -68280 -19246 -68263
rect -19146 -68263 -19130 -68246
rect -19004 -68246 -18872 -68230
rect -19004 -68263 -18988 -68246
rect -19146 -68280 -19096 -68263
rect -19296 -68318 -19096 -68280
rect -19038 -68280 -18988 -68263
rect -18888 -68263 -18872 -68246
rect -18746 -68246 -18614 -68230
rect -18746 -68263 -18730 -68246
rect -18888 -68280 -18838 -68263
rect -19038 -68318 -18838 -68280
rect -18780 -68280 -18730 -68263
rect -18630 -68263 -18614 -68246
rect -18488 -68246 -18356 -68230
rect -18488 -68263 -18472 -68246
rect -18630 -68280 -18580 -68263
rect -18780 -68318 -18580 -68280
rect -18522 -68280 -18472 -68263
rect -18372 -68263 -18356 -68246
rect -18230 -68246 -18098 -68230
rect -18230 -68263 -18214 -68246
rect -18372 -68280 -18322 -68263
rect -18522 -68318 -18322 -68280
rect -18264 -68280 -18214 -68263
rect -18114 -68263 -18098 -68246
rect -17972 -68246 -17840 -68230
rect -17972 -68263 -17956 -68246
rect -18114 -68280 -18064 -68263
rect -18264 -68318 -18064 -68280
rect -18006 -68280 -17956 -68263
rect -17856 -68263 -17840 -68246
rect -17856 -68280 -17806 -68263
rect -18006 -68318 -17806 -68280
rect -19296 -68756 -19096 -68718
rect -19296 -68773 -19246 -68756
rect -19262 -68790 -19246 -68773
rect -19146 -68773 -19096 -68756
rect -19038 -68756 -18838 -68718
rect -19038 -68773 -18988 -68756
rect -19146 -68790 -19130 -68773
rect -19262 -68806 -19130 -68790
rect -19004 -68790 -18988 -68773
rect -18888 -68773 -18838 -68756
rect -18780 -68756 -18580 -68718
rect -18780 -68773 -18730 -68756
rect -18888 -68790 -18872 -68773
rect -19004 -68806 -18872 -68790
rect -18746 -68790 -18730 -68773
rect -18630 -68773 -18580 -68756
rect -18522 -68756 -18322 -68718
rect -18522 -68773 -18472 -68756
rect -18630 -68790 -18614 -68773
rect -18746 -68806 -18614 -68790
rect -18488 -68790 -18472 -68773
rect -18372 -68773 -18322 -68756
rect -18264 -68756 -18064 -68718
rect -18264 -68773 -18214 -68756
rect -18372 -68790 -18356 -68773
rect -18488 -68806 -18356 -68790
rect -18230 -68790 -18214 -68773
rect -18114 -68773 -18064 -68756
rect -18006 -68756 -17806 -68718
rect -18006 -68773 -17956 -68756
rect -18114 -68790 -18098 -68773
rect -18230 -68806 -18098 -68790
rect -17972 -68790 -17956 -68773
rect -17856 -68773 -17806 -68756
rect -17856 -68790 -17840 -68773
rect -17972 -68806 -17840 -68790
rect -11952 -67805 -11922 -67779
rect -15262 -68246 -15130 -68230
rect -15262 -68263 -15246 -68246
rect -15296 -68280 -15246 -68263
rect -15146 -68263 -15130 -68246
rect -15004 -68246 -14872 -68230
rect -15004 -68263 -14988 -68246
rect -15146 -68280 -15096 -68263
rect -15296 -68318 -15096 -68280
rect -15038 -68280 -14988 -68263
rect -14888 -68263 -14872 -68246
rect -14746 -68246 -14614 -68230
rect -14746 -68263 -14730 -68246
rect -14888 -68280 -14838 -68263
rect -15038 -68318 -14838 -68280
rect -14780 -68280 -14730 -68263
rect -14630 -68263 -14614 -68246
rect -14488 -68246 -14356 -68230
rect -14488 -68263 -14472 -68246
rect -14630 -68280 -14580 -68263
rect -14780 -68318 -14580 -68280
rect -14522 -68280 -14472 -68263
rect -14372 -68263 -14356 -68246
rect -14230 -68246 -14098 -68230
rect -14230 -68263 -14214 -68246
rect -14372 -68280 -14322 -68263
rect -14522 -68318 -14322 -68280
rect -14264 -68280 -14214 -68263
rect -14114 -68263 -14098 -68246
rect -13972 -68246 -13840 -68230
rect -13972 -68263 -13956 -68246
rect -14114 -68280 -14064 -68263
rect -14264 -68318 -14064 -68280
rect -14006 -68280 -13956 -68263
rect -13856 -68263 -13840 -68246
rect -13856 -68280 -13806 -68263
rect -14006 -68318 -13806 -68280
rect -15296 -68756 -15096 -68718
rect -15296 -68773 -15246 -68756
rect -15262 -68790 -15246 -68773
rect -15146 -68773 -15096 -68756
rect -15038 -68756 -14838 -68718
rect -15038 -68773 -14988 -68756
rect -15146 -68790 -15130 -68773
rect -15262 -68806 -15130 -68790
rect -15004 -68790 -14988 -68773
rect -14888 -68773 -14838 -68756
rect -14780 -68756 -14580 -68718
rect -14780 -68773 -14730 -68756
rect -14888 -68790 -14872 -68773
rect -15004 -68806 -14872 -68790
rect -14746 -68790 -14730 -68773
rect -14630 -68773 -14580 -68756
rect -14522 -68756 -14322 -68718
rect -14522 -68773 -14472 -68756
rect -14630 -68790 -14614 -68773
rect -14746 -68806 -14614 -68790
rect -14488 -68790 -14472 -68773
rect -14372 -68773 -14322 -68756
rect -14264 -68756 -14064 -68718
rect -14264 -68773 -14214 -68756
rect -14372 -68790 -14356 -68773
rect -14488 -68806 -14356 -68790
rect -14230 -68790 -14214 -68773
rect -14114 -68773 -14064 -68756
rect -14006 -68756 -13806 -68718
rect -14006 -68773 -13956 -68756
rect -14114 -68790 -14098 -68773
rect -14230 -68806 -14098 -68790
rect -13972 -68790 -13956 -68773
rect -13856 -68773 -13806 -68756
rect -13856 -68790 -13840 -68773
rect -13972 -68806 -13840 -68790
rect -7952 -67805 -7922 -67779
rect -11262 -68246 -11130 -68230
rect -11262 -68263 -11246 -68246
rect -11296 -68280 -11246 -68263
rect -11146 -68263 -11130 -68246
rect -11004 -68246 -10872 -68230
rect -11004 -68263 -10988 -68246
rect -11146 -68280 -11096 -68263
rect -11296 -68318 -11096 -68280
rect -11038 -68280 -10988 -68263
rect -10888 -68263 -10872 -68246
rect -10746 -68246 -10614 -68230
rect -10746 -68263 -10730 -68246
rect -10888 -68280 -10838 -68263
rect -11038 -68318 -10838 -68280
rect -10780 -68280 -10730 -68263
rect -10630 -68263 -10614 -68246
rect -10488 -68246 -10356 -68230
rect -10488 -68263 -10472 -68246
rect -10630 -68280 -10580 -68263
rect -10780 -68318 -10580 -68280
rect -10522 -68280 -10472 -68263
rect -10372 -68263 -10356 -68246
rect -10230 -68246 -10098 -68230
rect -10230 -68263 -10214 -68246
rect -10372 -68280 -10322 -68263
rect -10522 -68318 -10322 -68280
rect -10264 -68280 -10214 -68263
rect -10114 -68263 -10098 -68246
rect -9972 -68246 -9840 -68230
rect -9972 -68263 -9956 -68246
rect -10114 -68280 -10064 -68263
rect -10264 -68318 -10064 -68280
rect -10006 -68280 -9956 -68263
rect -9856 -68263 -9840 -68246
rect -9856 -68280 -9806 -68263
rect -10006 -68318 -9806 -68280
rect -11296 -68756 -11096 -68718
rect -11296 -68773 -11246 -68756
rect -11262 -68790 -11246 -68773
rect -11146 -68773 -11096 -68756
rect -11038 -68756 -10838 -68718
rect -11038 -68773 -10988 -68756
rect -11146 -68790 -11130 -68773
rect -11262 -68806 -11130 -68790
rect -11004 -68790 -10988 -68773
rect -10888 -68773 -10838 -68756
rect -10780 -68756 -10580 -68718
rect -10780 -68773 -10730 -68756
rect -10888 -68790 -10872 -68773
rect -11004 -68806 -10872 -68790
rect -10746 -68790 -10730 -68773
rect -10630 -68773 -10580 -68756
rect -10522 -68756 -10322 -68718
rect -10522 -68773 -10472 -68756
rect -10630 -68790 -10614 -68773
rect -10746 -68806 -10614 -68790
rect -10488 -68790 -10472 -68773
rect -10372 -68773 -10322 -68756
rect -10264 -68756 -10064 -68718
rect -10264 -68773 -10214 -68756
rect -10372 -68790 -10356 -68773
rect -10488 -68806 -10356 -68790
rect -10230 -68790 -10214 -68773
rect -10114 -68773 -10064 -68756
rect -10006 -68756 -9806 -68718
rect -10006 -68773 -9956 -68756
rect -10114 -68790 -10098 -68773
rect -10230 -68806 -10098 -68790
rect -9972 -68790 -9956 -68773
rect -9856 -68773 -9806 -68756
rect -9856 -68790 -9840 -68773
rect -9972 -68806 -9840 -68790
rect -3952 -67805 -3922 -67779
rect -7262 -68246 -7130 -68230
rect -7262 -68263 -7246 -68246
rect -7296 -68280 -7246 -68263
rect -7146 -68263 -7130 -68246
rect -7004 -68246 -6872 -68230
rect -7004 -68263 -6988 -68246
rect -7146 -68280 -7096 -68263
rect -7296 -68318 -7096 -68280
rect -7038 -68280 -6988 -68263
rect -6888 -68263 -6872 -68246
rect -6746 -68246 -6614 -68230
rect -6746 -68263 -6730 -68246
rect -6888 -68280 -6838 -68263
rect -7038 -68318 -6838 -68280
rect -6780 -68280 -6730 -68263
rect -6630 -68263 -6614 -68246
rect -6488 -68246 -6356 -68230
rect -6488 -68263 -6472 -68246
rect -6630 -68280 -6580 -68263
rect -6780 -68318 -6580 -68280
rect -6522 -68280 -6472 -68263
rect -6372 -68263 -6356 -68246
rect -6230 -68246 -6098 -68230
rect -6230 -68263 -6214 -68246
rect -6372 -68280 -6322 -68263
rect -6522 -68318 -6322 -68280
rect -6264 -68280 -6214 -68263
rect -6114 -68263 -6098 -68246
rect -5972 -68246 -5840 -68230
rect -5972 -68263 -5956 -68246
rect -6114 -68280 -6064 -68263
rect -6264 -68318 -6064 -68280
rect -6006 -68280 -5956 -68263
rect -5856 -68263 -5840 -68246
rect -5856 -68280 -5806 -68263
rect -6006 -68318 -5806 -68280
rect -7296 -68756 -7096 -68718
rect -7296 -68773 -7246 -68756
rect -7262 -68790 -7246 -68773
rect -7146 -68773 -7096 -68756
rect -7038 -68756 -6838 -68718
rect -7038 -68773 -6988 -68756
rect -7146 -68790 -7130 -68773
rect -7262 -68806 -7130 -68790
rect -7004 -68790 -6988 -68773
rect -6888 -68773 -6838 -68756
rect -6780 -68756 -6580 -68718
rect -6780 -68773 -6730 -68756
rect -6888 -68790 -6872 -68773
rect -7004 -68806 -6872 -68790
rect -6746 -68790 -6730 -68773
rect -6630 -68773 -6580 -68756
rect -6522 -68756 -6322 -68718
rect -6522 -68773 -6472 -68756
rect -6630 -68790 -6614 -68773
rect -6746 -68806 -6614 -68790
rect -6488 -68790 -6472 -68773
rect -6372 -68773 -6322 -68756
rect -6264 -68756 -6064 -68718
rect -6264 -68773 -6214 -68756
rect -6372 -68790 -6356 -68773
rect -6488 -68806 -6356 -68790
rect -6230 -68790 -6214 -68773
rect -6114 -68773 -6064 -68756
rect -6006 -68756 -5806 -68718
rect -6006 -68773 -5956 -68756
rect -6114 -68790 -6098 -68773
rect -6230 -68806 -6098 -68790
rect -5972 -68790 -5956 -68773
rect -5856 -68773 -5806 -68756
rect -5856 -68790 -5840 -68773
rect -5972 -68806 -5840 -68790
rect 48 -67805 78 -67779
rect -3262 -68246 -3130 -68230
rect -3262 -68263 -3246 -68246
rect -3296 -68280 -3246 -68263
rect -3146 -68263 -3130 -68246
rect -3004 -68246 -2872 -68230
rect -3004 -68263 -2988 -68246
rect -3146 -68280 -3096 -68263
rect -3296 -68318 -3096 -68280
rect -3038 -68280 -2988 -68263
rect -2888 -68263 -2872 -68246
rect -2746 -68246 -2614 -68230
rect -2746 -68263 -2730 -68246
rect -2888 -68280 -2838 -68263
rect -3038 -68318 -2838 -68280
rect -2780 -68280 -2730 -68263
rect -2630 -68263 -2614 -68246
rect -2488 -68246 -2356 -68230
rect -2488 -68263 -2472 -68246
rect -2630 -68280 -2580 -68263
rect -2780 -68318 -2580 -68280
rect -2522 -68280 -2472 -68263
rect -2372 -68263 -2356 -68246
rect -2230 -68246 -2098 -68230
rect -2230 -68263 -2214 -68246
rect -2372 -68280 -2322 -68263
rect -2522 -68318 -2322 -68280
rect -2264 -68280 -2214 -68263
rect -2114 -68263 -2098 -68246
rect -1972 -68246 -1840 -68230
rect -1972 -68263 -1956 -68246
rect -2114 -68280 -2064 -68263
rect -2264 -68318 -2064 -68280
rect -2006 -68280 -1956 -68263
rect -1856 -68263 -1840 -68246
rect -1856 -68280 -1806 -68263
rect -2006 -68318 -1806 -68280
rect -3296 -68756 -3096 -68718
rect -3296 -68773 -3246 -68756
rect -3262 -68790 -3246 -68773
rect -3146 -68773 -3096 -68756
rect -3038 -68756 -2838 -68718
rect -3038 -68773 -2988 -68756
rect -3146 -68790 -3130 -68773
rect -3262 -68806 -3130 -68790
rect -3004 -68790 -2988 -68773
rect -2888 -68773 -2838 -68756
rect -2780 -68756 -2580 -68718
rect -2780 -68773 -2730 -68756
rect -2888 -68790 -2872 -68773
rect -3004 -68806 -2872 -68790
rect -2746 -68790 -2730 -68773
rect -2630 -68773 -2580 -68756
rect -2522 -68756 -2322 -68718
rect -2522 -68773 -2472 -68756
rect -2630 -68790 -2614 -68773
rect -2746 -68806 -2614 -68790
rect -2488 -68790 -2472 -68773
rect -2372 -68773 -2322 -68756
rect -2264 -68756 -2064 -68718
rect -2264 -68773 -2214 -68756
rect -2372 -68790 -2356 -68773
rect -2488 -68806 -2356 -68790
rect -2230 -68790 -2214 -68773
rect -2114 -68773 -2064 -68756
rect -2006 -68756 -1806 -68718
rect -2006 -68773 -1956 -68756
rect -2114 -68790 -2098 -68773
rect -2230 -68806 -2098 -68790
rect -1972 -68790 -1956 -68773
rect -1856 -68773 -1806 -68756
rect -1856 -68790 -1840 -68773
rect -1972 -68806 -1840 -68790
rect 4048 -67805 4078 -67779
rect 738 -68246 870 -68230
rect 738 -68263 754 -68246
rect 704 -68280 754 -68263
rect 854 -68263 870 -68246
rect 996 -68246 1128 -68230
rect 996 -68263 1012 -68246
rect 854 -68280 904 -68263
rect 704 -68318 904 -68280
rect 962 -68280 1012 -68263
rect 1112 -68263 1128 -68246
rect 1254 -68246 1386 -68230
rect 1254 -68263 1270 -68246
rect 1112 -68280 1162 -68263
rect 962 -68318 1162 -68280
rect 1220 -68280 1270 -68263
rect 1370 -68263 1386 -68246
rect 1512 -68246 1644 -68230
rect 1512 -68263 1528 -68246
rect 1370 -68280 1420 -68263
rect 1220 -68318 1420 -68280
rect 1478 -68280 1528 -68263
rect 1628 -68263 1644 -68246
rect 1770 -68246 1902 -68230
rect 1770 -68263 1786 -68246
rect 1628 -68280 1678 -68263
rect 1478 -68318 1678 -68280
rect 1736 -68280 1786 -68263
rect 1886 -68263 1902 -68246
rect 2028 -68246 2160 -68230
rect 2028 -68263 2044 -68246
rect 1886 -68280 1936 -68263
rect 1736 -68318 1936 -68280
rect 1994 -68280 2044 -68263
rect 2144 -68263 2160 -68246
rect 2144 -68280 2194 -68263
rect 1994 -68318 2194 -68280
rect 704 -68756 904 -68718
rect 704 -68773 754 -68756
rect 738 -68790 754 -68773
rect 854 -68773 904 -68756
rect 962 -68756 1162 -68718
rect 962 -68773 1012 -68756
rect 854 -68790 870 -68773
rect 738 -68806 870 -68790
rect 996 -68790 1012 -68773
rect 1112 -68773 1162 -68756
rect 1220 -68756 1420 -68718
rect 1220 -68773 1270 -68756
rect 1112 -68790 1128 -68773
rect 996 -68806 1128 -68790
rect 1254 -68790 1270 -68773
rect 1370 -68773 1420 -68756
rect 1478 -68756 1678 -68718
rect 1478 -68773 1528 -68756
rect 1370 -68790 1386 -68773
rect 1254 -68806 1386 -68790
rect 1512 -68790 1528 -68773
rect 1628 -68773 1678 -68756
rect 1736 -68756 1936 -68718
rect 1736 -68773 1786 -68756
rect 1628 -68790 1644 -68773
rect 1512 -68806 1644 -68790
rect 1770 -68790 1786 -68773
rect 1886 -68773 1936 -68756
rect 1994 -68756 2194 -68718
rect 1994 -68773 2044 -68756
rect 1886 -68790 1902 -68773
rect 1770 -68806 1902 -68790
rect 2028 -68790 2044 -68773
rect 2144 -68773 2194 -68756
rect 2144 -68790 2160 -68773
rect 2028 -68806 2160 -68790
rect 4738 -68246 4870 -68230
rect 4738 -68263 4754 -68246
rect 4704 -68280 4754 -68263
rect 4854 -68263 4870 -68246
rect 4996 -68246 5128 -68230
rect 4996 -68263 5012 -68246
rect 4854 -68280 4904 -68263
rect 4704 -68318 4904 -68280
rect 4962 -68280 5012 -68263
rect 5112 -68263 5128 -68246
rect 5254 -68246 5386 -68230
rect 5254 -68263 5270 -68246
rect 5112 -68280 5162 -68263
rect 4962 -68318 5162 -68280
rect 5220 -68280 5270 -68263
rect 5370 -68263 5386 -68246
rect 5512 -68246 5644 -68230
rect 5512 -68263 5528 -68246
rect 5370 -68280 5420 -68263
rect 5220 -68318 5420 -68280
rect 5478 -68280 5528 -68263
rect 5628 -68263 5644 -68246
rect 5770 -68246 5902 -68230
rect 5770 -68263 5786 -68246
rect 5628 -68280 5678 -68263
rect 5478 -68318 5678 -68280
rect 5736 -68280 5786 -68263
rect 5886 -68263 5902 -68246
rect 6028 -68246 6160 -68230
rect 6028 -68263 6044 -68246
rect 5886 -68280 5936 -68263
rect 5736 -68318 5936 -68280
rect 5994 -68280 6044 -68263
rect 6144 -68263 6160 -68246
rect 6144 -68280 6194 -68263
rect 5994 -68318 6194 -68280
rect 4704 -68756 4904 -68718
rect 4704 -68773 4754 -68756
rect 4738 -68790 4754 -68773
rect 4854 -68773 4904 -68756
rect 4962 -68756 5162 -68718
rect 4962 -68773 5012 -68756
rect 4854 -68790 4870 -68773
rect 4738 -68806 4870 -68790
rect 4996 -68790 5012 -68773
rect 5112 -68773 5162 -68756
rect 5220 -68756 5420 -68718
rect 5220 -68773 5270 -68756
rect 5112 -68790 5128 -68773
rect 4996 -68806 5128 -68790
rect 5254 -68790 5270 -68773
rect 5370 -68773 5420 -68756
rect 5478 -68756 5678 -68718
rect 5478 -68773 5528 -68756
rect 5370 -68790 5386 -68773
rect 5254 -68806 5386 -68790
rect 5512 -68790 5528 -68773
rect 5628 -68773 5678 -68756
rect 5736 -68756 5936 -68718
rect 5736 -68773 5786 -68756
rect 5628 -68790 5644 -68773
rect 5512 -68806 5644 -68790
rect 5770 -68790 5786 -68773
rect 5886 -68773 5936 -68756
rect 5994 -68756 6194 -68718
rect 5994 -68773 6044 -68756
rect 5886 -68790 5902 -68773
rect 5770 -68806 5902 -68790
rect 6028 -68790 6044 -68773
rect 6144 -68773 6194 -68756
rect 6144 -68790 6160 -68773
rect 6028 -68806 6160 -68790
rect -27262 -71406 -27130 -71390
rect -27262 -71423 -27246 -71406
rect -27296 -71440 -27246 -71423
rect -27146 -71423 -27130 -71406
rect -27004 -71406 -26872 -71390
rect -27004 -71423 -26988 -71406
rect -27146 -71440 -27096 -71423
rect -27296 -71478 -27096 -71440
rect -27038 -71440 -26988 -71423
rect -26888 -71423 -26872 -71406
rect -26746 -71406 -26614 -71390
rect -26746 -71423 -26730 -71406
rect -26888 -71440 -26838 -71423
rect -27038 -71478 -26838 -71440
rect -26780 -71440 -26730 -71423
rect -26630 -71423 -26614 -71406
rect -26488 -71406 -26356 -71390
rect -26488 -71423 -26472 -71406
rect -26630 -71440 -26580 -71423
rect -26780 -71478 -26580 -71440
rect -26522 -71440 -26472 -71423
rect -26372 -71423 -26356 -71406
rect -26230 -71406 -26098 -71390
rect -26230 -71423 -26214 -71406
rect -26372 -71440 -26322 -71423
rect -26522 -71478 -26322 -71440
rect -26264 -71440 -26214 -71423
rect -26114 -71423 -26098 -71406
rect -25972 -71406 -25840 -71390
rect -25972 -71423 -25956 -71406
rect -26114 -71440 -26064 -71423
rect -26264 -71478 -26064 -71440
rect -26006 -71440 -25956 -71423
rect -25856 -71423 -25840 -71406
rect -25856 -71440 -25806 -71423
rect -26006 -71478 -25806 -71440
rect -27296 -71916 -27096 -71878
rect -27296 -71933 -27246 -71916
rect -27262 -71950 -27246 -71933
rect -27146 -71933 -27096 -71916
rect -27038 -71916 -26838 -71878
rect -27038 -71933 -26988 -71916
rect -27146 -71950 -27130 -71933
rect -27262 -71966 -27130 -71950
rect -27004 -71950 -26988 -71933
rect -26888 -71933 -26838 -71916
rect -26780 -71916 -26580 -71878
rect -26780 -71933 -26730 -71916
rect -26888 -71950 -26872 -71933
rect -27004 -71966 -26872 -71950
rect -26746 -71950 -26730 -71933
rect -26630 -71933 -26580 -71916
rect -26522 -71916 -26322 -71878
rect -26522 -71933 -26472 -71916
rect -26630 -71950 -26614 -71933
rect -26746 -71966 -26614 -71950
rect -26488 -71950 -26472 -71933
rect -26372 -71933 -26322 -71916
rect -26264 -71916 -26064 -71878
rect -26264 -71933 -26214 -71916
rect -26372 -71950 -26356 -71933
rect -26488 -71966 -26356 -71950
rect -26230 -71950 -26214 -71933
rect -26114 -71933 -26064 -71916
rect -26006 -71916 -25806 -71878
rect -26006 -71933 -25956 -71916
rect -26114 -71950 -26098 -71933
rect -26230 -71966 -26098 -71950
rect -25972 -71950 -25956 -71933
rect -25856 -71933 -25806 -71916
rect -25856 -71950 -25840 -71933
rect -25972 -71966 -25840 -71950
rect -27952 -72417 -27922 -72391
rect -23262 -71406 -23130 -71390
rect -23262 -71423 -23246 -71406
rect -23296 -71440 -23246 -71423
rect -23146 -71423 -23130 -71406
rect -23004 -71406 -22872 -71390
rect -23004 -71423 -22988 -71406
rect -23146 -71440 -23096 -71423
rect -23296 -71478 -23096 -71440
rect -23038 -71440 -22988 -71423
rect -22888 -71423 -22872 -71406
rect -22746 -71406 -22614 -71390
rect -22746 -71423 -22730 -71406
rect -22888 -71440 -22838 -71423
rect -23038 -71478 -22838 -71440
rect -22780 -71440 -22730 -71423
rect -22630 -71423 -22614 -71406
rect -22488 -71406 -22356 -71390
rect -22488 -71423 -22472 -71406
rect -22630 -71440 -22580 -71423
rect -22780 -71478 -22580 -71440
rect -22522 -71440 -22472 -71423
rect -22372 -71423 -22356 -71406
rect -22230 -71406 -22098 -71390
rect -22230 -71423 -22214 -71406
rect -22372 -71440 -22322 -71423
rect -22522 -71478 -22322 -71440
rect -22264 -71440 -22214 -71423
rect -22114 -71423 -22098 -71406
rect -21972 -71406 -21840 -71390
rect -21972 -71423 -21956 -71406
rect -22114 -71440 -22064 -71423
rect -22264 -71478 -22064 -71440
rect -22006 -71440 -21956 -71423
rect -21856 -71423 -21840 -71406
rect -21856 -71440 -21806 -71423
rect -22006 -71478 -21806 -71440
rect -23296 -71916 -23096 -71878
rect -23296 -71933 -23246 -71916
rect -23262 -71950 -23246 -71933
rect -23146 -71933 -23096 -71916
rect -23038 -71916 -22838 -71878
rect -23038 -71933 -22988 -71916
rect -23146 -71950 -23130 -71933
rect -23262 -71966 -23130 -71950
rect -23004 -71950 -22988 -71933
rect -22888 -71933 -22838 -71916
rect -22780 -71916 -22580 -71878
rect -22780 -71933 -22730 -71916
rect -22888 -71950 -22872 -71933
rect -23004 -71966 -22872 -71950
rect -22746 -71950 -22730 -71933
rect -22630 -71933 -22580 -71916
rect -22522 -71916 -22322 -71878
rect -22522 -71933 -22472 -71916
rect -22630 -71950 -22614 -71933
rect -22746 -71966 -22614 -71950
rect -22488 -71950 -22472 -71933
rect -22372 -71933 -22322 -71916
rect -22264 -71916 -22064 -71878
rect -22264 -71933 -22214 -71916
rect -22372 -71950 -22356 -71933
rect -22488 -71966 -22356 -71950
rect -22230 -71950 -22214 -71933
rect -22114 -71933 -22064 -71916
rect -22006 -71916 -21806 -71878
rect -22006 -71933 -21956 -71916
rect -22114 -71950 -22098 -71933
rect -22230 -71966 -22098 -71950
rect -21972 -71950 -21956 -71933
rect -21856 -71933 -21806 -71916
rect -21856 -71950 -21840 -71933
rect -21972 -71966 -21840 -71950
rect -23952 -72417 -23922 -72391
rect -19262 -71406 -19130 -71390
rect -19262 -71423 -19246 -71406
rect -19296 -71440 -19246 -71423
rect -19146 -71423 -19130 -71406
rect -19004 -71406 -18872 -71390
rect -19004 -71423 -18988 -71406
rect -19146 -71440 -19096 -71423
rect -19296 -71478 -19096 -71440
rect -19038 -71440 -18988 -71423
rect -18888 -71423 -18872 -71406
rect -18746 -71406 -18614 -71390
rect -18746 -71423 -18730 -71406
rect -18888 -71440 -18838 -71423
rect -19038 -71478 -18838 -71440
rect -18780 -71440 -18730 -71423
rect -18630 -71423 -18614 -71406
rect -18488 -71406 -18356 -71390
rect -18488 -71423 -18472 -71406
rect -18630 -71440 -18580 -71423
rect -18780 -71478 -18580 -71440
rect -18522 -71440 -18472 -71423
rect -18372 -71423 -18356 -71406
rect -18230 -71406 -18098 -71390
rect -18230 -71423 -18214 -71406
rect -18372 -71440 -18322 -71423
rect -18522 -71478 -18322 -71440
rect -18264 -71440 -18214 -71423
rect -18114 -71423 -18098 -71406
rect -17972 -71406 -17840 -71390
rect -17972 -71423 -17956 -71406
rect -18114 -71440 -18064 -71423
rect -18264 -71478 -18064 -71440
rect -18006 -71440 -17956 -71423
rect -17856 -71423 -17840 -71406
rect -17856 -71440 -17806 -71423
rect -18006 -71478 -17806 -71440
rect -19296 -71916 -19096 -71878
rect -19296 -71933 -19246 -71916
rect -19262 -71950 -19246 -71933
rect -19146 -71933 -19096 -71916
rect -19038 -71916 -18838 -71878
rect -19038 -71933 -18988 -71916
rect -19146 -71950 -19130 -71933
rect -19262 -71966 -19130 -71950
rect -19004 -71950 -18988 -71933
rect -18888 -71933 -18838 -71916
rect -18780 -71916 -18580 -71878
rect -18780 -71933 -18730 -71916
rect -18888 -71950 -18872 -71933
rect -19004 -71966 -18872 -71950
rect -18746 -71950 -18730 -71933
rect -18630 -71933 -18580 -71916
rect -18522 -71916 -18322 -71878
rect -18522 -71933 -18472 -71916
rect -18630 -71950 -18614 -71933
rect -18746 -71966 -18614 -71950
rect -18488 -71950 -18472 -71933
rect -18372 -71933 -18322 -71916
rect -18264 -71916 -18064 -71878
rect -18264 -71933 -18214 -71916
rect -18372 -71950 -18356 -71933
rect -18488 -71966 -18356 -71950
rect -18230 -71950 -18214 -71933
rect -18114 -71933 -18064 -71916
rect -18006 -71916 -17806 -71878
rect -18006 -71933 -17956 -71916
rect -18114 -71950 -18098 -71933
rect -18230 -71966 -18098 -71950
rect -17972 -71950 -17956 -71933
rect -17856 -71933 -17806 -71916
rect -17856 -71950 -17840 -71933
rect -17972 -71966 -17840 -71950
rect -19952 -72417 -19922 -72391
rect -15262 -71406 -15130 -71390
rect -15262 -71423 -15246 -71406
rect -15296 -71440 -15246 -71423
rect -15146 -71423 -15130 -71406
rect -15004 -71406 -14872 -71390
rect -15004 -71423 -14988 -71406
rect -15146 -71440 -15096 -71423
rect -15296 -71478 -15096 -71440
rect -15038 -71440 -14988 -71423
rect -14888 -71423 -14872 -71406
rect -14746 -71406 -14614 -71390
rect -14746 -71423 -14730 -71406
rect -14888 -71440 -14838 -71423
rect -15038 -71478 -14838 -71440
rect -14780 -71440 -14730 -71423
rect -14630 -71423 -14614 -71406
rect -14488 -71406 -14356 -71390
rect -14488 -71423 -14472 -71406
rect -14630 -71440 -14580 -71423
rect -14780 -71478 -14580 -71440
rect -14522 -71440 -14472 -71423
rect -14372 -71423 -14356 -71406
rect -14230 -71406 -14098 -71390
rect -14230 -71423 -14214 -71406
rect -14372 -71440 -14322 -71423
rect -14522 -71478 -14322 -71440
rect -14264 -71440 -14214 -71423
rect -14114 -71423 -14098 -71406
rect -13972 -71406 -13840 -71390
rect -13972 -71423 -13956 -71406
rect -14114 -71440 -14064 -71423
rect -14264 -71478 -14064 -71440
rect -14006 -71440 -13956 -71423
rect -13856 -71423 -13840 -71406
rect -13856 -71440 -13806 -71423
rect -14006 -71478 -13806 -71440
rect -15296 -71916 -15096 -71878
rect -15296 -71933 -15246 -71916
rect -15262 -71950 -15246 -71933
rect -15146 -71933 -15096 -71916
rect -15038 -71916 -14838 -71878
rect -15038 -71933 -14988 -71916
rect -15146 -71950 -15130 -71933
rect -15262 -71966 -15130 -71950
rect -15004 -71950 -14988 -71933
rect -14888 -71933 -14838 -71916
rect -14780 -71916 -14580 -71878
rect -14780 -71933 -14730 -71916
rect -14888 -71950 -14872 -71933
rect -15004 -71966 -14872 -71950
rect -14746 -71950 -14730 -71933
rect -14630 -71933 -14580 -71916
rect -14522 -71916 -14322 -71878
rect -14522 -71933 -14472 -71916
rect -14630 -71950 -14614 -71933
rect -14746 -71966 -14614 -71950
rect -14488 -71950 -14472 -71933
rect -14372 -71933 -14322 -71916
rect -14264 -71916 -14064 -71878
rect -14264 -71933 -14214 -71916
rect -14372 -71950 -14356 -71933
rect -14488 -71966 -14356 -71950
rect -14230 -71950 -14214 -71933
rect -14114 -71933 -14064 -71916
rect -14006 -71916 -13806 -71878
rect -14006 -71933 -13956 -71916
rect -14114 -71950 -14098 -71933
rect -14230 -71966 -14098 -71950
rect -13972 -71950 -13956 -71933
rect -13856 -71933 -13806 -71916
rect -13856 -71950 -13840 -71933
rect -13972 -71966 -13840 -71950
rect -15952 -72417 -15922 -72391
rect -11262 -71406 -11130 -71390
rect -11262 -71423 -11246 -71406
rect -11296 -71440 -11246 -71423
rect -11146 -71423 -11130 -71406
rect -11004 -71406 -10872 -71390
rect -11004 -71423 -10988 -71406
rect -11146 -71440 -11096 -71423
rect -11296 -71478 -11096 -71440
rect -11038 -71440 -10988 -71423
rect -10888 -71423 -10872 -71406
rect -10746 -71406 -10614 -71390
rect -10746 -71423 -10730 -71406
rect -10888 -71440 -10838 -71423
rect -11038 -71478 -10838 -71440
rect -10780 -71440 -10730 -71423
rect -10630 -71423 -10614 -71406
rect -10488 -71406 -10356 -71390
rect -10488 -71423 -10472 -71406
rect -10630 -71440 -10580 -71423
rect -10780 -71478 -10580 -71440
rect -10522 -71440 -10472 -71423
rect -10372 -71423 -10356 -71406
rect -10230 -71406 -10098 -71390
rect -10230 -71423 -10214 -71406
rect -10372 -71440 -10322 -71423
rect -10522 -71478 -10322 -71440
rect -10264 -71440 -10214 -71423
rect -10114 -71423 -10098 -71406
rect -9972 -71406 -9840 -71390
rect -9972 -71423 -9956 -71406
rect -10114 -71440 -10064 -71423
rect -10264 -71478 -10064 -71440
rect -10006 -71440 -9956 -71423
rect -9856 -71423 -9840 -71406
rect -9856 -71440 -9806 -71423
rect -10006 -71478 -9806 -71440
rect -11296 -71916 -11096 -71878
rect -11296 -71933 -11246 -71916
rect -11262 -71950 -11246 -71933
rect -11146 -71933 -11096 -71916
rect -11038 -71916 -10838 -71878
rect -11038 -71933 -10988 -71916
rect -11146 -71950 -11130 -71933
rect -11262 -71966 -11130 -71950
rect -11004 -71950 -10988 -71933
rect -10888 -71933 -10838 -71916
rect -10780 -71916 -10580 -71878
rect -10780 -71933 -10730 -71916
rect -10888 -71950 -10872 -71933
rect -11004 -71966 -10872 -71950
rect -10746 -71950 -10730 -71933
rect -10630 -71933 -10580 -71916
rect -10522 -71916 -10322 -71878
rect -10522 -71933 -10472 -71916
rect -10630 -71950 -10614 -71933
rect -10746 -71966 -10614 -71950
rect -10488 -71950 -10472 -71933
rect -10372 -71933 -10322 -71916
rect -10264 -71916 -10064 -71878
rect -10264 -71933 -10214 -71916
rect -10372 -71950 -10356 -71933
rect -10488 -71966 -10356 -71950
rect -10230 -71950 -10214 -71933
rect -10114 -71933 -10064 -71916
rect -10006 -71916 -9806 -71878
rect -10006 -71933 -9956 -71916
rect -10114 -71950 -10098 -71933
rect -10230 -71966 -10098 -71950
rect -9972 -71950 -9956 -71933
rect -9856 -71933 -9806 -71916
rect -9856 -71950 -9840 -71933
rect -9972 -71966 -9840 -71950
rect -11952 -72417 -11922 -72391
rect -7262 -71406 -7130 -71390
rect -7262 -71423 -7246 -71406
rect -7296 -71440 -7246 -71423
rect -7146 -71423 -7130 -71406
rect -7004 -71406 -6872 -71390
rect -7004 -71423 -6988 -71406
rect -7146 -71440 -7096 -71423
rect -7296 -71478 -7096 -71440
rect -7038 -71440 -6988 -71423
rect -6888 -71423 -6872 -71406
rect -6746 -71406 -6614 -71390
rect -6746 -71423 -6730 -71406
rect -6888 -71440 -6838 -71423
rect -7038 -71478 -6838 -71440
rect -6780 -71440 -6730 -71423
rect -6630 -71423 -6614 -71406
rect -6488 -71406 -6356 -71390
rect -6488 -71423 -6472 -71406
rect -6630 -71440 -6580 -71423
rect -6780 -71478 -6580 -71440
rect -6522 -71440 -6472 -71423
rect -6372 -71423 -6356 -71406
rect -6230 -71406 -6098 -71390
rect -6230 -71423 -6214 -71406
rect -6372 -71440 -6322 -71423
rect -6522 -71478 -6322 -71440
rect -6264 -71440 -6214 -71423
rect -6114 -71423 -6098 -71406
rect -5972 -71406 -5840 -71390
rect -5972 -71423 -5956 -71406
rect -6114 -71440 -6064 -71423
rect -6264 -71478 -6064 -71440
rect -6006 -71440 -5956 -71423
rect -5856 -71423 -5840 -71406
rect -5856 -71440 -5806 -71423
rect -6006 -71478 -5806 -71440
rect -7296 -71916 -7096 -71878
rect -7296 -71933 -7246 -71916
rect -7262 -71950 -7246 -71933
rect -7146 -71933 -7096 -71916
rect -7038 -71916 -6838 -71878
rect -7038 -71933 -6988 -71916
rect -7146 -71950 -7130 -71933
rect -7262 -71966 -7130 -71950
rect -7004 -71950 -6988 -71933
rect -6888 -71933 -6838 -71916
rect -6780 -71916 -6580 -71878
rect -6780 -71933 -6730 -71916
rect -6888 -71950 -6872 -71933
rect -7004 -71966 -6872 -71950
rect -6746 -71950 -6730 -71933
rect -6630 -71933 -6580 -71916
rect -6522 -71916 -6322 -71878
rect -6522 -71933 -6472 -71916
rect -6630 -71950 -6614 -71933
rect -6746 -71966 -6614 -71950
rect -6488 -71950 -6472 -71933
rect -6372 -71933 -6322 -71916
rect -6264 -71916 -6064 -71878
rect -6264 -71933 -6214 -71916
rect -6372 -71950 -6356 -71933
rect -6488 -71966 -6356 -71950
rect -6230 -71950 -6214 -71933
rect -6114 -71933 -6064 -71916
rect -6006 -71916 -5806 -71878
rect -6006 -71933 -5956 -71916
rect -6114 -71950 -6098 -71933
rect -6230 -71966 -6098 -71950
rect -5972 -71950 -5956 -71933
rect -5856 -71933 -5806 -71916
rect -5856 -71950 -5840 -71933
rect -5972 -71966 -5840 -71950
rect -7952 -72417 -7922 -72391
rect -3262 -71406 -3130 -71390
rect -3262 -71423 -3246 -71406
rect -3296 -71440 -3246 -71423
rect -3146 -71423 -3130 -71406
rect -3004 -71406 -2872 -71390
rect -3004 -71423 -2988 -71406
rect -3146 -71440 -3096 -71423
rect -3296 -71478 -3096 -71440
rect -3038 -71440 -2988 -71423
rect -2888 -71423 -2872 -71406
rect -2746 -71406 -2614 -71390
rect -2746 -71423 -2730 -71406
rect -2888 -71440 -2838 -71423
rect -3038 -71478 -2838 -71440
rect -2780 -71440 -2730 -71423
rect -2630 -71423 -2614 -71406
rect -2488 -71406 -2356 -71390
rect -2488 -71423 -2472 -71406
rect -2630 -71440 -2580 -71423
rect -2780 -71478 -2580 -71440
rect -2522 -71440 -2472 -71423
rect -2372 -71423 -2356 -71406
rect -2230 -71406 -2098 -71390
rect -2230 -71423 -2214 -71406
rect -2372 -71440 -2322 -71423
rect -2522 -71478 -2322 -71440
rect -2264 -71440 -2214 -71423
rect -2114 -71423 -2098 -71406
rect -1972 -71406 -1840 -71390
rect -1972 -71423 -1956 -71406
rect -2114 -71440 -2064 -71423
rect -2264 -71478 -2064 -71440
rect -2006 -71440 -1956 -71423
rect -1856 -71423 -1840 -71406
rect -1856 -71440 -1806 -71423
rect -2006 -71478 -1806 -71440
rect -3296 -71916 -3096 -71878
rect -3296 -71933 -3246 -71916
rect -3262 -71950 -3246 -71933
rect -3146 -71933 -3096 -71916
rect -3038 -71916 -2838 -71878
rect -3038 -71933 -2988 -71916
rect -3146 -71950 -3130 -71933
rect -3262 -71966 -3130 -71950
rect -3004 -71950 -2988 -71933
rect -2888 -71933 -2838 -71916
rect -2780 -71916 -2580 -71878
rect -2780 -71933 -2730 -71916
rect -2888 -71950 -2872 -71933
rect -3004 -71966 -2872 -71950
rect -2746 -71950 -2730 -71933
rect -2630 -71933 -2580 -71916
rect -2522 -71916 -2322 -71878
rect -2522 -71933 -2472 -71916
rect -2630 -71950 -2614 -71933
rect -2746 -71966 -2614 -71950
rect -2488 -71950 -2472 -71933
rect -2372 -71933 -2322 -71916
rect -2264 -71916 -2064 -71878
rect -2264 -71933 -2214 -71916
rect -2372 -71950 -2356 -71933
rect -2488 -71966 -2356 -71950
rect -2230 -71950 -2214 -71933
rect -2114 -71933 -2064 -71916
rect -2006 -71916 -1806 -71878
rect -2006 -71933 -1956 -71916
rect -2114 -71950 -2098 -71933
rect -2230 -71966 -2098 -71950
rect -1972 -71950 -1956 -71933
rect -1856 -71933 -1806 -71916
rect -1856 -71950 -1840 -71933
rect -1972 -71966 -1840 -71950
rect -3952 -72417 -3922 -72391
rect 738 -71406 870 -71390
rect 738 -71423 754 -71406
rect 704 -71440 754 -71423
rect 854 -71423 870 -71406
rect 996 -71406 1128 -71390
rect 996 -71423 1012 -71406
rect 854 -71440 904 -71423
rect 704 -71478 904 -71440
rect 962 -71440 1012 -71423
rect 1112 -71423 1128 -71406
rect 1254 -71406 1386 -71390
rect 1254 -71423 1270 -71406
rect 1112 -71440 1162 -71423
rect 962 -71478 1162 -71440
rect 1220 -71440 1270 -71423
rect 1370 -71423 1386 -71406
rect 1512 -71406 1644 -71390
rect 1512 -71423 1528 -71406
rect 1370 -71440 1420 -71423
rect 1220 -71478 1420 -71440
rect 1478 -71440 1528 -71423
rect 1628 -71423 1644 -71406
rect 1770 -71406 1902 -71390
rect 1770 -71423 1786 -71406
rect 1628 -71440 1678 -71423
rect 1478 -71478 1678 -71440
rect 1736 -71440 1786 -71423
rect 1886 -71423 1902 -71406
rect 2028 -71406 2160 -71390
rect 2028 -71423 2044 -71406
rect 1886 -71440 1936 -71423
rect 1736 -71478 1936 -71440
rect 1994 -71440 2044 -71423
rect 2144 -71423 2160 -71406
rect 2144 -71440 2194 -71423
rect 1994 -71478 2194 -71440
rect 704 -71916 904 -71878
rect 704 -71933 754 -71916
rect 738 -71950 754 -71933
rect 854 -71933 904 -71916
rect 962 -71916 1162 -71878
rect 962 -71933 1012 -71916
rect 854 -71950 870 -71933
rect 738 -71966 870 -71950
rect 996 -71950 1012 -71933
rect 1112 -71933 1162 -71916
rect 1220 -71916 1420 -71878
rect 1220 -71933 1270 -71916
rect 1112 -71950 1128 -71933
rect 996 -71966 1128 -71950
rect 1254 -71950 1270 -71933
rect 1370 -71933 1420 -71916
rect 1478 -71916 1678 -71878
rect 1478 -71933 1528 -71916
rect 1370 -71950 1386 -71933
rect 1254 -71966 1386 -71950
rect 1512 -71950 1528 -71933
rect 1628 -71933 1678 -71916
rect 1736 -71916 1936 -71878
rect 1736 -71933 1786 -71916
rect 1628 -71950 1644 -71933
rect 1512 -71966 1644 -71950
rect 1770 -71950 1786 -71933
rect 1886 -71933 1936 -71916
rect 1994 -71916 2194 -71878
rect 1994 -71933 2044 -71916
rect 1886 -71950 1902 -71933
rect 1770 -71966 1902 -71950
rect 2028 -71950 2044 -71933
rect 2144 -71933 2194 -71916
rect 2144 -71950 2160 -71933
rect 2028 -71966 2160 -71950
rect 48 -72417 78 -72391
rect 4738 -71406 4870 -71390
rect 4738 -71423 4754 -71406
rect 4704 -71440 4754 -71423
rect 4854 -71423 4870 -71406
rect 4996 -71406 5128 -71390
rect 4996 -71423 5012 -71406
rect 4854 -71440 4904 -71423
rect 4704 -71478 4904 -71440
rect 4962 -71440 5012 -71423
rect 5112 -71423 5128 -71406
rect 5254 -71406 5386 -71390
rect 5254 -71423 5270 -71406
rect 5112 -71440 5162 -71423
rect 4962 -71478 5162 -71440
rect 5220 -71440 5270 -71423
rect 5370 -71423 5386 -71406
rect 5512 -71406 5644 -71390
rect 5512 -71423 5528 -71406
rect 5370 -71440 5420 -71423
rect 5220 -71478 5420 -71440
rect 5478 -71440 5528 -71423
rect 5628 -71423 5644 -71406
rect 5770 -71406 5902 -71390
rect 5770 -71423 5786 -71406
rect 5628 -71440 5678 -71423
rect 5478 -71478 5678 -71440
rect 5736 -71440 5786 -71423
rect 5886 -71423 5902 -71406
rect 6028 -71406 6160 -71390
rect 6028 -71423 6044 -71406
rect 5886 -71440 5936 -71423
rect 5736 -71478 5936 -71440
rect 5994 -71440 6044 -71423
rect 6144 -71423 6160 -71406
rect 6144 -71440 6194 -71423
rect 5994 -71478 6194 -71440
rect 4704 -71916 4904 -71878
rect 4704 -71933 4754 -71916
rect 4738 -71950 4754 -71933
rect 4854 -71933 4904 -71916
rect 4962 -71916 5162 -71878
rect 4962 -71933 5012 -71916
rect 4854 -71950 4870 -71933
rect 4738 -71966 4870 -71950
rect 4996 -71950 5012 -71933
rect 5112 -71933 5162 -71916
rect 5220 -71916 5420 -71878
rect 5220 -71933 5270 -71916
rect 5112 -71950 5128 -71933
rect 4996 -71966 5128 -71950
rect 5254 -71950 5270 -71933
rect 5370 -71933 5420 -71916
rect 5478 -71916 5678 -71878
rect 5478 -71933 5528 -71916
rect 5370 -71950 5386 -71933
rect 5254 -71966 5386 -71950
rect 5512 -71950 5528 -71933
rect 5628 -71933 5678 -71916
rect 5736 -71916 5936 -71878
rect 5736 -71933 5786 -71916
rect 5628 -71950 5644 -71933
rect 5512 -71966 5644 -71950
rect 5770 -71950 5786 -71933
rect 5886 -71933 5936 -71916
rect 5994 -71916 6194 -71878
rect 5994 -71933 6044 -71916
rect 5886 -71950 5902 -71933
rect 5770 -71966 5902 -71950
rect 6028 -71950 6044 -71933
rect 6144 -71933 6194 -71916
rect 6144 -71950 6160 -71933
rect 6028 -71966 6160 -71950
rect 4048 -72417 4078 -72391
rect -27952 -72569 -27922 -72547
rect -23952 -72569 -23922 -72547
rect -19952 -72569 -19922 -72547
rect -15952 -72569 -15922 -72547
rect -11952 -72569 -11922 -72547
rect -7952 -72569 -7922 -72547
rect -3952 -72569 -3922 -72547
rect 48 -72569 78 -72547
rect 4048 -72569 4078 -72547
rect -28008 -72585 -27922 -72569
rect -28008 -72619 -27992 -72585
rect -27958 -72619 -27922 -72585
rect -28008 -72635 -27922 -72619
rect -24008 -72585 -23922 -72569
rect -24008 -72619 -23992 -72585
rect -23958 -72619 -23922 -72585
rect -24008 -72635 -23922 -72619
rect -20008 -72585 -19922 -72569
rect -20008 -72619 -19992 -72585
rect -19958 -72619 -19922 -72585
rect -20008 -72635 -19922 -72619
rect -16008 -72585 -15922 -72569
rect -16008 -72619 -15992 -72585
rect -15958 -72619 -15922 -72585
rect -16008 -72635 -15922 -72619
rect -12008 -72585 -11922 -72569
rect -12008 -72619 -11992 -72585
rect -11958 -72619 -11922 -72585
rect -12008 -72635 -11922 -72619
rect -8008 -72585 -7922 -72569
rect -8008 -72619 -7992 -72585
rect -7958 -72619 -7922 -72585
rect -8008 -72635 -7922 -72619
rect -4008 -72585 -3922 -72569
rect -4008 -72619 -3992 -72585
rect -3958 -72619 -3922 -72585
rect -4008 -72635 -3922 -72619
rect -8 -72585 78 -72569
rect -8 -72619 8 -72585
rect 42 -72619 78 -72585
rect -8 -72635 78 -72619
rect 3992 -72585 4078 -72569
rect 3992 -72619 4008 -72585
rect 4042 -72619 4078 -72585
rect 3992 -72635 4078 -72619
rect -27952 -72667 -27922 -72635
rect -23952 -72667 -23922 -72635
rect -27952 -72893 -27922 -72867
rect -27257 -73230 -27125 -73214
rect -27257 -73247 -27241 -73230
rect -27291 -73264 -27241 -73247
rect -27141 -73247 -27125 -73230
rect -26999 -73230 -26867 -73214
rect -26999 -73247 -26983 -73230
rect -27141 -73264 -27091 -73247
rect -27291 -73311 -27091 -73264
rect -27033 -73264 -26983 -73247
rect -26883 -73247 -26867 -73230
rect -26741 -73230 -26609 -73214
rect -26741 -73247 -26725 -73230
rect -26883 -73264 -26833 -73247
rect -27033 -73311 -26833 -73264
rect -26775 -73264 -26725 -73247
rect -26625 -73247 -26609 -73230
rect -26483 -73230 -26351 -73214
rect -26483 -73247 -26467 -73230
rect -26625 -73264 -26575 -73247
rect -26775 -73311 -26575 -73264
rect -26517 -73264 -26467 -73247
rect -26367 -73247 -26351 -73230
rect -26225 -73230 -26093 -73214
rect -26225 -73247 -26209 -73230
rect -26367 -73264 -26317 -73247
rect -26517 -73311 -26317 -73264
rect -26259 -73264 -26209 -73247
rect -26109 -73247 -26093 -73230
rect -25967 -73230 -25835 -73214
rect -25967 -73247 -25951 -73230
rect -26109 -73264 -26059 -73247
rect -26259 -73311 -26059 -73264
rect -26001 -73264 -25951 -73247
rect -25851 -73247 -25835 -73230
rect -25851 -73264 -25801 -73247
rect -26001 -73311 -25801 -73264
rect -27291 -73758 -27091 -73711
rect -27291 -73775 -27241 -73758
rect -27257 -73792 -27241 -73775
rect -27141 -73775 -27091 -73758
rect -27033 -73758 -26833 -73711
rect -27033 -73775 -26983 -73758
rect -27141 -73792 -27125 -73775
rect -27257 -73808 -27125 -73792
rect -26999 -73792 -26983 -73775
rect -26883 -73775 -26833 -73758
rect -26775 -73758 -26575 -73711
rect -26775 -73775 -26725 -73758
rect -26883 -73792 -26867 -73775
rect -26999 -73808 -26867 -73792
rect -26741 -73792 -26725 -73775
rect -26625 -73775 -26575 -73758
rect -26517 -73758 -26317 -73711
rect -26517 -73775 -26467 -73758
rect -26625 -73792 -26609 -73775
rect -26741 -73808 -26609 -73792
rect -26483 -73792 -26467 -73775
rect -26367 -73775 -26317 -73758
rect -26259 -73758 -26059 -73711
rect -26259 -73775 -26209 -73758
rect -26367 -73792 -26351 -73775
rect -26483 -73808 -26351 -73792
rect -26225 -73792 -26209 -73775
rect -26109 -73775 -26059 -73758
rect -26001 -73758 -25801 -73711
rect -26001 -73775 -25951 -73758
rect -26109 -73792 -26093 -73775
rect -26225 -73808 -26093 -73792
rect -25967 -73792 -25951 -73775
rect -25851 -73775 -25801 -73758
rect -25851 -73792 -25835 -73775
rect -25967 -73808 -25835 -73792
rect -27257 -74090 -27125 -74074
rect -27257 -74107 -27241 -74090
rect -27291 -74124 -27241 -74107
rect -27141 -74107 -27125 -74090
rect -26999 -74090 -26867 -74074
rect -26999 -74107 -26983 -74090
rect -27141 -74124 -27091 -74107
rect -27291 -74171 -27091 -74124
rect -27033 -74124 -26983 -74107
rect -26883 -74107 -26867 -74090
rect -26741 -74090 -26609 -74074
rect -26741 -74107 -26725 -74090
rect -26883 -74124 -26833 -74107
rect -27033 -74171 -26833 -74124
rect -26775 -74124 -26725 -74107
rect -26625 -74107 -26609 -74090
rect -26483 -74090 -26351 -74074
rect -26483 -74107 -26467 -74090
rect -26625 -74124 -26575 -74107
rect -26775 -74171 -26575 -74124
rect -26517 -74124 -26467 -74107
rect -26367 -74107 -26351 -74090
rect -26225 -74090 -26093 -74074
rect -26225 -74107 -26209 -74090
rect -26367 -74124 -26317 -74107
rect -26517 -74171 -26317 -74124
rect -26259 -74124 -26209 -74107
rect -26109 -74107 -26093 -74090
rect -25967 -74090 -25835 -74074
rect -25967 -74107 -25951 -74090
rect -26109 -74124 -26059 -74107
rect -26259 -74171 -26059 -74124
rect -26001 -74124 -25951 -74107
rect -25851 -74107 -25835 -74090
rect -25851 -74124 -25801 -74107
rect -26001 -74171 -25801 -74124
rect -27291 -74618 -27091 -74571
rect -27291 -74635 -27241 -74618
rect -27257 -74652 -27241 -74635
rect -27141 -74635 -27091 -74618
rect -27033 -74618 -26833 -74571
rect -27033 -74635 -26983 -74618
rect -27141 -74652 -27125 -74635
rect -27257 -74668 -27125 -74652
rect -26999 -74652 -26983 -74635
rect -26883 -74635 -26833 -74618
rect -26775 -74618 -26575 -74571
rect -26775 -74635 -26725 -74618
rect -26883 -74652 -26867 -74635
rect -26999 -74668 -26867 -74652
rect -26741 -74652 -26725 -74635
rect -26625 -74635 -26575 -74618
rect -26517 -74618 -26317 -74571
rect -26517 -74635 -26467 -74618
rect -26625 -74652 -26609 -74635
rect -26741 -74668 -26609 -74652
rect -26483 -74652 -26467 -74635
rect -26367 -74635 -26317 -74618
rect -26259 -74618 -26059 -74571
rect -26259 -74635 -26209 -74618
rect -26367 -74652 -26351 -74635
rect -26483 -74668 -26351 -74652
rect -26225 -74652 -26209 -74635
rect -26109 -74635 -26059 -74618
rect -26001 -74618 -25801 -74571
rect -26001 -74635 -25951 -74618
rect -26109 -74652 -26093 -74635
rect -26225 -74668 -26093 -74652
rect -25967 -74652 -25951 -74635
rect -25851 -74635 -25801 -74618
rect -25851 -74652 -25835 -74635
rect -25967 -74668 -25835 -74652
rect -19952 -72667 -19922 -72635
rect -23952 -72893 -23922 -72867
rect -23257 -73230 -23125 -73214
rect -23257 -73247 -23241 -73230
rect -23291 -73264 -23241 -73247
rect -23141 -73247 -23125 -73230
rect -22999 -73230 -22867 -73214
rect -22999 -73247 -22983 -73230
rect -23141 -73264 -23091 -73247
rect -23291 -73311 -23091 -73264
rect -23033 -73264 -22983 -73247
rect -22883 -73247 -22867 -73230
rect -22741 -73230 -22609 -73214
rect -22741 -73247 -22725 -73230
rect -22883 -73264 -22833 -73247
rect -23033 -73311 -22833 -73264
rect -22775 -73264 -22725 -73247
rect -22625 -73247 -22609 -73230
rect -22483 -73230 -22351 -73214
rect -22483 -73247 -22467 -73230
rect -22625 -73264 -22575 -73247
rect -22775 -73311 -22575 -73264
rect -22517 -73264 -22467 -73247
rect -22367 -73247 -22351 -73230
rect -22225 -73230 -22093 -73214
rect -22225 -73247 -22209 -73230
rect -22367 -73264 -22317 -73247
rect -22517 -73311 -22317 -73264
rect -22259 -73264 -22209 -73247
rect -22109 -73247 -22093 -73230
rect -21967 -73230 -21835 -73214
rect -21967 -73247 -21951 -73230
rect -22109 -73264 -22059 -73247
rect -22259 -73311 -22059 -73264
rect -22001 -73264 -21951 -73247
rect -21851 -73247 -21835 -73230
rect -21851 -73264 -21801 -73247
rect -22001 -73311 -21801 -73264
rect -23291 -73758 -23091 -73711
rect -23291 -73775 -23241 -73758
rect -23257 -73792 -23241 -73775
rect -23141 -73775 -23091 -73758
rect -23033 -73758 -22833 -73711
rect -23033 -73775 -22983 -73758
rect -23141 -73792 -23125 -73775
rect -23257 -73808 -23125 -73792
rect -22999 -73792 -22983 -73775
rect -22883 -73775 -22833 -73758
rect -22775 -73758 -22575 -73711
rect -22775 -73775 -22725 -73758
rect -22883 -73792 -22867 -73775
rect -22999 -73808 -22867 -73792
rect -22741 -73792 -22725 -73775
rect -22625 -73775 -22575 -73758
rect -22517 -73758 -22317 -73711
rect -22517 -73775 -22467 -73758
rect -22625 -73792 -22609 -73775
rect -22741 -73808 -22609 -73792
rect -22483 -73792 -22467 -73775
rect -22367 -73775 -22317 -73758
rect -22259 -73758 -22059 -73711
rect -22259 -73775 -22209 -73758
rect -22367 -73792 -22351 -73775
rect -22483 -73808 -22351 -73792
rect -22225 -73792 -22209 -73775
rect -22109 -73775 -22059 -73758
rect -22001 -73758 -21801 -73711
rect -22001 -73775 -21951 -73758
rect -22109 -73792 -22093 -73775
rect -22225 -73808 -22093 -73792
rect -21967 -73792 -21951 -73775
rect -21851 -73775 -21801 -73758
rect -21851 -73792 -21835 -73775
rect -21967 -73808 -21835 -73792
rect -23257 -74090 -23125 -74074
rect -23257 -74107 -23241 -74090
rect -23291 -74124 -23241 -74107
rect -23141 -74107 -23125 -74090
rect -22999 -74090 -22867 -74074
rect -22999 -74107 -22983 -74090
rect -23141 -74124 -23091 -74107
rect -23291 -74171 -23091 -74124
rect -23033 -74124 -22983 -74107
rect -22883 -74107 -22867 -74090
rect -22741 -74090 -22609 -74074
rect -22741 -74107 -22725 -74090
rect -22883 -74124 -22833 -74107
rect -23033 -74171 -22833 -74124
rect -22775 -74124 -22725 -74107
rect -22625 -74107 -22609 -74090
rect -22483 -74090 -22351 -74074
rect -22483 -74107 -22467 -74090
rect -22625 -74124 -22575 -74107
rect -22775 -74171 -22575 -74124
rect -22517 -74124 -22467 -74107
rect -22367 -74107 -22351 -74090
rect -22225 -74090 -22093 -74074
rect -22225 -74107 -22209 -74090
rect -22367 -74124 -22317 -74107
rect -22517 -74171 -22317 -74124
rect -22259 -74124 -22209 -74107
rect -22109 -74107 -22093 -74090
rect -21967 -74090 -21835 -74074
rect -21967 -74107 -21951 -74090
rect -22109 -74124 -22059 -74107
rect -22259 -74171 -22059 -74124
rect -22001 -74124 -21951 -74107
rect -21851 -74107 -21835 -74090
rect -21851 -74124 -21801 -74107
rect -22001 -74171 -21801 -74124
rect -23291 -74618 -23091 -74571
rect -23291 -74635 -23241 -74618
rect -23257 -74652 -23241 -74635
rect -23141 -74635 -23091 -74618
rect -23033 -74618 -22833 -74571
rect -23033 -74635 -22983 -74618
rect -23141 -74652 -23125 -74635
rect -23257 -74668 -23125 -74652
rect -22999 -74652 -22983 -74635
rect -22883 -74635 -22833 -74618
rect -22775 -74618 -22575 -74571
rect -22775 -74635 -22725 -74618
rect -22883 -74652 -22867 -74635
rect -22999 -74668 -22867 -74652
rect -22741 -74652 -22725 -74635
rect -22625 -74635 -22575 -74618
rect -22517 -74618 -22317 -74571
rect -22517 -74635 -22467 -74618
rect -22625 -74652 -22609 -74635
rect -22741 -74668 -22609 -74652
rect -22483 -74652 -22467 -74635
rect -22367 -74635 -22317 -74618
rect -22259 -74618 -22059 -74571
rect -22259 -74635 -22209 -74618
rect -22367 -74652 -22351 -74635
rect -22483 -74668 -22351 -74652
rect -22225 -74652 -22209 -74635
rect -22109 -74635 -22059 -74618
rect -22001 -74618 -21801 -74571
rect -22001 -74635 -21951 -74618
rect -22109 -74652 -22093 -74635
rect -22225 -74668 -22093 -74652
rect -21967 -74652 -21951 -74635
rect -21851 -74635 -21801 -74618
rect -21851 -74652 -21835 -74635
rect -21967 -74668 -21835 -74652
rect -15952 -72667 -15922 -72635
rect -19952 -72893 -19922 -72867
rect -19257 -73230 -19125 -73214
rect -19257 -73247 -19241 -73230
rect -19291 -73264 -19241 -73247
rect -19141 -73247 -19125 -73230
rect -18999 -73230 -18867 -73214
rect -18999 -73247 -18983 -73230
rect -19141 -73264 -19091 -73247
rect -19291 -73311 -19091 -73264
rect -19033 -73264 -18983 -73247
rect -18883 -73247 -18867 -73230
rect -18741 -73230 -18609 -73214
rect -18741 -73247 -18725 -73230
rect -18883 -73264 -18833 -73247
rect -19033 -73311 -18833 -73264
rect -18775 -73264 -18725 -73247
rect -18625 -73247 -18609 -73230
rect -18483 -73230 -18351 -73214
rect -18483 -73247 -18467 -73230
rect -18625 -73264 -18575 -73247
rect -18775 -73311 -18575 -73264
rect -18517 -73264 -18467 -73247
rect -18367 -73247 -18351 -73230
rect -18225 -73230 -18093 -73214
rect -18225 -73247 -18209 -73230
rect -18367 -73264 -18317 -73247
rect -18517 -73311 -18317 -73264
rect -18259 -73264 -18209 -73247
rect -18109 -73247 -18093 -73230
rect -17967 -73230 -17835 -73214
rect -17967 -73247 -17951 -73230
rect -18109 -73264 -18059 -73247
rect -18259 -73311 -18059 -73264
rect -18001 -73264 -17951 -73247
rect -17851 -73247 -17835 -73230
rect -17851 -73264 -17801 -73247
rect -18001 -73311 -17801 -73264
rect -19291 -73758 -19091 -73711
rect -19291 -73775 -19241 -73758
rect -19257 -73792 -19241 -73775
rect -19141 -73775 -19091 -73758
rect -19033 -73758 -18833 -73711
rect -19033 -73775 -18983 -73758
rect -19141 -73792 -19125 -73775
rect -19257 -73808 -19125 -73792
rect -18999 -73792 -18983 -73775
rect -18883 -73775 -18833 -73758
rect -18775 -73758 -18575 -73711
rect -18775 -73775 -18725 -73758
rect -18883 -73792 -18867 -73775
rect -18999 -73808 -18867 -73792
rect -18741 -73792 -18725 -73775
rect -18625 -73775 -18575 -73758
rect -18517 -73758 -18317 -73711
rect -18517 -73775 -18467 -73758
rect -18625 -73792 -18609 -73775
rect -18741 -73808 -18609 -73792
rect -18483 -73792 -18467 -73775
rect -18367 -73775 -18317 -73758
rect -18259 -73758 -18059 -73711
rect -18259 -73775 -18209 -73758
rect -18367 -73792 -18351 -73775
rect -18483 -73808 -18351 -73792
rect -18225 -73792 -18209 -73775
rect -18109 -73775 -18059 -73758
rect -18001 -73758 -17801 -73711
rect -18001 -73775 -17951 -73758
rect -18109 -73792 -18093 -73775
rect -18225 -73808 -18093 -73792
rect -17967 -73792 -17951 -73775
rect -17851 -73775 -17801 -73758
rect -17851 -73792 -17835 -73775
rect -17967 -73808 -17835 -73792
rect -19257 -74090 -19125 -74074
rect -19257 -74107 -19241 -74090
rect -19291 -74124 -19241 -74107
rect -19141 -74107 -19125 -74090
rect -18999 -74090 -18867 -74074
rect -18999 -74107 -18983 -74090
rect -19141 -74124 -19091 -74107
rect -19291 -74171 -19091 -74124
rect -19033 -74124 -18983 -74107
rect -18883 -74107 -18867 -74090
rect -18741 -74090 -18609 -74074
rect -18741 -74107 -18725 -74090
rect -18883 -74124 -18833 -74107
rect -19033 -74171 -18833 -74124
rect -18775 -74124 -18725 -74107
rect -18625 -74107 -18609 -74090
rect -18483 -74090 -18351 -74074
rect -18483 -74107 -18467 -74090
rect -18625 -74124 -18575 -74107
rect -18775 -74171 -18575 -74124
rect -18517 -74124 -18467 -74107
rect -18367 -74107 -18351 -74090
rect -18225 -74090 -18093 -74074
rect -18225 -74107 -18209 -74090
rect -18367 -74124 -18317 -74107
rect -18517 -74171 -18317 -74124
rect -18259 -74124 -18209 -74107
rect -18109 -74107 -18093 -74090
rect -17967 -74090 -17835 -74074
rect -17967 -74107 -17951 -74090
rect -18109 -74124 -18059 -74107
rect -18259 -74171 -18059 -74124
rect -18001 -74124 -17951 -74107
rect -17851 -74107 -17835 -74090
rect -17851 -74124 -17801 -74107
rect -18001 -74171 -17801 -74124
rect -19291 -74618 -19091 -74571
rect -19291 -74635 -19241 -74618
rect -19257 -74652 -19241 -74635
rect -19141 -74635 -19091 -74618
rect -19033 -74618 -18833 -74571
rect -19033 -74635 -18983 -74618
rect -19141 -74652 -19125 -74635
rect -19257 -74668 -19125 -74652
rect -18999 -74652 -18983 -74635
rect -18883 -74635 -18833 -74618
rect -18775 -74618 -18575 -74571
rect -18775 -74635 -18725 -74618
rect -18883 -74652 -18867 -74635
rect -18999 -74668 -18867 -74652
rect -18741 -74652 -18725 -74635
rect -18625 -74635 -18575 -74618
rect -18517 -74618 -18317 -74571
rect -18517 -74635 -18467 -74618
rect -18625 -74652 -18609 -74635
rect -18741 -74668 -18609 -74652
rect -18483 -74652 -18467 -74635
rect -18367 -74635 -18317 -74618
rect -18259 -74618 -18059 -74571
rect -18259 -74635 -18209 -74618
rect -18367 -74652 -18351 -74635
rect -18483 -74668 -18351 -74652
rect -18225 -74652 -18209 -74635
rect -18109 -74635 -18059 -74618
rect -18001 -74618 -17801 -74571
rect -18001 -74635 -17951 -74618
rect -18109 -74652 -18093 -74635
rect -18225 -74668 -18093 -74652
rect -17967 -74652 -17951 -74635
rect -17851 -74635 -17801 -74618
rect -17851 -74652 -17835 -74635
rect -17967 -74668 -17835 -74652
rect -11952 -72667 -11922 -72635
rect -15952 -72893 -15922 -72867
rect -15257 -73230 -15125 -73214
rect -15257 -73247 -15241 -73230
rect -15291 -73264 -15241 -73247
rect -15141 -73247 -15125 -73230
rect -14999 -73230 -14867 -73214
rect -14999 -73247 -14983 -73230
rect -15141 -73264 -15091 -73247
rect -15291 -73311 -15091 -73264
rect -15033 -73264 -14983 -73247
rect -14883 -73247 -14867 -73230
rect -14741 -73230 -14609 -73214
rect -14741 -73247 -14725 -73230
rect -14883 -73264 -14833 -73247
rect -15033 -73311 -14833 -73264
rect -14775 -73264 -14725 -73247
rect -14625 -73247 -14609 -73230
rect -14483 -73230 -14351 -73214
rect -14483 -73247 -14467 -73230
rect -14625 -73264 -14575 -73247
rect -14775 -73311 -14575 -73264
rect -14517 -73264 -14467 -73247
rect -14367 -73247 -14351 -73230
rect -14225 -73230 -14093 -73214
rect -14225 -73247 -14209 -73230
rect -14367 -73264 -14317 -73247
rect -14517 -73311 -14317 -73264
rect -14259 -73264 -14209 -73247
rect -14109 -73247 -14093 -73230
rect -13967 -73230 -13835 -73214
rect -13967 -73247 -13951 -73230
rect -14109 -73264 -14059 -73247
rect -14259 -73311 -14059 -73264
rect -14001 -73264 -13951 -73247
rect -13851 -73247 -13835 -73230
rect -13851 -73264 -13801 -73247
rect -14001 -73311 -13801 -73264
rect -15291 -73758 -15091 -73711
rect -15291 -73775 -15241 -73758
rect -15257 -73792 -15241 -73775
rect -15141 -73775 -15091 -73758
rect -15033 -73758 -14833 -73711
rect -15033 -73775 -14983 -73758
rect -15141 -73792 -15125 -73775
rect -15257 -73808 -15125 -73792
rect -14999 -73792 -14983 -73775
rect -14883 -73775 -14833 -73758
rect -14775 -73758 -14575 -73711
rect -14775 -73775 -14725 -73758
rect -14883 -73792 -14867 -73775
rect -14999 -73808 -14867 -73792
rect -14741 -73792 -14725 -73775
rect -14625 -73775 -14575 -73758
rect -14517 -73758 -14317 -73711
rect -14517 -73775 -14467 -73758
rect -14625 -73792 -14609 -73775
rect -14741 -73808 -14609 -73792
rect -14483 -73792 -14467 -73775
rect -14367 -73775 -14317 -73758
rect -14259 -73758 -14059 -73711
rect -14259 -73775 -14209 -73758
rect -14367 -73792 -14351 -73775
rect -14483 -73808 -14351 -73792
rect -14225 -73792 -14209 -73775
rect -14109 -73775 -14059 -73758
rect -14001 -73758 -13801 -73711
rect -14001 -73775 -13951 -73758
rect -14109 -73792 -14093 -73775
rect -14225 -73808 -14093 -73792
rect -13967 -73792 -13951 -73775
rect -13851 -73775 -13801 -73758
rect -13851 -73792 -13835 -73775
rect -13967 -73808 -13835 -73792
rect -15257 -74090 -15125 -74074
rect -15257 -74107 -15241 -74090
rect -15291 -74124 -15241 -74107
rect -15141 -74107 -15125 -74090
rect -14999 -74090 -14867 -74074
rect -14999 -74107 -14983 -74090
rect -15141 -74124 -15091 -74107
rect -15291 -74171 -15091 -74124
rect -15033 -74124 -14983 -74107
rect -14883 -74107 -14867 -74090
rect -14741 -74090 -14609 -74074
rect -14741 -74107 -14725 -74090
rect -14883 -74124 -14833 -74107
rect -15033 -74171 -14833 -74124
rect -14775 -74124 -14725 -74107
rect -14625 -74107 -14609 -74090
rect -14483 -74090 -14351 -74074
rect -14483 -74107 -14467 -74090
rect -14625 -74124 -14575 -74107
rect -14775 -74171 -14575 -74124
rect -14517 -74124 -14467 -74107
rect -14367 -74107 -14351 -74090
rect -14225 -74090 -14093 -74074
rect -14225 -74107 -14209 -74090
rect -14367 -74124 -14317 -74107
rect -14517 -74171 -14317 -74124
rect -14259 -74124 -14209 -74107
rect -14109 -74107 -14093 -74090
rect -13967 -74090 -13835 -74074
rect -13967 -74107 -13951 -74090
rect -14109 -74124 -14059 -74107
rect -14259 -74171 -14059 -74124
rect -14001 -74124 -13951 -74107
rect -13851 -74107 -13835 -74090
rect -13851 -74124 -13801 -74107
rect -14001 -74171 -13801 -74124
rect -15291 -74618 -15091 -74571
rect -15291 -74635 -15241 -74618
rect -15257 -74652 -15241 -74635
rect -15141 -74635 -15091 -74618
rect -15033 -74618 -14833 -74571
rect -15033 -74635 -14983 -74618
rect -15141 -74652 -15125 -74635
rect -15257 -74668 -15125 -74652
rect -14999 -74652 -14983 -74635
rect -14883 -74635 -14833 -74618
rect -14775 -74618 -14575 -74571
rect -14775 -74635 -14725 -74618
rect -14883 -74652 -14867 -74635
rect -14999 -74668 -14867 -74652
rect -14741 -74652 -14725 -74635
rect -14625 -74635 -14575 -74618
rect -14517 -74618 -14317 -74571
rect -14517 -74635 -14467 -74618
rect -14625 -74652 -14609 -74635
rect -14741 -74668 -14609 -74652
rect -14483 -74652 -14467 -74635
rect -14367 -74635 -14317 -74618
rect -14259 -74618 -14059 -74571
rect -14259 -74635 -14209 -74618
rect -14367 -74652 -14351 -74635
rect -14483 -74668 -14351 -74652
rect -14225 -74652 -14209 -74635
rect -14109 -74635 -14059 -74618
rect -14001 -74618 -13801 -74571
rect -14001 -74635 -13951 -74618
rect -14109 -74652 -14093 -74635
rect -14225 -74668 -14093 -74652
rect -13967 -74652 -13951 -74635
rect -13851 -74635 -13801 -74618
rect -13851 -74652 -13835 -74635
rect -13967 -74668 -13835 -74652
rect -7952 -72667 -7922 -72635
rect -11952 -72893 -11922 -72867
rect -11257 -73230 -11125 -73214
rect -11257 -73247 -11241 -73230
rect -11291 -73264 -11241 -73247
rect -11141 -73247 -11125 -73230
rect -10999 -73230 -10867 -73214
rect -10999 -73247 -10983 -73230
rect -11141 -73264 -11091 -73247
rect -11291 -73311 -11091 -73264
rect -11033 -73264 -10983 -73247
rect -10883 -73247 -10867 -73230
rect -10741 -73230 -10609 -73214
rect -10741 -73247 -10725 -73230
rect -10883 -73264 -10833 -73247
rect -11033 -73311 -10833 -73264
rect -10775 -73264 -10725 -73247
rect -10625 -73247 -10609 -73230
rect -10483 -73230 -10351 -73214
rect -10483 -73247 -10467 -73230
rect -10625 -73264 -10575 -73247
rect -10775 -73311 -10575 -73264
rect -10517 -73264 -10467 -73247
rect -10367 -73247 -10351 -73230
rect -10225 -73230 -10093 -73214
rect -10225 -73247 -10209 -73230
rect -10367 -73264 -10317 -73247
rect -10517 -73311 -10317 -73264
rect -10259 -73264 -10209 -73247
rect -10109 -73247 -10093 -73230
rect -9967 -73230 -9835 -73214
rect -9967 -73247 -9951 -73230
rect -10109 -73264 -10059 -73247
rect -10259 -73311 -10059 -73264
rect -10001 -73264 -9951 -73247
rect -9851 -73247 -9835 -73230
rect -9851 -73264 -9801 -73247
rect -10001 -73311 -9801 -73264
rect -11291 -73758 -11091 -73711
rect -11291 -73775 -11241 -73758
rect -11257 -73792 -11241 -73775
rect -11141 -73775 -11091 -73758
rect -11033 -73758 -10833 -73711
rect -11033 -73775 -10983 -73758
rect -11141 -73792 -11125 -73775
rect -11257 -73808 -11125 -73792
rect -10999 -73792 -10983 -73775
rect -10883 -73775 -10833 -73758
rect -10775 -73758 -10575 -73711
rect -10775 -73775 -10725 -73758
rect -10883 -73792 -10867 -73775
rect -10999 -73808 -10867 -73792
rect -10741 -73792 -10725 -73775
rect -10625 -73775 -10575 -73758
rect -10517 -73758 -10317 -73711
rect -10517 -73775 -10467 -73758
rect -10625 -73792 -10609 -73775
rect -10741 -73808 -10609 -73792
rect -10483 -73792 -10467 -73775
rect -10367 -73775 -10317 -73758
rect -10259 -73758 -10059 -73711
rect -10259 -73775 -10209 -73758
rect -10367 -73792 -10351 -73775
rect -10483 -73808 -10351 -73792
rect -10225 -73792 -10209 -73775
rect -10109 -73775 -10059 -73758
rect -10001 -73758 -9801 -73711
rect -10001 -73775 -9951 -73758
rect -10109 -73792 -10093 -73775
rect -10225 -73808 -10093 -73792
rect -9967 -73792 -9951 -73775
rect -9851 -73775 -9801 -73758
rect -9851 -73792 -9835 -73775
rect -9967 -73808 -9835 -73792
rect -11257 -74090 -11125 -74074
rect -11257 -74107 -11241 -74090
rect -11291 -74124 -11241 -74107
rect -11141 -74107 -11125 -74090
rect -10999 -74090 -10867 -74074
rect -10999 -74107 -10983 -74090
rect -11141 -74124 -11091 -74107
rect -11291 -74171 -11091 -74124
rect -11033 -74124 -10983 -74107
rect -10883 -74107 -10867 -74090
rect -10741 -74090 -10609 -74074
rect -10741 -74107 -10725 -74090
rect -10883 -74124 -10833 -74107
rect -11033 -74171 -10833 -74124
rect -10775 -74124 -10725 -74107
rect -10625 -74107 -10609 -74090
rect -10483 -74090 -10351 -74074
rect -10483 -74107 -10467 -74090
rect -10625 -74124 -10575 -74107
rect -10775 -74171 -10575 -74124
rect -10517 -74124 -10467 -74107
rect -10367 -74107 -10351 -74090
rect -10225 -74090 -10093 -74074
rect -10225 -74107 -10209 -74090
rect -10367 -74124 -10317 -74107
rect -10517 -74171 -10317 -74124
rect -10259 -74124 -10209 -74107
rect -10109 -74107 -10093 -74090
rect -9967 -74090 -9835 -74074
rect -9967 -74107 -9951 -74090
rect -10109 -74124 -10059 -74107
rect -10259 -74171 -10059 -74124
rect -10001 -74124 -9951 -74107
rect -9851 -74107 -9835 -74090
rect -9851 -74124 -9801 -74107
rect -10001 -74171 -9801 -74124
rect -11291 -74618 -11091 -74571
rect -11291 -74635 -11241 -74618
rect -11257 -74652 -11241 -74635
rect -11141 -74635 -11091 -74618
rect -11033 -74618 -10833 -74571
rect -11033 -74635 -10983 -74618
rect -11141 -74652 -11125 -74635
rect -11257 -74668 -11125 -74652
rect -10999 -74652 -10983 -74635
rect -10883 -74635 -10833 -74618
rect -10775 -74618 -10575 -74571
rect -10775 -74635 -10725 -74618
rect -10883 -74652 -10867 -74635
rect -10999 -74668 -10867 -74652
rect -10741 -74652 -10725 -74635
rect -10625 -74635 -10575 -74618
rect -10517 -74618 -10317 -74571
rect -10517 -74635 -10467 -74618
rect -10625 -74652 -10609 -74635
rect -10741 -74668 -10609 -74652
rect -10483 -74652 -10467 -74635
rect -10367 -74635 -10317 -74618
rect -10259 -74618 -10059 -74571
rect -10259 -74635 -10209 -74618
rect -10367 -74652 -10351 -74635
rect -10483 -74668 -10351 -74652
rect -10225 -74652 -10209 -74635
rect -10109 -74635 -10059 -74618
rect -10001 -74618 -9801 -74571
rect -10001 -74635 -9951 -74618
rect -10109 -74652 -10093 -74635
rect -10225 -74668 -10093 -74652
rect -9967 -74652 -9951 -74635
rect -9851 -74635 -9801 -74618
rect -9851 -74652 -9835 -74635
rect -9967 -74668 -9835 -74652
rect -3952 -72667 -3922 -72635
rect -7952 -72893 -7922 -72867
rect -7257 -73230 -7125 -73214
rect -7257 -73247 -7241 -73230
rect -7291 -73264 -7241 -73247
rect -7141 -73247 -7125 -73230
rect -6999 -73230 -6867 -73214
rect -6999 -73247 -6983 -73230
rect -7141 -73264 -7091 -73247
rect -7291 -73311 -7091 -73264
rect -7033 -73264 -6983 -73247
rect -6883 -73247 -6867 -73230
rect -6741 -73230 -6609 -73214
rect -6741 -73247 -6725 -73230
rect -6883 -73264 -6833 -73247
rect -7033 -73311 -6833 -73264
rect -6775 -73264 -6725 -73247
rect -6625 -73247 -6609 -73230
rect -6483 -73230 -6351 -73214
rect -6483 -73247 -6467 -73230
rect -6625 -73264 -6575 -73247
rect -6775 -73311 -6575 -73264
rect -6517 -73264 -6467 -73247
rect -6367 -73247 -6351 -73230
rect -6225 -73230 -6093 -73214
rect -6225 -73247 -6209 -73230
rect -6367 -73264 -6317 -73247
rect -6517 -73311 -6317 -73264
rect -6259 -73264 -6209 -73247
rect -6109 -73247 -6093 -73230
rect -5967 -73230 -5835 -73214
rect -5967 -73247 -5951 -73230
rect -6109 -73264 -6059 -73247
rect -6259 -73311 -6059 -73264
rect -6001 -73264 -5951 -73247
rect -5851 -73247 -5835 -73230
rect -5851 -73264 -5801 -73247
rect -6001 -73311 -5801 -73264
rect -7291 -73758 -7091 -73711
rect -7291 -73775 -7241 -73758
rect -7257 -73792 -7241 -73775
rect -7141 -73775 -7091 -73758
rect -7033 -73758 -6833 -73711
rect -7033 -73775 -6983 -73758
rect -7141 -73792 -7125 -73775
rect -7257 -73808 -7125 -73792
rect -6999 -73792 -6983 -73775
rect -6883 -73775 -6833 -73758
rect -6775 -73758 -6575 -73711
rect -6775 -73775 -6725 -73758
rect -6883 -73792 -6867 -73775
rect -6999 -73808 -6867 -73792
rect -6741 -73792 -6725 -73775
rect -6625 -73775 -6575 -73758
rect -6517 -73758 -6317 -73711
rect -6517 -73775 -6467 -73758
rect -6625 -73792 -6609 -73775
rect -6741 -73808 -6609 -73792
rect -6483 -73792 -6467 -73775
rect -6367 -73775 -6317 -73758
rect -6259 -73758 -6059 -73711
rect -6259 -73775 -6209 -73758
rect -6367 -73792 -6351 -73775
rect -6483 -73808 -6351 -73792
rect -6225 -73792 -6209 -73775
rect -6109 -73775 -6059 -73758
rect -6001 -73758 -5801 -73711
rect -6001 -73775 -5951 -73758
rect -6109 -73792 -6093 -73775
rect -6225 -73808 -6093 -73792
rect -5967 -73792 -5951 -73775
rect -5851 -73775 -5801 -73758
rect -5851 -73792 -5835 -73775
rect -5967 -73808 -5835 -73792
rect -7257 -74090 -7125 -74074
rect -7257 -74107 -7241 -74090
rect -7291 -74124 -7241 -74107
rect -7141 -74107 -7125 -74090
rect -6999 -74090 -6867 -74074
rect -6999 -74107 -6983 -74090
rect -7141 -74124 -7091 -74107
rect -7291 -74171 -7091 -74124
rect -7033 -74124 -6983 -74107
rect -6883 -74107 -6867 -74090
rect -6741 -74090 -6609 -74074
rect -6741 -74107 -6725 -74090
rect -6883 -74124 -6833 -74107
rect -7033 -74171 -6833 -74124
rect -6775 -74124 -6725 -74107
rect -6625 -74107 -6609 -74090
rect -6483 -74090 -6351 -74074
rect -6483 -74107 -6467 -74090
rect -6625 -74124 -6575 -74107
rect -6775 -74171 -6575 -74124
rect -6517 -74124 -6467 -74107
rect -6367 -74107 -6351 -74090
rect -6225 -74090 -6093 -74074
rect -6225 -74107 -6209 -74090
rect -6367 -74124 -6317 -74107
rect -6517 -74171 -6317 -74124
rect -6259 -74124 -6209 -74107
rect -6109 -74107 -6093 -74090
rect -5967 -74090 -5835 -74074
rect -5967 -74107 -5951 -74090
rect -6109 -74124 -6059 -74107
rect -6259 -74171 -6059 -74124
rect -6001 -74124 -5951 -74107
rect -5851 -74107 -5835 -74090
rect -5851 -74124 -5801 -74107
rect -6001 -74171 -5801 -74124
rect -7291 -74618 -7091 -74571
rect -7291 -74635 -7241 -74618
rect -7257 -74652 -7241 -74635
rect -7141 -74635 -7091 -74618
rect -7033 -74618 -6833 -74571
rect -7033 -74635 -6983 -74618
rect -7141 -74652 -7125 -74635
rect -7257 -74668 -7125 -74652
rect -6999 -74652 -6983 -74635
rect -6883 -74635 -6833 -74618
rect -6775 -74618 -6575 -74571
rect -6775 -74635 -6725 -74618
rect -6883 -74652 -6867 -74635
rect -6999 -74668 -6867 -74652
rect -6741 -74652 -6725 -74635
rect -6625 -74635 -6575 -74618
rect -6517 -74618 -6317 -74571
rect -6517 -74635 -6467 -74618
rect -6625 -74652 -6609 -74635
rect -6741 -74668 -6609 -74652
rect -6483 -74652 -6467 -74635
rect -6367 -74635 -6317 -74618
rect -6259 -74618 -6059 -74571
rect -6259 -74635 -6209 -74618
rect -6367 -74652 -6351 -74635
rect -6483 -74668 -6351 -74652
rect -6225 -74652 -6209 -74635
rect -6109 -74635 -6059 -74618
rect -6001 -74618 -5801 -74571
rect -6001 -74635 -5951 -74618
rect -6109 -74652 -6093 -74635
rect -6225 -74668 -6093 -74652
rect -5967 -74652 -5951 -74635
rect -5851 -74635 -5801 -74618
rect -5851 -74652 -5835 -74635
rect -5967 -74668 -5835 -74652
rect 48 -72667 78 -72635
rect -3952 -72893 -3922 -72867
rect -3257 -73230 -3125 -73214
rect -3257 -73247 -3241 -73230
rect -3291 -73264 -3241 -73247
rect -3141 -73247 -3125 -73230
rect -2999 -73230 -2867 -73214
rect -2999 -73247 -2983 -73230
rect -3141 -73264 -3091 -73247
rect -3291 -73311 -3091 -73264
rect -3033 -73264 -2983 -73247
rect -2883 -73247 -2867 -73230
rect -2741 -73230 -2609 -73214
rect -2741 -73247 -2725 -73230
rect -2883 -73264 -2833 -73247
rect -3033 -73311 -2833 -73264
rect -2775 -73264 -2725 -73247
rect -2625 -73247 -2609 -73230
rect -2483 -73230 -2351 -73214
rect -2483 -73247 -2467 -73230
rect -2625 -73264 -2575 -73247
rect -2775 -73311 -2575 -73264
rect -2517 -73264 -2467 -73247
rect -2367 -73247 -2351 -73230
rect -2225 -73230 -2093 -73214
rect -2225 -73247 -2209 -73230
rect -2367 -73264 -2317 -73247
rect -2517 -73311 -2317 -73264
rect -2259 -73264 -2209 -73247
rect -2109 -73247 -2093 -73230
rect -1967 -73230 -1835 -73214
rect -1967 -73247 -1951 -73230
rect -2109 -73264 -2059 -73247
rect -2259 -73311 -2059 -73264
rect -2001 -73264 -1951 -73247
rect -1851 -73247 -1835 -73230
rect -1851 -73264 -1801 -73247
rect -2001 -73311 -1801 -73264
rect -3291 -73758 -3091 -73711
rect -3291 -73775 -3241 -73758
rect -3257 -73792 -3241 -73775
rect -3141 -73775 -3091 -73758
rect -3033 -73758 -2833 -73711
rect -3033 -73775 -2983 -73758
rect -3141 -73792 -3125 -73775
rect -3257 -73808 -3125 -73792
rect -2999 -73792 -2983 -73775
rect -2883 -73775 -2833 -73758
rect -2775 -73758 -2575 -73711
rect -2775 -73775 -2725 -73758
rect -2883 -73792 -2867 -73775
rect -2999 -73808 -2867 -73792
rect -2741 -73792 -2725 -73775
rect -2625 -73775 -2575 -73758
rect -2517 -73758 -2317 -73711
rect -2517 -73775 -2467 -73758
rect -2625 -73792 -2609 -73775
rect -2741 -73808 -2609 -73792
rect -2483 -73792 -2467 -73775
rect -2367 -73775 -2317 -73758
rect -2259 -73758 -2059 -73711
rect -2259 -73775 -2209 -73758
rect -2367 -73792 -2351 -73775
rect -2483 -73808 -2351 -73792
rect -2225 -73792 -2209 -73775
rect -2109 -73775 -2059 -73758
rect -2001 -73758 -1801 -73711
rect -2001 -73775 -1951 -73758
rect -2109 -73792 -2093 -73775
rect -2225 -73808 -2093 -73792
rect -1967 -73792 -1951 -73775
rect -1851 -73775 -1801 -73758
rect -1851 -73792 -1835 -73775
rect -1967 -73808 -1835 -73792
rect -3257 -74090 -3125 -74074
rect -3257 -74107 -3241 -74090
rect -3291 -74124 -3241 -74107
rect -3141 -74107 -3125 -74090
rect -2999 -74090 -2867 -74074
rect -2999 -74107 -2983 -74090
rect -3141 -74124 -3091 -74107
rect -3291 -74171 -3091 -74124
rect -3033 -74124 -2983 -74107
rect -2883 -74107 -2867 -74090
rect -2741 -74090 -2609 -74074
rect -2741 -74107 -2725 -74090
rect -2883 -74124 -2833 -74107
rect -3033 -74171 -2833 -74124
rect -2775 -74124 -2725 -74107
rect -2625 -74107 -2609 -74090
rect -2483 -74090 -2351 -74074
rect -2483 -74107 -2467 -74090
rect -2625 -74124 -2575 -74107
rect -2775 -74171 -2575 -74124
rect -2517 -74124 -2467 -74107
rect -2367 -74107 -2351 -74090
rect -2225 -74090 -2093 -74074
rect -2225 -74107 -2209 -74090
rect -2367 -74124 -2317 -74107
rect -2517 -74171 -2317 -74124
rect -2259 -74124 -2209 -74107
rect -2109 -74107 -2093 -74090
rect -1967 -74090 -1835 -74074
rect -1967 -74107 -1951 -74090
rect -2109 -74124 -2059 -74107
rect -2259 -74171 -2059 -74124
rect -2001 -74124 -1951 -74107
rect -1851 -74107 -1835 -74090
rect -1851 -74124 -1801 -74107
rect -2001 -74171 -1801 -74124
rect -3291 -74618 -3091 -74571
rect -3291 -74635 -3241 -74618
rect -3257 -74652 -3241 -74635
rect -3141 -74635 -3091 -74618
rect -3033 -74618 -2833 -74571
rect -3033 -74635 -2983 -74618
rect -3141 -74652 -3125 -74635
rect -3257 -74668 -3125 -74652
rect -2999 -74652 -2983 -74635
rect -2883 -74635 -2833 -74618
rect -2775 -74618 -2575 -74571
rect -2775 -74635 -2725 -74618
rect -2883 -74652 -2867 -74635
rect -2999 -74668 -2867 -74652
rect -2741 -74652 -2725 -74635
rect -2625 -74635 -2575 -74618
rect -2517 -74618 -2317 -74571
rect -2517 -74635 -2467 -74618
rect -2625 -74652 -2609 -74635
rect -2741 -74668 -2609 -74652
rect -2483 -74652 -2467 -74635
rect -2367 -74635 -2317 -74618
rect -2259 -74618 -2059 -74571
rect -2259 -74635 -2209 -74618
rect -2367 -74652 -2351 -74635
rect -2483 -74668 -2351 -74652
rect -2225 -74652 -2209 -74635
rect -2109 -74635 -2059 -74618
rect -2001 -74618 -1801 -74571
rect -2001 -74635 -1951 -74618
rect -2109 -74652 -2093 -74635
rect -2225 -74668 -2093 -74652
rect -1967 -74652 -1951 -74635
rect -1851 -74635 -1801 -74618
rect -1851 -74652 -1835 -74635
rect -1967 -74668 -1835 -74652
rect 4048 -72667 4078 -72635
rect 48 -72893 78 -72867
rect 743 -73230 875 -73214
rect 743 -73247 759 -73230
rect 709 -73264 759 -73247
rect 859 -73247 875 -73230
rect 1001 -73230 1133 -73214
rect 1001 -73247 1017 -73230
rect 859 -73264 909 -73247
rect 709 -73311 909 -73264
rect 967 -73264 1017 -73247
rect 1117 -73247 1133 -73230
rect 1259 -73230 1391 -73214
rect 1259 -73247 1275 -73230
rect 1117 -73264 1167 -73247
rect 967 -73311 1167 -73264
rect 1225 -73264 1275 -73247
rect 1375 -73247 1391 -73230
rect 1517 -73230 1649 -73214
rect 1517 -73247 1533 -73230
rect 1375 -73264 1425 -73247
rect 1225 -73311 1425 -73264
rect 1483 -73264 1533 -73247
rect 1633 -73247 1649 -73230
rect 1775 -73230 1907 -73214
rect 1775 -73247 1791 -73230
rect 1633 -73264 1683 -73247
rect 1483 -73311 1683 -73264
rect 1741 -73264 1791 -73247
rect 1891 -73247 1907 -73230
rect 2033 -73230 2165 -73214
rect 2033 -73247 2049 -73230
rect 1891 -73264 1941 -73247
rect 1741 -73311 1941 -73264
rect 1999 -73264 2049 -73247
rect 2149 -73247 2165 -73230
rect 2149 -73264 2199 -73247
rect 1999 -73311 2199 -73264
rect 709 -73758 909 -73711
rect 709 -73775 759 -73758
rect 743 -73792 759 -73775
rect 859 -73775 909 -73758
rect 967 -73758 1167 -73711
rect 967 -73775 1017 -73758
rect 859 -73792 875 -73775
rect 743 -73808 875 -73792
rect 1001 -73792 1017 -73775
rect 1117 -73775 1167 -73758
rect 1225 -73758 1425 -73711
rect 1225 -73775 1275 -73758
rect 1117 -73792 1133 -73775
rect 1001 -73808 1133 -73792
rect 1259 -73792 1275 -73775
rect 1375 -73775 1425 -73758
rect 1483 -73758 1683 -73711
rect 1483 -73775 1533 -73758
rect 1375 -73792 1391 -73775
rect 1259 -73808 1391 -73792
rect 1517 -73792 1533 -73775
rect 1633 -73775 1683 -73758
rect 1741 -73758 1941 -73711
rect 1741 -73775 1791 -73758
rect 1633 -73792 1649 -73775
rect 1517 -73808 1649 -73792
rect 1775 -73792 1791 -73775
rect 1891 -73775 1941 -73758
rect 1999 -73758 2199 -73711
rect 1999 -73775 2049 -73758
rect 1891 -73792 1907 -73775
rect 1775 -73808 1907 -73792
rect 2033 -73792 2049 -73775
rect 2149 -73775 2199 -73758
rect 2149 -73792 2165 -73775
rect 2033 -73808 2165 -73792
rect 743 -74090 875 -74074
rect 743 -74107 759 -74090
rect 709 -74124 759 -74107
rect 859 -74107 875 -74090
rect 1001 -74090 1133 -74074
rect 1001 -74107 1017 -74090
rect 859 -74124 909 -74107
rect 709 -74171 909 -74124
rect 967 -74124 1017 -74107
rect 1117 -74107 1133 -74090
rect 1259 -74090 1391 -74074
rect 1259 -74107 1275 -74090
rect 1117 -74124 1167 -74107
rect 967 -74171 1167 -74124
rect 1225 -74124 1275 -74107
rect 1375 -74107 1391 -74090
rect 1517 -74090 1649 -74074
rect 1517 -74107 1533 -74090
rect 1375 -74124 1425 -74107
rect 1225 -74171 1425 -74124
rect 1483 -74124 1533 -74107
rect 1633 -74107 1649 -74090
rect 1775 -74090 1907 -74074
rect 1775 -74107 1791 -74090
rect 1633 -74124 1683 -74107
rect 1483 -74171 1683 -74124
rect 1741 -74124 1791 -74107
rect 1891 -74107 1907 -74090
rect 2033 -74090 2165 -74074
rect 2033 -74107 2049 -74090
rect 1891 -74124 1941 -74107
rect 1741 -74171 1941 -74124
rect 1999 -74124 2049 -74107
rect 2149 -74107 2165 -74090
rect 2149 -74124 2199 -74107
rect 1999 -74171 2199 -74124
rect 709 -74618 909 -74571
rect 709 -74635 759 -74618
rect 743 -74652 759 -74635
rect 859 -74635 909 -74618
rect 967 -74618 1167 -74571
rect 967 -74635 1017 -74618
rect 859 -74652 875 -74635
rect 743 -74668 875 -74652
rect 1001 -74652 1017 -74635
rect 1117 -74635 1167 -74618
rect 1225 -74618 1425 -74571
rect 1225 -74635 1275 -74618
rect 1117 -74652 1133 -74635
rect 1001 -74668 1133 -74652
rect 1259 -74652 1275 -74635
rect 1375 -74635 1425 -74618
rect 1483 -74618 1683 -74571
rect 1483 -74635 1533 -74618
rect 1375 -74652 1391 -74635
rect 1259 -74668 1391 -74652
rect 1517 -74652 1533 -74635
rect 1633 -74635 1683 -74618
rect 1741 -74618 1941 -74571
rect 1741 -74635 1791 -74618
rect 1633 -74652 1649 -74635
rect 1517 -74668 1649 -74652
rect 1775 -74652 1791 -74635
rect 1891 -74635 1941 -74618
rect 1999 -74618 2199 -74571
rect 1999 -74635 2049 -74618
rect 1891 -74652 1907 -74635
rect 1775 -74668 1907 -74652
rect 2033 -74652 2049 -74635
rect 2149 -74635 2199 -74618
rect 2149 -74652 2165 -74635
rect 2033 -74668 2165 -74652
rect 4048 -72893 4078 -72867
rect 4743 -73230 4875 -73214
rect 4743 -73247 4759 -73230
rect 4709 -73264 4759 -73247
rect 4859 -73247 4875 -73230
rect 5001 -73230 5133 -73214
rect 5001 -73247 5017 -73230
rect 4859 -73264 4909 -73247
rect 4709 -73311 4909 -73264
rect 4967 -73264 5017 -73247
rect 5117 -73247 5133 -73230
rect 5259 -73230 5391 -73214
rect 5259 -73247 5275 -73230
rect 5117 -73264 5167 -73247
rect 4967 -73311 5167 -73264
rect 5225 -73264 5275 -73247
rect 5375 -73247 5391 -73230
rect 5517 -73230 5649 -73214
rect 5517 -73247 5533 -73230
rect 5375 -73264 5425 -73247
rect 5225 -73311 5425 -73264
rect 5483 -73264 5533 -73247
rect 5633 -73247 5649 -73230
rect 5775 -73230 5907 -73214
rect 5775 -73247 5791 -73230
rect 5633 -73264 5683 -73247
rect 5483 -73311 5683 -73264
rect 5741 -73264 5791 -73247
rect 5891 -73247 5907 -73230
rect 6033 -73230 6165 -73214
rect 6033 -73247 6049 -73230
rect 5891 -73264 5941 -73247
rect 5741 -73311 5941 -73264
rect 5999 -73264 6049 -73247
rect 6149 -73247 6165 -73230
rect 6149 -73264 6199 -73247
rect 5999 -73311 6199 -73264
rect 4709 -73758 4909 -73711
rect 4709 -73775 4759 -73758
rect 4743 -73792 4759 -73775
rect 4859 -73775 4909 -73758
rect 4967 -73758 5167 -73711
rect 4967 -73775 5017 -73758
rect 4859 -73792 4875 -73775
rect 4743 -73808 4875 -73792
rect 5001 -73792 5017 -73775
rect 5117 -73775 5167 -73758
rect 5225 -73758 5425 -73711
rect 5225 -73775 5275 -73758
rect 5117 -73792 5133 -73775
rect 5001 -73808 5133 -73792
rect 5259 -73792 5275 -73775
rect 5375 -73775 5425 -73758
rect 5483 -73758 5683 -73711
rect 5483 -73775 5533 -73758
rect 5375 -73792 5391 -73775
rect 5259 -73808 5391 -73792
rect 5517 -73792 5533 -73775
rect 5633 -73775 5683 -73758
rect 5741 -73758 5941 -73711
rect 5741 -73775 5791 -73758
rect 5633 -73792 5649 -73775
rect 5517 -73808 5649 -73792
rect 5775 -73792 5791 -73775
rect 5891 -73775 5941 -73758
rect 5999 -73758 6199 -73711
rect 5999 -73775 6049 -73758
rect 5891 -73792 5907 -73775
rect 5775 -73808 5907 -73792
rect 6033 -73792 6049 -73775
rect 6149 -73775 6199 -73758
rect 6149 -73792 6165 -73775
rect 6033 -73808 6165 -73792
rect 4743 -74090 4875 -74074
rect 4743 -74107 4759 -74090
rect 4709 -74124 4759 -74107
rect 4859 -74107 4875 -74090
rect 5001 -74090 5133 -74074
rect 5001 -74107 5017 -74090
rect 4859 -74124 4909 -74107
rect 4709 -74171 4909 -74124
rect 4967 -74124 5017 -74107
rect 5117 -74107 5133 -74090
rect 5259 -74090 5391 -74074
rect 5259 -74107 5275 -74090
rect 5117 -74124 5167 -74107
rect 4967 -74171 5167 -74124
rect 5225 -74124 5275 -74107
rect 5375 -74107 5391 -74090
rect 5517 -74090 5649 -74074
rect 5517 -74107 5533 -74090
rect 5375 -74124 5425 -74107
rect 5225 -74171 5425 -74124
rect 5483 -74124 5533 -74107
rect 5633 -74107 5649 -74090
rect 5775 -74090 5907 -74074
rect 5775 -74107 5791 -74090
rect 5633 -74124 5683 -74107
rect 5483 -74171 5683 -74124
rect 5741 -74124 5791 -74107
rect 5891 -74107 5907 -74090
rect 6033 -74090 6165 -74074
rect 6033 -74107 6049 -74090
rect 5891 -74124 5941 -74107
rect 5741 -74171 5941 -74124
rect 5999 -74124 6049 -74107
rect 6149 -74107 6165 -74090
rect 6149 -74124 6199 -74107
rect 5999 -74171 6199 -74124
rect 4709 -74618 4909 -74571
rect 4709 -74635 4759 -74618
rect 4743 -74652 4759 -74635
rect 4859 -74635 4909 -74618
rect 4967 -74618 5167 -74571
rect 4967 -74635 5017 -74618
rect 4859 -74652 4875 -74635
rect 4743 -74668 4875 -74652
rect 5001 -74652 5017 -74635
rect 5117 -74635 5167 -74618
rect 5225 -74618 5425 -74571
rect 5225 -74635 5275 -74618
rect 5117 -74652 5133 -74635
rect 5001 -74668 5133 -74652
rect 5259 -74652 5275 -74635
rect 5375 -74635 5425 -74618
rect 5483 -74618 5683 -74571
rect 5483 -74635 5533 -74618
rect 5375 -74652 5391 -74635
rect 5259 -74668 5391 -74652
rect 5517 -74652 5533 -74635
rect 5633 -74635 5683 -74618
rect 5741 -74618 5941 -74571
rect 5741 -74635 5791 -74618
rect 5633 -74652 5649 -74635
rect 5517 -74668 5649 -74652
rect 5775 -74652 5791 -74635
rect 5891 -74635 5941 -74618
rect 5999 -74618 6199 -74571
rect 5999 -74635 6049 -74618
rect 5891 -74652 5907 -74635
rect 5775 -74668 5907 -74652
rect 6033 -74652 6049 -74635
rect 6149 -74635 6199 -74618
rect 6149 -74652 6165 -74635
rect 6033 -74668 6165 -74652
<< polycont >>
rect 32180 -30457 32736 -30423
rect 33198 -30457 33754 -30423
rect 34216 -30457 34772 -30423
rect 35234 -30457 35790 -30423
rect 36252 -30457 36808 -30423
rect 37270 -30457 37826 -30423
rect 38288 -30457 38844 -30423
rect 39306 -30457 39862 -30423
rect 40324 -30457 40880 -30423
rect 41342 -30457 41898 -30423
rect 42360 -30457 42916 -30423
rect 43378 -30457 43934 -30423
rect 44396 -30457 44952 -30423
rect 45414 -30457 45970 -30423
rect 46432 -30457 46988 -30423
rect 47450 -30457 48006 -30423
rect 32180 -31185 32736 -31151
rect 33198 -31185 33754 -31151
rect 34216 -31185 34772 -31151
rect 35234 -31185 35790 -31151
rect 36252 -31185 36808 -31151
rect 37270 -31185 37826 -31151
rect 38288 -31185 38844 -31151
rect 39306 -31185 39862 -31151
rect 40324 -31185 40880 -31151
rect 41342 -31185 41898 -31151
rect 42360 -31185 42916 -31151
rect 43378 -31185 43934 -31151
rect 44396 -31185 44952 -31151
rect 45414 -31185 45970 -31151
rect 46432 -31185 46988 -31151
rect 47450 -31185 48006 -31151
rect 32180 -31593 32736 -31559
rect 33198 -31593 33754 -31559
rect 34216 -31593 34772 -31559
rect 35234 -31593 35790 -31559
rect 36252 -31593 36808 -31559
rect 37270 -31593 37826 -31559
rect 38288 -31593 38844 -31559
rect 39306 -31593 39862 -31559
rect 40324 -31593 40880 -31559
rect 41342 -31593 41898 -31559
rect 42360 -31593 42916 -31559
rect 43378 -31593 43934 -31559
rect 44396 -31593 44952 -31559
rect 45414 -31593 45970 -31559
rect 46432 -31593 46988 -31559
rect 47450 -31593 48006 -31559
rect 32180 -32321 32736 -32287
rect 33198 -32321 33754 -32287
rect 34216 -32321 34772 -32287
rect 35234 -32321 35790 -32287
rect 36252 -32321 36808 -32287
rect 37270 -32321 37826 -32287
rect 38288 -32321 38844 -32287
rect 39306 -32321 39862 -32287
rect 40324 -32321 40880 -32287
rect 41342 -32321 41898 -32287
rect 42360 -32321 42916 -32287
rect 43378 -32321 43934 -32287
rect 44396 -32321 44952 -32287
rect 45414 -32321 45970 -32287
rect 46432 -32321 46988 -32287
rect 47450 -32321 48006 -32287
rect 32180 -32729 32736 -32695
rect 33198 -32729 33754 -32695
rect 34216 -32729 34772 -32695
rect 35234 -32729 35790 -32695
rect 36252 -32729 36808 -32695
rect 37270 -32729 37826 -32695
rect 38288 -32729 38844 -32695
rect 39306 -32729 39862 -32695
rect 40324 -32729 40880 -32695
rect 41342 -32729 41898 -32695
rect 42360 -32729 42916 -32695
rect 43378 -32729 43934 -32695
rect 44396 -32729 44952 -32695
rect 45414 -32729 45970 -32695
rect 46432 -32729 46988 -32695
rect 47450 -32729 48006 -32695
rect 32180 -33457 32736 -33423
rect 33198 -33457 33754 -33423
rect 34216 -33457 34772 -33423
rect 35234 -33457 35790 -33423
rect 36252 -33457 36808 -33423
rect 37270 -33457 37826 -33423
rect 38288 -33457 38844 -33423
rect 39306 -33457 39862 -33423
rect 40324 -33457 40880 -33423
rect 41342 -33457 41898 -33423
rect 42360 -33457 42916 -33423
rect 43378 -33457 43934 -33423
rect 44396 -33457 44952 -33423
rect 45414 -33457 45970 -33423
rect 46432 -33457 46988 -33423
rect 47450 -33457 48006 -33423
rect 33374 -34367 33930 -34333
rect 34392 -34367 34948 -34333
rect 35410 -34367 35966 -34333
rect 36428 -34367 36984 -34333
rect 37446 -34367 38002 -34333
rect 38464 -34367 39020 -34333
rect 39482 -34367 40038 -34333
rect 40500 -34367 41056 -34333
rect 41518 -34367 42074 -34333
rect 42536 -34367 43092 -34333
rect 43554 -34367 44110 -34333
rect 44572 -34367 45128 -34333
rect 45590 -34367 46146 -34333
rect 46608 -34367 47164 -34333
rect 33374 -35095 33930 -35061
rect 34392 -35095 34948 -35061
rect 35410 -35095 35966 -35061
rect 36428 -35095 36984 -35061
rect 37446 -35095 38002 -35061
rect 38464 -35095 39020 -35061
rect 39482 -35095 40038 -35061
rect 40500 -35095 41056 -35061
rect 41518 -35095 42074 -35061
rect 42536 -35095 43092 -35061
rect 43554 -35095 44110 -35061
rect 44572 -35095 45128 -35061
rect 45590 -35095 46146 -35061
rect 46608 -35095 47164 -35061
rect 33374 -35399 33930 -35365
rect 34392 -35399 34948 -35365
rect 35410 -35399 35966 -35365
rect 36428 -35399 36984 -35365
rect 37446 -35399 38002 -35365
rect 38464 -35399 39020 -35365
rect 39482 -35399 40038 -35365
rect 40500 -35399 41056 -35365
rect 41518 -35399 42074 -35365
rect 42536 -35399 43092 -35365
rect 43554 -35399 44110 -35365
rect 44572 -35399 45128 -35365
rect 45590 -35399 46146 -35365
rect 46608 -35399 47164 -35365
rect 33374 -36127 33930 -36093
rect 34392 -36127 34948 -36093
rect 35410 -36127 35966 -36093
rect 36428 -36127 36984 -36093
rect 37446 -36127 38002 -36093
rect 38464 -36127 39020 -36093
rect 39482 -36127 40038 -36093
rect 40500 -36127 41056 -36093
rect 41518 -36127 42074 -36093
rect 42536 -36127 43092 -36093
rect 43554 -36127 44110 -36093
rect 44572 -36127 45128 -36093
rect 45590 -36127 46146 -36093
rect 46608 -36127 47164 -36093
rect 33166 -37003 33722 -36969
rect 34184 -37003 34740 -36969
rect 35202 -37003 35758 -36969
rect 36220 -37003 36776 -36969
rect 37238 -37003 37794 -36969
rect 38256 -37003 38812 -36969
rect 39274 -37003 39830 -36969
rect 40292 -37003 40848 -36969
rect 41310 -37003 41866 -36969
rect 42328 -37003 42884 -36969
rect 43346 -37003 43902 -36969
rect 44364 -37003 44920 -36969
rect 45382 -37003 45938 -36969
rect 46400 -37003 46956 -36969
rect 47418 -37003 47974 -36969
rect 27862 -37107 28418 -37073
rect 28880 -37107 29436 -37073
rect 29898 -37107 30454 -37073
rect 30916 -37107 31472 -37073
rect 33166 -37731 33722 -37697
rect 34184 -37731 34740 -37697
rect 35202 -37731 35758 -37697
rect 36220 -37731 36776 -37697
rect 37238 -37731 37794 -37697
rect 38256 -37731 38812 -37697
rect 39274 -37731 39830 -37697
rect 40292 -37731 40848 -37697
rect 41310 -37731 41866 -37697
rect 42328 -37731 42884 -37697
rect 43346 -37731 43902 -37697
rect 44364 -37731 44920 -37697
rect 45382 -37731 45938 -37697
rect 46400 -37731 46956 -37697
rect 47418 -37731 47974 -37697
rect 27862 -37835 28418 -37801
rect 28880 -37835 29436 -37801
rect 29898 -37835 30454 -37801
rect 30916 -37835 31472 -37801
rect 27862 -38139 28418 -38105
rect 28880 -38139 29436 -38105
rect 29898 -38139 30454 -38105
rect 30916 -38139 31472 -38105
rect 33166 -38259 33722 -38225
rect 34184 -38259 34740 -38225
rect 35202 -38259 35758 -38225
rect 36220 -38259 36776 -38225
rect 37238 -38259 37794 -38225
rect 38256 -38259 38812 -38225
rect 39274 -38259 39830 -38225
rect 40292 -38259 40848 -38225
rect 41310 -38259 41866 -38225
rect 42328 -38259 42884 -38225
rect 43346 -38259 43902 -38225
rect 44364 -38259 44920 -38225
rect 45382 -38259 45938 -38225
rect 46400 -38259 46956 -38225
rect 47418 -38259 47974 -38225
rect 27862 -38867 28418 -38833
rect 28880 -38867 29436 -38833
rect 29898 -38867 30454 -38833
rect 30916 -38867 31472 -38833
rect 33166 -38987 33722 -38953
rect 34184 -38987 34740 -38953
rect 35202 -38987 35758 -38953
rect 36220 -38987 36776 -38953
rect 37238 -38987 37794 -38953
rect 38256 -38987 38812 -38953
rect 39274 -38987 39830 -38953
rect 40292 -38987 40848 -38953
rect 41310 -38987 41866 -38953
rect 42328 -38987 42884 -38953
rect 43346 -38987 43902 -38953
rect 44364 -38987 44920 -38953
rect 45382 -38987 45938 -38953
rect 46400 -38987 46956 -38953
rect 47418 -38987 47974 -38953
rect 27862 -39171 28418 -39137
rect 28880 -39171 29436 -39137
rect 29898 -39171 30454 -39137
rect 30916 -39171 31472 -39137
rect 33166 -39515 33722 -39481
rect 34184 -39515 34740 -39481
rect 35202 -39515 35758 -39481
rect 36220 -39515 36776 -39481
rect 37238 -39515 37794 -39481
rect 38256 -39515 38812 -39481
rect 39274 -39515 39830 -39481
rect 40292 -39515 40848 -39481
rect 41310 -39515 41866 -39481
rect 42328 -39515 42884 -39481
rect 43346 -39515 43902 -39481
rect 44364 -39515 44920 -39481
rect 45382 -39515 45938 -39481
rect 46400 -39515 46956 -39481
rect 47418 -39515 47974 -39481
rect 27862 -39899 28418 -39865
rect 28880 -39899 29436 -39865
rect 29898 -39899 30454 -39865
rect 30916 -39899 31472 -39865
rect 27862 -40203 28418 -40169
rect 28880 -40203 29436 -40169
rect 29898 -40203 30454 -40169
rect 30916 -40203 31472 -40169
rect 33166 -40243 33722 -40209
rect 34184 -40243 34740 -40209
rect 35202 -40243 35758 -40209
rect 36220 -40243 36776 -40209
rect 37238 -40243 37794 -40209
rect 38256 -40243 38812 -40209
rect 39274 -40243 39830 -40209
rect 40292 -40243 40848 -40209
rect 41310 -40243 41866 -40209
rect 42328 -40243 42884 -40209
rect 43346 -40243 43902 -40209
rect 44364 -40243 44920 -40209
rect 45382 -40243 45938 -40209
rect 46400 -40243 46956 -40209
rect 47418 -40243 47974 -40209
rect 33166 -40771 33722 -40737
rect 34184 -40771 34740 -40737
rect 35202 -40771 35758 -40737
rect 36220 -40771 36776 -40737
rect 37238 -40771 37794 -40737
rect 38256 -40771 38812 -40737
rect 39274 -40771 39830 -40737
rect 40292 -40771 40848 -40737
rect 41310 -40771 41866 -40737
rect 42328 -40771 42884 -40737
rect 43346 -40771 43902 -40737
rect 44364 -40771 44920 -40737
rect 45382 -40771 45938 -40737
rect 46400 -40771 46956 -40737
rect 47418 -40771 47974 -40737
rect 27862 -40931 28418 -40897
rect 28880 -40931 29436 -40897
rect 29898 -40931 30454 -40897
rect 30916 -40931 31472 -40897
rect 33166 -41499 33722 -41465
rect 34184 -41499 34740 -41465
rect 35202 -41499 35758 -41465
rect 36220 -41499 36776 -41465
rect 37238 -41499 37794 -41465
rect 38256 -41499 38812 -41465
rect 39274 -41499 39830 -41465
rect 40292 -41499 40848 -41465
rect 41310 -41499 41866 -41465
rect 42328 -41499 42884 -41465
rect 43346 -41499 43902 -41465
rect 44364 -41499 44920 -41465
rect 45382 -41499 45938 -41465
rect 46400 -41499 46956 -41465
rect 47418 -41499 47974 -41465
rect 52578 -39633 52798 -39599
rect 53036 -39633 53256 -39599
rect 53494 -39633 53714 -39599
rect 53952 -39633 54172 -39599
rect 54410 -39633 54630 -39599
rect 54868 -39633 55088 -39599
rect 52578 -39961 52798 -39927
rect 53036 -39961 53256 -39927
rect 53494 -39961 53714 -39927
rect 53952 -39961 54172 -39927
rect 54410 -39961 54630 -39927
rect 54868 -39961 55088 -39927
rect 52597 -40516 52697 -40482
rect 52855 -40516 52955 -40482
rect 53113 -40516 53213 -40482
rect 53371 -40516 53471 -40482
rect 53629 -40516 53729 -40482
rect 53887 -40516 53987 -40482
rect 54145 -40516 54245 -40482
rect 54403 -40516 54503 -40482
rect 54661 -40516 54761 -40482
rect 54919 -40516 55019 -40482
rect 52597 -41044 52697 -41010
rect 52855 -41044 52955 -41010
rect 53113 -41044 53213 -41010
rect 53371 -41044 53471 -41010
rect 53629 -41044 53729 -41010
rect 53887 -41044 53987 -41010
rect 54145 -41044 54245 -41010
rect 54403 -41044 54503 -41010
rect 54661 -41044 54761 -41010
rect 54919 -41044 55019 -41010
rect 52597 -41376 52697 -41342
rect 52855 -41376 52955 -41342
rect 53113 -41376 53213 -41342
rect 53371 -41376 53471 -41342
rect 53629 -41376 53729 -41342
rect 53887 -41376 53987 -41342
rect 54145 -41376 54245 -41342
rect 54403 -41376 54503 -41342
rect 54661 -41376 54761 -41342
rect 54919 -41376 55019 -41342
rect 52597 -41904 52697 -41870
rect 52855 -41904 52955 -41870
rect 53113 -41904 53213 -41870
rect 53371 -41904 53471 -41870
rect 53629 -41904 53729 -41870
rect 53887 -41904 53987 -41870
rect 54145 -41904 54245 -41870
rect 54403 -41904 54503 -41870
rect 54661 -41904 54761 -41870
rect 54919 -41904 55019 -41870
rect 56166 -39833 56266 -39799
rect 56424 -39833 56524 -39799
rect 56682 -39833 56782 -39799
rect 56940 -39833 57040 -39799
rect 57198 -39833 57298 -39799
rect 57456 -39833 57556 -39799
rect 57714 -39833 57814 -39799
rect 56166 -40361 56266 -40327
rect 56424 -40361 56524 -40327
rect 56682 -40361 56782 -40327
rect 56940 -40361 57040 -40327
rect 57198 -40361 57298 -40327
rect 57456 -40361 57556 -40327
rect 57714 -40361 57814 -40327
rect 56166 -40693 56266 -40659
rect 56424 -40693 56524 -40659
rect 56682 -40693 56782 -40659
rect 56940 -40693 57040 -40659
rect 57198 -40693 57298 -40659
rect 57456 -40693 57556 -40659
rect 57714 -40693 57814 -40659
rect 56166 -41221 56266 -41187
rect 56424 -41221 56524 -41187
rect 56682 -41221 56782 -41187
rect 56940 -41221 57040 -41187
rect 57198 -41221 57298 -41187
rect 57456 -41221 57556 -41187
rect 57714 -41221 57814 -41187
rect 56184 -41921 56218 -41887
rect 56460 -41921 56494 -41887
rect 56692 -41921 56726 -41887
rect 56860 -41921 56894 -41887
rect 57156 -41921 57190 -41887
rect 57324 -41921 57358 -41887
rect 57556 -41921 57590 -41887
rect 57832 -41921 57866 -41887
rect 54402 -42537 54452 -42487
rect 54530 -42537 54580 -42487
rect 54658 -42537 54708 -42487
rect 54786 -42537 54836 -42487
rect 54914 -42537 54964 -42487
rect 55042 -42537 55092 -42487
rect 55170 -42537 55220 -42487
rect 54274 -42899 54324 -42849
rect 55298 -42899 55348 -42849
rect 56075 -42664 56109 -42630
rect 56736 -42552 56776 -42512
rect 56972 -42552 57012 -42512
rect 57090 -42552 57130 -42512
rect 57326 -42552 57366 -42512
rect 56558 -42916 56598 -42876
rect 56854 -42918 56894 -42878
rect 57208 -42918 57248 -42878
rect 57506 -42916 57546 -42876
rect 10506 -56875 10606 -56841
rect 10764 -56875 10864 -56841
rect 11022 -56875 11122 -56841
rect 11280 -56875 11380 -56841
rect 11538 -56875 11638 -56841
rect 11796 -56875 11896 -56841
rect 10506 -57403 10606 -57369
rect 10764 -57403 10864 -57369
rect 11022 -57403 11122 -57369
rect 11280 -57403 11380 -57369
rect 11538 -57403 11638 -57369
rect 11796 -57403 11896 -57369
rect 12342 -57587 12376 -57553
rect 10506 -57808 10606 -57774
rect 10764 -57808 10864 -57774
rect 11022 -57808 11122 -57774
rect 11280 -57808 11380 -57774
rect 11538 -57808 11638 -57774
rect 11796 -57808 11896 -57774
rect 10506 -58118 10606 -58084
rect 10764 -58118 10864 -58084
rect 11022 -58118 11122 -58084
rect 11280 -58118 11380 -58084
rect 11538 -58118 11638 -58084
rect 11796 -58118 11896 -58084
rect 28274 -43976 28830 -43942
rect 29292 -43976 29848 -43942
rect 30310 -43976 30866 -43942
rect 31328 -43976 31884 -43942
rect 32346 -43976 32902 -43942
rect 33364 -43976 33920 -43942
rect 34382 -43976 34938 -43942
rect 35400 -43976 35956 -43942
rect 36418 -43976 36974 -43942
rect 37436 -43976 37992 -43942
rect 38454 -43976 39010 -43942
rect 39472 -43976 40028 -43942
rect 40490 -43976 41046 -43942
rect 41508 -43976 42064 -43942
rect 42526 -43976 43082 -43942
rect 43544 -43976 44100 -43942
rect 44562 -43976 45118 -43942
rect 45580 -43976 46136 -43942
rect 46598 -43976 47154 -43942
rect 47616 -43976 48172 -43942
rect 16508 -44452 17064 -44418
rect 17526 -44452 18082 -44418
rect 18544 -44452 19100 -44418
rect 19562 -44452 20118 -44418
rect 20580 -44452 21136 -44418
rect 21598 -44452 22154 -44418
rect 22616 -44452 23172 -44418
rect 23634 -44452 24190 -44418
rect 24652 -44452 25208 -44418
rect 28274 -44686 28830 -44652
rect 29292 -44686 29848 -44652
rect 30310 -44686 30866 -44652
rect 31328 -44686 31884 -44652
rect 32346 -44686 32902 -44652
rect 33364 -44686 33920 -44652
rect 34382 -44686 34938 -44652
rect 35400 -44686 35956 -44652
rect 36418 -44686 36974 -44652
rect 37436 -44686 37992 -44652
rect 38454 -44686 39010 -44652
rect 39472 -44686 40028 -44652
rect 40490 -44686 41046 -44652
rect 41508 -44686 42064 -44652
rect 42526 -44686 43082 -44652
rect 43544 -44686 44100 -44652
rect 44562 -44686 45118 -44652
rect 45580 -44686 46136 -44652
rect 46598 -44686 47154 -44652
rect 47616 -44686 48172 -44652
rect 28274 -44794 28830 -44760
rect 29292 -44794 29848 -44760
rect 30310 -44794 30866 -44760
rect 31328 -44794 31884 -44760
rect 32346 -44794 32902 -44760
rect 33364 -44794 33920 -44760
rect 34382 -44794 34938 -44760
rect 35400 -44794 35956 -44760
rect 36418 -44794 36974 -44760
rect 37436 -44794 37992 -44760
rect 38454 -44794 39010 -44760
rect 39472 -44794 40028 -44760
rect 40490 -44794 41046 -44760
rect 41508 -44794 42064 -44760
rect 42526 -44794 43082 -44760
rect 43544 -44794 44100 -44760
rect 44562 -44794 45118 -44760
rect 45580 -44794 46136 -44760
rect 46598 -44794 47154 -44760
rect 47616 -44794 48172 -44760
rect 16508 -45162 17064 -45128
rect 17526 -45162 18082 -45128
rect 16508 -45270 17064 -45236
rect 18544 -45162 19100 -45128
rect 17526 -45270 18082 -45236
rect 19562 -45162 20118 -45128
rect 18544 -45270 19100 -45236
rect 20580 -45162 21136 -45128
rect 19562 -45270 20118 -45236
rect 21598 -45162 22154 -45128
rect 20580 -45270 21136 -45236
rect 22616 -45162 23172 -45128
rect 21598 -45270 22154 -45236
rect 23634 -45162 24190 -45128
rect 22616 -45270 23172 -45236
rect 24652 -45162 25208 -45128
rect 23634 -45270 24190 -45236
rect 24652 -45270 25208 -45236
rect 28274 -45504 28830 -45470
rect 29292 -45504 29848 -45470
rect 30310 -45504 30866 -45470
rect 31328 -45504 31884 -45470
rect 32346 -45504 32902 -45470
rect 33364 -45504 33920 -45470
rect 34382 -45504 34938 -45470
rect 35400 -45504 35956 -45470
rect 36418 -45504 36974 -45470
rect 37436 -45504 37992 -45470
rect 38454 -45504 39010 -45470
rect 39472 -45504 40028 -45470
rect 40490 -45504 41046 -45470
rect 41508 -45504 42064 -45470
rect 42526 -45504 43082 -45470
rect 43544 -45504 44100 -45470
rect 44562 -45504 45118 -45470
rect 45580 -45504 46136 -45470
rect 46598 -45504 47154 -45470
rect 47616 -45504 48172 -45470
rect 16508 -45980 17064 -45946
rect 17526 -45980 18082 -45946
rect 16508 -46088 17064 -46054
rect 18544 -45980 19100 -45946
rect 17526 -46088 18082 -46054
rect 19562 -45980 20118 -45946
rect 18544 -46088 19100 -46054
rect 20580 -45980 21136 -45946
rect 19562 -46088 20118 -46054
rect 21598 -45980 22154 -45946
rect 20580 -46088 21136 -46054
rect 22616 -45980 23172 -45946
rect 21598 -46088 22154 -46054
rect 23634 -45980 24190 -45946
rect 22616 -46088 23172 -46054
rect 24652 -45980 25208 -45946
rect 23634 -46088 24190 -46054
rect 24652 -46088 25208 -46054
rect 28274 -46172 28830 -46138
rect 29292 -46172 29848 -46138
rect 30310 -46172 30866 -46138
rect 31328 -46172 31884 -46138
rect 32346 -46172 32902 -46138
rect 33364 -46172 33920 -46138
rect 34382 -46172 34938 -46138
rect 35400 -46172 35956 -46138
rect 36418 -46172 36974 -46138
rect 37436 -46172 37992 -46138
rect 38454 -46172 39010 -46138
rect 39472 -46172 40028 -46138
rect 40490 -46172 41046 -46138
rect 41508 -46172 42064 -46138
rect 42526 -46172 43082 -46138
rect 43544 -46172 44100 -46138
rect 44562 -46172 45118 -46138
rect 45580 -46172 46136 -46138
rect 46598 -46172 47154 -46138
rect 47616 -46172 48172 -46138
rect 16508 -46798 17064 -46764
rect 17526 -46798 18082 -46764
rect 16508 -46906 17064 -46872
rect 18544 -46798 19100 -46764
rect 17526 -46906 18082 -46872
rect 19562 -46798 20118 -46764
rect 18544 -46906 19100 -46872
rect 20580 -46798 21136 -46764
rect 19562 -46906 20118 -46872
rect 21598 -46798 22154 -46764
rect 20580 -46906 21136 -46872
rect 22616 -46798 23172 -46764
rect 21598 -46906 22154 -46872
rect 23634 -46798 24190 -46764
rect 22616 -46906 23172 -46872
rect 24652 -46798 25208 -46764
rect 23634 -46906 24190 -46872
rect 24652 -46906 25208 -46872
rect 28274 -46882 28830 -46848
rect 29292 -46882 29848 -46848
rect 30310 -46882 30866 -46848
rect 31328 -46882 31884 -46848
rect 32346 -46882 32902 -46848
rect 33364 -46882 33920 -46848
rect 34382 -46882 34938 -46848
rect 35400 -46882 35956 -46848
rect 36418 -46882 36974 -46848
rect 37436 -46882 37992 -46848
rect 38454 -46882 39010 -46848
rect 39472 -46882 40028 -46848
rect 40490 -46882 41046 -46848
rect 41508 -46882 42064 -46848
rect 42526 -46882 43082 -46848
rect 43544 -46882 44100 -46848
rect 44562 -46882 45118 -46848
rect 45580 -46882 46136 -46848
rect 46598 -46882 47154 -46848
rect 47616 -46882 48172 -46848
rect 28274 -47404 28830 -47370
rect 29292 -47404 29848 -47370
rect 30310 -47404 30866 -47370
rect 31328 -47404 31884 -47370
rect 32346 -47404 32902 -47370
rect 33364 -47404 33920 -47370
rect 34382 -47404 34938 -47370
rect 35400 -47404 35956 -47370
rect 36418 -47404 36974 -47370
rect 37436 -47404 37992 -47370
rect 38454 -47404 39010 -47370
rect 39472 -47404 40028 -47370
rect 40490 -47404 41046 -47370
rect 41508 -47404 42064 -47370
rect 42526 -47404 43082 -47370
rect 43544 -47404 44100 -47370
rect 44562 -47404 45118 -47370
rect 45580 -47404 46136 -47370
rect 46598 -47404 47154 -47370
rect 47616 -47404 48172 -47370
rect 16508 -47616 17064 -47582
rect 17526 -47616 18082 -47582
rect 16508 -47724 17064 -47690
rect 18544 -47616 19100 -47582
rect 17526 -47724 18082 -47690
rect 19562 -47616 20118 -47582
rect 18544 -47724 19100 -47690
rect 20580 -47616 21136 -47582
rect 19562 -47724 20118 -47690
rect 21598 -47616 22154 -47582
rect 20580 -47724 21136 -47690
rect 22616 -47616 23172 -47582
rect 21598 -47724 22154 -47690
rect 23634 -47616 24190 -47582
rect 22616 -47724 23172 -47690
rect 24652 -47616 25208 -47582
rect 23634 -47724 24190 -47690
rect 24652 -47724 25208 -47690
rect 28274 -48114 28830 -48080
rect 29292 -48114 29848 -48080
rect 30310 -48114 30866 -48080
rect 31328 -48114 31884 -48080
rect 32346 -48114 32902 -48080
rect 33364 -48114 33920 -48080
rect 34382 -48114 34938 -48080
rect 35400 -48114 35956 -48080
rect 36418 -48114 36974 -48080
rect 37436 -48114 37992 -48080
rect 38454 -48114 39010 -48080
rect 39472 -48114 40028 -48080
rect 40490 -48114 41046 -48080
rect 41508 -48114 42064 -48080
rect 42526 -48114 43082 -48080
rect 43544 -48114 44100 -48080
rect 44562 -48114 45118 -48080
rect 45580 -48114 46136 -48080
rect 46598 -48114 47154 -48080
rect 47616 -48114 48172 -48080
rect 16508 -48434 17064 -48400
rect 17526 -48434 18082 -48400
rect 16508 -48542 17064 -48508
rect 18544 -48434 19100 -48400
rect 17526 -48542 18082 -48508
rect 19562 -48434 20118 -48400
rect 18544 -48542 19100 -48508
rect 20580 -48434 21136 -48400
rect 19562 -48542 20118 -48508
rect 21598 -48434 22154 -48400
rect 20580 -48542 21136 -48508
rect 22616 -48434 23172 -48400
rect 21598 -48542 22154 -48508
rect 23634 -48434 24190 -48400
rect 22616 -48542 23172 -48508
rect 24652 -48434 25208 -48400
rect 23634 -48542 24190 -48508
rect 24652 -48542 25208 -48508
rect 28272 -48638 28828 -48604
rect 29290 -48638 29846 -48604
rect 30308 -48638 30864 -48604
rect 31326 -48638 31882 -48604
rect 32344 -48638 32900 -48604
rect 33362 -48638 33918 -48604
rect 34380 -48638 34936 -48604
rect 35398 -48638 35954 -48604
rect 36416 -48638 36972 -48604
rect 37434 -48638 37990 -48604
rect 38452 -48638 39008 -48604
rect 39470 -48638 40026 -48604
rect 40488 -48638 41044 -48604
rect 41506 -48638 42062 -48604
rect 42524 -48638 43080 -48604
rect 43542 -48638 44098 -48604
rect 44560 -48638 45116 -48604
rect 45578 -48638 46134 -48604
rect 46596 -48638 47152 -48604
rect 47614 -48638 48170 -48604
rect 16508 -49252 17064 -49218
rect 17526 -49252 18082 -49218
rect 16508 -49360 17064 -49326
rect 18544 -49252 19100 -49218
rect 17526 -49360 18082 -49326
rect 19562 -49252 20118 -49218
rect 18544 -49360 19100 -49326
rect 20580 -49252 21136 -49218
rect 19562 -49360 20118 -49326
rect 21598 -49252 22154 -49218
rect 20580 -49360 21136 -49326
rect 22616 -49252 23172 -49218
rect 21598 -49360 22154 -49326
rect 23634 -49252 24190 -49218
rect 22616 -49360 23172 -49326
rect 24652 -49252 25208 -49218
rect 23634 -49360 24190 -49326
rect 24652 -49360 25208 -49326
rect 28272 -49348 28828 -49314
rect 29290 -49348 29846 -49314
rect 30308 -49348 30864 -49314
rect 31326 -49348 31882 -49314
rect 32344 -49348 32900 -49314
rect 33362 -49348 33918 -49314
rect 34380 -49348 34936 -49314
rect 35398 -49348 35954 -49314
rect 36416 -49348 36972 -49314
rect 37434 -49348 37990 -49314
rect 38452 -49348 39008 -49314
rect 39470 -49348 40026 -49314
rect 40488 -49348 41044 -49314
rect 41506 -49348 42062 -49314
rect 42524 -49348 43080 -49314
rect 43542 -49348 44098 -49314
rect 44560 -49348 45116 -49314
rect 45578 -49348 46134 -49314
rect 46596 -49348 47152 -49314
rect 47614 -49348 48170 -49314
rect 28272 -49872 28828 -49838
rect 29290 -49872 29846 -49838
rect 30308 -49872 30864 -49838
rect 31326 -49872 31882 -49838
rect 32344 -49872 32900 -49838
rect 33362 -49872 33918 -49838
rect 34380 -49872 34936 -49838
rect 35398 -49872 35954 -49838
rect 36416 -49872 36972 -49838
rect 37434 -49872 37990 -49838
rect 38452 -49872 39008 -49838
rect 39470 -49872 40026 -49838
rect 40488 -49872 41044 -49838
rect 41506 -49872 42062 -49838
rect 42524 -49872 43080 -49838
rect 43542 -49872 44098 -49838
rect 44560 -49872 45116 -49838
rect 45578 -49872 46134 -49838
rect 46596 -49872 47152 -49838
rect 47614 -49872 48170 -49838
rect 16508 -50070 17064 -50036
rect 17526 -50070 18082 -50036
rect 16508 -50178 17064 -50144
rect 18544 -50070 19100 -50036
rect 17526 -50178 18082 -50144
rect 19562 -50070 20118 -50036
rect 18544 -50178 19100 -50144
rect 20580 -50070 21136 -50036
rect 19562 -50178 20118 -50144
rect 21598 -50070 22154 -50036
rect 20580 -50178 21136 -50144
rect 22616 -50070 23172 -50036
rect 21598 -50178 22154 -50144
rect 23634 -50070 24190 -50036
rect 22616 -50178 23172 -50144
rect 24652 -50070 25208 -50036
rect 23634 -50178 24190 -50144
rect 24652 -50178 25208 -50144
rect 28272 -50582 28828 -50548
rect 29290 -50582 29846 -50548
rect 30308 -50582 30864 -50548
rect 31326 -50582 31882 -50548
rect 32344 -50582 32900 -50548
rect 33362 -50582 33918 -50548
rect 34380 -50582 34936 -50548
rect 35398 -50582 35954 -50548
rect 36416 -50582 36972 -50548
rect 37434 -50582 37990 -50548
rect 38452 -50582 39008 -50548
rect 39470 -50582 40026 -50548
rect 40488 -50582 41044 -50548
rect 41506 -50582 42062 -50548
rect 42524 -50582 43080 -50548
rect 43542 -50582 44098 -50548
rect 44560 -50582 45116 -50548
rect 45578 -50582 46134 -50548
rect 46596 -50582 47152 -50548
rect 47614 -50582 48170 -50548
rect 16508 -50888 17064 -50854
rect 17526 -50888 18082 -50854
rect 18544 -50888 19100 -50854
rect 19562 -50888 20118 -50854
rect 20580 -50888 21136 -50854
rect 21598 -50888 22154 -50854
rect 22616 -50888 23172 -50854
rect 23634 -50888 24190 -50854
rect 24652 -50888 25208 -50854
rect 28272 -51104 28828 -51070
rect 29290 -51104 29846 -51070
rect 30308 -51104 30864 -51070
rect 31326 -51104 31882 -51070
rect 32344 -51104 32900 -51070
rect 33362 -51104 33918 -51070
rect 34380 -51104 34936 -51070
rect 35398 -51104 35954 -51070
rect 36416 -51104 36972 -51070
rect 37434 -51104 37990 -51070
rect 38452 -51104 39008 -51070
rect 39470 -51104 40026 -51070
rect 40488 -51104 41044 -51070
rect 41506 -51104 42062 -51070
rect 42524 -51104 43080 -51070
rect 43542 -51104 44098 -51070
rect 44560 -51104 45116 -51070
rect 45578 -51104 46134 -51070
rect 46596 -51104 47152 -51070
rect 47614 -51104 48170 -51070
rect 28272 -51814 28828 -51780
rect 29290 -51814 29846 -51780
rect 30308 -51814 30864 -51780
rect 31326 -51814 31882 -51780
rect 32344 -51814 32900 -51780
rect 33362 -51814 33918 -51780
rect 34380 -51814 34936 -51780
rect 35398 -51814 35954 -51780
rect 36416 -51814 36972 -51780
rect 37434 -51814 37990 -51780
rect 38452 -51814 39008 -51780
rect 39470 -51814 40026 -51780
rect 40488 -51814 41044 -51780
rect 41506 -51814 42062 -51780
rect 42524 -51814 43080 -51780
rect 43542 -51814 44098 -51780
rect 44560 -51814 45116 -51780
rect 45578 -51814 46134 -51780
rect 46596 -51814 47152 -51780
rect 47614 -51814 48170 -51780
rect 15184 -52202 15740 -52168
rect 16202 -52202 16758 -52168
rect 17220 -52202 17776 -52168
rect 18238 -52202 18794 -52168
rect 19256 -52202 19812 -52168
rect 20274 -52202 20830 -52168
rect 21292 -52202 21848 -52168
rect 22310 -52202 22866 -52168
rect 23328 -52202 23884 -52168
rect 24346 -52202 24902 -52168
rect 25364 -52202 25920 -52168
rect 28272 -52338 28828 -52304
rect 29290 -52338 29846 -52304
rect 30308 -52338 30864 -52304
rect 31326 -52338 31882 -52304
rect 32344 -52338 32900 -52304
rect 33362 -52338 33918 -52304
rect 34380 -52338 34936 -52304
rect 35398 -52338 35954 -52304
rect 36416 -52338 36972 -52304
rect 37434 -52338 37990 -52304
rect 38452 -52338 39008 -52304
rect 39470 -52338 40026 -52304
rect 40488 -52338 41044 -52304
rect 41506 -52338 42062 -52304
rect 42524 -52338 43080 -52304
rect 43542 -52338 44098 -52304
rect 44560 -52338 45116 -52304
rect 45578 -52338 46134 -52304
rect 46596 -52338 47152 -52304
rect 47614 -52338 48170 -52304
rect 15184 -52912 15740 -52878
rect 16202 -52912 16758 -52878
rect 17220 -52912 17776 -52878
rect 18238 -52912 18794 -52878
rect 19256 -52912 19812 -52878
rect 20274 -52912 20830 -52878
rect 21292 -52912 21848 -52878
rect 22310 -52912 22866 -52878
rect 23328 -52912 23884 -52878
rect 24346 -52912 24902 -52878
rect 25364 -52912 25920 -52878
rect 28272 -53048 28828 -53014
rect 29290 -53048 29846 -53014
rect 30308 -53048 30864 -53014
rect 31326 -53048 31882 -53014
rect 32344 -53048 32900 -53014
rect 33362 -53048 33918 -53014
rect 34380 -53048 34936 -53014
rect 35398 -53048 35954 -53014
rect 36416 -53048 36972 -53014
rect 37434 -53048 37990 -53014
rect 38452 -53048 39008 -53014
rect 39470 -53048 40026 -53014
rect 40488 -53048 41044 -53014
rect 41506 -53048 42062 -53014
rect 42524 -53048 43080 -53014
rect 43542 -53048 44098 -53014
rect 44560 -53048 45116 -53014
rect 45578 -53048 46134 -53014
rect 46596 -53048 47152 -53014
rect 47614 -53048 48170 -53014
rect 15184 -53314 15740 -53280
rect 16202 -53314 16758 -53280
rect 17220 -53314 17776 -53280
rect 18238 -53314 18794 -53280
rect 19256 -53314 19812 -53280
rect 20274 -53314 20830 -53280
rect 21292 -53314 21848 -53280
rect 22310 -53314 22866 -53280
rect 23328 -53314 23884 -53280
rect 24346 -53314 24902 -53280
rect 25364 -53314 25920 -53280
rect 28272 -53572 28828 -53538
rect 29290 -53572 29846 -53538
rect 30308 -53572 30864 -53538
rect 31326 -53572 31882 -53538
rect 32344 -53572 32900 -53538
rect 33362 -53572 33918 -53538
rect 34380 -53572 34936 -53538
rect 35398 -53572 35954 -53538
rect 36416 -53572 36972 -53538
rect 37434 -53572 37990 -53538
rect 38452 -53572 39008 -53538
rect 39470 -53572 40026 -53538
rect 40488 -53572 41044 -53538
rect 41506 -53572 42062 -53538
rect 42524 -53572 43080 -53538
rect 43542 -53572 44098 -53538
rect 44560 -53572 45116 -53538
rect 45578 -53572 46134 -53538
rect 46596 -53572 47152 -53538
rect 47614 -53572 48170 -53538
rect 15184 -54024 15740 -53990
rect 16202 -54024 16758 -53990
rect 17220 -54024 17776 -53990
rect 18238 -54024 18794 -53990
rect 19256 -54024 19812 -53990
rect 20274 -54024 20830 -53990
rect 21292 -54024 21848 -53990
rect 22310 -54024 22866 -53990
rect 23328 -54024 23884 -53990
rect 24346 -54024 24902 -53990
rect 25364 -54024 25920 -53990
rect 28272 -54282 28828 -54248
rect 29290 -54282 29846 -54248
rect 30308 -54282 30864 -54248
rect 31326 -54282 31882 -54248
rect 32344 -54282 32900 -54248
rect 33362 -54282 33918 -54248
rect 34380 -54282 34936 -54248
rect 35398 -54282 35954 -54248
rect 36416 -54282 36972 -54248
rect 37434 -54282 37990 -54248
rect 38452 -54282 39008 -54248
rect 39470 -54282 40026 -54248
rect 40488 -54282 41044 -54248
rect 41506 -54282 42062 -54248
rect 42524 -54282 43080 -54248
rect 43542 -54282 44098 -54248
rect 44560 -54282 45116 -54248
rect 45578 -54282 46134 -54248
rect 46596 -54282 47152 -54248
rect 47614 -54282 48170 -54248
rect 15184 -54426 15740 -54392
rect 16202 -54426 16758 -54392
rect 17220 -54426 17776 -54392
rect 18238 -54426 18794 -54392
rect 19256 -54426 19812 -54392
rect 20274 -54426 20830 -54392
rect 21292 -54426 21848 -54392
rect 22310 -54426 22866 -54392
rect 23328 -54426 23884 -54392
rect 24346 -54426 24902 -54392
rect 25364 -54426 25920 -54392
rect 28272 -54804 28828 -54770
rect 29290 -54804 29846 -54770
rect 30308 -54804 30864 -54770
rect 31326 -54804 31882 -54770
rect 32344 -54804 32900 -54770
rect 33362 -54804 33918 -54770
rect 34380 -54804 34936 -54770
rect 35398 -54804 35954 -54770
rect 36416 -54804 36972 -54770
rect 37434 -54804 37990 -54770
rect 38452 -54804 39008 -54770
rect 39470 -54804 40026 -54770
rect 40488 -54804 41044 -54770
rect 41506 -54804 42062 -54770
rect 42524 -54804 43080 -54770
rect 43542 -54804 44098 -54770
rect 44560 -54804 45116 -54770
rect 45578 -54804 46134 -54770
rect 46596 -54804 47152 -54770
rect 47614 -54804 48170 -54770
rect 15184 -55136 15740 -55102
rect 16202 -55136 16758 -55102
rect 17220 -55136 17776 -55102
rect 18238 -55136 18794 -55102
rect 19256 -55136 19812 -55102
rect 20274 -55136 20830 -55102
rect 21292 -55136 21848 -55102
rect 22310 -55136 22866 -55102
rect 23328 -55136 23884 -55102
rect 24346 -55136 24902 -55102
rect 25364 -55136 25920 -55102
rect 15184 -55538 15740 -55504
rect 16202 -55538 16758 -55504
rect 17220 -55538 17776 -55504
rect 18238 -55538 18794 -55504
rect 19256 -55538 19812 -55504
rect 20274 -55538 20830 -55504
rect 21292 -55538 21848 -55504
rect 22310 -55538 22866 -55504
rect 23328 -55538 23884 -55504
rect 24346 -55538 24902 -55504
rect 25364 -55538 25920 -55504
rect 28272 -55514 28828 -55480
rect 29290 -55514 29846 -55480
rect 30308 -55514 30864 -55480
rect 31326 -55514 31882 -55480
rect 32344 -55514 32900 -55480
rect 33362 -55514 33918 -55480
rect 34380 -55514 34936 -55480
rect 35398 -55514 35954 -55480
rect 36416 -55514 36972 -55480
rect 37434 -55514 37990 -55480
rect 38452 -55514 39008 -55480
rect 39470 -55514 40026 -55480
rect 40488 -55514 41044 -55480
rect 41506 -55514 42062 -55480
rect 42524 -55514 43080 -55480
rect 43542 -55514 44098 -55480
rect 44560 -55514 45116 -55480
rect 45578 -55514 46134 -55480
rect 46596 -55514 47152 -55480
rect 47614 -55514 48170 -55480
rect 28272 -56038 28828 -56004
rect 29290 -56038 29846 -56004
rect 30308 -56038 30864 -56004
rect 31326 -56038 31882 -56004
rect 32344 -56038 32900 -56004
rect 33362 -56038 33918 -56004
rect 34380 -56038 34936 -56004
rect 35398 -56038 35954 -56004
rect 36416 -56038 36972 -56004
rect 37434 -56038 37990 -56004
rect 38452 -56038 39008 -56004
rect 39470 -56038 40026 -56004
rect 40488 -56038 41044 -56004
rect 41506 -56038 42062 -56004
rect 42524 -56038 43080 -56004
rect 43542 -56038 44098 -56004
rect 44560 -56038 45116 -56004
rect 45578 -56038 46134 -56004
rect 46596 -56038 47152 -56004
rect 47614 -56038 48170 -56004
rect 15184 -56248 15740 -56214
rect 16202 -56248 16758 -56214
rect 17220 -56248 17776 -56214
rect 18238 -56248 18794 -56214
rect 19256 -56248 19812 -56214
rect 20274 -56248 20830 -56214
rect 21292 -56248 21848 -56214
rect 22310 -56248 22866 -56214
rect 23328 -56248 23884 -56214
rect 24346 -56248 24902 -56214
rect 25364 -56248 25920 -56214
rect 28272 -56748 28828 -56714
rect 29290 -56748 29846 -56714
rect 30308 -56748 30864 -56714
rect 31326 -56748 31882 -56714
rect 32344 -56748 32900 -56714
rect 33362 -56748 33918 -56714
rect 34380 -56748 34936 -56714
rect 35398 -56748 35954 -56714
rect 36416 -56748 36972 -56714
rect 37434 -56748 37990 -56714
rect 38452 -56748 39008 -56714
rect 39470 -56748 40026 -56714
rect 40488 -56748 41044 -56714
rect 41506 -56748 42062 -56714
rect 42524 -56748 43080 -56714
rect 43542 -56748 44098 -56714
rect 44560 -56748 45116 -56714
rect 45578 -56748 46134 -56714
rect 46596 -56748 47152 -56714
rect 47614 -56748 48170 -56714
rect 15642 -57080 16198 -57046
rect 16660 -57080 17216 -57046
rect 17678 -57080 18234 -57046
rect 18696 -57080 19252 -57046
rect 19714 -57080 20270 -57046
rect 20732 -57080 21288 -57046
rect 21750 -57080 22306 -57046
rect 22768 -57080 23324 -57046
rect 23786 -57080 24342 -57046
rect 24804 -57080 25360 -57046
rect 28272 -57270 28828 -57236
rect 29290 -57270 29846 -57236
rect 30308 -57270 30864 -57236
rect 31326 -57270 31882 -57236
rect 32344 -57270 32900 -57236
rect 33362 -57270 33918 -57236
rect 34380 -57270 34936 -57236
rect 35398 -57270 35954 -57236
rect 36416 -57270 36972 -57236
rect 37434 -57270 37990 -57236
rect 38452 -57270 39008 -57236
rect 39470 -57270 40026 -57236
rect 40488 -57270 41044 -57236
rect 41506 -57270 42062 -57236
rect 42524 -57270 43080 -57236
rect 43542 -57270 44098 -57236
rect 44560 -57270 45116 -57236
rect 45578 -57270 46134 -57236
rect 46596 -57270 47152 -57236
rect 47614 -57270 48170 -57236
rect 15642 -57790 16198 -57756
rect 16660 -57790 17216 -57756
rect 17678 -57790 18234 -57756
rect 18696 -57790 19252 -57756
rect 19714 -57790 20270 -57756
rect 20732 -57790 21288 -57756
rect 21750 -57790 22306 -57756
rect 22768 -57790 23324 -57756
rect 23786 -57790 24342 -57756
rect 24804 -57790 25360 -57756
rect 28272 -57980 28828 -57946
rect 29290 -57980 29846 -57946
rect 30308 -57980 30864 -57946
rect 31326 -57980 31882 -57946
rect 32344 -57980 32900 -57946
rect 33362 -57980 33918 -57946
rect 34380 -57980 34936 -57946
rect 35398 -57980 35954 -57946
rect 36416 -57980 36972 -57946
rect 37434 -57980 37990 -57946
rect 38452 -57980 39008 -57946
rect 39470 -57980 40026 -57946
rect 40488 -57980 41044 -57946
rect 41506 -57980 42062 -57946
rect 42524 -57980 43080 -57946
rect 43542 -57980 44098 -57946
rect 44560 -57980 45116 -57946
rect 45578 -57980 46134 -57946
rect 46596 -57980 47152 -57946
rect 47614 -57980 48170 -57946
rect 57979 -42664 58013 -42630
rect -27241 -65578 -27141 -65544
rect -26983 -65578 -26883 -65544
rect -26725 -65578 -26625 -65544
rect -26467 -65578 -26367 -65544
rect -26209 -65578 -26109 -65544
rect -25951 -65578 -25851 -65544
rect -27241 -66106 -27141 -66072
rect -26983 -66106 -26883 -66072
rect -26725 -66106 -26625 -66072
rect -26467 -66106 -26367 -66072
rect -26209 -66106 -26109 -66072
rect -25951 -66106 -25851 -66072
rect -27241 -66438 -27141 -66404
rect -26983 -66438 -26883 -66404
rect -26725 -66438 -26625 -66404
rect -26467 -66438 -26367 -66404
rect -26209 -66438 -26109 -66404
rect -25951 -66438 -25851 -66404
rect -27241 -66966 -27141 -66932
rect -26983 -66966 -26883 -66932
rect -26725 -66966 -26625 -66932
rect -26467 -66966 -26367 -66932
rect -26209 -66966 -26109 -66932
rect -25951 -66966 -25851 -66932
rect -23241 -65578 -23141 -65544
rect -22983 -65578 -22883 -65544
rect -22725 -65578 -22625 -65544
rect -22467 -65578 -22367 -65544
rect -22209 -65578 -22109 -65544
rect -21951 -65578 -21851 -65544
rect -23241 -66106 -23141 -66072
rect -22983 -66106 -22883 -66072
rect -22725 -66106 -22625 -66072
rect -22467 -66106 -22367 -66072
rect -22209 -66106 -22109 -66072
rect -21951 -66106 -21851 -66072
rect -23241 -66438 -23141 -66404
rect -22983 -66438 -22883 -66404
rect -22725 -66438 -22625 -66404
rect -22467 -66438 -22367 -66404
rect -22209 -66438 -22109 -66404
rect -21951 -66438 -21851 -66404
rect -23241 -66966 -23141 -66932
rect -22983 -66966 -22883 -66932
rect -22725 -66966 -22625 -66932
rect -22467 -66966 -22367 -66932
rect -22209 -66966 -22109 -66932
rect -21951 -66966 -21851 -66932
rect -19241 -65578 -19141 -65544
rect -18983 -65578 -18883 -65544
rect -18725 -65578 -18625 -65544
rect -18467 -65578 -18367 -65544
rect -18209 -65578 -18109 -65544
rect -17951 -65578 -17851 -65544
rect -19241 -66106 -19141 -66072
rect -18983 -66106 -18883 -66072
rect -18725 -66106 -18625 -66072
rect -18467 -66106 -18367 -66072
rect -18209 -66106 -18109 -66072
rect -17951 -66106 -17851 -66072
rect -19241 -66438 -19141 -66404
rect -18983 -66438 -18883 -66404
rect -18725 -66438 -18625 -66404
rect -18467 -66438 -18367 -66404
rect -18209 -66438 -18109 -66404
rect -17951 -66438 -17851 -66404
rect -19241 -66966 -19141 -66932
rect -18983 -66966 -18883 -66932
rect -18725 -66966 -18625 -66932
rect -18467 -66966 -18367 -66932
rect -18209 -66966 -18109 -66932
rect -17951 -66966 -17851 -66932
rect -15241 -65578 -15141 -65544
rect -14983 -65578 -14883 -65544
rect -14725 -65578 -14625 -65544
rect -14467 -65578 -14367 -65544
rect -14209 -65578 -14109 -65544
rect -13951 -65578 -13851 -65544
rect -15241 -66106 -15141 -66072
rect -14983 -66106 -14883 -66072
rect -14725 -66106 -14625 -66072
rect -14467 -66106 -14367 -66072
rect -14209 -66106 -14109 -66072
rect -13951 -66106 -13851 -66072
rect -15241 -66438 -15141 -66404
rect -14983 -66438 -14883 -66404
rect -14725 -66438 -14625 -66404
rect -14467 -66438 -14367 -66404
rect -14209 -66438 -14109 -66404
rect -13951 -66438 -13851 -66404
rect -15241 -66966 -15141 -66932
rect -14983 -66966 -14883 -66932
rect -14725 -66966 -14625 -66932
rect -14467 -66966 -14367 -66932
rect -14209 -66966 -14109 -66932
rect -13951 -66966 -13851 -66932
rect -11241 -65578 -11141 -65544
rect -10983 -65578 -10883 -65544
rect -10725 -65578 -10625 -65544
rect -10467 -65578 -10367 -65544
rect -10209 -65578 -10109 -65544
rect -9951 -65578 -9851 -65544
rect -11241 -66106 -11141 -66072
rect -10983 -66106 -10883 -66072
rect -10725 -66106 -10625 -66072
rect -10467 -66106 -10367 -66072
rect -10209 -66106 -10109 -66072
rect -9951 -66106 -9851 -66072
rect -11241 -66438 -11141 -66404
rect -10983 -66438 -10883 -66404
rect -10725 -66438 -10625 -66404
rect -10467 -66438 -10367 -66404
rect -10209 -66438 -10109 -66404
rect -9951 -66438 -9851 -66404
rect -11241 -66966 -11141 -66932
rect -10983 -66966 -10883 -66932
rect -10725 -66966 -10625 -66932
rect -10467 -66966 -10367 -66932
rect -10209 -66966 -10109 -66932
rect -9951 -66966 -9851 -66932
rect -7241 -65578 -7141 -65544
rect -6983 -65578 -6883 -65544
rect -6725 -65578 -6625 -65544
rect -6467 -65578 -6367 -65544
rect -6209 -65578 -6109 -65544
rect -5951 -65578 -5851 -65544
rect -7241 -66106 -7141 -66072
rect -6983 -66106 -6883 -66072
rect -6725 -66106 -6625 -66072
rect -6467 -66106 -6367 -66072
rect -6209 -66106 -6109 -66072
rect -5951 -66106 -5851 -66072
rect -7241 -66438 -7141 -66404
rect -6983 -66438 -6883 -66404
rect -6725 -66438 -6625 -66404
rect -6467 -66438 -6367 -66404
rect -6209 -66438 -6109 -66404
rect -5951 -66438 -5851 -66404
rect -7241 -66966 -7141 -66932
rect -6983 -66966 -6883 -66932
rect -6725 -66966 -6625 -66932
rect -6467 -66966 -6367 -66932
rect -6209 -66966 -6109 -66932
rect -5951 -66966 -5851 -66932
rect -3241 -65578 -3141 -65544
rect -2983 -65578 -2883 -65544
rect -2725 -65578 -2625 -65544
rect -2467 -65578 -2367 -65544
rect -2209 -65578 -2109 -65544
rect -1951 -65578 -1851 -65544
rect -3241 -66106 -3141 -66072
rect -2983 -66106 -2883 -66072
rect -2725 -66106 -2625 -66072
rect -2467 -66106 -2367 -66072
rect -2209 -66106 -2109 -66072
rect -1951 -66106 -1851 -66072
rect -3241 -66438 -3141 -66404
rect -2983 -66438 -2883 -66404
rect -2725 -66438 -2625 -66404
rect -2467 -66438 -2367 -66404
rect -2209 -66438 -2109 -66404
rect -1951 -66438 -1851 -66404
rect -3241 -66966 -3141 -66932
rect -2983 -66966 -2883 -66932
rect -2725 -66966 -2625 -66932
rect -2467 -66966 -2367 -66932
rect -2209 -66966 -2109 -66932
rect -1951 -66966 -1851 -66932
rect 759 -65578 859 -65544
rect 1017 -65578 1117 -65544
rect 1275 -65578 1375 -65544
rect 1533 -65578 1633 -65544
rect 1791 -65578 1891 -65544
rect 2049 -65578 2149 -65544
rect 759 -66106 859 -66072
rect 1017 -66106 1117 -66072
rect 1275 -66106 1375 -66072
rect 1533 -66106 1633 -66072
rect 1791 -66106 1891 -66072
rect 2049 -66106 2149 -66072
rect 759 -66438 859 -66404
rect 1017 -66438 1117 -66404
rect 1275 -66438 1375 -66404
rect 1533 -66438 1633 -66404
rect 1791 -66438 1891 -66404
rect 2049 -66438 2149 -66404
rect 759 -66966 859 -66932
rect 1017 -66966 1117 -66932
rect 1275 -66966 1375 -66932
rect 1533 -66966 1633 -66932
rect 1791 -66966 1891 -66932
rect 2049 -66966 2149 -66932
rect 4759 -65578 4859 -65544
rect 5017 -65578 5117 -65544
rect 5275 -65578 5375 -65544
rect 5533 -65578 5633 -65544
rect 5791 -65578 5891 -65544
rect 6049 -65578 6149 -65544
rect 4759 -66106 4859 -66072
rect 5017 -66106 5117 -66072
rect 5275 -66106 5375 -66072
rect 5533 -66106 5633 -66072
rect 5791 -66106 5891 -66072
rect 6049 -66106 6149 -66072
rect 4759 -66438 4859 -66404
rect 5017 -66438 5117 -66404
rect 5275 -66438 5375 -66404
rect 5533 -66438 5633 -66404
rect 5791 -66438 5891 -66404
rect 6049 -66438 6149 -66404
rect 4759 -66966 4859 -66932
rect 5017 -66966 5117 -66932
rect 5275 -66966 5375 -66932
rect 5533 -66966 5633 -66932
rect 5791 -66966 5891 -66932
rect 6049 -66966 6149 -66932
rect -27992 -67611 -27958 -67577
rect -23992 -67611 -23958 -67577
rect -19992 -67611 -19958 -67577
rect -15992 -67611 -15958 -67577
rect -11992 -67611 -11958 -67577
rect -7992 -67611 -7958 -67577
rect -3992 -67611 -3958 -67577
rect 8 -67611 42 -67577
rect 4008 -67611 4042 -67577
rect -27246 -68280 -27146 -68246
rect -26988 -68280 -26888 -68246
rect -26730 -68280 -26630 -68246
rect -26472 -68280 -26372 -68246
rect -26214 -68280 -26114 -68246
rect -25956 -68280 -25856 -68246
rect -27246 -68790 -27146 -68756
rect -26988 -68790 -26888 -68756
rect -26730 -68790 -26630 -68756
rect -26472 -68790 -26372 -68756
rect -26214 -68790 -26114 -68756
rect -25956 -68790 -25856 -68756
rect -23246 -68280 -23146 -68246
rect -22988 -68280 -22888 -68246
rect -22730 -68280 -22630 -68246
rect -22472 -68280 -22372 -68246
rect -22214 -68280 -22114 -68246
rect -21956 -68280 -21856 -68246
rect -23246 -68790 -23146 -68756
rect -22988 -68790 -22888 -68756
rect -22730 -68790 -22630 -68756
rect -22472 -68790 -22372 -68756
rect -22214 -68790 -22114 -68756
rect -21956 -68790 -21856 -68756
rect -19246 -68280 -19146 -68246
rect -18988 -68280 -18888 -68246
rect -18730 -68280 -18630 -68246
rect -18472 -68280 -18372 -68246
rect -18214 -68280 -18114 -68246
rect -17956 -68280 -17856 -68246
rect -19246 -68790 -19146 -68756
rect -18988 -68790 -18888 -68756
rect -18730 -68790 -18630 -68756
rect -18472 -68790 -18372 -68756
rect -18214 -68790 -18114 -68756
rect -17956 -68790 -17856 -68756
rect -15246 -68280 -15146 -68246
rect -14988 -68280 -14888 -68246
rect -14730 -68280 -14630 -68246
rect -14472 -68280 -14372 -68246
rect -14214 -68280 -14114 -68246
rect -13956 -68280 -13856 -68246
rect -15246 -68790 -15146 -68756
rect -14988 -68790 -14888 -68756
rect -14730 -68790 -14630 -68756
rect -14472 -68790 -14372 -68756
rect -14214 -68790 -14114 -68756
rect -13956 -68790 -13856 -68756
rect -11246 -68280 -11146 -68246
rect -10988 -68280 -10888 -68246
rect -10730 -68280 -10630 -68246
rect -10472 -68280 -10372 -68246
rect -10214 -68280 -10114 -68246
rect -9956 -68280 -9856 -68246
rect -11246 -68790 -11146 -68756
rect -10988 -68790 -10888 -68756
rect -10730 -68790 -10630 -68756
rect -10472 -68790 -10372 -68756
rect -10214 -68790 -10114 -68756
rect -9956 -68790 -9856 -68756
rect -7246 -68280 -7146 -68246
rect -6988 -68280 -6888 -68246
rect -6730 -68280 -6630 -68246
rect -6472 -68280 -6372 -68246
rect -6214 -68280 -6114 -68246
rect -5956 -68280 -5856 -68246
rect -7246 -68790 -7146 -68756
rect -6988 -68790 -6888 -68756
rect -6730 -68790 -6630 -68756
rect -6472 -68790 -6372 -68756
rect -6214 -68790 -6114 -68756
rect -5956 -68790 -5856 -68756
rect -3246 -68280 -3146 -68246
rect -2988 -68280 -2888 -68246
rect -2730 -68280 -2630 -68246
rect -2472 -68280 -2372 -68246
rect -2214 -68280 -2114 -68246
rect -1956 -68280 -1856 -68246
rect -3246 -68790 -3146 -68756
rect -2988 -68790 -2888 -68756
rect -2730 -68790 -2630 -68756
rect -2472 -68790 -2372 -68756
rect -2214 -68790 -2114 -68756
rect -1956 -68790 -1856 -68756
rect 754 -68280 854 -68246
rect 1012 -68280 1112 -68246
rect 1270 -68280 1370 -68246
rect 1528 -68280 1628 -68246
rect 1786 -68280 1886 -68246
rect 2044 -68280 2144 -68246
rect 754 -68790 854 -68756
rect 1012 -68790 1112 -68756
rect 1270 -68790 1370 -68756
rect 1528 -68790 1628 -68756
rect 1786 -68790 1886 -68756
rect 2044 -68790 2144 -68756
rect 4754 -68280 4854 -68246
rect 5012 -68280 5112 -68246
rect 5270 -68280 5370 -68246
rect 5528 -68280 5628 -68246
rect 5786 -68280 5886 -68246
rect 6044 -68280 6144 -68246
rect 4754 -68790 4854 -68756
rect 5012 -68790 5112 -68756
rect 5270 -68790 5370 -68756
rect 5528 -68790 5628 -68756
rect 5786 -68790 5886 -68756
rect 6044 -68790 6144 -68756
rect -27246 -71440 -27146 -71406
rect -26988 -71440 -26888 -71406
rect -26730 -71440 -26630 -71406
rect -26472 -71440 -26372 -71406
rect -26214 -71440 -26114 -71406
rect -25956 -71440 -25856 -71406
rect -27246 -71950 -27146 -71916
rect -26988 -71950 -26888 -71916
rect -26730 -71950 -26630 -71916
rect -26472 -71950 -26372 -71916
rect -26214 -71950 -26114 -71916
rect -25956 -71950 -25856 -71916
rect -23246 -71440 -23146 -71406
rect -22988 -71440 -22888 -71406
rect -22730 -71440 -22630 -71406
rect -22472 -71440 -22372 -71406
rect -22214 -71440 -22114 -71406
rect -21956 -71440 -21856 -71406
rect -23246 -71950 -23146 -71916
rect -22988 -71950 -22888 -71916
rect -22730 -71950 -22630 -71916
rect -22472 -71950 -22372 -71916
rect -22214 -71950 -22114 -71916
rect -21956 -71950 -21856 -71916
rect -19246 -71440 -19146 -71406
rect -18988 -71440 -18888 -71406
rect -18730 -71440 -18630 -71406
rect -18472 -71440 -18372 -71406
rect -18214 -71440 -18114 -71406
rect -17956 -71440 -17856 -71406
rect -19246 -71950 -19146 -71916
rect -18988 -71950 -18888 -71916
rect -18730 -71950 -18630 -71916
rect -18472 -71950 -18372 -71916
rect -18214 -71950 -18114 -71916
rect -17956 -71950 -17856 -71916
rect -15246 -71440 -15146 -71406
rect -14988 -71440 -14888 -71406
rect -14730 -71440 -14630 -71406
rect -14472 -71440 -14372 -71406
rect -14214 -71440 -14114 -71406
rect -13956 -71440 -13856 -71406
rect -15246 -71950 -15146 -71916
rect -14988 -71950 -14888 -71916
rect -14730 -71950 -14630 -71916
rect -14472 -71950 -14372 -71916
rect -14214 -71950 -14114 -71916
rect -13956 -71950 -13856 -71916
rect -11246 -71440 -11146 -71406
rect -10988 -71440 -10888 -71406
rect -10730 -71440 -10630 -71406
rect -10472 -71440 -10372 -71406
rect -10214 -71440 -10114 -71406
rect -9956 -71440 -9856 -71406
rect -11246 -71950 -11146 -71916
rect -10988 -71950 -10888 -71916
rect -10730 -71950 -10630 -71916
rect -10472 -71950 -10372 -71916
rect -10214 -71950 -10114 -71916
rect -9956 -71950 -9856 -71916
rect -7246 -71440 -7146 -71406
rect -6988 -71440 -6888 -71406
rect -6730 -71440 -6630 -71406
rect -6472 -71440 -6372 -71406
rect -6214 -71440 -6114 -71406
rect -5956 -71440 -5856 -71406
rect -7246 -71950 -7146 -71916
rect -6988 -71950 -6888 -71916
rect -6730 -71950 -6630 -71916
rect -6472 -71950 -6372 -71916
rect -6214 -71950 -6114 -71916
rect -5956 -71950 -5856 -71916
rect -3246 -71440 -3146 -71406
rect -2988 -71440 -2888 -71406
rect -2730 -71440 -2630 -71406
rect -2472 -71440 -2372 -71406
rect -2214 -71440 -2114 -71406
rect -1956 -71440 -1856 -71406
rect -3246 -71950 -3146 -71916
rect -2988 -71950 -2888 -71916
rect -2730 -71950 -2630 -71916
rect -2472 -71950 -2372 -71916
rect -2214 -71950 -2114 -71916
rect -1956 -71950 -1856 -71916
rect 754 -71440 854 -71406
rect 1012 -71440 1112 -71406
rect 1270 -71440 1370 -71406
rect 1528 -71440 1628 -71406
rect 1786 -71440 1886 -71406
rect 2044 -71440 2144 -71406
rect 754 -71950 854 -71916
rect 1012 -71950 1112 -71916
rect 1270 -71950 1370 -71916
rect 1528 -71950 1628 -71916
rect 1786 -71950 1886 -71916
rect 2044 -71950 2144 -71916
rect 4754 -71440 4854 -71406
rect 5012 -71440 5112 -71406
rect 5270 -71440 5370 -71406
rect 5528 -71440 5628 -71406
rect 5786 -71440 5886 -71406
rect 6044 -71440 6144 -71406
rect 4754 -71950 4854 -71916
rect 5012 -71950 5112 -71916
rect 5270 -71950 5370 -71916
rect 5528 -71950 5628 -71916
rect 5786 -71950 5886 -71916
rect 6044 -71950 6144 -71916
rect -27992 -72619 -27958 -72585
rect -23992 -72619 -23958 -72585
rect -19992 -72619 -19958 -72585
rect -15992 -72619 -15958 -72585
rect -11992 -72619 -11958 -72585
rect -7992 -72619 -7958 -72585
rect -3992 -72619 -3958 -72585
rect 8 -72619 42 -72585
rect 4008 -72619 4042 -72585
rect -27241 -73264 -27141 -73230
rect -26983 -73264 -26883 -73230
rect -26725 -73264 -26625 -73230
rect -26467 -73264 -26367 -73230
rect -26209 -73264 -26109 -73230
rect -25951 -73264 -25851 -73230
rect -27241 -73792 -27141 -73758
rect -26983 -73792 -26883 -73758
rect -26725 -73792 -26625 -73758
rect -26467 -73792 -26367 -73758
rect -26209 -73792 -26109 -73758
rect -25951 -73792 -25851 -73758
rect -27241 -74124 -27141 -74090
rect -26983 -74124 -26883 -74090
rect -26725 -74124 -26625 -74090
rect -26467 -74124 -26367 -74090
rect -26209 -74124 -26109 -74090
rect -25951 -74124 -25851 -74090
rect -27241 -74652 -27141 -74618
rect -26983 -74652 -26883 -74618
rect -26725 -74652 -26625 -74618
rect -26467 -74652 -26367 -74618
rect -26209 -74652 -26109 -74618
rect -25951 -74652 -25851 -74618
rect -23241 -73264 -23141 -73230
rect -22983 -73264 -22883 -73230
rect -22725 -73264 -22625 -73230
rect -22467 -73264 -22367 -73230
rect -22209 -73264 -22109 -73230
rect -21951 -73264 -21851 -73230
rect -23241 -73792 -23141 -73758
rect -22983 -73792 -22883 -73758
rect -22725 -73792 -22625 -73758
rect -22467 -73792 -22367 -73758
rect -22209 -73792 -22109 -73758
rect -21951 -73792 -21851 -73758
rect -23241 -74124 -23141 -74090
rect -22983 -74124 -22883 -74090
rect -22725 -74124 -22625 -74090
rect -22467 -74124 -22367 -74090
rect -22209 -74124 -22109 -74090
rect -21951 -74124 -21851 -74090
rect -23241 -74652 -23141 -74618
rect -22983 -74652 -22883 -74618
rect -22725 -74652 -22625 -74618
rect -22467 -74652 -22367 -74618
rect -22209 -74652 -22109 -74618
rect -21951 -74652 -21851 -74618
rect -19241 -73264 -19141 -73230
rect -18983 -73264 -18883 -73230
rect -18725 -73264 -18625 -73230
rect -18467 -73264 -18367 -73230
rect -18209 -73264 -18109 -73230
rect -17951 -73264 -17851 -73230
rect -19241 -73792 -19141 -73758
rect -18983 -73792 -18883 -73758
rect -18725 -73792 -18625 -73758
rect -18467 -73792 -18367 -73758
rect -18209 -73792 -18109 -73758
rect -17951 -73792 -17851 -73758
rect -19241 -74124 -19141 -74090
rect -18983 -74124 -18883 -74090
rect -18725 -74124 -18625 -74090
rect -18467 -74124 -18367 -74090
rect -18209 -74124 -18109 -74090
rect -17951 -74124 -17851 -74090
rect -19241 -74652 -19141 -74618
rect -18983 -74652 -18883 -74618
rect -18725 -74652 -18625 -74618
rect -18467 -74652 -18367 -74618
rect -18209 -74652 -18109 -74618
rect -17951 -74652 -17851 -74618
rect -15241 -73264 -15141 -73230
rect -14983 -73264 -14883 -73230
rect -14725 -73264 -14625 -73230
rect -14467 -73264 -14367 -73230
rect -14209 -73264 -14109 -73230
rect -13951 -73264 -13851 -73230
rect -15241 -73792 -15141 -73758
rect -14983 -73792 -14883 -73758
rect -14725 -73792 -14625 -73758
rect -14467 -73792 -14367 -73758
rect -14209 -73792 -14109 -73758
rect -13951 -73792 -13851 -73758
rect -15241 -74124 -15141 -74090
rect -14983 -74124 -14883 -74090
rect -14725 -74124 -14625 -74090
rect -14467 -74124 -14367 -74090
rect -14209 -74124 -14109 -74090
rect -13951 -74124 -13851 -74090
rect -15241 -74652 -15141 -74618
rect -14983 -74652 -14883 -74618
rect -14725 -74652 -14625 -74618
rect -14467 -74652 -14367 -74618
rect -14209 -74652 -14109 -74618
rect -13951 -74652 -13851 -74618
rect -11241 -73264 -11141 -73230
rect -10983 -73264 -10883 -73230
rect -10725 -73264 -10625 -73230
rect -10467 -73264 -10367 -73230
rect -10209 -73264 -10109 -73230
rect -9951 -73264 -9851 -73230
rect -11241 -73792 -11141 -73758
rect -10983 -73792 -10883 -73758
rect -10725 -73792 -10625 -73758
rect -10467 -73792 -10367 -73758
rect -10209 -73792 -10109 -73758
rect -9951 -73792 -9851 -73758
rect -11241 -74124 -11141 -74090
rect -10983 -74124 -10883 -74090
rect -10725 -74124 -10625 -74090
rect -10467 -74124 -10367 -74090
rect -10209 -74124 -10109 -74090
rect -9951 -74124 -9851 -74090
rect -11241 -74652 -11141 -74618
rect -10983 -74652 -10883 -74618
rect -10725 -74652 -10625 -74618
rect -10467 -74652 -10367 -74618
rect -10209 -74652 -10109 -74618
rect -9951 -74652 -9851 -74618
rect -7241 -73264 -7141 -73230
rect -6983 -73264 -6883 -73230
rect -6725 -73264 -6625 -73230
rect -6467 -73264 -6367 -73230
rect -6209 -73264 -6109 -73230
rect -5951 -73264 -5851 -73230
rect -7241 -73792 -7141 -73758
rect -6983 -73792 -6883 -73758
rect -6725 -73792 -6625 -73758
rect -6467 -73792 -6367 -73758
rect -6209 -73792 -6109 -73758
rect -5951 -73792 -5851 -73758
rect -7241 -74124 -7141 -74090
rect -6983 -74124 -6883 -74090
rect -6725 -74124 -6625 -74090
rect -6467 -74124 -6367 -74090
rect -6209 -74124 -6109 -74090
rect -5951 -74124 -5851 -74090
rect -7241 -74652 -7141 -74618
rect -6983 -74652 -6883 -74618
rect -6725 -74652 -6625 -74618
rect -6467 -74652 -6367 -74618
rect -6209 -74652 -6109 -74618
rect -5951 -74652 -5851 -74618
rect -3241 -73264 -3141 -73230
rect -2983 -73264 -2883 -73230
rect -2725 -73264 -2625 -73230
rect -2467 -73264 -2367 -73230
rect -2209 -73264 -2109 -73230
rect -1951 -73264 -1851 -73230
rect -3241 -73792 -3141 -73758
rect -2983 -73792 -2883 -73758
rect -2725 -73792 -2625 -73758
rect -2467 -73792 -2367 -73758
rect -2209 -73792 -2109 -73758
rect -1951 -73792 -1851 -73758
rect -3241 -74124 -3141 -74090
rect -2983 -74124 -2883 -74090
rect -2725 -74124 -2625 -74090
rect -2467 -74124 -2367 -74090
rect -2209 -74124 -2109 -74090
rect -1951 -74124 -1851 -74090
rect -3241 -74652 -3141 -74618
rect -2983 -74652 -2883 -74618
rect -2725 -74652 -2625 -74618
rect -2467 -74652 -2367 -74618
rect -2209 -74652 -2109 -74618
rect -1951 -74652 -1851 -74618
rect 759 -73264 859 -73230
rect 1017 -73264 1117 -73230
rect 1275 -73264 1375 -73230
rect 1533 -73264 1633 -73230
rect 1791 -73264 1891 -73230
rect 2049 -73264 2149 -73230
rect 759 -73792 859 -73758
rect 1017 -73792 1117 -73758
rect 1275 -73792 1375 -73758
rect 1533 -73792 1633 -73758
rect 1791 -73792 1891 -73758
rect 2049 -73792 2149 -73758
rect 759 -74124 859 -74090
rect 1017 -74124 1117 -74090
rect 1275 -74124 1375 -74090
rect 1533 -74124 1633 -74090
rect 1791 -74124 1891 -74090
rect 2049 -74124 2149 -74090
rect 759 -74652 859 -74618
rect 1017 -74652 1117 -74618
rect 1275 -74652 1375 -74618
rect 1533 -74652 1633 -74618
rect 1791 -74652 1891 -74618
rect 2049 -74652 2149 -74618
rect 4759 -73264 4859 -73230
rect 5017 -73264 5117 -73230
rect 5275 -73264 5375 -73230
rect 5533 -73264 5633 -73230
rect 5791 -73264 5891 -73230
rect 6049 -73264 6149 -73230
rect 4759 -73792 4859 -73758
rect 5017 -73792 5117 -73758
rect 5275 -73792 5375 -73758
rect 5533 -73792 5633 -73758
rect 5791 -73792 5891 -73758
rect 6049 -73792 6149 -73758
rect 4759 -74124 4859 -74090
rect 5017 -74124 5117 -74090
rect 5275 -74124 5375 -74090
rect 5533 -74124 5633 -74090
rect 5791 -74124 5891 -74090
rect 6049 -74124 6149 -74090
rect 4759 -74652 4859 -74618
rect 5017 -74652 5117 -74618
rect 5275 -74652 5375 -74618
rect 5533 -74652 5633 -74618
rect 5791 -74652 5891 -74618
rect 6049 -74652 6149 -74618
<< locali >>
rect 25822 -27818 25922 -27656
rect 50166 -27818 50266 -27656
rect 32412 -30200 32502 -30170
rect 32412 -30234 32440 -30200
rect 32474 -30234 32502 -30200
rect 32412 -30262 32502 -30234
rect 33430 -30200 33520 -30170
rect 33430 -30234 33458 -30200
rect 33492 -30234 33520 -30200
rect 33430 -30262 33520 -30234
rect 34448 -30200 34538 -30170
rect 34448 -30234 34476 -30200
rect 34510 -30234 34538 -30200
rect 34448 -30262 34538 -30234
rect 35466 -30200 35556 -30170
rect 35466 -30234 35494 -30200
rect 35528 -30234 35556 -30200
rect 35466 -30262 35556 -30234
rect 36484 -30200 36574 -30170
rect 36484 -30234 36512 -30200
rect 36546 -30234 36574 -30200
rect 36484 -30262 36574 -30234
rect 37502 -30200 37592 -30170
rect 37502 -30234 37530 -30200
rect 37564 -30234 37592 -30200
rect 37502 -30262 37592 -30234
rect 38520 -30200 38610 -30170
rect 38520 -30234 38548 -30200
rect 38582 -30234 38610 -30200
rect 38520 -30262 38610 -30234
rect 39538 -30200 39628 -30170
rect 39538 -30234 39566 -30200
rect 39600 -30234 39628 -30200
rect 39538 -30262 39628 -30234
rect 40556 -30200 40646 -30170
rect 40556 -30234 40584 -30200
rect 40618 -30234 40646 -30200
rect 40556 -30262 40646 -30234
rect 41574 -30200 41664 -30170
rect 41574 -30234 41602 -30200
rect 41636 -30234 41664 -30200
rect 41574 -30262 41664 -30234
rect 42592 -30200 42682 -30170
rect 42592 -30234 42620 -30200
rect 42654 -30234 42682 -30200
rect 42592 -30262 42682 -30234
rect 43610 -30200 43700 -30170
rect 43610 -30234 43638 -30200
rect 43672 -30234 43700 -30200
rect 43610 -30262 43700 -30234
rect 44628 -30200 44718 -30170
rect 44628 -30234 44656 -30200
rect 44690 -30234 44718 -30200
rect 44628 -30262 44718 -30234
rect 45646 -30200 45736 -30170
rect 45646 -30234 45674 -30200
rect 45708 -30234 45736 -30200
rect 45646 -30262 45736 -30234
rect 46664 -30200 46754 -30170
rect 46664 -30234 46692 -30200
rect 46726 -30234 46754 -30200
rect 46664 -30262 46754 -30234
rect 47682 -30200 47772 -30170
rect 47682 -30234 47710 -30200
rect 47744 -30234 47772 -30200
rect 47682 -30262 47772 -30234
rect 32164 -30457 32180 -30423
rect 32736 -30457 32752 -30423
rect 33182 -30457 33198 -30423
rect 33754 -30457 33770 -30423
rect 34200 -30457 34216 -30423
rect 34772 -30457 34788 -30423
rect 35218 -30457 35234 -30423
rect 35790 -30457 35806 -30423
rect 36236 -30457 36252 -30423
rect 36808 -30457 36824 -30423
rect 37254 -30457 37270 -30423
rect 37826 -30457 37842 -30423
rect 38272 -30457 38288 -30423
rect 38844 -30457 38860 -30423
rect 39290 -30457 39306 -30423
rect 39862 -30457 39878 -30423
rect 40308 -30457 40324 -30423
rect 40880 -30457 40896 -30423
rect 41326 -30457 41342 -30423
rect 41898 -30457 41914 -30423
rect 42344 -30457 42360 -30423
rect 42916 -30457 42932 -30423
rect 43362 -30457 43378 -30423
rect 43934 -30457 43950 -30423
rect 44380 -30457 44396 -30423
rect 44952 -30457 44968 -30423
rect 45398 -30457 45414 -30423
rect 45970 -30457 45986 -30423
rect 46416 -30457 46432 -30423
rect 46988 -30457 47004 -30423
rect 47434 -30457 47450 -30423
rect 48006 -30457 48022 -30423
rect 31932 -30516 31966 -30500
rect 31932 -31108 31966 -31092
rect 32950 -30516 32984 -30500
rect 32950 -31108 32984 -31092
rect 33968 -30516 34002 -30500
rect 33968 -31108 34002 -31092
rect 34986 -30516 35020 -30500
rect 34986 -31108 35020 -31092
rect 36004 -30516 36038 -30500
rect 36004 -31108 36038 -31092
rect 37022 -30516 37056 -30500
rect 37022 -31108 37056 -31092
rect 38040 -30516 38074 -30500
rect 38040 -31108 38074 -31092
rect 39058 -30516 39092 -30500
rect 39058 -31108 39092 -31092
rect 40076 -30516 40110 -30500
rect 40076 -31108 40110 -31092
rect 41094 -30516 41128 -30500
rect 41094 -31108 41128 -31092
rect 42112 -30516 42146 -30500
rect 42112 -31108 42146 -31092
rect 43130 -30516 43164 -30500
rect 43130 -31108 43164 -31092
rect 44148 -30516 44182 -30500
rect 44148 -31108 44182 -31092
rect 45166 -30516 45200 -30500
rect 45166 -31108 45200 -31092
rect 46184 -30516 46218 -30500
rect 46184 -31108 46218 -31092
rect 47202 -30516 47236 -30500
rect 47202 -31108 47236 -31092
rect 48220 -30516 48254 -30500
rect 48220 -31108 48254 -31092
rect 32164 -31185 32180 -31151
rect 32736 -31185 32752 -31151
rect 33182 -31185 33198 -31151
rect 33754 -31185 33770 -31151
rect 34200 -31185 34216 -31151
rect 34772 -31185 34788 -31151
rect 35218 -31185 35234 -31151
rect 35790 -31185 35806 -31151
rect 36236 -31185 36252 -31151
rect 36808 -31185 36824 -31151
rect 37254 -31185 37270 -31151
rect 37826 -31185 37842 -31151
rect 38272 -31185 38288 -31151
rect 38844 -31185 38860 -31151
rect 39290 -31185 39306 -31151
rect 39862 -31185 39878 -31151
rect 40308 -31185 40324 -31151
rect 40880 -31185 40896 -31151
rect 41326 -31185 41342 -31151
rect 41898 -31185 41914 -31151
rect 42344 -31185 42360 -31151
rect 42916 -31185 42932 -31151
rect 43362 -31185 43378 -31151
rect 43934 -31185 43950 -31151
rect 44380 -31185 44396 -31151
rect 44952 -31185 44968 -31151
rect 45398 -31185 45414 -31151
rect 45970 -31185 45986 -31151
rect 46416 -31185 46432 -31151
rect 46988 -31185 47004 -31151
rect 47434 -31185 47450 -31151
rect 48006 -31185 48022 -31151
rect 32434 -31354 32524 -31324
rect 32434 -31388 32462 -31354
rect 32496 -31388 32524 -31354
rect 32434 -31416 32524 -31388
rect 33452 -31354 33542 -31324
rect 33452 -31388 33480 -31354
rect 33514 -31388 33542 -31354
rect 33452 -31416 33542 -31388
rect 34470 -31354 34560 -31324
rect 34470 -31388 34498 -31354
rect 34532 -31388 34560 -31354
rect 34470 -31416 34560 -31388
rect 35488 -31354 35578 -31324
rect 35488 -31388 35516 -31354
rect 35550 -31388 35578 -31354
rect 35488 -31416 35578 -31388
rect 36506 -31354 36596 -31324
rect 36506 -31388 36534 -31354
rect 36568 -31388 36596 -31354
rect 36506 -31416 36596 -31388
rect 37524 -31354 37614 -31324
rect 37524 -31388 37552 -31354
rect 37586 -31388 37614 -31354
rect 37524 -31416 37614 -31388
rect 38542 -31354 38632 -31324
rect 38542 -31388 38570 -31354
rect 38604 -31388 38632 -31354
rect 38542 -31416 38632 -31388
rect 39560 -31354 39650 -31324
rect 39560 -31388 39588 -31354
rect 39622 -31388 39650 -31354
rect 39560 -31416 39650 -31388
rect 40578 -31354 40668 -31324
rect 40578 -31388 40606 -31354
rect 40640 -31388 40668 -31354
rect 40578 -31416 40668 -31388
rect 41596 -31354 41686 -31324
rect 41596 -31388 41624 -31354
rect 41658 -31388 41686 -31354
rect 41596 -31416 41686 -31388
rect 42614 -31354 42704 -31324
rect 42614 -31388 42642 -31354
rect 42676 -31388 42704 -31354
rect 42614 -31416 42704 -31388
rect 43632 -31354 43722 -31324
rect 43632 -31388 43660 -31354
rect 43694 -31388 43722 -31354
rect 43632 -31416 43722 -31388
rect 44650 -31354 44740 -31324
rect 44650 -31388 44678 -31354
rect 44712 -31388 44740 -31354
rect 44650 -31416 44740 -31388
rect 45668 -31354 45758 -31324
rect 45668 -31388 45696 -31354
rect 45730 -31388 45758 -31354
rect 45668 -31416 45758 -31388
rect 46686 -31354 46776 -31324
rect 46686 -31388 46714 -31354
rect 46748 -31388 46776 -31354
rect 46686 -31416 46776 -31388
rect 47704 -31354 47794 -31324
rect 47704 -31388 47732 -31354
rect 47766 -31388 47794 -31354
rect 47704 -31416 47794 -31388
rect 32164 -31593 32180 -31559
rect 32736 -31593 32752 -31559
rect 33182 -31593 33198 -31559
rect 33754 -31593 33770 -31559
rect 34200 -31593 34216 -31559
rect 34772 -31593 34788 -31559
rect 35218 -31593 35234 -31559
rect 35790 -31593 35806 -31559
rect 36236 -31593 36252 -31559
rect 36808 -31593 36824 -31559
rect 37254 -31593 37270 -31559
rect 37826 -31593 37842 -31559
rect 38272 -31593 38288 -31559
rect 38844 -31593 38860 -31559
rect 39290 -31593 39306 -31559
rect 39862 -31593 39878 -31559
rect 40308 -31593 40324 -31559
rect 40880 -31593 40896 -31559
rect 41326 -31593 41342 -31559
rect 41898 -31593 41914 -31559
rect 42344 -31593 42360 -31559
rect 42916 -31593 42932 -31559
rect 43362 -31593 43378 -31559
rect 43934 -31593 43950 -31559
rect 44380 -31593 44396 -31559
rect 44952 -31593 44968 -31559
rect 45398 -31593 45414 -31559
rect 45970 -31593 45986 -31559
rect 46416 -31593 46432 -31559
rect 46988 -31593 47004 -31559
rect 47434 -31593 47450 -31559
rect 48006 -31593 48022 -31559
rect 31932 -31652 31966 -31636
rect 31932 -32244 31966 -32228
rect 32950 -31652 32984 -31636
rect 32950 -32244 32984 -32228
rect 33968 -31652 34002 -31636
rect 33968 -32244 34002 -32228
rect 34986 -31652 35020 -31636
rect 34986 -32244 35020 -32228
rect 36004 -31652 36038 -31636
rect 36004 -32244 36038 -32228
rect 37022 -31652 37056 -31636
rect 37022 -32244 37056 -32228
rect 38040 -31652 38074 -31636
rect 38040 -32244 38074 -32228
rect 39058 -31652 39092 -31636
rect 39058 -32244 39092 -32228
rect 40076 -31652 40110 -31636
rect 40076 -32244 40110 -32228
rect 41094 -31652 41128 -31636
rect 41094 -32244 41128 -32228
rect 42112 -31652 42146 -31636
rect 42112 -32244 42146 -32228
rect 43130 -31652 43164 -31636
rect 43130 -32244 43164 -32228
rect 44148 -31652 44182 -31636
rect 44148 -32244 44182 -32228
rect 45166 -31652 45200 -31636
rect 45166 -32244 45200 -32228
rect 46184 -31652 46218 -31636
rect 46184 -32244 46218 -32228
rect 47202 -31652 47236 -31636
rect 47202 -32244 47236 -32228
rect 48220 -31652 48254 -31636
rect 48220 -32244 48254 -32228
rect 32164 -32321 32180 -32287
rect 32736 -32321 32752 -32287
rect 33182 -32321 33198 -32287
rect 33754 -32321 33770 -32287
rect 34200 -32321 34216 -32287
rect 34772 -32321 34788 -32287
rect 35218 -32321 35234 -32287
rect 35790 -32321 35806 -32287
rect 36236 -32321 36252 -32287
rect 36808 -32321 36824 -32287
rect 37254 -32321 37270 -32287
rect 37826 -32321 37842 -32287
rect 38272 -32321 38288 -32287
rect 38844 -32321 38860 -32287
rect 39290 -32321 39306 -32287
rect 39862 -32321 39878 -32287
rect 40308 -32321 40324 -32287
rect 40880 -32321 40896 -32287
rect 41326 -32321 41342 -32287
rect 41898 -32321 41914 -32287
rect 42344 -32321 42360 -32287
rect 42916 -32321 42932 -32287
rect 43362 -32321 43378 -32287
rect 43934 -32321 43950 -32287
rect 44380 -32321 44396 -32287
rect 44952 -32321 44968 -32287
rect 45398 -32321 45414 -32287
rect 45970 -32321 45986 -32287
rect 46416 -32321 46432 -32287
rect 46988 -32321 47004 -32287
rect 47434 -32321 47450 -32287
rect 48006 -32321 48022 -32287
rect 32412 -32486 32502 -32456
rect 32412 -32520 32440 -32486
rect 32474 -32520 32502 -32486
rect 32412 -32548 32502 -32520
rect 33430 -32486 33520 -32456
rect 33430 -32520 33458 -32486
rect 33492 -32520 33520 -32486
rect 33430 -32548 33520 -32520
rect 34448 -32486 34538 -32456
rect 34448 -32520 34476 -32486
rect 34510 -32520 34538 -32486
rect 34448 -32548 34538 -32520
rect 35466 -32486 35556 -32456
rect 35466 -32520 35494 -32486
rect 35528 -32520 35556 -32486
rect 35466 -32548 35556 -32520
rect 36484 -32486 36574 -32456
rect 36484 -32520 36512 -32486
rect 36546 -32520 36574 -32486
rect 36484 -32548 36574 -32520
rect 37502 -32486 37592 -32456
rect 37502 -32520 37530 -32486
rect 37564 -32520 37592 -32486
rect 37502 -32548 37592 -32520
rect 38520 -32486 38610 -32456
rect 38520 -32520 38548 -32486
rect 38582 -32520 38610 -32486
rect 38520 -32548 38610 -32520
rect 39538 -32486 39628 -32456
rect 39538 -32520 39566 -32486
rect 39600 -32520 39628 -32486
rect 39538 -32548 39628 -32520
rect 40556 -32486 40646 -32456
rect 40556 -32520 40584 -32486
rect 40618 -32520 40646 -32486
rect 40556 -32548 40646 -32520
rect 41574 -32486 41664 -32456
rect 41574 -32520 41602 -32486
rect 41636 -32520 41664 -32486
rect 41574 -32548 41664 -32520
rect 42592 -32486 42682 -32456
rect 42592 -32520 42620 -32486
rect 42654 -32520 42682 -32486
rect 42592 -32548 42682 -32520
rect 43610 -32486 43700 -32456
rect 43610 -32520 43638 -32486
rect 43672 -32520 43700 -32486
rect 43610 -32548 43700 -32520
rect 44628 -32486 44718 -32456
rect 44628 -32520 44656 -32486
rect 44690 -32520 44718 -32486
rect 44628 -32548 44718 -32520
rect 45646 -32486 45736 -32456
rect 45646 -32520 45674 -32486
rect 45708 -32520 45736 -32486
rect 45646 -32548 45736 -32520
rect 46664 -32486 46754 -32456
rect 46664 -32520 46692 -32486
rect 46726 -32520 46754 -32486
rect 46664 -32548 46754 -32520
rect 47682 -32486 47772 -32456
rect 47682 -32520 47710 -32486
rect 47744 -32520 47772 -32486
rect 47682 -32548 47772 -32520
rect 32164 -32729 32180 -32695
rect 32736 -32729 32752 -32695
rect 33182 -32729 33198 -32695
rect 33754 -32729 33770 -32695
rect 34200 -32729 34216 -32695
rect 34772 -32729 34788 -32695
rect 35218 -32729 35234 -32695
rect 35790 -32729 35806 -32695
rect 36236 -32729 36252 -32695
rect 36808 -32729 36824 -32695
rect 37254 -32729 37270 -32695
rect 37826 -32729 37842 -32695
rect 38272 -32729 38288 -32695
rect 38844 -32729 38860 -32695
rect 39290 -32729 39306 -32695
rect 39862 -32729 39878 -32695
rect 40308 -32729 40324 -32695
rect 40880 -32729 40896 -32695
rect 41326 -32729 41342 -32695
rect 41898 -32729 41914 -32695
rect 42344 -32729 42360 -32695
rect 42916 -32729 42932 -32695
rect 43362 -32729 43378 -32695
rect 43934 -32729 43950 -32695
rect 44380 -32729 44396 -32695
rect 44952 -32729 44968 -32695
rect 45398 -32729 45414 -32695
rect 45970 -32729 45986 -32695
rect 46416 -32729 46432 -32695
rect 46988 -32729 47004 -32695
rect 47434 -32729 47450 -32695
rect 48006 -32729 48022 -32695
rect 31932 -32788 31966 -32772
rect 31932 -33380 31966 -33364
rect 32950 -32788 32984 -32772
rect 32950 -33380 32984 -33364
rect 33968 -32788 34002 -32772
rect 33968 -33380 34002 -33364
rect 34986 -32788 35020 -32772
rect 34986 -33380 35020 -33364
rect 36004 -32788 36038 -32772
rect 36004 -33380 36038 -33364
rect 37022 -32788 37056 -32772
rect 37022 -33380 37056 -33364
rect 38040 -32788 38074 -32772
rect 38040 -33380 38074 -33364
rect 39058 -32788 39092 -32772
rect 39058 -33380 39092 -33364
rect 40076 -32788 40110 -32772
rect 40076 -33380 40110 -33364
rect 41094 -32788 41128 -32772
rect 41094 -33380 41128 -33364
rect 42112 -32788 42146 -32772
rect 42112 -33380 42146 -33364
rect 43130 -32788 43164 -32772
rect 43130 -33380 43164 -33364
rect 44148 -32788 44182 -32772
rect 44148 -33380 44182 -33364
rect 45166 -32788 45200 -32772
rect 45166 -33380 45200 -33364
rect 46184 -32788 46218 -32772
rect 46184 -33380 46218 -33364
rect 47202 -32788 47236 -32772
rect 47202 -33380 47236 -33364
rect 48220 -32788 48254 -32772
rect 48220 -33380 48254 -33364
rect 32164 -33457 32180 -33423
rect 32736 -33457 32752 -33423
rect 33182 -33457 33198 -33423
rect 33754 -33457 33770 -33423
rect 34200 -33457 34216 -33423
rect 34772 -33457 34788 -33423
rect 35218 -33457 35234 -33423
rect 35790 -33457 35806 -33423
rect 36236 -33457 36252 -33423
rect 36808 -33457 36824 -33423
rect 37254 -33457 37270 -33423
rect 37826 -33457 37842 -33423
rect 38272 -33457 38288 -33423
rect 38844 -33457 38860 -33423
rect 39290 -33457 39306 -33423
rect 39862 -33457 39878 -33423
rect 40308 -33457 40324 -33423
rect 40880 -33457 40896 -33423
rect 41326 -33457 41342 -33423
rect 41898 -33457 41914 -33423
rect 42344 -33457 42360 -33423
rect 42916 -33457 42932 -33423
rect 43362 -33457 43378 -33423
rect 43934 -33457 43950 -33423
rect 44380 -33457 44396 -33423
rect 44952 -33457 44968 -33423
rect 45398 -33457 45414 -33423
rect 45970 -33457 45986 -33423
rect 46416 -33457 46432 -33423
rect 46988 -33457 47004 -33423
rect 47434 -33457 47450 -33423
rect 48006 -33457 48022 -33423
rect 32412 -33868 32502 -33838
rect 32412 -33902 32440 -33868
rect 32474 -33902 32502 -33868
rect 32412 -33930 32502 -33902
rect 33430 -33868 33520 -33838
rect 33430 -33902 33458 -33868
rect 33492 -33902 33520 -33868
rect 33430 -33930 33520 -33902
rect 34448 -33868 34538 -33838
rect 34448 -33902 34476 -33868
rect 34510 -33902 34538 -33868
rect 34448 -33930 34538 -33902
rect 35466 -33868 35556 -33838
rect 35466 -33902 35494 -33868
rect 35528 -33902 35556 -33868
rect 35466 -33930 35556 -33902
rect 36484 -33868 36574 -33838
rect 36484 -33902 36512 -33868
rect 36546 -33902 36574 -33868
rect 36484 -33930 36574 -33902
rect 37502 -33868 37592 -33838
rect 37502 -33902 37530 -33868
rect 37564 -33902 37592 -33868
rect 37502 -33930 37592 -33902
rect 38520 -33868 38610 -33838
rect 38520 -33902 38548 -33868
rect 38582 -33902 38610 -33868
rect 38520 -33930 38610 -33902
rect 39538 -33868 39628 -33838
rect 39538 -33902 39566 -33868
rect 39600 -33902 39628 -33868
rect 39538 -33930 39628 -33902
rect 40556 -33868 40646 -33838
rect 40556 -33902 40584 -33868
rect 40618 -33902 40646 -33868
rect 40556 -33930 40646 -33902
rect 41574 -33868 41664 -33838
rect 41574 -33902 41602 -33868
rect 41636 -33902 41664 -33868
rect 41574 -33930 41664 -33902
rect 42592 -33868 42682 -33838
rect 42592 -33902 42620 -33868
rect 42654 -33902 42682 -33868
rect 42592 -33930 42682 -33902
rect 43610 -33868 43700 -33838
rect 43610 -33902 43638 -33868
rect 43672 -33902 43700 -33868
rect 43610 -33930 43700 -33902
rect 44628 -33868 44718 -33838
rect 44628 -33902 44656 -33868
rect 44690 -33902 44718 -33868
rect 44628 -33930 44718 -33902
rect 45646 -33868 45736 -33838
rect 45646 -33902 45674 -33868
rect 45708 -33902 45736 -33868
rect 45646 -33930 45736 -33902
rect 46664 -33868 46754 -33838
rect 46664 -33902 46692 -33868
rect 46726 -33902 46754 -33868
rect 46664 -33930 46754 -33902
rect 47682 -33868 47772 -33838
rect 47682 -33902 47710 -33868
rect 47744 -33902 47772 -33868
rect 47682 -33930 47772 -33902
rect 33358 -34367 33374 -34333
rect 33930 -34367 33946 -34333
rect 34376 -34367 34392 -34333
rect 34948 -34367 34964 -34333
rect 35394 -34367 35410 -34333
rect 35966 -34367 35982 -34333
rect 36412 -34367 36428 -34333
rect 36984 -34367 37000 -34333
rect 37430 -34367 37446 -34333
rect 38002 -34367 38018 -34333
rect 38448 -34367 38464 -34333
rect 39020 -34367 39036 -34333
rect 39466 -34367 39482 -34333
rect 40038 -34367 40054 -34333
rect 40484 -34367 40500 -34333
rect 41056 -34367 41072 -34333
rect 41502 -34367 41518 -34333
rect 42074 -34367 42090 -34333
rect 42520 -34367 42536 -34333
rect 43092 -34367 43108 -34333
rect 43538 -34367 43554 -34333
rect 44110 -34367 44126 -34333
rect 44556 -34367 44572 -34333
rect 45128 -34367 45144 -34333
rect 45574 -34367 45590 -34333
rect 46146 -34367 46162 -34333
rect 46592 -34367 46608 -34333
rect 47164 -34367 47180 -34333
rect 33126 -34426 33160 -34410
rect 33126 -35018 33160 -35002
rect 34144 -34426 34178 -34410
rect 34144 -35018 34178 -35002
rect 35162 -34426 35196 -34410
rect 35162 -35018 35196 -35002
rect 36180 -34426 36214 -34410
rect 36180 -35018 36214 -35002
rect 37198 -34426 37232 -34410
rect 37198 -35018 37232 -35002
rect 38216 -34426 38250 -34410
rect 38216 -35018 38250 -35002
rect 39234 -34426 39268 -34410
rect 39234 -35018 39268 -35002
rect 40252 -34426 40286 -34410
rect 40252 -35018 40286 -35002
rect 41270 -34426 41304 -34410
rect 41270 -35018 41304 -35002
rect 42288 -34426 42322 -34410
rect 42288 -35018 42322 -35002
rect 43306 -34426 43340 -34410
rect 43306 -35018 43340 -35002
rect 44324 -34426 44358 -34410
rect 44324 -35018 44358 -35002
rect 45342 -34426 45376 -34410
rect 45342 -35018 45376 -35002
rect 46360 -34426 46394 -34410
rect 46360 -35018 46394 -35002
rect 47378 -34426 47412 -34410
rect 47378 -35018 47412 -35002
rect 33358 -35095 33374 -35061
rect 33930 -35095 33946 -35061
rect 34376 -35095 34392 -35061
rect 34948 -35095 34964 -35061
rect 35394 -35095 35410 -35061
rect 35966 -35095 35982 -35061
rect 36412 -35095 36428 -35061
rect 36984 -35095 37000 -35061
rect 37430 -35095 37446 -35061
rect 38002 -35095 38018 -35061
rect 38448 -35095 38464 -35061
rect 39020 -35095 39036 -35061
rect 39466 -35095 39482 -35061
rect 40038 -35095 40054 -35061
rect 40484 -35095 40500 -35061
rect 41056 -35095 41072 -35061
rect 41502 -35095 41518 -35061
rect 42074 -35095 42090 -35061
rect 42520 -35095 42536 -35061
rect 43092 -35095 43108 -35061
rect 43538 -35095 43554 -35061
rect 44110 -35095 44126 -35061
rect 44556 -35095 44572 -35061
rect 45128 -35095 45144 -35061
rect 45574 -35095 45590 -35061
rect 46146 -35095 46162 -35061
rect 46592 -35095 46608 -35061
rect 47164 -35095 47180 -35061
rect 33100 -35216 33190 -35186
rect 33100 -35250 33128 -35216
rect 33162 -35250 33190 -35216
rect 33100 -35278 33190 -35250
rect 34118 -35216 34208 -35186
rect 34118 -35250 34146 -35216
rect 34180 -35250 34208 -35216
rect 34118 -35278 34208 -35250
rect 35136 -35216 35226 -35186
rect 35136 -35250 35164 -35216
rect 35198 -35250 35226 -35216
rect 35136 -35278 35226 -35250
rect 36154 -35216 36244 -35186
rect 36154 -35250 36182 -35216
rect 36216 -35250 36244 -35216
rect 36154 -35278 36244 -35250
rect 37172 -35216 37262 -35186
rect 37172 -35250 37200 -35216
rect 37234 -35250 37262 -35216
rect 37172 -35278 37262 -35250
rect 38190 -35216 38280 -35186
rect 38190 -35250 38218 -35216
rect 38252 -35250 38280 -35216
rect 38190 -35278 38280 -35250
rect 39208 -35216 39298 -35186
rect 39208 -35250 39236 -35216
rect 39270 -35250 39298 -35216
rect 39208 -35278 39298 -35250
rect 40226 -35216 40316 -35186
rect 40226 -35250 40254 -35216
rect 40288 -35250 40316 -35216
rect 40226 -35278 40316 -35250
rect 41244 -35216 41334 -35186
rect 41244 -35250 41272 -35216
rect 41306 -35250 41334 -35216
rect 41244 -35278 41334 -35250
rect 42262 -35216 42352 -35186
rect 42262 -35250 42290 -35216
rect 42324 -35250 42352 -35216
rect 42262 -35278 42352 -35250
rect 43280 -35216 43370 -35186
rect 43280 -35250 43308 -35216
rect 43342 -35250 43370 -35216
rect 43280 -35278 43370 -35250
rect 44298 -35216 44388 -35186
rect 44298 -35250 44326 -35216
rect 44360 -35250 44388 -35216
rect 44298 -35278 44388 -35250
rect 45316 -35216 45406 -35186
rect 45316 -35250 45344 -35216
rect 45378 -35250 45406 -35216
rect 45316 -35278 45406 -35250
rect 46334 -35216 46424 -35186
rect 46334 -35250 46362 -35216
rect 46396 -35250 46424 -35216
rect 46334 -35278 46424 -35250
rect 47352 -35216 47442 -35186
rect 47352 -35250 47380 -35216
rect 47414 -35250 47442 -35216
rect 47352 -35278 47442 -35250
rect 33358 -35399 33374 -35365
rect 33930 -35399 33946 -35365
rect 34376 -35399 34392 -35365
rect 34948 -35399 34964 -35365
rect 35394 -35399 35410 -35365
rect 35966 -35399 35982 -35365
rect 36412 -35399 36428 -35365
rect 36984 -35399 37000 -35365
rect 37430 -35399 37446 -35365
rect 38002 -35399 38018 -35365
rect 38448 -35399 38464 -35365
rect 39020 -35399 39036 -35365
rect 39466 -35399 39482 -35365
rect 40038 -35399 40054 -35365
rect 40484 -35399 40500 -35365
rect 41056 -35399 41072 -35365
rect 41502 -35399 41518 -35365
rect 42074 -35399 42090 -35365
rect 42520 -35399 42536 -35365
rect 43092 -35399 43108 -35365
rect 43538 -35399 43554 -35365
rect 44110 -35399 44126 -35365
rect 44556 -35399 44572 -35365
rect 45128 -35399 45144 -35365
rect 45574 -35399 45590 -35365
rect 46146 -35399 46162 -35365
rect 46592 -35399 46608 -35365
rect 47164 -35399 47180 -35365
rect 33126 -35458 33160 -35442
rect 33126 -36050 33160 -36034
rect 34144 -35458 34178 -35442
rect 34144 -36050 34178 -36034
rect 35162 -35458 35196 -35442
rect 35162 -36050 35196 -36034
rect 36180 -35458 36214 -35442
rect 36180 -36050 36214 -36034
rect 37198 -35458 37232 -35442
rect 37198 -36050 37232 -36034
rect 38216 -35458 38250 -35442
rect 38216 -36050 38250 -36034
rect 39234 -35458 39268 -35442
rect 39234 -36050 39268 -36034
rect 40252 -35458 40286 -35442
rect 40252 -36050 40286 -36034
rect 41270 -35458 41304 -35442
rect 41270 -36050 41304 -36034
rect 42288 -35458 42322 -35442
rect 42288 -36050 42322 -36034
rect 43306 -35458 43340 -35442
rect 43306 -36050 43340 -36034
rect 44324 -35458 44358 -35442
rect 44324 -36050 44358 -36034
rect 45342 -35458 45376 -35442
rect 45342 -36050 45376 -36034
rect 46360 -35458 46394 -35442
rect 46360 -36050 46394 -36034
rect 47378 -35458 47412 -35442
rect 47378 -36050 47412 -36034
rect 33358 -36127 33374 -36093
rect 33930 -36127 33946 -36093
rect 34376 -36127 34392 -36093
rect 34948 -36127 34964 -36093
rect 35394 -36127 35410 -36093
rect 35966 -36127 35982 -36093
rect 36412 -36127 36428 -36093
rect 36984 -36127 37000 -36093
rect 37430 -36127 37446 -36093
rect 38002 -36127 38018 -36093
rect 38448 -36127 38464 -36093
rect 39020 -36127 39036 -36093
rect 39466 -36127 39482 -36093
rect 40038 -36127 40054 -36093
rect 40484 -36127 40500 -36093
rect 41056 -36127 41072 -36093
rect 41502 -36127 41518 -36093
rect 42074 -36127 42090 -36093
rect 42520 -36127 42536 -36093
rect 43092 -36127 43108 -36093
rect 43538 -36127 43554 -36093
rect 44110 -36127 44126 -36093
rect 44556 -36127 44572 -36093
rect 45128 -36127 45144 -36093
rect 45574 -36127 45590 -36093
rect 46146 -36127 46162 -36093
rect 46592 -36127 46608 -36093
rect 47164 -36127 47180 -36093
rect 32706 -36494 32796 -36464
rect 32706 -36528 32734 -36494
rect 32768 -36528 32796 -36494
rect 32706 -36556 32796 -36528
rect 33724 -36494 33814 -36464
rect 33724 -36528 33752 -36494
rect 33786 -36528 33814 -36494
rect 33724 -36556 33814 -36528
rect 34742 -36494 34832 -36464
rect 34742 -36528 34770 -36494
rect 34804 -36528 34832 -36494
rect 34742 -36556 34832 -36528
rect 35760 -36494 35850 -36464
rect 35760 -36528 35788 -36494
rect 35822 -36528 35850 -36494
rect 35760 -36556 35850 -36528
rect 36778 -36494 36868 -36464
rect 36778 -36528 36806 -36494
rect 36840 -36528 36868 -36494
rect 36778 -36556 36868 -36528
rect 37796 -36494 37886 -36464
rect 37796 -36528 37824 -36494
rect 37858 -36528 37886 -36494
rect 37796 -36556 37886 -36528
rect 38814 -36494 38904 -36464
rect 38814 -36528 38842 -36494
rect 38876 -36528 38904 -36494
rect 38814 -36556 38904 -36528
rect 39832 -36494 39922 -36464
rect 39832 -36528 39860 -36494
rect 39894 -36528 39922 -36494
rect 39832 -36556 39922 -36528
rect 40850 -36494 40940 -36464
rect 40850 -36528 40878 -36494
rect 40912 -36528 40940 -36494
rect 40850 -36556 40940 -36528
rect 41868 -36494 41958 -36464
rect 41868 -36528 41896 -36494
rect 41930 -36528 41958 -36494
rect 41868 -36556 41958 -36528
rect 42886 -36494 42976 -36464
rect 42886 -36528 42914 -36494
rect 42948 -36528 42976 -36494
rect 42886 -36556 42976 -36528
rect 43904 -36494 43994 -36464
rect 43904 -36528 43932 -36494
rect 43966 -36528 43994 -36494
rect 43904 -36556 43994 -36528
rect 44922 -36494 45012 -36464
rect 44922 -36528 44950 -36494
rect 44984 -36528 45012 -36494
rect 44922 -36556 45012 -36528
rect 45940 -36494 46030 -36464
rect 45940 -36528 45968 -36494
rect 46002 -36528 46030 -36494
rect 45940 -36556 46030 -36528
rect 46958 -36494 47048 -36464
rect 46958 -36528 46986 -36494
rect 47020 -36528 47048 -36494
rect 46958 -36556 47048 -36528
rect 47976 -36494 48066 -36464
rect 47976 -36528 48004 -36494
rect 48038 -36528 48066 -36494
rect 47976 -36556 48066 -36528
rect 28108 -36804 28198 -36774
rect 28108 -36838 28136 -36804
rect 28170 -36838 28198 -36804
rect 28108 -36866 28198 -36838
rect 29126 -36804 29216 -36774
rect 29126 -36838 29154 -36804
rect 29188 -36838 29216 -36804
rect 29126 -36866 29216 -36838
rect 30144 -36804 30234 -36774
rect 30144 -36838 30172 -36804
rect 30206 -36838 30234 -36804
rect 30144 -36866 30234 -36838
rect 31162 -36804 31252 -36774
rect 31162 -36838 31190 -36804
rect 31224 -36838 31252 -36804
rect 31162 -36866 31252 -36838
rect 33150 -37003 33166 -36969
rect 33722 -37003 33738 -36969
rect 34168 -37003 34184 -36969
rect 34740 -37003 34756 -36969
rect 35186 -37003 35202 -36969
rect 35758 -37003 35774 -36969
rect 36204 -37003 36220 -36969
rect 36776 -37003 36792 -36969
rect 37222 -37003 37238 -36969
rect 37794 -37003 37810 -36969
rect 38240 -37003 38256 -36969
rect 38812 -37003 38828 -36969
rect 39258 -37003 39274 -36969
rect 39830 -37003 39846 -36969
rect 40276 -37003 40292 -36969
rect 40848 -37003 40864 -36969
rect 41294 -37003 41310 -36969
rect 41866 -37003 41882 -36969
rect 42312 -37003 42328 -36969
rect 42884 -37003 42900 -36969
rect 43330 -37003 43346 -36969
rect 43902 -37003 43918 -36969
rect 44348 -37003 44364 -36969
rect 44920 -37003 44936 -36969
rect 45366 -37003 45382 -36969
rect 45938 -37003 45954 -36969
rect 46384 -37003 46400 -36969
rect 46956 -37003 46972 -36969
rect 47402 -37003 47418 -36969
rect 47974 -37003 47990 -36969
rect 32918 -37062 32952 -37046
rect 27846 -37107 27862 -37073
rect 28418 -37107 28434 -37073
rect 28864 -37107 28880 -37073
rect 29436 -37107 29452 -37073
rect 29882 -37107 29898 -37073
rect 30454 -37107 30470 -37073
rect 30900 -37107 30916 -37073
rect 31472 -37107 31488 -37073
rect 27614 -37166 27648 -37150
rect 27614 -37758 27648 -37742
rect 28632 -37166 28666 -37150
rect 28632 -37758 28666 -37742
rect 29650 -37166 29684 -37150
rect 29650 -37758 29684 -37742
rect 30668 -37166 30702 -37150
rect 30668 -37758 30702 -37742
rect 31686 -37166 31720 -37150
rect 32918 -37654 32952 -37638
rect 33936 -37062 33970 -37046
rect 33936 -37654 33970 -37638
rect 34954 -37062 34988 -37046
rect 34954 -37654 34988 -37638
rect 35972 -37062 36006 -37046
rect 35972 -37654 36006 -37638
rect 36990 -37062 37024 -37046
rect 36990 -37654 37024 -37638
rect 38008 -37062 38042 -37046
rect 38008 -37654 38042 -37638
rect 39026 -37062 39060 -37046
rect 39026 -37654 39060 -37638
rect 40044 -37062 40078 -37046
rect 40044 -37654 40078 -37638
rect 41062 -37062 41096 -37046
rect 41062 -37654 41096 -37638
rect 42080 -37062 42114 -37046
rect 42080 -37654 42114 -37638
rect 43098 -37062 43132 -37046
rect 43098 -37654 43132 -37638
rect 44116 -37062 44150 -37046
rect 44116 -37654 44150 -37638
rect 45134 -37062 45168 -37046
rect 45134 -37654 45168 -37638
rect 46152 -37062 46186 -37046
rect 46152 -37654 46186 -37638
rect 47170 -37062 47204 -37046
rect 47170 -37654 47204 -37638
rect 48188 -37062 48222 -37046
rect 48188 -37654 48222 -37638
rect 33150 -37731 33166 -37697
rect 33722 -37731 33738 -37697
rect 34168 -37731 34184 -37697
rect 34740 -37731 34756 -37697
rect 35186 -37731 35202 -37697
rect 35758 -37731 35774 -37697
rect 36204 -37731 36220 -37697
rect 36776 -37731 36792 -37697
rect 37222 -37731 37238 -37697
rect 37794 -37731 37810 -37697
rect 38240 -37731 38256 -37697
rect 38812 -37731 38828 -37697
rect 39258 -37731 39274 -37697
rect 39830 -37731 39846 -37697
rect 40276 -37731 40292 -37697
rect 40848 -37731 40864 -37697
rect 41294 -37731 41310 -37697
rect 41866 -37731 41882 -37697
rect 42312 -37731 42328 -37697
rect 42884 -37731 42900 -37697
rect 43330 -37731 43346 -37697
rect 43902 -37731 43918 -37697
rect 44348 -37731 44364 -37697
rect 44920 -37731 44936 -37697
rect 45366 -37731 45382 -37697
rect 45938 -37731 45954 -37697
rect 46384 -37731 46400 -37697
rect 46956 -37731 46972 -37697
rect 47402 -37731 47418 -37697
rect 47974 -37731 47990 -37697
rect 31686 -37758 31720 -37742
rect 27846 -37835 27862 -37801
rect 28418 -37835 28434 -37801
rect 28864 -37835 28880 -37801
rect 29436 -37835 29452 -37801
rect 29882 -37835 29898 -37801
rect 30454 -37835 30470 -37801
rect 30900 -37835 30916 -37801
rect 31472 -37835 31488 -37801
rect 27584 -37958 27674 -37928
rect 27584 -37992 27612 -37958
rect 27646 -37992 27674 -37958
rect 27584 -38020 27674 -37992
rect 28602 -37958 28692 -37928
rect 28602 -37992 28630 -37958
rect 28664 -37992 28692 -37958
rect 28602 -38020 28692 -37992
rect 29620 -37958 29710 -37928
rect 29620 -37992 29648 -37958
rect 29682 -37992 29710 -37958
rect 29620 -38020 29710 -37992
rect 30638 -37958 30728 -37928
rect 30638 -37992 30666 -37958
rect 30700 -37992 30728 -37958
rect 30638 -38020 30728 -37992
rect 32796 -37942 32886 -37912
rect 32796 -37976 32824 -37942
rect 32858 -37976 32886 -37942
rect 32796 -38004 32886 -37976
rect 33814 -37942 33904 -37912
rect 33814 -37976 33842 -37942
rect 33876 -37976 33904 -37942
rect 33814 -38004 33904 -37976
rect 34832 -37942 34922 -37912
rect 34832 -37976 34860 -37942
rect 34894 -37976 34922 -37942
rect 34832 -38004 34922 -37976
rect 35850 -37942 35940 -37912
rect 35850 -37976 35878 -37942
rect 35912 -37976 35940 -37942
rect 35850 -38004 35940 -37976
rect 36868 -37942 36958 -37912
rect 36868 -37976 36896 -37942
rect 36930 -37976 36958 -37942
rect 36868 -38004 36958 -37976
rect 37886 -37942 37976 -37912
rect 37886 -37976 37914 -37942
rect 37948 -37976 37976 -37942
rect 37886 -38004 37976 -37976
rect 38904 -37942 38994 -37912
rect 38904 -37976 38932 -37942
rect 38966 -37976 38994 -37942
rect 38904 -38004 38994 -37976
rect 39922 -37942 40012 -37912
rect 39922 -37976 39950 -37942
rect 39984 -37976 40012 -37942
rect 39922 -38004 40012 -37976
rect 40940 -37942 41030 -37912
rect 40940 -37976 40968 -37942
rect 41002 -37976 41030 -37942
rect 40940 -38004 41030 -37976
rect 41958 -37942 42048 -37912
rect 41958 -37976 41986 -37942
rect 42020 -37976 42048 -37942
rect 41958 -38004 42048 -37976
rect 42976 -37942 43066 -37912
rect 42976 -37976 43004 -37942
rect 43038 -37976 43066 -37942
rect 42976 -38004 43066 -37976
rect 43994 -37942 44084 -37912
rect 43994 -37976 44022 -37942
rect 44056 -37976 44084 -37942
rect 43994 -38004 44084 -37976
rect 45012 -37942 45102 -37912
rect 45012 -37976 45040 -37942
rect 45074 -37976 45102 -37942
rect 45012 -38004 45102 -37976
rect 46030 -37942 46120 -37912
rect 46030 -37976 46058 -37942
rect 46092 -37976 46120 -37942
rect 46030 -38004 46120 -37976
rect 47048 -37942 47138 -37912
rect 47048 -37976 47076 -37942
rect 47110 -37976 47138 -37942
rect 47048 -38004 47138 -37976
rect 48066 -37942 48156 -37912
rect 48066 -37976 48094 -37942
rect 48128 -37976 48156 -37942
rect 48066 -38004 48156 -37976
rect 27846 -38139 27862 -38105
rect 28418 -38139 28434 -38105
rect 28864 -38139 28880 -38105
rect 29436 -38139 29452 -38105
rect 29882 -38139 29898 -38105
rect 30454 -38139 30470 -38105
rect 30900 -38139 30916 -38105
rect 31472 -38139 31488 -38105
rect 27614 -38198 27648 -38182
rect 27614 -38790 27648 -38774
rect 28632 -38198 28666 -38182
rect 28632 -38790 28666 -38774
rect 29650 -38198 29684 -38182
rect 29650 -38790 29684 -38774
rect 30668 -38198 30702 -38182
rect 30668 -38790 30702 -38774
rect 31686 -38198 31720 -38182
rect 33150 -38259 33166 -38225
rect 33722 -38259 33738 -38225
rect 34168 -38259 34184 -38225
rect 34740 -38259 34756 -38225
rect 35186 -38259 35202 -38225
rect 35758 -38259 35774 -38225
rect 36204 -38259 36220 -38225
rect 36776 -38259 36792 -38225
rect 37222 -38259 37238 -38225
rect 37794 -38259 37810 -38225
rect 38240 -38259 38256 -38225
rect 38812 -38259 38828 -38225
rect 39258 -38259 39274 -38225
rect 39830 -38259 39846 -38225
rect 40276 -38259 40292 -38225
rect 40848 -38259 40864 -38225
rect 41294 -38259 41310 -38225
rect 41866 -38259 41882 -38225
rect 42312 -38259 42328 -38225
rect 42884 -38259 42900 -38225
rect 43330 -38259 43346 -38225
rect 43902 -38259 43918 -38225
rect 44348 -38259 44364 -38225
rect 44920 -38259 44936 -38225
rect 45366 -38259 45382 -38225
rect 45938 -38259 45954 -38225
rect 46384 -38259 46400 -38225
rect 46956 -38259 46972 -38225
rect 47402 -38259 47418 -38225
rect 47974 -38259 47990 -38225
rect 31686 -38790 31720 -38774
rect 32918 -38318 32952 -38302
rect 27846 -38867 27862 -38833
rect 28418 -38867 28434 -38833
rect 28864 -38867 28880 -38833
rect 29436 -38867 29452 -38833
rect 29882 -38867 29898 -38833
rect 30454 -38867 30470 -38833
rect 30900 -38867 30916 -38833
rect 31472 -38867 31488 -38833
rect 32918 -38910 32952 -38894
rect 33936 -38318 33970 -38302
rect 33936 -38910 33970 -38894
rect 34954 -38318 34988 -38302
rect 34954 -38910 34988 -38894
rect 35972 -38318 36006 -38302
rect 35972 -38910 36006 -38894
rect 36990 -38318 37024 -38302
rect 36990 -38910 37024 -38894
rect 38008 -38318 38042 -38302
rect 38008 -38910 38042 -38894
rect 39026 -38318 39060 -38302
rect 39026 -38910 39060 -38894
rect 40044 -38318 40078 -38302
rect 40044 -38910 40078 -38894
rect 41062 -38318 41096 -38302
rect 41062 -38910 41096 -38894
rect 42080 -38318 42114 -38302
rect 42080 -38910 42114 -38894
rect 43098 -38318 43132 -38302
rect 43098 -38910 43132 -38894
rect 44116 -38318 44150 -38302
rect 44116 -38910 44150 -38894
rect 45134 -38318 45168 -38302
rect 45134 -38910 45168 -38894
rect 46152 -38318 46186 -38302
rect 46152 -38910 46186 -38894
rect 47170 -38318 47204 -38302
rect 47170 -38910 47204 -38894
rect 48188 -38318 48222 -38302
rect 48188 -38910 48222 -38894
rect 27594 -38986 27684 -38956
rect 27594 -39020 27622 -38986
rect 27656 -39020 27684 -38986
rect 27594 -39048 27684 -39020
rect 28612 -38986 28702 -38956
rect 28612 -39020 28640 -38986
rect 28674 -39020 28702 -38986
rect 28612 -39048 28702 -39020
rect 29630 -38986 29720 -38956
rect 29630 -39020 29658 -38986
rect 29692 -39020 29720 -38986
rect 29630 -39048 29720 -39020
rect 30648 -38986 30738 -38956
rect 30648 -39020 30676 -38986
rect 30710 -39020 30738 -38986
rect 33150 -38987 33166 -38953
rect 33722 -38987 33738 -38953
rect 34168 -38987 34184 -38953
rect 34740 -38987 34756 -38953
rect 35186 -38987 35202 -38953
rect 35758 -38987 35774 -38953
rect 36204 -38987 36220 -38953
rect 36776 -38987 36792 -38953
rect 37222 -38987 37238 -38953
rect 37794 -38987 37810 -38953
rect 38240 -38987 38256 -38953
rect 38812 -38987 38828 -38953
rect 39258 -38987 39274 -38953
rect 39830 -38987 39846 -38953
rect 40276 -38987 40292 -38953
rect 40848 -38987 40864 -38953
rect 41294 -38987 41310 -38953
rect 41866 -38987 41882 -38953
rect 42312 -38987 42328 -38953
rect 42884 -38987 42900 -38953
rect 43330 -38987 43346 -38953
rect 43902 -38987 43918 -38953
rect 44348 -38987 44364 -38953
rect 44920 -38987 44936 -38953
rect 45366 -38987 45382 -38953
rect 45938 -38987 45954 -38953
rect 46384 -38987 46400 -38953
rect 46956 -38987 46972 -38953
rect 47402 -38987 47418 -38953
rect 47974 -38987 47990 -38953
rect 30648 -39048 30738 -39020
rect 27846 -39171 27862 -39137
rect 28418 -39171 28434 -39137
rect 28864 -39171 28880 -39137
rect 29436 -39171 29452 -39137
rect 29882 -39171 29898 -39137
rect 30454 -39171 30470 -39137
rect 30900 -39171 30916 -39137
rect 31472 -39171 31488 -39137
rect 32820 -39210 32910 -39180
rect 27614 -39230 27648 -39214
rect 27614 -39822 27648 -39806
rect 28632 -39230 28666 -39214
rect 28632 -39822 28666 -39806
rect 29650 -39230 29684 -39214
rect 29650 -39822 29684 -39806
rect 30668 -39230 30702 -39214
rect 30668 -39822 30702 -39806
rect 31686 -39230 31720 -39214
rect 32820 -39244 32848 -39210
rect 32882 -39244 32910 -39210
rect 32820 -39272 32910 -39244
rect 33838 -39210 33928 -39180
rect 33838 -39244 33866 -39210
rect 33900 -39244 33928 -39210
rect 33838 -39272 33928 -39244
rect 34856 -39210 34946 -39180
rect 34856 -39244 34884 -39210
rect 34918 -39244 34946 -39210
rect 34856 -39272 34946 -39244
rect 35874 -39210 35964 -39180
rect 35874 -39244 35902 -39210
rect 35936 -39244 35964 -39210
rect 35874 -39272 35964 -39244
rect 36892 -39210 36982 -39180
rect 36892 -39244 36920 -39210
rect 36954 -39244 36982 -39210
rect 36892 -39272 36982 -39244
rect 37910 -39210 38000 -39180
rect 37910 -39244 37938 -39210
rect 37972 -39244 38000 -39210
rect 37910 -39272 38000 -39244
rect 38928 -39210 39018 -39180
rect 38928 -39244 38956 -39210
rect 38990 -39244 39018 -39210
rect 38928 -39272 39018 -39244
rect 39946 -39210 40036 -39180
rect 39946 -39244 39974 -39210
rect 40008 -39244 40036 -39210
rect 39946 -39272 40036 -39244
rect 40964 -39210 41054 -39180
rect 40964 -39244 40992 -39210
rect 41026 -39244 41054 -39210
rect 40964 -39272 41054 -39244
rect 41982 -39210 42072 -39180
rect 41982 -39244 42010 -39210
rect 42044 -39244 42072 -39210
rect 41982 -39272 42072 -39244
rect 43000 -39210 43090 -39180
rect 43000 -39244 43028 -39210
rect 43062 -39244 43090 -39210
rect 43000 -39272 43090 -39244
rect 44018 -39210 44108 -39180
rect 44018 -39244 44046 -39210
rect 44080 -39244 44108 -39210
rect 44018 -39272 44108 -39244
rect 45036 -39210 45126 -39180
rect 45036 -39244 45064 -39210
rect 45098 -39244 45126 -39210
rect 45036 -39272 45126 -39244
rect 46054 -39210 46144 -39180
rect 46054 -39244 46082 -39210
rect 46116 -39244 46144 -39210
rect 46054 -39272 46144 -39244
rect 47072 -39210 47162 -39180
rect 47072 -39244 47100 -39210
rect 47134 -39244 47162 -39210
rect 47072 -39272 47162 -39244
rect 48090 -39210 48180 -39180
rect 48090 -39244 48118 -39210
rect 48152 -39244 48180 -39210
rect 48090 -39272 48180 -39244
rect 33150 -39515 33166 -39481
rect 33722 -39515 33738 -39481
rect 34168 -39515 34184 -39481
rect 34740 -39515 34756 -39481
rect 35186 -39515 35202 -39481
rect 35758 -39515 35774 -39481
rect 36204 -39515 36220 -39481
rect 36776 -39515 36792 -39481
rect 37222 -39515 37238 -39481
rect 37794 -39515 37810 -39481
rect 38240 -39515 38256 -39481
rect 38812 -39515 38828 -39481
rect 39258 -39515 39274 -39481
rect 39830 -39515 39846 -39481
rect 40276 -39515 40292 -39481
rect 40848 -39515 40864 -39481
rect 41294 -39515 41310 -39481
rect 41866 -39515 41882 -39481
rect 42312 -39515 42328 -39481
rect 42884 -39515 42900 -39481
rect 43330 -39515 43346 -39481
rect 43902 -39515 43918 -39481
rect 44348 -39515 44364 -39481
rect 44920 -39515 44936 -39481
rect 45366 -39515 45382 -39481
rect 45938 -39515 45954 -39481
rect 46384 -39515 46400 -39481
rect 46956 -39515 46972 -39481
rect 47402 -39515 47418 -39481
rect 47974 -39515 47990 -39481
rect 31686 -39822 31720 -39806
rect 32918 -39574 32952 -39558
rect 27846 -39899 27862 -39865
rect 28418 -39899 28434 -39865
rect 28864 -39899 28880 -39865
rect 29436 -39899 29452 -39865
rect 29882 -39899 29898 -39865
rect 30454 -39899 30470 -39865
rect 30900 -39899 30916 -39865
rect 31472 -39899 31488 -39865
rect 27584 -40014 27674 -39984
rect 27584 -40048 27612 -40014
rect 27646 -40048 27674 -40014
rect 27584 -40076 27674 -40048
rect 28602 -40014 28692 -39984
rect 28602 -40048 28630 -40014
rect 28664 -40048 28692 -40014
rect 28602 -40076 28692 -40048
rect 29620 -40014 29710 -39984
rect 29620 -40048 29648 -40014
rect 29682 -40048 29710 -40014
rect 29620 -40076 29710 -40048
rect 30638 -40014 30728 -39984
rect 30638 -40048 30666 -40014
rect 30700 -40048 30728 -40014
rect 30638 -40076 30728 -40048
rect 32918 -40166 32952 -40150
rect 33936 -39574 33970 -39558
rect 33936 -40166 33970 -40150
rect 34954 -39574 34988 -39558
rect 34954 -40166 34988 -40150
rect 35972 -39574 36006 -39558
rect 35972 -40166 36006 -40150
rect 36990 -39574 37024 -39558
rect 36990 -40166 37024 -40150
rect 38008 -39574 38042 -39558
rect 38008 -40166 38042 -40150
rect 39026 -39574 39060 -39558
rect 39026 -40166 39060 -40150
rect 40044 -39574 40078 -39558
rect 40044 -40166 40078 -40150
rect 41062 -39574 41096 -39558
rect 41062 -40166 41096 -40150
rect 42080 -39574 42114 -39558
rect 42080 -40166 42114 -40150
rect 43098 -39574 43132 -39558
rect 43098 -40166 43132 -40150
rect 44116 -39574 44150 -39558
rect 44116 -40166 44150 -40150
rect 45134 -39574 45168 -39558
rect 45134 -40166 45168 -40150
rect 46152 -39574 46186 -39558
rect 46152 -40166 46186 -40150
rect 47170 -39574 47204 -39558
rect 47170 -40166 47204 -40150
rect 48188 -39574 48222 -39558
rect 48188 -40166 48222 -40150
rect 27846 -40203 27862 -40169
rect 28418 -40203 28434 -40169
rect 28864 -40203 28880 -40169
rect 29436 -40203 29452 -40169
rect 29882 -40203 29898 -40169
rect 30454 -40203 30470 -40169
rect 30900 -40203 30916 -40169
rect 31472 -40203 31488 -40169
rect 33150 -40243 33166 -40209
rect 33722 -40243 33738 -40209
rect 34168 -40243 34184 -40209
rect 34740 -40243 34756 -40209
rect 35186 -40243 35202 -40209
rect 35758 -40243 35774 -40209
rect 36204 -40243 36220 -40209
rect 36776 -40243 36792 -40209
rect 37222 -40243 37238 -40209
rect 37794 -40243 37810 -40209
rect 38240 -40243 38256 -40209
rect 38812 -40243 38828 -40209
rect 39258 -40243 39274 -40209
rect 39830 -40243 39846 -40209
rect 40276 -40243 40292 -40209
rect 40848 -40243 40864 -40209
rect 41294 -40243 41310 -40209
rect 41866 -40243 41882 -40209
rect 42312 -40243 42328 -40209
rect 42884 -40243 42900 -40209
rect 43330 -40243 43346 -40209
rect 43902 -40243 43918 -40209
rect 44348 -40243 44364 -40209
rect 44920 -40243 44936 -40209
rect 45366 -40243 45382 -40209
rect 45938 -40243 45954 -40209
rect 46384 -40243 46400 -40209
rect 46956 -40243 46972 -40209
rect 47402 -40243 47418 -40209
rect 47974 -40243 47990 -40209
rect 27614 -40262 27648 -40246
rect 27614 -40854 27648 -40838
rect 28632 -40262 28666 -40246
rect 28632 -40854 28666 -40838
rect 29650 -40262 29684 -40246
rect 29650 -40854 29684 -40838
rect 30668 -40262 30702 -40246
rect 30668 -40854 30702 -40838
rect 31686 -40262 31720 -40246
rect 32684 -40454 32774 -40424
rect 32684 -40488 32712 -40454
rect 32746 -40488 32774 -40454
rect 32684 -40516 32774 -40488
rect 33702 -40454 33792 -40424
rect 33702 -40488 33730 -40454
rect 33764 -40488 33792 -40454
rect 33702 -40516 33792 -40488
rect 34720 -40454 34810 -40424
rect 34720 -40488 34748 -40454
rect 34782 -40488 34810 -40454
rect 34720 -40516 34810 -40488
rect 35738 -40454 35828 -40424
rect 35738 -40488 35766 -40454
rect 35800 -40488 35828 -40454
rect 35738 -40516 35828 -40488
rect 36756 -40454 36846 -40424
rect 36756 -40488 36784 -40454
rect 36818 -40488 36846 -40454
rect 36756 -40516 36846 -40488
rect 37774 -40454 37864 -40424
rect 37774 -40488 37802 -40454
rect 37836 -40488 37864 -40454
rect 37774 -40516 37864 -40488
rect 38792 -40454 38882 -40424
rect 38792 -40488 38820 -40454
rect 38854 -40488 38882 -40454
rect 38792 -40516 38882 -40488
rect 39810 -40454 39900 -40424
rect 39810 -40488 39838 -40454
rect 39872 -40488 39900 -40454
rect 39810 -40516 39900 -40488
rect 40828 -40454 40918 -40424
rect 40828 -40488 40856 -40454
rect 40890 -40488 40918 -40454
rect 40828 -40516 40918 -40488
rect 41846 -40454 41936 -40424
rect 41846 -40488 41874 -40454
rect 41908 -40488 41936 -40454
rect 41846 -40516 41936 -40488
rect 42864 -40454 42954 -40424
rect 42864 -40488 42892 -40454
rect 42926 -40488 42954 -40454
rect 42864 -40516 42954 -40488
rect 43882 -40454 43972 -40424
rect 43882 -40488 43910 -40454
rect 43944 -40488 43972 -40454
rect 43882 -40516 43972 -40488
rect 44900 -40454 44990 -40424
rect 44900 -40488 44928 -40454
rect 44962 -40488 44990 -40454
rect 44900 -40516 44990 -40488
rect 45918 -40454 46008 -40424
rect 45918 -40488 45946 -40454
rect 45980 -40488 46008 -40454
rect 45918 -40516 46008 -40488
rect 46936 -40454 47026 -40424
rect 46936 -40488 46964 -40454
rect 46998 -40488 47026 -40454
rect 46936 -40516 47026 -40488
rect 47954 -40454 48044 -40424
rect 47954 -40488 47982 -40454
rect 48016 -40488 48044 -40454
rect 47954 -40516 48044 -40488
rect 33150 -40771 33166 -40737
rect 33722 -40771 33738 -40737
rect 34168 -40771 34184 -40737
rect 34740 -40771 34756 -40737
rect 35186 -40771 35202 -40737
rect 35758 -40771 35774 -40737
rect 36204 -40771 36220 -40737
rect 36776 -40771 36792 -40737
rect 37222 -40771 37238 -40737
rect 37794 -40771 37810 -40737
rect 38240 -40771 38256 -40737
rect 38812 -40771 38828 -40737
rect 39258 -40771 39274 -40737
rect 39830 -40771 39846 -40737
rect 40276 -40771 40292 -40737
rect 40848 -40771 40864 -40737
rect 41294 -40771 41310 -40737
rect 41866 -40771 41882 -40737
rect 42312 -40771 42328 -40737
rect 42884 -40771 42900 -40737
rect 43330 -40771 43346 -40737
rect 43902 -40771 43918 -40737
rect 44348 -40771 44364 -40737
rect 44920 -40771 44936 -40737
rect 45366 -40771 45382 -40737
rect 45938 -40771 45954 -40737
rect 46384 -40771 46400 -40737
rect 46956 -40771 46972 -40737
rect 47402 -40771 47418 -40737
rect 47974 -40771 47990 -40737
rect 31686 -40854 31720 -40838
rect 32918 -40830 32952 -40814
rect 27846 -40931 27862 -40897
rect 28418 -40931 28434 -40897
rect 28864 -40931 28880 -40897
rect 29436 -40931 29452 -40897
rect 29882 -40931 29898 -40897
rect 30454 -40931 30470 -40897
rect 30900 -40931 30916 -40897
rect 31472 -40931 31488 -40897
rect 28108 -41166 28198 -41136
rect 28108 -41200 28136 -41166
rect 28170 -41200 28198 -41166
rect 28108 -41228 28198 -41200
rect 29126 -41166 29216 -41136
rect 29126 -41200 29154 -41166
rect 29188 -41200 29216 -41166
rect 29126 -41228 29216 -41200
rect 30144 -41166 30234 -41136
rect 30144 -41200 30172 -41166
rect 30206 -41200 30234 -41166
rect 30144 -41228 30234 -41200
rect 31162 -41166 31252 -41136
rect 31162 -41200 31190 -41166
rect 31224 -41200 31252 -41166
rect 31162 -41228 31252 -41200
rect 32918 -41422 32952 -41406
rect 33936 -40830 33970 -40814
rect 33936 -41422 33970 -41406
rect 34954 -40830 34988 -40814
rect 34954 -41422 34988 -41406
rect 35972 -40830 36006 -40814
rect 35972 -41422 36006 -41406
rect 36990 -40830 37024 -40814
rect 36990 -41422 37024 -41406
rect 38008 -40830 38042 -40814
rect 38008 -41422 38042 -41406
rect 39026 -40830 39060 -40814
rect 39026 -41422 39060 -41406
rect 40044 -40830 40078 -40814
rect 40044 -41422 40078 -41406
rect 41062 -40830 41096 -40814
rect 41062 -41422 41096 -41406
rect 42080 -40830 42114 -40814
rect 42080 -41422 42114 -41406
rect 43098 -40830 43132 -40814
rect 43098 -41422 43132 -41406
rect 44116 -40830 44150 -40814
rect 44116 -41422 44150 -41406
rect 45134 -40830 45168 -40814
rect 45134 -41422 45168 -41406
rect 46152 -40830 46186 -40814
rect 46152 -41422 46186 -41406
rect 47170 -40830 47204 -40814
rect 47170 -41422 47204 -41406
rect 48188 -40830 48222 -40814
rect 48188 -41422 48222 -41406
rect 33150 -41499 33166 -41465
rect 33722 -41499 33738 -41465
rect 34168 -41499 34184 -41465
rect 34740 -41499 34756 -41465
rect 35186 -41499 35202 -41465
rect 35758 -41499 35774 -41465
rect 36204 -41499 36220 -41465
rect 36776 -41499 36792 -41465
rect 37222 -41499 37238 -41465
rect 37794 -41499 37810 -41465
rect 38240 -41499 38256 -41465
rect 38812 -41499 38828 -41465
rect 39258 -41499 39274 -41465
rect 39830 -41499 39846 -41465
rect 40276 -41499 40292 -41465
rect 40848 -41499 40864 -41465
rect 41294 -41499 41310 -41465
rect 41866 -41499 41882 -41465
rect 42312 -41499 42328 -41465
rect 42884 -41499 42900 -41465
rect 43330 -41499 43346 -41465
rect 43902 -41499 43918 -41465
rect 44348 -41499 44364 -41465
rect 44920 -41499 44936 -41465
rect 45366 -41499 45382 -41465
rect 45938 -41499 45954 -41465
rect 46384 -41499 46400 -41465
rect 46956 -41499 46972 -41465
rect 47402 -41499 47418 -41465
rect 47974 -41499 47990 -41465
rect 25822 -42326 25922 -42164
rect 50166 -42326 50266 -42164
rect 52156 -39142 52256 -38980
rect 55420 -39142 55520 -38980
rect 52562 -39633 52578 -39599
rect 52798 -39633 52814 -39599
rect 53020 -39633 53036 -39599
rect 53256 -39633 53272 -39599
rect 53478 -39633 53494 -39599
rect 53714 -39633 53730 -39599
rect 53936 -39633 53952 -39599
rect 54172 -39633 54188 -39599
rect 54394 -39633 54410 -39599
rect 54630 -39633 54646 -39599
rect 54852 -39633 54868 -39599
rect 55088 -39633 55104 -39599
rect 52442 -39692 52476 -39676
rect 52442 -39884 52476 -39868
rect 52900 -39692 52934 -39676
rect 52900 -39884 52934 -39868
rect 53358 -39692 53392 -39676
rect 53358 -39884 53392 -39868
rect 53816 -39692 53850 -39676
rect 53816 -39884 53850 -39868
rect 54274 -39692 54308 -39676
rect 54274 -39884 54308 -39868
rect 54732 -39692 54766 -39676
rect 54732 -39884 54766 -39868
rect 55190 -39692 55224 -39676
rect 55190 -39884 55224 -39868
rect 52562 -39961 52578 -39927
rect 52798 -39961 52814 -39927
rect 53020 -39961 53036 -39927
rect 53256 -39961 53272 -39927
rect 53478 -39961 53494 -39927
rect 53714 -39961 53730 -39927
rect 53936 -39961 53952 -39927
rect 54172 -39961 54188 -39927
rect 54394 -39961 54410 -39927
rect 54630 -39961 54646 -39927
rect 54852 -39961 54868 -39927
rect 55088 -39961 55104 -39927
rect 52581 -40516 52597 -40482
rect 52697 -40516 52713 -40482
rect 52839 -40516 52855 -40482
rect 52955 -40516 52971 -40482
rect 53097 -40516 53113 -40482
rect 53213 -40516 53229 -40482
rect 53355 -40516 53371 -40482
rect 53471 -40516 53487 -40482
rect 53613 -40516 53629 -40482
rect 53729 -40516 53745 -40482
rect 53871 -40516 53887 -40482
rect 53987 -40516 54003 -40482
rect 54129 -40516 54145 -40482
rect 54245 -40516 54261 -40482
rect 54387 -40516 54403 -40482
rect 54503 -40516 54519 -40482
rect 54645 -40516 54661 -40482
rect 54761 -40516 54777 -40482
rect 54903 -40516 54919 -40482
rect 55019 -40516 55035 -40482
rect 52501 -40575 52535 -40559
rect 52501 -40967 52535 -40951
rect 52759 -40575 52793 -40559
rect 52759 -40967 52793 -40951
rect 53017 -40575 53051 -40559
rect 53017 -40967 53051 -40951
rect 53275 -40575 53309 -40559
rect 53275 -40967 53309 -40951
rect 53533 -40575 53567 -40559
rect 53533 -40967 53567 -40951
rect 53791 -40575 53825 -40559
rect 53791 -40967 53825 -40951
rect 54049 -40575 54083 -40559
rect 54049 -40967 54083 -40951
rect 54307 -40575 54341 -40559
rect 54307 -40967 54341 -40951
rect 54565 -40575 54599 -40559
rect 54565 -40967 54599 -40951
rect 54823 -40575 54857 -40559
rect 54823 -40967 54857 -40951
rect 55081 -40575 55115 -40559
rect 55081 -40967 55115 -40951
rect 52581 -41044 52597 -41010
rect 52697 -41044 52713 -41010
rect 52839 -41044 52855 -41010
rect 52955 -41044 52971 -41010
rect 53097 -41044 53113 -41010
rect 53213 -41044 53229 -41010
rect 53355 -41044 53371 -41010
rect 53471 -41044 53487 -41010
rect 53613 -41044 53629 -41010
rect 53729 -41044 53745 -41010
rect 53871 -41044 53887 -41010
rect 53987 -41044 54003 -41010
rect 54129 -41044 54145 -41010
rect 54245 -41044 54261 -41010
rect 54387 -41044 54403 -41010
rect 54503 -41044 54519 -41010
rect 54645 -41044 54661 -41010
rect 54761 -41044 54777 -41010
rect 54903 -41044 54919 -41010
rect 55019 -41044 55035 -41010
rect 52581 -41376 52597 -41342
rect 52697 -41376 52713 -41342
rect 52839 -41376 52855 -41342
rect 52955 -41376 52971 -41342
rect 53097 -41376 53113 -41342
rect 53213 -41376 53229 -41342
rect 53355 -41376 53371 -41342
rect 53471 -41376 53487 -41342
rect 53613 -41376 53629 -41342
rect 53729 -41376 53745 -41342
rect 53871 -41376 53887 -41342
rect 53987 -41376 54003 -41342
rect 54129 -41376 54145 -41342
rect 54245 -41376 54261 -41342
rect 54387 -41376 54403 -41342
rect 54503 -41376 54519 -41342
rect 54645 -41376 54661 -41342
rect 54761 -41376 54777 -41342
rect 54903 -41376 54919 -41342
rect 55019 -41376 55035 -41342
rect 52501 -41435 52535 -41419
rect 52501 -41827 52535 -41811
rect 52759 -41435 52793 -41419
rect 52759 -41827 52793 -41811
rect 53017 -41435 53051 -41419
rect 53017 -41827 53051 -41811
rect 53275 -41435 53309 -41419
rect 53275 -41827 53309 -41811
rect 53533 -41435 53567 -41419
rect 53533 -41827 53567 -41811
rect 53791 -41435 53825 -41419
rect 53791 -41827 53825 -41811
rect 54049 -41435 54083 -41419
rect 54049 -41827 54083 -41811
rect 54307 -41435 54341 -41419
rect 54307 -41827 54341 -41811
rect 54565 -41435 54599 -41419
rect 54565 -41827 54599 -41811
rect 54823 -41435 54857 -41419
rect 54823 -41827 54857 -41811
rect 55081 -41435 55115 -41419
rect 55081 -41827 55115 -41811
rect 52581 -41904 52597 -41870
rect 52697 -41904 52713 -41870
rect 52839 -41904 52855 -41870
rect 52955 -41904 52971 -41870
rect 53097 -41904 53113 -41870
rect 53213 -41904 53229 -41870
rect 53355 -41904 53371 -41870
rect 53471 -41904 53487 -41870
rect 53613 -41904 53629 -41870
rect 53729 -41904 53745 -41870
rect 53871 -41904 53887 -41870
rect 53987 -41904 54003 -41870
rect 54129 -41904 54145 -41870
rect 54245 -41904 54261 -41870
rect 54387 -41904 54403 -41870
rect 54503 -41904 54519 -41870
rect 54645 -41904 54661 -41870
rect 54761 -41904 54777 -41870
rect 54903 -41904 54919 -41870
rect 55019 -41904 55035 -41870
rect 52156 -42324 52256 -42162
rect 55858 -39142 55958 -38980
rect 58162 -39142 58262 -38980
rect 56150 -39833 56166 -39799
rect 56266 -39833 56282 -39799
rect 56408 -39833 56424 -39799
rect 56524 -39833 56540 -39799
rect 56666 -39833 56682 -39799
rect 56782 -39833 56798 -39799
rect 56924 -39833 56940 -39799
rect 57040 -39833 57056 -39799
rect 57182 -39833 57198 -39799
rect 57298 -39833 57314 -39799
rect 57440 -39833 57456 -39799
rect 57556 -39833 57572 -39799
rect 57698 -39833 57714 -39799
rect 57814 -39833 57830 -39799
rect 56070 -39892 56104 -39876
rect 56070 -40284 56104 -40268
rect 56328 -39892 56362 -39876
rect 56328 -40284 56362 -40268
rect 56586 -39892 56620 -39876
rect 56586 -40284 56620 -40268
rect 56844 -39892 56878 -39876
rect 56844 -40284 56878 -40268
rect 57102 -39892 57136 -39876
rect 57102 -40284 57136 -40268
rect 57360 -39892 57394 -39876
rect 57360 -40284 57394 -40268
rect 57618 -39892 57652 -39876
rect 57618 -40284 57652 -40268
rect 57876 -39892 57910 -39876
rect 57876 -40284 57910 -40268
rect 56150 -40361 56166 -40327
rect 56266 -40361 56282 -40327
rect 56408 -40361 56424 -40327
rect 56524 -40361 56540 -40327
rect 56666 -40361 56682 -40327
rect 56782 -40361 56798 -40327
rect 56924 -40361 56940 -40327
rect 57040 -40361 57056 -40327
rect 57182 -40361 57198 -40327
rect 57298 -40361 57314 -40327
rect 57440 -40361 57456 -40327
rect 57556 -40361 57572 -40327
rect 57698 -40361 57714 -40327
rect 57814 -40361 57830 -40327
rect 56150 -40693 56166 -40659
rect 56266 -40693 56282 -40659
rect 56408 -40693 56424 -40659
rect 56524 -40693 56540 -40659
rect 56666 -40693 56682 -40659
rect 56782 -40693 56798 -40659
rect 56924 -40693 56940 -40659
rect 57040 -40693 57056 -40659
rect 57182 -40693 57198 -40659
rect 57298 -40693 57314 -40659
rect 57440 -40693 57456 -40659
rect 57556 -40693 57572 -40659
rect 57698 -40693 57714 -40659
rect 57814 -40693 57830 -40659
rect 56070 -40752 56104 -40736
rect 56070 -41144 56104 -41128
rect 56328 -40752 56362 -40736
rect 56328 -41144 56362 -41128
rect 56586 -40752 56620 -40736
rect 56586 -41144 56620 -41128
rect 56844 -40752 56878 -40736
rect 56844 -41144 56878 -41128
rect 57102 -40752 57136 -40736
rect 57102 -41144 57136 -41128
rect 57360 -40752 57394 -40736
rect 57360 -41144 57394 -41128
rect 57618 -40752 57652 -40736
rect 57618 -41144 57652 -41128
rect 57876 -40752 57910 -40736
rect 57876 -41144 57910 -41128
rect 56150 -41221 56166 -41187
rect 56266 -41221 56282 -41187
rect 56408 -41221 56424 -41187
rect 56524 -41221 56540 -41187
rect 56666 -41221 56682 -41187
rect 56782 -41221 56798 -41187
rect 56924 -41221 56940 -41187
rect 57040 -41221 57056 -41187
rect 57182 -41221 57198 -41187
rect 57298 -41221 57314 -41187
rect 57440 -41221 57456 -41187
rect 57556 -41221 57572 -41187
rect 57698 -41221 57714 -41187
rect 57814 -41221 57830 -41187
rect 55858 -41530 55958 -41368
rect 58162 -41530 58262 -41368
rect 56104 -41609 56133 -41575
rect 56167 -41609 56225 -41575
rect 56259 -41609 56317 -41575
rect 56351 -41609 56409 -41575
rect 56443 -41609 56501 -41575
rect 56535 -41609 56593 -41575
rect 56627 -41609 56685 -41575
rect 56719 -41609 56777 -41575
rect 56811 -41609 56869 -41575
rect 56903 -41608 56958 -41575
rect 56992 -41608 57050 -41575
rect 57084 -41608 57147 -41575
rect 56903 -41609 57147 -41608
rect 57181 -41609 57239 -41575
rect 57273 -41609 57331 -41575
rect 57365 -41609 57423 -41575
rect 57457 -41609 57515 -41575
rect 57549 -41609 57607 -41575
rect 57641 -41609 57699 -41575
rect 57733 -41609 57791 -41575
rect 57825 -41609 57883 -41575
rect 57917 -41609 57946 -41575
rect 56172 -41651 56214 -41609
rect 56172 -41685 56180 -41651
rect 56172 -41719 56214 -41685
rect 56172 -41753 56180 -41719
rect 56172 -41787 56214 -41753
rect 56172 -41821 56180 -41787
rect 56172 -41837 56214 -41821
rect 56248 -41651 56314 -41643
rect 56248 -41685 56264 -41651
rect 56298 -41685 56314 -41651
rect 56248 -41719 56314 -41685
rect 56248 -41753 56264 -41719
rect 56298 -41753 56314 -41719
rect 56248 -41787 56314 -41753
rect 56248 -41821 56264 -41787
rect 56298 -41821 56314 -41787
rect 56248 -41839 56314 -41821
rect 56448 -41651 56490 -41609
rect 56448 -41685 56456 -41651
rect 56448 -41719 56490 -41685
rect 56448 -41753 56456 -41719
rect 56448 -41787 56490 -41753
rect 56448 -41821 56456 -41787
rect 56448 -41837 56490 -41821
rect 56524 -41651 56590 -41643
rect 56524 -41685 56540 -41651
rect 56574 -41685 56590 -41651
rect 56524 -41719 56590 -41685
rect 56524 -41753 56540 -41719
rect 56574 -41753 56590 -41719
rect 56524 -41787 56590 -41753
rect 56524 -41821 56540 -41787
rect 56574 -41821 56590 -41787
rect 56524 -41839 56590 -41821
rect 56673 -41651 56729 -41609
rect 56673 -41685 56695 -41651
rect 56673 -41719 56729 -41685
rect 56673 -41753 56695 -41719
rect 56673 -41787 56729 -41753
rect 56673 -41821 56695 -41787
rect 56673 -41837 56729 -41821
rect 56763 -41651 56829 -41643
rect 56763 -41685 56779 -41651
rect 56813 -41685 56829 -41651
rect 56763 -41719 56829 -41685
rect 56763 -41753 56779 -41719
rect 56813 -41753 56829 -41719
rect 56763 -41787 56829 -41753
rect 56763 -41821 56779 -41787
rect 56813 -41821 56829 -41787
rect 56763 -41839 56829 -41821
rect 56863 -41651 56915 -41609
rect 56897 -41685 56915 -41651
rect 56863 -41719 56915 -41685
rect 56897 -41753 56915 -41719
rect 56863 -41787 56915 -41753
rect 56897 -41821 56915 -41787
rect 56863 -41837 56915 -41821
rect 57135 -41651 57187 -41609
rect 57135 -41685 57153 -41651
rect 57135 -41719 57187 -41685
rect 57135 -41753 57153 -41719
rect 57135 -41787 57187 -41753
rect 57135 -41821 57153 -41787
rect 57135 -41837 57187 -41821
rect 57221 -41651 57287 -41643
rect 57221 -41685 57237 -41651
rect 57271 -41685 57287 -41651
rect 57221 -41719 57287 -41685
rect 57221 -41753 57237 -41719
rect 57271 -41753 57287 -41719
rect 57221 -41787 57287 -41753
rect 57221 -41821 57237 -41787
rect 57271 -41821 57287 -41787
rect 57221 -41839 57287 -41821
rect 57321 -41651 57377 -41609
rect 57355 -41685 57377 -41651
rect 57321 -41719 57377 -41685
rect 57355 -41753 57377 -41719
rect 57321 -41787 57377 -41753
rect 57355 -41821 57377 -41787
rect 57321 -41837 57377 -41821
rect 57460 -41651 57526 -41643
rect 57460 -41685 57476 -41651
rect 57510 -41685 57526 -41651
rect 57460 -41719 57526 -41685
rect 57460 -41753 57476 -41719
rect 57510 -41753 57526 -41719
rect 57460 -41787 57526 -41753
rect 57460 -41821 57476 -41787
rect 57510 -41821 57526 -41787
rect 57460 -41839 57526 -41821
rect 57560 -41651 57602 -41609
rect 57594 -41685 57602 -41651
rect 57560 -41719 57602 -41685
rect 57594 -41753 57602 -41719
rect 57560 -41787 57602 -41753
rect 57594 -41821 57602 -41787
rect 57560 -41837 57602 -41821
rect 57736 -41651 57802 -41643
rect 57736 -41685 57752 -41651
rect 57786 -41685 57802 -41651
rect 57736 -41719 57802 -41685
rect 57736 -41753 57752 -41719
rect 57786 -41753 57802 -41719
rect 57736 -41787 57802 -41753
rect 57736 -41821 57752 -41787
rect 57786 -41821 57802 -41787
rect 57736 -41839 57802 -41821
rect 57836 -41651 57878 -41609
rect 57870 -41685 57878 -41651
rect 57836 -41719 57878 -41685
rect 57870 -41753 57878 -41719
rect 57836 -41787 57878 -41753
rect 57870 -41821 57878 -41787
rect 57836 -41837 57878 -41821
rect 56268 -41872 56314 -41839
rect 56544 -41872 56590 -41839
rect 56675 -41872 56742 -41871
rect 56168 -41920 56170 -41873
rect 56168 -41921 56184 -41920
rect 56218 -41921 56234 -41873
rect 56268 -41920 56282 -41872
rect 56490 -41887 56510 -41873
rect 56168 -41971 56214 -41955
rect 56268 -41959 56314 -41920
rect 56444 -41921 56460 -41920
rect 56494 -41921 56510 -41887
rect 56544 -41920 56550 -41872
rect 56675 -41920 56682 -41872
rect 56730 -41920 56742 -41872
rect 56168 -42005 56180 -41971
rect 56168 -42039 56214 -42005
rect 56168 -42073 56180 -42039
rect 56168 -42119 56214 -42073
rect 56248 -41971 56314 -41959
rect 56248 -42005 56264 -41971
rect 56298 -42005 56314 -41971
rect 56248 -42039 56314 -42005
rect 56248 -42073 56264 -42039
rect 56298 -42073 56314 -42039
rect 56248 -42085 56314 -42073
rect 56444 -41971 56490 -41955
rect 56544 -41959 56590 -41920
rect 56675 -41921 56692 -41920
rect 56726 -41921 56742 -41920
rect 56675 -41925 56742 -41921
rect 56776 -41959 56810 -41839
rect 56844 -41872 56911 -41871
rect 56844 -41920 56856 -41872
rect 56904 -41920 56911 -41872
rect 56844 -41921 56860 -41920
rect 56894 -41921 56911 -41920
rect 57139 -41886 57206 -41871
rect 57139 -41920 57152 -41886
rect 57186 -41887 57206 -41886
rect 57139 -41921 57156 -41920
rect 57190 -41921 57206 -41887
rect 57240 -41959 57274 -41839
rect 57308 -41874 57375 -41871
rect 57460 -41874 57506 -41839
rect 57736 -41872 57782 -41839
rect 57308 -41887 57330 -41874
rect 57308 -41921 57324 -41887
rect 57308 -41922 57330 -41921
rect 57492 -41922 57506 -41874
rect 57540 -41887 57560 -41873
rect 57540 -41921 57556 -41887
rect 57768 -41920 57782 -41872
rect 57590 -41921 57606 -41920
rect 57308 -41925 57375 -41922
rect 57460 -41959 57506 -41922
rect 56444 -42005 56456 -41971
rect 56444 -42039 56490 -42005
rect 56444 -42073 56456 -42039
rect 56444 -42119 56490 -42073
rect 56524 -41971 56590 -41959
rect 56524 -42005 56540 -41971
rect 56574 -42005 56590 -41971
rect 56524 -42039 56590 -42005
rect 56524 -42073 56540 -42039
rect 56574 -42073 56590 -42039
rect 56524 -42085 56590 -42073
rect 56673 -41975 56735 -41959
rect 56673 -42009 56695 -41975
rect 56729 -42009 56735 -41975
rect 56673 -42043 56735 -42009
rect 56673 -42077 56695 -42043
rect 56729 -42077 56735 -42043
rect 56673 -42119 56735 -42077
rect 56776 -41975 56915 -41959
rect 56776 -41990 56863 -41975
rect 56897 -41990 56915 -41975
rect 56776 -42038 56862 -41990
rect 56910 -42038 56915 -41990
rect 56776 -42043 56915 -42038
rect 56776 -42077 56863 -42043
rect 56897 -42077 56915 -42043
rect 56776 -42085 56915 -42077
rect 57135 -41975 57274 -41959
rect 57135 -41990 57153 -41975
rect 57187 -41990 57274 -41975
rect 57135 -42038 57142 -41990
rect 57190 -42038 57274 -41990
rect 57135 -42043 57274 -42038
rect 57135 -42077 57153 -42043
rect 57187 -42077 57274 -42043
rect 57135 -42085 57274 -42077
rect 57315 -41975 57377 -41959
rect 57315 -42009 57321 -41975
rect 57355 -42009 57377 -41975
rect 57315 -42043 57377 -42009
rect 57315 -42077 57321 -42043
rect 57355 -42077 57377 -42043
rect 56104 -42153 56133 -42119
rect 56167 -42153 56225 -42119
rect 56259 -42153 56317 -42119
rect 56351 -42153 56409 -42119
rect 56443 -42153 56501 -42119
rect 56535 -42153 56593 -42119
rect 56627 -42153 56685 -42119
rect 56719 -42153 56777 -42119
rect 56811 -42153 56869 -42119
rect 56903 -42120 57050 -42119
rect 56903 -42153 56958 -42120
rect 56992 -42152 57050 -42120
rect 57315 -42119 57377 -42077
rect 57460 -41971 57526 -41959
rect 57460 -42005 57476 -41971
rect 57510 -42005 57526 -41971
rect 57460 -42039 57526 -42005
rect 57460 -42073 57476 -42039
rect 57510 -42073 57526 -42039
rect 57460 -42085 57526 -42073
rect 57560 -41971 57606 -41955
rect 57594 -42005 57606 -41971
rect 57560 -42039 57606 -42005
rect 57594 -42073 57606 -42039
rect 57560 -42119 57606 -42073
rect 57736 -41959 57782 -41920
rect 57816 -41921 57832 -41873
rect 57880 -41920 57882 -41873
rect 57866 -41921 57882 -41920
rect 57736 -41971 57802 -41959
rect 57736 -42005 57752 -41971
rect 57786 -42005 57802 -41971
rect 57736 -42039 57802 -42005
rect 57736 -42073 57752 -42039
rect 57786 -42073 57802 -42039
rect 57736 -42085 57802 -42073
rect 57836 -41971 57882 -41955
rect 57870 -42005 57882 -41971
rect 57836 -42039 57882 -42005
rect 57870 -42073 57882 -42039
rect 57836 -42119 57882 -42073
rect 57084 -42152 57147 -42119
rect 56992 -42153 57147 -42152
rect 57181 -42153 57239 -42119
rect 57273 -42153 57331 -42119
rect 57365 -42153 57423 -42119
rect 57457 -42153 57515 -42119
rect 57549 -42153 57607 -42119
rect 57641 -42153 57699 -42119
rect 57733 -42153 57791 -42119
rect 57825 -42153 57883 -42119
rect 57917 -42153 57946 -42119
rect 55420 -42324 55520 -42162
rect 54104 -42418 54200 -42384
rect 55424 -42418 55518 -42384
rect 54104 -42454 54138 -42418
rect 54402 -42482 54452 -42471
rect 54530 -42482 54580 -42471
rect 54658 -42482 54708 -42471
rect 54786 -42477 54836 -42471
rect 54914 -42477 54964 -42471
rect 55042 -42477 55092 -42471
rect 55170 -42477 55220 -42471
rect 55484 -42476 55518 -42418
rect 54776 -42482 55289 -42477
rect 54266 -42487 55289 -42482
rect 54266 -42537 54402 -42487
rect 54452 -42537 54530 -42487
rect 54580 -42537 54658 -42487
rect 54708 -42537 54786 -42487
rect 54836 -42537 54914 -42487
rect 54964 -42537 55042 -42487
rect 55092 -42537 55170 -42487
rect 55220 -42537 55289 -42487
rect 54266 -42542 55289 -42537
rect 54402 -42553 54452 -42542
rect 54530 -42553 54580 -42542
rect 54658 -42553 54708 -42542
rect 54776 -42547 55289 -42542
rect 54786 -42553 54836 -42547
rect 54914 -42553 54964 -42547
rect 55042 -42553 55092 -42547
rect 55170 -42553 55220 -42547
rect 56370 -42487 56470 -42346
rect 57628 -42486 57728 -42346
rect 56972 -42502 57130 -42496
rect 57326 -42502 57366 -42496
rect 54218 -42606 54252 -42590
rect 54201 -42782 54218 -42755
rect 54346 -42606 54380 -42590
rect 54252 -42782 54271 -42755
rect 54201 -42832 54271 -42782
rect 54346 -42798 54380 -42782
rect 54474 -42606 54508 -42590
rect 54474 -42798 54508 -42782
rect 54602 -42606 54636 -42590
rect 54602 -42798 54636 -42782
rect 54730 -42606 54764 -42590
rect 54730 -42798 54764 -42782
rect 54858 -42606 54892 -42590
rect 54858 -42798 54892 -42782
rect 54986 -42606 55020 -42590
rect 54986 -42798 55020 -42782
rect 55114 -42606 55148 -42590
rect 55114 -42798 55148 -42782
rect 55242 -42606 55276 -42590
rect 55370 -42606 55404 -42590
rect 55242 -42798 55276 -42782
rect 55353 -42782 55370 -42761
rect 55404 -42782 55423 -42761
rect 55353 -42832 55423 -42782
rect 54201 -42833 54290 -42832
rect 55346 -42833 55348 -42832
rect 54274 -42839 54324 -42833
rect 55298 -42839 55348 -42833
rect 54274 -42849 54334 -42839
rect 54324 -42899 54334 -42849
rect 54274 -42906 54334 -42899
rect 54201 -42909 54334 -42906
rect 55288 -42849 55348 -42839
rect 55288 -42899 55298 -42849
rect 55288 -42907 55348 -42899
rect 55288 -42909 55423 -42907
rect 54274 -42915 54324 -42909
rect 55298 -42915 55348 -42909
rect 54104 -42966 54138 -42922
rect 55484 -42966 55518 -42922
rect 54104 -43000 54198 -42966
rect 55422 -43000 55518 -42966
rect 55902 -42562 55998 -42528
rect 56186 -42562 56282 -42528
rect 55902 -42624 55936 -42562
rect 56248 -42624 56282 -42562
rect 56059 -42664 56075 -42630
rect 56109 -42664 56125 -42630
rect 56016 -42714 56050 -42698
rect 56016 -42906 56050 -42890
rect 56134 -42714 56168 -42698
rect 56134 -42906 56168 -42890
rect 55902 -42980 55936 -42918
rect 56248 -42980 56282 -42918
rect 55902 -43014 55998 -42980
rect 56186 -43014 56282 -42980
rect 56962 -42512 57140 -42502
rect 56720 -42552 56726 -42512
rect 56786 -42552 56792 -42512
rect 56962 -42552 56972 -42512
rect 57012 -42552 57090 -42512
rect 57130 -42552 57140 -42512
rect 56962 -42562 57140 -42552
rect 56972 -42568 57130 -42562
rect 57326 -42568 57366 -42562
rect 56562 -42628 56596 -42612
rect 56562 -42820 56596 -42804
rect 56680 -42628 56714 -42612
rect 56680 -42820 56714 -42804
rect 56798 -42628 56832 -42612
rect 56798 -42820 56832 -42804
rect 56916 -42628 56950 -42612
rect 57020 -42628 57080 -42568
rect 57020 -42652 57034 -42628
rect 56916 -42820 56950 -42804
rect 57068 -42652 57080 -42628
rect 57152 -42628 57186 -42612
rect 57034 -42820 57068 -42804
rect 57152 -42820 57186 -42804
rect 57270 -42628 57304 -42612
rect 57270 -42820 57304 -42804
rect 57388 -42628 57422 -42612
rect 57388 -42820 57422 -42804
rect 57506 -42628 57540 -42612
rect 57506 -42820 57540 -42804
rect 56558 -42866 56598 -42860
rect 56854 -42868 56894 -42862
rect 57208 -42868 57248 -42862
rect 57506 -42866 57546 -42860
rect 56844 -42874 56978 -42868
rect 56844 -42878 56924 -42874
rect 56844 -42918 56854 -42878
rect 56894 -42918 56924 -42878
rect 56844 -42922 56924 -42918
rect 56972 -42922 56978 -42874
rect 56558 -42932 56598 -42926
rect 56844 -42928 56978 -42922
rect 57142 -42874 57258 -42868
rect 57142 -42922 57144 -42874
rect 57192 -42878 57258 -42874
rect 57192 -42918 57208 -42878
rect 57248 -42918 57258 -42878
rect 57192 -42922 57258 -42918
rect 57142 -42928 57258 -42922
rect 56854 -42934 56894 -42928
rect 57208 -42934 57248 -42928
rect 57506 -42932 57546 -42926
rect 13122 -43318 13222 -43156
rect 50266 -43318 50366 -43156
rect 28530 -43762 28612 -43738
rect 28530 -43796 28554 -43762
rect 28588 -43796 28612 -43762
rect 28530 -43820 28612 -43796
rect 29548 -43762 29630 -43738
rect 29548 -43796 29572 -43762
rect 29606 -43796 29630 -43762
rect 29548 -43820 29630 -43796
rect 30566 -43762 30648 -43738
rect 30566 -43796 30590 -43762
rect 30624 -43796 30648 -43762
rect 30566 -43820 30648 -43796
rect 31584 -43762 31666 -43738
rect 31584 -43796 31608 -43762
rect 31642 -43796 31666 -43762
rect 31584 -43820 31666 -43796
rect 32602 -43762 32684 -43738
rect 32602 -43796 32626 -43762
rect 32660 -43796 32684 -43762
rect 32602 -43820 32684 -43796
rect 33620 -43762 33702 -43738
rect 33620 -43796 33644 -43762
rect 33678 -43796 33702 -43762
rect 33620 -43820 33702 -43796
rect 34638 -43762 34720 -43738
rect 34638 -43796 34662 -43762
rect 34696 -43796 34720 -43762
rect 34638 -43820 34720 -43796
rect 35656 -43762 35738 -43738
rect 35656 -43796 35680 -43762
rect 35714 -43796 35738 -43762
rect 35656 -43820 35738 -43796
rect 36674 -43762 36756 -43738
rect 36674 -43796 36698 -43762
rect 36732 -43796 36756 -43762
rect 36674 -43820 36756 -43796
rect 37692 -43762 37774 -43738
rect 37692 -43796 37716 -43762
rect 37750 -43796 37774 -43762
rect 37692 -43820 37774 -43796
rect 38710 -43762 38792 -43738
rect 38710 -43796 38734 -43762
rect 38768 -43796 38792 -43762
rect 38710 -43820 38792 -43796
rect 39728 -43762 39810 -43738
rect 39728 -43796 39752 -43762
rect 39786 -43796 39810 -43762
rect 39728 -43820 39810 -43796
rect 40746 -43762 40828 -43738
rect 40746 -43796 40770 -43762
rect 40804 -43796 40828 -43762
rect 40746 -43820 40828 -43796
rect 41764 -43762 41846 -43738
rect 41764 -43796 41788 -43762
rect 41822 -43796 41846 -43762
rect 41764 -43820 41846 -43796
rect 42782 -43762 42864 -43738
rect 42782 -43796 42806 -43762
rect 42840 -43796 42864 -43762
rect 42782 -43820 42864 -43796
rect 43800 -43762 43882 -43738
rect 43800 -43796 43824 -43762
rect 43858 -43796 43882 -43762
rect 43800 -43820 43882 -43796
rect 44818 -43762 44900 -43738
rect 44818 -43796 44842 -43762
rect 44876 -43796 44900 -43762
rect 44818 -43820 44900 -43796
rect 45836 -43762 45918 -43738
rect 45836 -43796 45860 -43762
rect 45894 -43796 45918 -43762
rect 45836 -43820 45918 -43796
rect 46854 -43762 46936 -43738
rect 46854 -43796 46878 -43762
rect 46912 -43796 46936 -43762
rect 46854 -43820 46936 -43796
rect 47872 -43762 47954 -43738
rect 47872 -43796 47896 -43762
rect 47930 -43796 47954 -43762
rect 47872 -43820 47954 -43796
rect 28258 -43976 28274 -43942
rect 28830 -43976 28846 -43942
rect 29276 -43976 29292 -43942
rect 29848 -43976 29864 -43942
rect 30294 -43976 30310 -43942
rect 30866 -43976 30882 -43942
rect 31312 -43976 31328 -43942
rect 31884 -43976 31900 -43942
rect 32330 -43976 32346 -43942
rect 32902 -43976 32918 -43942
rect 33348 -43976 33364 -43942
rect 33920 -43976 33936 -43942
rect 34366 -43976 34382 -43942
rect 34938 -43976 34954 -43942
rect 35384 -43976 35400 -43942
rect 35956 -43976 35972 -43942
rect 36402 -43976 36418 -43942
rect 36974 -43976 36990 -43942
rect 37420 -43976 37436 -43942
rect 37992 -43976 38008 -43942
rect 38438 -43976 38454 -43942
rect 39010 -43976 39026 -43942
rect 39456 -43976 39472 -43942
rect 40028 -43976 40044 -43942
rect 40474 -43976 40490 -43942
rect 41046 -43976 41062 -43942
rect 41492 -43976 41508 -43942
rect 42064 -43976 42080 -43942
rect 42510 -43976 42526 -43942
rect 43082 -43976 43098 -43942
rect 43528 -43976 43544 -43942
rect 44100 -43976 44116 -43942
rect 44546 -43976 44562 -43942
rect 45118 -43976 45134 -43942
rect 45564 -43976 45580 -43942
rect 46136 -43976 46152 -43942
rect 46582 -43976 46598 -43942
rect 47154 -43976 47170 -43942
rect 47600 -43976 47616 -43942
rect 48172 -43976 48188 -43942
rect 10296 -56772 10342 -56739
rect 12036 -56772 12106 -56739
rect 10296 -56773 10392 -56772
rect 12010 -56773 12106 -56772
rect 10296 -56835 10330 -56773
rect 12072 -56834 12106 -56773
rect 10490 -56875 10506 -56841
rect 10606 -56875 10622 -56841
rect 10748 -56875 10764 -56841
rect 10864 -56875 10880 -56841
rect 11006 -56875 11022 -56841
rect 11122 -56875 11138 -56841
rect 11264 -56875 11280 -56841
rect 11380 -56875 11396 -56841
rect 11522 -56875 11538 -56841
rect 11638 -56875 11654 -56841
rect 11780 -56875 11796 -56841
rect 11896 -56875 11912 -56841
rect 10410 -56934 10444 -56918
rect 10410 -57326 10444 -57310
rect 10668 -56934 10702 -56918
rect 10668 -57326 10702 -57310
rect 10926 -56934 10960 -56918
rect 10926 -57326 10960 -57310
rect 11184 -56934 11218 -56918
rect 11184 -57326 11218 -57310
rect 11442 -56934 11476 -56918
rect 11442 -57326 11476 -57310
rect 11700 -56934 11734 -56918
rect 11700 -57326 11734 -57310
rect 11958 -56934 11992 -56918
rect 11958 -57326 11992 -57310
rect 10490 -57403 10506 -57369
rect 10606 -57403 10622 -57369
rect 10748 -57403 10764 -57369
rect 10864 -57403 10880 -57369
rect 11006 -57403 11022 -57369
rect 11122 -57403 11138 -57369
rect 11264 -57403 11280 -57369
rect 11380 -57403 11396 -57369
rect 11522 -57403 11538 -57369
rect 11638 -57403 11654 -57369
rect 11780 -57403 11796 -57369
rect 11896 -57403 11912 -57369
rect 10296 -57471 10330 -57409
rect 12180 -57275 12209 -57241
rect 12243 -57275 12301 -57241
rect 12335 -57275 12393 -57241
rect 12427 -57275 12456 -57241
rect 12072 -57471 12106 -57410
rect 10296 -57472 10392 -57471
rect 10296 -57505 10342 -57472
rect 12036 -57504 12106 -57471
rect 12010 -57505 12106 -57504
rect 12246 -57317 12312 -57309
rect 12246 -57351 12262 -57317
rect 12296 -57351 12312 -57317
rect 12246 -57385 12312 -57351
rect 12246 -57419 12262 -57385
rect 12296 -57419 12312 -57385
rect 12246 -57453 12312 -57419
rect 12246 -57487 12262 -57453
rect 12296 -57487 12312 -57453
rect 12246 -57505 12312 -57487
rect 12346 -57317 12388 -57275
rect 12380 -57351 12388 -57317
rect 12346 -57385 12388 -57351
rect 12380 -57419 12388 -57385
rect 12346 -57453 12388 -57419
rect 12380 -57487 12388 -57453
rect 12346 -57503 12388 -57487
rect 12246 -57538 12292 -57505
rect 12286 -57586 12292 -57538
rect 12246 -57625 12292 -57586
rect 12326 -57587 12342 -57539
rect 12390 -57586 12392 -57539
rect 12376 -57587 12392 -57586
rect 12246 -57637 12312 -57625
rect 12246 -57671 12262 -57637
rect 12296 -57671 12312 -57637
rect 10296 -57706 10366 -57672
rect 12036 -57706 12106 -57672
rect 10296 -57768 10330 -57706
rect 12072 -57768 12106 -57706
rect 12246 -57705 12312 -57671
rect 12246 -57739 12262 -57705
rect 12296 -57739 12312 -57705
rect 12246 -57751 12312 -57739
rect 12346 -57637 12392 -57621
rect 12380 -57671 12392 -57637
rect 12346 -57705 12392 -57671
rect 12380 -57739 12392 -57705
rect 10490 -57808 10506 -57774
rect 10606 -57808 10622 -57774
rect 10748 -57808 10764 -57774
rect 10864 -57808 10880 -57774
rect 11006 -57808 11022 -57774
rect 11122 -57808 11138 -57774
rect 11264 -57808 11280 -57774
rect 11380 -57808 11396 -57774
rect 11522 -57808 11538 -57774
rect 11638 -57808 11654 -57774
rect 11780 -57808 11796 -57774
rect 11896 -57808 11912 -57774
rect 10410 -57858 10444 -57842
rect 10410 -58050 10444 -58034
rect 10668 -57858 10702 -57842
rect 10668 -58050 10702 -58034
rect 10926 -57858 10960 -57842
rect 10926 -58050 10960 -58034
rect 11184 -57858 11218 -57842
rect 11184 -58050 11218 -58034
rect 11442 -57858 11476 -57842
rect 11442 -58050 11476 -58034
rect 11700 -57858 11734 -57842
rect 11700 -58050 11734 -58034
rect 11958 -57858 11992 -57842
rect 11958 -58050 11992 -58034
rect 10490 -58118 10506 -58084
rect 10606 -58118 10622 -58084
rect 10748 -58118 10764 -58084
rect 10864 -58118 10880 -58084
rect 11006 -58118 11022 -58084
rect 11122 -58118 11138 -58084
rect 11264 -58118 11280 -58084
rect 11380 -58118 11396 -58084
rect 11522 -58118 11538 -58084
rect 11638 -58118 11654 -58084
rect 11780 -58118 11796 -58084
rect 11896 -58118 11912 -58084
rect 12346 -57785 12392 -57739
rect 12180 -57819 12209 -57785
rect 12243 -57819 12301 -57785
rect 12335 -57819 12393 -57785
rect 12427 -57819 12456 -57785
rect 10296 -58186 10330 -58124
rect 12072 -58186 12106 -58124
rect 10296 -58220 10364 -58186
rect 12038 -58220 12106 -58186
rect 28026 -44026 28060 -44010
rect 16236 -44364 16318 -44340
rect 16236 -44398 16260 -44364
rect 16294 -44398 16318 -44364
rect 16236 -44422 16318 -44398
rect 17254 -44364 17336 -44340
rect 17254 -44398 17278 -44364
rect 17312 -44398 17336 -44364
rect 16492 -44452 16508 -44418
rect 17064 -44452 17080 -44418
rect 17254 -44422 17336 -44398
rect 18272 -44364 18354 -44340
rect 18272 -44398 18296 -44364
rect 18330 -44398 18354 -44364
rect 17510 -44452 17526 -44418
rect 18082 -44452 18098 -44418
rect 18272 -44422 18354 -44398
rect 19290 -44364 19372 -44340
rect 19290 -44398 19314 -44364
rect 19348 -44398 19372 -44364
rect 18528 -44452 18544 -44418
rect 19100 -44452 19116 -44418
rect 19290 -44422 19372 -44398
rect 20308 -44364 20390 -44340
rect 20308 -44398 20332 -44364
rect 20366 -44398 20390 -44364
rect 19546 -44452 19562 -44418
rect 20118 -44452 20134 -44418
rect 20308 -44422 20390 -44398
rect 21326 -44364 21408 -44340
rect 21326 -44398 21350 -44364
rect 21384 -44398 21408 -44364
rect 20564 -44452 20580 -44418
rect 21136 -44452 21152 -44418
rect 21326 -44422 21408 -44398
rect 22344 -44364 22426 -44340
rect 22344 -44398 22368 -44364
rect 22402 -44398 22426 -44364
rect 21582 -44452 21598 -44418
rect 22154 -44452 22170 -44418
rect 22344 -44422 22426 -44398
rect 23362 -44364 23444 -44340
rect 23362 -44398 23386 -44364
rect 23420 -44398 23444 -44364
rect 22600 -44452 22616 -44418
rect 23172 -44452 23188 -44418
rect 23362 -44422 23444 -44398
rect 24380 -44364 24462 -44340
rect 24380 -44398 24404 -44364
rect 24438 -44398 24462 -44364
rect 23618 -44452 23634 -44418
rect 24190 -44452 24206 -44418
rect 24380 -44422 24462 -44398
rect 25408 -44364 25490 -44340
rect 25408 -44398 25432 -44364
rect 25466 -44398 25490 -44364
rect 24636 -44452 24652 -44418
rect 25208 -44452 25224 -44418
rect 25408 -44422 25490 -44398
rect 16260 -44502 16294 -44486
rect 16260 -45094 16294 -45078
rect 17278 -44502 17312 -44486
rect 17278 -45094 17312 -45078
rect 18296 -44502 18330 -44486
rect 18296 -45094 18330 -45078
rect 19314 -44502 19348 -44486
rect 19314 -45094 19348 -45078
rect 20332 -44502 20366 -44486
rect 20332 -45094 20366 -45078
rect 21350 -44502 21384 -44486
rect 21350 -45094 21384 -45078
rect 22368 -44502 22402 -44486
rect 22368 -45094 22402 -45078
rect 23386 -44502 23420 -44486
rect 23386 -45094 23420 -45078
rect 24404 -44502 24438 -44486
rect 24404 -45094 24438 -45078
rect 25422 -44502 25456 -44486
rect 28026 -44618 28060 -44602
rect 29044 -44026 29078 -44010
rect 29044 -44618 29078 -44602
rect 30062 -44026 30096 -44010
rect 30062 -44618 30096 -44602
rect 31080 -44026 31114 -44010
rect 31080 -44618 31114 -44602
rect 32098 -44026 32132 -44010
rect 32098 -44618 32132 -44602
rect 33116 -44026 33150 -44010
rect 33116 -44618 33150 -44602
rect 34134 -44026 34168 -44010
rect 34134 -44618 34168 -44602
rect 35152 -44026 35186 -44010
rect 35152 -44618 35186 -44602
rect 36170 -44026 36204 -44010
rect 36170 -44618 36204 -44602
rect 37188 -44026 37222 -44010
rect 37188 -44618 37222 -44602
rect 38206 -44026 38240 -44010
rect 38206 -44618 38240 -44602
rect 39224 -44026 39258 -44010
rect 39224 -44618 39258 -44602
rect 40242 -44026 40276 -44010
rect 40242 -44618 40276 -44602
rect 41260 -44026 41294 -44010
rect 41260 -44618 41294 -44602
rect 42278 -44026 42312 -44010
rect 42278 -44618 42312 -44602
rect 43296 -44026 43330 -44010
rect 43296 -44618 43330 -44602
rect 44314 -44026 44348 -44010
rect 44314 -44618 44348 -44602
rect 45332 -44026 45366 -44010
rect 45332 -44618 45366 -44602
rect 46350 -44026 46384 -44010
rect 46350 -44618 46384 -44602
rect 47368 -44026 47402 -44010
rect 47368 -44618 47402 -44602
rect 48386 -44026 48420 -44010
rect 48386 -44618 48420 -44602
rect 56370 -43704 56470 -43563
rect 57806 -42562 57902 -42528
rect 58090 -42562 58186 -42528
rect 57806 -42624 57840 -42562
rect 58152 -42624 58186 -42562
rect 57963 -42664 57979 -42630
rect 58013 -42664 58029 -42630
rect 57920 -42714 57954 -42698
rect 57920 -42906 57954 -42890
rect 58038 -42714 58072 -42698
rect 58038 -42906 58072 -42890
rect 57806 -42980 57840 -42918
rect 58152 -42980 58186 -42918
rect 57806 -43014 57902 -42980
rect 58090 -43014 58186 -42980
rect 57628 -43704 57728 -43563
rect 28258 -44686 28274 -44652
rect 28830 -44686 28846 -44652
rect 29276 -44686 29292 -44652
rect 29848 -44686 29864 -44652
rect 30294 -44686 30310 -44652
rect 30866 -44686 30882 -44652
rect 31312 -44686 31328 -44652
rect 31884 -44686 31900 -44652
rect 32330 -44686 32346 -44652
rect 32902 -44686 32918 -44652
rect 33348 -44686 33364 -44652
rect 33920 -44686 33936 -44652
rect 34366 -44686 34382 -44652
rect 34938 -44686 34954 -44652
rect 35384 -44686 35400 -44652
rect 35956 -44686 35972 -44652
rect 36402 -44686 36418 -44652
rect 36974 -44686 36990 -44652
rect 37420 -44686 37436 -44652
rect 37992 -44686 38008 -44652
rect 38438 -44686 38454 -44652
rect 39010 -44686 39026 -44652
rect 39456 -44686 39472 -44652
rect 40028 -44686 40044 -44652
rect 40474 -44686 40490 -44652
rect 41046 -44686 41062 -44652
rect 41492 -44686 41508 -44652
rect 42064 -44686 42080 -44652
rect 42510 -44686 42526 -44652
rect 43082 -44686 43098 -44652
rect 43528 -44686 43544 -44652
rect 44100 -44686 44116 -44652
rect 44546 -44686 44562 -44652
rect 45118 -44686 45134 -44652
rect 45564 -44686 45580 -44652
rect 46136 -44686 46152 -44652
rect 46582 -44686 46598 -44652
rect 47154 -44686 47170 -44652
rect 47600 -44686 47616 -44652
rect 48172 -44686 48188 -44652
rect 28258 -44794 28274 -44760
rect 28830 -44794 28846 -44760
rect 29276 -44794 29292 -44760
rect 29848 -44794 29864 -44760
rect 30294 -44794 30310 -44760
rect 30866 -44794 30882 -44760
rect 31312 -44794 31328 -44760
rect 31884 -44794 31900 -44760
rect 32330 -44794 32346 -44760
rect 32902 -44794 32918 -44760
rect 33348 -44794 33364 -44760
rect 33920 -44794 33936 -44760
rect 34366 -44794 34382 -44760
rect 34938 -44794 34954 -44760
rect 35384 -44794 35400 -44760
rect 35956 -44794 35972 -44760
rect 36402 -44794 36418 -44760
rect 36974 -44794 36990 -44760
rect 37420 -44794 37436 -44760
rect 37992 -44794 38008 -44760
rect 38438 -44794 38454 -44760
rect 39010 -44794 39026 -44760
rect 39456 -44794 39472 -44760
rect 40028 -44794 40044 -44760
rect 40474 -44794 40490 -44760
rect 41046 -44794 41062 -44760
rect 41492 -44794 41508 -44760
rect 42064 -44794 42080 -44760
rect 42510 -44794 42526 -44760
rect 43082 -44794 43098 -44760
rect 43528 -44794 43544 -44760
rect 44100 -44794 44116 -44760
rect 44546 -44794 44562 -44760
rect 45118 -44794 45134 -44760
rect 45564 -44794 45580 -44760
rect 46136 -44794 46152 -44760
rect 46582 -44794 46598 -44760
rect 47154 -44794 47170 -44760
rect 47600 -44794 47616 -44760
rect 48172 -44794 48188 -44760
rect 25422 -45094 25456 -45078
rect 28026 -44844 28060 -44828
rect 16236 -45182 16318 -45158
rect 16492 -45162 16508 -45128
rect 17064 -45162 17080 -45128
rect 16236 -45216 16260 -45182
rect 16294 -45216 16318 -45182
rect 16236 -45240 16318 -45216
rect 17254 -45182 17336 -45158
rect 17510 -45162 17526 -45128
rect 18082 -45162 18098 -45128
rect 17254 -45216 17278 -45182
rect 17312 -45216 17336 -45182
rect 16492 -45270 16508 -45236
rect 17064 -45270 17080 -45236
rect 17254 -45240 17336 -45216
rect 18272 -45182 18354 -45158
rect 18528 -45162 18544 -45128
rect 19100 -45162 19116 -45128
rect 18272 -45216 18296 -45182
rect 18330 -45216 18354 -45182
rect 17510 -45270 17526 -45236
rect 18082 -45270 18098 -45236
rect 18272 -45240 18354 -45216
rect 19290 -45182 19372 -45158
rect 19546 -45162 19562 -45128
rect 20118 -45162 20134 -45128
rect 19290 -45216 19314 -45182
rect 19348 -45216 19372 -45182
rect 18528 -45270 18544 -45236
rect 19100 -45270 19116 -45236
rect 19290 -45240 19372 -45216
rect 20308 -45182 20390 -45158
rect 20564 -45162 20580 -45128
rect 21136 -45162 21152 -45128
rect 20308 -45216 20332 -45182
rect 20366 -45216 20390 -45182
rect 19546 -45270 19562 -45236
rect 20118 -45270 20134 -45236
rect 20308 -45240 20390 -45216
rect 21326 -45182 21408 -45158
rect 21582 -45162 21598 -45128
rect 22154 -45162 22170 -45128
rect 21326 -45216 21350 -45182
rect 21384 -45216 21408 -45182
rect 20564 -45270 20580 -45236
rect 21136 -45270 21152 -45236
rect 21326 -45240 21408 -45216
rect 22344 -45182 22426 -45158
rect 22600 -45162 22616 -45128
rect 23172 -45162 23188 -45128
rect 22344 -45216 22368 -45182
rect 22402 -45216 22426 -45182
rect 21582 -45270 21598 -45236
rect 22154 -45270 22170 -45236
rect 22344 -45240 22426 -45216
rect 23362 -45182 23444 -45158
rect 23618 -45162 23634 -45128
rect 24190 -45162 24206 -45128
rect 23362 -45216 23386 -45182
rect 23420 -45216 23444 -45182
rect 22600 -45270 22616 -45236
rect 23172 -45270 23188 -45236
rect 23362 -45240 23444 -45216
rect 24380 -45182 24462 -45158
rect 24636 -45162 24652 -45128
rect 25208 -45162 25224 -45128
rect 24380 -45216 24404 -45182
rect 24438 -45216 24462 -45182
rect 23618 -45270 23634 -45236
rect 24190 -45270 24206 -45236
rect 24380 -45240 24462 -45216
rect 25408 -45182 25490 -45158
rect 25408 -45216 25432 -45182
rect 25466 -45216 25490 -45182
rect 24636 -45270 24652 -45236
rect 25208 -45270 25224 -45236
rect 25408 -45240 25490 -45216
rect 21852 -45272 21912 -45270
rect 16260 -45320 16294 -45304
rect 16260 -45912 16294 -45896
rect 17278 -45320 17312 -45304
rect 17278 -45912 17312 -45896
rect 18296 -45320 18330 -45304
rect 18296 -45912 18330 -45896
rect 19314 -45320 19348 -45304
rect 19314 -45912 19348 -45896
rect 20332 -45320 20366 -45304
rect 20332 -45912 20366 -45896
rect 21350 -45320 21384 -45304
rect 21350 -45912 21384 -45896
rect 22368 -45320 22402 -45304
rect 22368 -45912 22402 -45896
rect 23386 -45320 23420 -45304
rect 23386 -45912 23420 -45896
rect 24404 -45320 24438 -45304
rect 24404 -45912 24438 -45896
rect 25422 -45320 25456 -45304
rect 28026 -45436 28060 -45420
rect 29044 -44844 29078 -44828
rect 29044 -45436 29078 -45420
rect 30062 -44844 30096 -44828
rect 30062 -45436 30096 -45420
rect 31080 -44844 31114 -44828
rect 31080 -45436 31114 -45420
rect 32098 -44844 32132 -44828
rect 32098 -45436 32132 -45420
rect 33116 -44844 33150 -44828
rect 33116 -45436 33150 -45420
rect 34134 -44844 34168 -44828
rect 34134 -45436 34168 -45420
rect 35152 -44844 35186 -44828
rect 35152 -45436 35186 -45420
rect 36170 -44844 36204 -44828
rect 36170 -45436 36204 -45420
rect 37188 -44844 37222 -44828
rect 37188 -45436 37222 -45420
rect 38206 -44844 38240 -44828
rect 38206 -45436 38240 -45420
rect 39224 -44844 39258 -44828
rect 39224 -45436 39258 -45420
rect 40242 -44844 40276 -44828
rect 40242 -45436 40276 -45420
rect 41260 -44844 41294 -44828
rect 41260 -45436 41294 -45420
rect 42278 -44844 42312 -44828
rect 42278 -45436 42312 -45420
rect 43296 -44844 43330 -44828
rect 43296 -45436 43330 -45420
rect 44314 -44844 44348 -44828
rect 44314 -45436 44348 -45420
rect 45332 -44844 45366 -44828
rect 45332 -45436 45366 -45420
rect 46350 -44844 46384 -44828
rect 46350 -45436 46384 -45420
rect 47368 -44844 47402 -44828
rect 47368 -45436 47402 -45420
rect 48386 -44844 48420 -44828
rect 48386 -45436 48420 -45420
rect 28258 -45504 28274 -45470
rect 28830 -45504 28846 -45470
rect 29276 -45504 29292 -45470
rect 29848 -45504 29864 -45470
rect 30294 -45504 30310 -45470
rect 30866 -45504 30882 -45470
rect 31312 -45504 31328 -45470
rect 31884 -45504 31900 -45470
rect 32330 -45504 32346 -45470
rect 32902 -45504 32918 -45470
rect 33348 -45504 33364 -45470
rect 33920 -45504 33936 -45470
rect 34366 -45504 34382 -45470
rect 34938 -45504 34954 -45470
rect 35384 -45504 35400 -45470
rect 35956 -45504 35972 -45470
rect 36402 -45504 36418 -45470
rect 36974 -45504 36990 -45470
rect 37420 -45504 37436 -45470
rect 37992 -45504 38008 -45470
rect 38438 -45504 38454 -45470
rect 39010 -45504 39026 -45470
rect 39456 -45504 39472 -45470
rect 40028 -45504 40044 -45470
rect 40474 -45504 40490 -45470
rect 41046 -45504 41062 -45470
rect 41492 -45504 41508 -45470
rect 42064 -45504 42080 -45470
rect 42510 -45504 42526 -45470
rect 43082 -45504 43098 -45470
rect 43528 -45504 43544 -45470
rect 44100 -45504 44116 -45470
rect 44546 -45504 44562 -45470
rect 45118 -45504 45134 -45470
rect 45564 -45504 45580 -45470
rect 46136 -45504 46152 -45470
rect 46582 -45504 46598 -45470
rect 47154 -45504 47170 -45470
rect 47600 -45504 47616 -45470
rect 48172 -45504 48188 -45470
rect 28542 -45788 28624 -45764
rect 28542 -45822 28566 -45788
rect 28600 -45822 28624 -45788
rect 28542 -45846 28624 -45822
rect 29560 -45788 29642 -45764
rect 29560 -45822 29584 -45788
rect 29618 -45822 29642 -45788
rect 29560 -45846 29642 -45822
rect 30578 -45788 30660 -45764
rect 30578 -45822 30602 -45788
rect 30636 -45822 30660 -45788
rect 30578 -45846 30660 -45822
rect 31596 -45788 31678 -45764
rect 31596 -45822 31620 -45788
rect 31654 -45822 31678 -45788
rect 31596 -45846 31678 -45822
rect 32614 -45788 32696 -45764
rect 32614 -45822 32638 -45788
rect 32672 -45822 32696 -45788
rect 32614 -45846 32696 -45822
rect 33632 -45788 33714 -45764
rect 33632 -45822 33656 -45788
rect 33690 -45822 33714 -45788
rect 33632 -45846 33714 -45822
rect 34650 -45788 34732 -45764
rect 34650 -45822 34674 -45788
rect 34708 -45822 34732 -45788
rect 34650 -45846 34732 -45822
rect 35668 -45788 35750 -45764
rect 35668 -45822 35692 -45788
rect 35726 -45822 35750 -45788
rect 35668 -45846 35750 -45822
rect 36686 -45788 36768 -45764
rect 36686 -45822 36710 -45788
rect 36744 -45822 36768 -45788
rect 36686 -45846 36768 -45822
rect 37704 -45788 37786 -45764
rect 37704 -45822 37728 -45788
rect 37762 -45822 37786 -45788
rect 37704 -45846 37786 -45822
rect 38722 -45788 38804 -45764
rect 38722 -45822 38746 -45788
rect 38780 -45822 38804 -45788
rect 38722 -45846 38804 -45822
rect 39740 -45788 39822 -45764
rect 39740 -45822 39764 -45788
rect 39798 -45822 39822 -45788
rect 39740 -45846 39822 -45822
rect 40758 -45788 40840 -45764
rect 40758 -45822 40782 -45788
rect 40816 -45822 40840 -45788
rect 40758 -45846 40840 -45822
rect 41776 -45788 41858 -45764
rect 41776 -45822 41800 -45788
rect 41834 -45822 41858 -45788
rect 41776 -45846 41858 -45822
rect 42794 -45788 42876 -45764
rect 42794 -45822 42818 -45788
rect 42852 -45822 42876 -45788
rect 42794 -45846 42876 -45822
rect 43812 -45788 43894 -45764
rect 43812 -45822 43836 -45788
rect 43870 -45822 43894 -45788
rect 43812 -45846 43894 -45822
rect 44830 -45788 44912 -45764
rect 44830 -45822 44854 -45788
rect 44888 -45822 44912 -45788
rect 44830 -45846 44912 -45822
rect 45848 -45788 45930 -45764
rect 45848 -45822 45872 -45788
rect 45906 -45822 45930 -45788
rect 45848 -45846 45930 -45822
rect 46866 -45788 46948 -45764
rect 46866 -45822 46890 -45788
rect 46924 -45822 46948 -45788
rect 46866 -45846 46948 -45822
rect 47884 -45788 47966 -45764
rect 47884 -45822 47908 -45788
rect 47942 -45822 47966 -45788
rect 47884 -45846 47966 -45822
rect 25422 -45912 25456 -45896
rect 17784 -45946 17844 -45944
rect 18798 -45946 18858 -45944
rect 22872 -45946 22932 -45944
rect 23888 -45946 23948 -45944
rect 16236 -46000 16318 -45976
rect 16492 -45980 16508 -45946
rect 17064 -45980 17080 -45946
rect 16236 -46034 16260 -46000
rect 16294 -46034 16318 -46000
rect 16236 -46058 16318 -46034
rect 17254 -46000 17336 -45976
rect 17510 -45980 17526 -45946
rect 18082 -45980 18098 -45946
rect 17254 -46034 17278 -46000
rect 17312 -46034 17336 -46000
rect 16492 -46088 16508 -46054
rect 17064 -46088 17080 -46054
rect 17254 -46058 17336 -46034
rect 18272 -46000 18354 -45976
rect 18528 -45980 18544 -45946
rect 19100 -45980 19116 -45946
rect 18272 -46034 18296 -46000
rect 18330 -46034 18354 -46000
rect 17510 -46088 17526 -46054
rect 18082 -46088 18098 -46054
rect 18272 -46058 18354 -46034
rect 19290 -46000 19372 -45976
rect 19546 -45980 19562 -45946
rect 20118 -45980 20134 -45946
rect 19290 -46034 19314 -46000
rect 19348 -46034 19372 -46000
rect 18528 -46088 18544 -46054
rect 19100 -46088 19116 -46054
rect 19290 -46058 19372 -46034
rect 20308 -46000 20390 -45976
rect 20564 -45980 20580 -45946
rect 21136 -45980 21152 -45946
rect 20308 -46034 20332 -46000
rect 20366 -46034 20390 -46000
rect 19546 -46088 19562 -46054
rect 20118 -46088 20134 -46054
rect 20308 -46058 20390 -46034
rect 21326 -46000 21408 -45976
rect 21582 -45980 21598 -45946
rect 22154 -45980 22170 -45946
rect 21326 -46034 21350 -46000
rect 21384 -46034 21408 -46000
rect 20564 -46088 20580 -46054
rect 21136 -46088 21152 -46054
rect 21326 -46058 21408 -46034
rect 22344 -46000 22426 -45976
rect 22600 -45980 22616 -45946
rect 23172 -45980 23188 -45946
rect 22344 -46034 22368 -46000
rect 22402 -46034 22426 -46000
rect 21582 -46088 21598 -46054
rect 22154 -46088 22170 -46054
rect 22344 -46058 22426 -46034
rect 23362 -46000 23444 -45976
rect 23618 -45980 23634 -45946
rect 24190 -45980 24206 -45946
rect 23362 -46034 23386 -46000
rect 23420 -46034 23444 -46000
rect 22600 -46088 22616 -46054
rect 23172 -46088 23188 -46054
rect 23362 -46058 23444 -46034
rect 24380 -46000 24462 -45976
rect 24636 -45980 24652 -45946
rect 25208 -45980 25224 -45946
rect 24380 -46034 24404 -46000
rect 24438 -46034 24462 -46000
rect 23618 -46088 23634 -46054
rect 24190 -46088 24206 -46054
rect 24380 -46058 24462 -46034
rect 25408 -46000 25490 -45976
rect 25408 -46034 25432 -46000
rect 25466 -46034 25490 -46000
rect 24636 -46088 24652 -46054
rect 25208 -46088 25224 -46054
rect 25408 -46058 25490 -46034
rect 16260 -46138 16294 -46122
rect 16260 -46730 16294 -46714
rect 17278 -46138 17312 -46122
rect 17278 -46730 17312 -46714
rect 18296 -46138 18330 -46122
rect 18296 -46730 18330 -46714
rect 19314 -46138 19348 -46122
rect 19314 -46730 19348 -46714
rect 20332 -46138 20366 -46122
rect 20332 -46730 20366 -46714
rect 21350 -46138 21384 -46122
rect 21350 -46730 21384 -46714
rect 22368 -46138 22402 -46122
rect 22368 -46730 22402 -46714
rect 23386 -46138 23420 -46122
rect 23386 -46730 23420 -46714
rect 24404 -46138 24438 -46122
rect 24404 -46730 24438 -46714
rect 25422 -46138 25456 -46122
rect 28258 -46172 28274 -46138
rect 28830 -46172 28846 -46138
rect 29276 -46172 29292 -46138
rect 29848 -46172 29864 -46138
rect 30294 -46172 30310 -46138
rect 30866 -46172 30882 -46138
rect 31312 -46172 31328 -46138
rect 31884 -46172 31900 -46138
rect 32330 -46172 32346 -46138
rect 32902 -46172 32918 -46138
rect 33348 -46172 33364 -46138
rect 33920 -46172 33936 -46138
rect 34366 -46172 34382 -46138
rect 34938 -46172 34954 -46138
rect 35384 -46172 35400 -46138
rect 35956 -46172 35972 -46138
rect 36402 -46172 36418 -46138
rect 36974 -46172 36990 -46138
rect 37420 -46172 37436 -46138
rect 37992 -46172 38008 -46138
rect 38438 -46172 38454 -46138
rect 39010 -46172 39026 -46138
rect 39456 -46172 39472 -46138
rect 40028 -46172 40044 -46138
rect 40474 -46172 40490 -46138
rect 41046 -46172 41062 -46138
rect 41492 -46172 41508 -46138
rect 42064 -46172 42080 -46138
rect 42510 -46172 42526 -46138
rect 43082 -46172 43098 -46138
rect 43528 -46172 43544 -46138
rect 44100 -46172 44116 -46138
rect 44546 -46172 44562 -46138
rect 45118 -46172 45134 -46138
rect 45564 -46172 45580 -46138
rect 46136 -46172 46152 -46138
rect 46582 -46172 46598 -46138
rect 47154 -46172 47170 -46138
rect 47600 -46172 47616 -46138
rect 48172 -46172 48188 -46138
rect 37682 -46178 37742 -46172
rect 25422 -46730 25456 -46714
rect 28026 -46222 28060 -46206
rect 17788 -46764 17848 -46762
rect 18802 -46764 18862 -46762
rect 22876 -46764 22936 -46762
rect 23892 -46764 23952 -46762
rect 16236 -46818 16318 -46794
rect 16492 -46798 16508 -46764
rect 17064 -46798 17080 -46764
rect 16236 -46852 16260 -46818
rect 16294 -46852 16318 -46818
rect 16236 -46876 16318 -46852
rect 17254 -46818 17336 -46794
rect 17510 -46798 17526 -46764
rect 18082 -46798 18098 -46764
rect 17254 -46852 17278 -46818
rect 17312 -46852 17336 -46818
rect 16492 -46906 16508 -46872
rect 17064 -46906 17080 -46872
rect 17254 -46876 17336 -46852
rect 18272 -46818 18354 -46794
rect 18528 -46798 18544 -46764
rect 19100 -46798 19116 -46764
rect 18272 -46852 18296 -46818
rect 18330 -46852 18354 -46818
rect 17510 -46906 17526 -46872
rect 18082 -46906 18098 -46872
rect 18272 -46876 18354 -46852
rect 19290 -46818 19372 -46794
rect 19546 -46798 19562 -46764
rect 20118 -46798 20134 -46764
rect 19290 -46852 19314 -46818
rect 19348 -46852 19372 -46818
rect 18528 -46906 18544 -46872
rect 19100 -46906 19116 -46872
rect 19290 -46876 19372 -46852
rect 20308 -46818 20390 -46794
rect 20564 -46798 20580 -46764
rect 21136 -46798 21152 -46764
rect 20308 -46852 20332 -46818
rect 20366 -46852 20390 -46818
rect 19546 -46906 19562 -46872
rect 20118 -46906 20134 -46872
rect 20308 -46876 20390 -46852
rect 21326 -46818 21408 -46794
rect 21582 -46798 21598 -46764
rect 22154 -46798 22170 -46764
rect 21326 -46852 21350 -46818
rect 21384 -46852 21408 -46818
rect 20564 -46906 20580 -46872
rect 21136 -46906 21152 -46872
rect 21326 -46876 21408 -46852
rect 22344 -46818 22426 -46794
rect 22600 -46798 22616 -46764
rect 23172 -46798 23188 -46764
rect 22344 -46852 22368 -46818
rect 22402 -46852 22426 -46818
rect 21582 -46906 21598 -46872
rect 22154 -46906 22170 -46872
rect 22344 -46876 22426 -46852
rect 23362 -46818 23444 -46794
rect 23618 -46798 23634 -46764
rect 24190 -46798 24206 -46764
rect 23362 -46852 23386 -46818
rect 23420 -46852 23444 -46818
rect 22600 -46906 22616 -46872
rect 23172 -46906 23188 -46872
rect 23362 -46876 23444 -46852
rect 24380 -46818 24462 -46794
rect 24636 -46798 24652 -46764
rect 25208 -46798 25224 -46764
rect 24380 -46852 24404 -46818
rect 24438 -46852 24462 -46818
rect 23618 -46906 23634 -46872
rect 24190 -46906 24206 -46872
rect 24380 -46876 24462 -46852
rect 25408 -46818 25490 -46794
rect 28026 -46814 28060 -46798
rect 29044 -46222 29078 -46206
rect 29044 -46814 29078 -46798
rect 30062 -46222 30096 -46206
rect 30062 -46814 30096 -46798
rect 31080 -46222 31114 -46206
rect 31080 -46814 31114 -46798
rect 32098 -46222 32132 -46206
rect 32098 -46814 32132 -46798
rect 33116 -46222 33150 -46206
rect 33116 -46814 33150 -46798
rect 34134 -46222 34168 -46206
rect 34134 -46814 34168 -46798
rect 35152 -46222 35186 -46206
rect 35152 -46814 35186 -46798
rect 36170 -46222 36204 -46206
rect 36170 -46814 36204 -46798
rect 37188 -46222 37222 -46206
rect 37188 -46814 37222 -46798
rect 38206 -46222 38240 -46206
rect 38206 -46814 38240 -46798
rect 39224 -46222 39258 -46206
rect 39224 -46814 39258 -46798
rect 40242 -46222 40276 -46206
rect 40242 -46814 40276 -46798
rect 41260 -46222 41294 -46206
rect 41260 -46814 41294 -46798
rect 42278 -46222 42312 -46206
rect 42278 -46814 42312 -46798
rect 43296 -46222 43330 -46206
rect 43296 -46814 43330 -46798
rect 44314 -46222 44348 -46206
rect 44314 -46814 44348 -46798
rect 45332 -46222 45366 -46206
rect 45332 -46814 45366 -46798
rect 46350 -46222 46384 -46206
rect 46350 -46814 46384 -46798
rect 47368 -46222 47402 -46206
rect 47368 -46814 47402 -46798
rect 48386 -46222 48420 -46206
rect 48386 -46814 48420 -46798
rect 25408 -46852 25432 -46818
rect 25466 -46852 25490 -46818
rect 33610 -46848 33670 -46842
rect 35646 -46848 35706 -46842
rect 36666 -46848 36726 -46842
rect 41738 -46848 41798 -46842
rect 24636 -46906 24652 -46872
rect 25208 -46906 25224 -46872
rect 25408 -46876 25490 -46852
rect 28258 -46882 28274 -46848
rect 28830 -46882 28846 -46848
rect 29276 -46882 29292 -46848
rect 29848 -46882 29864 -46848
rect 30294 -46882 30310 -46848
rect 30866 -46882 30882 -46848
rect 31312 -46882 31328 -46848
rect 31884 -46882 31900 -46848
rect 32330 -46882 32346 -46848
rect 32902 -46882 32918 -46848
rect 33348 -46882 33364 -46848
rect 33920 -46882 33936 -46848
rect 34366 -46882 34382 -46848
rect 34938 -46882 34954 -46848
rect 35384 -46882 35400 -46848
rect 35956 -46882 35972 -46848
rect 36402 -46882 36418 -46848
rect 36974 -46882 36990 -46848
rect 37420 -46882 37436 -46848
rect 37992 -46882 38008 -46848
rect 38438 -46882 38454 -46848
rect 39010 -46882 39026 -46848
rect 39456 -46882 39472 -46848
rect 40028 -46882 40044 -46848
rect 40474 -46882 40490 -46848
rect 41046 -46882 41062 -46848
rect 41492 -46882 41508 -46848
rect 42064 -46882 42080 -46848
rect 42510 -46882 42526 -46848
rect 43082 -46882 43098 -46848
rect 43528 -46882 43544 -46848
rect 44100 -46882 44116 -46848
rect 44546 -46882 44562 -46848
rect 45118 -46882 45134 -46848
rect 45564 -46882 45580 -46848
rect 46136 -46882 46152 -46848
rect 46582 -46882 46598 -46848
rect 47154 -46882 47170 -46848
rect 47600 -46882 47616 -46848
rect 48172 -46882 48188 -46848
rect 16260 -46956 16294 -46940
rect 16260 -47548 16294 -47532
rect 17278 -46956 17312 -46940
rect 17278 -47548 17312 -47532
rect 18296 -46956 18330 -46940
rect 18296 -47548 18330 -47532
rect 19314 -46956 19348 -46940
rect 19314 -47548 19348 -47532
rect 20332 -46956 20366 -46940
rect 20332 -47548 20366 -47532
rect 21350 -46956 21384 -46940
rect 21350 -47548 21384 -47532
rect 22368 -46956 22402 -46940
rect 22368 -47548 22402 -47532
rect 23386 -46956 23420 -46940
rect 23386 -47548 23420 -47532
rect 24404 -46956 24438 -46940
rect 24404 -47548 24438 -47532
rect 25422 -46956 25456 -46940
rect 28530 -47094 28612 -47070
rect 28530 -47128 28554 -47094
rect 28588 -47128 28612 -47094
rect 28530 -47152 28612 -47128
rect 29548 -47094 29630 -47070
rect 29548 -47128 29572 -47094
rect 29606 -47128 29630 -47094
rect 29548 -47152 29630 -47128
rect 30566 -47094 30648 -47070
rect 30566 -47128 30590 -47094
rect 30624 -47128 30648 -47094
rect 30566 -47152 30648 -47128
rect 31584 -47094 31666 -47070
rect 31584 -47128 31608 -47094
rect 31642 -47128 31666 -47094
rect 31584 -47152 31666 -47128
rect 32602 -47094 32684 -47070
rect 32602 -47128 32626 -47094
rect 32660 -47128 32684 -47094
rect 32602 -47152 32684 -47128
rect 33620 -47094 33702 -47070
rect 33620 -47128 33644 -47094
rect 33678 -47128 33702 -47094
rect 33620 -47152 33702 -47128
rect 34638 -47094 34720 -47070
rect 34638 -47128 34662 -47094
rect 34696 -47128 34720 -47094
rect 34638 -47152 34720 -47128
rect 35656 -47094 35738 -47070
rect 35656 -47128 35680 -47094
rect 35714 -47128 35738 -47094
rect 35656 -47152 35738 -47128
rect 36674 -47094 36756 -47070
rect 36674 -47128 36698 -47094
rect 36732 -47128 36756 -47094
rect 36674 -47152 36756 -47128
rect 37692 -47094 37774 -47070
rect 37692 -47128 37716 -47094
rect 37750 -47128 37774 -47094
rect 37692 -47152 37774 -47128
rect 38710 -47094 38792 -47070
rect 38710 -47128 38734 -47094
rect 38768 -47128 38792 -47094
rect 38710 -47152 38792 -47128
rect 39728 -47094 39810 -47070
rect 39728 -47128 39752 -47094
rect 39786 -47128 39810 -47094
rect 39728 -47152 39810 -47128
rect 40746 -47094 40828 -47070
rect 40746 -47128 40770 -47094
rect 40804 -47128 40828 -47094
rect 40746 -47152 40828 -47128
rect 41764 -47094 41846 -47070
rect 41764 -47128 41788 -47094
rect 41822 -47128 41846 -47094
rect 41764 -47152 41846 -47128
rect 42782 -47094 42864 -47070
rect 42782 -47128 42806 -47094
rect 42840 -47128 42864 -47094
rect 42782 -47152 42864 -47128
rect 43800 -47094 43882 -47070
rect 43800 -47128 43824 -47094
rect 43858 -47128 43882 -47094
rect 43800 -47152 43882 -47128
rect 44818 -47094 44900 -47070
rect 44818 -47128 44842 -47094
rect 44876 -47128 44900 -47094
rect 44818 -47152 44900 -47128
rect 45836 -47094 45918 -47070
rect 45836 -47128 45860 -47094
rect 45894 -47128 45918 -47094
rect 45836 -47152 45918 -47128
rect 46854 -47094 46936 -47070
rect 46854 -47128 46878 -47094
rect 46912 -47128 46936 -47094
rect 46854 -47152 46936 -47128
rect 47872 -47094 47954 -47070
rect 47872 -47128 47896 -47094
rect 47930 -47128 47954 -47094
rect 47872 -47152 47954 -47128
rect 28258 -47404 28274 -47370
rect 28830 -47404 28846 -47370
rect 29276 -47404 29292 -47370
rect 29848 -47404 29864 -47370
rect 30294 -47404 30310 -47370
rect 30866 -47404 30882 -47370
rect 31312 -47404 31328 -47370
rect 31884 -47404 31900 -47370
rect 32330 -47404 32346 -47370
rect 32902 -47404 32918 -47370
rect 33348 -47404 33364 -47370
rect 33920 -47404 33936 -47370
rect 34366 -47404 34382 -47370
rect 34938 -47404 34954 -47370
rect 35384 -47404 35400 -47370
rect 35956 -47404 35972 -47370
rect 36402 -47404 36418 -47370
rect 36974 -47404 36990 -47370
rect 37420 -47404 37436 -47370
rect 37992 -47404 38008 -47370
rect 38438 -47404 38454 -47370
rect 39010 -47404 39026 -47370
rect 39456 -47404 39472 -47370
rect 40028 -47404 40044 -47370
rect 40474 -47404 40490 -47370
rect 41046 -47404 41062 -47370
rect 41492 -47404 41508 -47370
rect 42064 -47404 42080 -47370
rect 42510 -47404 42526 -47370
rect 43082 -47404 43098 -47370
rect 43528 -47404 43544 -47370
rect 44100 -47404 44116 -47370
rect 44546 -47404 44562 -47370
rect 45118 -47404 45134 -47370
rect 45564 -47404 45580 -47370
rect 46136 -47404 46152 -47370
rect 46582 -47404 46598 -47370
rect 47154 -47404 47170 -47370
rect 47600 -47404 47616 -47370
rect 48172 -47404 48188 -47370
rect 29544 -47408 29604 -47404
rect 30560 -47408 30620 -47404
rect 34636 -47412 34696 -47404
rect 38702 -47408 38762 -47404
rect 40736 -47408 40796 -47404
rect 46848 -47408 46908 -47404
rect 25422 -47548 25456 -47532
rect 28026 -47454 28060 -47438
rect 16236 -47636 16318 -47612
rect 16492 -47616 16508 -47582
rect 17064 -47616 17080 -47582
rect 16236 -47670 16260 -47636
rect 16294 -47670 16318 -47636
rect 16236 -47694 16318 -47670
rect 17254 -47636 17336 -47612
rect 17510 -47616 17526 -47582
rect 18082 -47616 18098 -47582
rect 17254 -47670 17278 -47636
rect 17312 -47670 17336 -47636
rect 16492 -47724 16508 -47690
rect 17064 -47724 17080 -47690
rect 17254 -47694 17336 -47670
rect 18272 -47636 18354 -47612
rect 18528 -47616 18544 -47582
rect 19100 -47616 19116 -47582
rect 18272 -47670 18296 -47636
rect 18330 -47670 18354 -47636
rect 17510 -47724 17526 -47690
rect 18082 -47724 18098 -47690
rect 18272 -47694 18354 -47670
rect 19290 -47636 19372 -47612
rect 19546 -47616 19562 -47582
rect 20118 -47616 20134 -47582
rect 19290 -47670 19314 -47636
rect 19348 -47670 19372 -47636
rect 18528 -47724 18544 -47690
rect 19100 -47724 19116 -47690
rect 19290 -47694 19372 -47670
rect 20308 -47636 20390 -47612
rect 20564 -47616 20580 -47582
rect 21136 -47616 21152 -47582
rect 20308 -47670 20332 -47636
rect 20366 -47670 20390 -47636
rect 19546 -47724 19562 -47690
rect 20118 -47724 20134 -47690
rect 20308 -47694 20390 -47670
rect 21326 -47636 21408 -47612
rect 21582 -47616 21598 -47582
rect 22154 -47616 22170 -47582
rect 21326 -47670 21350 -47636
rect 21384 -47670 21408 -47636
rect 20564 -47724 20580 -47690
rect 21136 -47724 21152 -47690
rect 21326 -47694 21408 -47670
rect 22344 -47636 22426 -47612
rect 22600 -47616 22616 -47582
rect 23172 -47616 23188 -47582
rect 22344 -47670 22368 -47636
rect 22402 -47670 22426 -47636
rect 21582 -47724 21598 -47690
rect 22154 -47724 22170 -47690
rect 22344 -47694 22426 -47670
rect 23362 -47636 23444 -47612
rect 23618 -47616 23634 -47582
rect 24190 -47616 24206 -47582
rect 23362 -47670 23386 -47636
rect 23420 -47670 23444 -47636
rect 22600 -47724 22616 -47690
rect 23172 -47724 23188 -47690
rect 23362 -47694 23444 -47670
rect 24380 -47636 24462 -47612
rect 24636 -47616 24652 -47582
rect 25208 -47616 25224 -47582
rect 24380 -47670 24404 -47636
rect 24438 -47670 24462 -47636
rect 23618 -47724 23634 -47690
rect 24190 -47724 24206 -47690
rect 24380 -47694 24462 -47670
rect 25408 -47636 25490 -47612
rect 25408 -47670 25432 -47636
rect 25466 -47670 25490 -47636
rect 24636 -47724 24652 -47690
rect 25208 -47724 25224 -47690
rect 25408 -47694 25490 -47670
rect 21848 -47726 21908 -47724
rect 16260 -47774 16294 -47758
rect 16260 -48366 16294 -48350
rect 17278 -47774 17312 -47758
rect 17278 -48366 17312 -48350
rect 18296 -47774 18330 -47758
rect 18296 -48366 18330 -48350
rect 19314 -47774 19348 -47758
rect 19314 -48366 19348 -48350
rect 20332 -47774 20366 -47758
rect 20332 -48366 20366 -48350
rect 21350 -47774 21384 -47758
rect 21350 -48366 21384 -48350
rect 22368 -47774 22402 -47758
rect 22368 -48366 22402 -48350
rect 23386 -47774 23420 -47758
rect 23386 -48366 23420 -48350
rect 24404 -47774 24438 -47758
rect 24404 -48366 24438 -48350
rect 25422 -47774 25456 -47758
rect 28026 -48046 28060 -48030
rect 29044 -47454 29078 -47438
rect 29044 -48046 29078 -48030
rect 30062 -47454 30096 -47438
rect 30062 -48046 30096 -48030
rect 31080 -47454 31114 -47438
rect 31080 -48046 31114 -48030
rect 32098 -47454 32132 -47438
rect 32098 -48046 32132 -48030
rect 33116 -47454 33150 -47438
rect 33116 -48046 33150 -48030
rect 34134 -47454 34168 -47438
rect 34134 -48046 34168 -48030
rect 35152 -47454 35186 -47438
rect 35152 -48046 35186 -48030
rect 36170 -47454 36204 -47438
rect 36170 -48046 36204 -48030
rect 37188 -47454 37222 -47438
rect 37188 -48046 37222 -48030
rect 38206 -47454 38240 -47438
rect 38206 -48046 38240 -48030
rect 39224 -47454 39258 -47438
rect 39224 -48046 39258 -48030
rect 40242 -47454 40276 -47438
rect 40242 -48046 40276 -48030
rect 41260 -47454 41294 -47438
rect 41260 -48046 41294 -48030
rect 42278 -47454 42312 -47438
rect 42278 -48046 42312 -48030
rect 43296 -47454 43330 -47438
rect 43296 -48046 43330 -48030
rect 44314 -47454 44348 -47438
rect 44314 -48046 44348 -48030
rect 45332 -47454 45366 -47438
rect 45332 -48046 45366 -48030
rect 46350 -47454 46384 -47438
rect 46350 -48046 46384 -48030
rect 47368 -47454 47402 -47438
rect 47368 -48046 47402 -48030
rect 48386 -47454 48420 -47438
rect 48420 -48030 48426 -47982
rect 48386 -48046 48420 -48030
rect 31570 -48080 31630 -48078
rect 28258 -48114 28274 -48080
rect 28830 -48114 28846 -48080
rect 29276 -48114 29292 -48080
rect 29848 -48114 29864 -48080
rect 30294 -48114 30310 -48080
rect 30866 -48114 30882 -48080
rect 31312 -48114 31328 -48080
rect 31884 -48114 31900 -48080
rect 32330 -48114 32346 -48080
rect 32902 -48114 32918 -48080
rect 33348 -48114 33364 -48080
rect 33920 -48114 33936 -48080
rect 34366 -48114 34382 -48080
rect 34938 -48114 34954 -48080
rect 35384 -48114 35400 -48080
rect 35956 -48114 35972 -48080
rect 36402 -48114 36418 -48080
rect 36974 -48114 36990 -48080
rect 37420 -48114 37436 -48080
rect 37992 -48114 38008 -48080
rect 38438 -48114 38454 -48080
rect 39010 -48114 39026 -48080
rect 39456 -48114 39472 -48080
rect 40028 -48114 40044 -48080
rect 40474 -48114 40490 -48080
rect 41046 -48114 41062 -48080
rect 41492 -48114 41508 -48080
rect 42064 -48114 42080 -48080
rect 42510 -48114 42526 -48080
rect 43082 -48114 43098 -48080
rect 43528 -48114 43544 -48080
rect 44100 -48114 44116 -48080
rect 44546 -48114 44562 -48080
rect 45118 -48114 45134 -48080
rect 45564 -48114 45580 -48080
rect 46136 -48114 46152 -48080
rect 46582 -48114 46598 -48080
rect 47154 -48114 47170 -48080
rect 47600 -48114 47616 -48080
rect 48172 -48114 48188 -48080
rect 33604 -48118 33664 -48114
rect 42762 -48128 42822 -48114
rect 43796 -48128 43856 -48114
rect 25422 -48366 25456 -48350
rect 28518 -48330 28600 -48306
rect 28518 -48364 28542 -48330
rect 28576 -48364 28600 -48330
rect 28518 -48388 28600 -48364
rect 29536 -48330 29618 -48306
rect 29536 -48364 29560 -48330
rect 29594 -48364 29618 -48330
rect 29536 -48388 29618 -48364
rect 30554 -48330 30636 -48306
rect 30554 -48364 30578 -48330
rect 30612 -48364 30636 -48330
rect 30554 -48388 30636 -48364
rect 31572 -48330 31654 -48306
rect 31572 -48364 31596 -48330
rect 31630 -48364 31654 -48330
rect 31572 -48388 31654 -48364
rect 32590 -48330 32672 -48306
rect 32590 -48364 32614 -48330
rect 32648 -48364 32672 -48330
rect 32590 -48388 32672 -48364
rect 33608 -48330 33690 -48306
rect 33608 -48364 33632 -48330
rect 33666 -48364 33690 -48330
rect 33608 -48388 33690 -48364
rect 34626 -48330 34708 -48306
rect 34626 -48364 34650 -48330
rect 34684 -48364 34708 -48330
rect 34626 -48388 34708 -48364
rect 35644 -48330 35726 -48306
rect 35644 -48364 35668 -48330
rect 35702 -48364 35726 -48330
rect 35644 -48388 35726 -48364
rect 36662 -48330 36744 -48306
rect 36662 -48364 36686 -48330
rect 36720 -48364 36744 -48330
rect 36662 -48388 36744 -48364
rect 37680 -48330 37762 -48306
rect 37680 -48364 37704 -48330
rect 37738 -48364 37762 -48330
rect 37680 -48388 37762 -48364
rect 38698 -48330 38780 -48306
rect 38698 -48364 38722 -48330
rect 38756 -48364 38780 -48330
rect 38698 -48388 38780 -48364
rect 39716 -48330 39798 -48306
rect 39716 -48364 39740 -48330
rect 39774 -48364 39798 -48330
rect 39716 -48388 39798 -48364
rect 40734 -48330 40816 -48306
rect 40734 -48364 40758 -48330
rect 40792 -48364 40816 -48330
rect 40734 -48388 40816 -48364
rect 41752 -48330 41834 -48306
rect 41752 -48364 41776 -48330
rect 41810 -48364 41834 -48330
rect 41752 -48388 41834 -48364
rect 42770 -48330 42852 -48306
rect 42770 -48364 42794 -48330
rect 42828 -48364 42852 -48330
rect 42770 -48388 42852 -48364
rect 43788 -48330 43870 -48306
rect 43788 -48364 43812 -48330
rect 43846 -48364 43870 -48330
rect 43788 -48388 43870 -48364
rect 44806 -48330 44888 -48306
rect 44806 -48364 44830 -48330
rect 44864 -48364 44888 -48330
rect 44806 -48388 44888 -48364
rect 45824 -48330 45906 -48306
rect 45824 -48364 45848 -48330
rect 45882 -48364 45906 -48330
rect 45824 -48388 45906 -48364
rect 46842 -48330 46924 -48306
rect 46842 -48364 46866 -48330
rect 46900 -48364 46924 -48330
rect 46842 -48388 46924 -48364
rect 47860 -48330 47942 -48306
rect 47860 -48364 47884 -48330
rect 47918 -48364 47942 -48330
rect 47860 -48388 47942 -48364
rect 17774 -48400 17834 -48398
rect 18788 -48400 18848 -48398
rect 22862 -48400 22922 -48398
rect 23878 -48400 23938 -48398
rect 16236 -48454 16318 -48430
rect 16492 -48434 16508 -48400
rect 17064 -48434 17080 -48400
rect 16236 -48488 16260 -48454
rect 16294 -48488 16318 -48454
rect 16236 -48512 16318 -48488
rect 17254 -48454 17336 -48430
rect 17510 -48434 17526 -48400
rect 18082 -48434 18098 -48400
rect 17254 -48488 17278 -48454
rect 17312 -48488 17336 -48454
rect 16492 -48542 16508 -48508
rect 17064 -48542 17080 -48508
rect 17254 -48512 17336 -48488
rect 18272 -48454 18354 -48430
rect 18528 -48434 18544 -48400
rect 19100 -48434 19116 -48400
rect 18272 -48488 18296 -48454
rect 18330 -48488 18354 -48454
rect 17510 -48542 17526 -48508
rect 18082 -48542 18098 -48508
rect 18272 -48512 18354 -48488
rect 19290 -48454 19372 -48430
rect 19546 -48434 19562 -48400
rect 20118 -48434 20134 -48400
rect 19290 -48488 19314 -48454
rect 19348 -48488 19372 -48454
rect 18528 -48542 18544 -48508
rect 19100 -48542 19116 -48508
rect 19290 -48512 19372 -48488
rect 20308 -48454 20390 -48430
rect 20564 -48434 20580 -48400
rect 21136 -48434 21152 -48400
rect 20308 -48488 20332 -48454
rect 20366 -48488 20390 -48454
rect 19546 -48542 19562 -48508
rect 20118 -48542 20134 -48508
rect 20308 -48512 20390 -48488
rect 21326 -48454 21408 -48430
rect 21582 -48434 21598 -48400
rect 22154 -48434 22170 -48400
rect 21326 -48488 21350 -48454
rect 21384 -48488 21408 -48454
rect 20564 -48542 20580 -48508
rect 21136 -48542 21152 -48508
rect 21326 -48512 21408 -48488
rect 22344 -48454 22426 -48430
rect 22600 -48434 22616 -48400
rect 23172 -48434 23188 -48400
rect 22344 -48488 22368 -48454
rect 22402 -48488 22426 -48454
rect 21582 -48542 21598 -48508
rect 22154 -48542 22170 -48508
rect 22344 -48512 22426 -48488
rect 23362 -48454 23444 -48430
rect 23618 -48434 23634 -48400
rect 24190 -48434 24206 -48400
rect 23362 -48488 23386 -48454
rect 23420 -48488 23444 -48454
rect 22600 -48542 22616 -48508
rect 23172 -48542 23188 -48508
rect 23362 -48512 23444 -48488
rect 24380 -48454 24462 -48430
rect 24636 -48434 24652 -48400
rect 25208 -48434 25224 -48400
rect 24380 -48488 24404 -48454
rect 24438 -48488 24462 -48454
rect 23618 -48542 23634 -48508
rect 24190 -48542 24206 -48508
rect 24380 -48512 24462 -48488
rect 25408 -48454 25490 -48430
rect 25408 -48488 25432 -48454
rect 25466 -48488 25490 -48454
rect 24636 -48542 24652 -48508
rect 25208 -48542 25224 -48508
rect 25408 -48512 25490 -48488
rect 16260 -48592 16294 -48576
rect 16260 -49184 16294 -49168
rect 17278 -48592 17312 -48576
rect 17278 -49184 17312 -49168
rect 18296 -48592 18330 -48576
rect 18296 -49184 18330 -49168
rect 19314 -48592 19348 -48576
rect 19314 -49184 19348 -49168
rect 20332 -48592 20366 -48576
rect 20332 -49184 20366 -49168
rect 21350 -48592 21384 -48576
rect 21350 -49184 21384 -49168
rect 22368 -48592 22402 -48576
rect 22368 -49184 22402 -49168
rect 23386 -48592 23420 -48576
rect 23386 -49184 23420 -49168
rect 24404 -48592 24438 -48576
rect 24404 -49184 24438 -49168
rect 25422 -48592 25456 -48576
rect 28256 -48638 28272 -48604
rect 28828 -48638 28844 -48604
rect 29274 -48638 29290 -48604
rect 29846 -48638 29862 -48604
rect 30292 -48638 30308 -48604
rect 30864 -48638 30880 -48604
rect 31310 -48638 31326 -48604
rect 31882 -48638 31898 -48604
rect 32328 -48638 32344 -48604
rect 32900 -48638 32916 -48604
rect 33346 -48638 33362 -48604
rect 33918 -48638 33934 -48604
rect 34364 -48638 34380 -48604
rect 34936 -48638 34952 -48604
rect 35382 -48638 35398 -48604
rect 35954 -48638 35970 -48604
rect 36400 -48638 36416 -48604
rect 36972 -48638 36988 -48604
rect 37418 -48638 37434 -48604
rect 37990 -48638 38006 -48604
rect 38436 -48638 38452 -48604
rect 39008 -48638 39024 -48604
rect 39454 -48638 39470 -48604
rect 40026 -48638 40042 -48604
rect 40472 -48638 40488 -48604
rect 41044 -48638 41060 -48604
rect 41490 -48638 41506 -48604
rect 42062 -48638 42078 -48604
rect 42508 -48638 42524 -48604
rect 43080 -48638 43096 -48604
rect 43526 -48638 43542 -48604
rect 44098 -48638 44114 -48604
rect 44544 -48638 44560 -48604
rect 45116 -48638 45132 -48604
rect 45562 -48638 45578 -48604
rect 46134 -48638 46150 -48604
rect 46580 -48638 46596 -48604
rect 47152 -48638 47168 -48604
rect 47598 -48638 47614 -48604
rect 48170 -48638 48186 -48604
rect 30566 -48642 30626 -48638
rect 25422 -49184 25456 -49168
rect 28024 -48688 28058 -48672
rect 17778 -49218 17838 -49216
rect 18792 -49218 18852 -49216
rect 22866 -49218 22926 -49216
rect 23882 -49218 23942 -49216
rect 16236 -49272 16318 -49248
rect 16492 -49252 16508 -49218
rect 17064 -49252 17080 -49218
rect 16236 -49306 16260 -49272
rect 16294 -49306 16318 -49272
rect 16236 -49330 16318 -49306
rect 17254 -49272 17336 -49248
rect 17510 -49252 17526 -49218
rect 18082 -49252 18098 -49218
rect 17254 -49306 17278 -49272
rect 17312 -49306 17336 -49272
rect 16492 -49360 16508 -49326
rect 17064 -49360 17080 -49326
rect 17254 -49330 17336 -49306
rect 18272 -49272 18354 -49248
rect 18528 -49252 18544 -49218
rect 19100 -49252 19116 -49218
rect 18272 -49306 18296 -49272
rect 18330 -49306 18354 -49272
rect 17510 -49360 17526 -49326
rect 18082 -49360 18098 -49326
rect 18272 -49330 18354 -49306
rect 19290 -49272 19372 -49248
rect 19546 -49252 19562 -49218
rect 20118 -49252 20134 -49218
rect 19290 -49306 19314 -49272
rect 19348 -49306 19372 -49272
rect 18528 -49360 18544 -49326
rect 19100 -49360 19116 -49326
rect 19290 -49330 19372 -49306
rect 20308 -49272 20390 -49248
rect 20564 -49252 20580 -49218
rect 21136 -49252 21152 -49218
rect 20308 -49306 20332 -49272
rect 20366 -49306 20390 -49272
rect 19546 -49360 19562 -49326
rect 20118 -49360 20134 -49326
rect 20308 -49330 20390 -49306
rect 21326 -49272 21408 -49248
rect 21582 -49252 21598 -49218
rect 22154 -49252 22170 -49218
rect 21326 -49306 21350 -49272
rect 21384 -49306 21408 -49272
rect 20564 -49360 20580 -49326
rect 21136 -49360 21152 -49326
rect 21326 -49330 21408 -49306
rect 22344 -49272 22426 -49248
rect 22600 -49252 22616 -49218
rect 23172 -49252 23188 -49218
rect 22344 -49306 22368 -49272
rect 22402 -49306 22426 -49272
rect 21582 -49360 21598 -49326
rect 22154 -49360 22170 -49326
rect 22344 -49330 22426 -49306
rect 23362 -49272 23444 -49248
rect 23618 -49252 23634 -49218
rect 24190 -49252 24206 -49218
rect 23362 -49306 23386 -49272
rect 23420 -49306 23444 -49272
rect 22600 -49360 22616 -49326
rect 23172 -49360 23188 -49326
rect 23362 -49330 23444 -49306
rect 24380 -49272 24462 -49248
rect 24636 -49252 24652 -49218
rect 25208 -49252 25224 -49218
rect 24380 -49306 24404 -49272
rect 24438 -49306 24462 -49272
rect 23618 -49360 23634 -49326
rect 24190 -49360 24206 -49326
rect 24380 -49330 24462 -49306
rect 25408 -49272 25490 -49248
rect 25408 -49306 25432 -49272
rect 25466 -49306 25490 -49272
rect 28024 -49280 28058 -49264
rect 29042 -48688 29076 -48672
rect 29042 -49280 29076 -49264
rect 30060 -48688 30094 -48672
rect 30060 -49280 30094 -49264
rect 31078 -48688 31112 -48672
rect 31078 -49280 31112 -49264
rect 32096 -48688 32130 -48672
rect 32096 -49280 32130 -49264
rect 33114 -48688 33148 -48672
rect 33114 -49280 33148 -49264
rect 34132 -48688 34166 -48672
rect 34132 -49280 34166 -49264
rect 35150 -48688 35184 -48672
rect 35150 -49280 35184 -49264
rect 36168 -48688 36202 -48672
rect 36168 -49280 36202 -49264
rect 37186 -48688 37220 -48672
rect 37186 -49280 37220 -49264
rect 38204 -48688 38238 -48672
rect 38204 -49280 38238 -49264
rect 39222 -48688 39256 -48672
rect 39222 -49280 39256 -49264
rect 40240 -48688 40274 -48672
rect 40240 -49280 40274 -49264
rect 41258 -48688 41292 -48672
rect 41258 -49280 41292 -49264
rect 42276 -48688 42310 -48672
rect 42276 -49280 42310 -49264
rect 43294 -48688 43328 -48672
rect 43294 -49280 43328 -49264
rect 44312 -48688 44346 -48672
rect 44312 -49280 44346 -49264
rect 45330 -48688 45364 -48672
rect 45330 -49280 45364 -49264
rect 46348 -48688 46382 -48672
rect 46348 -49280 46382 -49264
rect 47366 -48688 47400 -48672
rect 47366 -49280 47400 -49264
rect 48384 -48688 48418 -48672
rect 48384 -49280 48418 -49264
rect 24636 -49360 24652 -49326
rect 25208 -49360 25224 -49326
rect 25408 -49330 25490 -49306
rect 35634 -49314 35694 -49310
rect 36662 -49314 36722 -49312
rect 38706 -49314 38766 -49310
rect 28256 -49348 28272 -49314
rect 28828 -49348 28844 -49314
rect 29274 -49348 29290 -49314
rect 29846 -49348 29862 -49314
rect 30292 -49348 30308 -49314
rect 30864 -49348 30880 -49314
rect 31310 -49348 31326 -49314
rect 31882 -49348 31898 -49314
rect 32328 -49348 32344 -49314
rect 32900 -49348 32916 -49314
rect 33346 -49348 33362 -49314
rect 33918 -49348 33934 -49314
rect 34364 -49348 34380 -49314
rect 34936 -49348 34952 -49314
rect 35382 -49348 35398 -49314
rect 35954 -49348 35970 -49314
rect 36400 -49348 36416 -49314
rect 36972 -49348 36988 -49314
rect 37418 -49348 37434 -49314
rect 37990 -49348 38006 -49314
rect 38436 -49348 38452 -49314
rect 39008 -49348 39024 -49314
rect 39454 -49348 39470 -49314
rect 40026 -49348 40042 -49314
rect 40472 -49348 40488 -49314
rect 41044 -49348 41060 -49314
rect 41490 -49348 41506 -49314
rect 42062 -49348 42078 -49314
rect 42508 -49348 42524 -49314
rect 43080 -49348 43096 -49314
rect 43526 -49348 43542 -49314
rect 44098 -49348 44114 -49314
rect 44544 -49348 44560 -49314
rect 45116 -49348 45132 -49314
rect 45562 -49348 45578 -49314
rect 46134 -49348 46150 -49314
rect 46580 -49348 46596 -49314
rect 47152 -49348 47168 -49314
rect 47598 -49348 47614 -49314
rect 48170 -49348 48186 -49314
rect 16260 -49410 16294 -49394
rect 16260 -50002 16294 -49986
rect 17278 -49410 17312 -49394
rect 17278 -50002 17312 -49986
rect 18296 -49410 18330 -49394
rect 18296 -50002 18330 -49986
rect 19314 -49410 19348 -49394
rect 19314 -50002 19348 -49986
rect 20332 -49410 20366 -49394
rect 20332 -50002 20366 -49986
rect 21350 -49410 21384 -49394
rect 21350 -50002 21384 -49986
rect 22368 -49410 22402 -49394
rect 22368 -50002 22402 -49986
rect 23386 -49410 23420 -49394
rect 23386 -50002 23420 -49986
rect 24404 -49410 24438 -49394
rect 24404 -50002 24438 -49986
rect 25422 -49410 25456 -49394
rect 28518 -49554 28600 -49530
rect 28518 -49588 28542 -49554
rect 28576 -49588 28600 -49554
rect 28518 -49612 28600 -49588
rect 29536 -49554 29618 -49530
rect 29536 -49588 29560 -49554
rect 29594 -49588 29618 -49554
rect 29536 -49612 29618 -49588
rect 30554 -49554 30636 -49530
rect 30554 -49588 30578 -49554
rect 30612 -49588 30636 -49554
rect 30554 -49612 30636 -49588
rect 31572 -49554 31654 -49530
rect 31572 -49588 31596 -49554
rect 31630 -49588 31654 -49554
rect 31572 -49612 31654 -49588
rect 32590 -49554 32672 -49530
rect 32590 -49588 32614 -49554
rect 32648 -49588 32672 -49554
rect 32590 -49612 32672 -49588
rect 33608 -49554 33690 -49530
rect 33608 -49588 33632 -49554
rect 33666 -49588 33690 -49554
rect 33608 -49612 33690 -49588
rect 34626 -49554 34708 -49530
rect 34626 -49588 34650 -49554
rect 34684 -49588 34708 -49554
rect 34626 -49612 34708 -49588
rect 35644 -49554 35726 -49530
rect 35644 -49588 35668 -49554
rect 35702 -49588 35726 -49554
rect 35644 -49612 35726 -49588
rect 36662 -49554 36744 -49530
rect 36662 -49588 36686 -49554
rect 36720 -49588 36744 -49554
rect 36662 -49612 36744 -49588
rect 37680 -49554 37762 -49530
rect 37680 -49588 37704 -49554
rect 37738 -49588 37762 -49554
rect 37680 -49612 37762 -49588
rect 38698 -49554 38780 -49530
rect 38698 -49588 38722 -49554
rect 38756 -49588 38780 -49554
rect 38698 -49612 38780 -49588
rect 39716 -49554 39798 -49530
rect 39716 -49588 39740 -49554
rect 39774 -49588 39798 -49554
rect 39716 -49612 39798 -49588
rect 40734 -49554 40816 -49530
rect 40734 -49588 40758 -49554
rect 40792 -49588 40816 -49554
rect 40734 -49612 40816 -49588
rect 41752 -49554 41834 -49530
rect 41752 -49588 41776 -49554
rect 41810 -49588 41834 -49554
rect 41752 -49612 41834 -49588
rect 42770 -49554 42852 -49530
rect 42770 -49588 42794 -49554
rect 42828 -49588 42852 -49554
rect 42770 -49612 42852 -49588
rect 43788 -49554 43870 -49530
rect 43788 -49588 43812 -49554
rect 43846 -49588 43870 -49554
rect 43788 -49612 43870 -49588
rect 44806 -49554 44888 -49530
rect 44806 -49588 44830 -49554
rect 44864 -49588 44888 -49554
rect 44806 -49612 44888 -49588
rect 45824 -49554 45906 -49530
rect 45824 -49588 45848 -49554
rect 45882 -49588 45906 -49554
rect 45824 -49612 45906 -49588
rect 46842 -49554 46924 -49530
rect 46842 -49588 46866 -49554
rect 46900 -49588 46924 -49554
rect 46842 -49612 46924 -49588
rect 47860 -49554 47942 -49530
rect 47860 -49588 47884 -49554
rect 47918 -49588 47942 -49554
rect 47860 -49612 47942 -49588
rect 28256 -49872 28272 -49838
rect 28828 -49872 28844 -49838
rect 29274 -49872 29290 -49838
rect 29846 -49872 29862 -49838
rect 30292 -49872 30308 -49838
rect 30864 -49872 30880 -49838
rect 31310 -49872 31326 -49838
rect 31882 -49872 31898 -49838
rect 32328 -49872 32344 -49838
rect 32900 -49872 32916 -49838
rect 33346 -49872 33362 -49838
rect 33918 -49872 33934 -49838
rect 34364 -49872 34380 -49838
rect 34936 -49872 34952 -49838
rect 35382 -49872 35398 -49838
rect 35954 -49872 35970 -49838
rect 36400 -49872 36416 -49838
rect 36972 -49872 36988 -49838
rect 37418 -49872 37434 -49838
rect 37990 -49872 38006 -49838
rect 38436 -49872 38452 -49838
rect 39008 -49872 39024 -49838
rect 39454 -49872 39470 -49838
rect 40026 -49872 40042 -49838
rect 40472 -49872 40488 -49838
rect 41044 -49872 41060 -49838
rect 41490 -49872 41506 -49838
rect 42062 -49872 42078 -49838
rect 42508 -49872 42524 -49838
rect 43080 -49872 43096 -49838
rect 43526 -49872 43542 -49838
rect 44098 -49872 44114 -49838
rect 44544 -49872 44560 -49838
rect 45116 -49872 45132 -49838
rect 45562 -49872 45578 -49838
rect 46134 -49872 46150 -49838
rect 46580 -49872 46596 -49838
rect 47152 -49872 47168 -49838
rect 47598 -49872 47614 -49838
rect 48170 -49872 48186 -49838
rect 25422 -50002 25456 -49986
rect 28024 -49922 28058 -49906
rect 16752 -50036 16812 -50034
rect 17778 -50036 17838 -50032
rect 18792 -50036 18852 -50032
rect 19812 -50036 19872 -50034
rect 20834 -50036 20894 -50034
rect 22866 -50036 22926 -50032
rect 23882 -50036 23942 -50032
rect 24902 -50036 24962 -50034
rect 16236 -50090 16318 -50066
rect 16492 -50070 16508 -50036
rect 17064 -50070 17080 -50036
rect 16236 -50124 16260 -50090
rect 16294 -50124 16318 -50090
rect 16236 -50148 16318 -50124
rect 17254 -50090 17336 -50066
rect 17510 -50070 17526 -50036
rect 18082 -50070 18098 -50036
rect 17254 -50124 17278 -50090
rect 17312 -50124 17336 -50090
rect 16492 -50178 16508 -50144
rect 17064 -50178 17080 -50144
rect 17254 -50148 17336 -50124
rect 18272 -50090 18354 -50066
rect 18528 -50070 18544 -50036
rect 19100 -50070 19116 -50036
rect 18272 -50124 18296 -50090
rect 18330 -50124 18354 -50090
rect 17510 -50178 17526 -50144
rect 18082 -50178 18098 -50144
rect 18272 -50148 18354 -50124
rect 19290 -50090 19372 -50066
rect 19546 -50070 19562 -50036
rect 20118 -50070 20134 -50036
rect 19290 -50124 19314 -50090
rect 19348 -50124 19372 -50090
rect 18528 -50178 18544 -50144
rect 19100 -50178 19116 -50144
rect 19290 -50148 19372 -50124
rect 20308 -50090 20390 -50066
rect 20564 -50070 20580 -50036
rect 21136 -50070 21152 -50036
rect 20308 -50124 20332 -50090
rect 20366 -50124 20390 -50090
rect 19546 -50178 19562 -50144
rect 20118 -50178 20134 -50144
rect 20308 -50148 20390 -50124
rect 21326 -50090 21408 -50066
rect 21582 -50070 21598 -50036
rect 22154 -50070 22170 -50036
rect 21326 -50124 21350 -50090
rect 21384 -50124 21408 -50090
rect 20564 -50178 20580 -50144
rect 21136 -50178 21152 -50144
rect 21326 -50148 21408 -50124
rect 22344 -50090 22426 -50066
rect 22600 -50070 22616 -50036
rect 23172 -50070 23188 -50036
rect 22344 -50124 22368 -50090
rect 22402 -50124 22426 -50090
rect 21582 -50178 21598 -50144
rect 22154 -50178 22170 -50144
rect 22344 -50148 22426 -50124
rect 23362 -50090 23444 -50066
rect 23618 -50070 23634 -50036
rect 24190 -50070 24206 -50036
rect 23362 -50124 23386 -50090
rect 23420 -50124 23444 -50090
rect 22600 -50178 22616 -50144
rect 23172 -50178 23188 -50144
rect 23362 -50148 23444 -50124
rect 24380 -50090 24462 -50066
rect 24636 -50070 24652 -50036
rect 25208 -50070 25224 -50036
rect 24380 -50124 24404 -50090
rect 24438 -50124 24462 -50090
rect 23618 -50178 23634 -50144
rect 24190 -50178 24206 -50144
rect 24380 -50148 24462 -50124
rect 25408 -50090 25490 -50066
rect 25408 -50124 25432 -50090
rect 25466 -50124 25490 -50090
rect 24636 -50178 24652 -50144
rect 25208 -50178 25224 -50144
rect 25408 -50148 25490 -50124
rect 16260 -50228 16294 -50212
rect 16260 -50820 16294 -50804
rect 17278 -50228 17312 -50212
rect 17278 -50820 17312 -50804
rect 18296 -50228 18330 -50212
rect 18296 -50820 18330 -50804
rect 19314 -50228 19348 -50212
rect 19314 -50820 19348 -50804
rect 20332 -50228 20366 -50212
rect 20332 -50820 20366 -50804
rect 21350 -50228 21384 -50212
rect 21350 -50820 21384 -50804
rect 22368 -50228 22402 -50212
rect 22368 -50820 22402 -50804
rect 23386 -50228 23420 -50212
rect 23386 -50820 23420 -50804
rect 24404 -50228 24438 -50212
rect 24404 -50820 24438 -50804
rect 25422 -50228 25456 -50212
rect 28024 -50514 28058 -50498
rect 29042 -49922 29076 -49906
rect 29042 -50514 29076 -50498
rect 30060 -49922 30094 -49906
rect 30060 -50514 30094 -50498
rect 31078 -49922 31112 -49906
rect 31078 -50514 31112 -50498
rect 32096 -49922 32130 -49906
rect 32096 -50514 32130 -50498
rect 33114 -49922 33148 -49906
rect 33114 -50514 33148 -50498
rect 34132 -49922 34166 -49906
rect 34132 -50514 34166 -50498
rect 35150 -49922 35184 -49906
rect 35150 -50514 35184 -50498
rect 36168 -49922 36202 -49906
rect 36168 -50514 36202 -50498
rect 37186 -49922 37220 -49906
rect 37186 -50514 37220 -50498
rect 38204 -49922 38238 -49906
rect 38204 -50514 38238 -50498
rect 39222 -49922 39256 -49906
rect 39222 -50514 39256 -50498
rect 40240 -49922 40274 -49906
rect 40240 -50514 40274 -50498
rect 41258 -49922 41292 -49906
rect 41258 -50514 41292 -50498
rect 42276 -49922 42310 -49906
rect 42276 -50514 42310 -50498
rect 43294 -49922 43328 -49906
rect 43294 -50514 43328 -50498
rect 44312 -49922 44346 -49906
rect 44312 -50514 44346 -50498
rect 45330 -49922 45364 -49906
rect 45330 -50514 45364 -50498
rect 46348 -49922 46382 -49906
rect 46348 -50514 46382 -50498
rect 47366 -49922 47400 -49906
rect 47366 -50514 47400 -50498
rect 48384 -49922 48418 -49906
rect 48384 -50514 48418 -50498
rect 28256 -50582 28272 -50548
rect 28828 -50582 28844 -50548
rect 29274 -50582 29290 -50548
rect 29846 -50582 29862 -50548
rect 30292 -50582 30308 -50548
rect 30864 -50582 30880 -50548
rect 31310 -50582 31326 -50548
rect 31882 -50582 31898 -50548
rect 32328 -50582 32344 -50548
rect 32900 -50582 32916 -50548
rect 33346 -50582 33362 -50548
rect 33918 -50582 33934 -50548
rect 34364 -50582 34380 -50548
rect 34936 -50582 34952 -50548
rect 35382 -50582 35398 -50548
rect 35954 -50582 35970 -50548
rect 36400 -50582 36416 -50548
rect 36972 -50582 36988 -50548
rect 37418 -50582 37434 -50548
rect 37990 -50582 38006 -50548
rect 38436 -50582 38452 -50548
rect 39008 -50582 39024 -50548
rect 39454 -50582 39470 -50548
rect 40026 -50582 40042 -50548
rect 40472 -50582 40488 -50548
rect 41044 -50582 41060 -50548
rect 41490 -50582 41506 -50548
rect 42062 -50582 42078 -50548
rect 42508 -50582 42524 -50548
rect 43080 -50582 43096 -50548
rect 43526 -50582 43542 -50548
rect 44098 -50582 44114 -50548
rect 44544 -50582 44560 -50548
rect 45116 -50582 45132 -50548
rect 45562 -50582 45578 -50548
rect 46134 -50582 46150 -50548
rect 46580 -50582 46596 -50548
rect 47152 -50582 47168 -50548
rect 47598 -50582 47614 -50548
rect 48170 -50582 48186 -50548
rect 25422 -50820 25456 -50804
rect 28530 -50790 28612 -50766
rect 28530 -50824 28554 -50790
rect 28588 -50824 28612 -50790
rect 28530 -50848 28612 -50824
rect 29548 -50790 29630 -50766
rect 29548 -50824 29572 -50790
rect 29606 -50824 29630 -50790
rect 29548 -50848 29630 -50824
rect 30566 -50790 30648 -50766
rect 30566 -50824 30590 -50790
rect 30624 -50824 30648 -50790
rect 30566 -50848 30648 -50824
rect 31584 -50790 31666 -50766
rect 31584 -50824 31608 -50790
rect 31642 -50824 31666 -50790
rect 31584 -50848 31666 -50824
rect 32602 -50790 32684 -50766
rect 32602 -50824 32626 -50790
rect 32660 -50824 32684 -50790
rect 32602 -50848 32684 -50824
rect 33620 -50790 33702 -50766
rect 33620 -50824 33644 -50790
rect 33678 -50824 33702 -50790
rect 33620 -50848 33702 -50824
rect 34638 -50790 34720 -50766
rect 34638 -50824 34662 -50790
rect 34696 -50824 34720 -50790
rect 34638 -50848 34720 -50824
rect 35656 -50790 35738 -50766
rect 35656 -50824 35680 -50790
rect 35714 -50824 35738 -50790
rect 35656 -50848 35738 -50824
rect 36674 -50790 36756 -50766
rect 36674 -50824 36698 -50790
rect 36732 -50824 36756 -50790
rect 36674 -50848 36756 -50824
rect 37692 -50790 37774 -50766
rect 37692 -50824 37716 -50790
rect 37750 -50824 37774 -50790
rect 37692 -50848 37774 -50824
rect 38710 -50790 38792 -50766
rect 38710 -50824 38734 -50790
rect 38768 -50824 38792 -50790
rect 38710 -50848 38792 -50824
rect 39728 -50790 39810 -50766
rect 39728 -50824 39752 -50790
rect 39786 -50824 39810 -50790
rect 39728 -50848 39810 -50824
rect 40746 -50790 40828 -50766
rect 40746 -50824 40770 -50790
rect 40804 -50824 40828 -50790
rect 40746 -50848 40828 -50824
rect 41764 -50790 41846 -50766
rect 41764 -50824 41788 -50790
rect 41822 -50824 41846 -50790
rect 41764 -50848 41846 -50824
rect 42782 -50790 42864 -50766
rect 42782 -50824 42806 -50790
rect 42840 -50824 42864 -50790
rect 42782 -50848 42864 -50824
rect 43800 -50790 43882 -50766
rect 43800 -50824 43824 -50790
rect 43858 -50824 43882 -50790
rect 43800 -50848 43882 -50824
rect 44818 -50790 44900 -50766
rect 44818 -50824 44842 -50790
rect 44876 -50824 44900 -50790
rect 44818 -50848 44900 -50824
rect 45836 -50790 45918 -50766
rect 45836 -50824 45860 -50790
rect 45894 -50824 45918 -50790
rect 45836 -50848 45918 -50824
rect 46854 -50790 46936 -50766
rect 46854 -50824 46878 -50790
rect 46912 -50824 46936 -50790
rect 46854 -50848 46936 -50824
rect 47872 -50790 47954 -50766
rect 47872 -50824 47896 -50790
rect 47930 -50824 47954 -50790
rect 47872 -50848 47954 -50824
rect 16492 -50888 16508 -50854
rect 17064 -50888 17080 -50854
rect 17510 -50888 17526 -50854
rect 18082 -50888 18098 -50854
rect 18528 -50888 18544 -50854
rect 19100 -50888 19116 -50854
rect 19546 -50888 19562 -50854
rect 20118 -50888 20134 -50854
rect 20564 -50888 20580 -50854
rect 21136 -50888 21152 -50854
rect 21582 -50888 21598 -50854
rect 22154 -50888 22170 -50854
rect 22600 -50888 22616 -50854
rect 23172 -50888 23188 -50854
rect 23618 -50888 23634 -50854
rect 24190 -50888 24206 -50854
rect 24636 -50888 24652 -50854
rect 25208 -50888 25224 -50854
rect 16224 -50984 16306 -50960
rect 16224 -51018 16248 -50984
rect 16282 -51018 16306 -50984
rect 16224 -51042 16306 -51018
rect 17242 -50984 17324 -50960
rect 17242 -51018 17266 -50984
rect 17300 -51018 17324 -50984
rect 17242 -51042 17324 -51018
rect 18260 -50984 18342 -50960
rect 18260 -51018 18284 -50984
rect 18318 -51018 18342 -50984
rect 18260 -51042 18342 -51018
rect 19278 -50984 19360 -50960
rect 19278 -51018 19302 -50984
rect 19336 -51018 19360 -50984
rect 19278 -51042 19360 -51018
rect 20296 -50984 20378 -50960
rect 20296 -51018 20320 -50984
rect 20354 -51018 20378 -50984
rect 20296 -51042 20378 -51018
rect 21314 -50984 21396 -50960
rect 21314 -51018 21338 -50984
rect 21372 -51018 21396 -50984
rect 21314 -51042 21396 -51018
rect 22332 -50984 22414 -50960
rect 22332 -51018 22356 -50984
rect 22390 -51018 22414 -50984
rect 22332 -51042 22414 -51018
rect 23350 -50984 23432 -50960
rect 23350 -51018 23374 -50984
rect 23408 -51018 23432 -50984
rect 23350 -51042 23432 -51018
rect 24368 -50984 24450 -50960
rect 24368 -51018 24392 -50984
rect 24426 -51018 24450 -50984
rect 24368 -51042 24450 -51018
rect 25396 -50984 25478 -50960
rect 25396 -51018 25420 -50984
rect 25454 -51018 25478 -50984
rect 25396 -51042 25478 -51018
rect 28256 -51104 28272 -51070
rect 28828 -51104 28844 -51070
rect 29274 -51104 29290 -51070
rect 29846 -51104 29862 -51070
rect 30292 -51104 30308 -51070
rect 30864 -51104 30880 -51070
rect 31310 -51104 31326 -51070
rect 31882 -51104 31898 -51070
rect 32328 -51104 32344 -51070
rect 32900 -51104 32916 -51070
rect 33346 -51104 33362 -51070
rect 33918 -51104 33934 -51070
rect 34364 -51104 34380 -51070
rect 34936 -51104 34952 -51070
rect 35382 -51104 35398 -51070
rect 35954 -51104 35970 -51070
rect 36400 -51104 36416 -51070
rect 36972 -51104 36988 -51070
rect 37418 -51104 37434 -51070
rect 37990 -51104 38006 -51070
rect 38436 -51104 38452 -51070
rect 39008 -51104 39024 -51070
rect 39454 -51104 39470 -51070
rect 40026 -51104 40042 -51070
rect 40472 -51104 40488 -51070
rect 41044 -51104 41060 -51070
rect 41490 -51104 41506 -51070
rect 42062 -51104 42078 -51070
rect 42508 -51104 42524 -51070
rect 43080 -51104 43096 -51070
rect 43526 -51104 43542 -51070
rect 44098 -51104 44114 -51070
rect 44544 -51104 44560 -51070
rect 45116 -51104 45132 -51070
rect 45562 -51104 45578 -51070
rect 46134 -51104 46150 -51070
rect 46580 -51104 46596 -51070
rect 47152 -51104 47168 -51070
rect 47598 -51104 47614 -51070
rect 48170 -51104 48186 -51070
rect 28024 -51154 28058 -51138
rect 28024 -51746 28058 -51730
rect 29042 -51154 29076 -51138
rect 29042 -51746 29076 -51730
rect 30060 -51154 30094 -51138
rect 30060 -51746 30094 -51730
rect 31078 -51154 31112 -51138
rect 31078 -51746 31112 -51730
rect 32096 -51154 32130 -51138
rect 32096 -51746 32130 -51730
rect 33114 -51154 33148 -51138
rect 33114 -51746 33148 -51730
rect 34132 -51154 34166 -51138
rect 34132 -51746 34166 -51730
rect 35150 -51154 35184 -51138
rect 35150 -51746 35184 -51730
rect 36168 -51154 36202 -51138
rect 36168 -51746 36202 -51730
rect 37186 -51154 37220 -51138
rect 37186 -51746 37220 -51730
rect 38204 -51154 38238 -51138
rect 38204 -51746 38238 -51730
rect 39222 -51154 39256 -51138
rect 39222 -51746 39256 -51730
rect 40240 -51154 40274 -51138
rect 40240 -51746 40274 -51730
rect 41258 -51154 41292 -51138
rect 41258 -51746 41292 -51730
rect 42276 -51154 42310 -51138
rect 42276 -51746 42310 -51730
rect 43294 -51154 43328 -51138
rect 43294 -51746 43328 -51730
rect 44312 -51154 44346 -51138
rect 44312 -51746 44346 -51730
rect 45330 -51154 45364 -51138
rect 45330 -51746 45364 -51730
rect 46348 -51154 46382 -51138
rect 46348 -51746 46382 -51730
rect 47366 -51154 47400 -51138
rect 47366 -51746 47400 -51730
rect 48384 -51154 48418 -51138
rect 48384 -51746 48418 -51730
rect 36674 -51780 36734 -51778
rect 38718 -51780 38778 -51776
rect 46852 -51780 46912 -51778
rect 28256 -51814 28272 -51780
rect 28828 -51814 28844 -51780
rect 29274 -51814 29290 -51780
rect 29846 -51814 29862 -51780
rect 30292 -51814 30308 -51780
rect 30864 -51814 30880 -51780
rect 31310 -51814 31326 -51780
rect 31882 -51814 31898 -51780
rect 32328 -51814 32344 -51780
rect 32900 -51814 32916 -51780
rect 33346 -51814 33362 -51780
rect 33918 -51814 33934 -51780
rect 34364 -51814 34380 -51780
rect 34936 -51814 34952 -51780
rect 35382 -51814 35398 -51780
rect 35954 -51814 35970 -51780
rect 36400 -51814 36416 -51780
rect 36972 -51814 36988 -51780
rect 37418 -51814 37434 -51780
rect 37990 -51814 38006 -51780
rect 38436 -51814 38452 -51780
rect 39008 -51814 39024 -51780
rect 39454 -51814 39470 -51780
rect 40026 -51814 40042 -51780
rect 40472 -51814 40488 -51780
rect 41044 -51814 41060 -51780
rect 41490 -51814 41506 -51780
rect 42062 -51814 42078 -51780
rect 42508 -51814 42524 -51780
rect 43080 -51814 43096 -51780
rect 43526 -51814 43542 -51780
rect 44098 -51814 44114 -51780
rect 44544 -51814 44560 -51780
rect 45116 -51814 45132 -51780
rect 45562 -51814 45578 -51780
rect 46134 -51814 46150 -51780
rect 46580 -51814 46596 -51780
rect 47152 -51814 47168 -51780
rect 47598 -51814 47614 -51780
rect 48170 -51814 48186 -51780
rect 15428 -51932 15510 -51908
rect 15428 -51966 15452 -51932
rect 15486 -51966 15510 -51932
rect 15428 -51990 15510 -51966
rect 16446 -51932 16528 -51908
rect 16446 -51966 16470 -51932
rect 16504 -51966 16528 -51932
rect 16446 -51990 16528 -51966
rect 17464 -51932 17546 -51908
rect 17464 -51966 17488 -51932
rect 17522 -51966 17546 -51932
rect 17464 -51990 17546 -51966
rect 18482 -51932 18564 -51908
rect 18482 -51966 18506 -51932
rect 18540 -51966 18564 -51932
rect 18482 -51990 18564 -51966
rect 19500 -51932 19582 -51908
rect 19500 -51966 19524 -51932
rect 19558 -51966 19582 -51932
rect 19500 -51990 19582 -51966
rect 20518 -51932 20600 -51908
rect 20518 -51966 20542 -51932
rect 20576 -51966 20600 -51932
rect 20518 -51990 20600 -51966
rect 21536 -51932 21618 -51908
rect 21536 -51966 21560 -51932
rect 21594 -51966 21618 -51932
rect 21536 -51990 21618 -51966
rect 22554 -51932 22636 -51908
rect 22554 -51966 22578 -51932
rect 22612 -51966 22636 -51932
rect 22554 -51990 22636 -51966
rect 23572 -51932 23654 -51908
rect 23572 -51966 23596 -51932
rect 23630 -51966 23654 -51932
rect 23572 -51990 23654 -51966
rect 24590 -51932 24672 -51908
rect 24590 -51966 24614 -51932
rect 24648 -51966 24672 -51932
rect 24590 -51990 24672 -51966
rect 25608 -51932 25690 -51908
rect 25608 -51966 25632 -51932
rect 25666 -51966 25690 -51932
rect 25608 -51990 25690 -51966
rect 28530 -52038 28612 -52014
rect 28530 -52072 28554 -52038
rect 28588 -52072 28612 -52038
rect 28530 -52096 28612 -52072
rect 29548 -52038 29630 -52014
rect 29548 -52072 29572 -52038
rect 29606 -52072 29630 -52038
rect 29548 -52096 29630 -52072
rect 30566 -52038 30648 -52014
rect 30566 -52072 30590 -52038
rect 30624 -52072 30648 -52038
rect 30566 -52096 30648 -52072
rect 31584 -52038 31666 -52014
rect 31584 -52072 31608 -52038
rect 31642 -52072 31666 -52038
rect 31584 -52096 31666 -52072
rect 32602 -52038 32684 -52014
rect 32602 -52072 32626 -52038
rect 32660 -52072 32684 -52038
rect 32602 -52096 32684 -52072
rect 33620 -52038 33702 -52014
rect 33620 -52072 33644 -52038
rect 33678 -52072 33702 -52038
rect 33620 -52096 33702 -52072
rect 34638 -52038 34720 -52014
rect 34638 -52072 34662 -52038
rect 34696 -52072 34720 -52038
rect 34638 -52096 34720 -52072
rect 35656 -52038 35738 -52014
rect 35656 -52072 35680 -52038
rect 35714 -52072 35738 -52038
rect 35656 -52096 35738 -52072
rect 36674 -52038 36756 -52014
rect 36674 -52072 36698 -52038
rect 36732 -52072 36756 -52038
rect 36674 -52096 36756 -52072
rect 37692 -52038 37774 -52014
rect 37692 -52072 37716 -52038
rect 37750 -52072 37774 -52038
rect 37692 -52096 37774 -52072
rect 38710 -52038 38792 -52014
rect 38710 -52072 38734 -52038
rect 38768 -52072 38792 -52038
rect 38710 -52096 38792 -52072
rect 39728 -52038 39810 -52014
rect 39728 -52072 39752 -52038
rect 39786 -52072 39810 -52038
rect 39728 -52096 39810 -52072
rect 40746 -52038 40828 -52014
rect 40746 -52072 40770 -52038
rect 40804 -52072 40828 -52038
rect 40746 -52096 40828 -52072
rect 41764 -52038 41846 -52014
rect 41764 -52072 41788 -52038
rect 41822 -52072 41846 -52038
rect 41764 -52096 41846 -52072
rect 42782 -52038 42864 -52014
rect 42782 -52072 42806 -52038
rect 42840 -52072 42864 -52038
rect 42782 -52096 42864 -52072
rect 43800 -52038 43882 -52014
rect 43800 -52072 43824 -52038
rect 43858 -52072 43882 -52038
rect 43800 -52096 43882 -52072
rect 44818 -52038 44900 -52014
rect 44818 -52072 44842 -52038
rect 44876 -52072 44900 -52038
rect 44818 -52096 44900 -52072
rect 45836 -52038 45918 -52014
rect 45836 -52072 45860 -52038
rect 45894 -52072 45918 -52038
rect 45836 -52096 45918 -52072
rect 46854 -52038 46936 -52014
rect 46854 -52072 46878 -52038
rect 46912 -52072 46936 -52038
rect 46854 -52096 46936 -52072
rect 47872 -52038 47954 -52014
rect 47872 -52072 47896 -52038
rect 47930 -52072 47954 -52038
rect 47872 -52096 47954 -52072
rect 15168 -52202 15184 -52168
rect 15740 -52202 15756 -52168
rect 16186 -52202 16202 -52168
rect 16758 -52202 16774 -52168
rect 17204 -52202 17220 -52168
rect 17776 -52202 17792 -52168
rect 18222 -52202 18238 -52168
rect 18794 -52202 18810 -52168
rect 19240 -52202 19256 -52168
rect 19812 -52202 19828 -52168
rect 20258 -52202 20274 -52168
rect 20830 -52202 20846 -52168
rect 21276 -52202 21292 -52168
rect 21848 -52202 21864 -52168
rect 22294 -52202 22310 -52168
rect 22866 -52202 22882 -52168
rect 23312 -52202 23328 -52168
rect 23884 -52202 23900 -52168
rect 24330 -52202 24346 -52168
rect 24902 -52202 24918 -52168
rect 25348 -52202 25364 -52168
rect 25920 -52202 25936 -52168
rect 14936 -52252 14970 -52236
rect 14936 -52844 14970 -52828
rect 15954 -52252 15988 -52236
rect 15954 -52844 15988 -52828
rect 16972 -52252 17006 -52236
rect 16972 -52844 17006 -52828
rect 17990 -52252 18024 -52236
rect 17990 -52844 18024 -52828
rect 19008 -52252 19042 -52236
rect 19008 -52844 19042 -52828
rect 20026 -52252 20060 -52236
rect 20026 -52844 20060 -52828
rect 21044 -52252 21078 -52236
rect 21044 -52844 21078 -52828
rect 22062 -52252 22096 -52236
rect 22062 -52844 22096 -52828
rect 23080 -52252 23114 -52236
rect 23080 -52844 23114 -52828
rect 24098 -52252 24132 -52236
rect 24098 -52844 24132 -52828
rect 25116 -52252 25150 -52236
rect 25116 -52844 25150 -52828
rect 26134 -52252 26168 -52236
rect 28256 -52338 28272 -52304
rect 28828 -52338 28844 -52304
rect 29274 -52338 29290 -52304
rect 29846 -52338 29862 -52304
rect 30292 -52338 30308 -52304
rect 30864 -52338 30880 -52304
rect 31310 -52338 31326 -52304
rect 31882 -52338 31898 -52304
rect 32328 -52338 32344 -52304
rect 32900 -52338 32916 -52304
rect 33346 -52338 33362 -52304
rect 33918 -52338 33934 -52304
rect 34364 -52338 34380 -52304
rect 34936 -52338 34952 -52304
rect 35382 -52338 35398 -52304
rect 35954 -52338 35970 -52304
rect 36400 -52338 36416 -52304
rect 36972 -52338 36988 -52304
rect 37418 -52338 37434 -52304
rect 37990 -52338 38006 -52304
rect 38436 -52338 38452 -52304
rect 39008 -52338 39024 -52304
rect 39454 -52338 39470 -52304
rect 40026 -52338 40042 -52304
rect 40472 -52338 40488 -52304
rect 41044 -52338 41060 -52304
rect 41490 -52338 41506 -52304
rect 42062 -52338 42078 -52304
rect 42508 -52338 42524 -52304
rect 43080 -52338 43096 -52304
rect 43526 -52338 43542 -52304
rect 44098 -52338 44114 -52304
rect 44544 -52338 44560 -52304
rect 45116 -52338 45132 -52304
rect 45562 -52338 45578 -52304
rect 46134 -52338 46150 -52304
rect 46580 -52338 46596 -52304
rect 47152 -52338 47168 -52304
rect 47598 -52338 47614 -52304
rect 48170 -52338 48186 -52304
rect 26134 -52844 26168 -52828
rect 28024 -52388 28058 -52372
rect 15168 -52912 15184 -52878
rect 15740 -52912 15756 -52878
rect 16186 -52912 16202 -52878
rect 16758 -52912 16774 -52878
rect 17204 -52912 17220 -52878
rect 17776 -52912 17792 -52878
rect 18222 -52912 18238 -52878
rect 18794 -52912 18810 -52878
rect 19240 -52912 19256 -52878
rect 19812 -52912 19828 -52878
rect 20258 -52912 20274 -52878
rect 20830 -52912 20846 -52878
rect 21276 -52912 21292 -52878
rect 21848 -52912 21864 -52878
rect 22294 -52912 22310 -52878
rect 22866 -52912 22882 -52878
rect 23312 -52912 23328 -52878
rect 23884 -52912 23900 -52878
rect 24330 -52912 24346 -52878
rect 24902 -52912 24918 -52878
rect 25348 -52912 25364 -52878
rect 25920 -52912 25936 -52878
rect 28024 -52980 28058 -52964
rect 29042 -52388 29076 -52372
rect 29042 -52980 29076 -52964
rect 30060 -52388 30094 -52372
rect 30060 -52980 30094 -52964
rect 31078 -52388 31112 -52372
rect 31078 -52980 31112 -52964
rect 32096 -52388 32130 -52372
rect 32096 -52980 32130 -52964
rect 33114 -52388 33148 -52372
rect 33114 -52980 33148 -52964
rect 34132 -52388 34166 -52372
rect 34132 -52980 34166 -52964
rect 35150 -52388 35184 -52372
rect 35150 -52980 35184 -52964
rect 36168 -52388 36202 -52372
rect 36168 -52980 36202 -52964
rect 37186 -52388 37220 -52372
rect 37186 -52980 37220 -52964
rect 38204 -52388 38238 -52372
rect 38204 -52980 38238 -52964
rect 39222 -52388 39256 -52372
rect 39222 -52980 39256 -52964
rect 40240 -52388 40274 -52372
rect 40240 -52980 40274 -52964
rect 41258 -52388 41292 -52372
rect 41258 -52980 41292 -52964
rect 42276 -52388 42310 -52372
rect 42276 -52980 42310 -52964
rect 43294 -52388 43328 -52372
rect 43294 -52980 43328 -52964
rect 44312 -52388 44346 -52372
rect 44312 -52980 44346 -52964
rect 45330 -52388 45364 -52372
rect 45330 -52980 45364 -52964
rect 46348 -52388 46382 -52372
rect 46348 -52980 46382 -52964
rect 47366 -52388 47400 -52372
rect 47366 -52980 47400 -52964
rect 48384 -52388 48418 -52372
rect 48384 -52980 48418 -52964
rect 30550 -53014 30610 -53010
rect 28256 -53048 28272 -53014
rect 28828 -53048 28844 -53014
rect 29274 -53048 29290 -53014
rect 29846 -53048 29862 -53014
rect 30292 -53048 30308 -53014
rect 30864 -53048 30880 -53014
rect 31310 -53048 31326 -53014
rect 31882 -53048 31898 -53014
rect 32328 -53048 32344 -53014
rect 32900 -53048 32916 -53014
rect 33346 -53048 33362 -53014
rect 33918 -53048 33934 -53014
rect 34364 -53048 34380 -53014
rect 34936 -53048 34952 -53014
rect 35382 -53048 35398 -53014
rect 35954 -53048 35970 -53014
rect 36400 -53048 36416 -53014
rect 36972 -53048 36988 -53014
rect 37418 -53048 37434 -53014
rect 37990 -53048 38006 -53014
rect 38436 -53048 38452 -53014
rect 39008 -53048 39024 -53014
rect 39454 -53048 39470 -53014
rect 40026 -53048 40042 -53014
rect 40472 -53048 40488 -53014
rect 41044 -53048 41060 -53014
rect 41490 -53048 41506 -53014
rect 42062 -53048 42078 -53014
rect 42508 -53048 42524 -53014
rect 43080 -53048 43096 -53014
rect 43526 -53048 43542 -53014
rect 44098 -53048 44114 -53014
rect 44544 -53048 44560 -53014
rect 45116 -53048 45132 -53014
rect 45562 -53048 45578 -53014
rect 46134 -53048 46150 -53014
rect 46580 -53048 46596 -53014
rect 47152 -53048 47168 -53014
rect 47598 -53048 47614 -53014
rect 48170 -53048 48186 -53014
rect 15440 -53074 15522 -53050
rect 15440 -53108 15464 -53074
rect 15498 -53108 15522 -53074
rect 15440 -53132 15522 -53108
rect 16458 -53074 16540 -53050
rect 16458 -53108 16482 -53074
rect 16516 -53108 16540 -53074
rect 16458 -53132 16540 -53108
rect 17476 -53074 17558 -53050
rect 17476 -53108 17500 -53074
rect 17534 -53108 17558 -53074
rect 17476 -53132 17558 -53108
rect 18494 -53074 18576 -53050
rect 18494 -53108 18518 -53074
rect 18552 -53108 18576 -53074
rect 18494 -53132 18576 -53108
rect 19512 -53074 19594 -53050
rect 19512 -53108 19536 -53074
rect 19570 -53108 19594 -53074
rect 19512 -53132 19594 -53108
rect 20530 -53074 20612 -53050
rect 20530 -53108 20554 -53074
rect 20588 -53108 20612 -53074
rect 20530 -53132 20612 -53108
rect 21548 -53074 21630 -53050
rect 21548 -53108 21572 -53074
rect 21606 -53108 21630 -53074
rect 21548 -53132 21630 -53108
rect 22566 -53074 22648 -53050
rect 22566 -53108 22590 -53074
rect 22624 -53108 22648 -53074
rect 22566 -53132 22648 -53108
rect 23584 -53074 23666 -53050
rect 23584 -53108 23608 -53074
rect 23642 -53108 23666 -53074
rect 23584 -53132 23666 -53108
rect 24602 -53074 24684 -53050
rect 24602 -53108 24626 -53074
rect 24660 -53108 24684 -53074
rect 24602 -53132 24684 -53108
rect 25620 -53074 25702 -53050
rect 25620 -53108 25644 -53074
rect 25678 -53108 25702 -53074
rect 25620 -53132 25702 -53108
rect 28506 -53274 28588 -53250
rect 15168 -53314 15184 -53280
rect 15740 -53314 15756 -53280
rect 16186 -53314 16202 -53280
rect 16758 -53314 16774 -53280
rect 17204 -53314 17220 -53280
rect 17776 -53314 17792 -53280
rect 18222 -53314 18238 -53280
rect 18794 -53314 18810 -53280
rect 19240 -53314 19256 -53280
rect 19812 -53314 19828 -53280
rect 20258 -53314 20274 -53280
rect 20830 -53314 20846 -53280
rect 21276 -53314 21292 -53280
rect 21848 -53314 21864 -53280
rect 22294 -53314 22310 -53280
rect 22866 -53314 22882 -53280
rect 23312 -53314 23328 -53280
rect 23884 -53314 23900 -53280
rect 24330 -53314 24346 -53280
rect 24902 -53314 24918 -53280
rect 25348 -53314 25364 -53280
rect 25920 -53314 25936 -53280
rect 28506 -53308 28530 -53274
rect 28564 -53308 28588 -53274
rect 28506 -53332 28588 -53308
rect 29524 -53274 29606 -53250
rect 29524 -53308 29548 -53274
rect 29582 -53308 29606 -53274
rect 29524 -53332 29606 -53308
rect 30542 -53274 30624 -53250
rect 30542 -53308 30566 -53274
rect 30600 -53308 30624 -53274
rect 30542 -53332 30624 -53308
rect 31560 -53274 31642 -53250
rect 31560 -53308 31584 -53274
rect 31618 -53308 31642 -53274
rect 31560 -53332 31642 -53308
rect 32578 -53274 32660 -53250
rect 32578 -53308 32602 -53274
rect 32636 -53308 32660 -53274
rect 32578 -53332 32660 -53308
rect 33596 -53274 33678 -53250
rect 33596 -53308 33620 -53274
rect 33654 -53308 33678 -53274
rect 33596 -53332 33678 -53308
rect 34614 -53274 34696 -53250
rect 34614 -53308 34638 -53274
rect 34672 -53308 34696 -53274
rect 34614 -53332 34696 -53308
rect 35632 -53274 35714 -53250
rect 35632 -53308 35656 -53274
rect 35690 -53308 35714 -53274
rect 35632 -53332 35714 -53308
rect 36650 -53274 36732 -53250
rect 36650 -53308 36674 -53274
rect 36708 -53308 36732 -53274
rect 36650 -53332 36732 -53308
rect 37668 -53274 37750 -53250
rect 37668 -53308 37692 -53274
rect 37726 -53308 37750 -53274
rect 37668 -53332 37750 -53308
rect 38686 -53274 38768 -53250
rect 38686 -53308 38710 -53274
rect 38744 -53308 38768 -53274
rect 38686 -53332 38768 -53308
rect 39704 -53274 39786 -53250
rect 39704 -53308 39728 -53274
rect 39762 -53308 39786 -53274
rect 39704 -53332 39786 -53308
rect 40722 -53274 40804 -53250
rect 40722 -53308 40746 -53274
rect 40780 -53308 40804 -53274
rect 40722 -53332 40804 -53308
rect 41740 -53274 41822 -53250
rect 41740 -53308 41764 -53274
rect 41798 -53308 41822 -53274
rect 41740 -53332 41822 -53308
rect 42758 -53274 42840 -53250
rect 42758 -53308 42782 -53274
rect 42816 -53308 42840 -53274
rect 42758 -53332 42840 -53308
rect 43776 -53274 43858 -53250
rect 43776 -53308 43800 -53274
rect 43834 -53308 43858 -53274
rect 43776 -53332 43858 -53308
rect 44794 -53274 44876 -53250
rect 44794 -53308 44818 -53274
rect 44852 -53308 44876 -53274
rect 44794 -53332 44876 -53308
rect 45812 -53274 45894 -53250
rect 45812 -53308 45836 -53274
rect 45870 -53308 45894 -53274
rect 45812 -53332 45894 -53308
rect 46830 -53274 46912 -53250
rect 46830 -53308 46854 -53274
rect 46888 -53308 46912 -53274
rect 46830 -53332 46912 -53308
rect 47848 -53274 47930 -53250
rect 47848 -53308 47872 -53274
rect 47906 -53308 47930 -53274
rect 47848 -53332 47930 -53308
rect 14936 -53364 14970 -53348
rect 14936 -53956 14970 -53940
rect 15954 -53364 15988 -53348
rect 15954 -53956 15988 -53940
rect 16972 -53364 17006 -53348
rect 16972 -53956 17006 -53940
rect 17990 -53364 18024 -53348
rect 17990 -53956 18024 -53940
rect 19008 -53364 19042 -53348
rect 19008 -53956 19042 -53940
rect 20026 -53364 20060 -53348
rect 20026 -53956 20060 -53940
rect 21044 -53364 21078 -53348
rect 21044 -53956 21078 -53940
rect 22062 -53364 22096 -53348
rect 22062 -53956 22096 -53940
rect 23080 -53364 23114 -53348
rect 23080 -53956 23114 -53940
rect 24098 -53364 24132 -53348
rect 24098 -53956 24132 -53940
rect 25116 -53364 25150 -53348
rect 25116 -53956 25150 -53940
rect 26134 -53364 26168 -53348
rect 28256 -53572 28272 -53538
rect 28828 -53572 28844 -53538
rect 29274 -53572 29290 -53538
rect 29846 -53572 29862 -53538
rect 30292 -53572 30308 -53538
rect 30864 -53572 30880 -53538
rect 31310 -53572 31326 -53538
rect 31882 -53572 31898 -53538
rect 32328 -53572 32344 -53538
rect 32900 -53572 32916 -53538
rect 33346 -53572 33362 -53538
rect 33918 -53572 33934 -53538
rect 34364 -53572 34380 -53538
rect 34936 -53572 34952 -53538
rect 35382 -53572 35398 -53538
rect 35954 -53572 35970 -53538
rect 36400 -53572 36416 -53538
rect 36972 -53572 36988 -53538
rect 37418 -53572 37434 -53538
rect 37990 -53572 38006 -53538
rect 38436 -53572 38452 -53538
rect 39008 -53572 39024 -53538
rect 39454 -53572 39470 -53538
rect 40026 -53572 40042 -53538
rect 40472 -53572 40488 -53538
rect 41044 -53572 41060 -53538
rect 41490 -53572 41506 -53538
rect 42062 -53572 42078 -53538
rect 42508 -53572 42524 -53538
rect 43080 -53572 43096 -53538
rect 43526 -53572 43542 -53538
rect 44098 -53572 44114 -53538
rect 44544 -53572 44560 -53538
rect 45116 -53572 45132 -53538
rect 45562 -53572 45578 -53538
rect 46134 -53572 46150 -53538
rect 46580 -53572 46596 -53538
rect 47152 -53572 47168 -53538
rect 47598 -53572 47614 -53538
rect 48170 -53572 48186 -53538
rect 26134 -53956 26168 -53940
rect 28024 -53622 28058 -53606
rect 15168 -54024 15184 -53990
rect 15740 -54024 15756 -53990
rect 16186 -54024 16202 -53990
rect 16758 -54024 16774 -53990
rect 17204 -54024 17220 -53990
rect 17776 -54024 17792 -53990
rect 18222 -54024 18238 -53990
rect 18794 -54024 18810 -53990
rect 19240 -54024 19256 -53990
rect 19812 -54024 19828 -53990
rect 20258 -54024 20274 -53990
rect 20830 -54024 20846 -53990
rect 21276 -54024 21292 -53990
rect 21848 -54024 21864 -53990
rect 22294 -54024 22310 -53990
rect 22866 -54024 22882 -53990
rect 23312 -54024 23328 -53990
rect 23884 -54024 23900 -53990
rect 24330 -54024 24346 -53990
rect 24902 -54024 24918 -53990
rect 25348 -54024 25364 -53990
rect 25920 -54024 25936 -53990
rect 15418 -54182 15500 -54158
rect 15418 -54216 15442 -54182
rect 15476 -54216 15500 -54182
rect 15418 -54240 15500 -54216
rect 16436 -54182 16518 -54158
rect 16436 -54216 16460 -54182
rect 16494 -54216 16518 -54182
rect 16436 -54240 16518 -54216
rect 17454 -54182 17536 -54158
rect 17454 -54216 17478 -54182
rect 17512 -54216 17536 -54182
rect 17454 -54240 17536 -54216
rect 18472 -54182 18554 -54158
rect 18472 -54216 18496 -54182
rect 18530 -54216 18554 -54182
rect 18472 -54240 18554 -54216
rect 19490 -54182 19572 -54158
rect 19490 -54216 19514 -54182
rect 19548 -54216 19572 -54182
rect 19490 -54240 19572 -54216
rect 20508 -54182 20590 -54158
rect 20508 -54216 20532 -54182
rect 20566 -54216 20590 -54182
rect 20508 -54240 20590 -54216
rect 21526 -54182 21608 -54158
rect 21526 -54216 21550 -54182
rect 21584 -54216 21608 -54182
rect 21526 -54240 21608 -54216
rect 22544 -54182 22626 -54158
rect 22544 -54216 22568 -54182
rect 22602 -54216 22626 -54182
rect 22544 -54240 22626 -54216
rect 23562 -54182 23644 -54158
rect 23562 -54216 23586 -54182
rect 23620 -54216 23644 -54182
rect 23562 -54240 23644 -54216
rect 24580 -54182 24662 -54158
rect 24580 -54216 24604 -54182
rect 24638 -54216 24662 -54182
rect 24580 -54240 24662 -54216
rect 25598 -54182 25680 -54158
rect 25598 -54216 25622 -54182
rect 25656 -54216 25680 -54182
rect 28024 -54214 28058 -54198
rect 29042 -53622 29076 -53606
rect 29042 -54214 29076 -54198
rect 30060 -53622 30094 -53606
rect 30060 -54214 30094 -54198
rect 31078 -53622 31112 -53606
rect 31078 -54214 31112 -54198
rect 32096 -53622 32130 -53606
rect 32096 -54214 32130 -54198
rect 33114 -53622 33148 -53606
rect 33114 -54214 33148 -54198
rect 34132 -53622 34166 -53606
rect 34132 -54214 34166 -54198
rect 35150 -53622 35184 -53606
rect 35150 -54214 35184 -54198
rect 36168 -53622 36202 -53606
rect 36168 -54214 36202 -54198
rect 37186 -53622 37220 -53606
rect 37186 -54214 37220 -54198
rect 38204 -53622 38238 -53606
rect 38204 -54214 38238 -54198
rect 39222 -53622 39256 -53606
rect 39222 -54214 39256 -54198
rect 40240 -53622 40274 -53606
rect 40240 -54214 40274 -54198
rect 41258 -53622 41292 -53606
rect 41258 -54214 41292 -54198
rect 42276 -53622 42310 -53606
rect 42276 -54214 42310 -54198
rect 43294 -53622 43328 -53606
rect 43294 -54214 43328 -54198
rect 44312 -53622 44346 -53606
rect 44312 -54214 44346 -54198
rect 45330 -53622 45364 -53606
rect 45330 -54214 45364 -54198
rect 46348 -53622 46382 -53606
rect 46348 -54214 46382 -54198
rect 47366 -53622 47400 -53606
rect 47366 -54214 47400 -54198
rect 48384 -53622 48418 -53606
rect 48384 -54214 48418 -54198
rect 25598 -54240 25680 -54216
rect 36674 -54248 36734 -54246
rect 38718 -54248 38778 -54244
rect 41756 -54248 41816 -54244
rect 28256 -54282 28272 -54248
rect 28828 -54282 28844 -54248
rect 29274 -54282 29290 -54248
rect 29846 -54282 29862 -54248
rect 30292 -54282 30308 -54248
rect 30864 -54282 30880 -54248
rect 31310 -54282 31326 -54248
rect 31882 -54282 31898 -54248
rect 32328 -54282 32344 -54248
rect 32900 -54282 32916 -54248
rect 33346 -54282 33362 -54248
rect 33918 -54282 33934 -54248
rect 34364 -54282 34380 -54248
rect 34936 -54282 34952 -54248
rect 35382 -54282 35398 -54248
rect 35954 -54282 35970 -54248
rect 36400 -54282 36416 -54248
rect 36972 -54282 36988 -54248
rect 37418 -54282 37434 -54248
rect 37990 -54282 38006 -54248
rect 38436 -54282 38452 -54248
rect 39008 -54282 39024 -54248
rect 39454 -54282 39470 -54248
rect 40026 -54282 40042 -54248
rect 40472 -54282 40488 -54248
rect 41044 -54282 41060 -54248
rect 41490 -54282 41506 -54248
rect 42062 -54282 42078 -54248
rect 42508 -54282 42524 -54248
rect 43080 -54282 43096 -54248
rect 43526 -54282 43542 -54248
rect 44098 -54282 44114 -54248
rect 44544 -54282 44560 -54248
rect 45116 -54282 45132 -54248
rect 45562 -54282 45578 -54248
rect 46134 -54282 46150 -54248
rect 46580 -54282 46596 -54248
rect 47152 -54282 47168 -54248
rect 47598 -54282 47614 -54248
rect 48170 -54282 48186 -54248
rect 15168 -54426 15184 -54392
rect 15740 -54426 15756 -54392
rect 16186 -54426 16202 -54392
rect 16758 -54426 16774 -54392
rect 17204 -54426 17220 -54392
rect 17776 -54426 17792 -54392
rect 18222 -54426 18238 -54392
rect 18794 -54426 18810 -54392
rect 19240 -54426 19256 -54392
rect 19812 -54426 19828 -54392
rect 20258 -54426 20274 -54392
rect 20830 -54426 20846 -54392
rect 21276 -54426 21292 -54392
rect 21848 -54426 21864 -54392
rect 22294 -54426 22310 -54392
rect 22866 -54426 22882 -54392
rect 23312 -54426 23328 -54392
rect 23884 -54426 23900 -54392
rect 24330 -54426 24346 -54392
rect 24902 -54426 24918 -54392
rect 25348 -54426 25364 -54392
rect 25920 -54426 25936 -54392
rect 14936 -54476 14970 -54460
rect 14936 -55068 14970 -55052
rect 15954 -54476 15988 -54460
rect 15954 -55068 15988 -55052
rect 16972 -54476 17006 -54460
rect 16972 -55068 17006 -55052
rect 17990 -54476 18024 -54460
rect 17990 -55068 18024 -55052
rect 19008 -54476 19042 -54460
rect 19008 -55068 19042 -55052
rect 20026 -54476 20060 -54460
rect 20026 -55068 20060 -55052
rect 21044 -54476 21078 -54460
rect 21044 -55068 21078 -55052
rect 22062 -54476 22096 -54460
rect 22062 -55068 22096 -55052
rect 23080 -54476 23114 -54460
rect 23080 -55068 23114 -55052
rect 24098 -54476 24132 -54460
rect 24098 -55068 24132 -55052
rect 25116 -54476 25150 -54460
rect 25116 -55068 25150 -55052
rect 26134 -54476 26168 -54460
rect 28518 -54498 28600 -54474
rect 28518 -54532 28542 -54498
rect 28576 -54532 28600 -54498
rect 28518 -54556 28600 -54532
rect 29536 -54498 29618 -54474
rect 29536 -54532 29560 -54498
rect 29594 -54532 29618 -54498
rect 29536 -54556 29618 -54532
rect 30554 -54498 30636 -54474
rect 30554 -54532 30578 -54498
rect 30612 -54532 30636 -54498
rect 30554 -54556 30636 -54532
rect 31572 -54498 31654 -54474
rect 31572 -54532 31596 -54498
rect 31630 -54532 31654 -54498
rect 31572 -54556 31654 -54532
rect 32590 -54498 32672 -54474
rect 32590 -54532 32614 -54498
rect 32648 -54532 32672 -54498
rect 32590 -54556 32672 -54532
rect 33608 -54498 33690 -54474
rect 33608 -54532 33632 -54498
rect 33666 -54532 33690 -54498
rect 33608 -54556 33690 -54532
rect 34626 -54498 34708 -54474
rect 34626 -54532 34650 -54498
rect 34684 -54532 34708 -54498
rect 34626 -54556 34708 -54532
rect 35644 -54498 35726 -54474
rect 35644 -54532 35668 -54498
rect 35702 -54532 35726 -54498
rect 35644 -54556 35726 -54532
rect 36662 -54498 36744 -54474
rect 36662 -54532 36686 -54498
rect 36720 -54532 36744 -54498
rect 36662 -54556 36744 -54532
rect 37680 -54498 37762 -54474
rect 37680 -54532 37704 -54498
rect 37738 -54532 37762 -54498
rect 37680 -54556 37762 -54532
rect 38698 -54498 38780 -54474
rect 38698 -54532 38722 -54498
rect 38756 -54532 38780 -54498
rect 38698 -54556 38780 -54532
rect 39716 -54498 39798 -54474
rect 39716 -54532 39740 -54498
rect 39774 -54532 39798 -54498
rect 39716 -54556 39798 -54532
rect 40734 -54498 40816 -54474
rect 40734 -54532 40758 -54498
rect 40792 -54532 40816 -54498
rect 40734 -54556 40816 -54532
rect 41752 -54498 41834 -54474
rect 41752 -54532 41776 -54498
rect 41810 -54532 41834 -54498
rect 41752 -54556 41834 -54532
rect 42770 -54498 42852 -54474
rect 42770 -54532 42794 -54498
rect 42828 -54532 42852 -54498
rect 42770 -54556 42852 -54532
rect 43788 -54498 43870 -54474
rect 43788 -54532 43812 -54498
rect 43846 -54532 43870 -54498
rect 43788 -54556 43870 -54532
rect 44806 -54498 44888 -54474
rect 44806 -54532 44830 -54498
rect 44864 -54532 44888 -54498
rect 44806 -54556 44888 -54532
rect 45824 -54498 45906 -54474
rect 45824 -54532 45848 -54498
rect 45882 -54532 45906 -54498
rect 45824 -54556 45906 -54532
rect 46842 -54498 46924 -54474
rect 46842 -54532 46866 -54498
rect 46900 -54532 46924 -54498
rect 46842 -54556 46924 -54532
rect 47860 -54498 47942 -54474
rect 47860 -54532 47884 -54498
rect 47918 -54532 47942 -54498
rect 47860 -54556 47942 -54532
rect 28256 -54804 28272 -54770
rect 28828 -54804 28844 -54770
rect 29274 -54804 29290 -54770
rect 29846 -54804 29862 -54770
rect 30292 -54804 30308 -54770
rect 30864 -54804 30880 -54770
rect 31310 -54804 31326 -54770
rect 31882 -54804 31898 -54770
rect 32328 -54804 32344 -54770
rect 32900 -54804 32916 -54770
rect 33346 -54804 33362 -54770
rect 33918 -54804 33934 -54770
rect 34364 -54804 34380 -54770
rect 34936 -54804 34952 -54770
rect 35382 -54804 35398 -54770
rect 35954 -54804 35970 -54770
rect 36400 -54804 36416 -54770
rect 36972 -54804 36988 -54770
rect 37418 -54804 37434 -54770
rect 37990 -54804 38006 -54770
rect 38436 -54804 38452 -54770
rect 39008 -54804 39024 -54770
rect 39454 -54804 39470 -54770
rect 40026 -54804 40042 -54770
rect 40472 -54804 40488 -54770
rect 41044 -54804 41060 -54770
rect 41490 -54804 41506 -54770
rect 42062 -54804 42078 -54770
rect 42508 -54804 42524 -54770
rect 43080 -54804 43096 -54770
rect 43526 -54804 43542 -54770
rect 44098 -54804 44114 -54770
rect 44544 -54804 44560 -54770
rect 45116 -54804 45132 -54770
rect 45562 -54804 45578 -54770
rect 46134 -54804 46150 -54770
rect 46580 -54804 46596 -54770
rect 47152 -54804 47168 -54770
rect 47598 -54804 47614 -54770
rect 48170 -54804 48186 -54770
rect 31578 -54806 31638 -54804
rect 26134 -55068 26168 -55052
rect 28024 -54854 28058 -54838
rect 15168 -55136 15184 -55102
rect 15740 -55136 15756 -55102
rect 16186 -55136 16202 -55102
rect 16758 -55136 16774 -55102
rect 17204 -55136 17220 -55102
rect 17776 -55136 17792 -55102
rect 18222 -55136 18238 -55102
rect 18794 -55136 18810 -55102
rect 19240 -55136 19256 -55102
rect 19812 -55136 19828 -55102
rect 20258 -55136 20274 -55102
rect 20830 -55136 20846 -55102
rect 21276 -55136 21292 -55102
rect 21848 -55136 21864 -55102
rect 22294 -55136 22310 -55102
rect 22866 -55136 22882 -55102
rect 23312 -55136 23328 -55102
rect 23884 -55136 23900 -55102
rect 24330 -55136 24346 -55102
rect 24902 -55136 24918 -55102
rect 25348 -55136 25364 -55102
rect 25920 -55136 25936 -55102
rect 15418 -55288 15500 -55264
rect 15418 -55322 15442 -55288
rect 15476 -55322 15500 -55288
rect 15418 -55346 15500 -55322
rect 16436 -55288 16518 -55264
rect 16436 -55322 16460 -55288
rect 16494 -55322 16518 -55288
rect 16436 -55346 16518 -55322
rect 17454 -55288 17536 -55264
rect 17454 -55322 17478 -55288
rect 17512 -55322 17536 -55288
rect 17454 -55346 17536 -55322
rect 18472 -55288 18554 -55264
rect 18472 -55322 18496 -55288
rect 18530 -55322 18554 -55288
rect 18472 -55346 18554 -55322
rect 19490 -55288 19572 -55264
rect 19490 -55322 19514 -55288
rect 19548 -55322 19572 -55288
rect 19490 -55346 19572 -55322
rect 20508 -55288 20590 -55264
rect 20508 -55322 20532 -55288
rect 20566 -55322 20590 -55288
rect 20508 -55346 20590 -55322
rect 21526 -55288 21608 -55264
rect 21526 -55322 21550 -55288
rect 21584 -55322 21608 -55288
rect 21526 -55346 21608 -55322
rect 22544 -55288 22626 -55264
rect 22544 -55322 22568 -55288
rect 22602 -55322 22626 -55288
rect 22544 -55346 22626 -55322
rect 23562 -55288 23644 -55264
rect 23562 -55322 23586 -55288
rect 23620 -55322 23644 -55288
rect 23562 -55346 23644 -55322
rect 24580 -55288 24662 -55264
rect 24580 -55322 24604 -55288
rect 24638 -55322 24662 -55288
rect 24580 -55346 24662 -55322
rect 25598 -55288 25680 -55264
rect 25598 -55322 25622 -55288
rect 25656 -55322 25680 -55288
rect 25598 -55346 25680 -55322
rect 28024 -55446 28058 -55430
rect 29042 -54854 29076 -54838
rect 29042 -55446 29076 -55430
rect 30060 -54854 30094 -54838
rect 30060 -55446 30094 -55430
rect 31078 -54854 31112 -54838
rect 31078 -55446 31112 -55430
rect 32096 -54854 32130 -54838
rect 32096 -55446 32130 -55430
rect 33114 -54854 33148 -54838
rect 33114 -55446 33148 -55430
rect 34132 -54854 34166 -54838
rect 34132 -55446 34166 -55430
rect 35150 -54854 35184 -54838
rect 35150 -55446 35184 -55430
rect 36168 -54854 36202 -54838
rect 36168 -55446 36202 -55430
rect 37186 -54854 37220 -54838
rect 37186 -55446 37220 -55430
rect 38204 -54854 38238 -54838
rect 38204 -55446 38238 -55430
rect 39222 -54854 39256 -54838
rect 39222 -55446 39256 -55430
rect 40240 -54854 40274 -54838
rect 40240 -55446 40274 -55430
rect 41258 -54854 41292 -54838
rect 41258 -55446 41292 -55430
rect 42276 -54854 42310 -54838
rect 42276 -55446 42310 -55430
rect 43294 -54854 43328 -54838
rect 43294 -55446 43328 -55430
rect 44312 -54854 44346 -54838
rect 44312 -55446 44346 -55430
rect 45330 -54854 45364 -54838
rect 45330 -55446 45364 -55430
rect 46348 -54854 46382 -54838
rect 46348 -55446 46382 -55430
rect 47366 -54854 47400 -54838
rect 47366 -55446 47400 -55430
rect 48384 -54854 48418 -54838
rect 48384 -55446 48418 -55430
rect 35650 -55480 35710 -55470
rect 15168 -55538 15184 -55504
rect 15740 -55538 15756 -55504
rect 16186 -55538 16202 -55504
rect 16758 -55538 16774 -55504
rect 17204 -55538 17220 -55504
rect 17776 -55538 17792 -55504
rect 18222 -55538 18238 -55504
rect 18794 -55538 18810 -55504
rect 19240 -55538 19256 -55504
rect 19812 -55538 19828 -55504
rect 20258 -55538 20274 -55504
rect 20830 -55538 20846 -55504
rect 21276 -55538 21292 -55504
rect 21848 -55538 21864 -55504
rect 22294 -55538 22310 -55504
rect 22866 -55538 22882 -55504
rect 23312 -55538 23328 -55504
rect 23884 -55538 23900 -55504
rect 24330 -55538 24346 -55504
rect 24902 -55538 24918 -55504
rect 25348 -55538 25364 -55504
rect 25920 -55538 25936 -55504
rect 28256 -55514 28272 -55480
rect 28828 -55514 28844 -55480
rect 29274 -55514 29290 -55480
rect 29846 -55514 29862 -55480
rect 30292 -55514 30308 -55480
rect 30864 -55514 30880 -55480
rect 31310 -55514 31326 -55480
rect 31882 -55514 31898 -55480
rect 32328 -55514 32344 -55480
rect 32900 -55514 32916 -55480
rect 33346 -55514 33362 -55480
rect 33918 -55514 33934 -55480
rect 34364 -55514 34380 -55480
rect 34936 -55514 34952 -55480
rect 35382 -55514 35398 -55480
rect 35954 -55514 35970 -55480
rect 36400 -55514 36416 -55480
rect 36972 -55514 36988 -55480
rect 37418 -55514 37434 -55480
rect 37990 -55514 38006 -55480
rect 38436 -55514 38452 -55480
rect 39008 -55514 39024 -55480
rect 39454 -55514 39470 -55480
rect 40026 -55514 40042 -55480
rect 40472 -55514 40488 -55480
rect 41044 -55514 41060 -55480
rect 41490 -55514 41506 -55480
rect 42062 -55514 42078 -55480
rect 42508 -55514 42524 -55480
rect 43080 -55514 43096 -55480
rect 43526 -55514 43542 -55480
rect 44098 -55514 44114 -55480
rect 44544 -55514 44560 -55480
rect 45116 -55514 45132 -55480
rect 45562 -55514 45578 -55480
rect 46134 -55514 46150 -55480
rect 46580 -55514 46596 -55480
rect 47152 -55514 47168 -55480
rect 47598 -55514 47614 -55480
rect 48170 -55514 48186 -55480
rect 14936 -55588 14970 -55572
rect 14936 -56180 14970 -56164
rect 15954 -55588 15988 -55572
rect 15954 -56180 15988 -56164
rect 16972 -55588 17006 -55572
rect 16972 -56180 17006 -56164
rect 17990 -55588 18024 -55572
rect 17990 -56180 18024 -56164
rect 19008 -55588 19042 -55572
rect 19008 -56180 19042 -56164
rect 20026 -55588 20060 -55572
rect 20026 -56180 20060 -56164
rect 21044 -55588 21078 -55572
rect 21044 -56180 21078 -56164
rect 22062 -55588 22096 -55572
rect 22062 -56180 22096 -56164
rect 23080 -55588 23114 -55572
rect 23080 -56180 23114 -56164
rect 24098 -55588 24132 -55572
rect 24098 -56180 24132 -56164
rect 25116 -55588 25150 -55572
rect 25116 -56180 25150 -56164
rect 26134 -55588 26168 -55572
rect 28518 -55734 28600 -55710
rect 28518 -55768 28542 -55734
rect 28576 -55768 28600 -55734
rect 28518 -55792 28600 -55768
rect 29536 -55734 29618 -55710
rect 29536 -55768 29560 -55734
rect 29594 -55768 29618 -55734
rect 29536 -55792 29618 -55768
rect 30554 -55734 30636 -55710
rect 30554 -55768 30578 -55734
rect 30612 -55768 30636 -55734
rect 30554 -55792 30636 -55768
rect 31572 -55734 31654 -55710
rect 31572 -55768 31596 -55734
rect 31630 -55768 31654 -55734
rect 31572 -55792 31654 -55768
rect 32590 -55734 32672 -55710
rect 32590 -55768 32614 -55734
rect 32648 -55768 32672 -55734
rect 32590 -55792 32672 -55768
rect 33608 -55734 33690 -55710
rect 33608 -55768 33632 -55734
rect 33666 -55768 33690 -55734
rect 33608 -55792 33690 -55768
rect 34626 -55734 34708 -55710
rect 34626 -55768 34650 -55734
rect 34684 -55768 34708 -55734
rect 34626 -55792 34708 -55768
rect 35644 -55734 35726 -55710
rect 35644 -55768 35668 -55734
rect 35702 -55768 35726 -55734
rect 35644 -55792 35726 -55768
rect 36662 -55734 36744 -55710
rect 36662 -55768 36686 -55734
rect 36720 -55768 36744 -55734
rect 36662 -55792 36744 -55768
rect 37680 -55734 37762 -55710
rect 37680 -55768 37704 -55734
rect 37738 -55768 37762 -55734
rect 37680 -55792 37762 -55768
rect 38698 -55734 38780 -55710
rect 38698 -55768 38722 -55734
rect 38756 -55768 38780 -55734
rect 38698 -55792 38780 -55768
rect 39716 -55734 39798 -55710
rect 39716 -55768 39740 -55734
rect 39774 -55768 39798 -55734
rect 39716 -55792 39798 -55768
rect 40734 -55734 40816 -55710
rect 40734 -55768 40758 -55734
rect 40792 -55768 40816 -55734
rect 40734 -55792 40816 -55768
rect 41752 -55734 41834 -55710
rect 41752 -55768 41776 -55734
rect 41810 -55768 41834 -55734
rect 41752 -55792 41834 -55768
rect 42770 -55734 42852 -55710
rect 42770 -55768 42794 -55734
rect 42828 -55768 42852 -55734
rect 42770 -55792 42852 -55768
rect 43788 -55734 43870 -55710
rect 43788 -55768 43812 -55734
rect 43846 -55768 43870 -55734
rect 43788 -55792 43870 -55768
rect 44806 -55734 44888 -55710
rect 44806 -55768 44830 -55734
rect 44864 -55768 44888 -55734
rect 44806 -55792 44888 -55768
rect 45824 -55734 45906 -55710
rect 45824 -55768 45848 -55734
rect 45882 -55768 45906 -55734
rect 45824 -55792 45906 -55768
rect 46842 -55734 46924 -55710
rect 46842 -55768 46866 -55734
rect 46900 -55768 46924 -55734
rect 46842 -55792 46924 -55768
rect 47860 -55734 47942 -55710
rect 47860 -55768 47884 -55734
rect 47918 -55768 47942 -55734
rect 47860 -55792 47942 -55768
rect 28256 -56038 28272 -56004
rect 28828 -56038 28844 -56004
rect 29274 -56038 29290 -56004
rect 29846 -56038 29862 -56004
rect 30292 -56038 30308 -56004
rect 30864 -56038 30880 -56004
rect 31310 -56038 31326 -56004
rect 31882 -56038 31898 -56004
rect 32328 -56038 32344 -56004
rect 32900 -56038 32916 -56004
rect 33346 -56038 33362 -56004
rect 33918 -56038 33934 -56004
rect 34364 -56038 34380 -56004
rect 34936 -56038 34952 -56004
rect 35382 -56038 35398 -56004
rect 35954 -56038 35970 -56004
rect 36400 -56038 36416 -56004
rect 36972 -56038 36988 -56004
rect 37418 -56038 37434 -56004
rect 37990 -56038 38006 -56004
rect 38436 -56038 38452 -56004
rect 39008 -56038 39024 -56004
rect 39454 -56038 39470 -56004
rect 40026 -56038 40042 -56004
rect 40472 -56038 40488 -56004
rect 41044 -56038 41060 -56004
rect 41490 -56038 41506 -56004
rect 42062 -56038 42078 -56004
rect 42508 -56038 42524 -56004
rect 43080 -56038 43096 -56004
rect 43526 -56038 43542 -56004
rect 44098 -56038 44114 -56004
rect 44544 -56038 44560 -56004
rect 45116 -56038 45132 -56004
rect 45562 -56038 45578 -56004
rect 46134 -56038 46150 -56004
rect 46580 -56038 46596 -56004
rect 47152 -56038 47168 -56004
rect 47598 -56038 47614 -56004
rect 48170 -56038 48186 -56004
rect 31564 -56040 31624 -56038
rect 26134 -56180 26168 -56164
rect 28024 -56088 28058 -56072
rect 15168 -56248 15184 -56214
rect 15740 -56248 15756 -56214
rect 16186 -56248 16202 -56214
rect 16758 -56248 16774 -56214
rect 17204 -56248 17220 -56214
rect 17776 -56248 17792 -56214
rect 18222 -56248 18238 -56214
rect 18794 -56248 18810 -56214
rect 19240 -56248 19256 -56214
rect 19812 -56248 19828 -56214
rect 20258 -56248 20274 -56214
rect 20830 -56248 20846 -56214
rect 21276 -56248 21292 -56214
rect 21848 -56248 21864 -56214
rect 22294 -56248 22310 -56214
rect 22866 -56248 22882 -56214
rect 23312 -56248 23328 -56214
rect 23884 -56248 23900 -56214
rect 24330 -56248 24346 -56214
rect 24902 -56248 24918 -56214
rect 25348 -56248 25364 -56214
rect 25920 -56248 25936 -56214
rect 15418 -56630 15500 -56606
rect 15418 -56664 15442 -56630
rect 15476 -56664 15500 -56630
rect 15418 -56688 15500 -56664
rect 16436 -56630 16518 -56606
rect 16436 -56664 16460 -56630
rect 16494 -56664 16518 -56630
rect 16436 -56688 16518 -56664
rect 17454 -56630 17536 -56606
rect 17454 -56664 17478 -56630
rect 17512 -56664 17536 -56630
rect 17454 -56688 17536 -56664
rect 18472 -56630 18554 -56606
rect 18472 -56664 18496 -56630
rect 18530 -56664 18554 -56630
rect 18472 -56688 18554 -56664
rect 19490 -56630 19572 -56606
rect 19490 -56664 19514 -56630
rect 19548 -56664 19572 -56630
rect 19490 -56688 19572 -56664
rect 20508 -56630 20590 -56606
rect 20508 -56664 20532 -56630
rect 20566 -56664 20590 -56630
rect 20508 -56688 20590 -56664
rect 21526 -56630 21608 -56606
rect 21526 -56664 21550 -56630
rect 21584 -56664 21608 -56630
rect 21526 -56688 21608 -56664
rect 22544 -56630 22626 -56606
rect 22544 -56664 22568 -56630
rect 22602 -56664 22626 -56630
rect 22544 -56688 22626 -56664
rect 23562 -56630 23644 -56606
rect 23562 -56664 23586 -56630
rect 23620 -56664 23644 -56630
rect 23562 -56688 23644 -56664
rect 24580 -56630 24662 -56606
rect 24580 -56664 24604 -56630
rect 24638 -56664 24662 -56630
rect 24580 -56688 24662 -56664
rect 25598 -56630 25680 -56606
rect 25598 -56664 25622 -56630
rect 25656 -56664 25680 -56630
rect 25598 -56688 25680 -56664
rect 28024 -56680 28058 -56664
rect 29042 -56088 29076 -56072
rect 29042 -56680 29076 -56664
rect 30060 -56088 30094 -56072
rect 30060 -56680 30094 -56664
rect 31078 -56088 31112 -56072
rect 31078 -56680 31112 -56664
rect 32096 -56088 32130 -56072
rect 32096 -56680 32130 -56664
rect 33114 -56088 33148 -56072
rect 33114 -56680 33148 -56664
rect 34132 -56088 34166 -56072
rect 34132 -56680 34166 -56664
rect 35150 -56088 35184 -56072
rect 35150 -56680 35184 -56664
rect 36168 -56088 36202 -56072
rect 36168 -56680 36202 -56664
rect 37186 -56088 37220 -56072
rect 37186 -56680 37220 -56664
rect 38204 -56088 38238 -56072
rect 38204 -56680 38238 -56664
rect 39222 -56088 39256 -56072
rect 39222 -56680 39256 -56664
rect 40240 -56088 40274 -56072
rect 40240 -56680 40274 -56664
rect 41258 -56088 41292 -56072
rect 41258 -56680 41292 -56664
rect 42276 -56088 42310 -56072
rect 42276 -56680 42310 -56664
rect 43294 -56088 43328 -56072
rect 43294 -56680 43328 -56664
rect 44312 -56088 44346 -56072
rect 44312 -56680 44346 -56664
rect 45330 -56088 45364 -56072
rect 45330 -56680 45364 -56664
rect 46348 -56088 46382 -56072
rect 46348 -56680 46382 -56664
rect 47366 -56088 47400 -56072
rect 47366 -56680 47400 -56664
rect 48384 -56088 48418 -56072
rect 48384 -56680 48418 -56664
rect 29532 -56714 29592 -56712
rect 35644 -56714 35704 -56712
rect 37678 -56714 37738 -56712
rect 41744 -56714 41804 -56708
rect 45820 -56714 45880 -56712
rect 46836 -56714 46896 -56712
rect 28256 -56748 28272 -56714
rect 28828 -56748 28844 -56714
rect 29274 -56748 29290 -56714
rect 29846 -56748 29862 -56714
rect 30292 -56748 30308 -56714
rect 30864 -56748 30880 -56714
rect 31310 -56748 31326 -56714
rect 31882 -56748 31898 -56714
rect 32328 -56748 32344 -56714
rect 32900 -56748 32916 -56714
rect 33346 -56748 33362 -56714
rect 33918 -56748 33934 -56714
rect 34364 -56748 34380 -56714
rect 34936 -56748 34952 -56714
rect 35382 -56748 35398 -56714
rect 35954 -56748 35970 -56714
rect 36400 -56748 36416 -56714
rect 36972 -56748 36988 -56714
rect 37418 -56748 37434 -56714
rect 37990 -56748 38006 -56714
rect 38436 -56748 38452 -56714
rect 39008 -56748 39024 -56714
rect 39454 -56748 39470 -56714
rect 40026 -56748 40042 -56714
rect 40472 -56748 40488 -56714
rect 41044 -56748 41060 -56714
rect 41490 -56748 41506 -56714
rect 42062 -56748 42078 -56714
rect 42508 -56748 42524 -56714
rect 43080 -56748 43096 -56714
rect 43526 -56748 43542 -56714
rect 44098 -56748 44114 -56714
rect 44544 -56748 44560 -56714
rect 45116 -56748 45132 -56714
rect 45562 -56748 45578 -56714
rect 46134 -56748 46150 -56714
rect 46580 -56748 46596 -56714
rect 47152 -56748 47168 -56714
rect 47598 -56748 47614 -56714
rect 48170 -56748 48186 -56714
rect 28530 -56980 28612 -56956
rect 28530 -57014 28554 -56980
rect 28588 -57014 28612 -56980
rect 28530 -57038 28612 -57014
rect 29548 -56980 29630 -56956
rect 29548 -57014 29572 -56980
rect 29606 -57014 29630 -56980
rect 29548 -57038 29630 -57014
rect 30566 -56980 30648 -56956
rect 30566 -57014 30590 -56980
rect 30624 -57014 30648 -56980
rect 30566 -57038 30648 -57014
rect 31584 -56980 31666 -56956
rect 31584 -57014 31608 -56980
rect 31642 -57014 31666 -56980
rect 31584 -57038 31666 -57014
rect 32602 -56980 32684 -56956
rect 32602 -57014 32626 -56980
rect 32660 -57014 32684 -56980
rect 32602 -57038 32684 -57014
rect 33620 -56980 33702 -56956
rect 33620 -57014 33644 -56980
rect 33678 -57014 33702 -56980
rect 33620 -57038 33702 -57014
rect 34638 -56980 34720 -56956
rect 34638 -57014 34662 -56980
rect 34696 -57014 34720 -56980
rect 34638 -57038 34720 -57014
rect 35656 -56980 35738 -56956
rect 35656 -57014 35680 -56980
rect 35714 -57014 35738 -56980
rect 35656 -57038 35738 -57014
rect 36674 -56980 36756 -56956
rect 36674 -57014 36698 -56980
rect 36732 -57014 36756 -56980
rect 36674 -57038 36756 -57014
rect 37692 -56980 37774 -56956
rect 37692 -57014 37716 -56980
rect 37750 -57014 37774 -56980
rect 37692 -57038 37774 -57014
rect 38710 -56980 38792 -56956
rect 38710 -57014 38734 -56980
rect 38768 -57014 38792 -56980
rect 38710 -57038 38792 -57014
rect 39728 -56980 39810 -56956
rect 39728 -57014 39752 -56980
rect 39786 -57014 39810 -56980
rect 39728 -57038 39810 -57014
rect 40746 -56980 40828 -56956
rect 40746 -57014 40770 -56980
rect 40804 -57014 40828 -56980
rect 40746 -57038 40828 -57014
rect 41764 -56980 41846 -56956
rect 41764 -57014 41788 -56980
rect 41822 -57014 41846 -56980
rect 41764 -57038 41846 -57014
rect 42782 -56980 42864 -56956
rect 42782 -57014 42806 -56980
rect 42840 -57014 42864 -56980
rect 42782 -57038 42864 -57014
rect 43800 -56980 43882 -56956
rect 43800 -57014 43824 -56980
rect 43858 -57014 43882 -56980
rect 43800 -57038 43882 -57014
rect 44818 -56980 44900 -56956
rect 44818 -57014 44842 -56980
rect 44876 -57014 44900 -56980
rect 44818 -57038 44900 -57014
rect 45836 -56980 45918 -56956
rect 45836 -57014 45860 -56980
rect 45894 -57014 45918 -56980
rect 45836 -57038 45918 -57014
rect 46854 -56980 46936 -56956
rect 46854 -57014 46878 -56980
rect 46912 -57014 46936 -56980
rect 46854 -57038 46936 -57014
rect 47872 -56980 47954 -56956
rect 47872 -57014 47896 -56980
rect 47930 -57014 47954 -56980
rect 47872 -57038 47954 -57014
rect 15626 -57080 15642 -57046
rect 16198 -57080 16214 -57046
rect 16644 -57080 16660 -57046
rect 17216 -57080 17232 -57046
rect 17662 -57080 17678 -57046
rect 18234 -57080 18250 -57046
rect 18680 -57080 18696 -57046
rect 19252 -57080 19268 -57046
rect 19698 -57080 19714 -57046
rect 20270 -57080 20286 -57046
rect 20716 -57080 20732 -57046
rect 21288 -57080 21304 -57046
rect 21734 -57080 21750 -57046
rect 22306 -57080 22322 -57046
rect 22752 -57080 22768 -57046
rect 23324 -57080 23340 -57046
rect 23770 -57080 23786 -57046
rect 24342 -57080 24358 -57046
rect 24788 -57080 24804 -57046
rect 25360 -57080 25376 -57046
rect 15394 -57130 15428 -57114
rect 15394 -57722 15428 -57706
rect 16412 -57130 16446 -57114
rect 16412 -57722 16446 -57706
rect 17430 -57130 17464 -57114
rect 17430 -57722 17464 -57706
rect 18448 -57130 18482 -57114
rect 18448 -57722 18482 -57706
rect 19466 -57130 19500 -57114
rect 19466 -57722 19500 -57706
rect 20484 -57130 20518 -57114
rect 20484 -57722 20518 -57706
rect 21502 -57130 21536 -57114
rect 21502 -57722 21536 -57706
rect 22520 -57130 22554 -57114
rect 22520 -57722 22554 -57706
rect 23538 -57130 23572 -57114
rect 23538 -57722 23572 -57706
rect 24556 -57130 24590 -57114
rect 24556 -57722 24590 -57706
rect 25574 -57130 25608 -57114
rect 28256 -57270 28272 -57236
rect 28828 -57270 28844 -57236
rect 29274 -57270 29290 -57236
rect 29846 -57270 29862 -57236
rect 30292 -57270 30308 -57236
rect 30864 -57270 30880 -57236
rect 31310 -57270 31326 -57236
rect 31882 -57270 31898 -57236
rect 32328 -57270 32344 -57236
rect 32900 -57270 32916 -57236
rect 33346 -57270 33362 -57236
rect 33918 -57270 33934 -57236
rect 34364 -57270 34380 -57236
rect 34936 -57270 34952 -57236
rect 35382 -57270 35398 -57236
rect 35954 -57270 35970 -57236
rect 36400 -57270 36416 -57236
rect 36972 -57270 36988 -57236
rect 37418 -57270 37434 -57236
rect 37990 -57270 38006 -57236
rect 38436 -57270 38452 -57236
rect 39008 -57270 39024 -57236
rect 39454 -57270 39470 -57236
rect 40026 -57270 40042 -57236
rect 40472 -57270 40488 -57236
rect 41044 -57270 41060 -57236
rect 41490 -57270 41506 -57236
rect 42062 -57270 42078 -57236
rect 42508 -57270 42524 -57236
rect 43080 -57270 43096 -57236
rect 43526 -57270 43542 -57236
rect 44098 -57270 44114 -57236
rect 44544 -57270 44560 -57236
rect 45116 -57270 45132 -57236
rect 45562 -57270 45578 -57236
rect 46134 -57270 46150 -57236
rect 46580 -57270 46596 -57236
rect 47152 -57270 47168 -57236
rect 47598 -57270 47614 -57236
rect 48170 -57270 48186 -57236
rect 25574 -57722 25608 -57706
rect 28024 -57320 28058 -57304
rect 15626 -57790 15642 -57756
rect 16198 -57790 16214 -57756
rect 16644 -57790 16660 -57756
rect 17216 -57790 17232 -57756
rect 17662 -57790 17678 -57756
rect 18234 -57790 18250 -57756
rect 18680 -57790 18696 -57756
rect 19252 -57790 19268 -57756
rect 19698 -57790 19714 -57756
rect 20270 -57790 20286 -57756
rect 20716 -57790 20732 -57756
rect 21288 -57790 21304 -57756
rect 21734 -57790 21750 -57756
rect 22306 -57790 22322 -57756
rect 22752 -57790 22768 -57756
rect 23324 -57790 23340 -57756
rect 23770 -57790 23786 -57756
rect 24342 -57790 24358 -57756
rect 24788 -57790 24804 -57756
rect 25360 -57790 25376 -57756
rect 28024 -57912 28058 -57896
rect 29042 -57320 29076 -57304
rect 29042 -57912 29076 -57896
rect 30060 -57320 30094 -57304
rect 30060 -57912 30094 -57896
rect 31078 -57320 31112 -57304
rect 31078 -57912 31112 -57896
rect 32096 -57320 32130 -57304
rect 32096 -57912 32130 -57896
rect 33114 -57320 33148 -57304
rect 33114 -57912 33148 -57896
rect 34132 -57320 34166 -57304
rect 34132 -57912 34166 -57896
rect 35150 -57320 35184 -57304
rect 35150 -57912 35184 -57896
rect 36168 -57320 36202 -57304
rect 36168 -57912 36202 -57896
rect 37186 -57320 37220 -57304
rect 37186 -57912 37220 -57896
rect 38204 -57320 38238 -57304
rect 38204 -57912 38238 -57896
rect 39222 -57320 39256 -57304
rect 39222 -57912 39256 -57896
rect 40240 -57320 40274 -57304
rect 40240 -57912 40274 -57896
rect 41258 -57320 41292 -57304
rect 41258 -57912 41292 -57896
rect 42276 -57320 42310 -57304
rect 42276 -57912 42310 -57896
rect 43294 -57320 43328 -57304
rect 43294 -57912 43328 -57896
rect 44312 -57320 44346 -57304
rect 44312 -57912 44346 -57896
rect 45330 -57320 45364 -57304
rect 45330 -57912 45364 -57896
rect 46348 -57320 46382 -57304
rect 46348 -57912 46382 -57896
rect 47366 -57320 47400 -57304
rect 47366 -57912 47400 -57896
rect 48384 -57320 48418 -57304
rect 48384 -57912 48418 -57896
rect 28256 -57980 28272 -57946
rect 28828 -57980 28844 -57946
rect 29274 -57980 29290 -57946
rect 29846 -57980 29862 -57946
rect 30292 -57980 30308 -57946
rect 30864 -57980 30880 -57946
rect 31310 -57980 31326 -57946
rect 31882 -57980 31898 -57946
rect 32328 -57980 32344 -57946
rect 32900 -57980 32916 -57946
rect 33346 -57980 33362 -57946
rect 33918 -57980 33934 -57946
rect 34364 -57980 34380 -57946
rect 34936 -57980 34952 -57946
rect 35382 -57980 35398 -57946
rect 35954 -57980 35970 -57946
rect 36400 -57980 36416 -57946
rect 36972 -57980 36988 -57946
rect 37418 -57980 37434 -57946
rect 37990 -57980 38006 -57946
rect 38436 -57980 38452 -57946
rect 39008 -57980 39024 -57946
rect 39454 -57980 39470 -57946
rect 40026 -57980 40042 -57946
rect 40472 -57980 40488 -57946
rect 41044 -57980 41060 -57946
rect 41490 -57980 41506 -57946
rect 42062 -57980 42078 -57946
rect 42508 -57980 42524 -57946
rect 43080 -57980 43096 -57946
rect 43526 -57980 43542 -57946
rect 44098 -57980 44114 -57946
rect 44544 -57980 44560 -57946
rect 45116 -57980 45132 -57946
rect 45562 -57980 45578 -57946
rect 46134 -57980 46150 -57946
rect 46580 -57980 46596 -57946
rect 47152 -57980 47168 -57946
rect 47598 -57980 47614 -57946
rect 48170 -57980 48186 -57946
rect 15228 -58076 15310 -58052
rect 15228 -58110 15252 -58076
rect 15286 -58110 15310 -58076
rect 15228 -58134 15310 -58110
rect 16246 -58076 16328 -58052
rect 16246 -58110 16270 -58076
rect 16304 -58110 16328 -58076
rect 16246 -58134 16328 -58110
rect 17264 -58076 17346 -58052
rect 17264 -58110 17288 -58076
rect 17322 -58110 17346 -58076
rect 17264 -58134 17346 -58110
rect 18282 -58076 18364 -58052
rect 18282 -58110 18306 -58076
rect 18340 -58110 18364 -58076
rect 18282 -58134 18364 -58110
rect 19300 -58076 19382 -58052
rect 19300 -58110 19324 -58076
rect 19358 -58110 19382 -58076
rect 19300 -58134 19382 -58110
rect 20318 -58076 20400 -58052
rect 20318 -58110 20342 -58076
rect 20376 -58110 20400 -58076
rect 20318 -58134 20400 -58110
rect 21336 -58076 21418 -58052
rect 21336 -58110 21360 -58076
rect 21394 -58110 21418 -58076
rect 21336 -58134 21418 -58110
rect 22354 -58076 22436 -58052
rect 22354 -58110 22378 -58076
rect 22412 -58110 22436 -58076
rect 22354 -58134 22436 -58110
rect 23372 -58076 23454 -58052
rect 23372 -58110 23396 -58076
rect 23430 -58110 23454 -58076
rect 23372 -58134 23454 -58110
rect 24390 -58076 24472 -58052
rect 24390 -58110 24414 -58076
rect 24448 -58110 24472 -58076
rect 24390 -58134 24472 -58110
rect 25408 -58076 25490 -58052
rect 25408 -58110 25432 -58076
rect 25466 -58110 25490 -58076
rect 25408 -58134 25490 -58110
rect 28518 -58158 28600 -58134
rect 28518 -58192 28542 -58158
rect 28576 -58192 28600 -58158
rect 28518 -58216 28600 -58192
rect 29536 -58158 29618 -58134
rect 29536 -58192 29560 -58158
rect 29594 -58192 29618 -58158
rect 29536 -58216 29618 -58192
rect 30554 -58158 30636 -58134
rect 30554 -58192 30578 -58158
rect 30612 -58192 30636 -58158
rect 30554 -58216 30636 -58192
rect 31572 -58158 31654 -58134
rect 31572 -58192 31596 -58158
rect 31630 -58192 31654 -58158
rect 31572 -58216 31654 -58192
rect 32590 -58158 32672 -58134
rect 32590 -58192 32614 -58158
rect 32648 -58192 32672 -58158
rect 32590 -58216 32672 -58192
rect 33608 -58158 33690 -58134
rect 33608 -58192 33632 -58158
rect 33666 -58192 33690 -58158
rect 33608 -58216 33690 -58192
rect 34626 -58158 34708 -58134
rect 34626 -58192 34650 -58158
rect 34684 -58192 34708 -58158
rect 34626 -58216 34708 -58192
rect 35644 -58158 35726 -58134
rect 35644 -58192 35668 -58158
rect 35702 -58192 35726 -58158
rect 35644 -58216 35726 -58192
rect 36662 -58158 36744 -58134
rect 36662 -58192 36686 -58158
rect 36720 -58192 36744 -58158
rect 36662 -58216 36744 -58192
rect 37680 -58158 37762 -58134
rect 37680 -58192 37704 -58158
rect 37738 -58192 37762 -58158
rect 37680 -58216 37762 -58192
rect 38698 -58158 38780 -58134
rect 38698 -58192 38722 -58158
rect 38756 -58192 38780 -58158
rect 38698 -58216 38780 -58192
rect 39716 -58158 39798 -58134
rect 39716 -58192 39740 -58158
rect 39774 -58192 39798 -58158
rect 39716 -58216 39798 -58192
rect 40734 -58158 40816 -58134
rect 40734 -58192 40758 -58158
rect 40792 -58192 40816 -58158
rect 40734 -58216 40816 -58192
rect 41752 -58158 41834 -58134
rect 41752 -58192 41776 -58158
rect 41810 -58192 41834 -58158
rect 41752 -58216 41834 -58192
rect 42770 -58158 42852 -58134
rect 42770 -58192 42794 -58158
rect 42828 -58192 42852 -58158
rect 42770 -58216 42852 -58192
rect 43788 -58158 43870 -58134
rect 43788 -58192 43812 -58158
rect 43846 -58192 43870 -58158
rect 43788 -58216 43870 -58192
rect 44806 -58158 44888 -58134
rect 44806 -58192 44830 -58158
rect 44864 -58192 44888 -58158
rect 44806 -58216 44888 -58192
rect 45824 -58158 45906 -58134
rect 45824 -58192 45848 -58158
rect 45882 -58192 45906 -58158
rect 45824 -58216 45906 -58192
rect 46842 -58158 46924 -58134
rect 46842 -58192 46866 -58158
rect 46900 -58192 46924 -58158
rect 46842 -58216 46924 -58192
rect 47860 -58158 47942 -58134
rect 47860 -58192 47884 -58158
rect 47918 -58192 47942 -58158
rect 47860 -58216 47942 -58192
rect 13122 -59200 13222 -59038
rect 50266 -59200 50366 -59038
rect -27684 -64588 -27584 -64426
rect -28072 -67299 -28043 -67265
rect -28009 -67299 -27951 -67265
rect -27917 -67299 -27859 -67265
rect -27825 -67299 -27796 -67265
rect -25460 -64588 -25360 -64426
rect -27257 -65578 -27241 -65544
rect -27141 -65578 -27125 -65544
rect -26999 -65578 -26983 -65544
rect -26883 -65578 -26867 -65544
rect -26741 -65578 -26725 -65544
rect -26625 -65578 -26609 -65544
rect -26483 -65578 -26467 -65544
rect -26367 -65578 -26351 -65544
rect -26225 -65578 -26209 -65544
rect -26109 -65578 -26093 -65544
rect -25967 -65578 -25951 -65544
rect -25851 -65578 -25835 -65544
rect -27337 -65637 -27303 -65621
rect -27337 -66029 -27303 -66013
rect -27079 -65637 -27045 -65621
rect -27079 -66029 -27045 -66013
rect -26821 -65637 -26787 -65621
rect -26821 -66029 -26787 -66013
rect -26563 -65637 -26529 -65621
rect -26563 -66029 -26529 -66013
rect -26305 -65637 -26271 -65621
rect -26305 -66029 -26271 -66013
rect -26047 -65637 -26013 -65621
rect -26047 -66029 -26013 -66013
rect -25789 -65637 -25755 -65621
rect -25789 -66029 -25755 -66013
rect -27257 -66106 -27241 -66072
rect -27141 -66106 -27125 -66072
rect -26999 -66106 -26983 -66072
rect -26883 -66106 -26867 -66072
rect -26741 -66106 -26725 -66072
rect -26625 -66106 -26609 -66072
rect -26483 -66106 -26467 -66072
rect -26367 -66106 -26351 -66072
rect -26225 -66106 -26209 -66072
rect -26109 -66106 -26093 -66072
rect -25967 -66106 -25951 -66072
rect -25851 -66106 -25835 -66072
rect -27257 -66438 -27241 -66404
rect -27141 -66438 -27125 -66404
rect -26999 -66438 -26983 -66404
rect -26883 -66438 -26867 -66404
rect -26741 -66438 -26725 -66404
rect -26625 -66438 -26609 -66404
rect -26483 -66438 -26467 -66404
rect -26367 -66438 -26351 -66404
rect -26225 -66438 -26209 -66404
rect -26109 -66438 -26093 -66404
rect -25967 -66438 -25951 -66404
rect -25851 -66438 -25835 -66404
rect -27337 -66497 -27303 -66481
rect -27337 -66889 -27303 -66873
rect -27079 -66497 -27045 -66481
rect -27079 -66889 -27045 -66873
rect -26821 -66497 -26787 -66481
rect -26821 -66889 -26787 -66873
rect -26563 -66497 -26529 -66481
rect -26563 -66889 -26529 -66873
rect -26305 -66497 -26271 -66481
rect -26305 -66889 -26271 -66873
rect -26047 -66497 -26013 -66481
rect -26047 -66889 -26013 -66873
rect -25789 -66497 -25755 -66481
rect -25789 -66889 -25755 -66873
rect -27257 -66966 -27241 -66932
rect -27141 -66966 -27125 -66932
rect -26999 -66966 -26983 -66932
rect -26883 -66966 -26867 -66932
rect -26741 -66966 -26725 -66932
rect -26625 -66966 -26609 -66932
rect -26483 -66966 -26467 -66932
rect -26367 -66966 -26351 -66932
rect -26225 -66966 -26209 -66932
rect -26109 -66966 -26093 -66932
rect -25967 -66966 -25951 -66932
rect -25851 -66966 -25835 -66932
rect -28004 -67341 -27962 -67299
rect -28004 -67375 -27996 -67341
rect -28004 -67409 -27962 -67375
rect -28004 -67443 -27996 -67409
rect -28004 -67477 -27962 -67443
rect -28004 -67511 -27996 -67477
rect -28004 -67527 -27962 -67511
rect -27928 -67341 -27862 -67333
rect -27928 -67375 -27912 -67341
rect -27878 -67375 -27862 -67341
rect -27928 -67409 -27862 -67375
rect -27928 -67443 -27912 -67409
rect -27878 -67443 -27862 -67409
rect -27928 -67477 -27862 -67443
rect -27928 -67511 -27912 -67477
rect -27878 -67511 -27862 -67477
rect -27928 -67529 -27862 -67511
rect -28008 -67610 -28004 -67563
rect -27956 -67610 -27942 -67563
rect -28008 -67611 -27992 -67610
rect -27958 -67611 -27942 -67610
rect -27908 -67620 -27862 -67529
rect -27684 -67530 -27584 -67368
rect -23684 -64588 -23584 -64426
rect -24072 -67299 -24043 -67265
rect -24009 -67299 -23951 -67265
rect -23917 -67299 -23859 -67265
rect -23825 -67299 -23796 -67265
rect -21460 -64588 -21360 -64426
rect -23257 -65578 -23241 -65544
rect -23141 -65578 -23125 -65544
rect -22999 -65578 -22983 -65544
rect -22883 -65578 -22867 -65544
rect -22741 -65578 -22725 -65544
rect -22625 -65578 -22609 -65544
rect -22483 -65578 -22467 -65544
rect -22367 -65578 -22351 -65544
rect -22225 -65578 -22209 -65544
rect -22109 -65578 -22093 -65544
rect -21967 -65578 -21951 -65544
rect -21851 -65578 -21835 -65544
rect -23337 -65637 -23303 -65621
rect -23337 -66029 -23303 -66013
rect -23079 -65637 -23045 -65621
rect -23079 -66029 -23045 -66013
rect -22821 -65637 -22787 -65621
rect -22821 -66029 -22787 -66013
rect -22563 -65637 -22529 -65621
rect -22563 -66029 -22529 -66013
rect -22305 -65637 -22271 -65621
rect -22305 -66029 -22271 -66013
rect -22047 -65637 -22013 -65621
rect -22047 -66029 -22013 -66013
rect -21789 -65637 -21755 -65621
rect -21789 -66029 -21755 -66013
rect -23257 -66106 -23241 -66072
rect -23141 -66106 -23125 -66072
rect -22999 -66106 -22983 -66072
rect -22883 -66106 -22867 -66072
rect -22741 -66106 -22725 -66072
rect -22625 -66106 -22609 -66072
rect -22483 -66106 -22467 -66072
rect -22367 -66106 -22351 -66072
rect -22225 -66106 -22209 -66072
rect -22109 -66106 -22093 -66072
rect -21967 -66106 -21951 -66072
rect -21851 -66106 -21835 -66072
rect -23257 -66438 -23241 -66404
rect -23141 -66438 -23125 -66404
rect -22999 -66438 -22983 -66404
rect -22883 -66438 -22867 -66404
rect -22741 -66438 -22725 -66404
rect -22625 -66438 -22609 -66404
rect -22483 -66438 -22467 -66404
rect -22367 -66438 -22351 -66404
rect -22225 -66438 -22209 -66404
rect -22109 -66438 -22093 -66404
rect -21967 -66438 -21951 -66404
rect -21851 -66438 -21835 -66404
rect -23337 -66497 -23303 -66481
rect -23337 -66889 -23303 -66873
rect -23079 -66497 -23045 -66481
rect -23079 -66889 -23045 -66873
rect -22821 -66497 -22787 -66481
rect -22821 -66889 -22787 -66873
rect -22563 -66497 -22529 -66481
rect -22563 -66889 -22529 -66873
rect -22305 -66497 -22271 -66481
rect -22305 -66889 -22271 -66873
rect -22047 -66497 -22013 -66481
rect -22047 -66889 -22013 -66873
rect -21789 -66497 -21755 -66481
rect -21789 -66889 -21755 -66873
rect -23257 -66966 -23241 -66932
rect -23141 -66966 -23125 -66932
rect -22999 -66966 -22983 -66932
rect -22883 -66966 -22867 -66932
rect -22741 -66966 -22725 -66932
rect -22625 -66966 -22609 -66932
rect -22483 -66966 -22467 -66932
rect -22367 -66966 -22351 -66932
rect -22225 -66966 -22209 -66932
rect -22109 -66966 -22093 -66932
rect -21967 -66966 -21951 -66932
rect -21851 -66966 -21835 -66932
rect -25460 -67530 -25360 -67368
rect -24004 -67341 -23962 -67299
rect -24004 -67375 -23996 -67341
rect -24004 -67409 -23962 -67375
rect -24004 -67443 -23996 -67409
rect -24004 -67477 -23962 -67443
rect -24004 -67511 -23996 -67477
rect -24004 -67527 -23962 -67511
rect -23928 -67341 -23862 -67333
rect -23928 -67375 -23912 -67341
rect -23878 -67375 -23862 -67341
rect -23928 -67409 -23862 -67375
rect -23928 -67443 -23912 -67409
rect -23878 -67443 -23862 -67409
rect -23928 -67477 -23862 -67443
rect -23928 -67511 -23912 -67477
rect -23878 -67511 -23862 -67477
rect -23928 -67529 -23862 -67511
rect -24008 -67610 -24004 -67563
rect -23956 -67610 -23942 -67563
rect -24008 -67611 -23992 -67610
rect -23958 -67611 -23942 -67610
rect -23908 -67620 -23862 -67529
rect -23684 -67530 -23584 -67368
rect -19684 -64588 -19584 -64426
rect -20072 -67299 -20043 -67265
rect -20009 -67299 -19951 -67265
rect -19917 -67299 -19859 -67265
rect -19825 -67299 -19796 -67265
rect -17460 -64588 -17360 -64426
rect -19257 -65578 -19241 -65544
rect -19141 -65578 -19125 -65544
rect -18999 -65578 -18983 -65544
rect -18883 -65578 -18867 -65544
rect -18741 -65578 -18725 -65544
rect -18625 -65578 -18609 -65544
rect -18483 -65578 -18467 -65544
rect -18367 -65578 -18351 -65544
rect -18225 -65578 -18209 -65544
rect -18109 -65578 -18093 -65544
rect -17967 -65578 -17951 -65544
rect -17851 -65578 -17835 -65544
rect -19337 -65637 -19303 -65621
rect -19337 -66029 -19303 -66013
rect -19079 -65637 -19045 -65621
rect -19079 -66029 -19045 -66013
rect -18821 -65637 -18787 -65621
rect -18821 -66029 -18787 -66013
rect -18563 -65637 -18529 -65621
rect -18563 -66029 -18529 -66013
rect -18305 -65637 -18271 -65621
rect -18305 -66029 -18271 -66013
rect -18047 -65637 -18013 -65621
rect -18047 -66029 -18013 -66013
rect -17789 -65637 -17755 -65621
rect -17789 -66029 -17755 -66013
rect -19257 -66106 -19241 -66072
rect -19141 -66106 -19125 -66072
rect -18999 -66106 -18983 -66072
rect -18883 -66106 -18867 -66072
rect -18741 -66106 -18725 -66072
rect -18625 -66106 -18609 -66072
rect -18483 -66106 -18467 -66072
rect -18367 -66106 -18351 -66072
rect -18225 -66106 -18209 -66072
rect -18109 -66106 -18093 -66072
rect -17967 -66106 -17951 -66072
rect -17851 -66106 -17835 -66072
rect -19257 -66438 -19241 -66404
rect -19141 -66438 -19125 -66404
rect -18999 -66438 -18983 -66404
rect -18883 -66438 -18867 -66404
rect -18741 -66438 -18725 -66404
rect -18625 -66438 -18609 -66404
rect -18483 -66438 -18467 -66404
rect -18367 -66438 -18351 -66404
rect -18225 -66438 -18209 -66404
rect -18109 -66438 -18093 -66404
rect -17967 -66438 -17951 -66404
rect -17851 -66438 -17835 -66404
rect -19337 -66497 -19303 -66481
rect -19337 -66889 -19303 -66873
rect -19079 -66497 -19045 -66481
rect -19079 -66889 -19045 -66873
rect -18821 -66497 -18787 -66481
rect -18821 -66889 -18787 -66873
rect -18563 -66497 -18529 -66481
rect -18563 -66889 -18529 -66873
rect -18305 -66497 -18271 -66481
rect -18305 -66889 -18271 -66873
rect -18047 -66497 -18013 -66481
rect -18047 -66889 -18013 -66873
rect -17789 -66497 -17755 -66481
rect -17789 -66889 -17755 -66873
rect -19257 -66966 -19241 -66932
rect -19141 -66966 -19125 -66932
rect -18999 -66966 -18983 -66932
rect -18883 -66966 -18867 -66932
rect -18741 -66966 -18725 -66932
rect -18625 -66966 -18609 -66932
rect -18483 -66966 -18467 -66932
rect -18367 -66966 -18351 -66932
rect -18225 -66966 -18209 -66932
rect -18109 -66966 -18093 -66932
rect -17967 -66966 -17951 -66932
rect -17851 -66966 -17835 -66932
rect -21460 -67530 -21360 -67368
rect -20004 -67341 -19962 -67299
rect -20004 -67375 -19996 -67341
rect -20004 -67409 -19962 -67375
rect -20004 -67443 -19996 -67409
rect -20004 -67477 -19962 -67443
rect -20004 -67511 -19996 -67477
rect -20004 -67527 -19962 -67511
rect -19928 -67341 -19862 -67333
rect -19928 -67375 -19912 -67341
rect -19878 -67375 -19862 -67341
rect -19928 -67409 -19862 -67375
rect -19928 -67443 -19912 -67409
rect -19878 -67443 -19862 -67409
rect -19928 -67477 -19862 -67443
rect -19928 -67511 -19912 -67477
rect -19878 -67511 -19862 -67477
rect -19928 -67529 -19862 -67511
rect -20008 -67610 -20004 -67563
rect -19956 -67610 -19942 -67563
rect -20008 -67611 -19992 -67610
rect -19958 -67611 -19942 -67610
rect -19908 -67620 -19862 -67529
rect -19684 -67530 -19584 -67368
rect -15684 -64588 -15584 -64426
rect -16072 -67299 -16043 -67265
rect -16009 -67299 -15951 -67265
rect -15917 -67299 -15859 -67265
rect -15825 -67299 -15796 -67265
rect -13460 -64588 -13360 -64426
rect -15257 -65578 -15241 -65544
rect -15141 -65578 -15125 -65544
rect -14999 -65578 -14983 -65544
rect -14883 -65578 -14867 -65544
rect -14741 -65578 -14725 -65544
rect -14625 -65578 -14609 -65544
rect -14483 -65578 -14467 -65544
rect -14367 -65578 -14351 -65544
rect -14225 -65578 -14209 -65544
rect -14109 -65578 -14093 -65544
rect -13967 -65578 -13951 -65544
rect -13851 -65578 -13835 -65544
rect -15337 -65637 -15303 -65621
rect -15337 -66029 -15303 -66013
rect -15079 -65637 -15045 -65621
rect -15079 -66029 -15045 -66013
rect -14821 -65637 -14787 -65621
rect -14821 -66029 -14787 -66013
rect -14563 -65637 -14529 -65621
rect -14563 -66029 -14529 -66013
rect -14305 -65637 -14271 -65621
rect -14305 -66029 -14271 -66013
rect -14047 -65637 -14013 -65621
rect -14047 -66029 -14013 -66013
rect -13789 -65637 -13755 -65621
rect -13789 -66029 -13755 -66013
rect -15257 -66106 -15241 -66072
rect -15141 -66106 -15125 -66072
rect -14999 -66106 -14983 -66072
rect -14883 -66106 -14867 -66072
rect -14741 -66106 -14725 -66072
rect -14625 -66106 -14609 -66072
rect -14483 -66106 -14467 -66072
rect -14367 -66106 -14351 -66072
rect -14225 -66106 -14209 -66072
rect -14109 -66106 -14093 -66072
rect -13967 -66106 -13951 -66072
rect -13851 -66106 -13835 -66072
rect -15257 -66438 -15241 -66404
rect -15141 -66438 -15125 -66404
rect -14999 -66438 -14983 -66404
rect -14883 -66438 -14867 -66404
rect -14741 -66438 -14725 -66404
rect -14625 -66438 -14609 -66404
rect -14483 -66438 -14467 -66404
rect -14367 -66438 -14351 -66404
rect -14225 -66438 -14209 -66404
rect -14109 -66438 -14093 -66404
rect -13967 -66438 -13951 -66404
rect -13851 -66438 -13835 -66404
rect -15337 -66497 -15303 -66481
rect -15337 -66889 -15303 -66873
rect -15079 -66497 -15045 -66481
rect -15079 -66889 -15045 -66873
rect -14821 -66497 -14787 -66481
rect -14821 -66889 -14787 -66873
rect -14563 -66497 -14529 -66481
rect -14563 -66889 -14529 -66873
rect -14305 -66497 -14271 -66481
rect -14305 -66889 -14271 -66873
rect -14047 -66497 -14013 -66481
rect -14047 -66889 -14013 -66873
rect -13789 -66497 -13755 -66481
rect -13789 -66889 -13755 -66873
rect -15257 -66966 -15241 -66932
rect -15141 -66966 -15125 -66932
rect -14999 -66966 -14983 -66932
rect -14883 -66966 -14867 -66932
rect -14741 -66966 -14725 -66932
rect -14625 -66966 -14609 -66932
rect -14483 -66966 -14467 -66932
rect -14367 -66966 -14351 -66932
rect -14225 -66966 -14209 -66932
rect -14109 -66966 -14093 -66932
rect -13967 -66966 -13951 -66932
rect -13851 -66966 -13835 -66932
rect -17460 -67530 -17360 -67368
rect -16004 -67341 -15962 -67299
rect -16004 -67375 -15996 -67341
rect -16004 -67409 -15962 -67375
rect -16004 -67443 -15996 -67409
rect -16004 -67477 -15962 -67443
rect -16004 -67511 -15996 -67477
rect -16004 -67527 -15962 -67511
rect -15928 -67341 -15862 -67333
rect -15928 -67375 -15912 -67341
rect -15878 -67375 -15862 -67341
rect -15928 -67409 -15862 -67375
rect -15928 -67443 -15912 -67409
rect -15878 -67443 -15862 -67409
rect -15928 -67477 -15862 -67443
rect -15928 -67511 -15912 -67477
rect -15878 -67511 -15862 -67477
rect -15928 -67529 -15862 -67511
rect -16008 -67610 -16004 -67563
rect -15956 -67610 -15942 -67563
rect -16008 -67611 -15992 -67610
rect -15958 -67611 -15942 -67610
rect -15908 -67620 -15862 -67529
rect -15684 -67530 -15584 -67368
rect -11684 -64588 -11584 -64426
rect -12072 -67299 -12043 -67265
rect -12009 -67299 -11951 -67265
rect -11917 -67299 -11859 -67265
rect -11825 -67299 -11796 -67265
rect -9460 -64588 -9360 -64426
rect -11257 -65578 -11241 -65544
rect -11141 -65578 -11125 -65544
rect -10999 -65578 -10983 -65544
rect -10883 -65578 -10867 -65544
rect -10741 -65578 -10725 -65544
rect -10625 -65578 -10609 -65544
rect -10483 -65578 -10467 -65544
rect -10367 -65578 -10351 -65544
rect -10225 -65578 -10209 -65544
rect -10109 -65578 -10093 -65544
rect -9967 -65578 -9951 -65544
rect -9851 -65578 -9835 -65544
rect -11337 -65637 -11303 -65621
rect -11337 -66029 -11303 -66013
rect -11079 -65637 -11045 -65621
rect -11079 -66029 -11045 -66013
rect -10821 -65637 -10787 -65621
rect -10821 -66029 -10787 -66013
rect -10563 -65637 -10529 -65621
rect -10563 -66029 -10529 -66013
rect -10305 -65637 -10271 -65621
rect -10305 -66029 -10271 -66013
rect -10047 -65637 -10013 -65621
rect -10047 -66029 -10013 -66013
rect -9789 -65637 -9755 -65621
rect -9789 -66029 -9755 -66013
rect -11257 -66106 -11241 -66072
rect -11141 -66106 -11125 -66072
rect -10999 -66106 -10983 -66072
rect -10883 -66106 -10867 -66072
rect -10741 -66106 -10725 -66072
rect -10625 -66106 -10609 -66072
rect -10483 -66106 -10467 -66072
rect -10367 -66106 -10351 -66072
rect -10225 -66106 -10209 -66072
rect -10109 -66106 -10093 -66072
rect -9967 -66106 -9951 -66072
rect -9851 -66106 -9835 -66072
rect -11257 -66438 -11241 -66404
rect -11141 -66438 -11125 -66404
rect -10999 -66438 -10983 -66404
rect -10883 -66438 -10867 -66404
rect -10741 -66438 -10725 -66404
rect -10625 -66438 -10609 -66404
rect -10483 -66438 -10467 -66404
rect -10367 -66438 -10351 -66404
rect -10225 -66438 -10209 -66404
rect -10109 -66438 -10093 -66404
rect -9967 -66438 -9951 -66404
rect -9851 -66438 -9835 -66404
rect -11337 -66497 -11303 -66481
rect -11337 -66889 -11303 -66873
rect -11079 -66497 -11045 -66481
rect -11079 -66889 -11045 -66873
rect -10821 -66497 -10787 -66481
rect -10821 -66889 -10787 -66873
rect -10563 -66497 -10529 -66481
rect -10563 -66889 -10529 -66873
rect -10305 -66497 -10271 -66481
rect -10305 -66889 -10271 -66873
rect -10047 -66497 -10013 -66481
rect -10047 -66889 -10013 -66873
rect -9789 -66497 -9755 -66481
rect -9789 -66889 -9755 -66873
rect -11257 -66966 -11241 -66932
rect -11141 -66966 -11125 -66932
rect -10999 -66966 -10983 -66932
rect -10883 -66966 -10867 -66932
rect -10741 -66966 -10725 -66932
rect -10625 -66966 -10609 -66932
rect -10483 -66966 -10467 -66932
rect -10367 -66966 -10351 -66932
rect -10225 -66966 -10209 -66932
rect -10109 -66966 -10093 -66932
rect -9967 -66966 -9951 -66932
rect -9851 -66966 -9835 -66932
rect -13460 -67530 -13360 -67368
rect -12004 -67341 -11962 -67299
rect -12004 -67375 -11996 -67341
rect -12004 -67409 -11962 -67375
rect -12004 -67443 -11996 -67409
rect -12004 -67477 -11962 -67443
rect -12004 -67511 -11996 -67477
rect -12004 -67527 -11962 -67511
rect -11928 -67341 -11862 -67333
rect -11928 -67375 -11912 -67341
rect -11878 -67375 -11862 -67341
rect -11928 -67409 -11862 -67375
rect -11928 -67443 -11912 -67409
rect -11878 -67443 -11862 -67409
rect -11928 -67477 -11862 -67443
rect -11928 -67511 -11912 -67477
rect -11878 -67511 -11862 -67477
rect -11928 -67529 -11862 -67511
rect -12008 -67610 -12004 -67563
rect -11956 -67610 -11942 -67563
rect -12008 -67611 -11992 -67610
rect -11958 -67611 -11942 -67610
rect -11908 -67620 -11862 -67529
rect -11684 -67530 -11584 -67368
rect -7684 -64588 -7584 -64426
rect -8072 -67299 -8043 -67265
rect -8009 -67299 -7951 -67265
rect -7917 -67299 -7859 -67265
rect -7825 -67299 -7796 -67265
rect -5460 -64588 -5360 -64426
rect -7257 -65578 -7241 -65544
rect -7141 -65578 -7125 -65544
rect -6999 -65578 -6983 -65544
rect -6883 -65578 -6867 -65544
rect -6741 -65578 -6725 -65544
rect -6625 -65578 -6609 -65544
rect -6483 -65578 -6467 -65544
rect -6367 -65578 -6351 -65544
rect -6225 -65578 -6209 -65544
rect -6109 -65578 -6093 -65544
rect -5967 -65578 -5951 -65544
rect -5851 -65578 -5835 -65544
rect -7337 -65637 -7303 -65621
rect -7337 -66029 -7303 -66013
rect -7079 -65637 -7045 -65621
rect -7079 -66029 -7045 -66013
rect -6821 -65637 -6787 -65621
rect -6821 -66029 -6787 -66013
rect -6563 -65637 -6529 -65621
rect -6563 -66029 -6529 -66013
rect -6305 -65637 -6271 -65621
rect -6305 -66029 -6271 -66013
rect -6047 -65637 -6013 -65621
rect -6047 -66029 -6013 -66013
rect -5789 -65637 -5755 -65621
rect -5789 -66029 -5755 -66013
rect -7257 -66106 -7241 -66072
rect -7141 -66106 -7125 -66072
rect -6999 -66106 -6983 -66072
rect -6883 -66106 -6867 -66072
rect -6741 -66106 -6725 -66072
rect -6625 -66106 -6609 -66072
rect -6483 -66106 -6467 -66072
rect -6367 -66106 -6351 -66072
rect -6225 -66106 -6209 -66072
rect -6109 -66106 -6093 -66072
rect -5967 -66106 -5951 -66072
rect -5851 -66106 -5835 -66072
rect -7257 -66438 -7241 -66404
rect -7141 -66438 -7125 -66404
rect -6999 -66438 -6983 -66404
rect -6883 -66438 -6867 -66404
rect -6741 -66438 -6725 -66404
rect -6625 -66438 -6609 -66404
rect -6483 -66438 -6467 -66404
rect -6367 -66438 -6351 -66404
rect -6225 -66438 -6209 -66404
rect -6109 -66438 -6093 -66404
rect -5967 -66438 -5951 -66404
rect -5851 -66438 -5835 -66404
rect -7337 -66497 -7303 -66481
rect -7337 -66889 -7303 -66873
rect -7079 -66497 -7045 -66481
rect -7079 -66889 -7045 -66873
rect -6821 -66497 -6787 -66481
rect -6821 -66889 -6787 -66873
rect -6563 -66497 -6529 -66481
rect -6563 -66889 -6529 -66873
rect -6305 -66497 -6271 -66481
rect -6305 -66889 -6271 -66873
rect -6047 -66497 -6013 -66481
rect -6047 -66889 -6013 -66873
rect -5789 -66497 -5755 -66481
rect -5789 -66889 -5755 -66873
rect -7257 -66966 -7241 -66932
rect -7141 -66966 -7125 -66932
rect -6999 -66966 -6983 -66932
rect -6883 -66966 -6867 -66932
rect -6741 -66966 -6725 -66932
rect -6625 -66966 -6609 -66932
rect -6483 -66966 -6467 -66932
rect -6367 -66966 -6351 -66932
rect -6225 -66966 -6209 -66932
rect -6109 -66966 -6093 -66932
rect -5967 -66966 -5951 -66932
rect -5851 -66966 -5835 -66932
rect -9460 -67530 -9360 -67368
rect -8004 -67341 -7962 -67299
rect -8004 -67375 -7996 -67341
rect -8004 -67409 -7962 -67375
rect -8004 -67443 -7996 -67409
rect -8004 -67477 -7962 -67443
rect -8004 -67511 -7996 -67477
rect -8004 -67527 -7962 -67511
rect -7928 -67341 -7862 -67333
rect -7928 -67375 -7912 -67341
rect -7878 -67375 -7862 -67341
rect -7928 -67409 -7862 -67375
rect -7928 -67443 -7912 -67409
rect -7878 -67443 -7862 -67409
rect -7928 -67477 -7862 -67443
rect -7928 -67511 -7912 -67477
rect -7878 -67511 -7862 -67477
rect -7928 -67529 -7862 -67511
rect -8008 -67610 -8004 -67563
rect -7956 -67610 -7942 -67563
rect -8008 -67611 -7992 -67610
rect -7958 -67611 -7942 -67610
rect -7908 -67620 -7862 -67529
rect -7684 -67530 -7584 -67368
rect -3684 -64588 -3584 -64426
rect -4072 -67299 -4043 -67265
rect -4009 -67299 -3951 -67265
rect -3917 -67299 -3859 -67265
rect -3825 -67299 -3796 -67265
rect -1460 -64588 -1360 -64426
rect -3257 -65578 -3241 -65544
rect -3141 -65578 -3125 -65544
rect -2999 -65578 -2983 -65544
rect -2883 -65578 -2867 -65544
rect -2741 -65578 -2725 -65544
rect -2625 -65578 -2609 -65544
rect -2483 -65578 -2467 -65544
rect -2367 -65578 -2351 -65544
rect -2225 -65578 -2209 -65544
rect -2109 -65578 -2093 -65544
rect -1967 -65578 -1951 -65544
rect -1851 -65578 -1835 -65544
rect -3337 -65637 -3303 -65621
rect -3337 -66029 -3303 -66013
rect -3079 -65637 -3045 -65621
rect -3079 -66029 -3045 -66013
rect -2821 -65637 -2787 -65621
rect -2821 -66029 -2787 -66013
rect -2563 -65637 -2529 -65621
rect -2563 -66029 -2529 -66013
rect -2305 -65637 -2271 -65621
rect -2305 -66029 -2271 -66013
rect -2047 -65637 -2013 -65621
rect -2047 -66029 -2013 -66013
rect -1789 -65637 -1755 -65621
rect -1789 -66029 -1755 -66013
rect -3257 -66106 -3241 -66072
rect -3141 -66106 -3125 -66072
rect -2999 -66106 -2983 -66072
rect -2883 -66106 -2867 -66072
rect -2741 -66106 -2725 -66072
rect -2625 -66106 -2609 -66072
rect -2483 -66106 -2467 -66072
rect -2367 -66106 -2351 -66072
rect -2225 -66106 -2209 -66072
rect -2109 -66106 -2093 -66072
rect -1967 -66106 -1951 -66072
rect -1851 -66106 -1835 -66072
rect -3257 -66438 -3241 -66404
rect -3141 -66438 -3125 -66404
rect -2999 -66438 -2983 -66404
rect -2883 -66438 -2867 -66404
rect -2741 -66438 -2725 -66404
rect -2625 -66438 -2609 -66404
rect -2483 -66438 -2467 -66404
rect -2367 -66438 -2351 -66404
rect -2225 -66438 -2209 -66404
rect -2109 -66438 -2093 -66404
rect -1967 -66438 -1951 -66404
rect -1851 -66438 -1835 -66404
rect -3337 -66497 -3303 -66481
rect -3337 -66889 -3303 -66873
rect -3079 -66497 -3045 -66481
rect -3079 -66889 -3045 -66873
rect -2821 -66497 -2787 -66481
rect -2821 -66889 -2787 -66873
rect -2563 -66497 -2529 -66481
rect -2563 -66889 -2529 -66873
rect -2305 -66497 -2271 -66481
rect -2305 -66889 -2271 -66873
rect -2047 -66497 -2013 -66481
rect -2047 -66889 -2013 -66873
rect -1789 -66497 -1755 -66481
rect -1789 -66889 -1755 -66873
rect -3257 -66966 -3241 -66932
rect -3141 -66966 -3125 -66932
rect -2999 -66966 -2983 -66932
rect -2883 -66966 -2867 -66932
rect -2741 -66966 -2725 -66932
rect -2625 -66966 -2609 -66932
rect -2483 -66966 -2467 -66932
rect -2367 -66966 -2351 -66932
rect -2225 -66966 -2209 -66932
rect -2109 -66966 -2093 -66932
rect -1967 -66966 -1951 -66932
rect -1851 -66966 -1835 -66932
rect -5460 -67530 -5360 -67368
rect -4004 -67341 -3962 -67299
rect -4004 -67375 -3996 -67341
rect -4004 -67409 -3962 -67375
rect -4004 -67443 -3996 -67409
rect -4004 -67477 -3962 -67443
rect -4004 -67511 -3996 -67477
rect -4004 -67527 -3962 -67511
rect -3928 -67341 -3862 -67333
rect -3928 -67375 -3912 -67341
rect -3878 -67375 -3862 -67341
rect -3928 -67409 -3862 -67375
rect -3928 -67443 -3912 -67409
rect -3878 -67443 -3862 -67409
rect -3928 -67477 -3862 -67443
rect -3928 -67511 -3912 -67477
rect -3878 -67511 -3862 -67477
rect -3928 -67529 -3862 -67511
rect -4008 -67610 -4004 -67563
rect -3956 -67610 -3942 -67563
rect -4008 -67611 -3992 -67610
rect -3958 -67611 -3942 -67610
rect -3908 -67620 -3862 -67529
rect -3684 -67530 -3584 -67368
rect 316 -64588 416 -64426
rect -72 -67299 -43 -67265
rect -9 -67299 49 -67265
rect 83 -67299 141 -67265
rect 175 -67299 204 -67265
rect 2540 -64588 2640 -64426
rect 743 -65578 759 -65544
rect 859 -65578 875 -65544
rect 1001 -65578 1017 -65544
rect 1117 -65578 1133 -65544
rect 1259 -65578 1275 -65544
rect 1375 -65578 1391 -65544
rect 1517 -65578 1533 -65544
rect 1633 -65578 1649 -65544
rect 1775 -65578 1791 -65544
rect 1891 -65578 1907 -65544
rect 2033 -65578 2049 -65544
rect 2149 -65578 2165 -65544
rect 663 -65637 697 -65621
rect 663 -66029 697 -66013
rect 921 -65637 955 -65621
rect 921 -66029 955 -66013
rect 1179 -65637 1213 -65621
rect 1179 -66029 1213 -66013
rect 1437 -65637 1471 -65621
rect 1437 -66029 1471 -66013
rect 1695 -65637 1729 -65621
rect 1695 -66029 1729 -66013
rect 1953 -65637 1987 -65621
rect 1953 -66029 1987 -66013
rect 2211 -65637 2245 -65621
rect 2211 -66029 2245 -66013
rect 743 -66106 759 -66072
rect 859 -66106 875 -66072
rect 1001 -66106 1017 -66072
rect 1117 -66106 1133 -66072
rect 1259 -66106 1275 -66072
rect 1375 -66106 1391 -66072
rect 1517 -66106 1533 -66072
rect 1633 -66106 1649 -66072
rect 1775 -66106 1791 -66072
rect 1891 -66106 1907 -66072
rect 2033 -66106 2049 -66072
rect 2149 -66106 2165 -66072
rect 743 -66438 759 -66404
rect 859 -66438 875 -66404
rect 1001 -66438 1017 -66404
rect 1117 -66438 1133 -66404
rect 1259 -66438 1275 -66404
rect 1375 -66438 1391 -66404
rect 1517 -66438 1533 -66404
rect 1633 -66438 1649 -66404
rect 1775 -66438 1791 -66404
rect 1891 -66438 1907 -66404
rect 2033 -66438 2049 -66404
rect 2149 -66438 2165 -66404
rect 663 -66497 697 -66481
rect 663 -66889 697 -66873
rect 921 -66497 955 -66481
rect 921 -66889 955 -66873
rect 1179 -66497 1213 -66481
rect 1179 -66889 1213 -66873
rect 1437 -66497 1471 -66481
rect 1437 -66889 1471 -66873
rect 1695 -66497 1729 -66481
rect 1695 -66889 1729 -66873
rect 1953 -66497 1987 -66481
rect 1953 -66889 1987 -66873
rect 2211 -66497 2245 -66481
rect 2211 -66889 2245 -66873
rect 743 -66966 759 -66932
rect 859 -66966 875 -66932
rect 1001 -66966 1017 -66932
rect 1117 -66966 1133 -66932
rect 1259 -66966 1275 -66932
rect 1375 -66966 1391 -66932
rect 1517 -66966 1533 -66932
rect 1633 -66966 1649 -66932
rect 1775 -66966 1791 -66932
rect 1891 -66966 1907 -66932
rect 2033 -66966 2049 -66932
rect 2149 -66966 2165 -66932
rect -1460 -67530 -1360 -67368
rect -4 -67341 38 -67299
rect -4 -67375 4 -67341
rect -4 -67409 38 -67375
rect -4 -67443 4 -67409
rect -4 -67477 38 -67443
rect -4 -67511 4 -67477
rect -4 -67527 38 -67511
rect 72 -67341 138 -67333
rect 72 -67375 88 -67341
rect 122 -67375 138 -67341
rect 72 -67409 138 -67375
rect 72 -67443 88 -67409
rect 122 -67443 138 -67409
rect 72 -67477 138 -67443
rect 72 -67511 88 -67477
rect 122 -67511 138 -67477
rect 72 -67529 138 -67511
rect -8 -67610 -4 -67563
rect 44 -67610 58 -67563
rect -8 -67611 8 -67610
rect 42 -67611 58 -67610
rect 92 -67620 138 -67529
rect 316 -67530 416 -67368
rect 4316 -64588 4416 -64426
rect 3928 -67299 3957 -67265
rect 3991 -67299 4049 -67265
rect 4083 -67299 4141 -67265
rect 4175 -67299 4204 -67265
rect 6540 -64588 6640 -64426
rect 4743 -65578 4759 -65544
rect 4859 -65578 4875 -65544
rect 5001 -65578 5017 -65544
rect 5117 -65578 5133 -65544
rect 5259 -65578 5275 -65544
rect 5375 -65578 5391 -65544
rect 5517 -65578 5533 -65544
rect 5633 -65578 5649 -65544
rect 5775 -65578 5791 -65544
rect 5891 -65578 5907 -65544
rect 6033 -65578 6049 -65544
rect 6149 -65578 6165 -65544
rect 4663 -65637 4697 -65621
rect 4663 -66029 4697 -66013
rect 4921 -65637 4955 -65621
rect 4921 -66029 4955 -66013
rect 5179 -65637 5213 -65621
rect 5179 -66029 5213 -66013
rect 5437 -65637 5471 -65621
rect 5437 -66029 5471 -66013
rect 5695 -65637 5729 -65621
rect 5695 -66029 5729 -66013
rect 5953 -65637 5987 -65621
rect 5953 -66029 5987 -66013
rect 6211 -65637 6245 -65621
rect 6211 -66029 6245 -66013
rect 4743 -66106 4759 -66072
rect 4859 -66106 4875 -66072
rect 5001 -66106 5017 -66072
rect 5117 -66106 5133 -66072
rect 5259 -66106 5275 -66072
rect 5375 -66106 5391 -66072
rect 5517 -66106 5533 -66072
rect 5633 -66106 5649 -66072
rect 5775 -66106 5791 -66072
rect 5891 -66106 5907 -66072
rect 6033 -66106 6049 -66072
rect 6149 -66106 6165 -66072
rect 4743 -66438 4759 -66404
rect 4859 -66438 4875 -66404
rect 5001 -66438 5017 -66404
rect 5117 -66438 5133 -66404
rect 5259 -66438 5275 -66404
rect 5375 -66438 5391 -66404
rect 5517 -66438 5533 -66404
rect 5633 -66438 5649 -66404
rect 5775 -66438 5791 -66404
rect 5891 -66438 5907 -66404
rect 6033 -66438 6049 -66404
rect 6149 -66438 6165 -66404
rect 4663 -66497 4697 -66481
rect 4663 -66889 4697 -66873
rect 4921 -66497 4955 -66481
rect 4921 -66889 4955 -66873
rect 5179 -66497 5213 -66481
rect 5179 -66889 5213 -66873
rect 5437 -66497 5471 -66481
rect 5437 -66889 5471 -66873
rect 5695 -66497 5729 -66481
rect 5695 -66889 5729 -66873
rect 5953 -66497 5987 -66481
rect 5953 -66889 5987 -66873
rect 6211 -66497 6245 -66481
rect 6211 -66889 6245 -66873
rect 4743 -66966 4759 -66932
rect 4859 -66966 4875 -66932
rect 5001 -66966 5017 -66932
rect 5117 -66966 5133 -66932
rect 5259 -66966 5275 -66932
rect 5375 -66966 5391 -66932
rect 5517 -66966 5533 -66932
rect 5633 -66966 5649 -66932
rect 5775 -66966 5791 -66932
rect 5891 -66966 5907 -66932
rect 6033 -66966 6049 -66932
rect 6149 -66966 6165 -66932
rect 2540 -67530 2640 -67368
rect 3996 -67341 4038 -67299
rect 3996 -67375 4004 -67341
rect 3996 -67409 4038 -67375
rect 3996 -67443 4004 -67409
rect 3996 -67477 4038 -67443
rect 3996 -67511 4004 -67477
rect 3996 -67527 4038 -67511
rect 4072 -67341 4138 -67333
rect 4072 -67375 4088 -67341
rect 4122 -67375 4138 -67341
rect 4072 -67409 4138 -67375
rect 4072 -67443 4088 -67409
rect 4122 -67443 4138 -67409
rect 4072 -67477 4138 -67443
rect 4072 -67511 4088 -67477
rect 4122 -67511 4138 -67477
rect 4072 -67529 4138 -67511
rect 3992 -67610 3996 -67563
rect 4044 -67610 4058 -67563
rect 3992 -67611 4008 -67610
rect 4042 -67611 4058 -67610
rect 4092 -67620 4138 -67529
rect 4316 -67530 4416 -67368
rect 6540 -67530 6640 -67368
rect -28008 -67661 -27962 -67645
rect -27908 -67649 -27902 -67620
rect -28008 -67695 -27996 -67661
rect -28008 -67729 -27962 -67695
rect -28008 -67763 -27996 -67729
rect -28008 -67809 -27962 -67763
rect -27928 -67661 -27902 -67649
rect -27928 -67695 -27912 -67661
rect -24008 -67661 -23962 -67645
rect -23908 -67649 -23902 -67620
rect -27878 -67695 -27862 -67668
rect -27928 -67729 -27862 -67695
rect -27928 -67763 -27912 -67729
rect -27878 -67763 -27862 -67729
rect -27928 -67775 -27862 -67763
rect -24008 -67695 -23996 -67661
rect -24008 -67729 -23962 -67695
rect -24008 -67763 -23996 -67729
rect -28072 -67843 -28043 -67809
rect -28009 -67843 -27951 -67809
rect -27917 -67843 -27859 -67809
rect -27825 -67843 -27796 -67809
rect -27684 -67928 -27584 -67766
rect -25460 -67928 -25360 -67766
rect -24008 -67809 -23962 -67763
rect -23928 -67661 -23902 -67649
rect -23928 -67695 -23912 -67661
rect -20008 -67661 -19962 -67645
rect -19908 -67649 -19902 -67620
rect -23878 -67695 -23862 -67668
rect -23928 -67729 -23862 -67695
rect -23928 -67763 -23912 -67729
rect -23878 -67763 -23862 -67729
rect -23928 -67775 -23862 -67763
rect -20008 -67695 -19996 -67661
rect -20008 -67729 -19962 -67695
rect -20008 -67763 -19996 -67729
rect -24072 -67843 -24043 -67809
rect -24009 -67843 -23951 -67809
rect -23917 -67843 -23859 -67809
rect -23825 -67843 -23796 -67809
rect -27262 -68280 -27246 -68246
rect -27146 -68280 -27130 -68246
rect -27004 -68280 -26988 -68246
rect -26888 -68280 -26872 -68246
rect -26746 -68280 -26730 -68246
rect -26630 -68280 -26614 -68246
rect -26488 -68280 -26472 -68246
rect -26372 -68280 -26356 -68246
rect -26230 -68280 -26214 -68246
rect -26114 -68280 -26098 -68246
rect -25972 -68280 -25956 -68246
rect -25856 -68280 -25840 -68246
rect -27342 -68330 -27308 -68314
rect -27342 -68722 -27308 -68706
rect -27084 -68330 -27050 -68314
rect -27084 -68722 -27050 -68706
rect -26826 -68330 -26792 -68314
rect -26826 -68722 -26792 -68706
rect -26568 -68330 -26534 -68314
rect -26568 -68722 -26534 -68706
rect -26310 -68330 -26276 -68314
rect -26310 -68722 -26276 -68706
rect -26052 -68330 -26018 -68314
rect -26052 -68722 -26018 -68706
rect -25794 -68330 -25760 -68314
rect -25794 -68722 -25760 -68706
rect -27262 -68790 -27246 -68756
rect -27146 -68790 -27130 -68756
rect -27004 -68790 -26988 -68756
rect -26888 -68790 -26872 -68756
rect -26746 -68790 -26730 -68756
rect -26630 -68790 -26614 -68756
rect -26488 -68790 -26472 -68756
rect -26372 -68790 -26356 -68756
rect -26230 -68790 -26214 -68756
rect -26114 -68790 -26098 -68756
rect -25972 -68790 -25956 -68756
rect -25856 -68790 -25840 -68756
rect -27684 -69810 -27584 -69648
rect -25460 -69810 -25360 -69648
rect -23684 -67928 -23584 -67766
rect -21460 -67928 -21360 -67766
rect -20008 -67809 -19962 -67763
rect -19928 -67661 -19902 -67649
rect -19928 -67695 -19912 -67661
rect -16008 -67661 -15962 -67645
rect -15908 -67649 -15902 -67620
rect -19878 -67695 -19862 -67668
rect -19928 -67729 -19862 -67695
rect -19928 -67763 -19912 -67729
rect -19878 -67763 -19862 -67729
rect -19928 -67775 -19862 -67763
rect -16008 -67695 -15996 -67661
rect -16008 -67729 -15962 -67695
rect -16008 -67763 -15996 -67729
rect -20072 -67843 -20043 -67809
rect -20009 -67843 -19951 -67809
rect -19917 -67843 -19859 -67809
rect -19825 -67843 -19796 -67809
rect -23262 -68280 -23246 -68246
rect -23146 -68280 -23130 -68246
rect -23004 -68280 -22988 -68246
rect -22888 -68280 -22872 -68246
rect -22746 -68280 -22730 -68246
rect -22630 -68280 -22614 -68246
rect -22488 -68280 -22472 -68246
rect -22372 -68280 -22356 -68246
rect -22230 -68280 -22214 -68246
rect -22114 -68280 -22098 -68246
rect -21972 -68280 -21956 -68246
rect -21856 -68280 -21840 -68246
rect -23342 -68330 -23308 -68314
rect -23342 -68722 -23308 -68706
rect -23084 -68330 -23050 -68314
rect -23084 -68722 -23050 -68706
rect -22826 -68330 -22792 -68314
rect -22826 -68722 -22792 -68706
rect -22568 -68330 -22534 -68314
rect -22568 -68722 -22534 -68706
rect -22310 -68330 -22276 -68314
rect -22310 -68722 -22276 -68706
rect -22052 -68330 -22018 -68314
rect -22052 -68722 -22018 -68706
rect -21794 -68330 -21760 -68314
rect -21794 -68722 -21760 -68706
rect -23262 -68790 -23246 -68756
rect -23146 -68790 -23130 -68756
rect -23004 -68790 -22988 -68756
rect -22888 -68790 -22872 -68756
rect -22746 -68790 -22730 -68756
rect -22630 -68790 -22614 -68756
rect -22488 -68790 -22472 -68756
rect -22372 -68790 -22356 -68756
rect -22230 -68790 -22214 -68756
rect -22114 -68790 -22098 -68756
rect -21972 -68790 -21956 -68756
rect -21856 -68790 -21840 -68756
rect -23684 -69810 -23584 -69648
rect -21460 -69810 -21360 -69648
rect -19684 -67928 -19584 -67766
rect -17460 -67928 -17360 -67766
rect -16008 -67809 -15962 -67763
rect -15928 -67661 -15902 -67649
rect -15928 -67695 -15912 -67661
rect -12008 -67661 -11962 -67645
rect -11908 -67649 -11902 -67620
rect -15878 -67695 -15862 -67668
rect -15928 -67729 -15862 -67695
rect -15928 -67763 -15912 -67729
rect -15878 -67763 -15862 -67729
rect -15928 -67775 -15862 -67763
rect -12008 -67695 -11996 -67661
rect -12008 -67729 -11962 -67695
rect -12008 -67763 -11996 -67729
rect -16072 -67843 -16043 -67809
rect -16009 -67843 -15951 -67809
rect -15917 -67843 -15859 -67809
rect -15825 -67843 -15796 -67809
rect -19262 -68280 -19246 -68246
rect -19146 -68280 -19130 -68246
rect -19004 -68280 -18988 -68246
rect -18888 -68280 -18872 -68246
rect -18746 -68280 -18730 -68246
rect -18630 -68280 -18614 -68246
rect -18488 -68280 -18472 -68246
rect -18372 -68280 -18356 -68246
rect -18230 -68280 -18214 -68246
rect -18114 -68280 -18098 -68246
rect -17972 -68280 -17956 -68246
rect -17856 -68280 -17840 -68246
rect -19342 -68330 -19308 -68314
rect -19342 -68722 -19308 -68706
rect -19084 -68330 -19050 -68314
rect -19084 -68722 -19050 -68706
rect -18826 -68330 -18792 -68314
rect -18826 -68722 -18792 -68706
rect -18568 -68330 -18534 -68314
rect -18568 -68722 -18534 -68706
rect -18310 -68330 -18276 -68314
rect -18310 -68722 -18276 -68706
rect -18052 -68330 -18018 -68314
rect -18052 -68722 -18018 -68706
rect -17794 -68330 -17760 -68314
rect -17794 -68722 -17760 -68706
rect -19262 -68790 -19246 -68756
rect -19146 -68790 -19130 -68756
rect -19004 -68790 -18988 -68756
rect -18888 -68790 -18872 -68756
rect -18746 -68790 -18730 -68756
rect -18630 -68790 -18614 -68756
rect -18488 -68790 -18472 -68756
rect -18372 -68790 -18356 -68756
rect -18230 -68790 -18214 -68756
rect -18114 -68790 -18098 -68756
rect -17972 -68790 -17956 -68756
rect -17856 -68790 -17840 -68756
rect -19684 -69810 -19584 -69648
rect -17460 -69810 -17360 -69648
rect -15684 -67928 -15584 -67766
rect -13460 -67928 -13360 -67766
rect -12008 -67809 -11962 -67763
rect -11928 -67661 -11902 -67649
rect -11928 -67695 -11912 -67661
rect -8008 -67661 -7962 -67645
rect -7908 -67649 -7902 -67620
rect -11878 -67695 -11862 -67668
rect -11928 -67729 -11862 -67695
rect -11928 -67763 -11912 -67729
rect -11878 -67763 -11862 -67729
rect -11928 -67775 -11862 -67763
rect -8008 -67695 -7996 -67661
rect -8008 -67729 -7962 -67695
rect -8008 -67763 -7996 -67729
rect -12072 -67843 -12043 -67809
rect -12009 -67843 -11951 -67809
rect -11917 -67843 -11859 -67809
rect -11825 -67843 -11796 -67809
rect -15262 -68280 -15246 -68246
rect -15146 -68280 -15130 -68246
rect -15004 -68280 -14988 -68246
rect -14888 -68280 -14872 -68246
rect -14746 -68280 -14730 -68246
rect -14630 -68280 -14614 -68246
rect -14488 -68280 -14472 -68246
rect -14372 -68280 -14356 -68246
rect -14230 -68280 -14214 -68246
rect -14114 -68280 -14098 -68246
rect -13972 -68280 -13956 -68246
rect -13856 -68280 -13840 -68246
rect -15342 -68330 -15308 -68314
rect -15342 -68722 -15308 -68706
rect -15084 -68330 -15050 -68314
rect -15084 -68722 -15050 -68706
rect -14826 -68330 -14792 -68314
rect -14826 -68722 -14792 -68706
rect -14568 -68330 -14534 -68314
rect -14568 -68722 -14534 -68706
rect -14310 -68330 -14276 -68314
rect -14310 -68722 -14276 -68706
rect -14052 -68330 -14018 -68314
rect -14052 -68722 -14018 -68706
rect -13794 -68330 -13760 -68314
rect -13794 -68722 -13760 -68706
rect -15262 -68790 -15246 -68756
rect -15146 -68790 -15130 -68756
rect -15004 -68790 -14988 -68756
rect -14888 -68790 -14872 -68756
rect -14746 -68790 -14730 -68756
rect -14630 -68790 -14614 -68756
rect -14488 -68790 -14472 -68756
rect -14372 -68790 -14356 -68756
rect -14230 -68790 -14214 -68756
rect -14114 -68790 -14098 -68756
rect -13972 -68790 -13956 -68756
rect -13856 -68790 -13840 -68756
rect -15684 -69810 -15584 -69648
rect -13460 -69810 -13360 -69648
rect -11684 -67928 -11584 -67766
rect -9460 -67928 -9360 -67766
rect -8008 -67809 -7962 -67763
rect -7928 -67661 -7902 -67649
rect -7928 -67695 -7912 -67661
rect -4008 -67661 -3962 -67645
rect -3908 -67649 -3902 -67620
rect -7878 -67695 -7862 -67668
rect -7928 -67729 -7862 -67695
rect -7928 -67763 -7912 -67729
rect -7878 -67763 -7862 -67729
rect -7928 -67775 -7862 -67763
rect -4008 -67695 -3996 -67661
rect -4008 -67729 -3962 -67695
rect -4008 -67763 -3996 -67729
rect -8072 -67843 -8043 -67809
rect -8009 -67843 -7951 -67809
rect -7917 -67843 -7859 -67809
rect -7825 -67843 -7796 -67809
rect -11262 -68280 -11246 -68246
rect -11146 -68280 -11130 -68246
rect -11004 -68280 -10988 -68246
rect -10888 -68280 -10872 -68246
rect -10746 -68280 -10730 -68246
rect -10630 -68280 -10614 -68246
rect -10488 -68280 -10472 -68246
rect -10372 -68280 -10356 -68246
rect -10230 -68280 -10214 -68246
rect -10114 -68280 -10098 -68246
rect -9972 -68280 -9956 -68246
rect -9856 -68280 -9840 -68246
rect -11342 -68330 -11308 -68314
rect -11342 -68722 -11308 -68706
rect -11084 -68330 -11050 -68314
rect -11084 -68722 -11050 -68706
rect -10826 -68330 -10792 -68314
rect -10826 -68722 -10792 -68706
rect -10568 -68330 -10534 -68314
rect -10568 -68722 -10534 -68706
rect -10310 -68330 -10276 -68314
rect -10310 -68722 -10276 -68706
rect -10052 -68330 -10018 -68314
rect -10052 -68722 -10018 -68706
rect -9794 -68330 -9760 -68314
rect -9794 -68722 -9760 -68706
rect -11262 -68790 -11246 -68756
rect -11146 -68790 -11130 -68756
rect -11004 -68790 -10988 -68756
rect -10888 -68790 -10872 -68756
rect -10746 -68790 -10730 -68756
rect -10630 -68790 -10614 -68756
rect -10488 -68790 -10472 -68756
rect -10372 -68790 -10356 -68756
rect -10230 -68790 -10214 -68756
rect -10114 -68790 -10098 -68756
rect -9972 -68790 -9956 -68756
rect -9856 -68790 -9840 -68756
rect -11684 -69810 -11584 -69648
rect -9460 -69810 -9360 -69648
rect -7684 -67928 -7584 -67766
rect -5460 -67928 -5360 -67766
rect -4008 -67809 -3962 -67763
rect -3928 -67661 -3902 -67649
rect -3928 -67695 -3912 -67661
rect -8 -67661 38 -67645
rect 92 -67649 98 -67620
rect -3878 -67695 -3862 -67668
rect -3928 -67729 -3862 -67695
rect -3928 -67763 -3912 -67729
rect -3878 -67763 -3862 -67729
rect -3928 -67775 -3862 -67763
rect -8 -67695 4 -67661
rect -8 -67729 38 -67695
rect -8 -67763 4 -67729
rect -4072 -67843 -4043 -67809
rect -4009 -67843 -3951 -67809
rect -3917 -67843 -3859 -67809
rect -3825 -67843 -3796 -67809
rect -7262 -68280 -7246 -68246
rect -7146 -68280 -7130 -68246
rect -7004 -68280 -6988 -68246
rect -6888 -68280 -6872 -68246
rect -6746 -68280 -6730 -68246
rect -6630 -68280 -6614 -68246
rect -6488 -68280 -6472 -68246
rect -6372 -68280 -6356 -68246
rect -6230 -68280 -6214 -68246
rect -6114 -68280 -6098 -68246
rect -5972 -68280 -5956 -68246
rect -5856 -68280 -5840 -68246
rect -7342 -68330 -7308 -68314
rect -7342 -68722 -7308 -68706
rect -7084 -68330 -7050 -68314
rect -7084 -68722 -7050 -68706
rect -6826 -68330 -6792 -68314
rect -6826 -68722 -6792 -68706
rect -6568 -68330 -6534 -68314
rect -6568 -68722 -6534 -68706
rect -6310 -68330 -6276 -68314
rect -6310 -68722 -6276 -68706
rect -6052 -68330 -6018 -68314
rect -6052 -68722 -6018 -68706
rect -5794 -68330 -5760 -68314
rect -5794 -68722 -5760 -68706
rect -7262 -68790 -7246 -68756
rect -7146 -68790 -7130 -68756
rect -7004 -68790 -6988 -68756
rect -6888 -68790 -6872 -68756
rect -6746 -68790 -6730 -68756
rect -6630 -68790 -6614 -68756
rect -6488 -68790 -6472 -68756
rect -6372 -68790 -6356 -68756
rect -6230 -68790 -6214 -68756
rect -6114 -68790 -6098 -68756
rect -5972 -68790 -5956 -68756
rect -5856 -68790 -5840 -68756
rect -7684 -69810 -7584 -69648
rect -5460 -69810 -5360 -69648
rect -3684 -67928 -3584 -67766
rect -1460 -67928 -1360 -67766
rect -8 -67809 38 -67763
rect 72 -67661 98 -67649
rect 72 -67695 88 -67661
rect 3992 -67661 4038 -67645
rect 4092 -67649 4098 -67620
rect 122 -67695 138 -67668
rect 72 -67729 138 -67695
rect 72 -67763 88 -67729
rect 122 -67763 138 -67729
rect 72 -67775 138 -67763
rect 3992 -67695 4004 -67661
rect 3992 -67729 4038 -67695
rect 3992 -67763 4004 -67729
rect -72 -67843 -43 -67809
rect -9 -67843 49 -67809
rect 83 -67843 141 -67809
rect 175 -67843 204 -67809
rect -3262 -68280 -3246 -68246
rect -3146 -68280 -3130 -68246
rect -3004 -68280 -2988 -68246
rect -2888 -68280 -2872 -68246
rect -2746 -68280 -2730 -68246
rect -2630 -68280 -2614 -68246
rect -2488 -68280 -2472 -68246
rect -2372 -68280 -2356 -68246
rect -2230 -68280 -2214 -68246
rect -2114 -68280 -2098 -68246
rect -1972 -68280 -1956 -68246
rect -1856 -68280 -1840 -68246
rect -3342 -68330 -3308 -68314
rect -3342 -68722 -3308 -68706
rect -3084 -68330 -3050 -68314
rect -3084 -68722 -3050 -68706
rect -2826 -68330 -2792 -68314
rect -2826 -68722 -2792 -68706
rect -2568 -68330 -2534 -68314
rect -2568 -68722 -2534 -68706
rect -2310 -68330 -2276 -68314
rect -2310 -68722 -2276 -68706
rect -2052 -68330 -2018 -68314
rect -2052 -68722 -2018 -68706
rect -1794 -68330 -1760 -68314
rect -1794 -68722 -1760 -68706
rect -3262 -68790 -3246 -68756
rect -3146 -68790 -3130 -68756
rect -3004 -68790 -2988 -68756
rect -2888 -68790 -2872 -68756
rect -2746 -68790 -2730 -68756
rect -2630 -68790 -2614 -68756
rect -2488 -68790 -2472 -68756
rect -2372 -68790 -2356 -68756
rect -2230 -68790 -2214 -68756
rect -2114 -68790 -2098 -68756
rect -1972 -68790 -1956 -68756
rect -1856 -68790 -1840 -68756
rect -3684 -69810 -3584 -69648
rect -1460 -69810 -1360 -69648
rect 316 -67928 416 -67766
rect 2540 -67928 2640 -67766
rect 3992 -67809 4038 -67763
rect 4072 -67661 4098 -67649
rect 4072 -67695 4088 -67661
rect 4122 -67695 4138 -67668
rect 4072 -67729 4138 -67695
rect 4072 -67763 4088 -67729
rect 4122 -67763 4138 -67729
rect 4072 -67775 4138 -67763
rect 3928 -67843 3957 -67809
rect 3991 -67843 4049 -67809
rect 4083 -67843 4141 -67809
rect 4175 -67843 4204 -67809
rect 738 -68280 754 -68246
rect 854 -68280 870 -68246
rect 996 -68280 1012 -68246
rect 1112 -68280 1128 -68246
rect 1254 -68280 1270 -68246
rect 1370 -68280 1386 -68246
rect 1512 -68280 1528 -68246
rect 1628 -68280 1644 -68246
rect 1770 -68280 1786 -68246
rect 1886 -68280 1902 -68246
rect 2028 -68280 2044 -68246
rect 2144 -68280 2160 -68246
rect 658 -68330 692 -68314
rect 658 -68722 692 -68706
rect 916 -68330 950 -68314
rect 916 -68722 950 -68706
rect 1174 -68330 1208 -68314
rect 1174 -68722 1208 -68706
rect 1432 -68330 1466 -68314
rect 1432 -68722 1466 -68706
rect 1690 -68330 1724 -68314
rect 1690 -68722 1724 -68706
rect 1948 -68330 1982 -68314
rect 1948 -68722 1982 -68706
rect 2206 -68330 2240 -68314
rect 2206 -68722 2240 -68706
rect 738 -68790 754 -68756
rect 854 -68790 870 -68756
rect 996 -68790 1012 -68756
rect 1112 -68790 1128 -68756
rect 1254 -68790 1270 -68756
rect 1370 -68790 1386 -68756
rect 1512 -68790 1528 -68756
rect 1628 -68790 1644 -68756
rect 1770 -68790 1786 -68756
rect 1886 -68790 1902 -68756
rect 2028 -68790 2044 -68756
rect 2144 -68790 2160 -68756
rect 316 -69810 416 -69648
rect 2540 -69810 2640 -69648
rect 4316 -67928 4416 -67766
rect 6540 -67928 6640 -67766
rect 4738 -68280 4754 -68246
rect 4854 -68280 4870 -68246
rect 4996 -68280 5012 -68246
rect 5112 -68280 5128 -68246
rect 5254 -68280 5270 -68246
rect 5370 -68280 5386 -68246
rect 5512 -68280 5528 -68246
rect 5628 -68280 5644 -68246
rect 5770 -68280 5786 -68246
rect 5886 -68280 5902 -68246
rect 6028 -68280 6044 -68246
rect 6144 -68280 6160 -68246
rect 4658 -68330 4692 -68314
rect 4658 -68722 4692 -68706
rect 4916 -68330 4950 -68314
rect 4916 -68722 4950 -68706
rect 5174 -68330 5208 -68314
rect 5174 -68722 5208 -68706
rect 5432 -68330 5466 -68314
rect 5432 -68722 5466 -68706
rect 5690 -68330 5724 -68314
rect 5690 -68722 5724 -68706
rect 5948 -68330 5982 -68314
rect 5948 -68722 5982 -68706
rect 6206 -68330 6240 -68314
rect 6206 -68722 6240 -68706
rect 4738 -68790 4754 -68756
rect 4854 -68790 4870 -68756
rect 4996 -68790 5012 -68756
rect 5112 -68790 5128 -68756
rect 5254 -68790 5270 -68756
rect 5370 -68790 5386 -68756
rect 5512 -68790 5528 -68756
rect 5628 -68790 5644 -68756
rect 5770 -68790 5786 -68756
rect 5886 -68790 5902 -68756
rect 6028 -68790 6044 -68756
rect 6144 -68790 6160 -68756
rect 4316 -69810 4416 -69648
rect 6540 -69810 6640 -69648
rect -27684 -70548 -27584 -70386
rect -25460 -70548 -25360 -70386
rect -27262 -71440 -27246 -71406
rect -27146 -71440 -27130 -71406
rect -27004 -71440 -26988 -71406
rect -26888 -71440 -26872 -71406
rect -26746 -71440 -26730 -71406
rect -26630 -71440 -26614 -71406
rect -26488 -71440 -26472 -71406
rect -26372 -71440 -26356 -71406
rect -26230 -71440 -26214 -71406
rect -26114 -71440 -26098 -71406
rect -25972 -71440 -25956 -71406
rect -25856 -71440 -25840 -71406
rect -27342 -71490 -27308 -71474
rect -27342 -71882 -27308 -71866
rect -27084 -71490 -27050 -71474
rect -27084 -71882 -27050 -71866
rect -26826 -71490 -26792 -71474
rect -26826 -71882 -26792 -71866
rect -26568 -71490 -26534 -71474
rect -26568 -71882 -26534 -71866
rect -26310 -71490 -26276 -71474
rect -26310 -71882 -26276 -71866
rect -26052 -71490 -26018 -71474
rect -26052 -71882 -26018 -71866
rect -25794 -71490 -25760 -71474
rect -25794 -71882 -25760 -71866
rect -27262 -71950 -27246 -71916
rect -27146 -71950 -27130 -71916
rect -27004 -71950 -26988 -71916
rect -26888 -71950 -26872 -71916
rect -26746 -71950 -26730 -71916
rect -26630 -71950 -26614 -71916
rect -26488 -71950 -26472 -71916
rect -26372 -71950 -26356 -71916
rect -26230 -71950 -26214 -71916
rect -26114 -71950 -26098 -71916
rect -25972 -71950 -25956 -71916
rect -25856 -71950 -25840 -71916
rect -28072 -72387 -28043 -72353
rect -28009 -72387 -27951 -72353
rect -27917 -72387 -27859 -72353
rect -27825 -72387 -27796 -72353
rect -28008 -72433 -27962 -72387
rect -28008 -72467 -27996 -72433
rect -28008 -72501 -27962 -72467
rect -28008 -72535 -27996 -72501
rect -28008 -72551 -27962 -72535
rect -27928 -72433 -27862 -72421
rect -27684 -72430 -27584 -72268
rect -25460 -72430 -25360 -72268
rect -23684 -70548 -23584 -70386
rect -21460 -70548 -21360 -70386
rect -23262 -71440 -23246 -71406
rect -23146 -71440 -23130 -71406
rect -23004 -71440 -22988 -71406
rect -22888 -71440 -22872 -71406
rect -22746 -71440 -22730 -71406
rect -22630 -71440 -22614 -71406
rect -22488 -71440 -22472 -71406
rect -22372 -71440 -22356 -71406
rect -22230 -71440 -22214 -71406
rect -22114 -71440 -22098 -71406
rect -21972 -71440 -21956 -71406
rect -21856 -71440 -21840 -71406
rect -23342 -71490 -23308 -71474
rect -23342 -71882 -23308 -71866
rect -23084 -71490 -23050 -71474
rect -23084 -71882 -23050 -71866
rect -22826 -71490 -22792 -71474
rect -22826 -71882 -22792 -71866
rect -22568 -71490 -22534 -71474
rect -22568 -71882 -22534 -71866
rect -22310 -71490 -22276 -71474
rect -22310 -71882 -22276 -71866
rect -22052 -71490 -22018 -71474
rect -22052 -71882 -22018 -71866
rect -21794 -71490 -21760 -71474
rect -21794 -71882 -21760 -71866
rect -23262 -71950 -23246 -71916
rect -23146 -71950 -23130 -71916
rect -23004 -71950 -22988 -71916
rect -22888 -71950 -22872 -71916
rect -22746 -71950 -22730 -71916
rect -22630 -71950 -22614 -71916
rect -22488 -71950 -22472 -71916
rect -22372 -71950 -22356 -71916
rect -22230 -71950 -22214 -71916
rect -22114 -71950 -22098 -71916
rect -21972 -71950 -21956 -71916
rect -21856 -71950 -21840 -71916
rect -24072 -72387 -24043 -72353
rect -24009 -72387 -23951 -72353
rect -23917 -72387 -23859 -72353
rect -23825 -72387 -23796 -72353
rect -27928 -72467 -27912 -72433
rect -27878 -72467 -27862 -72433
rect -27928 -72501 -27862 -72467
rect -27928 -72535 -27912 -72501
rect -27878 -72528 -27862 -72501
rect -24008 -72433 -23962 -72387
rect -24008 -72467 -23996 -72433
rect -24008 -72501 -23962 -72467
rect -27928 -72547 -27902 -72535
rect -27908 -72576 -27902 -72547
rect -24008 -72535 -23996 -72501
rect -24008 -72551 -23962 -72535
rect -23928 -72433 -23862 -72421
rect -23684 -72430 -23584 -72268
rect -21460 -72430 -21360 -72268
rect -19684 -70548 -19584 -70386
rect -17460 -70548 -17360 -70386
rect -19262 -71440 -19246 -71406
rect -19146 -71440 -19130 -71406
rect -19004 -71440 -18988 -71406
rect -18888 -71440 -18872 -71406
rect -18746 -71440 -18730 -71406
rect -18630 -71440 -18614 -71406
rect -18488 -71440 -18472 -71406
rect -18372 -71440 -18356 -71406
rect -18230 -71440 -18214 -71406
rect -18114 -71440 -18098 -71406
rect -17972 -71440 -17956 -71406
rect -17856 -71440 -17840 -71406
rect -19342 -71490 -19308 -71474
rect -19342 -71882 -19308 -71866
rect -19084 -71490 -19050 -71474
rect -19084 -71882 -19050 -71866
rect -18826 -71490 -18792 -71474
rect -18826 -71882 -18792 -71866
rect -18568 -71490 -18534 -71474
rect -18568 -71882 -18534 -71866
rect -18310 -71490 -18276 -71474
rect -18310 -71882 -18276 -71866
rect -18052 -71490 -18018 -71474
rect -18052 -71882 -18018 -71866
rect -17794 -71490 -17760 -71474
rect -17794 -71882 -17760 -71866
rect -19262 -71950 -19246 -71916
rect -19146 -71950 -19130 -71916
rect -19004 -71950 -18988 -71916
rect -18888 -71950 -18872 -71916
rect -18746 -71950 -18730 -71916
rect -18630 -71950 -18614 -71916
rect -18488 -71950 -18472 -71916
rect -18372 -71950 -18356 -71916
rect -18230 -71950 -18214 -71916
rect -18114 -71950 -18098 -71916
rect -17972 -71950 -17956 -71916
rect -17856 -71950 -17840 -71916
rect -20072 -72387 -20043 -72353
rect -20009 -72387 -19951 -72353
rect -19917 -72387 -19859 -72353
rect -19825 -72387 -19796 -72353
rect -23928 -72467 -23912 -72433
rect -23878 -72467 -23862 -72433
rect -23928 -72501 -23862 -72467
rect -23928 -72535 -23912 -72501
rect -23878 -72528 -23862 -72501
rect -20008 -72433 -19962 -72387
rect -20008 -72467 -19996 -72433
rect -20008 -72501 -19962 -72467
rect -23928 -72547 -23902 -72535
rect -23908 -72576 -23902 -72547
rect -20008 -72535 -19996 -72501
rect -20008 -72551 -19962 -72535
rect -19928 -72433 -19862 -72421
rect -19684 -72430 -19584 -72268
rect -17460 -72430 -17360 -72268
rect -15684 -70548 -15584 -70386
rect -13460 -70548 -13360 -70386
rect -15262 -71440 -15246 -71406
rect -15146 -71440 -15130 -71406
rect -15004 -71440 -14988 -71406
rect -14888 -71440 -14872 -71406
rect -14746 -71440 -14730 -71406
rect -14630 -71440 -14614 -71406
rect -14488 -71440 -14472 -71406
rect -14372 -71440 -14356 -71406
rect -14230 -71440 -14214 -71406
rect -14114 -71440 -14098 -71406
rect -13972 -71440 -13956 -71406
rect -13856 -71440 -13840 -71406
rect -15342 -71490 -15308 -71474
rect -15342 -71882 -15308 -71866
rect -15084 -71490 -15050 -71474
rect -15084 -71882 -15050 -71866
rect -14826 -71490 -14792 -71474
rect -14826 -71882 -14792 -71866
rect -14568 -71490 -14534 -71474
rect -14568 -71882 -14534 -71866
rect -14310 -71490 -14276 -71474
rect -14310 -71882 -14276 -71866
rect -14052 -71490 -14018 -71474
rect -14052 -71882 -14018 -71866
rect -13794 -71490 -13760 -71474
rect -13794 -71882 -13760 -71866
rect -15262 -71950 -15246 -71916
rect -15146 -71950 -15130 -71916
rect -15004 -71950 -14988 -71916
rect -14888 -71950 -14872 -71916
rect -14746 -71950 -14730 -71916
rect -14630 -71950 -14614 -71916
rect -14488 -71950 -14472 -71916
rect -14372 -71950 -14356 -71916
rect -14230 -71950 -14214 -71916
rect -14114 -71950 -14098 -71916
rect -13972 -71950 -13956 -71916
rect -13856 -71950 -13840 -71916
rect -16072 -72387 -16043 -72353
rect -16009 -72387 -15951 -72353
rect -15917 -72387 -15859 -72353
rect -15825 -72387 -15796 -72353
rect -19928 -72467 -19912 -72433
rect -19878 -72467 -19862 -72433
rect -19928 -72501 -19862 -72467
rect -19928 -72535 -19912 -72501
rect -19878 -72528 -19862 -72501
rect -16008 -72433 -15962 -72387
rect -16008 -72467 -15996 -72433
rect -16008 -72501 -15962 -72467
rect -19928 -72547 -19902 -72535
rect -19908 -72576 -19902 -72547
rect -16008 -72535 -15996 -72501
rect -16008 -72551 -15962 -72535
rect -15928 -72433 -15862 -72421
rect -15684 -72430 -15584 -72268
rect -13460 -72430 -13360 -72268
rect -11684 -70548 -11584 -70386
rect -9460 -70548 -9360 -70386
rect -11262 -71440 -11246 -71406
rect -11146 -71440 -11130 -71406
rect -11004 -71440 -10988 -71406
rect -10888 -71440 -10872 -71406
rect -10746 -71440 -10730 -71406
rect -10630 -71440 -10614 -71406
rect -10488 -71440 -10472 -71406
rect -10372 -71440 -10356 -71406
rect -10230 -71440 -10214 -71406
rect -10114 -71440 -10098 -71406
rect -9972 -71440 -9956 -71406
rect -9856 -71440 -9840 -71406
rect -11342 -71490 -11308 -71474
rect -11342 -71882 -11308 -71866
rect -11084 -71490 -11050 -71474
rect -11084 -71882 -11050 -71866
rect -10826 -71490 -10792 -71474
rect -10826 -71882 -10792 -71866
rect -10568 -71490 -10534 -71474
rect -10568 -71882 -10534 -71866
rect -10310 -71490 -10276 -71474
rect -10310 -71882 -10276 -71866
rect -10052 -71490 -10018 -71474
rect -10052 -71882 -10018 -71866
rect -9794 -71490 -9760 -71474
rect -9794 -71882 -9760 -71866
rect -11262 -71950 -11246 -71916
rect -11146 -71950 -11130 -71916
rect -11004 -71950 -10988 -71916
rect -10888 -71950 -10872 -71916
rect -10746 -71950 -10730 -71916
rect -10630 -71950 -10614 -71916
rect -10488 -71950 -10472 -71916
rect -10372 -71950 -10356 -71916
rect -10230 -71950 -10214 -71916
rect -10114 -71950 -10098 -71916
rect -9972 -71950 -9956 -71916
rect -9856 -71950 -9840 -71916
rect -12072 -72387 -12043 -72353
rect -12009 -72387 -11951 -72353
rect -11917 -72387 -11859 -72353
rect -11825 -72387 -11796 -72353
rect -15928 -72467 -15912 -72433
rect -15878 -72467 -15862 -72433
rect -15928 -72501 -15862 -72467
rect -15928 -72535 -15912 -72501
rect -15878 -72528 -15862 -72501
rect -12008 -72433 -11962 -72387
rect -12008 -72467 -11996 -72433
rect -12008 -72501 -11962 -72467
rect -15928 -72547 -15902 -72535
rect -15908 -72576 -15902 -72547
rect -12008 -72535 -11996 -72501
rect -12008 -72551 -11962 -72535
rect -11928 -72433 -11862 -72421
rect -11684 -72430 -11584 -72268
rect -9460 -72430 -9360 -72268
rect -7684 -70548 -7584 -70386
rect -5460 -70548 -5360 -70386
rect -7262 -71440 -7246 -71406
rect -7146 -71440 -7130 -71406
rect -7004 -71440 -6988 -71406
rect -6888 -71440 -6872 -71406
rect -6746 -71440 -6730 -71406
rect -6630 -71440 -6614 -71406
rect -6488 -71440 -6472 -71406
rect -6372 -71440 -6356 -71406
rect -6230 -71440 -6214 -71406
rect -6114 -71440 -6098 -71406
rect -5972 -71440 -5956 -71406
rect -5856 -71440 -5840 -71406
rect -7342 -71490 -7308 -71474
rect -7342 -71882 -7308 -71866
rect -7084 -71490 -7050 -71474
rect -7084 -71882 -7050 -71866
rect -6826 -71490 -6792 -71474
rect -6826 -71882 -6792 -71866
rect -6568 -71490 -6534 -71474
rect -6568 -71882 -6534 -71866
rect -6310 -71490 -6276 -71474
rect -6310 -71882 -6276 -71866
rect -6052 -71490 -6018 -71474
rect -6052 -71882 -6018 -71866
rect -5794 -71490 -5760 -71474
rect -5794 -71882 -5760 -71866
rect -7262 -71950 -7246 -71916
rect -7146 -71950 -7130 -71916
rect -7004 -71950 -6988 -71916
rect -6888 -71950 -6872 -71916
rect -6746 -71950 -6730 -71916
rect -6630 -71950 -6614 -71916
rect -6488 -71950 -6472 -71916
rect -6372 -71950 -6356 -71916
rect -6230 -71950 -6214 -71916
rect -6114 -71950 -6098 -71916
rect -5972 -71950 -5956 -71916
rect -5856 -71950 -5840 -71916
rect -8072 -72387 -8043 -72353
rect -8009 -72387 -7951 -72353
rect -7917 -72387 -7859 -72353
rect -7825 -72387 -7796 -72353
rect -11928 -72467 -11912 -72433
rect -11878 -72467 -11862 -72433
rect -11928 -72501 -11862 -72467
rect -11928 -72535 -11912 -72501
rect -11878 -72528 -11862 -72501
rect -8008 -72433 -7962 -72387
rect -8008 -72467 -7996 -72433
rect -8008 -72501 -7962 -72467
rect -11928 -72547 -11902 -72535
rect -11908 -72576 -11902 -72547
rect -8008 -72535 -7996 -72501
rect -8008 -72551 -7962 -72535
rect -7928 -72433 -7862 -72421
rect -7684 -72430 -7584 -72268
rect -5460 -72430 -5360 -72268
rect -3684 -70548 -3584 -70386
rect -1460 -70548 -1360 -70386
rect -3262 -71440 -3246 -71406
rect -3146 -71440 -3130 -71406
rect -3004 -71440 -2988 -71406
rect -2888 -71440 -2872 -71406
rect -2746 -71440 -2730 -71406
rect -2630 -71440 -2614 -71406
rect -2488 -71440 -2472 -71406
rect -2372 -71440 -2356 -71406
rect -2230 -71440 -2214 -71406
rect -2114 -71440 -2098 -71406
rect -1972 -71440 -1956 -71406
rect -1856 -71440 -1840 -71406
rect -3342 -71490 -3308 -71474
rect -3342 -71882 -3308 -71866
rect -3084 -71490 -3050 -71474
rect -3084 -71882 -3050 -71866
rect -2826 -71490 -2792 -71474
rect -2826 -71882 -2792 -71866
rect -2568 -71490 -2534 -71474
rect -2568 -71882 -2534 -71866
rect -2310 -71490 -2276 -71474
rect -2310 -71882 -2276 -71866
rect -2052 -71490 -2018 -71474
rect -2052 -71882 -2018 -71866
rect -1794 -71490 -1760 -71474
rect -1794 -71882 -1760 -71866
rect -3262 -71950 -3246 -71916
rect -3146 -71950 -3130 -71916
rect -3004 -71950 -2988 -71916
rect -2888 -71950 -2872 -71916
rect -2746 -71950 -2730 -71916
rect -2630 -71950 -2614 -71916
rect -2488 -71950 -2472 -71916
rect -2372 -71950 -2356 -71916
rect -2230 -71950 -2214 -71916
rect -2114 -71950 -2098 -71916
rect -1972 -71950 -1956 -71916
rect -1856 -71950 -1840 -71916
rect -4072 -72387 -4043 -72353
rect -4009 -72387 -3951 -72353
rect -3917 -72387 -3859 -72353
rect -3825 -72387 -3796 -72353
rect -7928 -72467 -7912 -72433
rect -7878 -72467 -7862 -72433
rect -7928 -72501 -7862 -72467
rect -7928 -72535 -7912 -72501
rect -7878 -72528 -7862 -72501
rect -4008 -72433 -3962 -72387
rect -4008 -72467 -3996 -72433
rect -4008 -72501 -3962 -72467
rect -7928 -72547 -7902 -72535
rect -7908 -72576 -7902 -72547
rect -4008 -72535 -3996 -72501
rect -4008 -72551 -3962 -72535
rect -3928 -72433 -3862 -72421
rect -3684 -72430 -3584 -72268
rect -1460 -72430 -1360 -72268
rect 316 -70548 416 -70386
rect 2540 -70548 2640 -70386
rect 738 -71440 754 -71406
rect 854 -71440 870 -71406
rect 996 -71440 1012 -71406
rect 1112 -71440 1128 -71406
rect 1254 -71440 1270 -71406
rect 1370 -71440 1386 -71406
rect 1512 -71440 1528 -71406
rect 1628 -71440 1644 -71406
rect 1770 -71440 1786 -71406
rect 1886 -71440 1902 -71406
rect 2028 -71440 2044 -71406
rect 2144 -71440 2160 -71406
rect 658 -71490 692 -71474
rect 658 -71882 692 -71866
rect 916 -71490 950 -71474
rect 916 -71882 950 -71866
rect 1174 -71490 1208 -71474
rect 1174 -71882 1208 -71866
rect 1432 -71490 1466 -71474
rect 1432 -71882 1466 -71866
rect 1690 -71490 1724 -71474
rect 1690 -71882 1724 -71866
rect 1948 -71490 1982 -71474
rect 1948 -71882 1982 -71866
rect 2206 -71490 2240 -71474
rect 2206 -71882 2240 -71866
rect 738 -71950 754 -71916
rect 854 -71950 870 -71916
rect 996 -71950 1012 -71916
rect 1112 -71950 1128 -71916
rect 1254 -71950 1270 -71916
rect 1370 -71950 1386 -71916
rect 1512 -71950 1528 -71916
rect 1628 -71950 1644 -71916
rect 1770 -71950 1786 -71916
rect 1886 -71950 1902 -71916
rect 2028 -71950 2044 -71916
rect 2144 -71950 2160 -71916
rect -72 -72387 -43 -72353
rect -9 -72387 49 -72353
rect 83 -72387 141 -72353
rect 175 -72387 204 -72353
rect -3928 -72467 -3912 -72433
rect -3878 -72467 -3862 -72433
rect -3928 -72501 -3862 -72467
rect -3928 -72535 -3912 -72501
rect -3878 -72528 -3862 -72501
rect -8 -72433 38 -72387
rect -8 -72467 4 -72433
rect -8 -72501 38 -72467
rect -3928 -72547 -3902 -72535
rect -3908 -72576 -3902 -72547
rect -8 -72535 4 -72501
rect -8 -72551 38 -72535
rect 72 -72433 138 -72421
rect 316 -72430 416 -72268
rect 2540 -72430 2640 -72268
rect 4316 -70548 4416 -70386
rect 6540 -70548 6640 -70386
rect 4738 -71440 4754 -71406
rect 4854 -71440 4870 -71406
rect 4996 -71440 5012 -71406
rect 5112 -71440 5128 -71406
rect 5254 -71440 5270 -71406
rect 5370 -71440 5386 -71406
rect 5512 -71440 5528 -71406
rect 5628 -71440 5644 -71406
rect 5770 -71440 5786 -71406
rect 5886 -71440 5902 -71406
rect 6028 -71440 6044 -71406
rect 6144 -71440 6160 -71406
rect 4658 -71490 4692 -71474
rect 4658 -71882 4692 -71866
rect 4916 -71490 4950 -71474
rect 4916 -71882 4950 -71866
rect 5174 -71490 5208 -71474
rect 5174 -71882 5208 -71866
rect 5432 -71490 5466 -71474
rect 5432 -71882 5466 -71866
rect 5690 -71490 5724 -71474
rect 5690 -71882 5724 -71866
rect 5948 -71490 5982 -71474
rect 5948 -71882 5982 -71866
rect 6206 -71490 6240 -71474
rect 6206 -71882 6240 -71866
rect 4738 -71950 4754 -71916
rect 4854 -71950 4870 -71916
rect 4996 -71950 5012 -71916
rect 5112 -71950 5128 -71916
rect 5254 -71950 5270 -71916
rect 5370 -71950 5386 -71916
rect 5512 -71950 5528 -71916
rect 5628 -71950 5644 -71916
rect 5770 -71950 5786 -71916
rect 5886 -71950 5902 -71916
rect 6028 -71950 6044 -71916
rect 6144 -71950 6160 -71916
rect 3928 -72387 3957 -72353
rect 3991 -72387 4049 -72353
rect 4083 -72387 4141 -72353
rect 4175 -72387 4204 -72353
rect 72 -72467 88 -72433
rect 122 -72467 138 -72433
rect 72 -72501 138 -72467
rect 72 -72535 88 -72501
rect 122 -72528 138 -72501
rect 3992 -72433 4038 -72387
rect 3992 -72467 4004 -72433
rect 3992 -72501 4038 -72467
rect 72 -72547 98 -72535
rect 92 -72576 98 -72547
rect 3992 -72535 4004 -72501
rect 3992 -72551 4038 -72535
rect 4072 -72433 4138 -72421
rect 4316 -72430 4416 -72268
rect 6540 -72430 6640 -72268
rect 4072 -72467 4088 -72433
rect 4122 -72467 4138 -72433
rect 4072 -72501 4138 -72467
rect 4072 -72535 4088 -72501
rect 4122 -72528 4138 -72501
rect 4072 -72547 4098 -72535
rect 4092 -72576 4098 -72547
rect -28008 -72586 -27992 -72585
rect -27958 -72586 -27942 -72585
rect -28008 -72633 -28004 -72586
rect -27956 -72633 -27942 -72586
rect -27908 -72667 -27862 -72576
rect -24008 -72586 -23992 -72585
rect -23958 -72586 -23942 -72585
rect -24008 -72633 -24004 -72586
rect -23956 -72633 -23942 -72586
rect -28004 -72685 -27962 -72669
rect -28004 -72719 -27996 -72685
rect -28004 -72753 -27962 -72719
rect -28004 -72787 -27996 -72753
rect -28004 -72821 -27962 -72787
rect -28004 -72855 -27996 -72821
rect -28004 -72897 -27962 -72855
rect -27928 -72685 -27862 -72667
rect -27928 -72719 -27912 -72685
rect -27878 -72719 -27862 -72685
rect -27928 -72753 -27862 -72719
rect -27928 -72787 -27912 -72753
rect -27878 -72787 -27862 -72753
rect -27928 -72821 -27862 -72787
rect -27928 -72855 -27912 -72821
rect -27878 -72855 -27862 -72821
rect -27928 -72863 -27862 -72855
rect -27684 -72828 -27584 -72666
rect -28072 -72931 -28043 -72897
rect -28009 -72931 -27951 -72897
rect -27917 -72931 -27859 -72897
rect -27825 -72931 -27796 -72897
rect -25460 -72828 -25360 -72666
rect -23908 -72667 -23862 -72576
rect -20008 -72586 -19992 -72585
rect -19958 -72586 -19942 -72585
rect -20008 -72633 -20004 -72586
rect -19956 -72633 -19942 -72586
rect -24004 -72685 -23962 -72669
rect -24004 -72719 -23996 -72685
rect -24004 -72753 -23962 -72719
rect -24004 -72787 -23996 -72753
rect -24004 -72821 -23962 -72787
rect -24004 -72855 -23996 -72821
rect -24004 -72897 -23962 -72855
rect -23928 -72685 -23862 -72667
rect -23928 -72719 -23912 -72685
rect -23878 -72719 -23862 -72685
rect -23928 -72753 -23862 -72719
rect -23928 -72787 -23912 -72753
rect -23878 -72787 -23862 -72753
rect -23928 -72821 -23862 -72787
rect -23928 -72855 -23912 -72821
rect -23878 -72855 -23862 -72821
rect -23928 -72863 -23862 -72855
rect -23684 -72828 -23584 -72666
rect -27257 -73264 -27241 -73230
rect -27141 -73264 -27125 -73230
rect -26999 -73264 -26983 -73230
rect -26883 -73264 -26867 -73230
rect -26741 -73264 -26725 -73230
rect -26625 -73264 -26609 -73230
rect -26483 -73264 -26467 -73230
rect -26367 -73264 -26351 -73230
rect -26225 -73264 -26209 -73230
rect -26109 -73264 -26093 -73230
rect -25967 -73264 -25951 -73230
rect -25851 -73264 -25835 -73230
rect -27337 -73323 -27303 -73307
rect -27337 -73715 -27303 -73699
rect -27079 -73323 -27045 -73307
rect -27079 -73715 -27045 -73699
rect -26821 -73323 -26787 -73307
rect -26821 -73715 -26787 -73699
rect -26563 -73323 -26529 -73307
rect -26563 -73715 -26529 -73699
rect -26305 -73323 -26271 -73307
rect -26305 -73715 -26271 -73699
rect -26047 -73323 -26013 -73307
rect -26047 -73715 -26013 -73699
rect -25789 -73323 -25755 -73307
rect -25789 -73715 -25755 -73699
rect -27257 -73792 -27241 -73758
rect -27141 -73792 -27125 -73758
rect -26999 -73792 -26983 -73758
rect -26883 -73792 -26867 -73758
rect -26741 -73792 -26725 -73758
rect -26625 -73792 -26609 -73758
rect -26483 -73792 -26467 -73758
rect -26367 -73792 -26351 -73758
rect -26225 -73792 -26209 -73758
rect -26109 -73792 -26093 -73758
rect -25967 -73792 -25951 -73758
rect -25851 -73792 -25835 -73758
rect -27257 -74124 -27241 -74090
rect -27141 -74124 -27125 -74090
rect -26999 -74124 -26983 -74090
rect -26883 -74124 -26867 -74090
rect -26741 -74124 -26725 -74090
rect -26625 -74124 -26609 -74090
rect -26483 -74124 -26467 -74090
rect -26367 -74124 -26351 -74090
rect -26225 -74124 -26209 -74090
rect -26109 -74124 -26093 -74090
rect -25967 -74124 -25951 -74090
rect -25851 -74124 -25835 -74090
rect -27337 -74183 -27303 -74167
rect -27337 -74575 -27303 -74559
rect -27079 -74183 -27045 -74167
rect -27079 -74575 -27045 -74559
rect -26821 -74183 -26787 -74167
rect -26821 -74575 -26787 -74559
rect -26563 -74183 -26529 -74167
rect -26563 -74575 -26529 -74559
rect -26305 -74183 -26271 -74167
rect -26305 -74575 -26271 -74559
rect -26047 -74183 -26013 -74167
rect -26047 -74575 -26013 -74559
rect -25789 -74183 -25755 -74167
rect -25789 -74575 -25755 -74559
rect -27257 -74652 -27241 -74618
rect -27141 -74652 -27125 -74618
rect -26999 -74652 -26983 -74618
rect -26883 -74652 -26867 -74618
rect -26741 -74652 -26725 -74618
rect -26625 -74652 -26609 -74618
rect -26483 -74652 -26467 -74618
rect -26367 -74652 -26351 -74618
rect -26225 -74652 -26209 -74618
rect -26109 -74652 -26093 -74618
rect -25967 -74652 -25951 -74618
rect -25851 -74652 -25835 -74618
rect -27684 -75770 -27584 -75608
rect -24072 -72931 -24043 -72897
rect -24009 -72931 -23951 -72897
rect -23917 -72931 -23859 -72897
rect -23825 -72931 -23796 -72897
rect -25460 -75770 -25360 -75608
rect -21460 -72828 -21360 -72666
rect -19908 -72667 -19862 -72576
rect -16008 -72586 -15992 -72585
rect -15958 -72586 -15942 -72585
rect -16008 -72633 -16004 -72586
rect -15956 -72633 -15942 -72586
rect -20004 -72685 -19962 -72669
rect -20004 -72719 -19996 -72685
rect -20004 -72753 -19962 -72719
rect -20004 -72787 -19996 -72753
rect -20004 -72821 -19962 -72787
rect -20004 -72855 -19996 -72821
rect -20004 -72897 -19962 -72855
rect -19928 -72685 -19862 -72667
rect -19928 -72719 -19912 -72685
rect -19878 -72719 -19862 -72685
rect -19928 -72753 -19862 -72719
rect -19928 -72787 -19912 -72753
rect -19878 -72787 -19862 -72753
rect -19928 -72821 -19862 -72787
rect -19928 -72855 -19912 -72821
rect -19878 -72855 -19862 -72821
rect -19928 -72863 -19862 -72855
rect -19684 -72828 -19584 -72666
rect -23257 -73264 -23241 -73230
rect -23141 -73264 -23125 -73230
rect -22999 -73264 -22983 -73230
rect -22883 -73264 -22867 -73230
rect -22741 -73264 -22725 -73230
rect -22625 -73264 -22609 -73230
rect -22483 -73264 -22467 -73230
rect -22367 -73264 -22351 -73230
rect -22225 -73264 -22209 -73230
rect -22109 -73264 -22093 -73230
rect -21967 -73264 -21951 -73230
rect -21851 -73264 -21835 -73230
rect -23337 -73323 -23303 -73307
rect -23337 -73715 -23303 -73699
rect -23079 -73323 -23045 -73307
rect -23079 -73715 -23045 -73699
rect -22821 -73323 -22787 -73307
rect -22821 -73715 -22787 -73699
rect -22563 -73323 -22529 -73307
rect -22563 -73715 -22529 -73699
rect -22305 -73323 -22271 -73307
rect -22305 -73715 -22271 -73699
rect -22047 -73323 -22013 -73307
rect -22047 -73715 -22013 -73699
rect -21789 -73323 -21755 -73307
rect -21789 -73715 -21755 -73699
rect -23257 -73792 -23241 -73758
rect -23141 -73792 -23125 -73758
rect -22999 -73792 -22983 -73758
rect -22883 -73792 -22867 -73758
rect -22741 -73792 -22725 -73758
rect -22625 -73792 -22609 -73758
rect -22483 -73792 -22467 -73758
rect -22367 -73792 -22351 -73758
rect -22225 -73792 -22209 -73758
rect -22109 -73792 -22093 -73758
rect -21967 -73792 -21951 -73758
rect -21851 -73792 -21835 -73758
rect -23257 -74124 -23241 -74090
rect -23141 -74124 -23125 -74090
rect -22999 -74124 -22983 -74090
rect -22883 -74124 -22867 -74090
rect -22741 -74124 -22725 -74090
rect -22625 -74124 -22609 -74090
rect -22483 -74124 -22467 -74090
rect -22367 -74124 -22351 -74090
rect -22225 -74124 -22209 -74090
rect -22109 -74124 -22093 -74090
rect -21967 -74124 -21951 -74090
rect -21851 -74124 -21835 -74090
rect -23337 -74183 -23303 -74167
rect -23337 -74575 -23303 -74559
rect -23079 -74183 -23045 -74167
rect -23079 -74575 -23045 -74559
rect -22821 -74183 -22787 -74167
rect -22821 -74575 -22787 -74559
rect -22563 -74183 -22529 -74167
rect -22563 -74575 -22529 -74559
rect -22305 -74183 -22271 -74167
rect -22305 -74575 -22271 -74559
rect -22047 -74183 -22013 -74167
rect -22047 -74575 -22013 -74559
rect -21789 -74183 -21755 -74167
rect -21789 -74575 -21755 -74559
rect -23257 -74652 -23241 -74618
rect -23141 -74652 -23125 -74618
rect -22999 -74652 -22983 -74618
rect -22883 -74652 -22867 -74618
rect -22741 -74652 -22725 -74618
rect -22625 -74652 -22609 -74618
rect -22483 -74652 -22467 -74618
rect -22367 -74652 -22351 -74618
rect -22225 -74652 -22209 -74618
rect -22109 -74652 -22093 -74618
rect -21967 -74652 -21951 -74618
rect -21851 -74652 -21835 -74618
rect -23684 -75770 -23584 -75608
rect -20072 -72931 -20043 -72897
rect -20009 -72931 -19951 -72897
rect -19917 -72931 -19859 -72897
rect -19825 -72931 -19796 -72897
rect -21460 -75770 -21360 -75608
rect -17460 -72828 -17360 -72666
rect -15908 -72667 -15862 -72576
rect -12008 -72586 -11992 -72585
rect -11958 -72586 -11942 -72585
rect -12008 -72633 -12004 -72586
rect -11956 -72633 -11942 -72586
rect -16004 -72685 -15962 -72669
rect -16004 -72719 -15996 -72685
rect -16004 -72753 -15962 -72719
rect -16004 -72787 -15996 -72753
rect -16004 -72821 -15962 -72787
rect -16004 -72855 -15996 -72821
rect -16004 -72897 -15962 -72855
rect -15928 -72685 -15862 -72667
rect -15928 -72719 -15912 -72685
rect -15878 -72719 -15862 -72685
rect -15928 -72753 -15862 -72719
rect -15928 -72787 -15912 -72753
rect -15878 -72787 -15862 -72753
rect -15928 -72821 -15862 -72787
rect -15928 -72855 -15912 -72821
rect -15878 -72855 -15862 -72821
rect -15928 -72863 -15862 -72855
rect -15684 -72828 -15584 -72666
rect -19257 -73264 -19241 -73230
rect -19141 -73264 -19125 -73230
rect -18999 -73264 -18983 -73230
rect -18883 -73264 -18867 -73230
rect -18741 -73264 -18725 -73230
rect -18625 -73264 -18609 -73230
rect -18483 -73264 -18467 -73230
rect -18367 -73264 -18351 -73230
rect -18225 -73264 -18209 -73230
rect -18109 -73264 -18093 -73230
rect -17967 -73264 -17951 -73230
rect -17851 -73264 -17835 -73230
rect -19337 -73323 -19303 -73307
rect -19337 -73715 -19303 -73699
rect -19079 -73323 -19045 -73307
rect -19079 -73715 -19045 -73699
rect -18821 -73323 -18787 -73307
rect -18821 -73715 -18787 -73699
rect -18563 -73323 -18529 -73307
rect -18563 -73715 -18529 -73699
rect -18305 -73323 -18271 -73307
rect -18305 -73715 -18271 -73699
rect -18047 -73323 -18013 -73307
rect -18047 -73715 -18013 -73699
rect -17789 -73323 -17755 -73307
rect -17789 -73715 -17755 -73699
rect -19257 -73792 -19241 -73758
rect -19141 -73792 -19125 -73758
rect -18999 -73792 -18983 -73758
rect -18883 -73792 -18867 -73758
rect -18741 -73792 -18725 -73758
rect -18625 -73792 -18609 -73758
rect -18483 -73792 -18467 -73758
rect -18367 -73792 -18351 -73758
rect -18225 -73792 -18209 -73758
rect -18109 -73792 -18093 -73758
rect -17967 -73792 -17951 -73758
rect -17851 -73792 -17835 -73758
rect -19257 -74124 -19241 -74090
rect -19141 -74124 -19125 -74090
rect -18999 -74124 -18983 -74090
rect -18883 -74124 -18867 -74090
rect -18741 -74124 -18725 -74090
rect -18625 -74124 -18609 -74090
rect -18483 -74124 -18467 -74090
rect -18367 -74124 -18351 -74090
rect -18225 -74124 -18209 -74090
rect -18109 -74124 -18093 -74090
rect -17967 -74124 -17951 -74090
rect -17851 -74124 -17835 -74090
rect -19337 -74183 -19303 -74167
rect -19337 -74575 -19303 -74559
rect -19079 -74183 -19045 -74167
rect -19079 -74575 -19045 -74559
rect -18821 -74183 -18787 -74167
rect -18821 -74575 -18787 -74559
rect -18563 -74183 -18529 -74167
rect -18563 -74575 -18529 -74559
rect -18305 -74183 -18271 -74167
rect -18305 -74575 -18271 -74559
rect -18047 -74183 -18013 -74167
rect -18047 -74575 -18013 -74559
rect -17789 -74183 -17755 -74167
rect -17789 -74575 -17755 -74559
rect -19257 -74652 -19241 -74618
rect -19141 -74652 -19125 -74618
rect -18999 -74652 -18983 -74618
rect -18883 -74652 -18867 -74618
rect -18741 -74652 -18725 -74618
rect -18625 -74652 -18609 -74618
rect -18483 -74652 -18467 -74618
rect -18367 -74652 -18351 -74618
rect -18225 -74652 -18209 -74618
rect -18109 -74652 -18093 -74618
rect -17967 -74652 -17951 -74618
rect -17851 -74652 -17835 -74618
rect -19684 -75770 -19584 -75608
rect -16072 -72931 -16043 -72897
rect -16009 -72931 -15951 -72897
rect -15917 -72931 -15859 -72897
rect -15825 -72931 -15796 -72897
rect -17460 -75770 -17360 -75608
rect -13460 -72828 -13360 -72666
rect -11908 -72667 -11862 -72576
rect -8008 -72586 -7992 -72585
rect -7958 -72586 -7942 -72585
rect -8008 -72633 -8004 -72586
rect -7956 -72633 -7942 -72586
rect -12004 -72685 -11962 -72669
rect -12004 -72719 -11996 -72685
rect -12004 -72753 -11962 -72719
rect -12004 -72787 -11996 -72753
rect -12004 -72821 -11962 -72787
rect -12004 -72855 -11996 -72821
rect -12004 -72897 -11962 -72855
rect -11928 -72685 -11862 -72667
rect -11928 -72719 -11912 -72685
rect -11878 -72719 -11862 -72685
rect -11928 -72753 -11862 -72719
rect -11928 -72787 -11912 -72753
rect -11878 -72787 -11862 -72753
rect -11928 -72821 -11862 -72787
rect -11928 -72855 -11912 -72821
rect -11878 -72855 -11862 -72821
rect -11928 -72863 -11862 -72855
rect -11684 -72828 -11584 -72666
rect -15257 -73264 -15241 -73230
rect -15141 -73264 -15125 -73230
rect -14999 -73264 -14983 -73230
rect -14883 -73264 -14867 -73230
rect -14741 -73264 -14725 -73230
rect -14625 -73264 -14609 -73230
rect -14483 -73264 -14467 -73230
rect -14367 -73264 -14351 -73230
rect -14225 -73264 -14209 -73230
rect -14109 -73264 -14093 -73230
rect -13967 -73264 -13951 -73230
rect -13851 -73264 -13835 -73230
rect -15337 -73323 -15303 -73307
rect -15337 -73715 -15303 -73699
rect -15079 -73323 -15045 -73307
rect -15079 -73715 -15045 -73699
rect -14821 -73323 -14787 -73307
rect -14821 -73715 -14787 -73699
rect -14563 -73323 -14529 -73307
rect -14563 -73715 -14529 -73699
rect -14305 -73323 -14271 -73307
rect -14305 -73715 -14271 -73699
rect -14047 -73323 -14013 -73307
rect -14047 -73715 -14013 -73699
rect -13789 -73323 -13755 -73307
rect -13789 -73715 -13755 -73699
rect -15257 -73792 -15241 -73758
rect -15141 -73792 -15125 -73758
rect -14999 -73792 -14983 -73758
rect -14883 -73792 -14867 -73758
rect -14741 -73792 -14725 -73758
rect -14625 -73792 -14609 -73758
rect -14483 -73792 -14467 -73758
rect -14367 -73792 -14351 -73758
rect -14225 -73792 -14209 -73758
rect -14109 -73792 -14093 -73758
rect -13967 -73792 -13951 -73758
rect -13851 -73792 -13835 -73758
rect -15257 -74124 -15241 -74090
rect -15141 -74124 -15125 -74090
rect -14999 -74124 -14983 -74090
rect -14883 -74124 -14867 -74090
rect -14741 -74124 -14725 -74090
rect -14625 -74124 -14609 -74090
rect -14483 -74124 -14467 -74090
rect -14367 -74124 -14351 -74090
rect -14225 -74124 -14209 -74090
rect -14109 -74124 -14093 -74090
rect -13967 -74124 -13951 -74090
rect -13851 -74124 -13835 -74090
rect -15337 -74183 -15303 -74167
rect -15337 -74575 -15303 -74559
rect -15079 -74183 -15045 -74167
rect -15079 -74575 -15045 -74559
rect -14821 -74183 -14787 -74167
rect -14821 -74575 -14787 -74559
rect -14563 -74183 -14529 -74167
rect -14563 -74575 -14529 -74559
rect -14305 -74183 -14271 -74167
rect -14305 -74575 -14271 -74559
rect -14047 -74183 -14013 -74167
rect -14047 -74575 -14013 -74559
rect -13789 -74183 -13755 -74167
rect -13789 -74575 -13755 -74559
rect -15257 -74652 -15241 -74618
rect -15141 -74652 -15125 -74618
rect -14999 -74652 -14983 -74618
rect -14883 -74652 -14867 -74618
rect -14741 -74652 -14725 -74618
rect -14625 -74652 -14609 -74618
rect -14483 -74652 -14467 -74618
rect -14367 -74652 -14351 -74618
rect -14225 -74652 -14209 -74618
rect -14109 -74652 -14093 -74618
rect -13967 -74652 -13951 -74618
rect -13851 -74652 -13835 -74618
rect -15684 -75770 -15584 -75608
rect -12072 -72931 -12043 -72897
rect -12009 -72931 -11951 -72897
rect -11917 -72931 -11859 -72897
rect -11825 -72931 -11796 -72897
rect -13460 -75770 -13360 -75608
rect -9460 -72828 -9360 -72666
rect -7908 -72667 -7862 -72576
rect -4008 -72586 -3992 -72585
rect -3958 -72586 -3942 -72585
rect -4008 -72633 -4004 -72586
rect -3956 -72633 -3942 -72586
rect -8004 -72685 -7962 -72669
rect -8004 -72719 -7996 -72685
rect -8004 -72753 -7962 -72719
rect -8004 -72787 -7996 -72753
rect -8004 -72821 -7962 -72787
rect -8004 -72855 -7996 -72821
rect -8004 -72897 -7962 -72855
rect -7928 -72685 -7862 -72667
rect -7928 -72719 -7912 -72685
rect -7878 -72719 -7862 -72685
rect -7928 -72753 -7862 -72719
rect -7928 -72787 -7912 -72753
rect -7878 -72787 -7862 -72753
rect -7928 -72821 -7862 -72787
rect -7928 -72855 -7912 -72821
rect -7878 -72855 -7862 -72821
rect -7928 -72863 -7862 -72855
rect -7684 -72828 -7584 -72666
rect -11257 -73264 -11241 -73230
rect -11141 -73264 -11125 -73230
rect -10999 -73264 -10983 -73230
rect -10883 -73264 -10867 -73230
rect -10741 -73264 -10725 -73230
rect -10625 -73264 -10609 -73230
rect -10483 -73264 -10467 -73230
rect -10367 -73264 -10351 -73230
rect -10225 -73264 -10209 -73230
rect -10109 -73264 -10093 -73230
rect -9967 -73264 -9951 -73230
rect -9851 -73264 -9835 -73230
rect -11337 -73323 -11303 -73307
rect -11337 -73715 -11303 -73699
rect -11079 -73323 -11045 -73307
rect -11079 -73715 -11045 -73699
rect -10821 -73323 -10787 -73307
rect -10821 -73715 -10787 -73699
rect -10563 -73323 -10529 -73307
rect -10563 -73715 -10529 -73699
rect -10305 -73323 -10271 -73307
rect -10305 -73715 -10271 -73699
rect -10047 -73323 -10013 -73307
rect -10047 -73715 -10013 -73699
rect -9789 -73323 -9755 -73307
rect -9789 -73715 -9755 -73699
rect -11257 -73792 -11241 -73758
rect -11141 -73792 -11125 -73758
rect -10999 -73792 -10983 -73758
rect -10883 -73792 -10867 -73758
rect -10741 -73792 -10725 -73758
rect -10625 -73792 -10609 -73758
rect -10483 -73792 -10467 -73758
rect -10367 -73792 -10351 -73758
rect -10225 -73792 -10209 -73758
rect -10109 -73792 -10093 -73758
rect -9967 -73792 -9951 -73758
rect -9851 -73792 -9835 -73758
rect -11257 -74124 -11241 -74090
rect -11141 -74124 -11125 -74090
rect -10999 -74124 -10983 -74090
rect -10883 -74124 -10867 -74090
rect -10741 -74124 -10725 -74090
rect -10625 -74124 -10609 -74090
rect -10483 -74124 -10467 -74090
rect -10367 -74124 -10351 -74090
rect -10225 -74124 -10209 -74090
rect -10109 -74124 -10093 -74090
rect -9967 -74124 -9951 -74090
rect -9851 -74124 -9835 -74090
rect -11337 -74183 -11303 -74167
rect -11337 -74575 -11303 -74559
rect -11079 -74183 -11045 -74167
rect -11079 -74575 -11045 -74559
rect -10821 -74183 -10787 -74167
rect -10821 -74575 -10787 -74559
rect -10563 -74183 -10529 -74167
rect -10563 -74575 -10529 -74559
rect -10305 -74183 -10271 -74167
rect -10305 -74575 -10271 -74559
rect -10047 -74183 -10013 -74167
rect -10047 -74575 -10013 -74559
rect -9789 -74183 -9755 -74167
rect -9789 -74575 -9755 -74559
rect -11257 -74652 -11241 -74618
rect -11141 -74652 -11125 -74618
rect -10999 -74652 -10983 -74618
rect -10883 -74652 -10867 -74618
rect -10741 -74652 -10725 -74618
rect -10625 -74652 -10609 -74618
rect -10483 -74652 -10467 -74618
rect -10367 -74652 -10351 -74618
rect -10225 -74652 -10209 -74618
rect -10109 -74652 -10093 -74618
rect -9967 -74652 -9951 -74618
rect -9851 -74652 -9835 -74618
rect -11684 -75770 -11584 -75608
rect -8072 -72931 -8043 -72897
rect -8009 -72931 -7951 -72897
rect -7917 -72931 -7859 -72897
rect -7825 -72931 -7796 -72897
rect -9460 -75770 -9360 -75608
rect -5460 -72828 -5360 -72666
rect -3908 -72667 -3862 -72576
rect -8 -72586 8 -72585
rect 42 -72586 58 -72585
rect -8 -72633 -4 -72586
rect 44 -72633 58 -72586
rect -4004 -72685 -3962 -72669
rect -4004 -72719 -3996 -72685
rect -4004 -72753 -3962 -72719
rect -4004 -72787 -3996 -72753
rect -4004 -72821 -3962 -72787
rect -4004 -72855 -3996 -72821
rect -4004 -72897 -3962 -72855
rect -3928 -72685 -3862 -72667
rect -3928 -72719 -3912 -72685
rect -3878 -72719 -3862 -72685
rect -3928 -72753 -3862 -72719
rect -3928 -72787 -3912 -72753
rect -3878 -72787 -3862 -72753
rect -3928 -72821 -3862 -72787
rect -3928 -72855 -3912 -72821
rect -3878 -72855 -3862 -72821
rect -3928 -72863 -3862 -72855
rect -3684 -72828 -3584 -72666
rect -7257 -73264 -7241 -73230
rect -7141 -73264 -7125 -73230
rect -6999 -73264 -6983 -73230
rect -6883 -73264 -6867 -73230
rect -6741 -73264 -6725 -73230
rect -6625 -73264 -6609 -73230
rect -6483 -73264 -6467 -73230
rect -6367 -73264 -6351 -73230
rect -6225 -73264 -6209 -73230
rect -6109 -73264 -6093 -73230
rect -5967 -73264 -5951 -73230
rect -5851 -73264 -5835 -73230
rect -7337 -73323 -7303 -73307
rect -7337 -73715 -7303 -73699
rect -7079 -73323 -7045 -73307
rect -7079 -73715 -7045 -73699
rect -6821 -73323 -6787 -73307
rect -6821 -73715 -6787 -73699
rect -6563 -73323 -6529 -73307
rect -6563 -73715 -6529 -73699
rect -6305 -73323 -6271 -73307
rect -6305 -73715 -6271 -73699
rect -6047 -73323 -6013 -73307
rect -6047 -73715 -6013 -73699
rect -5789 -73323 -5755 -73307
rect -5789 -73715 -5755 -73699
rect -7257 -73792 -7241 -73758
rect -7141 -73792 -7125 -73758
rect -6999 -73792 -6983 -73758
rect -6883 -73792 -6867 -73758
rect -6741 -73792 -6725 -73758
rect -6625 -73792 -6609 -73758
rect -6483 -73792 -6467 -73758
rect -6367 -73792 -6351 -73758
rect -6225 -73792 -6209 -73758
rect -6109 -73792 -6093 -73758
rect -5967 -73792 -5951 -73758
rect -5851 -73792 -5835 -73758
rect -7257 -74124 -7241 -74090
rect -7141 -74124 -7125 -74090
rect -6999 -74124 -6983 -74090
rect -6883 -74124 -6867 -74090
rect -6741 -74124 -6725 -74090
rect -6625 -74124 -6609 -74090
rect -6483 -74124 -6467 -74090
rect -6367 -74124 -6351 -74090
rect -6225 -74124 -6209 -74090
rect -6109 -74124 -6093 -74090
rect -5967 -74124 -5951 -74090
rect -5851 -74124 -5835 -74090
rect -7337 -74183 -7303 -74167
rect -7337 -74575 -7303 -74559
rect -7079 -74183 -7045 -74167
rect -7079 -74575 -7045 -74559
rect -6821 -74183 -6787 -74167
rect -6821 -74575 -6787 -74559
rect -6563 -74183 -6529 -74167
rect -6563 -74575 -6529 -74559
rect -6305 -74183 -6271 -74167
rect -6305 -74575 -6271 -74559
rect -6047 -74183 -6013 -74167
rect -6047 -74575 -6013 -74559
rect -5789 -74183 -5755 -74167
rect -5789 -74575 -5755 -74559
rect -7257 -74652 -7241 -74618
rect -7141 -74652 -7125 -74618
rect -6999 -74652 -6983 -74618
rect -6883 -74652 -6867 -74618
rect -6741 -74652 -6725 -74618
rect -6625 -74652 -6609 -74618
rect -6483 -74652 -6467 -74618
rect -6367 -74652 -6351 -74618
rect -6225 -74652 -6209 -74618
rect -6109 -74652 -6093 -74618
rect -5967 -74652 -5951 -74618
rect -5851 -74652 -5835 -74618
rect -7684 -75770 -7584 -75608
rect -4072 -72931 -4043 -72897
rect -4009 -72931 -3951 -72897
rect -3917 -72931 -3859 -72897
rect -3825 -72931 -3796 -72897
rect -5460 -75770 -5360 -75608
rect -1460 -72828 -1360 -72666
rect 92 -72667 138 -72576
rect 3992 -72586 4008 -72585
rect 4042 -72586 4058 -72585
rect 3992 -72633 3996 -72586
rect 4044 -72633 4058 -72586
rect -4 -72685 38 -72669
rect -4 -72719 4 -72685
rect -4 -72753 38 -72719
rect -4 -72787 4 -72753
rect -4 -72821 38 -72787
rect -4 -72855 4 -72821
rect -4 -72897 38 -72855
rect 72 -72685 138 -72667
rect 72 -72719 88 -72685
rect 122 -72719 138 -72685
rect 72 -72753 138 -72719
rect 72 -72787 88 -72753
rect 122 -72787 138 -72753
rect 72 -72821 138 -72787
rect 72 -72855 88 -72821
rect 122 -72855 138 -72821
rect 72 -72863 138 -72855
rect 316 -72828 416 -72666
rect -3257 -73264 -3241 -73230
rect -3141 -73264 -3125 -73230
rect -2999 -73264 -2983 -73230
rect -2883 -73264 -2867 -73230
rect -2741 -73264 -2725 -73230
rect -2625 -73264 -2609 -73230
rect -2483 -73264 -2467 -73230
rect -2367 -73264 -2351 -73230
rect -2225 -73264 -2209 -73230
rect -2109 -73264 -2093 -73230
rect -1967 -73264 -1951 -73230
rect -1851 -73264 -1835 -73230
rect -3337 -73323 -3303 -73307
rect -3337 -73715 -3303 -73699
rect -3079 -73323 -3045 -73307
rect -3079 -73715 -3045 -73699
rect -2821 -73323 -2787 -73307
rect -2821 -73715 -2787 -73699
rect -2563 -73323 -2529 -73307
rect -2563 -73715 -2529 -73699
rect -2305 -73323 -2271 -73307
rect -2305 -73715 -2271 -73699
rect -2047 -73323 -2013 -73307
rect -2047 -73715 -2013 -73699
rect -1789 -73323 -1755 -73307
rect -1789 -73715 -1755 -73699
rect -3257 -73792 -3241 -73758
rect -3141 -73792 -3125 -73758
rect -2999 -73792 -2983 -73758
rect -2883 -73792 -2867 -73758
rect -2741 -73792 -2725 -73758
rect -2625 -73792 -2609 -73758
rect -2483 -73792 -2467 -73758
rect -2367 -73792 -2351 -73758
rect -2225 -73792 -2209 -73758
rect -2109 -73792 -2093 -73758
rect -1967 -73792 -1951 -73758
rect -1851 -73792 -1835 -73758
rect -3257 -74124 -3241 -74090
rect -3141 -74124 -3125 -74090
rect -2999 -74124 -2983 -74090
rect -2883 -74124 -2867 -74090
rect -2741 -74124 -2725 -74090
rect -2625 -74124 -2609 -74090
rect -2483 -74124 -2467 -74090
rect -2367 -74124 -2351 -74090
rect -2225 -74124 -2209 -74090
rect -2109 -74124 -2093 -74090
rect -1967 -74124 -1951 -74090
rect -1851 -74124 -1835 -74090
rect -3337 -74183 -3303 -74167
rect -3337 -74575 -3303 -74559
rect -3079 -74183 -3045 -74167
rect -3079 -74575 -3045 -74559
rect -2821 -74183 -2787 -74167
rect -2821 -74575 -2787 -74559
rect -2563 -74183 -2529 -74167
rect -2563 -74575 -2529 -74559
rect -2305 -74183 -2271 -74167
rect -2305 -74575 -2271 -74559
rect -2047 -74183 -2013 -74167
rect -2047 -74575 -2013 -74559
rect -1789 -74183 -1755 -74167
rect -1789 -74575 -1755 -74559
rect -3257 -74652 -3241 -74618
rect -3141 -74652 -3125 -74618
rect -2999 -74652 -2983 -74618
rect -2883 -74652 -2867 -74618
rect -2741 -74652 -2725 -74618
rect -2625 -74652 -2609 -74618
rect -2483 -74652 -2467 -74618
rect -2367 -74652 -2351 -74618
rect -2225 -74652 -2209 -74618
rect -2109 -74652 -2093 -74618
rect -1967 -74652 -1951 -74618
rect -1851 -74652 -1835 -74618
rect -3684 -75770 -3584 -75608
rect -72 -72931 -43 -72897
rect -9 -72931 49 -72897
rect 83 -72931 141 -72897
rect 175 -72931 204 -72897
rect -1460 -75770 -1360 -75608
rect 2540 -72828 2640 -72666
rect 4092 -72667 4138 -72576
rect 3996 -72685 4038 -72669
rect 3996 -72719 4004 -72685
rect 3996 -72753 4038 -72719
rect 3996 -72787 4004 -72753
rect 3996 -72821 4038 -72787
rect 3996 -72855 4004 -72821
rect 3996 -72897 4038 -72855
rect 4072 -72685 4138 -72667
rect 4072 -72719 4088 -72685
rect 4122 -72719 4138 -72685
rect 4072 -72753 4138 -72719
rect 4072 -72787 4088 -72753
rect 4122 -72787 4138 -72753
rect 4072 -72821 4138 -72787
rect 4072 -72855 4088 -72821
rect 4122 -72855 4138 -72821
rect 4072 -72863 4138 -72855
rect 4316 -72828 4416 -72666
rect 743 -73264 759 -73230
rect 859 -73264 875 -73230
rect 1001 -73264 1017 -73230
rect 1117 -73264 1133 -73230
rect 1259 -73264 1275 -73230
rect 1375 -73264 1391 -73230
rect 1517 -73264 1533 -73230
rect 1633 -73264 1649 -73230
rect 1775 -73264 1791 -73230
rect 1891 -73264 1907 -73230
rect 2033 -73264 2049 -73230
rect 2149 -73264 2165 -73230
rect 663 -73323 697 -73307
rect 663 -73715 697 -73699
rect 921 -73323 955 -73307
rect 921 -73715 955 -73699
rect 1179 -73323 1213 -73307
rect 1179 -73715 1213 -73699
rect 1437 -73323 1471 -73307
rect 1437 -73715 1471 -73699
rect 1695 -73323 1729 -73307
rect 1695 -73715 1729 -73699
rect 1953 -73323 1987 -73307
rect 1953 -73715 1987 -73699
rect 2211 -73323 2245 -73307
rect 2211 -73715 2245 -73699
rect 743 -73792 759 -73758
rect 859 -73792 875 -73758
rect 1001 -73792 1017 -73758
rect 1117 -73792 1133 -73758
rect 1259 -73792 1275 -73758
rect 1375 -73792 1391 -73758
rect 1517 -73792 1533 -73758
rect 1633 -73792 1649 -73758
rect 1775 -73792 1791 -73758
rect 1891 -73792 1907 -73758
rect 2033 -73792 2049 -73758
rect 2149 -73792 2165 -73758
rect 743 -74124 759 -74090
rect 859 -74124 875 -74090
rect 1001 -74124 1017 -74090
rect 1117 -74124 1133 -74090
rect 1259 -74124 1275 -74090
rect 1375 -74124 1391 -74090
rect 1517 -74124 1533 -74090
rect 1633 -74124 1649 -74090
rect 1775 -74124 1791 -74090
rect 1891 -74124 1907 -74090
rect 2033 -74124 2049 -74090
rect 2149 -74124 2165 -74090
rect 663 -74183 697 -74167
rect 663 -74575 697 -74559
rect 921 -74183 955 -74167
rect 921 -74575 955 -74559
rect 1179 -74183 1213 -74167
rect 1179 -74575 1213 -74559
rect 1437 -74183 1471 -74167
rect 1437 -74575 1471 -74559
rect 1695 -74183 1729 -74167
rect 1695 -74575 1729 -74559
rect 1953 -74183 1987 -74167
rect 1953 -74575 1987 -74559
rect 2211 -74183 2245 -74167
rect 2211 -74575 2245 -74559
rect 743 -74652 759 -74618
rect 859 -74652 875 -74618
rect 1001 -74652 1017 -74618
rect 1117 -74652 1133 -74618
rect 1259 -74652 1275 -74618
rect 1375 -74652 1391 -74618
rect 1517 -74652 1533 -74618
rect 1633 -74652 1649 -74618
rect 1775 -74652 1791 -74618
rect 1891 -74652 1907 -74618
rect 2033 -74652 2049 -74618
rect 2149 -74652 2165 -74618
rect 316 -75770 416 -75608
rect 3928 -72931 3957 -72897
rect 3991 -72931 4049 -72897
rect 4083 -72931 4141 -72897
rect 4175 -72931 4204 -72897
rect 2540 -75770 2640 -75608
rect 6540 -72828 6640 -72666
rect 4743 -73264 4759 -73230
rect 4859 -73264 4875 -73230
rect 5001 -73264 5017 -73230
rect 5117 -73264 5133 -73230
rect 5259 -73264 5275 -73230
rect 5375 -73264 5391 -73230
rect 5517 -73264 5533 -73230
rect 5633 -73264 5649 -73230
rect 5775 -73264 5791 -73230
rect 5891 -73264 5907 -73230
rect 6033 -73264 6049 -73230
rect 6149 -73264 6165 -73230
rect 4663 -73323 4697 -73307
rect 4663 -73715 4697 -73699
rect 4921 -73323 4955 -73307
rect 4921 -73715 4955 -73699
rect 5179 -73323 5213 -73307
rect 5179 -73715 5213 -73699
rect 5437 -73323 5471 -73307
rect 5437 -73715 5471 -73699
rect 5695 -73323 5729 -73307
rect 5695 -73715 5729 -73699
rect 5953 -73323 5987 -73307
rect 5953 -73715 5987 -73699
rect 6211 -73323 6245 -73307
rect 6211 -73715 6245 -73699
rect 4743 -73792 4759 -73758
rect 4859 -73792 4875 -73758
rect 5001 -73792 5017 -73758
rect 5117 -73792 5133 -73758
rect 5259 -73792 5275 -73758
rect 5375 -73792 5391 -73758
rect 5517 -73792 5533 -73758
rect 5633 -73792 5649 -73758
rect 5775 -73792 5791 -73758
rect 5891 -73792 5907 -73758
rect 6033 -73792 6049 -73758
rect 6149 -73792 6165 -73758
rect 4743 -74124 4759 -74090
rect 4859 -74124 4875 -74090
rect 5001 -74124 5017 -74090
rect 5117 -74124 5133 -74090
rect 5259 -74124 5275 -74090
rect 5375 -74124 5391 -74090
rect 5517 -74124 5533 -74090
rect 5633 -74124 5649 -74090
rect 5775 -74124 5791 -74090
rect 5891 -74124 5907 -74090
rect 6033 -74124 6049 -74090
rect 6149 -74124 6165 -74090
rect 4663 -74183 4697 -74167
rect 4663 -74575 4697 -74559
rect 4921 -74183 4955 -74167
rect 4921 -74575 4955 -74559
rect 5179 -74183 5213 -74167
rect 5179 -74575 5213 -74559
rect 5437 -74183 5471 -74167
rect 5437 -74575 5471 -74559
rect 5695 -74183 5729 -74167
rect 5695 -74575 5729 -74559
rect 5953 -74183 5987 -74167
rect 5953 -74575 5987 -74559
rect 6211 -74183 6245 -74167
rect 6211 -74575 6245 -74559
rect 4743 -74652 4759 -74618
rect 4859 -74652 4875 -74618
rect 5001 -74652 5017 -74618
rect 5117 -74652 5133 -74618
rect 5259 -74652 5275 -74618
rect 5375 -74652 5391 -74618
rect 5517 -74652 5533 -74618
rect 5633 -74652 5649 -74618
rect 5775 -74652 5791 -74618
rect 5891 -74652 5907 -74618
rect 6033 -74652 6049 -74618
rect 6149 -74652 6165 -74618
rect 4316 -75770 4416 -75608
rect 6540 -75770 6640 -75608
<< viali >>
rect 25922 -27756 25984 -27656
rect 25984 -27756 50104 -27656
rect 50104 -27756 50166 -27656
rect 25822 -41706 25922 -28276
rect 32226 -30457 32690 -30423
rect 33244 -30457 33708 -30423
rect 34262 -30457 34726 -30423
rect 35280 -30457 35744 -30423
rect 36298 -30457 36762 -30423
rect 37316 -30457 37780 -30423
rect 38334 -30457 38798 -30423
rect 39352 -30457 39816 -30423
rect 40370 -30457 40834 -30423
rect 41388 -30457 41852 -30423
rect 42406 -30457 42870 -30423
rect 43424 -30457 43888 -30423
rect 44442 -30457 44906 -30423
rect 45460 -30457 45924 -30423
rect 46478 -30457 46942 -30423
rect 47496 -30457 47960 -30423
rect 31932 -31092 31966 -30516
rect 32950 -31092 32984 -30516
rect 33968 -31092 34002 -30516
rect 34986 -31092 35020 -30516
rect 36004 -31092 36038 -30516
rect 37022 -31092 37056 -30516
rect 38040 -31092 38074 -30516
rect 39058 -31092 39092 -30516
rect 40076 -31092 40110 -30516
rect 41094 -31092 41128 -30516
rect 42112 -31092 42146 -30516
rect 43130 -31092 43164 -30516
rect 44148 -31092 44182 -30516
rect 45166 -31092 45200 -30516
rect 46184 -31092 46218 -30516
rect 47202 -31092 47236 -30516
rect 48220 -31092 48254 -30516
rect 32226 -31185 32690 -31151
rect 33244 -31185 33708 -31151
rect 34262 -31185 34726 -31151
rect 35280 -31185 35744 -31151
rect 36298 -31185 36762 -31151
rect 37316 -31185 37780 -31151
rect 38334 -31185 38798 -31151
rect 39352 -31185 39816 -31151
rect 40370 -31185 40834 -31151
rect 41388 -31185 41852 -31151
rect 42406 -31185 42870 -31151
rect 43424 -31185 43888 -31151
rect 44442 -31185 44906 -31151
rect 45460 -31185 45924 -31151
rect 46478 -31185 46942 -31151
rect 47496 -31185 47960 -31151
rect 32226 -31593 32690 -31559
rect 33244 -31593 33708 -31559
rect 34262 -31593 34726 -31559
rect 35280 -31593 35744 -31559
rect 36298 -31593 36762 -31559
rect 37316 -31593 37780 -31559
rect 38334 -31593 38798 -31559
rect 39352 -31593 39816 -31559
rect 40370 -31593 40834 -31559
rect 41388 -31593 41852 -31559
rect 42406 -31593 42870 -31559
rect 43424 -31593 43888 -31559
rect 44442 -31593 44906 -31559
rect 45460 -31593 45924 -31559
rect 46478 -31593 46942 -31559
rect 47496 -31593 47960 -31559
rect 31932 -32228 31966 -31652
rect 32950 -32228 32984 -31652
rect 33968 -32228 34002 -31652
rect 34986 -32228 35020 -31652
rect 36004 -32228 36038 -31652
rect 37022 -32228 37056 -31652
rect 38040 -32228 38074 -31652
rect 39058 -32228 39092 -31652
rect 40076 -32228 40110 -31652
rect 41094 -32228 41128 -31652
rect 42112 -32228 42146 -31652
rect 43130 -32228 43164 -31652
rect 44148 -32228 44182 -31652
rect 45166 -32228 45200 -31652
rect 46184 -32228 46218 -31652
rect 47202 -32228 47236 -31652
rect 48220 -32228 48254 -31652
rect 32226 -32321 32690 -32287
rect 33244 -32321 33708 -32287
rect 34262 -32321 34726 -32287
rect 35280 -32321 35744 -32287
rect 36298 -32321 36762 -32287
rect 37316 -32321 37780 -32287
rect 38334 -32321 38798 -32287
rect 39352 -32321 39816 -32287
rect 40370 -32321 40834 -32287
rect 41388 -32321 41852 -32287
rect 42406 -32321 42870 -32287
rect 43424 -32321 43888 -32287
rect 44442 -32321 44906 -32287
rect 45460 -32321 45924 -32287
rect 46478 -32321 46942 -32287
rect 47496 -32321 47960 -32287
rect 32226 -32729 32690 -32695
rect 33244 -32729 33708 -32695
rect 34262 -32729 34726 -32695
rect 35280 -32729 35744 -32695
rect 36298 -32729 36762 -32695
rect 37316 -32729 37780 -32695
rect 38334 -32729 38798 -32695
rect 39352 -32729 39816 -32695
rect 40370 -32729 40834 -32695
rect 41388 -32729 41852 -32695
rect 42406 -32729 42870 -32695
rect 43424 -32729 43888 -32695
rect 44442 -32729 44906 -32695
rect 45460 -32729 45924 -32695
rect 46478 -32729 46942 -32695
rect 47496 -32729 47960 -32695
rect 31932 -33364 31966 -32788
rect 32950 -33364 32984 -32788
rect 33968 -33364 34002 -32788
rect 34986 -33364 35020 -32788
rect 36004 -33364 36038 -32788
rect 37022 -33364 37056 -32788
rect 38040 -33364 38074 -32788
rect 39058 -33364 39092 -32788
rect 40076 -33364 40110 -32788
rect 41094 -33364 41128 -32788
rect 42112 -33364 42146 -32788
rect 43130 -33364 43164 -32788
rect 44148 -33364 44182 -32788
rect 45166 -33364 45200 -32788
rect 46184 -33364 46218 -32788
rect 47202 -33364 47236 -32788
rect 48220 -33364 48254 -32788
rect 32226 -33457 32690 -33423
rect 33244 -33457 33708 -33423
rect 34262 -33457 34726 -33423
rect 35280 -33457 35744 -33423
rect 36298 -33457 36762 -33423
rect 37316 -33457 37780 -33423
rect 38334 -33457 38798 -33423
rect 39352 -33457 39816 -33423
rect 40370 -33457 40834 -33423
rect 41388 -33457 41852 -33423
rect 42406 -33457 42870 -33423
rect 43424 -33457 43888 -33423
rect 44442 -33457 44906 -33423
rect 45460 -33457 45924 -33423
rect 46478 -33457 46942 -33423
rect 47496 -33457 47960 -33423
rect 33420 -34367 33884 -34333
rect 34438 -34367 34902 -34333
rect 35456 -34367 35920 -34333
rect 36474 -34367 36938 -34333
rect 37492 -34367 37956 -34333
rect 38510 -34367 38974 -34333
rect 39528 -34367 39992 -34333
rect 40546 -34367 41010 -34333
rect 41564 -34367 42028 -34333
rect 42582 -34367 43046 -34333
rect 43600 -34367 44064 -34333
rect 44618 -34367 45082 -34333
rect 45636 -34367 46100 -34333
rect 46654 -34367 47118 -34333
rect 33126 -35002 33160 -34426
rect 34144 -35002 34178 -34426
rect 35162 -35002 35196 -34426
rect 36180 -35002 36214 -34426
rect 37198 -35002 37232 -34426
rect 38216 -35002 38250 -34426
rect 39234 -35002 39268 -34426
rect 40252 -35002 40286 -34426
rect 41270 -35002 41304 -34426
rect 42288 -35002 42322 -34426
rect 43306 -35002 43340 -34426
rect 44324 -35002 44358 -34426
rect 45342 -35002 45376 -34426
rect 46360 -35002 46394 -34426
rect 47378 -35002 47412 -34426
rect 33420 -35095 33884 -35061
rect 34438 -35095 34902 -35061
rect 35456 -35095 35920 -35061
rect 36474 -35095 36938 -35061
rect 37492 -35095 37956 -35061
rect 38510 -35095 38974 -35061
rect 39528 -35095 39992 -35061
rect 40546 -35095 41010 -35061
rect 41564 -35095 42028 -35061
rect 42582 -35095 43046 -35061
rect 43600 -35095 44064 -35061
rect 44618 -35095 45082 -35061
rect 45636 -35095 46100 -35061
rect 46654 -35095 47118 -35061
rect 33420 -35399 33884 -35365
rect 34438 -35399 34902 -35365
rect 35456 -35399 35920 -35365
rect 36474 -35399 36938 -35365
rect 37492 -35399 37956 -35365
rect 38510 -35399 38974 -35365
rect 39528 -35399 39992 -35365
rect 40546 -35399 41010 -35365
rect 41564 -35399 42028 -35365
rect 42582 -35399 43046 -35365
rect 43600 -35399 44064 -35365
rect 44618 -35399 45082 -35365
rect 45636 -35399 46100 -35365
rect 46654 -35399 47118 -35365
rect 33126 -36034 33160 -35458
rect 34144 -36034 34178 -35458
rect 35162 -36034 35196 -35458
rect 36180 -36034 36214 -35458
rect 37198 -36034 37232 -35458
rect 38216 -36034 38250 -35458
rect 39234 -36034 39268 -35458
rect 40252 -36034 40286 -35458
rect 41270 -36034 41304 -35458
rect 42288 -36034 42322 -35458
rect 43306 -36034 43340 -35458
rect 44324 -36034 44358 -35458
rect 45342 -36034 45376 -35458
rect 46360 -36034 46394 -35458
rect 47378 -36034 47412 -35458
rect 33420 -36127 33884 -36093
rect 34438 -36127 34902 -36093
rect 35456 -36127 35920 -36093
rect 36474 -36127 36938 -36093
rect 37492 -36127 37956 -36093
rect 38510 -36127 38974 -36093
rect 39528 -36127 39992 -36093
rect 40546 -36127 41010 -36093
rect 41564 -36127 42028 -36093
rect 42582 -36127 43046 -36093
rect 43600 -36127 44064 -36093
rect 44618 -36127 45082 -36093
rect 45636 -36127 46100 -36093
rect 46654 -36127 47118 -36093
rect 33212 -37003 33676 -36969
rect 34230 -37003 34694 -36969
rect 35248 -37003 35712 -36969
rect 36266 -37003 36730 -36969
rect 37284 -37003 37748 -36969
rect 38302 -37003 38766 -36969
rect 39320 -37003 39784 -36969
rect 40338 -37003 40802 -36969
rect 41356 -37003 41820 -36969
rect 42374 -37003 42838 -36969
rect 43392 -37003 43856 -36969
rect 44410 -37003 44874 -36969
rect 45428 -37003 45892 -36969
rect 46446 -37003 46910 -36969
rect 47464 -37003 47928 -36969
rect 27908 -37107 28372 -37073
rect 28926 -37107 29390 -37073
rect 29944 -37107 30408 -37073
rect 30962 -37107 31426 -37073
rect 27614 -37742 27648 -37166
rect 28632 -37742 28666 -37166
rect 29650 -37742 29684 -37166
rect 30668 -37742 30702 -37166
rect 31686 -37742 31720 -37166
rect 32918 -37638 32952 -37062
rect 33936 -37638 33970 -37062
rect 34954 -37638 34988 -37062
rect 35972 -37638 36006 -37062
rect 36990 -37638 37024 -37062
rect 38008 -37638 38042 -37062
rect 39026 -37638 39060 -37062
rect 40044 -37638 40078 -37062
rect 41062 -37638 41096 -37062
rect 42080 -37638 42114 -37062
rect 43098 -37638 43132 -37062
rect 44116 -37638 44150 -37062
rect 45134 -37638 45168 -37062
rect 46152 -37638 46186 -37062
rect 47170 -37638 47204 -37062
rect 48188 -37638 48222 -37062
rect 33212 -37731 33676 -37697
rect 34230 -37731 34694 -37697
rect 35248 -37731 35712 -37697
rect 36266 -37731 36730 -37697
rect 37284 -37731 37748 -37697
rect 38302 -37731 38766 -37697
rect 39320 -37731 39784 -37697
rect 40338 -37731 40802 -37697
rect 41356 -37731 41820 -37697
rect 42374 -37731 42838 -37697
rect 43392 -37731 43856 -37697
rect 44410 -37731 44874 -37697
rect 45428 -37731 45892 -37697
rect 46446 -37731 46910 -37697
rect 47464 -37731 47928 -37697
rect 27908 -37835 28372 -37801
rect 28926 -37835 29390 -37801
rect 29944 -37835 30408 -37801
rect 30962 -37835 31426 -37801
rect 27908 -38139 28372 -38105
rect 28926 -38139 29390 -38105
rect 29944 -38139 30408 -38105
rect 30962 -38139 31426 -38105
rect 27614 -38774 27648 -38198
rect 28632 -38774 28666 -38198
rect 29650 -38774 29684 -38198
rect 30668 -38774 30702 -38198
rect 31686 -38774 31720 -38198
rect 33212 -38259 33676 -38225
rect 34230 -38259 34694 -38225
rect 35248 -38259 35712 -38225
rect 36266 -38259 36730 -38225
rect 37284 -38259 37748 -38225
rect 38302 -38259 38766 -38225
rect 39320 -38259 39784 -38225
rect 40338 -38259 40802 -38225
rect 41356 -38259 41820 -38225
rect 42374 -38259 42838 -38225
rect 43392 -38259 43856 -38225
rect 44410 -38259 44874 -38225
rect 45428 -38259 45892 -38225
rect 46446 -38259 46910 -38225
rect 47464 -38259 47928 -38225
rect 27908 -38867 28372 -38833
rect 28926 -38867 29390 -38833
rect 29944 -38867 30408 -38833
rect 30962 -38867 31426 -38833
rect 32918 -38894 32952 -38318
rect 33936 -38894 33970 -38318
rect 34954 -38894 34988 -38318
rect 35972 -38894 36006 -38318
rect 36990 -38894 37024 -38318
rect 38008 -38894 38042 -38318
rect 39026 -38894 39060 -38318
rect 40044 -38894 40078 -38318
rect 41062 -38894 41096 -38318
rect 42080 -38894 42114 -38318
rect 43098 -38894 43132 -38318
rect 44116 -38894 44150 -38318
rect 45134 -38894 45168 -38318
rect 46152 -38894 46186 -38318
rect 47170 -38894 47204 -38318
rect 48188 -38894 48222 -38318
rect 33212 -38987 33676 -38953
rect 34230 -38987 34694 -38953
rect 35248 -38987 35712 -38953
rect 36266 -38987 36730 -38953
rect 37284 -38987 37748 -38953
rect 38302 -38987 38766 -38953
rect 39320 -38987 39784 -38953
rect 40338 -38987 40802 -38953
rect 41356 -38987 41820 -38953
rect 42374 -38987 42838 -38953
rect 43392 -38987 43856 -38953
rect 44410 -38987 44874 -38953
rect 45428 -38987 45892 -38953
rect 46446 -38987 46910 -38953
rect 47464 -38987 47928 -38953
rect 27908 -39171 28372 -39137
rect 28926 -39171 29390 -39137
rect 29944 -39171 30408 -39137
rect 30962 -39171 31426 -39137
rect 27614 -39806 27648 -39230
rect 28632 -39806 28666 -39230
rect 29650 -39806 29684 -39230
rect 30668 -39806 30702 -39230
rect 31686 -39806 31720 -39230
rect 33212 -39515 33676 -39481
rect 34230 -39515 34694 -39481
rect 35248 -39515 35712 -39481
rect 36266 -39515 36730 -39481
rect 37284 -39515 37748 -39481
rect 38302 -39515 38766 -39481
rect 39320 -39515 39784 -39481
rect 40338 -39515 40802 -39481
rect 41356 -39515 41820 -39481
rect 42374 -39515 42838 -39481
rect 43392 -39515 43856 -39481
rect 44410 -39515 44874 -39481
rect 45428 -39515 45892 -39481
rect 46446 -39515 46910 -39481
rect 47464 -39515 47928 -39481
rect 27908 -39899 28372 -39865
rect 28926 -39899 29390 -39865
rect 29944 -39899 30408 -39865
rect 30962 -39899 31426 -39865
rect 32918 -40150 32952 -39574
rect 33936 -40150 33970 -39574
rect 34954 -40150 34988 -39574
rect 35972 -40150 36006 -39574
rect 36990 -40150 37024 -39574
rect 38008 -40150 38042 -39574
rect 39026 -40150 39060 -39574
rect 40044 -40150 40078 -39574
rect 41062 -40150 41096 -39574
rect 42080 -40150 42114 -39574
rect 43098 -40150 43132 -39574
rect 44116 -40150 44150 -39574
rect 45134 -40150 45168 -39574
rect 46152 -40150 46186 -39574
rect 47170 -40150 47204 -39574
rect 48188 -40150 48222 -39574
rect 27908 -40203 28372 -40169
rect 28926 -40203 29390 -40169
rect 29944 -40203 30408 -40169
rect 30962 -40203 31426 -40169
rect 33212 -40243 33676 -40209
rect 34230 -40243 34694 -40209
rect 35248 -40243 35712 -40209
rect 36266 -40243 36730 -40209
rect 37284 -40243 37748 -40209
rect 38302 -40243 38766 -40209
rect 39320 -40243 39784 -40209
rect 40338 -40243 40802 -40209
rect 41356 -40243 41820 -40209
rect 42374 -40243 42838 -40209
rect 43392 -40243 43856 -40209
rect 44410 -40243 44874 -40209
rect 45428 -40243 45892 -40209
rect 46446 -40243 46910 -40209
rect 47464 -40243 47928 -40209
rect 27614 -40838 27648 -40262
rect 28632 -40838 28666 -40262
rect 29650 -40838 29684 -40262
rect 30668 -40838 30702 -40262
rect 31686 -40838 31720 -40262
rect 33212 -40771 33676 -40737
rect 34230 -40771 34694 -40737
rect 35248 -40771 35712 -40737
rect 36266 -40771 36730 -40737
rect 37284 -40771 37748 -40737
rect 38302 -40771 38766 -40737
rect 39320 -40771 39784 -40737
rect 40338 -40771 40802 -40737
rect 41356 -40771 41820 -40737
rect 42374 -40771 42838 -40737
rect 43392 -40771 43856 -40737
rect 44410 -40771 44874 -40737
rect 45428 -40771 45892 -40737
rect 46446 -40771 46910 -40737
rect 47464 -40771 47928 -40737
rect 27908 -40931 28372 -40897
rect 28926 -40931 29390 -40897
rect 29944 -40931 30408 -40897
rect 30962 -40931 31426 -40897
rect 32918 -41406 32952 -40830
rect 33936 -41406 33970 -40830
rect 34954 -41406 34988 -40830
rect 35972 -41406 36006 -40830
rect 36990 -41406 37024 -40830
rect 38008 -41406 38042 -40830
rect 39026 -41406 39060 -40830
rect 40044 -41406 40078 -40830
rect 41062 -41406 41096 -40830
rect 42080 -41406 42114 -40830
rect 43098 -41406 43132 -40830
rect 44116 -41406 44150 -40830
rect 45134 -41406 45168 -40830
rect 46152 -41406 46186 -40830
rect 47170 -41406 47204 -40830
rect 48188 -41406 48222 -40830
rect 33212 -41499 33676 -41465
rect 34230 -41499 34694 -41465
rect 35248 -41499 35712 -41465
rect 36266 -41499 36730 -41465
rect 37284 -41499 37748 -41465
rect 38302 -41499 38766 -41465
rect 39320 -41499 39784 -41465
rect 40338 -41499 40802 -41465
rect 41356 -41499 41820 -41465
rect 42374 -41499 42838 -41465
rect 43392 -41499 43856 -41465
rect 44410 -41499 44874 -41465
rect 45428 -41499 45892 -41465
rect 46446 -41499 46910 -41465
rect 47464 -41499 47928 -41465
rect 50166 -41706 50266 -28276
rect 25922 -42326 25984 -42226
rect 25984 -42326 50104 -42226
rect 50104 -42326 50166 -42226
rect 52256 -39080 52318 -38980
rect 52318 -39080 55358 -38980
rect 55358 -39080 55420 -38980
rect 52156 -42087 52256 -39217
rect 52596 -39633 52780 -39599
rect 53054 -39633 53238 -39599
rect 53512 -39633 53696 -39599
rect 53970 -39633 54154 -39599
rect 54428 -39633 54612 -39599
rect 54886 -39633 55070 -39599
rect 52442 -39868 52476 -39692
rect 52900 -39868 52934 -39692
rect 53358 -39868 53392 -39692
rect 53816 -39868 53850 -39692
rect 54274 -39868 54308 -39692
rect 54732 -39868 54766 -39692
rect 55190 -39868 55224 -39692
rect 52596 -39961 52780 -39927
rect 53054 -39961 53238 -39927
rect 53512 -39961 53696 -39927
rect 53970 -39961 54154 -39927
rect 54428 -39961 54612 -39927
rect 54886 -39961 55070 -39927
rect 52605 -40516 52689 -40482
rect 52863 -40516 52947 -40482
rect 53121 -40516 53205 -40482
rect 53379 -40516 53463 -40482
rect 53637 -40516 53721 -40482
rect 53895 -40516 53979 -40482
rect 54153 -40516 54237 -40482
rect 54411 -40516 54495 -40482
rect 54669 -40516 54753 -40482
rect 54927 -40516 55011 -40482
rect 52501 -40951 52535 -40575
rect 52759 -40951 52793 -40575
rect 53017 -40951 53051 -40575
rect 53275 -40951 53309 -40575
rect 53533 -40951 53567 -40575
rect 53791 -40951 53825 -40575
rect 54049 -40951 54083 -40575
rect 54307 -40951 54341 -40575
rect 54565 -40951 54599 -40575
rect 54823 -40951 54857 -40575
rect 55081 -40951 55115 -40575
rect 52605 -41044 52689 -41010
rect 52863 -41044 52947 -41010
rect 53121 -41044 53205 -41010
rect 53379 -41044 53463 -41010
rect 53637 -41044 53721 -41010
rect 53895 -41044 53979 -41010
rect 54153 -41044 54237 -41010
rect 54411 -41044 54495 -41010
rect 54669 -41044 54753 -41010
rect 54927 -41044 55011 -41010
rect 52605 -41376 52689 -41342
rect 52863 -41376 52947 -41342
rect 53121 -41376 53205 -41342
rect 53379 -41376 53463 -41342
rect 53637 -41376 53721 -41342
rect 53895 -41376 53979 -41342
rect 54153 -41376 54237 -41342
rect 54411 -41376 54495 -41342
rect 54669 -41376 54753 -41342
rect 54927 -41376 55011 -41342
rect 52501 -41811 52535 -41435
rect 52759 -41811 52793 -41435
rect 53017 -41811 53051 -41435
rect 53275 -41811 53309 -41435
rect 53533 -41811 53567 -41435
rect 53791 -41811 53825 -41435
rect 54049 -41811 54083 -41435
rect 54307 -41811 54341 -41435
rect 54565 -41811 54599 -41435
rect 54823 -41811 54857 -41435
rect 55081 -41811 55115 -41435
rect 52605 -41904 52689 -41870
rect 52863 -41904 52947 -41870
rect 53121 -41904 53205 -41870
rect 53379 -41904 53463 -41870
rect 53637 -41904 53721 -41870
rect 53895 -41904 53979 -41870
rect 54153 -41904 54237 -41870
rect 54411 -41904 54495 -41870
rect 54669 -41904 54753 -41870
rect 54927 -41904 55011 -41870
rect 55420 -42087 55520 -39217
rect 55958 -39080 56020 -38980
rect 56020 -39080 58100 -38980
rect 58100 -39080 58162 -38980
rect 55858 -41338 55958 -39172
rect 58166 -39406 58262 -39172
rect 56174 -39833 56258 -39799
rect 56432 -39833 56516 -39799
rect 56690 -39833 56774 -39799
rect 56948 -39833 57032 -39799
rect 57206 -39833 57290 -39799
rect 57464 -39833 57548 -39799
rect 57722 -39833 57806 -39799
rect 56070 -40268 56104 -39892
rect 56328 -40268 56362 -39892
rect 56586 -40268 56620 -39892
rect 56844 -40268 56878 -39892
rect 57102 -40268 57136 -39892
rect 57360 -40268 57394 -39892
rect 57618 -40268 57652 -39892
rect 57876 -40268 57910 -39892
rect 56174 -40361 56258 -40327
rect 56432 -40361 56516 -40327
rect 56690 -40361 56774 -40327
rect 56948 -40361 57032 -40327
rect 57206 -40361 57290 -40327
rect 57464 -40361 57548 -40327
rect 57722 -40361 57806 -40327
rect 56174 -40693 56258 -40659
rect 56432 -40693 56516 -40659
rect 56690 -40693 56774 -40659
rect 56948 -40693 57032 -40659
rect 57206 -40693 57290 -40659
rect 57464 -40693 57548 -40659
rect 57722 -40693 57806 -40659
rect 56070 -41128 56104 -40752
rect 56328 -41128 56362 -40752
rect 56586 -41128 56620 -40752
rect 56844 -41128 56878 -40752
rect 57102 -41128 57136 -40752
rect 57360 -41128 57394 -40752
rect 57618 -41128 57652 -40752
rect 57876 -41128 57910 -40752
rect 56174 -41221 56258 -41187
rect 56432 -41221 56516 -41187
rect 56690 -41221 56774 -41187
rect 56948 -41221 57032 -41187
rect 57206 -41221 57290 -41187
rect 57464 -41221 57548 -41187
rect 57722 -41221 57806 -41187
rect 58162 -41338 58262 -39406
rect 55958 -41530 56020 -41430
rect 56020 -41530 58100 -41430
rect 58100 -41530 58162 -41430
rect 56133 -41609 56167 -41575
rect 56225 -41609 56259 -41575
rect 56317 -41609 56351 -41575
rect 56409 -41609 56443 -41575
rect 56501 -41609 56535 -41575
rect 56593 -41609 56627 -41575
rect 56685 -41609 56719 -41575
rect 56777 -41609 56811 -41575
rect 56869 -41609 56903 -41575
rect 56958 -41608 56992 -41574
rect 57050 -41608 57084 -41574
rect 57147 -41609 57181 -41575
rect 57239 -41609 57273 -41575
rect 57331 -41609 57365 -41575
rect 57423 -41609 57457 -41575
rect 57515 -41609 57549 -41575
rect 57607 -41609 57641 -41575
rect 57699 -41609 57733 -41575
rect 57791 -41609 57825 -41575
rect 57883 -41609 57917 -41575
rect 56170 -41887 56218 -41872
rect 56170 -41920 56184 -41887
rect 56184 -41920 56218 -41887
rect 56282 -41920 56330 -41872
rect 56442 -41887 56490 -41872
rect 56442 -41920 56460 -41887
rect 56460 -41920 56490 -41887
rect 56550 -41920 56598 -41872
rect 56682 -41887 56730 -41872
rect 56682 -41920 56692 -41887
rect 56692 -41920 56726 -41887
rect 56726 -41920 56730 -41887
rect 56856 -41887 56904 -41872
rect 56856 -41920 56860 -41887
rect 56860 -41920 56894 -41887
rect 56894 -41920 56904 -41887
rect 57152 -41887 57186 -41886
rect 57152 -41920 57156 -41887
rect 57156 -41920 57186 -41887
rect 57330 -41887 57378 -41874
rect 57330 -41921 57358 -41887
rect 57358 -41921 57378 -41887
rect 57330 -41922 57378 -41921
rect 57444 -41922 57492 -41874
rect 57560 -41887 57608 -41872
rect 57560 -41920 57590 -41887
rect 57590 -41920 57608 -41887
rect 57720 -41920 57768 -41872
rect 56862 -42009 56863 -41990
rect 56863 -42009 56897 -41990
rect 56897 -42009 56910 -41990
rect 56862 -42038 56910 -42009
rect 57142 -42009 57153 -41990
rect 57153 -42009 57187 -41990
rect 57187 -42009 57190 -41990
rect 57142 -42038 57190 -42009
rect 56133 -42153 56167 -42119
rect 56225 -42153 56259 -42119
rect 56317 -42153 56351 -42119
rect 56409 -42153 56443 -42119
rect 56501 -42153 56535 -42119
rect 56593 -42153 56627 -42119
rect 56685 -42153 56719 -42119
rect 56777 -42153 56811 -42119
rect 56869 -42153 56903 -42119
rect 56958 -42154 56992 -42120
rect 57050 -42152 57084 -42118
rect 57832 -41887 57880 -41872
rect 57832 -41920 57866 -41887
rect 57866 -41920 57880 -41887
rect 57147 -42153 57181 -42119
rect 57239 -42153 57273 -42119
rect 57331 -42153 57365 -42119
rect 57423 -42153 57457 -42119
rect 57515 -42153 57549 -42119
rect 57607 -42153 57641 -42119
rect 57699 -42153 57733 -42119
rect 57791 -42153 57825 -42119
rect 57883 -42153 57917 -42119
rect 52256 -42324 52318 -42224
rect 52318 -42324 55358 -42224
rect 55358 -42324 55420 -42224
rect 54200 -42418 55422 -42384
rect 55422 -42418 55424 -42384
rect 54104 -42578 54138 -42454
rect 54206 -42542 54266 -42482
rect 55289 -42547 55359 -42477
rect 54104 -42810 54138 -42578
rect 55484 -42578 55518 -42476
rect 56470 -42446 56532 -42346
rect 56532 -42446 57516 -42346
rect 57516 -42446 57628 -42346
rect 56370 -42508 56470 -42487
rect 54104 -42922 54138 -42810
rect 54218 -42782 54252 -42606
rect 54346 -42782 54380 -42606
rect 54474 -42782 54508 -42606
rect 54602 -42782 54636 -42606
rect 54730 -42782 54764 -42606
rect 54858 -42782 54892 -42606
rect 54986 -42782 55020 -42606
rect 55114 -42782 55148 -42606
rect 55242 -42782 55276 -42606
rect 55370 -42782 55404 -42606
rect 54201 -42906 54274 -42833
rect 55348 -42907 55423 -42832
rect 55484 -42810 55518 -42578
rect 55484 -42922 55518 -42810
rect 54198 -43000 54200 -42966
rect 54200 -43000 55422 -42966
rect 55902 -42918 55936 -42624
rect 56075 -42664 56109 -42630
rect 56016 -42890 56050 -42714
rect 56134 -42890 56168 -42714
rect 56248 -42918 56282 -42624
rect 56370 -43070 56470 -42508
rect 56726 -42512 56786 -42502
rect 56726 -42552 56736 -42512
rect 56736 -42552 56776 -42512
rect 56776 -42552 56786 -42512
rect 56726 -42562 56786 -42552
rect 57316 -42512 57376 -42502
rect 57316 -42552 57326 -42512
rect 57326 -42552 57366 -42512
rect 57366 -42552 57376 -42512
rect 57316 -42562 57376 -42552
rect 57628 -42510 57728 -42486
rect 56562 -42804 56596 -42628
rect 56680 -42804 56714 -42628
rect 56798 -42804 56832 -42628
rect 56916 -42804 56950 -42628
rect 57034 -42804 57068 -42628
rect 57152 -42804 57186 -42628
rect 57270 -42804 57304 -42628
rect 57388 -42804 57422 -42628
rect 57506 -42804 57540 -42628
rect 56548 -42876 56608 -42866
rect 56548 -42916 56558 -42876
rect 56558 -42916 56598 -42876
rect 56598 -42916 56608 -42876
rect 56548 -42926 56608 -42916
rect 56924 -42922 56972 -42874
rect 57144 -42922 57192 -42874
rect 57496 -42876 57556 -42866
rect 57496 -42916 57506 -42876
rect 57506 -42916 57546 -42876
rect 57546 -42916 57556 -42876
rect 57496 -42926 57556 -42916
rect 13222 -43256 13284 -43156
rect 13284 -43256 50204 -43156
rect 50204 -43256 50266 -43156
rect 28320 -43976 28784 -43942
rect 29338 -43976 29802 -43942
rect 30356 -43976 30820 -43942
rect 31374 -43976 31838 -43942
rect 32392 -43976 32856 -43942
rect 33410 -43976 33874 -43942
rect 34428 -43976 34892 -43942
rect 35446 -43976 35910 -43942
rect 36464 -43976 36928 -43942
rect 37482 -43976 37946 -43942
rect 38500 -43976 38964 -43942
rect 39518 -43976 39982 -43942
rect 40536 -43976 41000 -43942
rect 41554 -43976 42018 -43942
rect 42572 -43976 43036 -43942
rect 43590 -43976 44054 -43942
rect 44608 -43976 45072 -43942
rect 45626 -43976 46090 -43942
rect 46644 -43976 47108 -43942
rect 47662 -43976 48126 -43942
rect 10342 -56739 10562 -56738
rect 11834 -56739 12036 -56738
rect 10342 -56772 10392 -56739
rect 10392 -56772 10562 -56739
rect 11834 -56772 12010 -56739
rect 12010 -56772 12036 -56739
rect 12070 -56835 12106 -56834
rect 10294 -57408 10296 -56836
rect 10296 -57408 10330 -56836
rect 10330 -57408 10332 -56836
rect 10514 -56875 10598 -56841
rect 10772 -56875 10856 -56841
rect 11030 -56875 11114 -56841
rect 11288 -56875 11372 -56841
rect 11546 -56875 11630 -56841
rect 11804 -56875 11888 -56841
rect 10410 -57310 10444 -56934
rect 10668 -57310 10702 -56934
rect 10926 -57310 10960 -56934
rect 11184 -57310 11218 -56934
rect 11442 -57310 11476 -56934
rect 11700 -57310 11734 -56934
rect 11958 -57310 11992 -56934
rect 10514 -57403 10598 -57369
rect 10772 -57403 10856 -57369
rect 11030 -57403 11114 -57369
rect 11288 -57403 11372 -57369
rect 11546 -57403 11630 -57369
rect 11804 -57403 11888 -57369
rect 12070 -57409 12072 -56835
rect 12072 -57409 12106 -56835
rect 12209 -57275 12243 -57241
rect 12301 -57275 12335 -57241
rect 12393 -57275 12427 -57241
rect 12070 -57410 12106 -57409
rect 11834 -57471 12036 -57470
rect 10342 -57505 10392 -57472
rect 10392 -57505 10562 -57472
rect 11834 -57504 12010 -57471
rect 12010 -57504 12036 -57471
rect 10342 -57506 10562 -57505
rect 12238 -57586 12286 -57538
rect 12342 -57553 12390 -57538
rect 12342 -57586 12376 -57553
rect 12376 -57586 12390 -57553
rect 10366 -57672 10574 -57670
rect 11838 -57672 12036 -57668
rect 10366 -57706 10392 -57672
rect 10392 -57706 10574 -57672
rect 11838 -57706 12010 -57672
rect 12010 -57706 12036 -57672
rect 10366 -57708 10574 -57706
rect 10294 -58124 10296 -57768
rect 10296 -58124 10330 -57768
rect 10514 -57808 10598 -57774
rect 10772 -57808 10856 -57774
rect 11030 -57808 11114 -57774
rect 11288 -57808 11372 -57774
rect 11546 -57808 11630 -57774
rect 11804 -57808 11888 -57774
rect 10410 -58034 10444 -57858
rect 10668 -58034 10702 -57858
rect 10926 -58034 10960 -57858
rect 11184 -58034 11218 -57858
rect 11442 -58034 11476 -57858
rect 11700 -58034 11734 -57858
rect 11958 -58034 11992 -57858
rect 10514 -58118 10598 -58084
rect 10772 -58118 10856 -58084
rect 11030 -58118 11114 -58084
rect 11288 -58118 11372 -58084
rect 11546 -58118 11630 -58084
rect 11804 -58118 11888 -58084
rect 12070 -58124 12072 -57768
rect 12072 -58124 12106 -57768
rect 12106 -58124 12108 -57768
rect 12209 -57819 12243 -57785
rect 12301 -57819 12335 -57785
rect 12393 -57819 12427 -57785
rect 10364 -58186 10572 -58184
rect 10364 -58220 10392 -58186
rect 10392 -58220 10572 -58186
rect 11836 -58220 12010 -58186
rect 12010 -58220 12038 -58186
rect 11836 -58222 12038 -58220
rect 13122 -58308 13222 -44048
rect 16554 -44452 17018 -44418
rect 17572 -44452 18036 -44418
rect 18590 -44452 19054 -44418
rect 19608 -44452 20072 -44418
rect 20626 -44452 21090 -44418
rect 21644 -44452 22108 -44418
rect 22662 -44452 23126 -44418
rect 23680 -44452 24144 -44418
rect 24698 -44452 25162 -44418
rect 16260 -45078 16294 -44502
rect 17278 -45078 17312 -44502
rect 18296 -45078 18330 -44502
rect 19314 -45078 19348 -44502
rect 20332 -45078 20366 -44502
rect 21350 -45078 21384 -44502
rect 22368 -45078 22402 -44502
rect 23386 -45078 23420 -44502
rect 24404 -45078 24438 -44502
rect 25422 -45078 25456 -44502
rect 28026 -44602 28060 -44026
rect 29044 -44602 29078 -44026
rect 30062 -44602 30096 -44026
rect 31080 -44602 31114 -44026
rect 32098 -44602 32132 -44026
rect 33116 -44602 33150 -44026
rect 34134 -44602 34168 -44026
rect 35152 -44602 35186 -44026
rect 36170 -44602 36204 -44026
rect 37188 -44602 37222 -44026
rect 38206 -44602 38240 -44026
rect 39224 -44602 39258 -44026
rect 40242 -44602 40276 -44026
rect 41260 -44602 41294 -44026
rect 42278 -44602 42312 -44026
rect 43296 -44602 43330 -44026
rect 44314 -44602 44348 -44026
rect 45332 -44602 45366 -44026
rect 46350 -44602 46384 -44026
rect 47368 -44602 47402 -44026
rect 48386 -44602 48420 -44026
rect 56370 -43563 56470 -43070
rect 57628 -43144 57728 -42510
rect 57806 -42918 57840 -42624
rect 57979 -42664 58013 -42630
rect 57920 -42890 57954 -42714
rect 58038 -42890 58072 -42714
rect 58152 -42918 58186 -42624
rect 57628 -43563 57728 -43144
rect 56470 -43704 56526 -43604
rect 56526 -43704 57510 -43604
rect 57510 -43704 57628 -43604
rect 28320 -44686 28784 -44652
rect 29338 -44686 29802 -44652
rect 30356 -44686 30820 -44652
rect 31374 -44686 31838 -44652
rect 32392 -44686 32856 -44652
rect 33410 -44686 33874 -44652
rect 34428 -44686 34892 -44652
rect 35446 -44686 35910 -44652
rect 36464 -44686 36928 -44652
rect 37482 -44686 37946 -44652
rect 38500 -44686 38964 -44652
rect 39518 -44686 39982 -44652
rect 40536 -44686 41000 -44652
rect 41554 -44686 42018 -44652
rect 42572 -44686 43036 -44652
rect 43590 -44686 44054 -44652
rect 44608 -44686 45072 -44652
rect 45626 -44686 46090 -44652
rect 46644 -44686 47108 -44652
rect 47662 -44686 48126 -44652
rect 28320 -44794 28784 -44760
rect 29338 -44794 29802 -44760
rect 30356 -44794 30820 -44760
rect 31374 -44794 31838 -44760
rect 32392 -44794 32856 -44760
rect 33410 -44794 33874 -44760
rect 34428 -44794 34892 -44760
rect 35446 -44794 35910 -44760
rect 36464 -44794 36928 -44760
rect 37482 -44794 37946 -44760
rect 38500 -44794 38964 -44760
rect 39518 -44794 39982 -44760
rect 40536 -44794 41000 -44760
rect 41554 -44794 42018 -44760
rect 42572 -44794 43036 -44760
rect 43590 -44794 44054 -44760
rect 44608 -44794 45072 -44760
rect 45626 -44794 46090 -44760
rect 46644 -44794 47108 -44760
rect 47662 -44794 48126 -44760
rect 16554 -45162 17018 -45128
rect 17572 -45162 18036 -45128
rect 16554 -45270 17018 -45236
rect 18590 -45162 19054 -45128
rect 17572 -45270 18036 -45236
rect 19608 -45162 20072 -45128
rect 18590 -45270 19054 -45236
rect 20626 -45162 21090 -45128
rect 19608 -45270 20072 -45236
rect 21644 -45162 22108 -45128
rect 20626 -45270 21090 -45236
rect 22662 -45162 23126 -45128
rect 21644 -45270 22108 -45236
rect 23680 -45162 24144 -45128
rect 22662 -45270 23126 -45236
rect 24698 -45162 25162 -45128
rect 23680 -45270 24144 -45236
rect 24698 -45270 25162 -45236
rect 16260 -45896 16294 -45320
rect 17278 -45896 17312 -45320
rect 18296 -45896 18330 -45320
rect 19314 -45896 19348 -45320
rect 20332 -45896 20366 -45320
rect 21350 -45896 21384 -45320
rect 22368 -45896 22402 -45320
rect 23386 -45896 23420 -45320
rect 24404 -45896 24438 -45320
rect 25422 -45896 25456 -45320
rect 28026 -45420 28060 -44844
rect 29044 -45420 29078 -44844
rect 30062 -45420 30096 -44844
rect 31080 -45420 31114 -44844
rect 32098 -45420 32132 -44844
rect 33116 -45420 33150 -44844
rect 34134 -45420 34168 -44844
rect 35152 -45420 35186 -44844
rect 36170 -45420 36204 -44844
rect 37188 -45420 37222 -44844
rect 38206 -45420 38240 -44844
rect 39224 -45420 39258 -44844
rect 40242 -45420 40276 -44844
rect 41260 -45420 41294 -44844
rect 42278 -45420 42312 -44844
rect 43296 -45420 43330 -44844
rect 44314 -45420 44348 -44844
rect 45332 -45420 45366 -44844
rect 46350 -45420 46384 -44844
rect 47368 -45420 47402 -44844
rect 48386 -45420 48420 -44844
rect 28320 -45504 28784 -45470
rect 29338 -45504 29802 -45470
rect 30356 -45504 30820 -45470
rect 31374 -45504 31838 -45470
rect 32392 -45504 32856 -45470
rect 33410 -45504 33874 -45470
rect 34428 -45504 34892 -45470
rect 35446 -45504 35910 -45470
rect 36464 -45504 36928 -45470
rect 37482 -45504 37946 -45470
rect 38500 -45504 38964 -45470
rect 39518 -45504 39982 -45470
rect 40536 -45504 41000 -45470
rect 41554 -45504 42018 -45470
rect 42572 -45504 43036 -45470
rect 43590 -45504 44054 -45470
rect 44608 -45504 45072 -45470
rect 45626 -45504 46090 -45470
rect 46644 -45504 47108 -45470
rect 47662 -45504 48126 -45470
rect 16554 -45980 17018 -45946
rect 17572 -45980 18036 -45946
rect 16554 -46088 17018 -46054
rect 18590 -45980 19054 -45946
rect 17572 -46088 18036 -46054
rect 19608 -45980 20072 -45946
rect 18590 -46088 19054 -46054
rect 20626 -45980 21090 -45946
rect 19608 -46088 20072 -46054
rect 21644 -45980 22108 -45946
rect 20626 -46088 21090 -46054
rect 22662 -45980 23126 -45946
rect 21644 -46088 22108 -46054
rect 23680 -45980 24144 -45946
rect 22662 -46088 23126 -46054
rect 24698 -45980 25162 -45946
rect 23680 -46088 24144 -46054
rect 24698 -46088 25162 -46054
rect 16260 -46714 16294 -46138
rect 17278 -46714 17312 -46138
rect 18296 -46714 18330 -46138
rect 19314 -46714 19348 -46138
rect 20332 -46714 20366 -46138
rect 21350 -46714 21384 -46138
rect 22368 -46714 22402 -46138
rect 23386 -46714 23420 -46138
rect 24404 -46714 24438 -46138
rect 25422 -46714 25456 -46138
rect 28320 -46172 28784 -46138
rect 29338 -46172 29802 -46138
rect 30356 -46172 30820 -46138
rect 31374 -46172 31838 -46138
rect 32392 -46172 32856 -46138
rect 33410 -46172 33874 -46138
rect 34428 -46172 34892 -46138
rect 35446 -46172 35910 -46138
rect 36464 -46172 36928 -46138
rect 37482 -46172 37946 -46138
rect 38500 -46172 38964 -46138
rect 39518 -46172 39982 -46138
rect 40536 -46172 41000 -46138
rect 41554 -46172 42018 -46138
rect 42572 -46172 43036 -46138
rect 43590 -46172 44054 -46138
rect 44608 -46172 45072 -46138
rect 45626 -46172 46090 -46138
rect 46644 -46172 47108 -46138
rect 47662 -46172 48126 -46138
rect 16554 -46798 17018 -46764
rect 17572 -46798 18036 -46764
rect 16554 -46906 17018 -46872
rect 18590 -46798 19054 -46764
rect 17572 -46906 18036 -46872
rect 19608 -46798 20072 -46764
rect 18590 -46906 19054 -46872
rect 20626 -46798 21090 -46764
rect 19608 -46906 20072 -46872
rect 21644 -46798 22108 -46764
rect 20626 -46906 21090 -46872
rect 22662 -46798 23126 -46764
rect 21644 -46906 22108 -46872
rect 23680 -46798 24144 -46764
rect 22662 -46906 23126 -46872
rect 24698 -46798 25162 -46764
rect 23680 -46906 24144 -46872
rect 28026 -46798 28060 -46222
rect 29044 -46798 29078 -46222
rect 30062 -46798 30096 -46222
rect 31080 -46798 31114 -46222
rect 32098 -46798 32132 -46222
rect 33116 -46798 33150 -46222
rect 34134 -46798 34168 -46222
rect 35152 -46798 35186 -46222
rect 36170 -46798 36204 -46222
rect 37188 -46798 37222 -46222
rect 38206 -46798 38240 -46222
rect 39224 -46798 39258 -46222
rect 40242 -46798 40276 -46222
rect 41260 -46798 41294 -46222
rect 42278 -46798 42312 -46222
rect 43296 -46798 43330 -46222
rect 44314 -46798 44348 -46222
rect 45332 -46798 45366 -46222
rect 46350 -46798 46384 -46222
rect 47368 -46798 47402 -46222
rect 48386 -46798 48420 -46222
rect 24698 -46906 25162 -46872
rect 28320 -46882 28784 -46848
rect 29338 -46882 29802 -46848
rect 30356 -46882 30820 -46848
rect 31374 -46882 31838 -46848
rect 32392 -46882 32856 -46848
rect 33410 -46882 33874 -46848
rect 34428 -46882 34892 -46848
rect 35446 -46882 35910 -46848
rect 36464 -46882 36928 -46848
rect 37482 -46882 37946 -46848
rect 38500 -46882 38964 -46848
rect 39518 -46882 39982 -46848
rect 40536 -46882 41000 -46848
rect 41554 -46882 42018 -46848
rect 42572 -46882 43036 -46848
rect 43590 -46882 44054 -46848
rect 44608 -46882 45072 -46848
rect 45626 -46882 46090 -46848
rect 46644 -46882 47108 -46848
rect 47662 -46882 48126 -46848
rect 16260 -47532 16294 -46956
rect 17278 -47532 17312 -46956
rect 18296 -47532 18330 -46956
rect 19314 -47532 19348 -46956
rect 20332 -47532 20366 -46956
rect 21350 -47532 21384 -46956
rect 22368 -47532 22402 -46956
rect 23386 -47532 23420 -46956
rect 24404 -47532 24438 -46956
rect 25422 -47532 25456 -46956
rect 28320 -47404 28784 -47370
rect 29338 -47404 29802 -47370
rect 30356 -47404 30820 -47370
rect 31374 -47404 31838 -47370
rect 32392 -47404 32856 -47370
rect 33410 -47404 33874 -47370
rect 34428 -47404 34892 -47370
rect 35446 -47404 35910 -47370
rect 36464 -47404 36928 -47370
rect 37482 -47404 37946 -47370
rect 38500 -47404 38964 -47370
rect 39518 -47404 39982 -47370
rect 40536 -47404 41000 -47370
rect 41554 -47404 42018 -47370
rect 42572 -47404 43036 -47370
rect 43590 -47404 44054 -47370
rect 44608 -47404 45072 -47370
rect 45626 -47404 46090 -47370
rect 46644 -47404 47108 -47370
rect 47662 -47404 48126 -47370
rect 16554 -47616 17018 -47582
rect 17572 -47616 18036 -47582
rect 16554 -47724 17018 -47690
rect 18590 -47616 19054 -47582
rect 17572 -47724 18036 -47690
rect 19608 -47616 20072 -47582
rect 18590 -47724 19054 -47690
rect 20626 -47616 21090 -47582
rect 19608 -47724 20072 -47690
rect 21644 -47616 22108 -47582
rect 20626 -47724 21090 -47690
rect 22662 -47616 23126 -47582
rect 21644 -47724 22108 -47690
rect 23680 -47616 24144 -47582
rect 22662 -47724 23126 -47690
rect 24698 -47616 25162 -47582
rect 23680 -47724 24144 -47690
rect 24698 -47724 25162 -47690
rect 16260 -48350 16294 -47774
rect 17278 -48350 17312 -47774
rect 18296 -48350 18330 -47774
rect 19314 -48350 19348 -47774
rect 20332 -48350 20366 -47774
rect 21350 -48350 21384 -47774
rect 22368 -48350 22402 -47774
rect 23386 -48350 23420 -47774
rect 24404 -48350 24438 -47774
rect 25422 -48350 25456 -47774
rect 28026 -48030 28060 -47454
rect 29044 -48030 29078 -47454
rect 30062 -48030 30096 -47454
rect 31080 -48030 31114 -47454
rect 32098 -48030 32132 -47454
rect 33116 -48030 33150 -47454
rect 34134 -48030 34168 -47454
rect 35152 -48030 35186 -47454
rect 36170 -48030 36204 -47454
rect 37188 -48030 37222 -47454
rect 38206 -48030 38240 -47454
rect 39224 -48030 39258 -47454
rect 40242 -48030 40276 -47454
rect 41260 -48030 41294 -47454
rect 42278 -48030 42312 -47454
rect 43296 -48030 43330 -47454
rect 44314 -48030 44348 -47454
rect 45332 -48030 45366 -47454
rect 46350 -48030 46384 -47454
rect 47368 -48030 47402 -47454
rect 48386 -48030 48420 -47454
rect 28320 -48114 28784 -48080
rect 29338 -48114 29802 -48080
rect 30356 -48114 30820 -48080
rect 31374 -48114 31838 -48080
rect 32392 -48114 32856 -48080
rect 33410 -48114 33874 -48080
rect 34428 -48114 34892 -48080
rect 35446 -48114 35910 -48080
rect 36464 -48114 36928 -48080
rect 37482 -48114 37946 -48080
rect 38500 -48114 38964 -48080
rect 39518 -48114 39982 -48080
rect 40536 -48114 41000 -48080
rect 41554 -48114 42018 -48080
rect 42572 -48114 43036 -48080
rect 43590 -48114 44054 -48080
rect 44608 -48114 45072 -48080
rect 45626 -48114 46090 -48080
rect 46644 -48114 47108 -48080
rect 47662 -48114 48126 -48080
rect 16554 -48434 17018 -48400
rect 17572 -48434 18036 -48400
rect 16554 -48542 17018 -48508
rect 18590 -48434 19054 -48400
rect 17572 -48542 18036 -48508
rect 19608 -48434 20072 -48400
rect 18590 -48542 19054 -48508
rect 20626 -48434 21090 -48400
rect 19608 -48542 20072 -48508
rect 21644 -48434 22108 -48400
rect 20626 -48542 21090 -48508
rect 22662 -48434 23126 -48400
rect 21644 -48542 22108 -48508
rect 23680 -48434 24144 -48400
rect 22662 -48542 23126 -48508
rect 24698 -48434 25162 -48400
rect 23680 -48542 24144 -48508
rect 24698 -48542 25162 -48508
rect 16260 -49168 16294 -48592
rect 17278 -49168 17312 -48592
rect 18296 -49168 18330 -48592
rect 19314 -49168 19348 -48592
rect 20332 -49168 20366 -48592
rect 21350 -49168 21384 -48592
rect 22368 -49168 22402 -48592
rect 23386 -49168 23420 -48592
rect 24404 -49168 24438 -48592
rect 25422 -49168 25456 -48592
rect 28318 -48638 28782 -48604
rect 29336 -48638 29800 -48604
rect 30354 -48638 30818 -48604
rect 31372 -48638 31836 -48604
rect 32390 -48638 32854 -48604
rect 33408 -48638 33872 -48604
rect 34426 -48638 34890 -48604
rect 35444 -48638 35908 -48604
rect 36462 -48638 36926 -48604
rect 37480 -48638 37944 -48604
rect 38498 -48638 38962 -48604
rect 39516 -48638 39980 -48604
rect 40534 -48638 40998 -48604
rect 41552 -48638 42016 -48604
rect 42570 -48638 43034 -48604
rect 43588 -48638 44052 -48604
rect 44606 -48638 45070 -48604
rect 45624 -48638 46088 -48604
rect 46642 -48638 47106 -48604
rect 47660 -48638 48124 -48604
rect 16554 -49252 17018 -49218
rect 17572 -49252 18036 -49218
rect 16554 -49360 17018 -49326
rect 18590 -49252 19054 -49218
rect 17572 -49360 18036 -49326
rect 19608 -49252 20072 -49218
rect 18590 -49360 19054 -49326
rect 20626 -49252 21090 -49218
rect 19608 -49360 20072 -49326
rect 21644 -49252 22108 -49218
rect 20626 -49360 21090 -49326
rect 22662 -49252 23126 -49218
rect 21644 -49360 22108 -49326
rect 23680 -49252 24144 -49218
rect 22662 -49360 23126 -49326
rect 24698 -49252 25162 -49218
rect 23680 -49360 24144 -49326
rect 28024 -49264 28058 -48688
rect 29042 -49264 29076 -48688
rect 30060 -49264 30094 -48688
rect 31078 -49264 31112 -48688
rect 32096 -49264 32130 -48688
rect 33114 -49264 33148 -48688
rect 34132 -49264 34166 -48688
rect 35150 -49264 35184 -48688
rect 36168 -49264 36202 -48688
rect 37186 -49264 37220 -48688
rect 38204 -49264 38238 -48688
rect 39222 -49264 39256 -48688
rect 40240 -49264 40274 -48688
rect 41258 -49264 41292 -48688
rect 42276 -49264 42310 -48688
rect 43294 -49264 43328 -48688
rect 44312 -49264 44346 -48688
rect 45330 -49264 45364 -48688
rect 46348 -49264 46382 -48688
rect 47366 -49264 47400 -48688
rect 48384 -49264 48418 -48688
rect 24698 -49360 25162 -49326
rect 28318 -49348 28782 -49314
rect 29336 -49348 29800 -49314
rect 30354 -49348 30818 -49314
rect 31372 -49348 31836 -49314
rect 32390 -49348 32854 -49314
rect 33408 -49348 33872 -49314
rect 34426 -49348 34890 -49314
rect 35444 -49348 35908 -49314
rect 36462 -49348 36926 -49314
rect 37480 -49348 37944 -49314
rect 38498 -49348 38962 -49314
rect 39516 -49348 39980 -49314
rect 40534 -49348 40998 -49314
rect 41552 -49348 42016 -49314
rect 42570 -49348 43034 -49314
rect 43588 -49348 44052 -49314
rect 44606 -49348 45070 -49314
rect 45624 -49348 46088 -49314
rect 46642 -49348 47106 -49314
rect 47660 -49348 48124 -49314
rect 16260 -49986 16294 -49410
rect 17278 -49986 17312 -49410
rect 18296 -49986 18330 -49410
rect 19314 -49986 19348 -49410
rect 20332 -49986 20366 -49410
rect 21350 -49986 21384 -49410
rect 22368 -49986 22402 -49410
rect 23386 -49986 23420 -49410
rect 24404 -49986 24438 -49410
rect 25422 -49986 25456 -49410
rect 28318 -49872 28782 -49838
rect 29336 -49872 29800 -49838
rect 30354 -49872 30818 -49838
rect 31372 -49872 31836 -49838
rect 32390 -49872 32854 -49838
rect 33408 -49872 33872 -49838
rect 34426 -49872 34890 -49838
rect 35444 -49872 35908 -49838
rect 36462 -49872 36926 -49838
rect 37480 -49872 37944 -49838
rect 38498 -49872 38962 -49838
rect 39516 -49872 39980 -49838
rect 40534 -49872 40998 -49838
rect 41552 -49872 42016 -49838
rect 42570 -49872 43034 -49838
rect 43588 -49872 44052 -49838
rect 44606 -49872 45070 -49838
rect 45624 -49872 46088 -49838
rect 46642 -49872 47106 -49838
rect 47660 -49872 48124 -49838
rect 16554 -50070 17018 -50036
rect 17572 -50070 18036 -50036
rect 16554 -50178 17018 -50144
rect 18590 -50070 19054 -50036
rect 17572 -50178 18036 -50144
rect 19608 -50070 20072 -50036
rect 18590 -50178 19054 -50144
rect 20626 -50070 21090 -50036
rect 19608 -50178 20072 -50144
rect 21644 -50070 22108 -50036
rect 20626 -50178 21090 -50144
rect 22662 -50070 23126 -50036
rect 21644 -50178 22108 -50144
rect 23680 -50070 24144 -50036
rect 22662 -50178 23126 -50144
rect 24698 -50070 25162 -50036
rect 23680 -50178 24144 -50144
rect 24698 -50178 25162 -50144
rect 16260 -50804 16294 -50228
rect 17278 -50804 17312 -50228
rect 18296 -50804 18330 -50228
rect 19314 -50804 19348 -50228
rect 20332 -50804 20366 -50228
rect 21350 -50804 21384 -50228
rect 22368 -50804 22402 -50228
rect 23386 -50804 23420 -50228
rect 24404 -50804 24438 -50228
rect 25422 -50804 25456 -50228
rect 28024 -50498 28058 -49922
rect 29042 -50498 29076 -49922
rect 30060 -50498 30094 -49922
rect 31078 -50498 31112 -49922
rect 32096 -50498 32130 -49922
rect 33114 -50498 33148 -49922
rect 34132 -50498 34166 -49922
rect 35150 -50498 35184 -49922
rect 36168 -50498 36202 -49922
rect 37186 -50498 37220 -49922
rect 38204 -50498 38238 -49922
rect 39222 -50498 39256 -49922
rect 40240 -50498 40274 -49922
rect 41258 -50498 41292 -49922
rect 42276 -50498 42310 -49922
rect 43294 -50498 43328 -49922
rect 44312 -50498 44346 -49922
rect 45330 -50498 45364 -49922
rect 46348 -50498 46382 -49922
rect 47366 -50498 47400 -49922
rect 48384 -50498 48418 -49922
rect 28318 -50582 28782 -50548
rect 29336 -50582 29800 -50548
rect 30354 -50582 30818 -50548
rect 31372 -50582 31836 -50548
rect 32390 -50582 32854 -50548
rect 33408 -50582 33872 -50548
rect 34426 -50582 34890 -50548
rect 35444 -50582 35908 -50548
rect 36462 -50582 36926 -50548
rect 37480 -50582 37944 -50548
rect 38498 -50582 38962 -50548
rect 39516 -50582 39980 -50548
rect 40534 -50582 40998 -50548
rect 41552 -50582 42016 -50548
rect 42570 -50582 43034 -50548
rect 43588 -50582 44052 -50548
rect 44606 -50582 45070 -50548
rect 45624 -50582 46088 -50548
rect 46642 -50582 47106 -50548
rect 47660 -50582 48124 -50548
rect 16554 -50888 17018 -50854
rect 17572 -50888 18036 -50854
rect 18590 -50888 19054 -50854
rect 19608 -50888 20072 -50854
rect 20626 -50888 21090 -50854
rect 21644 -50888 22108 -50854
rect 22662 -50888 23126 -50854
rect 23680 -50888 24144 -50854
rect 24698 -50888 25162 -50854
rect 28318 -51104 28782 -51070
rect 29336 -51104 29800 -51070
rect 30354 -51104 30818 -51070
rect 31372 -51104 31836 -51070
rect 32390 -51104 32854 -51070
rect 33408 -51104 33872 -51070
rect 34426 -51104 34890 -51070
rect 35444 -51104 35908 -51070
rect 36462 -51104 36926 -51070
rect 37480 -51104 37944 -51070
rect 38498 -51104 38962 -51070
rect 39516 -51104 39980 -51070
rect 40534 -51104 40998 -51070
rect 41552 -51104 42016 -51070
rect 42570 -51104 43034 -51070
rect 43588 -51104 44052 -51070
rect 44606 -51104 45070 -51070
rect 45624 -51104 46088 -51070
rect 46642 -51104 47106 -51070
rect 47660 -51104 48124 -51070
rect 28024 -51730 28058 -51154
rect 29042 -51730 29076 -51154
rect 30060 -51730 30094 -51154
rect 31078 -51730 31112 -51154
rect 32096 -51730 32130 -51154
rect 33114 -51730 33148 -51154
rect 34132 -51730 34166 -51154
rect 35150 -51730 35184 -51154
rect 36168 -51730 36202 -51154
rect 37186 -51730 37220 -51154
rect 38204 -51730 38238 -51154
rect 39222 -51730 39256 -51154
rect 40240 -51730 40274 -51154
rect 41258 -51730 41292 -51154
rect 42276 -51730 42310 -51154
rect 43294 -51730 43328 -51154
rect 44312 -51730 44346 -51154
rect 45330 -51730 45364 -51154
rect 46348 -51730 46382 -51154
rect 47366 -51730 47400 -51154
rect 48384 -51730 48418 -51154
rect 28318 -51814 28782 -51780
rect 29336 -51814 29800 -51780
rect 30354 -51814 30818 -51780
rect 31372 -51814 31836 -51780
rect 32390 -51814 32854 -51780
rect 33408 -51814 33872 -51780
rect 34426 -51814 34890 -51780
rect 35444 -51814 35908 -51780
rect 36462 -51814 36926 -51780
rect 37480 -51814 37944 -51780
rect 38498 -51814 38962 -51780
rect 39516 -51814 39980 -51780
rect 40534 -51814 40998 -51780
rect 41552 -51814 42016 -51780
rect 42570 -51814 43034 -51780
rect 43588 -51814 44052 -51780
rect 44606 -51814 45070 -51780
rect 45624 -51814 46088 -51780
rect 46642 -51814 47106 -51780
rect 47660 -51814 48124 -51780
rect 15230 -52202 15694 -52168
rect 16248 -52202 16712 -52168
rect 17266 -52202 17730 -52168
rect 18284 -52202 18748 -52168
rect 19302 -52202 19766 -52168
rect 20320 -52202 20784 -52168
rect 21338 -52202 21802 -52168
rect 22356 -52202 22820 -52168
rect 23374 -52202 23838 -52168
rect 24392 -52202 24856 -52168
rect 25410 -52202 25874 -52168
rect 14936 -52828 14970 -52252
rect 15954 -52828 15988 -52252
rect 16972 -52828 17006 -52252
rect 17990 -52828 18024 -52252
rect 19008 -52828 19042 -52252
rect 20026 -52828 20060 -52252
rect 21044 -52828 21078 -52252
rect 22062 -52828 22096 -52252
rect 23080 -52828 23114 -52252
rect 24098 -52828 24132 -52252
rect 25116 -52828 25150 -52252
rect 26134 -52828 26168 -52252
rect 28318 -52338 28782 -52304
rect 29336 -52338 29800 -52304
rect 30354 -52338 30818 -52304
rect 31372 -52338 31836 -52304
rect 32390 -52338 32854 -52304
rect 33408 -52338 33872 -52304
rect 34426 -52338 34890 -52304
rect 35444 -52338 35908 -52304
rect 36462 -52338 36926 -52304
rect 37480 -52338 37944 -52304
rect 38498 -52338 38962 -52304
rect 39516 -52338 39980 -52304
rect 40534 -52338 40998 -52304
rect 41552 -52338 42016 -52304
rect 42570 -52338 43034 -52304
rect 43588 -52338 44052 -52304
rect 44606 -52338 45070 -52304
rect 45624 -52338 46088 -52304
rect 46642 -52338 47106 -52304
rect 47660 -52338 48124 -52304
rect 15230 -52912 15694 -52878
rect 16248 -52912 16712 -52878
rect 17266 -52912 17730 -52878
rect 18284 -52912 18748 -52878
rect 19302 -52912 19766 -52878
rect 20320 -52912 20784 -52878
rect 21338 -52912 21802 -52878
rect 22356 -52912 22820 -52878
rect 23374 -52912 23838 -52878
rect 24392 -52912 24856 -52878
rect 25410 -52912 25874 -52878
rect 28024 -52964 28058 -52388
rect 29042 -52964 29076 -52388
rect 30060 -52964 30094 -52388
rect 31078 -52964 31112 -52388
rect 32096 -52964 32130 -52388
rect 33114 -52964 33148 -52388
rect 34132 -52964 34166 -52388
rect 35150 -52964 35184 -52388
rect 36168 -52964 36202 -52388
rect 37186 -52964 37220 -52388
rect 38204 -52964 38238 -52388
rect 39222 -52964 39256 -52388
rect 40240 -52964 40274 -52388
rect 41258 -52964 41292 -52388
rect 42276 -52964 42310 -52388
rect 43294 -52964 43328 -52388
rect 44312 -52964 44346 -52388
rect 45330 -52964 45364 -52388
rect 46348 -52964 46382 -52388
rect 47366 -52964 47400 -52388
rect 48384 -52964 48418 -52388
rect 28318 -53048 28782 -53014
rect 29336 -53048 29800 -53014
rect 30354 -53048 30818 -53014
rect 31372 -53048 31836 -53014
rect 32390 -53048 32854 -53014
rect 33408 -53048 33872 -53014
rect 34426 -53048 34890 -53014
rect 35444 -53048 35908 -53014
rect 36462 -53048 36926 -53014
rect 37480 -53048 37944 -53014
rect 38498 -53048 38962 -53014
rect 39516 -53048 39980 -53014
rect 40534 -53048 40998 -53014
rect 41552 -53048 42016 -53014
rect 42570 -53048 43034 -53014
rect 43588 -53048 44052 -53014
rect 44606 -53048 45070 -53014
rect 45624 -53048 46088 -53014
rect 46642 -53048 47106 -53014
rect 47660 -53048 48124 -53014
rect 15230 -53314 15694 -53280
rect 16248 -53314 16712 -53280
rect 17266 -53314 17730 -53280
rect 18284 -53314 18748 -53280
rect 19302 -53314 19766 -53280
rect 20320 -53314 20784 -53280
rect 21338 -53314 21802 -53280
rect 22356 -53314 22820 -53280
rect 23374 -53314 23838 -53280
rect 24392 -53314 24856 -53280
rect 25410 -53314 25874 -53280
rect 14936 -53940 14970 -53364
rect 15954 -53940 15988 -53364
rect 16972 -53940 17006 -53364
rect 17990 -53940 18024 -53364
rect 19008 -53940 19042 -53364
rect 20026 -53940 20060 -53364
rect 21044 -53940 21078 -53364
rect 22062 -53940 22096 -53364
rect 23080 -53940 23114 -53364
rect 24098 -53940 24132 -53364
rect 25116 -53940 25150 -53364
rect 26134 -53940 26168 -53364
rect 28318 -53572 28782 -53538
rect 29336 -53572 29800 -53538
rect 30354 -53572 30818 -53538
rect 31372 -53572 31836 -53538
rect 32390 -53572 32854 -53538
rect 33408 -53572 33872 -53538
rect 34426 -53572 34890 -53538
rect 35444 -53572 35908 -53538
rect 36462 -53572 36926 -53538
rect 37480 -53572 37944 -53538
rect 38498 -53572 38962 -53538
rect 39516 -53572 39980 -53538
rect 40534 -53572 40998 -53538
rect 41552 -53572 42016 -53538
rect 42570 -53572 43034 -53538
rect 43588 -53572 44052 -53538
rect 44606 -53572 45070 -53538
rect 45624 -53572 46088 -53538
rect 46642 -53572 47106 -53538
rect 47660 -53572 48124 -53538
rect 15230 -54024 15694 -53990
rect 16248 -54024 16712 -53990
rect 17266 -54024 17730 -53990
rect 18284 -54024 18748 -53990
rect 19302 -54024 19766 -53990
rect 20320 -54024 20784 -53990
rect 21338 -54024 21802 -53990
rect 22356 -54024 22820 -53990
rect 23374 -54024 23838 -53990
rect 24392 -54024 24856 -53990
rect 25410 -54024 25874 -53990
rect 28024 -54198 28058 -53622
rect 29042 -54198 29076 -53622
rect 30060 -54198 30094 -53622
rect 31078 -54198 31112 -53622
rect 32096 -54198 32130 -53622
rect 33114 -54198 33148 -53622
rect 34132 -54198 34166 -53622
rect 35150 -54198 35184 -53622
rect 36168 -54198 36202 -53622
rect 37186 -54198 37220 -53622
rect 38204 -54198 38238 -53622
rect 39222 -54198 39256 -53622
rect 40240 -54198 40274 -53622
rect 41258 -54198 41292 -53622
rect 42276 -54198 42310 -53622
rect 43294 -54198 43328 -53622
rect 44312 -54198 44346 -53622
rect 45330 -54198 45364 -53622
rect 46348 -54198 46382 -53622
rect 47366 -54198 47400 -53622
rect 48384 -54198 48418 -53622
rect 28318 -54282 28782 -54248
rect 29336 -54282 29800 -54248
rect 30354 -54282 30818 -54248
rect 31372 -54282 31836 -54248
rect 32390 -54282 32854 -54248
rect 33408 -54282 33872 -54248
rect 34426 -54282 34890 -54248
rect 35444 -54282 35908 -54248
rect 36462 -54282 36926 -54248
rect 37480 -54282 37944 -54248
rect 38498 -54282 38962 -54248
rect 39516 -54282 39980 -54248
rect 40534 -54282 40998 -54248
rect 41552 -54282 42016 -54248
rect 42570 -54282 43034 -54248
rect 43588 -54282 44052 -54248
rect 44606 -54282 45070 -54248
rect 45624 -54282 46088 -54248
rect 46642 -54282 47106 -54248
rect 47660 -54282 48124 -54248
rect 15230 -54426 15694 -54392
rect 16248 -54426 16712 -54392
rect 17266 -54426 17730 -54392
rect 18284 -54426 18748 -54392
rect 19302 -54426 19766 -54392
rect 20320 -54426 20784 -54392
rect 21338 -54426 21802 -54392
rect 22356 -54426 22820 -54392
rect 23374 -54426 23838 -54392
rect 24392 -54426 24856 -54392
rect 25410 -54426 25874 -54392
rect 14936 -55052 14970 -54476
rect 15954 -55052 15988 -54476
rect 16972 -55052 17006 -54476
rect 17990 -55052 18024 -54476
rect 19008 -55052 19042 -54476
rect 20026 -55052 20060 -54476
rect 21044 -55052 21078 -54476
rect 22062 -55052 22096 -54476
rect 23080 -55052 23114 -54476
rect 24098 -55052 24132 -54476
rect 25116 -55052 25150 -54476
rect 26134 -55052 26168 -54476
rect 28318 -54804 28782 -54770
rect 29336 -54804 29800 -54770
rect 30354 -54804 30818 -54770
rect 31372 -54804 31836 -54770
rect 32390 -54804 32854 -54770
rect 33408 -54804 33872 -54770
rect 34426 -54804 34890 -54770
rect 35444 -54804 35908 -54770
rect 36462 -54804 36926 -54770
rect 37480 -54804 37944 -54770
rect 38498 -54804 38962 -54770
rect 39516 -54804 39980 -54770
rect 40534 -54804 40998 -54770
rect 41552 -54804 42016 -54770
rect 42570 -54804 43034 -54770
rect 43588 -54804 44052 -54770
rect 44606 -54804 45070 -54770
rect 45624 -54804 46088 -54770
rect 46642 -54804 47106 -54770
rect 47660 -54804 48124 -54770
rect 15230 -55136 15694 -55102
rect 16248 -55136 16712 -55102
rect 17266 -55136 17730 -55102
rect 18284 -55136 18748 -55102
rect 19302 -55136 19766 -55102
rect 20320 -55136 20784 -55102
rect 21338 -55136 21802 -55102
rect 22356 -55136 22820 -55102
rect 23374 -55136 23838 -55102
rect 24392 -55136 24856 -55102
rect 25410 -55136 25874 -55102
rect 28024 -55430 28058 -54854
rect 29042 -55430 29076 -54854
rect 30060 -55430 30094 -54854
rect 31078 -55430 31112 -54854
rect 32096 -55430 32130 -54854
rect 33114 -55430 33148 -54854
rect 34132 -55430 34166 -54854
rect 35150 -55430 35184 -54854
rect 36168 -55430 36202 -54854
rect 37186 -55430 37220 -54854
rect 38204 -55430 38238 -54854
rect 39222 -55430 39256 -54854
rect 40240 -55430 40274 -54854
rect 41258 -55430 41292 -54854
rect 42276 -55430 42310 -54854
rect 43294 -55430 43328 -54854
rect 44312 -55430 44346 -54854
rect 45330 -55430 45364 -54854
rect 46348 -55430 46382 -54854
rect 47366 -55430 47400 -54854
rect 48384 -55430 48418 -54854
rect 15230 -55538 15694 -55504
rect 16248 -55538 16712 -55504
rect 17266 -55538 17730 -55504
rect 18284 -55538 18748 -55504
rect 19302 -55538 19766 -55504
rect 20320 -55538 20784 -55504
rect 21338 -55538 21802 -55504
rect 22356 -55538 22820 -55504
rect 23374 -55538 23838 -55504
rect 24392 -55538 24856 -55504
rect 25410 -55538 25874 -55504
rect 28318 -55514 28782 -55480
rect 29336 -55514 29800 -55480
rect 30354 -55514 30818 -55480
rect 31372 -55514 31836 -55480
rect 32390 -55514 32854 -55480
rect 33408 -55514 33872 -55480
rect 34426 -55514 34890 -55480
rect 35444 -55514 35908 -55480
rect 36462 -55514 36926 -55480
rect 37480 -55514 37944 -55480
rect 38498 -55514 38962 -55480
rect 39516 -55514 39980 -55480
rect 40534 -55514 40998 -55480
rect 41552 -55514 42016 -55480
rect 42570 -55514 43034 -55480
rect 43588 -55514 44052 -55480
rect 44606 -55514 45070 -55480
rect 45624 -55514 46088 -55480
rect 46642 -55514 47106 -55480
rect 47660 -55514 48124 -55480
rect 14936 -56164 14970 -55588
rect 15954 -56164 15988 -55588
rect 16972 -56164 17006 -55588
rect 17990 -56164 18024 -55588
rect 19008 -56164 19042 -55588
rect 20026 -56164 20060 -55588
rect 21044 -56164 21078 -55588
rect 22062 -56164 22096 -55588
rect 23080 -56164 23114 -55588
rect 24098 -56164 24132 -55588
rect 25116 -56164 25150 -55588
rect 26134 -56164 26168 -55588
rect 28318 -56038 28782 -56004
rect 29336 -56038 29800 -56004
rect 30354 -56038 30818 -56004
rect 31372 -56038 31836 -56004
rect 32390 -56038 32854 -56004
rect 33408 -56038 33872 -56004
rect 34426 -56038 34890 -56004
rect 35444 -56038 35908 -56004
rect 36462 -56038 36926 -56004
rect 37480 -56038 37944 -56004
rect 38498 -56038 38962 -56004
rect 39516 -56038 39980 -56004
rect 40534 -56038 40998 -56004
rect 41552 -56038 42016 -56004
rect 42570 -56038 43034 -56004
rect 43588 -56038 44052 -56004
rect 44606 -56038 45070 -56004
rect 45624 -56038 46088 -56004
rect 46642 -56038 47106 -56004
rect 47660 -56038 48124 -56004
rect 15230 -56248 15694 -56214
rect 16248 -56248 16712 -56214
rect 17266 -56248 17730 -56214
rect 18284 -56248 18748 -56214
rect 19302 -56248 19766 -56214
rect 20320 -56248 20784 -56214
rect 21338 -56248 21802 -56214
rect 22356 -56248 22820 -56214
rect 23374 -56248 23838 -56214
rect 24392 -56248 24856 -56214
rect 25410 -56248 25874 -56214
rect 28024 -56664 28058 -56088
rect 29042 -56664 29076 -56088
rect 30060 -56664 30094 -56088
rect 31078 -56664 31112 -56088
rect 32096 -56664 32130 -56088
rect 33114 -56664 33148 -56088
rect 34132 -56664 34166 -56088
rect 35150 -56664 35184 -56088
rect 36168 -56664 36202 -56088
rect 37186 -56664 37220 -56088
rect 38204 -56664 38238 -56088
rect 39222 -56664 39256 -56088
rect 40240 -56664 40274 -56088
rect 41258 -56664 41292 -56088
rect 42276 -56664 42310 -56088
rect 43294 -56664 43328 -56088
rect 44312 -56664 44346 -56088
rect 45330 -56664 45364 -56088
rect 46348 -56664 46382 -56088
rect 47366 -56664 47400 -56088
rect 48384 -56664 48418 -56088
rect 28318 -56748 28782 -56714
rect 29336 -56748 29800 -56714
rect 30354 -56748 30818 -56714
rect 31372 -56748 31836 -56714
rect 32390 -56748 32854 -56714
rect 33408 -56748 33872 -56714
rect 34426 -56748 34890 -56714
rect 35444 -56748 35908 -56714
rect 36462 -56748 36926 -56714
rect 37480 -56748 37944 -56714
rect 38498 -56748 38962 -56714
rect 39516 -56748 39980 -56714
rect 40534 -56748 40998 -56714
rect 41552 -56748 42016 -56714
rect 42570 -56748 43034 -56714
rect 43588 -56748 44052 -56714
rect 44606 -56748 45070 -56714
rect 45624 -56748 46088 -56714
rect 46642 -56748 47106 -56714
rect 47660 -56748 48124 -56714
rect 15688 -57080 16152 -57046
rect 16706 -57080 17170 -57046
rect 17724 -57080 18188 -57046
rect 18742 -57080 19206 -57046
rect 19760 -57080 20224 -57046
rect 20778 -57080 21242 -57046
rect 21796 -57080 22260 -57046
rect 22814 -57080 23278 -57046
rect 23832 -57080 24296 -57046
rect 24850 -57080 25314 -57046
rect 15394 -57706 15428 -57130
rect 16412 -57706 16446 -57130
rect 17430 -57706 17464 -57130
rect 18448 -57706 18482 -57130
rect 19466 -57706 19500 -57130
rect 20484 -57706 20518 -57130
rect 21502 -57706 21536 -57130
rect 22520 -57706 22554 -57130
rect 23538 -57706 23572 -57130
rect 24556 -57706 24590 -57130
rect 25574 -57706 25608 -57130
rect 28318 -57270 28782 -57236
rect 29336 -57270 29800 -57236
rect 30354 -57270 30818 -57236
rect 31372 -57270 31836 -57236
rect 32390 -57270 32854 -57236
rect 33408 -57270 33872 -57236
rect 34426 -57270 34890 -57236
rect 35444 -57270 35908 -57236
rect 36462 -57270 36926 -57236
rect 37480 -57270 37944 -57236
rect 38498 -57270 38962 -57236
rect 39516 -57270 39980 -57236
rect 40534 -57270 40998 -57236
rect 41552 -57270 42016 -57236
rect 42570 -57270 43034 -57236
rect 43588 -57270 44052 -57236
rect 44606 -57270 45070 -57236
rect 45624 -57270 46088 -57236
rect 46642 -57270 47106 -57236
rect 47660 -57270 48124 -57236
rect 15688 -57790 16152 -57756
rect 16706 -57790 17170 -57756
rect 17724 -57790 18188 -57756
rect 18742 -57790 19206 -57756
rect 19760 -57790 20224 -57756
rect 20778 -57790 21242 -57756
rect 21796 -57790 22260 -57756
rect 22814 -57790 23278 -57756
rect 23832 -57790 24296 -57756
rect 24850 -57790 25314 -57756
rect 28024 -57896 28058 -57320
rect 29042 -57896 29076 -57320
rect 30060 -57896 30094 -57320
rect 31078 -57896 31112 -57320
rect 32096 -57896 32130 -57320
rect 33114 -57896 33148 -57320
rect 34132 -57896 34166 -57320
rect 35150 -57896 35184 -57320
rect 36168 -57896 36202 -57320
rect 37186 -57896 37220 -57320
rect 38204 -57896 38238 -57320
rect 39222 -57896 39256 -57320
rect 40240 -57896 40274 -57320
rect 41258 -57896 41292 -57320
rect 42276 -57896 42310 -57320
rect 43294 -57896 43328 -57320
rect 44312 -57896 44346 -57320
rect 45330 -57896 45364 -57320
rect 46348 -57896 46382 -57320
rect 47366 -57896 47400 -57320
rect 48384 -57896 48418 -57320
rect 28318 -57980 28782 -57946
rect 29336 -57980 29800 -57946
rect 30354 -57980 30818 -57946
rect 31372 -57980 31836 -57946
rect 32390 -57980 32854 -57946
rect 33408 -57980 33872 -57946
rect 34426 -57980 34890 -57946
rect 35444 -57980 35908 -57946
rect 36462 -57980 36926 -57946
rect 37480 -57980 37944 -57946
rect 38498 -57980 38962 -57946
rect 39516 -57980 39980 -57946
rect 40534 -57980 40998 -57946
rect 41552 -57980 42016 -57946
rect 42570 -57980 43034 -57946
rect 43588 -57980 44052 -57946
rect 44606 -57980 45070 -57946
rect 45624 -57980 46088 -57946
rect 46642 -57980 47106 -57946
rect 47660 -57980 48124 -57946
rect 50266 -58308 50366 -44048
rect 13222 -59200 13284 -59100
rect 13284 -59200 50204 -59100
rect 50204 -59200 50266 -59100
rect -27584 -64526 -27522 -64426
rect -27522 -64526 -25522 -64426
rect -25522 -64526 -25460 -64426
rect -28043 -67299 -28009 -67265
rect -27951 -67299 -27917 -67265
rect -27859 -67299 -27825 -67265
rect -27684 -67290 -27584 -64666
rect -27233 -65578 -27149 -65544
rect -26975 -65578 -26891 -65544
rect -26717 -65578 -26633 -65544
rect -26459 -65578 -26375 -65544
rect -26201 -65578 -26117 -65544
rect -25943 -65578 -25859 -65544
rect -27337 -66013 -27303 -65637
rect -27079 -66013 -27045 -65637
rect -26821 -66013 -26787 -65637
rect -26563 -66013 -26529 -65637
rect -26305 -66013 -26271 -65637
rect -26047 -66013 -26013 -65637
rect -25789 -66013 -25755 -65637
rect -27233 -66106 -27149 -66072
rect -26975 -66106 -26891 -66072
rect -26717 -66106 -26633 -66072
rect -26459 -66106 -26375 -66072
rect -26201 -66106 -26117 -66072
rect -25943 -66106 -25859 -66072
rect -27233 -66438 -27149 -66404
rect -26975 -66438 -26891 -66404
rect -26717 -66438 -26633 -66404
rect -26459 -66438 -26375 -66404
rect -26201 -66438 -26117 -66404
rect -25943 -66438 -25859 -66404
rect -27337 -66873 -27303 -66497
rect -27079 -66873 -27045 -66497
rect -26821 -66873 -26787 -66497
rect -26563 -66873 -26529 -66497
rect -26305 -66873 -26271 -66497
rect -26047 -66873 -26013 -66497
rect -25789 -66873 -25755 -66497
rect -27233 -66966 -27149 -66932
rect -26975 -66966 -26891 -66932
rect -26717 -66966 -26633 -66932
rect -26459 -66966 -26375 -66932
rect -26201 -66966 -26117 -66932
rect -25943 -66966 -25859 -66932
rect -28004 -67577 -27956 -67562
rect -28004 -67610 -27992 -67577
rect -27992 -67610 -27958 -67577
rect -27958 -67610 -27956 -67577
rect -25460 -67290 -25360 -64666
rect -23584 -64526 -23522 -64426
rect -23522 -64526 -21522 -64426
rect -21522 -64526 -21460 -64426
rect -24043 -67299 -24009 -67265
rect -23951 -67299 -23917 -67265
rect -23859 -67299 -23825 -67265
rect -23684 -67290 -23584 -64666
rect -23233 -65578 -23149 -65544
rect -22975 -65578 -22891 -65544
rect -22717 -65578 -22633 -65544
rect -22459 -65578 -22375 -65544
rect -22201 -65578 -22117 -65544
rect -21943 -65578 -21859 -65544
rect -23337 -66013 -23303 -65637
rect -23079 -66013 -23045 -65637
rect -22821 -66013 -22787 -65637
rect -22563 -66013 -22529 -65637
rect -22305 -66013 -22271 -65637
rect -22047 -66013 -22013 -65637
rect -21789 -66013 -21755 -65637
rect -23233 -66106 -23149 -66072
rect -22975 -66106 -22891 -66072
rect -22717 -66106 -22633 -66072
rect -22459 -66106 -22375 -66072
rect -22201 -66106 -22117 -66072
rect -21943 -66106 -21859 -66072
rect -23233 -66438 -23149 -66404
rect -22975 -66438 -22891 -66404
rect -22717 -66438 -22633 -66404
rect -22459 -66438 -22375 -66404
rect -22201 -66438 -22117 -66404
rect -21943 -66438 -21859 -66404
rect -23337 -66873 -23303 -66497
rect -23079 -66873 -23045 -66497
rect -22821 -66873 -22787 -66497
rect -22563 -66873 -22529 -66497
rect -22305 -66873 -22271 -66497
rect -22047 -66873 -22013 -66497
rect -21789 -66873 -21755 -66497
rect -23233 -66966 -23149 -66932
rect -22975 -66966 -22891 -66932
rect -22717 -66966 -22633 -66932
rect -22459 -66966 -22375 -66932
rect -22201 -66966 -22117 -66932
rect -21943 -66966 -21859 -66932
rect -27584 -67530 -27522 -67430
rect -27522 -67530 -25522 -67430
rect -25522 -67530 -25460 -67430
rect -24004 -67577 -23956 -67562
rect -24004 -67610 -23992 -67577
rect -23992 -67610 -23958 -67577
rect -23958 -67610 -23956 -67577
rect -21460 -67290 -21360 -64666
rect -19584 -64526 -19522 -64426
rect -19522 -64526 -17522 -64426
rect -17522 -64526 -17460 -64426
rect -20043 -67299 -20009 -67265
rect -19951 -67299 -19917 -67265
rect -19859 -67299 -19825 -67265
rect -19684 -67290 -19584 -64666
rect -19233 -65578 -19149 -65544
rect -18975 -65578 -18891 -65544
rect -18717 -65578 -18633 -65544
rect -18459 -65578 -18375 -65544
rect -18201 -65578 -18117 -65544
rect -17943 -65578 -17859 -65544
rect -19337 -66013 -19303 -65637
rect -19079 -66013 -19045 -65637
rect -18821 -66013 -18787 -65637
rect -18563 -66013 -18529 -65637
rect -18305 -66013 -18271 -65637
rect -18047 -66013 -18013 -65637
rect -17789 -66013 -17755 -65637
rect -19233 -66106 -19149 -66072
rect -18975 -66106 -18891 -66072
rect -18717 -66106 -18633 -66072
rect -18459 -66106 -18375 -66072
rect -18201 -66106 -18117 -66072
rect -17943 -66106 -17859 -66072
rect -19233 -66438 -19149 -66404
rect -18975 -66438 -18891 -66404
rect -18717 -66438 -18633 -66404
rect -18459 -66438 -18375 -66404
rect -18201 -66438 -18117 -66404
rect -17943 -66438 -17859 -66404
rect -19337 -66873 -19303 -66497
rect -19079 -66873 -19045 -66497
rect -18821 -66873 -18787 -66497
rect -18563 -66873 -18529 -66497
rect -18305 -66873 -18271 -66497
rect -18047 -66873 -18013 -66497
rect -17789 -66873 -17755 -66497
rect -19233 -66966 -19149 -66932
rect -18975 -66966 -18891 -66932
rect -18717 -66966 -18633 -66932
rect -18459 -66966 -18375 -66932
rect -18201 -66966 -18117 -66932
rect -17943 -66966 -17859 -66932
rect -23584 -67530 -23522 -67430
rect -23522 -67530 -21522 -67430
rect -21522 -67530 -21460 -67430
rect -20004 -67577 -19956 -67562
rect -20004 -67610 -19992 -67577
rect -19992 -67610 -19958 -67577
rect -19958 -67610 -19956 -67577
rect -17460 -67290 -17360 -64666
rect -15584 -64526 -15522 -64426
rect -15522 -64526 -13522 -64426
rect -13522 -64526 -13460 -64426
rect -16043 -67299 -16009 -67265
rect -15951 -67299 -15917 -67265
rect -15859 -67299 -15825 -67265
rect -15684 -67290 -15584 -64666
rect -15233 -65578 -15149 -65544
rect -14975 -65578 -14891 -65544
rect -14717 -65578 -14633 -65544
rect -14459 -65578 -14375 -65544
rect -14201 -65578 -14117 -65544
rect -13943 -65578 -13859 -65544
rect -15337 -66013 -15303 -65637
rect -15079 -66013 -15045 -65637
rect -14821 -66013 -14787 -65637
rect -14563 -66013 -14529 -65637
rect -14305 -66013 -14271 -65637
rect -14047 -66013 -14013 -65637
rect -13789 -66013 -13755 -65637
rect -15233 -66106 -15149 -66072
rect -14975 -66106 -14891 -66072
rect -14717 -66106 -14633 -66072
rect -14459 -66106 -14375 -66072
rect -14201 -66106 -14117 -66072
rect -13943 -66106 -13859 -66072
rect -15233 -66438 -15149 -66404
rect -14975 -66438 -14891 -66404
rect -14717 -66438 -14633 -66404
rect -14459 -66438 -14375 -66404
rect -14201 -66438 -14117 -66404
rect -13943 -66438 -13859 -66404
rect -15337 -66873 -15303 -66497
rect -15079 -66873 -15045 -66497
rect -14821 -66873 -14787 -66497
rect -14563 -66873 -14529 -66497
rect -14305 -66873 -14271 -66497
rect -14047 -66873 -14013 -66497
rect -13789 -66873 -13755 -66497
rect -15233 -66966 -15149 -66932
rect -14975 -66966 -14891 -66932
rect -14717 -66966 -14633 -66932
rect -14459 -66966 -14375 -66932
rect -14201 -66966 -14117 -66932
rect -13943 -66966 -13859 -66932
rect -19584 -67530 -19522 -67430
rect -19522 -67530 -17522 -67430
rect -17522 -67530 -17460 -67430
rect -16004 -67577 -15956 -67562
rect -16004 -67610 -15992 -67577
rect -15992 -67610 -15958 -67577
rect -15958 -67610 -15956 -67577
rect -13460 -67290 -13360 -64666
rect -11584 -64526 -11522 -64426
rect -11522 -64526 -9522 -64426
rect -9522 -64526 -9460 -64426
rect -12043 -67299 -12009 -67265
rect -11951 -67299 -11917 -67265
rect -11859 -67299 -11825 -67265
rect -11684 -67290 -11584 -64666
rect -11233 -65578 -11149 -65544
rect -10975 -65578 -10891 -65544
rect -10717 -65578 -10633 -65544
rect -10459 -65578 -10375 -65544
rect -10201 -65578 -10117 -65544
rect -9943 -65578 -9859 -65544
rect -11337 -66013 -11303 -65637
rect -11079 -66013 -11045 -65637
rect -10821 -66013 -10787 -65637
rect -10563 -66013 -10529 -65637
rect -10305 -66013 -10271 -65637
rect -10047 -66013 -10013 -65637
rect -9789 -66013 -9755 -65637
rect -11233 -66106 -11149 -66072
rect -10975 -66106 -10891 -66072
rect -10717 -66106 -10633 -66072
rect -10459 -66106 -10375 -66072
rect -10201 -66106 -10117 -66072
rect -9943 -66106 -9859 -66072
rect -11233 -66438 -11149 -66404
rect -10975 -66438 -10891 -66404
rect -10717 -66438 -10633 -66404
rect -10459 -66438 -10375 -66404
rect -10201 -66438 -10117 -66404
rect -9943 -66438 -9859 -66404
rect -11337 -66873 -11303 -66497
rect -11079 -66873 -11045 -66497
rect -10821 -66873 -10787 -66497
rect -10563 -66873 -10529 -66497
rect -10305 -66873 -10271 -66497
rect -10047 -66873 -10013 -66497
rect -9789 -66873 -9755 -66497
rect -11233 -66966 -11149 -66932
rect -10975 -66966 -10891 -66932
rect -10717 -66966 -10633 -66932
rect -10459 -66966 -10375 -66932
rect -10201 -66966 -10117 -66932
rect -9943 -66966 -9859 -66932
rect -15584 -67530 -15522 -67430
rect -15522 -67530 -13522 -67430
rect -13522 -67530 -13460 -67430
rect -12004 -67577 -11956 -67562
rect -12004 -67610 -11992 -67577
rect -11992 -67610 -11958 -67577
rect -11958 -67610 -11956 -67577
rect -9460 -67290 -9360 -64666
rect -7584 -64526 -7522 -64426
rect -7522 -64526 -5522 -64426
rect -5522 -64526 -5460 -64426
rect -8043 -67299 -8009 -67265
rect -7951 -67299 -7917 -67265
rect -7859 -67299 -7825 -67265
rect -7684 -67290 -7584 -64666
rect -7233 -65578 -7149 -65544
rect -6975 -65578 -6891 -65544
rect -6717 -65578 -6633 -65544
rect -6459 -65578 -6375 -65544
rect -6201 -65578 -6117 -65544
rect -5943 -65578 -5859 -65544
rect -7337 -66013 -7303 -65637
rect -7079 -66013 -7045 -65637
rect -6821 -66013 -6787 -65637
rect -6563 -66013 -6529 -65637
rect -6305 -66013 -6271 -65637
rect -6047 -66013 -6013 -65637
rect -5789 -66013 -5755 -65637
rect -7233 -66106 -7149 -66072
rect -6975 -66106 -6891 -66072
rect -6717 -66106 -6633 -66072
rect -6459 -66106 -6375 -66072
rect -6201 -66106 -6117 -66072
rect -5943 -66106 -5859 -66072
rect -7233 -66438 -7149 -66404
rect -6975 -66438 -6891 -66404
rect -6717 -66438 -6633 -66404
rect -6459 -66438 -6375 -66404
rect -6201 -66438 -6117 -66404
rect -5943 -66438 -5859 -66404
rect -7337 -66873 -7303 -66497
rect -7079 -66873 -7045 -66497
rect -6821 -66873 -6787 -66497
rect -6563 -66873 -6529 -66497
rect -6305 -66873 -6271 -66497
rect -6047 -66873 -6013 -66497
rect -5789 -66873 -5755 -66497
rect -7233 -66966 -7149 -66932
rect -6975 -66966 -6891 -66932
rect -6717 -66966 -6633 -66932
rect -6459 -66966 -6375 -66932
rect -6201 -66966 -6117 -66932
rect -5943 -66966 -5859 -66932
rect -11584 -67530 -11522 -67430
rect -11522 -67530 -9522 -67430
rect -9522 -67530 -9460 -67430
rect -8004 -67577 -7956 -67562
rect -8004 -67610 -7992 -67577
rect -7992 -67610 -7958 -67577
rect -7958 -67610 -7956 -67577
rect -5460 -67290 -5360 -64666
rect -3584 -64526 -3522 -64426
rect -3522 -64526 -1522 -64426
rect -1522 -64526 -1460 -64426
rect -4043 -67299 -4009 -67265
rect -3951 -67299 -3917 -67265
rect -3859 -67299 -3825 -67265
rect -3684 -67290 -3584 -64666
rect -3233 -65578 -3149 -65544
rect -2975 -65578 -2891 -65544
rect -2717 -65578 -2633 -65544
rect -2459 -65578 -2375 -65544
rect -2201 -65578 -2117 -65544
rect -1943 -65578 -1859 -65544
rect -3337 -66013 -3303 -65637
rect -3079 -66013 -3045 -65637
rect -2821 -66013 -2787 -65637
rect -2563 -66013 -2529 -65637
rect -2305 -66013 -2271 -65637
rect -2047 -66013 -2013 -65637
rect -1789 -66013 -1755 -65637
rect -3233 -66106 -3149 -66072
rect -2975 -66106 -2891 -66072
rect -2717 -66106 -2633 -66072
rect -2459 -66106 -2375 -66072
rect -2201 -66106 -2117 -66072
rect -1943 -66106 -1859 -66072
rect -3233 -66438 -3149 -66404
rect -2975 -66438 -2891 -66404
rect -2717 -66438 -2633 -66404
rect -2459 -66438 -2375 -66404
rect -2201 -66438 -2117 -66404
rect -1943 -66438 -1859 -66404
rect -3337 -66873 -3303 -66497
rect -3079 -66873 -3045 -66497
rect -2821 -66873 -2787 -66497
rect -2563 -66873 -2529 -66497
rect -2305 -66873 -2271 -66497
rect -2047 -66873 -2013 -66497
rect -1789 -66873 -1755 -66497
rect -3233 -66966 -3149 -66932
rect -2975 -66966 -2891 -66932
rect -2717 -66966 -2633 -66932
rect -2459 -66966 -2375 -66932
rect -2201 -66966 -2117 -66932
rect -1943 -66966 -1859 -66932
rect -7584 -67530 -7522 -67430
rect -7522 -67530 -5522 -67430
rect -5522 -67530 -5460 -67430
rect -4004 -67577 -3956 -67562
rect -4004 -67610 -3992 -67577
rect -3992 -67610 -3958 -67577
rect -3958 -67610 -3956 -67577
rect -1460 -67290 -1360 -64666
rect 416 -64526 478 -64426
rect 478 -64526 2478 -64426
rect 2478 -64526 2540 -64426
rect -43 -67299 -9 -67265
rect 49 -67299 83 -67265
rect 141 -67299 175 -67265
rect 316 -67290 416 -64666
rect 767 -65578 851 -65544
rect 1025 -65578 1109 -65544
rect 1283 -65578 1367 -65544
rect 1541 -65578 1625 -65544
rect 1799 -65578 1883 -65544
rect 2057 -65578 2141 -65544
rect 663 -66013 697 -65637
rect 921 -66013 955 -65637
rect 1179 -66013 1213 -65637
rect 1437 -66013 1471 -65637
rect 1695 -66013 1729 -65637
rect 1953 -66013 1987 -65637
rect 2211 -66013 2245 -65637
rect 767 -66106 851 -66072
rect 1025 -66106 1109 -66072
rect 1283 -66106 1367 -66072
rect 1541 -66106 1625 -66072
rect 1799 -66106 1883 -66072
rect 2057 -66106 2141 -66072
rect 767 -66438 851 -66404
rect 1025 -66438 1109 -66404
rect 1283 -66438 1367 -66404
rect 1541 -66438 1625 -66404
rect 1799 -66438 1883 -66404
rect 2057 -66438 2141 -66404
rect 663 -66873 697 -66497
rect 921 -66873 955 -66497
rect 1179 -66873 1213 -66497
rect 1437 -66873 1471 -66497
rect 1695 -66873 1729 -66497
rect 1953 -66873 1987 -66497
rect 2211 -66873 2245 -66497
rect 767 -66966 851 -66932
rect 1025 -66966 1109 -66932
rect 1283 -66966 1367 -66932
rect 1541 -66966 1625 -66932
rect 1799 -66966 1883 -66932
rect 2057 -66966 2141 -66932
rect -3584 -67530 -3522 -67430
rect -3522 -67530 -1522 -67430
rect -1522 -67530 -1460 -67430
rect -4 -67577 44 -67562
rect -4 -67610 8 -67577
rect 8 -67610 42 -67577
rect 42 -67610 44 -67577
rect 2540 -67290 2640 -64666
rect 4416 -64526 4478 -64426
rect 4478 -64526 6478 -64426
rect 6478 -64526 6540 -64426
rect 3957 -67299 3991 -67265
rect 4049 -67299 4083 -67265
rect 4141 -67299 4175 -67265
rect 4316 -67290 4416 -64666
rect 4767 -65578 4851 -65544
rect 5025 -65578 5109 -65544
rect 5283 -65578 5367 -65544
rect 5541 -65578 5625 -65544
rect 5799 -65578 5883 -65544
rect 6057 -65578 6141 -65544
rect 4663 -66013 4697 -65637
rect 4921 -66013 4955 -65637
rect 5179 -66013 5213 -65637
rect 5437 -66013 5471 -65637
rect 5695 -66013 5729 -65637
rect 5953 -66013 5987 -65637
rect 6211 -66013 6245 -65637
rect 4767 -66106 4851 -66072
rect 5025 -66106 5109 -66072
rect 5283 -66106 5367 -66072
rect 5541 -66106 5625 -66072
rect 5799 -66106 5883 -66072
rect 6057 -66106 6141 -66072
rect 4767 -66438 4851 -66404
rect 5025 -66438 5109 -66404
rect 5283 -66438 5367 -66404
rect 5541 -66438 5625 -66404
rect 5799 -66438 5883 -66404
rect 6057 -66438 6141 -66404
rect 4663 -66873 4697 -66497
rect 4921 -66873 4955 -66497
rect 5179 -66873 5213 -66497
rect 5437 -66873 5471 -66497
rect 5695 -66873 5729 -66497
rect 5953 -66873 5987 -66497
rect 6211 -66873 6245 -66497
rect 4767 -66966 4851 -66932
rect 5025 -66966 5109 -66932
rect 5283 -66966 5367 -66932
rect 5541 -66966 5625 -66932
rect 5799 -66966 5883 -66932
rect 6057 -66966 6141 -66932
rect 416 -67530 478 -67430
rect 478 -67530 2478 -67430
rect 2478 -67530 2540 -67430
rect 3996 -67577 4044 -67562
rect 3996 -67610 4008 -67577
rect 4008 -67610 4042 -67577
rect 4042 -67610 4044 -67577
rect 6540 -67290 6640 -64666
rect 4416 -67530 4478 -67430
rect 4478 -67530 6478 -67430
rect 6478 -67530 6540 -67430
rect -27902 -67661 -27854 -67620
rect -27902 -67668 -27878 -67661
rect -27878 -67668 -27854 -67661
rect -28043 -67843 -28009 -67809
rect -27951 -67843 -27917 -67809
rect -27859 -67843 -27825 -67809
rect -27584 -67866 -27522 -67766
rect -27522 -67866 -25522 -67766
rect -25522 -67866 -25460 -67766
rect -27684 -69618 -27584 -67958
rect -23902 -67661 -23854 -67620
rect -23902 -67668 -23878 -67661
rect -23878 -67668 -23854 -67661
rect -24043 -67843 -24009 -67809
rect -23951 -67843 -23917 -67809
rect -23859 -67843 -23825 -67809
rect -27238 -68280 -27154 -68246
rect -26980 -68280 -26896 -68246
rect -26722 -68280 -26638 -68246
rect -26464 -68280 -26380 -68246
rect -26206 -68280 -26122 -68246
rect -25948 -68280 -25864 -68246
rect -27342 -68706 -27308 -68330
rect -27084 -68706 -27050 -68330
rect -26826 -68706 -26792 -68330
rect -26568 -68706 -26534 -68330
rect -26310 -68706 -26276 -68330
rect -26052 -68706 -26018 -68330
rect -25794 -68706 -25760 -68330
rect -27238 -68790 -27154 -68756
rect -26980 -68790 -26896 -68756
rect -26722 -68790 -26638 -68756
rect -26464 -68790 -26380 -68756
rect -26206 -68790 -26122 -68756
rect -25948 -68790 -25864 -68756
rect -25460 -69618 -25360 -67958
rect -27584 -69810 -27522 -69710
rect -27522 -69810 -25522 -69710
rect -25522 -69810 -25460 -69710
rect -23584 -67866 -23522 -67766
rect -23522 -67866 -21522 -67766
rect -21522 -67866 -21460 -67766
rect -23684 -69618 -23584 -67958
rect -19902 -67661 -19854 -67620
rect -19902 -67668 -19878 -67661
rect -19878 -67668 -19854 -67661
rect -20043 -67843 -20009 -67809
rect -19951 -67843 -19917 -67809
rect -19859 -67843 -19825 -67809
rect -23238 -68280 -23154 -68246
rect -22980 -68280 -22896 -68246
rect -22722 -68280 -22638 -68246
rect -22464 -68280 -22380 -68246
rect -22206 -68280 -22122 -68246
rect -21948 -68280 -21864 -68246
rect -23342 -68706 -23308 -68330
rect -23084 -68706 -23050 -68330
rect -22826 -68706 -22792 -68330
rect -22568 -68706 -22534 -68330
rect -22310 -68706 -22276 -68330
rect -22052 -68706 -22018 -68330
rect -21794 -68706 -21760 -68330
rect -23238 -68790 -23154 -68756
rect -22980 -68790 -22896 -68756
rect -22722 -68790 -22638 -68756
rect -22464 -68790 -22380 -68756
rect -22206 -68790 -22122 -68756
rect -21948 -68790 -21864 -68756
rect -21460 -69618 -21360 -67958
rect -23584 -69810 -23522 -69710
rect -23522 -69810 -21522 -69710
rect -21522 -69810 -21460 -69710
rect -19584 -67866 -19522 -67766
rect -19522 -67866 -17522 -67766
rect -17522 -67866 -17460 -67766
rect -19684 -69618 -19584 -67958
rect -15902 -67661 -15854 -67620
rect -15902 -67668 -15878 -67661
rect -15878 -67668 -15854 -67661
rect -16043 -67843 -16009 -67809
rect -15951 -67843 -15917 -67809
rect -15859 -67843 -15825 -67809
rect -19238 -68280 -19154 -68246
rect -18980 -68280 -18896 -68246
rect -18722 -68280 -18638 -68246
rect -18464 -68280 -18380 -68246
rect -18206 -68280 -18122 -68246
rect -17948 -68280 -17864 -68246
rect -19342 -68706 -19308 -68330
rect -19084 -68706 -19050 -68330
rect -18826 -68706 -18792 -68330
rect -18568 -68706 -18534 -68330
rect -18310 -68706 -18276 -68330
rect -18052 -68706 -18018 -68330
rect -17794 -68706 -17760 -68330
rect -19238 -68790 -19154 -68756
rect -18980 -68790 -18896 -68756
rect -18722 -68790 -18638 -68756
rect -18464 -68790 -18380 -68756
rect -18206 -68790 -18122 -68756
rect -17948 -68790 -17864 -68756
rect -17460 -69618 -17360 -67958
rect -19584 -69810 -19522 -69710
rect -19522 -69810 -17522 -69710
rect -17522 -69810 -17460 -69710
rect -15584 -67866 -15522 -67766
rect -15522 -67866 -13522 -67766
rect -13522 -67866 -13460 -67766
rect -15684 -69618 -15584 -67958
rect -11902 -67661 -11854 -67620
rect -11902 -67668 -11878 -67661
rect -11878 -67668 -11854 -67661
rect -12043 -67843 -12009 -67809
rect -11951 -67843 -11917 -67809
rect -11859 -67843 -11825 -67809
rect -15238 -68280 -15154 -68246
rect -14980 -68280 -14896 -68246
rect -14722 -68280 -14638 -68246
rect -14464 -68280 -14380 -68246
rect -14206 -68280 -14122 -68246
rect -13948 -68280 -13864 -68246
rect -15342 -68706 -15308 -68330
rect -15084 -68706 -15050 -68330
rect -14826 -68706 -14792 -68330
rect -14568 -68706 -14534 -68330
rect -14310 -68706 -14276 -68330
rect -14052 -68706 -14018 -68330
rect -13794 -68706 -13760 -68330
rect -15238 -68790 -15154 -68756
rect -14980 -68790 -14896 -68756
rect -14722 -68790 -14638 -68756
rect -14464 -68790 -14380 -68756
rect -14206 -68790 -14122 -68756
rect -13948 -68790 -13864 -68756
rect -13460 -69618 -13360 -67958
rect -15584 -69810 -15522 -69710
rect -15522 -69810 -13522 -69710
rect -13522 -69810 -13460 -69710
rect -11584 -67866 -11522 -67766
rect -11522 -67866 -9522 -67766
rect -9522 -67866 -9460 -67766
rect -11684 -69618 -11584 -67958
rect -7902 -67661 -7854 -67620
rect -7902 -67668 -7878 -67661
rect -7878 -67668 -7854 -67661
rect -8043 -67843 -8009 -67809
rect -7951 -67843 -7917 -67809
rect -7859 -67843 -7825 -67809
rect -11238 -68280 -11154 -68246
rect -10980 -68280 -10896 -68246
rect -10722 -68280 -10638 -68246
rect -10464 -68280 -10380 -68246
rect -10206 -68280 -10122 -68246
rect -9948 -68280 -9864 -68246
rect -11342 -68706 -11308 -68330
rect -11084 -68706 -11050 -68330
rect -10826 -68706 -10792 -68330
rect -10568 -68706 -10534 -68330
rect -10310 -68706 -10276 -68330
rect -10052 -68706 -10018 -68330
rect -9794 -68706 -9760 -68330
rect -11238 -68790 -11154 -68756
rect -10980 -68790 -10896 -68756
rect -10722 -68790 -10638 -68756
rect -10464 -68790 -10380 -68756
rect -10206 -68790 -10122 -68756
rect -9948 -68790 -9864 -68756
rect -9460 -69618 -9360 -67958
rect -11584 -69810 -11522 -69710
rect -11522 -69810 -9522 -69710
rect -9522 -69810 -9460 -69710
rect -7584 -67866 -7522 -67766
rect -7522 -67866 -5522 -67766
rect -5522 -67866 -5460 -67766
rect -7684 -69618 -7584 -67958
rect -3902 -67661 -3854 -67620
rect -3902 -67668 -3878 -67661
rect -3878 -67668 -3854 -67661
rect -4043 -67843 -4009 -67809
rect -3951 -67843 -3917 -67809
rect -3859 -67843 -3825 -67809
rect -7238 -68280 -7154 -68246
rect -6980 -68280 -6896 -68246
rect -6722 -68280 -6638 -68246
rect -6464 -68280 -6380 -68246
rect -6206 -68280 -6122 -68246
rect -5948 -68280 -5864 -68246
rect -7342 -68706 -7308 -68330
rect -7084 -68706 -7050 -68330
rect -6826 -68706 -6792 -68330
rect -6568 -68706 -6534 -68330
rect -6310 -68706 -6276 -68330
rect -6052 -68706 -6018 -68330
rect -5794 -68706 -5760 -68330
rect -7238 -68790 -7154 -68756
rect -6980 -68790 -6896 -68756
rect -6722 -68790 -6638 -68756
rect -6464 -68790 -6380 -68756
rect -6206 -68790 -6122 -68756
rect -5948 -68790 -5864 -68756
rect -5460 -69618 -5360 -67958
rect -7584 -69810 -7522 -69710
rect -7522 -69810 -5522 -69710
rect -5522 -69810 -5460 -69710
rect -3584 -67866 -3522 -67766
rect -3522 -67866 -1522 -67766
rect -1522 -67866 -1460 -67766
rect -3684 -69618 -3584 -67958
rect 98 -67661 146 -67620
rect 98 -67668 122 -67661
rect 122 -67668 146 -67661
rect -43 -67843 -9 -67809
rect 49 -67843 83 -67809
rect 141 -67843 175 -67809
rect -3238 -68280 -3154 -68246
rect -2980 -68280 -2896 -68246
rect -2722 -68280 -2638 -68246
rect -2464 -68280 -2380 -68246
rect -2206 -68280 -2122 -68246
rect -1948 -68280 -1864 -68246
rect -3342 -68706 -3308 -68330
rect -3084 -68706 -3050 -68330
rect -2826 -68706 -2792 -68330
rect -2568 -68706 -2534 -68330
rect -2310 -68706 -2276 -68330
rect -2052 -68706 -2018 -68330
rect -1794 -68706 -1760 -68330
rect -3238 -68790 -3154 -68756
rect -2980 -68790 -2896 -68756
rect -2722 -68790 -2638 -68756
rect -2464 -68790 -2380 -68756
rect -2206 -68790 -2122 -68756
rect -1948 -68790 -1864 -68756
rect -1460 -69618 -1360 -67958
rect -3584 -69810 -3522 -69710
rect -3522 -69810 -1522 -69710
rect -1522 -69810 -1460 -69710
rect 416 -67866 478 -67766
rect 478 -67866 2478 -67766
rect 2478 -67866 2540 -67766
rect 316 -69618 416 -67958
rect 4098 -67661 4146 -67620
rect 4098 -67668 4122 -67661
rect 4122 -67668 4146 -67661
rect 3957 -67843 3991 -67809
rect 4049 -67843 4083 -67809
rect 4141 -67843 4175 -67809
rect 762 -68280 846 -68246
rect 1020 -68280 1104 -68246
rect 1278 -68280 1362 -68246
rect 1536 -68280 1620 -68246
rect 1794 -68280 1878 -68246
rect 2052 -68280 2136 -68246
rect 658 -68706 692 -68330
rect 916 -68706 950 -68330
rect 1174 -68706 1208 -68330
rect 1432 -68706 1466 -68330
rect 1690 -68706 1724 -68330
rect 1948 -68706 1982 -68330
rect 2206 -68706 2240 -68330
rect 762 -68790 846 -68756
rect 1020 -68790 1104 -68756
rect 1278 -68790 1362 -68756
rect 1536 -68790 1620 -68756
rect 1794 -68790 1878 -68756
rect 2052 -68790 2136 -68756
rect 2540 -69618 2640 -67958
rect 416 -69810 478 -69710
rect 478 -69810 2478 -69710
rect 2478 -69810 2540 -69710
rect 4416 -67866 4478 -67766
rect 4478 -67866 6478 -67766
rect 6478 -67866 6540 -67766
rect 4316 -69618 4416 -67958
rect 4762 -68280 4846 -68246
rect 5020 -68280 5104 -68246
rect 5278 -68280 5362 -68246
rect 5536 -68280 5620 -68246
rect 5794 -68280 5878 -68246
rect 6052 -68280 6136 -68246
rect 4658 -68706 4692 -68330
rect 4916 -68706 4950 -68330
rect 5174 -68706 5208 -68330
rect 5432 -68706 5466 -68330
rect 5690 -68706 5724 -68330
rect 5948 -68706 5982 -68330
rect 6206 -68706 6240 -68330
rect 4762 -68790 4846 -68756
rect 5020 -68790 5104 -68756
rect 5278 -68790 5362 -68756
rect 5536 -68790 5620 -68756
rect 5794 -68790 5878 -68756
rect 6052 -68790 6136 -68756
rect 6540 -69618 6640 -67958
rect 4416 -69810 4478 -69710
rect 4478 -69810 6478 -69710
rect 6478 -69810 6540 -69710
rect -27584 -70486 -27522 -70386
rect -27522 -70486 -25522 -70386
rect -25522 -70486 -25460 -70386
rect -27684 -72238 -27584 -70578
rect -27238 -71440 -27154 -71406
rect -26980 -71440 -26896 -71406
rect -26722 -71440 -26638 -71406
rect -26464 -71440 -26380 -71406
rect -26206 -71440 -26122 -71406
rect -25948 -71440 -25864 -71406
rect -27342 -71866 -27308 -71490
rect -27084 -71866 -27050 -71490
rect -26826 -71866 -26792 -71490
rect -26568 -71866 -26534 -71490
rect -26310 -71866 -26276 -71490
rect -26052 -71866 -26018 -71490
rect -25794 -71866 -25760 -71490
rect -27238 -71950 -27154 -71916
rect -26980 -71950 -26896 -71916
rect -26722 -71950 -26638 -71916
rect -26464 -71950 -26380 -71916
rect -26206 -71950 -26122 -71916
rect -25948 -71950 -25864 -71916
rect -28043 -72387 -28009 -72353
rect -27951 -72387 -27917 -72353
rect -27859 -72387 -27825 -72353
rect -25460 -72238 -25360 -70578
rect -27584 -72430 -27522 -72330
rect -27522 -72430 -25522 -72330
rect -25522 -72430 -25460 -72330
rect -23584 -70486 -23522 -70386
rect -23522 -70486 -21522 -70386
rect -21522 -70486 -21460 -70386
rect -23684 -72238 -23584 -70578
rect -23238 -71440 -23154 -71406
rect -22980 -71440 -22896 -71406
rect -22722 -71440 -22638 -71406
rect -22464 -71440 -22380 -71406
rect -22206 -71440 -22122 -71406
rect -21948 -71440 -21864 -71406
rect -23342 -71866 -23308 -71490
rect -23084 -71866 -23050 -71490
rect -22826 -71866 -22792 -71490
rect -22568 -71866 -22534 -71490
rect -22310 -71866 -22276 -71490
rect -22052 -71866 -22018 -71490
rect -21794 -71866 -21760 -71490
rect -23238 -71950 -23154 -71916
rect -22980 -71950 -22896 -71916
rect -22722 -71950 -22638 -71916
rect -22464 -71950 -22380 -71916
rect -22206 -71950 -22122 -71916
rect -21948 -71950 -21864 -71916
rect -24043 -72387 -24009 -72353
rect -23951 -72387 -23917 -72353
rect -23859 -72387 -23825 -72353
rect -27902 -72535 -27878 -72528
rect -27878 -72535 -27854 -72528
rect -27902 -72576 -27854 -72535
rect -21460 -72238 -21360 -70578
rect -23584 -72430 -23522 -72330
rect -23522 -72430 -21522 -72330
rect -21522 -72430 -21460 -72330
rect -19584 -70486 -19522 -70386
rect -19522 -70486 -17522 -70386
rect -17522 -70486 -17460 -70386
rect -19684 -72238 -19584 -70578
rect -19238 -71440 -19154 -71406
rect -18980 -71440 -18896 -71406
rect -18722 -71440 -18638 -71406
rect -18464 -71440 -18380 -71406
rect -18206 -71440 -18122 -71406
rect -17948 -71440 -17864 -71406
rect -19342 -71866 -19308 -71490
rect -19084 -71866 -19050 -71490
rect -18826 -71866 -18792 -71490
rect -18568 -71866 -18534 -71490
rect -18310 -71866 -18276 -71490
rect -18052 -71866 -18018 -71490
rect -17794 -71866 -17760 -71490
rect -19238 -71950 -19154 -71916
rect -18980 -71950 -18896 -71916
rect -18722 -71950 -18638 -71916
rect -18464 -71950 -18380 -71916
rect -18206 -71950 -18122 -71916
rect -17948 -71950 -17864 -71916
rect -20043 -72387 -20009 -72353
rect -19951 -72387 -19917 -72353
rect -19859 -72387 -19825 -72353
rect -23902 -72535 -23878 -72528
rect -23878 -72535 -23854 -72528
rect -23902 -72576 -23854 -72535
rect -17460 -72238 -17360 -70578
rect -19584 -72430 -19522 -72330
rect -19522 -72430 -17522 -72330
rect -17522 -72430 -17460 -72330
rect -15584 -70486 -15522 -70386
rect -15522 -70486 -13522 -70386
rect -13522 -70486 -13460 -70386
rect -15684 -72238 -15584 -70578
rect -15238 -71440 -15154 -71406
rect -14980 -71440 -14896 -71406
rect -14722 -71440 -14638 -71406
rect -14464 -71440 -14380 -71406
rect -14206 -71440 -14122 -71406
rect -13948 -71440 -13864 -71406
rect -15342 -71866 -15308 -71490
rect -15084 -71866 -15050 -71490
rect -14826 -71866 -14792 -71490
rect -14568 -71866 -14534 -71490
rect -14310 -71866 -14276 -71490
rect -14052 -71866 -14018 -71490
rect -13794 -71866 -13760 -71490
rect -15238 -71950 -15154 -71916
rect -14980 -71950 -14896 -71916
rect -14722 -71950 -14638 -71916
rect -14464 -71950 -14380 -71916
rect -14206 -71950 -14122 -71916
rect -13948 -71950 -13864 -71916
rect -16043 -72387 -16009 -72353
rect -15951 -72387 -15917 -72353
rect -15859 -72387 -15825 -72353
rect -19902 -72535 -19878 -72528
rect -19878 -72535 -19854 -72528
rect -19902 -72576 -19854 -72535
rect -13460 -72238 -13360 -70578
rect -15584 -72430 -15522 -72330
rect -15522 -72430 -13522 -72330
rect -13522 -72430 -13460 -72330
rect -11584 -70486 -11522 -70386
rect -11522 -70486 -9522 -70386
rect -9522 -70486 -9460 -70386
rect -11684 -72238 -11584 -70578
rect -11238 -71440 -11154 -71406
rect -10980 -71440 -10896 -71406
rect -10722 -71440 -10638 -71406
rect -10464 -71440 -10380 -71406
rect -10206 -71440 -10122 -71406
rect -9948 -71440 -9864 -71406
rect -11342 -71866 -11308 -71490
rect -11084 -71866 -11050 -71490
rect -10826 -71866 -10792 -71490
rect -10568 -71866 -10534 -71490
rect -10310 -71866 -10276 -71490
rect -10052 -71866 -10018 -71490
rect -9794 -71866 -9760 -71490
rect -11238 -71950 -11154 -71916
rect -10980 -71950 -10896 -71916
rect -10722 -71950 -10638 -71916
rect -10464 -71950 -10380 -71916
rect -10206 -71950 -10122 -71916
rect -9948 -71950 -9864 -71916
rect -12043 -72387 -12009 -72353
rect -11951 -72387 -11917 -72353
rect -11859 -72387 -11825 -72353
rect -15902 -72535 -15878 -72528
rect -15878 -72535 -15854 -72528
rect -15902 -72576 -15854 -72535
rect -9460 -72238 -9360 -70578
rect -11584 -72430 -11522 -72330
rect -11522 -72430 -9522 -72330
rect -9522 -72430 -9460 -72330
rect -7584 -70486 -7522 -70386
rect -7522 -70486 -5522 -70386
rect -5522 -70486 -5460 -70386
rect -7684 -72238 -7584 -70578
rect -7238 -71440 -7154 -71406
rect -6980 -71440 -6896 -71406
rect -6722 -71440 -6638 -71406
rect -6464 -71440 -6380 -71406
rect -6206 -71440 -6122 -71406
rect -5948 -71440 -5864 -71406
rect -7342 -71866 -7308 -71490
rect -7084 -71866 -7050 -71490
rect -6826 -71866 -6792 -71490
rect -6568 -71866 -6534 -71490
rect -6310 -71866 -6276 -71490
rect -6052 -71866 -6018 -71490
rect -5794 -71866 -5760 -71490
rect -7238 -71950 -7154 -71916
rect -6980 -71950 -6896 -71916
rect -6722 -71950 -6638 -71916
rect -6464 -71950 -6380 -71916
rect -6206 -71950 -6122 -71916
rect -5948 -71950 -5864 -71916
rect -8043 -72387 -8009 -72353
rect -7951 -72387 -7917 -72353
rect -7859 -72387 -7825 -72353
rect -11902 -72535 -11878 -72528
rect -11878 -72535 -11854 -72528
rect -11902 -72576 -11854 -72535
rect -5460 -72238 -5360 -70578
rect -7584 -72430 -7522 -72330
rect -7522 -72430 -5522 -72330
rect -5522 -72430 -5460 -72330
rect -3584 -70486 -3522 -70386
rect -3522 -70486 -1522 -70386
rect -1522 -70486 -1460 -70386
rect -3684 -72238 -3584 -70578
rect -3238 -71440 -3154 -71406
rect -2980 -71440 -2896 -71406
rect -2722 -71440 -2638 -71406
rect -2464 -71440 -2380 -71406
rect -2206 -71440 -2122 -71406
rect -1948 -71440 -1864 -71406
rect -3342 -71866 -3308 -71490
rect -3084 -71866 -3050 -71490
rect -2826 -71866 -2792 -71490
rect -2568 -71866 -2534 -71490
rect -2310 -71866 -2276 -71490
rect -2052 -71866 -2018 -71490
rect -1794 -71866 -1760 -71490
rect -3238 -71950 -3154 -71916
rect -2980 -71950 -2896 -71916
rect -2722 -71950 -2638 -71916
rect -2464 -71950 -2380 -71916
rect -2206 -71950 -2122 -71916
rect -1948 -71950 -1864 -71916
rect -4043 -72387 -4009 -72353
rect -3951 -72387 -3917 -72353
rect -3859 -72387 -3825 -72353
rect -7902 -72535 -7878 -72528
rect -7878 -72535 -7854 -72528
rect -7902 -72576 -7854 -72535
rect -1460 -72238 -1360 -70578
rect -3584 -72430 -3522 -72330
rect -3522 -72430 -1522 -72330
rect -1522 -72430 -1460 -72330
rect 416 -70486 478 -70386
rect 478 -70486 2478 -70386
rect 2478 -70486 2540 -70386
rect 316 -72238 416 -70578
rect 762 -71440 846 -71406
rect 1020 -71440 1104 -71406
rect 1278 -71440 1362 -71406
rect 1536 -71440 1620 -71406
rect 1794 -71440 1878 -71406
rect 2052 -71440 2136 -71406
rect 658 -71866 692 -71490
rect 916 -71866 950 -71490
rect 1174 -71866 1208 -71490
rect 1432 -71866 1466 -71490
rect 1690 -71866 1724 -71490
rect 1948 -71866 1982 -71490
rect 2206 -71866 2240 -71490
rect 762 -71950 846 -71916
rect 1020 -71950 1104 -71916
rect 1278 -71950 1362 -71916
rect 1536 -71950 1620 -71916
rect 1794 -71950 1878 -71916
rect 2052 -71950 2136 -71916
rect -43 -72387 -9 -72353
rect 49 -72387 83 -72353
rect 141 -72387 175 -72353
rect -3902 -72535 -3878 -72528
rect -3878 -72535 -3854 -72528
rect -3902 -72576 -3854 -72535
rect 2540 -72238 2640 -70578
rect 416 -72430 478 -72330
rect 478 -72430 2478 -72330
rect 2478 -72430 2540 -72330
rect 4416 -70486 4478 -70386
rect 4478 -70486 6478 -70386
rect 6478 -70486 6540 -70386
rect 4316 -72238 4416 -70578
rect 4762 -71440 4846 -71406
rect 5020 -71440 5104 -71406
rect 5278 -71440 5362 -71406
rect 5536 -71440 5620 -71406
rect 5794 -71440 5878 -71406
rect 6052 -71440 6136 -71406
rect 4658 -71866 4692 -71490
rect 4916 -71866 4950 -71490
rect 5174 -71866 5208 -71490
rect 5432 -71866 5466 -71490
rect 5690 -71866 5724 -71490
rect 5948 -71866 5982 -71490
rect 6206 -71866 6240 -71490
rect 4762 -71950 4846 -71916
rect 5020 -71950 5104 -71916
rect 5278 -71950 5362 -71916
rect 5536 -71950 5620 -71916
rect 5794 -71950 5878 -71916
rect 6052 -71950 6136 -71916
rect 3957 -72387 3991 -72353
rect 4049 -72387 4083 -72353
rect 4141 -72387 4175 -72353
rect 98 -72535 122 -72528
rect 122 -72535 146 -72528
rect 98 -72576 146 -72535
rect 6540 -72238 6640 -70578
rect 4416 -72430 4478 -72330
rect 4478 -72430 6478 -72330
rect 6478 -72430 6540 -72330
rect 4098 -72535 4122 -72528
rect 4122 -72535 4146 -72528
rect 4098 -72576 4146 -72535
rect -28004 -72619 -27992 -72586
rect -27992 -72619 -27958 -72586
rect -27958 -72619 -27956 -72586
rect -28004 -72634 -27956 -72619
rect -24004 -72619 -23992 -72586
rect -23992 -72619 -23958 -72586
rect -23958 -72619 -23956 -72586
rect -24004 -72634 -23956 -72619
rect -27584 -72766 -27522 -72666
rect -27522 -72766 -25522 -72666
rect -25522 -72766 -25460 -72666
rect -28043 -72931 -28009 -72897
rect -27951 -72931 -27917 -72897
rect -27859 -72931 -27825 -72897
rect -27684 -75530 -27584 -72906
rect -20004 -72619 -19992 -72586
rect -19992 -72619 -19958 -72586
rect -19958 -72619 -19956 -72586
rect -20004 -72634 -19956 -72619
rect -23584 -72766 -23522 -72666
rect -23522 -72766 -21522 -72666
rect -21522 -72766 -21460 -72666
rect -27233 -73264 -27149 -73230
rect -26975 -73264 -26891 -73230
rect -26717 -73264 -26633 -73230
rect -26459 -73264 -26375 -73230
rect -26201 -73264 -26117 -73230
rect -25943 -73264 -25859 -73230
rect -27337 -73699 -27303 -73323
rect -27079 -73699 -27045 -73323
rect -26821 -73699 -26787 -73323
rect -26563 -73699 -26529 -73323
rect -26305 -73699 -26271 -73323
rect -26047 -73699 -26013 -73323
rect -25789 -73699 -25755 -73323
rect -27233 -73792 -27149 -73758
rect -26975 -73792 -26891 -73758
rect -26717 -73792 -26633 -73758
rect -26459 -73792 -26375 -73758
rect -26201 -73792 -26117 -73758
rect -25943 -73792 -25859 -73758
rect -27233 -74124 -27149 -74090
rect -26975 -74124 -26891 -74090
rect -26717 -74124 -26633 -74090
rect -26459 -74124 -26375 -74090
rect -26201 -74124 -26117 -74090
rect -25943 -74124 -25859 -74090
rect -27337 -74559 -27303 -74183
rect -27079 -74559 -27045 -74183
rect -26821 -74559 -26787 -74183
rect -26563 -74559 -26529 -74183
rect -26305 -74559 -26271 -74183
rect -26047 -74559 -26013 -74183
rect -25789 -74559 -25755 -74183
rect -27233 -74652 -27149 -74618
rect -26975 -74652 -26891 -74618
rect -26717 -74652 -26633 -74618
rect -26459 -74652 -26375 -74618
rect -26201 -74652 -26117 -74618
rect -25943 -74652 -25859 -74618
rect -25460 -75530 -25360 -72906
rect -24043 -72931 -24009 -72897
rect -23951 -72931 -23917 -72897
rect -23859 -72931 -23825 -72897
rect -27584 -75770 -27522 -75670
rect -27522 -75770 -25522 -75670
rect -25522 -75770 -25460 -75670
rect -23684 -75530 -23584 -72906
rect -16004 -72619 -15992 -72586
rect -15992 -72619 -15958 -72586
rect -15958 -72619 -15956 -72586
rect -16004 -72634 -15956 -72619
rect -19584 -72766 -19522 -72666
rect -19522 -72766 -17522 -72666
rect -17522 -72766 -17460 -72666
rect -23233 -73264 -23149 -73230
rect -22975 -73264 -22891 -73230
rect -22717 -73264 -22633 -73230
rect -22459 -73264 -22375 -73230
rect -22201 -73264 -22117 -73230
rect -21943 -73264 -21859 -73230
rect -23337 -73699 -23303 -73323
rect -23079 -73699 -23045 -73323
rect -22821 -73699 -22787 -73323
rect -22563 -73699 -22529 -73323
rect -22305 -73699 -22271 -73323
rect -22047 -73699 -22013 -73323
rect -21789 -73699 -21755 -73323
rect -23233 -73792 -23149 -73758
rect -22975 -73792 -22891 -73758
rect -22717 -73792 -22633 -73758
rect -22459 -73792 -22375 -73758
rect -22201 -73792 -22117 -73758
rect -21943 -73792 -21859 -73758
rect -23233 -74124 -23149 -74090
rect -22975 -74124 -22891 -74090
rect -22717 -74124 -22633 -74090
rect -22459 -74124 -22375 -74090
rect -22201 -74124 -22117 -74090
rect -21943 -74124 -21859 -74090
rect -23337 -74559 -23303 -74183
rect -23079 -74559 -23045 -74183
rect -22821 -74559 -22787 -74183
rect -22563 -74559 -22529 -74183
rect -22305 -74559 -22271 -74183
rect -22047 -74559 -22013 -74183
rect -21789 -74559 -21755 -74183
rect -23233 -74652 -23149 -74618
rect -22975 -74652 -22891 -74618
rect -22717 -74652 -22633 -74618
rect -22459 -74652 -22375 -74618
rect -22201 -74652 -22117 -74618
rect -21943 -74652 -21859 -74618
rect -21460 -75530 -21360 -72906
rect -20043 -72931 -20009 -72897
rect -19951 -72931 -19917 -72897
rect -19859 -72931 -19825 -72897
rect -23584 -75770 -23522 -75670
rect -23522 -75770 -21522 -75670
rect -21522 -75770 -21460 -75670
rect -19684 -75530 -19584 -72906
rect -12004 -72619 -11992 -72586
rect -11992 -72619 -11958 -72586
rect -11958 -72619 -11956 -72586
rect -12004 -72634 -11956 -72619
rect -15584 -72766 -15522 -72666
rect -15522 -72766 -13522 -72666
rect -13522 -72766 -13460 -72666
rect -19233 -73264 -19149 -73230
rect -18975 -73264 -18891 -73230
rect -18717 -73264 -18633 -73230
rect -18459 -73264 -18375 -73230
rect -18201 -73264 -18117 -73230
rect -17943 -73264 -17859 -73230
rect -19337 -73699 -19303 -73323
rect -19079 -73699 -19045 -73323
rect -18821 -73699 -18787 -73323
rect -18563 -73699 -18529 -73323
rect -18305 -73699 -18271 -73323
rect -18047 -73699 -18013 -73323
rect -17789 -73699 -17755 -73323
rect -19233 -73792 -19149 -73758
rect -18975 -73792 -18891 -73758
rect -18717 -73792 -18633 -73758
rect -18459 -73792 -18375 -73758
rect -18201 -73792 -18117 -73758
rect -17943 -73792 -17859 -73758
rect -19233 -74124 -19149 -74090
rect -18975 -74124 -18891 -74090
rect -18717 -74124 -18633 -74090
rect -18459 -74124 -18375 -74090
rect -18201 -74124 -18117 -74090
rect -17943 -74124 -17859 -74090
rect -19337 -74559 -19303 -74183
rect -19079 -74559 -19045 -74183
rect -18821 -74559 -18787 -74183
rect -18563 -74559 -18529 -74183
rect -18305 -74559 -18271 -74183
rect -18047 -74559 -18013 -74183
rect -17789 -74559 -17755 -74183
rect -19233 -74652 -19149 -74618
rect -18975 -74652 -18891 -74618
rect -18717 -74652 -18633 -74618
rect -18459 -74652 -18375 -74618
rect -18201 -74652 -18117 -74618
rect -17943 -74652 -17859 -74618
rect -17460 -75530 -17360 -72906
rect -16043 -72931 -16009 -72897
rect -15951 -72931 -15917 -72897
rect -15859 -72931 -15825 -72897
rect -19584 -75770 -19522 -75670
rect -19522 -75770 -17522 -75670
rect -17522 -75770 -17460 -75670
rect -15684 -75530 -15584 -72906
rect -8004 -72619 -7992 -72586
rect -7992 -72619 -7958 -72586
rect -7958 -72619 -7956 -72586
rect -8004 -72634 -7956 -72619
rect -11584 -72766 -11522 -72666
rect -11522 -72766 -9522 -72666
rect -9522 -72766 -9460 -72666
rect -15233 -73264 -15149 -73230
rect -14975 -73264 -14891 -73230
rect -14717 -73264 -14633 -73230
rect -14459 -73264 -14375 -73230
rect -14201 -73264 -14117 -73230
rect -13943 -73264 -13859 -73230
rect -15337 -73699 -15303 -73323
rect -15079 -73699 -15045 -73323
rect -14821 -73699 -14787 -73323
rect -14563 -73699 -14529 -73323
rect -14305 -73699 -14271 -73323
rect -14047 -73699 -14013 -73323
rect -13789 -73699 -13755 -73323
rect -15233 -73792 -15149 -73758
rect -14975 -73792 -14891 -73758
rect -14717 -73792 -14633 -73758
rect -14459 -73792 -14375 -73758
rect -14201 -73792 -14117 -73758
rect -13943 -73792 -13859 -73758
rect -15233 -74124 -15149 -74090
rect -14975 -74124 -14891 -74090
rect -14717 -74124 -14633 -74090
rect -14459 -74124 -14375 -74090
rect -14201 -74124 -14117 -74090
rect -13943 -74124 -13859 -74090
rect -15337 -74559 -15303 -74183
rect -15079 -74559 -15045 -74183
rect -14821 -74559 -14787 -74183
rect -14563 -74559 -14529 -74183
rect -14305 -74559 -14271 -74183
rect -14047 -74559 -14013 -74183
rect -13789 -74559 -13755 -74183
rect -15233 -74652 -15149 -74618
rect -14975 -74652 -14891 -74618
rect -14717 -74652 -14633 -74618
rect -14459 -74652 -14375 -74618
rect -14201 -74652 -14117 -74618
rect -13943 -74652 -13859 -74618
rect -13460 -75530 -13360 -72906
rect -12043 -72931 -12009 -72897
rect -11951 -72931 -11917 -72897
rect -11859 -72931 -11825 -72897
rect -15584 -75770 -15522 -75670
rect -15522 -75770 -13522 -75670
rect -13522 -75770 -13460 -75670
rect -11684 -75530 -11584 -72906
rect -4004 -72619 -3992 -72586
rect -3992 -72619 -3958 -72586
rect -3958 -72619 -3956 -72586
rect -4004 -72634 -3956 -72619
rect -7584 -72766 -7522 -72666
rect -7522 -72766 -5522 -72666
rect -5522 -72766 -5460 -72666
rect -11233 -73264 -11149 -73230
rect -10975 -73264 -10891 -73230
rect -10717 -73264 -10633 -73230
rect -10459 -73264 -10375 -73230
rect -10201 -73264 -10117 -73230
rect -9943 -73264 -9859 -73230
rect -11337 -73699 -11303 -73323
rect -11079 -73699 -11045 -73323
rect -10821 -73699 -10787 -73323
rect -10563 -73699 -10529 -73323
rect -10305 -73699 -10271 -73323
rect -10047 -73699 -10013 -73323
rect -9789 -73699 -9755 -73323
rect -11233 -73792 -11149 -73758
rect -10975 -73792 -10891 -73758
rect -10717 -73792 -10633 -73758
rect -10459 -73792 -10375 -73758
rect -10201 -73792 -10117 -73758
rect -9943 -73792 -9859 -73758
rect -11233 -74124 -11149 -74090
rect -10975 -74124 -10891 -74090
rect -10717 -74124 -10633 -74090
rect -10459 -74124 -10375 -74090
rect -10201 -74124 -10117 -74090
rect -9943 -74124 -9859 -74090
rect -11337 -74559 -11303 -74183
rect -11079 -74559 -11045 -74183
rect -10821 -74559 -10787 -74183
rect -10563 -74559 -10529 -74183
rect -10305 -74559 -10271 -74183
rect -10047 -74559 -10013 -74183
rect -9789 -74559 -9755 -74183
rect -11233 -74652 -11149 -74618
rect -10975 -74652 -10891 -74618
rect -10717 -74652 -10633 -74618
rect -10459 -74652 -10375 -74618
rect -10201 -74652 -10117 -74618
rect -9943 -74652 -9859 -74618
rect -9460 -75530 -9360 -72906
rect -8043 -72931 -8009 -72897
rect -7951 -72931 -7917 -72897
rect -7859 -72931 -7825 -72897
rect -11584 -75770 -11522 -75670
rect -11522 -75770 -9522 -75670
rect -9522 -75770 -9460 -75670
rect -7684 -75530 -7584 -72906
rect -4 -72619 8 -72586
rect 8 -72619 42 -72586
rect 42 -72619 44 -72586
rect -4 -72634 44 -72619
rect -3584 -72766 -3522 -72666
rect -3522 -72766 -1522 -72666
rect -1522 -72766 -1460 -72666
rect -7233 -73264 -7149 -73230
rect -6975 -73264 -6891 -73230
rect -6717 -73264 -6633 -73230
rect -6459 -73264 -6375 -73230
rect -6201 -73264 -6117 -73230
rect -5943 -73264 -5859 -73230
rect -7337 -73699 -7303 -73323
rect -7079 -73699 -7045 -73323
rect -6821 -73699 -6787 -73323
rect -6563 -73699 -6529 -73323
rect -6305 -73699 -6271 -73323
rect -6047 -73699 -6013 -73323
rect -5789 -73699 -5755 -73323
rect -7233 -73792 -7149 -73758
rect -6975 -73792 -6891 -73758
rect -6717 -73792 -6633 -73758
rect -6459 -73792 -6375 -73758
rect -6201 -73792 -6117 -73758
rect -5943 -73792 -5859 -73758
rect -7233 -74124 -7149 -74090
rect -6975 -74124 -6891 -74090
rect -6717 -74124 -6633 -74090
rect -6459 -74124 -6375 -74090
rect -6201 -74124 -6117 -74090
rect -5943 -74124 -5859 -74090
rect -7337 -74559 -7303 -74183
rect -7079 -74559 -7045 -74183
rect -6821 -74559 -6787 -74183
rect -6563 -74559 -6529 -74183
rect -6305 -74559 -6271 -74183
rect -6047 -74559 -6013 -74183
rect -5789 -74559 -5755 -74183
rect -7233 -74652 -7149 -74618
rect -6975 -74652 -6891 -74618
rect -6717 -74652 -6633 -74618
rect -6459 -74652 -6375 -74618
rect -6201 -74652 -6117 -74618
rect -5943 -74652 -5859 -74618
rect -5460 -75530 -5360 -72906
rect -4043 -72931 -4009 -72897
rect -3951 -72931 -3917 -72897
rect -3859 -72931 -3825 -72897
rect -7584 -75770 -7522 -75670
rect -7522 -75770 -5522 -75670
rect -5522 -75770 -5460 -75670
rect -3684 -75530 -3584 -72906
rect 3996 -72619 4008 -72586
rect 4008 -72619 4042 -72586
rect 4042 -72619 4044 -72586
rect 3996 -72634 4044 -72619
rect 416 -72766 478 -72666
rect 478 -72766 2478 -72666
rect 2478 -72766 2540 -72666
rect -3233 -73264 -3149 -73230
rect -2975 -73264 -2891 -73230
rect -2717 -73264 -2633 -73230
rect -2459 -73264 -2375 -73230
rect -2201 -73264 -2117 -73230
rect -1943 -73264 -1859 -73230
rect -3337 -73699 -3303 -73323
rect -3079 -73699 -3045 -73323
rect -2821 -73699 -2787 -73323
rect -2563 -73699 -2529 -73323
rect -2305 -73699 -2271 -73323
rect -2047 -73699 -2013 -73323
rect -1789 -73699 -1755 -73323
rect -3233 -73792 -3149 -73758
rect -2975 -73792 -2891 -73758
rect -2717 -73792 -2633 -73758
rect -2459 -73792 -2375 -73758
rect -2201 -73792 -2117 -73758
rect -1943 -73792 -1859 -73758
rect -3233 -74124 -3149 -74090
rect -2975 -74124 -2891 -74090
rect -2717 -74124 -2633 -74090
rect -2459 -74124 -2375 -74090
rect -2201 -74124 -2117 -74090
rect -1943 -74124 -1859 -74090
rect -3337 -74559 -3303 -74183
rect -3079 -74559 -3045 -74183
rect -2821 -74559 -2787 -74183
rect -2563 -74559 -2529 -74183
rect -2305 -74559 -2271 -74183
rect -2047 -74559 -2013 -74183
rect -1789 -74559 -1755 -74183
rect -3233 -74652 -3149 -74618
rect -2975 -74652 -2891 -74618
rect -2717 -74652 -2633 -74618
rect -2459 -74652 -2375 -74618
rect -2201 -74652 -2117 -74618
rect -1943 -74652 -1859 -74618
rect -1460 -75530 -1360 -72906
rect -43 -72931 -9 -72897
rect 49 -72931 83 -72897
rect 141 -72931 175 -72897
rect -3584 -75770 -3522 -75670
rect -3522 -75770 -1522 -75670
rect -1522 -75770 -1460 -75670
rect 316 -75530 416 -72906
rect 4416 -72766 4478 -72666
rect 4478 -72766 6478 -72666
rect 6478 -72766 6540 -72666
rect 767 -73264 851 -73230
rect 1025 -73264 1109 -73230
rect 1283 -73264 1367 -73230
rect 1541 -73264 1625 -73230
rect 1799 -73264 1883 -73230
rect 2057 -73264 2141 -73230
rect 663 -73699 697 -73323
rect 921 -73699 955 -73323
rect 1179 -73699 1213 -73323
rect 1437 -73699 1471 -73323
rect 1695 -73699 1729 -73323
rect 1953 -73699 1987 -73323
rect 2211 -73699 2245 -73323
rect 767 -73792 851 -73758
rect 1025 -73792 1109 -73758
rect 1283 -73792 1367 -73758
rect 1541 -73792 1625 -73758
rect 1799 -73792 1883 -73758
rect 2057 -73792 2141 -73758
rect 767 -74124 851 -74090
rect 1025 -74124 1109 -74090
rect 1283 -74124 1367 -74090
rect 1541 -74124 1625 -74090
rect 1799 -74124 1883 -74090
rect 2057 -74124 2141 -74090
rect 663 -74559 697 -74183
rect 921 -74559 955 -74183
rect 1179 -74559 1213 -74183
rect 1437 -74559 1471 -74183
rect 1695 -74559 1729 -74183
rect 1953 -74559 1987 -74183
rect 2211 -74559 2245 -74183
rect 767 -74652 851 -74618
rect 1025 -74652 1109 -74618
rect 1283 -74652 1367 -74618
rect 1541 -74652 1625 -74618
rect 1799 -74652 1883 -74618
rect 2057 -74652 2141 -74618
rect 2540 -75530 2640 -72906
rect 3957 -72931 3991 -72897
rect 4049 -72931 4083 -72897
rect 4141 -72931 4175 -72897
rect 416 -75770 478 -75670
rect 478 -75770 2478 -75670
rect 2478 -75770 2540 -75670
rect 4316 -75530 4416 -72906
rect 4767 -73264 4851 -73230
rect 5025 -73264 5109 -73230
rect 5283 -73264 5367 -73230
rect 5541 -73264 5625 -73230
rect 5799 -73264 5883 -73230
rect 6057 -73264 6141 -73230
rect 4663 -73699 4697 -73323
rect 4921 -73699 4955 -73323
rect 5179 -73699 5213 -73323
rect 5437 -73699 5471 -73323
rect 5695 -73699 5729 -73323
rect 5953 -73699 5987 -73323
rect 6211 -73699 6245 -73323
rect 4767 -73792 4851 -73758
rect 5025 -73792 5109 -73758
rect 5283 -73792 5367 -73758
rect 5541 -73792 5625 -73758
rect 5799 -73792 5883 -73758
rect 6057 -73792 6141 -73758
rect 4767 -74124 4851 -74090
rect 5025 -74124 5109 -74090
rect 5283 -74124 5367 -74090
rect 5541 -74124 5625 -74090
rect 5799 -74124 5883 -74090
rect 6057 -74124 6141 -74090
rect 4663 -74559 4697 -74183
rect 4921 -74559 4955 -74183
rect 5179 -74559 5213 -74183
rect 5437 -74559 5471 -74183
rect 5695 -74559 5729 -74183
rect 5953 -74559 5987 -74183
rect 6211 -74559 6245 -74183
rect 4767 -74652 4851 -74618
rect 5025 -74652 5109 -74618
rect 5283 -74652 5367 -74618
rect 5541 -74652 5625 -74618
rect 5799 -74652 5883 -74618
rect 6057 -74652 6141 -74618
rect 6540 -75530 6640 -72906
rect 4416 -75770 4478 -75670
rect 4478 -75770 6478 -75670
rect 6478 -75770 6540 -75670
<< metal1 >>
rect -74 -48 106 12
rect 25816 -27656 50272 -27650
rect 25816 -27756 25922 -27656
rect 50166 -27756 50272 -27656
rect 25816 -27762 50272 -27756
rect 25816 -28276 25928 -27762
rect 26528 -28062 26538 -27762
rect 49550 -28062 49560 -27762
rect 25816 -41706 25822 -28276
rect 25922 -41706 25928 -28276
rect 29442 -28144 46322 -28112
rect 29442 -28358 29505 -28144
rect 46290 -28358 46322 -28144
rect 29442 -28380 29492 -28358
rect 29552 -28380 29928 -28358
rect 29988 -28380 30366 -28358
rect 30426 -28380 30800 -28358
rect 30860 -28378 46322 -28358
rect 50160 -28276 50272 -27762
rect 30860 -28380 33796 -28378
rect 33956 -29854 34016 -28378
rect 35992 -29854 36052 -28378
rect 36496 -29854 36556 -28378
rect 37004 -29854 37064 -28378
rect 37516 -29854 37576 -28378
rect 38030 -29854 38090 -28378
rect 40062 -29854 40122 -28378
rect 42102 -29854 42162 -28378
rect 42592 -29854 42652 -28378
rect 43112 -29854 43172 -28378
rect 43620 -29854 43680 -28378
rect 44134 -29854 44194 -28378
rect 46170 -29854 46230 -28378
rect 33956 -29914 46230 -29854
rect 33424 -30120 33430 -30060
rect 33490 -30120 33496 -30060
rect 31918 -30336 32996 -30276
rect 31918 -30516 31978 -30336
rect 32422 -30417 32482 -30336
rect 32214 -30423 32702 -30417
rect 32214 -30457 32226 -30423
rect 32690 -30457 32702 -30423
rect 32214 -30463 32702 -30457
rect 31918 -30556 31932 -30516
rect 31926 -31092 31932 -30556
rect 31966 -30556 31978 -30516
rect 32936 -30516 32996 -30336
rect 33430 -30417 33490 -30120
rect 33956 -30306 34016 -29914
rect 34506 -30120 34512 -30060
rect 34572 -30120 34578 -30060
rect 35464 -30120 35470 -30060
rect 35530 -30120 35536 -30060
rect 33950 -30366 33956 -30306
rect 34016 -30366 34022 -30306
rect 33232 -30423 33720 -30417
rect 33232 -30457 33244 -30423
rect 33708 -30457 33720 -30423
rect 33232 -30463 33720 -30457
rect 32936 -30542 32950 -30516
rect 31966 -31092 31972 -30556
rect 32944 -31056 32950 -30542
rect 31926 -31104 31972 -31092
rect 32938 -31092 32950 -31056
rect 32984 -30542 32996 -30516
rect 33956 -30516 34016 -30366
rect 34512 -30417 34572 -30120
rect 35470 -30417 35530 -30120
rect 35992 -30306 36052 -29914
rect 35986 -30366 35992 -30306
rect 36052 -30366 36058 -30306
rect 34250 -30423 34738 -30417
rect 34250 -30457 34262 -30423
rect 34726 -30457 34738 -30423
rect 34250 -30463 34738 -30457
rect 35268 -30423 35756 -30417
rect 35268 -30457 35280 -30423
rect 35744 -30457 35756 -30423
rect 35268 -30463 35756 -30457
rect 35470 -30466 35530 -30463
rect 33956 -30540 33968 -30516
rect 32984 -31056 32990 -30542
rect 33962 -31052 33968 -30540
rect 32984 -31092 32998 -31056
rect 32214 -31151 32702 -31145
rect 32214 -31185 32226 -31151
rect 32690 -31185 32702 -31151
rect 32214 -31191 32702 -31185
rect 32938 -31238 32998 -31092
rect 33958 -31092 33968 -31052
rect 34002 -30540 34016 -30516
rect 34980 -30516 35026 -30504
rect 34002 -31052 34008 -30540
rect 34002 -31092 34018 -31052
rect 34980 -31064 34986 -30516
rect 33442 -31145 33502 -31144
rect 33232 -31151 33720 -31145
rect 33232 -31185 33244 -31151
rect 33708 -31185 33720 -31151
rect 33232 -31191 33720 -31185
rect 31768 -31298 31774 -31238
rect 31834 -31298 31840 -31238
rect 32932 -31298 32938 -31238
rect 32998 -31298 33004 -31238
rect 31638 -31502 31644 -31442
rect 31704 -31502 31710 -31442
rect 29630 -33686 29636 -33626
rect 29696 -33686 29702 -33626
rect 27458 -37002 28680 -36942
rect 27458 -38918 27518 -37002
rect 27600 -37166 27660 -37002
rect 28112 -37067 28172 -37002
rect 27896 -37073 28384 -37067
rect 27896 -37107 27908 -37073
rect 28372 -37107 28384 -37073
rect 27896 -37113 28384 -37107
rect 27600 -37216 27614 -37166
rect 27608 -37742 27614 -37216
rect 27648 -37216 27660 -37166
rect 28620 -37166 28680 -37002
rect 28914 -37073 29402 -37067
rect 28914 -37107 28926 -37073
rect 29390 -37107 29402 -37073
rect 28914 -37113 29402 -37107
rect 27648 -37742 27654 -37216
rect 28620 -37218 28632 -37166
rect 27608 -37754 27654 -37742
rect 28626 -37742 28632 -37218
rect 28666 -37218 28680 -37166
rect 29636 -37166 29696 -33686
rect 31644 -34058 31704 -31502
rect 31774 -33912 31834 -31298
rect 32932 -31502 32938 -31442
rect 32998 -31502 33004 -31442
rect 32214 -31559 32702 -31553
rect 32214 -31593 32226 -31559
rect 32690 -31593 32702 -31559
rect 32214 -31599 32702 -31593
rect 31926 -31652 31972 -31640
rect 31926 -32192 31932 -31652
rect 31920 -32228 31932 -32192
rect 31966 -32192 31972 -31652
rect 32938 -31652 32998 -31502
rect 33442 -31553 33502 -31191
rect 33232 -31559 33720 -31553
rect 33232 -31593 33244 -31559
rect 33708 -31593 33720 -31559
rect 33232 -31599 33720 -31593
rect 33442 -31602 33502 -31599
rect 32938 -31690 32950 -31652
rect 31966 -32228 31980 -32192
rect 32944 -32198 32950 -31690
rect 31920 -32378 31980 -32228
rect 32938 -32228 32950 -32198
rect 32984 -31690 32998 -31652
rect 33958 -31652 34018 -31092
rect 34974 -31092 34986 -31064
rect 35020 -31064 35026 -30516
rect 35992 -30516 36052 -30366
rect 36496 -30417 36556 -29914
rect 36286 -30423 36774 -30417
rect 36286 -30457 36298 -30423
rect 36762 -30457 36774 -30423
rect 36286 -30463 36774 -30457
rect 35992 -30540 36004 -30516
rect 35998 -31034 36004 -30540
rect 35020 -31092 35034 -31064
rect 34250 -31151 34738 -31145
rect 34250 -31185 34262 -31151
rect 34726 -31185 34738 -31151
rect 34250 -31191 34738 -31185
rect 34974 -31342 35034 -31092
rect 35982 -31092 36004 -31034
rect 36038 -30540 36052 -30516
rect 37004 -30516 37064 -29914
rect 37516 -30417 37576 -29914
rect 38030 -30304 38090 -29914
rect 38528 -30120 38534 -30060
rect 38594 -30120 38600 -30060
rect 39546 -30120 39552 -30060
rect 39612 -30120 39618 -30060
rect 38024 -30364 38030 -30304
rect 38090 -30364 38096 -30304
rect 37304 -30423 37792 -30417
rect 37304 -30457 37316 -30423
rect 37780 -30457 37792 -30423
rect 37304 -30463 37792 -30457
rect 36038 -31034 36044 -30540
rect 37004 -30586 37022 -30516
rect 36038 -31092 36046 -31034
rect 35268 -31151 35756 -31145
rect 35268 -31185 35280 -31151
rect 35744 -31185 35756 -31151
rect 35268 -31191 35756 -31185
rect 34968 -31402 34974 -31342
rect 35034 -31402 35040 -31342
rect 34250 -31559 34738 -31553
rect 34250 -31593 34262 -31559
rect 34726 -31593 34738 -31559
rect 34250 -31599 34738 -31593
rect 35268 -31559 35756 -31553
rect 35268 -31593 35280 -31559
rect 35744 -31593 35756 -31559
rect 35268 -31599 35756 -31593
rect 32984 -32198 32990 -31690
rect 33958 -31692 33968 -31652
rect 32984 -32228 32998 -32198
rect 33962 -32202 33968 -31692
rect 32214 -32287 32702 -32281
rect 32214 -32321 32226 -32287
rect 32690 -32321 32702 -32287
rect 32214 -32327 32702 -32321
rect 32432 -32378 32492 -32327
rect 32938 -32378 32998 -32228
rect 33954 -32228 33968 -32202
rect 34002 -31692 34018 -31652
rect 34980 -31652 35026 -31640
rect 34002 -32202 34008 -31692
rect 34002 -32228 34014 -32202
rect 34980 -32208 34986 -31652
rect 33424 -32281 33484 -32274
rect 33232 -32287 33720 -32281
rect 33232 -32321 33244 -32287
rect 33708 -32321 33720 -32287
rect 33232 -32327 33720 -32321
rect 31920 -32438 32998 -32378
rect 32932 -32582 32992 -32580
rect 31922 -32642 32992 -32582
rect 31922 -32788 31982 -32642
rect 32432 -32689 32492 -32642
rect 32214 -32695 32702 -32689
rect 32214 -32729 32226 -32695
rect 32690 -32729 32702 -32695
rect 32214 -32735 32702 -32729
rect 31922 -32820 31932 -32788
rect 31926 -33364 31932 -32820
rect 31966 -32820 31982 -32788
rect 32932 -32788 32992 -32642
rect 33424 -32592 33484 -32327
rect 33424 -32689 33484 -32652
rect 33954 -32374 34014 -32228
rect 34972 -32228 34986 -32208
rect 35020 -32208 35026 -31652
rect 35982 -31652 36046 -31092
rect 37016 -31092 37022 -30586
rect 37056 -30586 37064 -30516
rect 38030 -30516 38090 -30364
rect 38534 -30417 38594 -30120
rect 39552 -30417 39612 -30120
rect 40062 -30304 40122 -29914
rect 40570 -30120 40576 -30060
rect 40636 -30120 40642 -30060
rect 41582 -30120 41588 -30060
rect 41648 -30120 41654 -30060
rect 40054 -30364 40060 -30304
rect 40120 -30364 40126 -30304
rect 38322 -30423 38810 -30417
rect 38322 -30457 38334 -30423
rect 38798 -30457 38810 -30423
rect 38322 -30463 38810 -30457
rect 39340 -30423 39828 -30417
rect 39340 -30457 39352 -30423
rect 39816 -30457 39828 -30423
rect 39340 -30463 39828 -30457
rect 38030 -30556 38040 -30516
rect 37056 -31092 37062 -30586
rect 38034 -31038 38040 -30556
rect 37016 -31104 37062 -31092
rect 38018 -31092 38040 -31038
rect 38074 -30556 38090 -30516
rect 39052 -30516 39098 -30504
rect 38074 -31038 38080 -30556
rect 38074 -31092 38082 -31038
rect 39052 -31052 39058 -30516
rect 36286 -31151 36774 -31145
rect 36286 -31185 36298 -31151
rect 36762 -31185 36774 -31151
rect 36286 -31191 36774 -31185
rect 37304 -31151 37792 -31145
rect 37304 -31185 37316 -31151
rect 37780 -31185 37792 -31151
rect 37304 -31191 37792 -31185
rect 37004 -31402 37010 -31342
rect 37070 -31402 37076 -31342
rect 36286 -31559 36774 -31553
rect 36286 -31593 36298 -31559
rect 36762 -31593 36774 -31559
rect 36286 -31599 36774 -31593
rect 35982 -31682 36004 -31652
rect 35998 -32200 36004 -31682
rect 35020 -32228 35032 -32208
rect 34452 -32281 34512 -32280
rect 34250 -32287 34738 -32281
rect 34250 -32321 34262 -32287
rect 34726 -32321 34738 -32287
rect 34250 -32327 34738 -32321
rect 34452 -32374 34512 -32327
rect 34972 -32374 35032 -32228
rect 35990 -32228 36004 -32200
rect 36038 -31682 36046 -31652
rect 37010 -31652 37070 -31402
rect 37304 -31559 37792 -31553
rect 37304 -31593 37316 -31559
rect 37780 -31593 37792 -31559
rect 37304 -31599 37792 -31593
rect 36038 -32200 36044 -31682
rect 37010 -31690 37022 -31652
rect 37016 -32192 37022 -31690
rect 36038 -32202 36050 -32200
rect 36038 -32228 36054 -32202
rect 35480 -32281 35540 -32276
rect 35268 -32287 35756 -32281
rect 35268 -32321 35280 -32287
rect 35744 -32321 35756 -32287
rect 35268 -32327 35756 -32321
rect 35480 -32374 35540 -32327
rect 33954 -32376 35540 -32374
rect 35990 -32376 36054 -32228
rect 37008 -32228 37022 -32192
rect 37056 -31690 37070 -31652
rect 38018 -31652 38082 -31092
rect 39048 -31092 39058 -31052
rect 39092 -31052 39098 -30516
rect 40062 -30516 40122 -30364
rect 40576 -30417 40636 -30120
rect 41588 -30417 41648 -30120
rect 42102 -30302 42162 -29914
rect 42096 -30362 42102 -30302
rect 42162 -30362 42168 -30302
rect 40358 -30423 40846 -30417
rect 40358 -30457 40370 -30423
rect 40834 -30457 40846 -30423
rect 40358 -30463 40846 -30457
rect 41376 -30423 41864 -30417
rect 41376 -30457 41388 -30423
rect 41852 -30457 41864 -30423
rect 41376 -30463 41864 -30457
rect 40062 -30556 40076 -30516
rect 40070 -31036 40076 -30556
rect 39092 -31092 39108 -31052
rect 38536 -31145 38596 -31142
rect 38322 -31151 38810 -31145
rect 38322 -31185 38334 -31151
rect 38798 -31185 38810 -31151
rect 38322 -31191 38810 -31185
rect 38536 -31553 38596 -31191
rect 39048 -31238 39108 -31092
rect 40060 -31092 40076 -31036
rect 40110 -30556 40122 -30516
rect 41088 -30516 41134 -30504
rect 40110 -31036 40116 -30556
rect 40110 -31092 40124 -31036
rect 41088 -31054 41094 -30516
rect 39554 -31145 39614 -31136
rect 39340 -31151 39828 -31145
rect 39340 -31185 39352 -31151
rect 39816 -31185 39828 -31151
rect 39340 -31191 39828 -31185
rect 39042 -31298 39048 -31238
rect 39108 -31298 39114 -31238
rect 39038 -31502 39044 -31442
rect 39104 -31502 39110 -31442
rect 38322 -31559 38810 -31553
rect 38322 -31593 38334 -31559
rect 38798 -31593 38810 -31559
rect 38322 -31599 38810 -31593
rect 38536 -31600 38596 -31599
rect 38018 -31686 38040 -31652
rect 37056 -32192 37062 -31690
rect 38034 -32192 38040 -31686
rect 37056 -32228 37072 -32192
rect 36286 -32287 36774 -32281
rect 36286 -32321 36298 -32287
rect 36762 -32321 36774 -32287
rect 36286 -32327 36774 -32321
rect 33954 -32434 35480 -32376
rect 33232 -32695 33720 -32689
rect 33232 -32729 33244 -32695
rect 33708 -32729 33720 -32695
rect 33232 -32735 33720 -32729
rect 32932 -32820 32950 -32788
rect 31966 -33364 31972 -32820
rect 32944 -33322 32950 -32820
rect 31926 -33376 31972 -33364
rect 32932 -33364 32950 -33322
rect 32984 -32820 32992 -32788
rect 33954 -32788 34014 -32434
rect 35984 -32436 35990 -32376
rect 36050 -32436 36056 -32376
rect 35480 -32442 35540 -32436
rect 34966 -32538 34972 -32474
rect 35036 -32538 35042 -32474
rect 34456 -32652 34462 -32592
rect 34522 -32652 34528 -32592
rect 34972 -32632 35036 -32538
rect 34462 -32689 34522 -32652
rect 34250 -32695 34738 -32689
rect 34250 -32729 34262 -32695
rect 34726 -32729 34738 -32695
rect 34250 -32735 34738 -32729
rect 32984 -33322 32990 -32820
rect 33954 -32840 33968 -32788
rect 32984 -33364 32996 -33322
rect 33962 -33328 33968 -32840
rect 32214 -33423 32702 -33417
rect 32214 -33457 32226 -33423
rect 32690 -33457 32702 -33423
rect 32214 -33463 32702 -33457
rect 32932 -33572 32996 -33364
rect 33954 -33364 33968 -33328
rect 34002 -32840 34014 -32788
rect 34972 -32788 35038 -32632
rect 35468 -32652 35474 -32592
rect 35534 -32652 35540 -32592
rect 35474 -32689 35534 -32652
rect 35268 -32695 35756 -32689
rect 35268 -32729 35280 -32695
rect 35744 -32729 35756 -32695
rect 35268 -32735 35756 -32729
rect 35474 -32736 35534 -32735
rect 34972 -32838 34986 -32788
rect 34002 -33328 34008 -32840
rect 34002 -33364 34014 -33328
rect 34980 -33340 34986 -32838
rect 33232 -33423 33720 -33417
rect 33232 -33457 33244 -33423
rect 33708 -33457 33720 -33423
rect 33232 -33463 33720 -33457
rect 32488 -33632 32996 -33572
rect 31768 -33972 31774 -33912
rect 31834 -33972 31840 -33912
rect 31644 -34118 32064 -34058
rect 32004 -36930 32064 -34118
rect 32124 -36380 32130 -36320
rect 32190 -36380 32196 -36320
rect 30654 -36998 31864 -36938
rect 31998 -36990 32004 -36930
rect 32064 -36990 32070 -36930
rect 29932 -37073 30420 -37067
rect 29932 -37107 29944 -37073
rect 30408 -37107 30420 -37073
rect 29932 -37113 30420 -37107
rect 28666 -37742 28672 -37218
rect 28626 -37754 28672 -37742
rect 29636 -37742 29650 -37166
rect 29684 -37742 29696 -37166
rect 30654 -37166 30714 -36998
rect 31166 -37067 31226 -36998
rect 30950 -37073 31438 -37067
rect 30950 -37107 30962 -37073
rect 31426 -37107 31438 -37073
rect 30950 -37113 31438 -37107
rect 30654 -37214 30668 -37166
rect 27896 -37801 28384 -37795
rect 27896 -37835 27908 -37801
rect 28372 -37835 28384 -37801
rect 27896 -37841 28384 -37835
rect 28914 -37801 29402 -37795
rect 28914 -37835 28926 -37801
rect 29390 -37835 29402 -37801
rect 28914 -37841 29402 -37835
rect 29120 -37884 29180 -37841
rect 29114 -37944 29120 -37884
rect 29180 -37944 29186 -37884
rect 29222 -38056 29228 -37996
rect 29288 -38056 29294 -37996
rect 29228 -38099 29288 -38056
rect 27896 -38105 28384 -38099
rect 27896 -38139 27908 -38105
rect 28372 -38139 28384 -38105
rect 27896 -38145 28384 -38139
rect 28914 -38105 29402 -38099
rect 28914 -38139 28926 -38105
rect 29390 -38139 29402 -38105
rect 28914 -38145 29402 -38139
rect 27608 -38198 27654 -38186
rect 27608 -38716 27614 -38198
rect 27598 -38774 27614 -38716
rect 27648 -38716 27654 -38198
rect 28626 -38198 28672 -38186
rect 27648 -38774 27658 -38716
rect 28626 -38724 28632 -38198
rect 27452 -38978 27458 -38918
rect 27518 -38978 27524 -38918
rect 27332 -40006 27392 -40000
rect 27458 -40006 27518 -38978
rect 27598 -39028 27658 -38774
rect 28618 -38774 28632 -38724
rect 28666 -38724 28672 -38198
rect 29636 -38198 29696 -37742
rect 30662 -37742 30668 -37214
rect 30702 -37214 30714 -37166
rect 31672 -37166 31732 -36998
rect 31672 -37212 31686 -37166
rect 30702 -37742 30708 -37214
rect 30662 -37754 30708 -37742
rect 31680 -37742 31686 -37212
rect 31720 -37212 31732 -37166
rect 31720 -37742 31726 -37212
rect 31680 -37754 31726 -37742
rect 29932 -37801 30420 -37795
rect 29932 -37835 29944 -37801
rect 30408 -37835 30420 -37801
rect 29932 -37841 30420 -37835
rect 30950 -37801 31438 -37795
rect 30950 -37835 30962 -37801
rect 31426 -37835 31438 -37801
rect 30950 -37841 31438 -37835
rect 30012 -37996 30072 -37841
rect 30136 -37944 30142 -37884
rect 30202 -37944 30208 -37884
rect 30006 -38056 30012 -37996
rect 30072 -38056 30078 -37996
rect 30142 -38099 30202 -37944
rect 29932 -38105 30420 -38099
rect 29932 -38139 29944 -38105
rect 30408 -38139 30420 -38105
rect 29932 -38145 30420 -38139
rect 30950 -38105 31438 -38099
rect 30950 -38139 30962 -38105
rect 31426 -38139 31438 -38105
rect 30950 -38145 31438 -38139
rect 28666 -38774 28678 -38724
rect 27896 -38833 28384 -38827
rect 27896 -38867 27908 -38833
rect 28372 -38867 28384 -38833
rect 27896 -38873 28384 -38867
rect 28100 -39028 28160 -38873
rect 28618 -39028 28678 -38774
rect 29636 -38774 29650 -38198
rect 29684 -38774 29696 -38198
rect 30662 -38198 30708 -38186
rect 30662 -38688 30668 -38198
rect 28914 -38833 29402 -38827
rect 28914 -38867 28926 -38833
rect 29390 -38867 29402 -38833
rect 28914 -38873 29402 -38867
rect 27598 -39088 28618 -39028
rect 28678 -39088 28684 -39028
rect 27598 -39230 27658 -39088
rect 28100 -39131 28160 -39088
rect 27896 -39137 28384 -39131
rect 27896 -39171 27908 -39137
rect 28372 -39171 28384 -39137
rect 27896 -39177 28384 -39171
rect 27598 -39290 27614 -39230
rect 27608 -39806 27614 -39290
rect 27648 -39290 27658 -39230
rect 28618 -39230 28678 -39088
rect 29128 -39131 29188 -38873
rect 28914 -39137 29402 -39131
rect 28914 -39171 28926 -39137
rect 29390 -39171 29402 -39137
rect 28914 -39177 29402 -39171
rect 27648 -39806 27654 -39290
rect 28618 -39294 28632 -39230
rect 27608 -39818 27654 -39806
rect 28626 -39806 28632 -39294
rect 28666 -39294 28678 -39230
rect 29636 -39230 29696 -38774
rect 30652 -38774 30668 -38688
rect 30702 -38688 30708 -38198
rect 31680 -38198 31726 -38186
rect 30702 -38774 30712 -38688
rect 31680 -38728 31686 -38198
rect 29932 -38833 30420 -38827
rect 29932 -38867 29944 -38833
rect 30408 -38867 30420 -38833
rect 29932 -38873 30420 -38867
rect 30146 -39131 30206 -38873
rect 30652 -38918 30712 -38774
rect 31672 -38774 31686 -38728
rect 31720 -38728 31726 -38198
rect 31720 -38774 31732 -38728
rect 30950 -38833 31438 -38827
rect 30950 -38867 30962 -38833
rect 31426 -38867 31438 -38833
rect 30950 -38873 31438 -38867
rect 31166 -38918 31226 -38873
rect 31672 -38918 31732 -38774
rect 30646 -38978 30652 -38918
rect 30712 -38978 31732 -38918
rect 29932 -39137 30420 -39131
rect 29932 -39171 29944 -39137
rect 30408 -39171 30420 -39137
rect 29932 -39177 30420 -39171
rect 28666 -39806 28672 -39294
rect 28626 -39818 28672 -39806
rect 29636 -39806 29650 -39230
rect 29684 -39806 29696 -39230
rect 30652 -39230 30712 -38978
rect 31166 -39131 31226 -38978
rect 30950 -39137 31438 -39131
rect 30950 -39171 30962 -39137
rect 31426 -39171 31438 -39137
rect 30950 -39177 31438 -39171
rect 30652 -39286 30668 -39230
rect 27896 -39865 28384 -39859
rect 27896 -39899 27908 -39865
rect 28372 -39899 28384 -39865
rect 27896 -39905 28384 -39899
rect 28914 -39865 29402 -39859
rect 28914 -39899 28926 -39865
rect 29390 -39899 29402 -39865
rect 28914 -39905 29402 -39899
rect 29134 -39952 29194 -39905
rect 27392 -40066 28682 -40006
rect 29128 -40012 29134 -39952
rect 29194 -40012 29200 -39952
rect 27332 -40072 27392 -40066
rect 27596 -40262 27656 -40066
rect 28104 -40163 28164 -40066
rect 27896 -40169 28384 -40163
rect 27896 -40203 27908 -40169
rect 28372 -40203 28384 -40169
rect 27896 -40209 28384 -40203
rect 27596 -40314 27614 -40262
rect 27608 -40838 27614 -40314
rect 27648 -40314 27656 -40262
rect 28622 -40262 28682 -40066
rect 29234 -40112 29240 -40052
rect 29300 -40112 29306 -40052
rect 29240 -40163 29300 -40112
rect 28914 -40169 29402 -40163
rect 28914 -40203 28926 -40169
rect 29390 -40203 29402 -40169
rect 28914 -40209 29402 -40203
rect 28622 -40310 28632 -40262
rect 27648 -40838 27654 -40314
rect 27608 -40850 27654 -40838
rect 28626 -40838 28632 -40310
rect 28666 -40310 28682 -40262
rect 29636 -40262 29696 -39806
rect 30662 -39806 30668 -39286
rect 30702 -39286 30712 -39230
rect 31672 -39230 31732 -38978
rect 31804 -39028 31864 -36998
rect 31798 -39088 31804 -39028
rect 31864 -39088 31870 -39028
rect 31672 -39266 31686 -39230
rect 30702 -39806 30708 -39286
rect 30662 -39818 30708 -39806
rect 31680 -39806 31686 -39266
rect 31720 -39266 31732 -39230
rect 31720 -39806 31726 -39266
rect 31680 -39818 31726 -39806
rect 29932 -39865 30420 -39859
rect 29932 -39899 29944 -39865
rect 30408 -39899 30420 -39865
rect 29932 -39905 30420 -39899
rect 30950 -39865 31438 -39859
rect 30950 -39899 30962 -39865
rect 31426 -39899 31438 -39865
rect 30950 -39905 31438 -39899
rect 30026 -40052 30086 -39905
rect 30138 -40012 30144 -39952
rect 30204 -40012 30210 -39952
rect 31804 -40006 31864 -39088
rect 31990 -39216 31996 -39156
rect 32056 -39216 32062 -39156
rect 30020 -40112 30026 -40052
rect 30086 -40112 30092 -40052
rect 30144 -40163 30204 -40012
rect 30652 -40066 31864 -40006
rect 29932 -40169 30420 -40163
rect 29932 -40203 29944 -40169
rect 30408 -40203 30420 -40169
rect 29932 -40209 30420 -40203
rect 28666 -40838 28672 -40310
rect 29636 -40336 29650 -40262
rect 28626 -40850 28672 -40838
rect 29644 -40838 29650 -40336
rect 29684 -40336 29696 -40262
rect 30652 -40262 30712 -40066
rect 31154 -40163 31214 -40066
rect 30950 -40169 31438 -40163
rect 30950 -40203 30962 -40169
rect 31426 -40203 31438 -40169
rect 30950 -40209 31438 -40203
rect 30652 -40292 30668 -40262
rect 29684 -40838 29690 -40336
rect 30662 -40756 30668 -40292
rect 29644 -40850 29690 -40838
rect 30654 -40838 30668 -40756
rect 30702 -40292 30712 -40262
rect 31672 -40262 31732 -40066
rect 30702 -40756 30708 -40292
rect 31672 -40330 31686 -40262
rect 30702 -40838 30714 -40756
rect 30132 -40891 30192 -40887
rect 27896 -40897 28384 -40891
rect 27896 -40931 27908 -40897
rect 28372 -40931 28384 -40897
rect 27896 -40937 28384 -40931
rect 28914 -40897 29402 -40891
rect 28914 -40931 28926 -40897
rect 29390 -40931 29402 -40897
rect 28914 -40937 29402 -40931
rect 29932 -40897 30420 -40891
rect 29932 -40931 29944 -40897
rect 30408 -40931 30420 -40897
rect 29932 -40937 30420 -40931
rect 26846 -41062 26906 -41056
rect 29126 -41062 29186 -40937
rect 26906 -41122 29186 -41062
rect 26846 -41128 26906 -41122
rect 26986 -41238 27046 -41232
rect 30132 -41238 30192 -40937
rect 27046 -41240 30192 -41238
rect 27046 -41298 30132 -41240
rect 26986 -41304 27046 -41298
rect 30132 -41306 30192 -41300
rect 27886 -41412 27946 -41406
rect 30654 -41412 30714 -40838
rect 31680 -40838 31686 -40330
rect 31720 -40330 31732 -40262
rect 31720 -40838 31726 -40330
rect 31680 -40850 31726 -40838
rect 30950 -40897 31438 -40891
rect 30950 -40931 30962 -40897
rect 31426 -40931 31438 -40897
rect 30950 -40937 31438 -40931
rect 27946 -41472 30714 -41412
rect 27886 -41478 27946 -41472
rect 26726 -41562 26786 -41556
rect 31996 -41562 32056 -39216
rect 32130 -40308 32190 -36380
rect 32240 -36990 32246 -36930
rect 32306 -36990 32312 -36930
rect 32246 -39052 32306 -36990
rect 32488 -37894 32548 -33632
rect 32932 -33762 32996 -33632
rect 32926 -33826 32932 -33762
rect 32996 -33826 33002 -33762
rect 32756 -33912 32816 -33906
rect 32756 -36848 32816 -33972
rect 33434 -34018 33494 -33463
rect 33954 -33514 34014 -33364
rect 34970 -33364 34986 -33340
rect 35020 -32834 35038 -32788
rect 35990 -32788 36054 -32436
rect 36484 -32584 36544 -32327
rect 37008 -32474 37072 -32228
rect 38024 -32228 38040 -32192
rect 38074 -31686 38082 -31652
rect 39044 -31652 39104 -31502
rect 39554 -31553 39614 -31191
rect 39340 -31559 39828 -31553
rect 39340 -31593 39352 -31559
rect 39816 -31593 39828 -31559
rect 39340 -31599 39828 -31593
rect 39044 -31678 39058 -31652
rect 38074 -32192 38080 -31686
rect 38074 -32194 38084 -32192
rect 38074 -32228 38088 -32194
rect 37304 -32287 37792 -32281
rect 37304 -32321 37316 -32287
rect 37780 -32321 37792 -32287
rect 37304 -32327 37792 -32321
rect 36842 -32538 36848 -32474
rect 36912 -32538 37072 -32474
rect 37508 -32584 37568 -32327
rect 38024 -32376 38088 -32228
rect 39052 -32228 39058 -31678
rect 39092 -31678 39104 -31652
rect 40060 -31652 40124 -31092
rect 41082 -31092 41094 -31054
rect 41128 -31054 41134 -30516
rect 42102 -30516 42162 -30362
rect 42592 -30417 42652 -29914
rect 43112 -30302 43172 -29914
rect 43106 -30362 43112 -30302
rect 43172 -30362 43178 -30302
rect 42394 -30423 42882 -30417
rect 42394 -30457 42406 -30423
rect 42870 -30457 42882 -30423
rect 42394 -30463 42882 -30457
rect 42102 -30554 42112 -30516
rect 42106 -31052 42112 -30554
rect 41128 -31092 41142 -31054
rect 40570 -31145 40630 -31139
rect 40358 -31151 40846 -31145
rect 40358 -31185 40370 -31151
rect 40834 -31185 40846 -31151
rect 40358 -31191 40846 -31185
rect 40570 -31553 40630 -31191
rect 41082 -31238 41142 -31092
rect 42098 -31092 42112 -31052
rect 42146 -30554 42162 -30516
rect 43112 -30516 43172 -30362
rect 43620 -30417 43680 -29914
rect 44134 -30302 44194 -29914
rect 44640 -30120 44646 -30060
rect 44706 -30120 44712 -30060
rect 45652 -30120 45658 -30060
rect 45718 -30120 45724 -30060
rect 44128 -30362 44134 -30302
rect 44194 -30362 44200 -30302
rect 43412 -30423 43900 -30417
rect 43412 -30457 43424 -30423
rect 43888 -30457 43900 -30423
rect 43412 -30463 43900 -30457
rect 43620 -30466 43680 -30463
rect 42146 -31052 42152 -30554
rect 43112 -30586 43130 -30516
rect 42146 -31092 42162 -31052
rect 41582 -31145 41642 -31139
rect 41376 -31151 41864 -31145
rect 41376 -31185 41388 -31151
rect 41852 -31185 41864 -31151
rect 41376 -31191 41864 -31185
rect 41076 -31298 41082 -31238
rect 41142 -31298 41148 -31238
rect 41582 -31442 41642 -31191
rect 41074 -31502 41080 -31442
rect 41140 -31502 41146 -31442
rect 41576 -31502 41582 -31442
rect 41642 -31502 41648 -31442
rect 40358 -31559 40846 -31553
rect 40358 -31593 40370 -31559
rect 40834 -31593 40846 -31559
rect 40358 -31599 40846 -31593
rect 40570 -31602 40630 -31599
rect 39092 -32228 39098 -31678
rect 40060 -31684 40076 -31652
rect 40070 -32180 40076 -31684
rect 39052 -32240 39098 -32228
rect 40062 -32228 40076 -32180
rect 40110 -31684 40124 -31652
rect 41080 -31652 41140 -31502
rect 41582 -31553 41642 -31502
rect 41376 -31559 41864 -31553
rect 41376 -31593 41388 -31559
rect 41852 -31593 41864 -31559
rect 41376 -31599 41864 -31593
rect 41582 -31602 41642 -31599
rect 41080 -31684 41094 -31652
rect 40110 -32180 40116 -31684
rect 40110 -32182 40122 -32180
rect 40110 -32228 40126 -32182
rect 41088 -32198 41094 -31684
rect 38536 -32281 38596 -32274
rect 38322 -32287 38810 -32281
rect 38322 -32321 38334 -32287
rect 38798 -32321 38810 -32287
rect 38322 -32327 38810 -32321
rect 39340 -32287 39828 -32281
rect 39340 -32321 39352 -32287
rect 39816 -32321 39828 -32287
rect 39340 -32327 39828 -32321
rect 38018 -32436 38024 -32376
rect 38084 -32436 38090 -32376
rect 36478 -32644 36484 -32584
rect 36544 -32644 36550 -32584
rect 37502 -32644 37508 -32584
rect 37568 -32644 37574 -32584
rect 36286 -32695 36774 -32689
rect 36286 -32729 36298 -32695
rect 36762 -32729 36774 -32695
rect 36286 -32735 36774 -32729
rect 37304 -32695 37792 -32689
rect 37304 -32729 37316 -32695
rect 37780 -32729 37792 -32695
rect 37304 -32735 37792 -32729
rect 35020 -32838 35036 -32834
rect 35990 -32836 36004 -32788
rect 35020 -33340 35026 -32838
rect 35998 -33338 36004 -32836
rect 35020 -33364 35034 -33340
rect 34250 -33423 34738 -33417
rect 34250 -33457 34262 -33423
rect 34726 -33457 34738 -33423
rect 34250 -33463 34738 -33457
rect 33948 -33574 33954 -33514
rect 34014 -33574 34020 -33514
rect 34476 -34018 34536 -33463
rect 34970 -33624 35034 -33364
rect 35990 -33364 36004 -33338
rect 36038 -32836 36054 -32788
rect 37016 -32788 37062 -32776
rect 36038 -33338 36044 -32836
rect 37016 -33308 37022 -32788
rect 36038 -33340 36050 -33338
rect 36038 -33364 36054 -33340
rect 35268 -33423 35756 -33417
rect 35268 -33457 35280 -33423
rect 35744 -33457 35756 -33423
rect 35268 -33463 35756 -33457
rect 34964 -33688 34970 -33624
rect 35034 -33688 35040 -33624
rect 35476 -34018 35536 -33463
rect 35990 -33514 36054 -33364
rect 37010 -33364 37022 -33308
rect 37056 -33308 37062 -32788
rect 38024 -32788 38088 -32436
rect 38536 -32584 38596 -32327
rect 38530 -32644 38536 -32584
rect 38596 -32644 38602 -32584
rect 38536 -32689 38596 -32644
rect 39564 -32689 39624 -32327
rect 40062 -32378 40126 -32228
rect 41082 -32228 41094 -32198
rect 41128 -31684 41140 -31652
rect 42098 -31652 42162 -31092
rect 43124 -31092 43130 -30586
rect 43164 -30586 43172 -30516
rect 44134 -30516 44194 -30362
rect 44646 -30417 44706 -30120
rect 45658 -30417 45718 -30120
rect 46170 -30302 46230 -29914
rect 46670 -30120 46676 -30060
rect 46736 -30120 46742 -30060
rect 46164 -30362 46170 -30302
rect 46230 -30362 46236 -30302
rect 44430 -30423 44918 -30417
rect 44430 -30457 44442 -30423
rect 44906 -30457 44918 -30423
rect 44430 -30463 44918 -30457
rect 45448 -30423 45936 -30417
rect 45448 -30457 45460 -30423
rect 45924 -30457 45936 -30423
rect 45448 -30463 45936 -30457
rect 44134 -30544 44148 -30516
rect 43164 -31092 43170 -30586
rect 44142 -31044 44148 -30544
rect 43124 -31104 43170 -31092
rect 44134 -31092 44148 -31044
rect 44182 -30544 44194 -30516
rect 45160 -30516 45206 -30504
rect 44182 -31044 44188 -30544
rect 44182 -31092 44194 -31044
rect 45160 -31060 45166 -30516
rect 42394 -31151 42882 -31145
rect 42394 -31185 42406 -31151
rect 42870 -31185 42882 -31151
rect 42394 -31191 42882 -31185
rect 43412 -31151 43900 -31145
rect 43412 -31185 43424 -31151
rect 43888 -31185 43900 -31151
rect 43412 -31191 43900 -31185
rect 43110 -31402 43116 -31342
rect 43176 -31402 43182 -31342
rect 42596 -31502 42602 -31442
rect 42662 -31502 42668 -31442
rect 42602 -31553 42662 -31502
rect 42394 -31559 42882 -31553
rect 42394 -31593 42406 -31559
rect 42870 -31593 42882 -31559
rect 42394 -31599 42882 -31593
rect 41128 -32198 41134 -31684
rect 42098 -31700 42112 -31652
rect 42106 -32184 42112 -31700
rect 41128 -32228 41142 -32198
rect 40582 -32281 40642 -32269
rect 40358 -32287 40846 -32281
rect 40358 -32321 40370 -32287
rect 40834 -32321 40846 -32287
rect 40358 -32327 40846 -32321
rect 40056 -32438 40062 -32378
rect 40122 -32438 40128 -32378
rect 38322 -32695 38810 -32689
rect 38322 -32729 38334 -32695
rect 38798 -32729 38810 -32695
rect 38322 -32735 38810 -32729
rect 39340 -32695 39828 -32689
rect 39340 -32729 39352 -32695
rect 39816 -32729 39828 -32695
rect 39340 -32735 39828 -32729
rect 39564 -32742 39624 -32735
rect 38024 -32848 38040 -32788
rect 37056 -33364 37070 -33308
rect 38034 -33330 38040 -32848
rect 36512 -33417 36572 -33414
rect 36286 -33423 36774 -33417
rect 36286 -33457 36298 -33423
rect 36762 -33457 36774 -33423
rect 36286 -33463 36774 -33457
rect 36512 -33514 36572 -33463
rect 37010 -33514 37070 -33364
rect 38024 -33364 38040 -33330
rect 38074 -32848 38088 -32788
rect 39052 -32788 39098 -32776
rect 38074 -33330 38080 -32848
rect 38074 -33332 38084 -33330
rect 39052 -33332 39058 -32788
rect 38074 -33364 38088 -33332
rect 37304 -33423 37792 -33417
rect 37304 -33457 37316 -33423
rect 37780 -33457 37792 -33423
rect 37304 -33463 37792 -33457
rect 35984 -33574 35990 -33514
rect 36050 -33574 36056 -33514
rect 36506 -33574 36512 -33514
rect 36572 -33574 36578 -33514
rect 37004 -33574 37010 -33514
rect 37070 -33574 37076 -33514
rect 37484 -33518 37544 -33463
rect 38024 -33510 38088 -33364
rect 39042 -33364 39058 -33332
rect 39092 -33332 39098 -32788
rect 40062 -32788 40126 -32438
rect 40582 -32689 40642 -32327
rect 41082 -32476 41142 -32228
rect 42098 -32228 42112 -32184
rect 42146 -31700 42162 -31652
rect 43116 -31652 43176 -31402
rect 43622 -31502 43628 -31442
rect 43688 -31502 43694 -31442
rect 44134 -31446 44194 -31092
rect 45150 -31092 45166 -31060
rect 45200 -31060 45206 -30516
rect 46170 -30516 46230 -30362
rect 46676 -30417 46736 -30120
rect 47190 -30354 48270 -30294
rect 46466 -30423 46954 -30417
rect 46466 -30457 46478 -30423
rect 46942 -30457 46954 -30423
rect 46466 -30463 46954 -30457
rect 46170 -30548 46184 -30516
rect 46178 -31054 46184 -30548
rect 45200 -31092 45210 -31060
rect 44430 -31151 44918 -31145
rect 44430 -31185 44442 -31151
rect 44906 -31185 44918 -31151
rect 44430 -31191 44918 -31185
rect 45150 -31342 45210 -31092
rect 46174 -31092 46184 -31054
rect 46218 -30548 46230 -30516
rect 47190 -30516 47250 -30354
rect 47692 -30417 47752 -30354
rect 47484 -30423 47972 -30417
rect 47484 -30457 47496 -30423
rect 47960 -30457 47972 -30423
rect 47484 -30463 47972 -30457
rect 47190 -30546 47202 -30516
rect 46218 -31054 46224 -30548
rect 47196 -31052 47202 -30546
rect 46218 -31092 46234 -31054
rect 45448 -31151 45936 -31145
rect 45448 -31185 45460 -31151
rect 45924 -31185 45936 -31151
rect 45448 -31191 45936 -31185
rect 45144 -31402 45150 -31342
rect 45210 -31402 45216 -31342
rect 46174 -31440 46234 -31092
rect 47190 -31092 47202 -31052
rect 47236 -30546 47250 -30516
rect 48210 -30516 48270 -30354
rect 47236 -31052 47242 -30546
rect 48210 -30562 48220 -30516
rect 47236 -31092 47250 -31052
rect 46654 -31145 46714 -31133
rect 46466 -31151 46954 -31145
rect 46466 -31185 46478 -31151
rect 46942 -31185 46954 -31151
rect 46466 -31191 46954 -31185
rect 46174 -31446 46238 -31440
rect 43628 -31553 43688 -31502
rect 44128 -31506 44134 -31446
rect 44194 -31506 44200 -31446
rect 44642 -31506 44648 -31446
rect 44708 -31506 44714 -31446
rect 45146 -31506 45152 -31446
rect 45212 -31506 45218 -31446
rect 45652 -31506 45658 -31446
rect 45718 -31506 45724 -31446
rect 46174 -31506 46178 -31446
rect 43412 -31559 43900 -31553
rect 43412 -31593 43424 -31559
rect 43888 -31593 43900 -31559
rect 43412 -31599 43900 -31593
rect 43116 -31676 43130 -31652
rect 42146 -32184 42152 -31700
rect 42146 -32186 42158 -32184
rect 42146 -32228 42162 -32186
rect 41582 -32281 41642 -32273
rect 41376 -32287 41864 -32281
rect 41376 -32321 41388 -32287
rect 41852 -32321 41864 -32287
rect 41376 -32327 41864 -32321
rect 41076 -32536 41082 -32476
rect 41142 -32536 41148 -32476
rect 41582 -32689 41642 -32327
rect 42098 -32378 42162 -32228
rect 43124 -32228 43130 -31676
rect 43164 -31676 43176 -31652
rect 44134 -31652 44194 -31506
rect 44648 -31553 44708 -31506
rect 44430 -31559 44918 -31553
rect 44430 -31593 44442 -31559
rect 44906 -31593 44918 -31559
rect 44430 -31599 44918 -31593
rect 43164 -32228 43170 -31676
rect 44134 -31696 44148 -31652
rect 44142 -32192 44148 -31696
rect 43124 -32240 43170 -32228
rect 44134 -32228 44148 -32192
rect 44182 -31696 44194 -31652
rect 45152 -31652 45212 -31506
rect 45658 -31553 45718 -31506
rect 46174 -31512 46238 -31506
rect 45448 -31559 45936 -31553
rect 45448 -31593 45460 -31559
rect 45924 -31593 45936 -31559
rect 45448 -31599 45936 -31593
rect 45152 -31680 45166 -31652
rect 44182 -32192 44188 -31696
rect 45160 -32158 45166 -31680
rect 44182 -32228 44194 -32192
rect 42394 -32287 42882 -32281
rect 42394 -32321 42406 -32287
rect 42870 -32321 42882 -32287
rect 42394 -32327 42882 -32321
rect 43412 -32287 43900 -32281
rect 43412 -32321 43424 -32287
rect 43888 -32321 43900 -32287
rect 43412 -32327 43900 -32321
rect 44134 -32378 44194 -32228
rect 45150 -32228 45166 -32158
rect 45200 -31680 45212 -31652
rect 46174 -31652 46234 -31512
rect 46654 -31553 46714 -31191
rect 47190 -31238 47250 -31092
rect 48214 -31092 48220 -30562
rect 48254 -30562 48270 -30516
rect 48254 -31092 48260 -30562
rect 48214 -31104 48260 -31092
rect 47484 -31151 47972 -31145
rect 47484 -31185 47496 -31151
rect 47960 -31185 47972 -31151
rect 47484 -31191 47972 -31185
rect 47184 -31298 47190 -31238
rect 47250 -31298 47256 -31238
rect 48434 -31298 48440 -31238
rect 48500 -31298 48506 -31238
rect 47194 -31514 48264 -31454
rect 46466 -31559 46954 -31553
rect 46466 -31593 46478 -31559
rect 46942 -31593 46954 -31559
rect 46466 -31599 46954 -31593
rect 45200 -32158 45206 -31680
rect 46174 -31688 46184 -31652
rect 45200 -32228 45210 -32158
rect 46178 -32196 46184 -31688
rect 44430 -32287 44918 -32281
rect 44430 -32321 44442 -32287
rect 44906 -32321 44918 -32287
rect 44430 -32327 44918 -32321
rect 44636 -32378 44696 -32327
rect 42092 -32438 42098 -32378
rect 42158 -32438 42164 -32378
rect 42592 -32438 42598 -32378
rect 42658 -32438 42664 -32378
rect 43106 -32438 43112 -32378
rect 43172 -32438 43178 -32378
rect 43630 -32438 43636 -32378
rect 43696 -32438 43702 -32378
rect 44128 -32438 44134 -32378
rect 44194 -32438 44200 -32378
rect 44630 -32438 44636 -32378
rect 44696 -32438 44702 -32378
rect 45150 -32380 45210 -32228
rect 46168 -32228 46184 -32196
rect 46218 -31688 46234 -31652
rect 47194 -31652 47254 -31514
rect 47700 -31553 47760 -31514
rect 47484 -31559 47972 -31553
rect 47484 -31593 47496 -31559
rect 47960 -31593 47972 -31559
rect 47484 -31599 47972 -31593
rect 47194 -31680 47202 -31652
rect 46218 -32196 46224 -31688
rect 46218 -32198 46228 -32196
rect 47196 -32198 47202 -31680
rect 46218 -32228 46232 -32198
rect 45658 -32281 45718 -32274
rect 45448 -32287 45936 -32281
rect 45448 -32321 45460 -32287
rect 45924 -32321 45936 -32287
rect 45448 -32327 45936 -32321
rect 45658 -32380 45718 -32327
rect 46168 -32380 46232 -32228
rect 47190 -32228 47202 -32198
rect 47236 -31680 47254 -31652
rect 48204 -31652 48264 -31514
rect 47236 -32198 47242 -31680
rect 48204 -31686 48220 -31652
rect 47236 -32228 47250 -32198
rect 46654 -32281 46714 -32275
rect 46466 -32287 46954 -32281
rect 46466 -32321 46478 -32287
rect 46942 -32321 46954 -32287
rect 46466 -32327 46954 -32321
rect 40358 -32695 40846 -32689
rect 40358 -32729 40370 -32695
rect 40834 -32729 40846 -32695
rect 40358 -32735 40846 -32729
rect 41376 -32695 41864 -32689
rect 41376 -32729 41388 -32695
rect 41852 -32729 41864 -32695
rect 41376 -32735 41864 -32729
rect 41582 -32736 41642 -32735
rect 40062 -32828 40076 -32788
rect 40070 -33304 40076 -32828
rect 39092 -33364 39106 -33332
rect 38322 -33423 38810 -33417
rect 38322 -33457 38334 -33423
rect 38798 -33457 38810 -33423
rect 38322 -33463 38810 -33457
rect 32866 -34078 32872 -34018
rect 32932 -34078 32938 -34018
rect 33428 -34078 33434 -34018
rect 33494 -34078 33500 -34018
rect 34470 -34078 34476 -34018
rect 34536 -34078 34542 -34018
rect 35470 -34078 35476 -34018
rect 35536 -34078 35542 -34018
rect 32872 -36660 32932 -34078
rect 37484 -34116 37544 -33578
rect 37992 -33514 38088 -33510
rect 37992 -33516 38024 -33514
rect 38084 -33574 38090 -33514
rect 38478 -33574 38484 -33514
rect 38544 -33574 38550 -33514
rect 37992 -34116 38052 -33576
rect 38484 -34116 38544 -33574
rect 38638 -34018 38698 -33463
rect 39042 -33766 39106 -33364
rect 40060 -33364 40076 -33304
rect 40110 -32828 40126 -32788
rect 41088 -32788 41134 -32776
rect 40110 -33304 40116 -32828
rect 40110 -33364 40120 -33304
rect 41088 -33328 41094 -32788
rect 39340 -33423 39828 -33417
rect 39340 -33457 39352 -33423
rect 39816 -33457 39828 -33423
rect 39340 -33463 39828 -33457
rect 39042 -33836 39106 -33830
rect 39528 -33512 39588 -33506
rect 38632 -34078 38638 -34018
rect 38698 -34078 38704 -34018
rect 39528 -34116 39588 -33572
rect 39648 -34018 39708 -33463
rect 40060 -33514 40120 -33364
rect 41078 -33364 41094 -33328
rect 41128 -33328 41134 -32788
rect 42098 -32788 42162 -32438
rect 42598 -32689 42658 -32438
rect 42394 -32695 42882 -32689
rect 42394 -32729 42406 -32695
rect 42870 -32729 42882 -32695
rect 42394 -32735 42882 -32729
rect 42098 -32840 42112 -32788
rect 42106 -33322 42112 -32840
rect 41128 -33364 41142 -33328
rect 40358 -33423 40846 -33417
rect 40358 -33457 40370 -33423
rect 40834 -33457 40846 -33423
rect 40358 -33463 40846 -33457
rect 40054 -33574 40060 -33514
rect 40120 -33574 40126 -33514
rect 40590 -34018 40650 -33463
rect 41078 -33908 41142 -33364
rect 42098 -33364 42112 -33322
rect 42146 -32840 42162 -32788
rect 43112 -32788 43172 -32438
rect 43636 -32689 43696 -32438
rect 43412 -32695 43900 -32689
rect 43412 -32729 43424 -32695
rect 43888 -32729 43900 -32695
rect 43412 -32735 43900 -32729
rect 42146 -33322 42152 -32840
rect 43112 -32842 43130 -32788
rect 43124 -32918 43130 -32842
rect 42146 -33324 42158 -33322
rect 42146 -33364 42162 -33324
rect 41376 -33423 41864 -33417
rect 41376 -33457 41388 -33423
rect 41852 -33457 41864 -33423
rect 41376 -33463 41864 -33457
rect 41572 -33512 41632 -33506
rect 42098 -33512 42162 -33364
rect 43116 -33364 43130 -32918
rect 43164 -32842 43172 -32788
rect 44134 -32788 44194 -32438
rect 45144 -32440 45150 -32380
rect 45210 -32440 45216 -32380
rect 45652 -32440 45658 -32380
rect 45718 -32440 45724 -32380
rect 46162 -32440 46168 -32380
rect 46228 -32440 46234 -32380
rect 44634 -32652 44640 -32592
rect 44700 -32652 44706 -32592
rect 45646 -32652 45652 -32592
rect 45712 -32652 45718 -32592
rect 44640 -32689 44700 -32652
rect 45652 -32689 45712 -32652
rect 44430 -32695 44918 -32689
rect 44430 -32729 44442 -32695
rect 44906 -32729 44918 -32695
rect 44430 -32735 44918 -32729
rect 45448 -32695 45936 -32689
rect 45448 -32729 45460 -32695
rect 45924 -32729 45936 -32695
rect 45448 -32735 45936 -32729
rect 44134 -32842 44148 -32788
rect 43164 -32918 43170 -32842
rect 43164 -33364 43176 -32918
rect 44142 -33334 44148 -32842
rect 42594 -33417 42654 -33408
rect 42394 -33423 42882 -33417
rect 42394 -33457 42406 -33423
rect 42870 -33457 42882 -33423
rect 42394 -33463 42882 -33457
rect 41072 -33972 41078 -33908
rect 41142 -33972 41148 -33908
rect 39642 -34078 39648 -34018
rect 39708 -34078 39714 -34018
rect 40584 -34078 40590 -34018
rect 40650 -34078 40656 -34018
rect 41572 -34116 41632 -33572
rect 42066 -33516 42162 -33512
rect 42066 -33518 42098 -33516
rect 42158 -33576 42164 -33516
rect 42594 -33522 42654 -33463
rect 43116 -33512 43176 -33364
rect 44134 -33364 44148 -33334
rect 44182 -32842 44194 -32788
rect 45160 -32788 45206 -32776
rect 44182 -33334 44188 -32842
rect 45160 -33330 45166 -32788
rect 44182 -33336 44194 -33334
rect 44182 -33364 44198 -33336
rect 43594 -33417 43654 -33414
rect 43412 -33423 43900 -33417
rect 43412 -33457 43424 -33423
rect 43888 -33457 43900 -33423
rect 43412 -33463 43900 -33457
rect 42066 -34116 42126 -33578
rect 42594 -34116 42654 -33582
rect 43082 -33518 43176 -33512
rect 43142 -33520 43176 -33518
rect 43082 -33580 43116 -33578
rect 43082 -33586 43176 -33580
rect 43594 -33522 43654 -33463
rect 44134 -33518 44198 -33364
rect 45150 -33364 45166 -33330
rect 45200 -33330 45206 -32788
rect 46168 -32788 46232 -32440
rect 46654 -32592 46714 -32327
rect 47190 -32476 47250 -32228
rect 48214 -32228 48220 -31686
rect 48254 -31686 48264 -31652
rect 48254 -32228 48260 -31686
rect 48214 -32240 48260 -32228
rect 47484 -32287 47972 -32281
rect 47484 -32321 47496 -32287
rect 47960 -32321 47972 -32287
rect 47484 -32327 47972 -32321
rect 47184 -32536 47190 -32476
rect 47250 -32536 47256 -32476
rect 47192 -32590 47252 -32588
rect 46648 -32652 46654 -32592
rect 46714 -32652 46720 -32592
rect 47192 -32650 48264 -32590
rect 46654 -32689 46714 -32652
rect 46466 -32695 46954 -32689
rect 46466 -32729 46478 -32695
rect 46942 -32729 46954 -32695
rect 46466 -32735 46954 -32729
rect 46654 -32738 46714 -32735
rect 46168 -32834 46184 -32788
rect 45200 -33364 45214 -33330
rect 46178 -33334 46184 -32834
rect 44430 -33423 44918 -33417
rect 44430 -33457 44442 -33423
rect 44906 -33457 44918 -33423
rect 44430 -33463 44918 -33457
rect 44128 -33578 44134 -33518
rect 44194 -33578 44200 -33518
rect 43082 -34116 43142 -33586
rect 43594 -34116 43654 -33582
rect 45150 -33624 45214 -33364
rect 46168 -33364 46184 -33334
rect 46218 -32834 46232 -32788
rect 47192 -32788 47252 -32650
rect 47696 -32689 47756 -32650
rect 47484 -32695 47972 -32689
rect 47484 -32729 47496 -32695
rect 47960 -32729 47972 -32695
rect 47484 -32735 47972 -32729
rect 47192 -32814 47202 -32788
rect 46218 -33334 46224 -32834
rect 47196 -33276 47202 -32814
rect 46218 -33336 46228 -33334
rect 46218 -33364 46232 -33336
rect 45448 -33423 45936 -33417
rect 45448 -33457 45460 -33423
rect 45924 -33457 45936 -33423
rect 45448 -33463 45936 -33457
rect 46168 -33518 46232 -33364
rect 47184 -33364 47202 -33276
rect 47236 -32814 47252 -32788
rect 48204 -32788 48264 -32650
rect 47236 -33276 47242 -32814
rect 48204 -32838 48220 -32788
rect 47236 -33364 47244 -33276
rect 46466 -33423 46954 -33417
rect 46466 -33457 46478 -33423
rect 46942 -33457 46954 -33423
rect 46466 -33463 46954 -33457
rect 46162 -33578 46168 -33518
rect 46228 -33578 46234 -33518
rect 45144 -33688 45150 -33624
rect 45214 -33688 45220 -33624
rect 47184 -33912 47244 -33364
rect 48214 -33364 48220 -32838
rect 48254 -32838 48264 -32788
rect 48254 -33364 48260 -32838
rect 48214 -33376 48260 -33364
rect 47484 -33423 47972 -33417
rect 47484 -33457 47496 -33423
rect 47960 -33457 47972 -33423
rect 47484 -33463 47972 -33457
rect 48440 -33756 48500 -31298
rect 48436 -33762 48500 -33756
rect 48436 -33832 48500 -33826
rect 47178 -33972 47184 -33912
rect 47244 -33972 47250 -33912
rect 35148 -34176 45388 -34116
rect 32980 -34280 32986 -34220
rect 33046 -34280 33052 -34220
rect 32986 -36194 33046 -34280
rect 33408 -34333 33896 -34327
rect 33408 -34367 33420 -34333
rect 33884 -34367 33896 -34333
rect 33408 -34373 33896 -34367
rect 34426 -34333 34914 -34327
rect 34426 -34367 34438 -34333
rect 34902 -34367 34914 -34333
rect 34426 -34373 34914 -34367
rect 33120 -34426 33166 -34414
rect 33120 -34972 33126 -34426
rect 33112 -35002 33126 -34972
rect 33160 -34972 33166 -34426
rect 34138 -34426 34184 -34414
rect 33160 -35002 33172 -34972
rect 34138 -34978 34144 -34426
rect 33112 -35154 33172 -35002
rect 34130 -35002 34144 -34978
rect 34178 -34978 34184 -34426
rect 35148 -34426 35208 -34176
rect 36158 -34280 36164 -34220
rect 36224 -34280 36230 -34220
rect 35444 -34333 35932 -34327
rect 35444 -34367 35456 -34333
rect 35920 -34367 35932 -34333
rect 35444 -34373 35932 -34367
rect 34178 -35002 34190 -34978
rect 33408 -35061 33896 -35055
rect 33408 -35095 33420 -35061
rect 33884 -35095 33896 -35061
rect 33408 -35101 33896 -35095
rect 33624 -35154 33684 -35101
rect 34130 -35154 34190 -35002
rect 35148 -35002 35162 -34426
rect 35196 -35002 35208 -34426
rect 36164 -34426 36224 -34280
rect 36462 -34333 36950 -34327
rect 36462 -34367 36474 -34333
rect 36938 -34367 36950 -34333
rect 36462 -34373 36950 -34367
rect 36164 -34490 36180 -34426
rect 34426 -35061 34914 -35055
rect 34426 -35095 34438 -35061
rect 34902 -35095 34914 -35061
rect 34426 -35101 34914 -35095
rect 33112 -35156 34190 -35154
rect 33112 -35214 34130 -35156
rect 34124 -35216 34130 -35214
rect 34190 -35216 34196 -35156
rect 34634 -35264 34694 -35101
rect 34628 -35324 34634 -35264
rect 34694 -35324 34700 -35264
rect 34634 -35359 34694 -35324
rect 33408 -35365 33896 -35359
rect 33408 -35399 33420 -35365
rect 33884 -35399 33896 -35365
rect 33408 -35405 33896 -35399
rect 34426 -35365 34914 -35359
rect 34426 -35399 34438 -35365
rect 34902 -35399 34914 -35365
rect 34426 -35405 34914 -35399
rect 33120 -35458 33166 -35446
rect 33120 -35978 33126 -35458
rect 33112 -36034 33126 -35978
rect 33160 -35978 33166 -35458
rect 34138 -35458 34184 -35446
rect 33160 -36034 33172 -35978
rect 34138 -36004 34144 -35458
rect 33112 -36194 33172 -36034
rect 34126 -36034 34144 -36004
rect 34178 -36004 34184 -35458
rect 35148 -35458 35208 -35002
rect 36174 -35002 36180 -34490
rect 36214 -34490 36224 -34426
rect 37186 -34426 37246 -34176
rect 37480 -34333 37968 -34327
rect 37480 -34367 37492 -34333
rect 37956 -34367 37968 -34333
rect 37480 -34373 37968 -34367
rect 38498 -34333 38986 -34327
rect 38498 -34367 38510 -34333
rect 38974 -34367 38986 -34333
rect 38498 -34373 38986 -34367
rect 36214 -35002 36220 -34490
rect 36174 -35014 36220 -35002
rect 37186 -35002 37198 -34426
rect 37232 -35002 37246 -34426
rect 38210 -34426 38256 -34414
rect 38210 -34938 38216 -34426
rect 35654 -35055 35714 -35049
rect 35444 -35061 35932 -35055
rect 35444 -35095 35456 -35061
rect 35920 -35095 35932 -35061
rect 35444 -35101 35932 -35095
rect 36462 -35061 36950 -35055
rect 36462 -35095 36474 -35061
rect 36938 -35095 36950 -35061
rect 36462 -35101 36950 -35095
rect 35654 -35258 35714 -35101
rect 36158 -35216 36164 -35156
rect 36224 -35216 36230 -35156
rect 35654 -35264 35716 -35258
rect 35654 -35324 35656 -35264
rect 35654 -35330 35716 -35324
rect 35654 -35359 35714 -35330
rect 35444 -35365 35932 -35359
rect 35444 -35399 35456 -35365
rect 35920 -35399 35932 -35365
rect 35444 -35405 35932 -35399
rect 34178 -36034 34186 -36004
rect 33408 -36093 33896 -36087
rect 33408 -36127 33420 -36093
rect 33884 -36127 33896 -36093
rect 33408 -36133 33896 -36127
rect 33614 -36194 33674 -36133
rect 34126 -36188 34186 -36034
rect 35148 -36034 35162 -35458
rect 35196 -36034 35208 -35458
rect 36164 -35458 36224 -35216
rect 36676 -35258 36736 -35101
rect 36674 -35264 36736 -35258
rect 36734 -35324 36736 -35264
rect 36674 -35330 36736 -35324
rect 36676 -35359 36736 -35330
rect 36462 -35365 36950 -35359
rect 36462 -35399 36474 -35365
rect 36938 -35399 36950 -35365
rect 36462 -35405 36950 -35399
rect 36676 -35412 36736 -35405
rect 36164 -35504 36180 -35458
rect 34426 -36093 34914 -36087
rect 34426 -36127 34438 -36093
rect 34902 -36127 34914 -36093
rect 34426 -36133 34914 -36127
rect 34120 -36194 34126 -36188
rect 32986 -36248 34126 -36194
rect 34186 -36248 34192 -36188
rect 32986 -36254 34192 -36248
rect 34632 -36322 34692 -36133
rect 34632 -36388 34692 -36382
rect 35148 -36530 35208 -36034
rect 36174 -36034 36180 -35504
rect 36214 -35504 36224 -35458
rect 37186 -35458 37246 -35002
rect 38206 -35002 38216 -34938
rect 38250 -34938 38256 -34426
rect 39224 -34426 39284 -34176
rect 40226 -34280 40232 -34220
rect 40292 -34280 40298 -34220
rect 39516 -34333 40004 -34327
rect 39516 -34367 39528 -34333
rect 39992 -34367 40004 -34333
rect 39516 -34373 40004 -34367
rect 38250 -35002 38266 -34938
rect 37480 -35061 37968 -35055
rect 37480 -35095 37492 -35061
rect 37956 -35095 37968 -35061
rect 37480 -35101 37968 -35095
rect 37696 -35258 37756 -35101
rect 38206 -35156 38266 -35002
rect 39224 -35002 39234 -34426
rect 39268 -35002 39284 -34426
rect 40232 -34426 40292 -34280
rect 40534 -34333 41022 -34327
rect 40534 -34367 40546 -34333
rect 41010 -34367 41022 -34333
rect 40534 -34373 41022 -34367
rect 40232 -34500 40252 -34426
rect 38712 -35055 38772 -35053
rect 38498 -35061 38986 -35055
rect 38498 -35095 38510 -35061
rect 38974 -35095 38986 -35061
rect 38498 -35101 38986 -35095
rect 38200 -35216 38206 -35156
rect 38266 -35216 38272 -35156
rect 37696 -35264 37758 -35258
rect 37696 -35324 37698 -35264
rect 37696 -35330 37758 -35324
rect 38712 -35264 38772 -35101
rect 37696 -35359 37756 -35330
rect 38712 -35359 38772 -35324
rect 37480 -35365 37968 -35359
rect 37480 -35399 37492 -35365
rect 37956 -35399 37968 -35365
rect 37480 -35405 37968 -35399
rect 38498 -35365 38986 -35359
rect 38498 -35399 38510 -35365
rect 38974 -35399 38986 -35365
rect 38498 -35405 38986 -35399
rect 36214 -36034 36220 -35504
rect 36174 -36046 36220 -36034
rect 37186 -36034 37198 -35458
rect 37232 -36034 37246 -35458
rect 38210 -35458 38256 -35446
rect 38210 -35968 38216 -35458
rect 35646 -36087 35706 -36084
rect 35444 -36093 35932 -36087
rect 35444 -36127 35456 -36093
rect 35920 -36127 35932 -36093
rect 35444 -36133 35932 -36127
rect 36462 -36093 36950 -36087
rect 36462 -36127 36474 -36093
rect 36938 -36127 36950 -36093
rect 36462 -36133 36950 -36127
rect 35646 -36326 35706 -36133
rect 36678 -36318 36738 -36133
rect 36678 -36384 36738 -36378
rect 35646 -36392 35706 -36386
rect 37186 -36530 37246 -36034
rect 38206 -36034 38216 -35968
rect 38250 -35968 38256 -35458
rect 39224 -35458 39284 -35002
rect 40246 -35002 40252 -34500
rect 40286 -35002 40292 -34426
rect 40246 -35014 40292 -35002
rect 41260 -34426 41320 -34176
rect 41552 -34333 42040 -34327
rect 41552 -34367 41564 -34333
rect 42028 -34367 42040 -34333
rect 41552 -34373 42040 -34367
rect 42570 -34333 43058 -34327
rect 42570 -34367 42582 -34333
rect 43046 -34367 43058 -34333
rect 42570 -34373 43058 -34367
rect 41260 -35002 41270 -34426
rect 41304 -35002 41320 -34426
rect 42282 -34426 42328 -34414
rect 42282 -34938 42288 -34426
rect 39516 -35061 40004 -35055
rect 39516 -35095 39528 -35061
rect 39992 -35095 40004 -35061
rect 39516 -35101 40004 -35095
rect 40534 -35061 41022 -35055
rect 40534 -35095 40546 -35061
rect 41010 -35095 41022 -35061
rect 40534 -35101 41022 -35095
rect 39728 -35258 39788 -35101
rect 40226 -35216 40232 -35156
rect 40292 -35216 40298 -35156
rect 39728 -35264 39790 -35258
rect 39728 -35324 39730 -35264
rect 39728 -35330 39790 -35324
rect 39728 -35359 39788 -35330
rect 39516 -35365 40004 -35359
rect 39516 -35399 39528 -35365
rect 39992 -35399 40004 -35365
rect 39516 -35405 40004 -35399
rect 38250 -36034 38266 -35968
rect 37480 -36093 37968 -36087
rect 37480 -36127 37492 -36093
rect 37956 -36127 37968 -36093
rect 37480 -36133 37968 -36127
rect 37676 -36318 37736 -36133
rect 38206 -36188 38266 -36034
rect 39224 -36034 39234 -35458
rect 39268 -36034 39284 -35458
rect 40232 -35458 40292 -35216
rect 40738 -35258 40798 -35101
rect 40738 -35264 40800 -35258
rect 40738 -35324 40740 -35264
rect 40738 -35330 40800 -35324
rect 40738 -35359 40798 -35330
rect 40534 -35365 41022 -35359
rect 40534 -35399 40546 -35365
rect 41010 -35399 41022 -35365
rect 40534 -35405 41022 -35399
rect 40232 -35520 40252 -35458
rect 40246 -35942 40252 -35520
rect 38720 -36087 38780 -36074
rect 38498 -36093 38986 -36087
rect 38498 -36127 38510 -36093
rect 38974 -36127 38986 -36093
rect 38498 -36133 38986 -36127
rect 38200 -36248 38206 -36188
rect 38266 -36248 38272 -36188
rect 37676 -36384 37736 -36378
rect 38720 -36318 38780 -36133
rect 38720 -36384 38780 -36378
rect 39224 -36530 39284 -36034
rect 40242 -36034 40252 -35942
rect 40286 -35942 40292 -35458
rect 41260 -35458 41320 -35002
rect 42274 -35002 42288 -34938
rect 42322 -34938 42328 -34426
rect 43290 -34426 43350 -34176
rect 44302 -34280 44308 -34220
rect 44368 -34280 44374 -34220
rect 43588 -34333 44076 -34327
rect 43588 -34367 43600 -34333
rect 44064 -34367 44076 -34333
rect 43588 -34373 44076 -34367
rect 43290 -34836 43306 -34426
rect 43300 -34930 43306 -34836
rect 42322 -35002 42334 -34938
rect 41760 -35055 41820 -35053
rect 41552 -35061 42040 -35055
rect 41552 -35095 41564 -35061
rect 42028 -35095 42040 -35061
rect 41552 -35101 42040 -35095
rect 41760 -35258 41820 -35101
rect 42274 -35156 42334 -35002
rect 43290 -35002 43306 -34930
rect 43340 -34836 43350 -34426
rect 44308 -34426 44368 -34280
rect 44606 -34333 45094 -34327
rect 44606 -34367 44618 -34333
rect 45082 -34367 45094 -34333
rect 44606 -34373 45094 -34367
rect 44308 -34490 44324 -34426
rect 43340 -34930 43346 -34836
rect 43340 -35002 43350 -34930
rect 42774 -35055 42834 -35053
rect 42570 -35061 43058 -35055
rect 42570 -35095 42582 -35061
rect 43046 -35095 43058 -35061
rect 42570 -35101 43058 -35095
rect 42268 -35216 42274 -35156
rect 42334 -35216 42340 -35156
rect 42774 -35258 42834 -35101
rect 41760 -35264 41822 -35258
rect 41760 -35324 41762 -35264
rect 41760 -35330 41822 -35324
rect 42774 -35264 42836 -35258
rect 42774 -35324 42776 -35264
rect 42774 -35330 42836 -35324
rect 41760 -35359 41820 -35330
rect 42774 -35359 42834 -35330
rect 41552 -35365 42040 -35359
rect 41552 -35399 41564 -35365
rect 42028 -35399 42040 -35365
rect 41552 -35405 42040 -35399
rect 42570 -35365 43058 -35359
rect 42570 -35399 42582 -35365
rect 43046 -35399 43058 -35365
rect 42570 -35405 43058 -35399
rect 40286 -36034 40302 -35942
rect 39724 -36087 39784 -36084
rect 39516 -36093 40004 -36087
rect 39516 -36127 39528 -36093
rect 39992 -36127 40004 -36093
rect 39516 -36133 40004 -36127
rect 39724 -36322 39784 -36133
rect 39724 -36388 39784 -36382
rect 40242 -36438 40302 -36034
rect 41260 -36034 41270 -35458
rect 41304 -36034 41320 -35458
rect 42282 -35458 42328 -35446
rect 42282 -35952 42288 -35458
rect 40740 -36087 40800 -36080
rect 40534 -36093 41022 -36087
rect 40534 -36127 40546 -36093
rect 41010 -36127 41022 -36093
rect 40534 -36133 41022 -36127
rect 40740 -36322 40800 -36133
rect 40740 -36388 40800 -36382
rect 40032 -36498 40302 -36438
rect 35148 -36590 39524 -36530
rect 39584 -36590 39590 -36530
rect 32872 -36720 37040 -36660
rect 32750 -36908 32756 -36848
rect 32816 -36908 32822 -36848
rect 33916 -36908 33922 -36848
rect 33982 -36908 33988 -36848
rect 32482 -37954 32488 -37894
rect 32548 -37954 32554 -37894
rect 32240 -39112 32246 -39052
rect 32306 -39112 32312 -39052
rect 32236 -39326 32242 -39266
rect 32302 -39326 32308 -39266
rect 32124 -40368 32130 -40308
rect 32190 -40368 32196 -40308
rect 26786 -41622 32056 -41562
rect 26726 -41628 26786 -41622
rect 11452 -42356 22722 -42100
rect 25816 -42220 25928 -41706
rect 27780 -41824 27840 -41818
rect 30132 -41822 30192 -41816
rect 27776 -41884 27780 -41824
rect 27840 -41882 30132 -41824
rect 32242 -41824 32302 -39326
rect 32488 -41566 32548 -37954
rect 32618 -38052 32624 -37992
rect 32684 -38052 32690 -37992
rect 32482 -41626 32488 -41566
rect 32548 -41626 32554 -41566
rect 32624 -41696 32684 -38052
rect 32756 -40516 32816 -36908
rect 33200 -36969 33688 -36963
rect 33200 -37003 33212 -36969
rect 33676 -37003 33688 -36969
rect 33200 -37009 33688 -37003
rect 32912 -37062 32958 -37050
rect 32912 -37602 32918 -37062
rect 32904 -37638 32918 -37602
rect 32952 -37602 32958 -37062
rect 33922 -37062 33982 -36908
rect 34218 -36969 34706 -36963
rect 34218 -37003 34230 -36969
rect 34694 -37003 34706 -36969
rect 34218 -37009 34706 -37003
rect 33922 -37088 33936 -37062
rect 32952 -37638 32964 -37602
rect 33930 -37614 33936 -37088
rect 32904 -37796 32964 -37638
rect 33920 -37638 33936 -37614
rect 33970 -37088 33982 -37062
rect 34938 -37062 34998 -36720
rect 35952 -36908 35958 -36848
rect 36018 -36908 36024 -36848
rect 35236 -36969 35724 -36963
rect 35236 -37003 35248 -36969
rect 35712 -37003 35724 -36969
rect 35236 -37009 35724 -37003
rect 33970 -37614 33976 -37088
rect 34938 -37108 34954 -37062
rect 34948 -37614 34954 -37108
rect 33970 -37638 33980 -37614
rect 33200 -37697 33688 -37691
rect 33200 -37731 33212 -37697
rect 33676 -37731 33688 -37697
rect 33200 -37737 33688 -37731
rect 33418 -37796 33478 -37737
rect 33920 -37796 33980 -37638
rect 34940 -37638 34954 -37614
rect 34988 -37108 34998 -37062
rect 35958 -37062 36018 -36908
rect 36460 -36912 36466 -36848
rect 36530 -36912 36536 -36848
rect 36466 -36963 36530 -36912
rect 36254 -36969 36742 -36963
rect 36254 -37003 36266 -36969
rect 36730 -37003 36742 -36969
rect 36254 -37009 36742 -37003
rect 35958 -37086 35972 -37062
rect 34988 -37614 34994 -37108
rect 34988 -37638 35000 -37614
rect 34218 -37697 34706 -37691
rect 34218 -37731 34230 -37697
rect 34694 -37731 34706 -37697
rect 34218 -37737 34706 -37731
rect 32904 -37856 33980 -37796
rect 34410 -38098 34470 -37737
rect 34940 -37796 35000 -37638
rect 35966 -37638 35972 -37086
rect 36006 -37086 36018 -37062
rect 36980 -37062 37040 -36720
rect 37484 -36963 37544 -36590
rect 37272 -36969 37760 -36963
rect 37272 -37003 37284 -36969
rect 37748 -37003 37760 -36969
rect 37272 -37009 37760 -37003
rect 36006 -37638 36012 -37086
rect 36980 -37116 36990 -37062
rect 36984 -37610 36990 -37116
rect 35966 -37650 36012 -37638
rect 36976 -37638 36990 -37610
rect 37024 -37116 37040 -37062
rect 37992 -37062 38052 -36590
rect 38484 -36963 38544 -36590
rect 39522 -36963 39582 -36590
rect 38290 -36969 38778 -36963
rect 38290 -37003 38302 -36969
rect 38766 -37003 38778 -36969
rect 38290 -37009 38778 -37003
rect 39308 -36969 39796 -36963
rect 39308 -37003 39320 -36969
rect 39784 -37003 39796 -36969
rect 39308 -37009 39796 -37003
rect 37024 -37610 37030 -37116
rect 37024 -37638 37036 -37610
rect 35236 -37697 35724 -37691
rect 35236 -37731 35248 -37697
rect 35712 -37731 35724 -37697
rect 35236 -37737 35724 -37731
rect 36254 -37697 36742 -37691
rect 36254 -37731 36266 -37697
rect 36730 -37731 36742 -37697
rect 36254 -37737 36742 -37731
rect 34934 -37856 34940 -37796
rect 35000 -37856 35006 -37796
rect 35448 -37850 35508 -37737
rect 36454 -37850 36514 -37737
rect 36976 -37796 37036 -37638
rect 37992 -37638 38008 -37062
rect 38042 -37638 38052 -37062
rect 39020 -37062 39066 -37050
rect 39020 -37614 39026 -37062
rect 37272 -37697 37760 -37691
rect 37272 -37731 37284 -37697
rect 37748 -37731 37760 -37697
rect 37272 -37737 37760 -37731
rect 37486 -37792 37546 -37737
rect 37992 -37792 38052 -37638
rect 39012 -37638 39026 -37614
rect 39060 -37614 39066 -37062
rect 40032 -37062 40092 -36498
rect 41260 -36530 41320 -36034
rect 42274 -36034 42288 -35952
rect 42322 -35952 42328 -35458
rect 43290 -35458 43350 -35002
rect 44318 -35002 44324 -34490
rect 44358 -34490 44368 -34426
rect 45328 -34426 45388 -34176
rect 47498 -34280 47504 -34220
rect 47564 -34280 47570 -34220
rect 45624 -34333 46112 -34327
rect 45624 -34367 45636 -34333
rect 46100 -34367 46112 -34333
rect 45624 -34373 46112 -34367
rect 46642 -34333 47130 -34327
rect 46642 -34367 46654 -34333
rect 47118 -34367 47130 -34333
rect 46642 -34373 47130 -34367
rect 44358 -35002 44364 -34490
rect 44318 -35014 44364 -35002
rect 45328 -35002 45342 -34426
rect 45376 -35002 45388 -34426
rect 46354 -34426 46400 -34414
rect 46354 -34926 46360 -34426
rect 43806 -35055 43866 -35053
rect 44816 -35055 44876 -35053
rect 43588 -35061 44076 -35055
rect 43588 -35095 43600 -35061
rect 44064 -35095 44076 -35061
rect 43588 -35101 44076 -35095
rect 44606 -35061 45094 -35055
rect 44606 -35095 44618 -35061
rect 45082 -35095 45094 -35061
rect 44606 -35101 45094 -35095
rect 43806 -35258 43866 -35101
rect 44304 -35216 44310 -35156
rect 44370 -35216 44376 -35156
rect 43806 -35264 43868 -35258
rect 43806 -35324 43808 -35264
rect 43806 -35330 43868 -35324
rect 43806 -35359 43866 -35330
rect 43588 -35365 44076 -35359
rect 43588 -35399 43600 -35365
rect 44064 -35399 44076 -35365
rect 43588 -35405 44076 -35399
rect 42322 -36034 42334 -35952
rect 41552 -36093 42040 -36087
rect 41552 -36127 41564 -36093
rect 42028 -36127 42040 -36093
rect 41552 -36133 42040 -36127
rect 41744 -36322 41804 -36133
rect 42274 -36188 42334 -36034
rect 43290 -36034 43306 -35458
rect 43340 -36034 43350 -35458
rect 44310 -35458 44370 -35216
rect 44816 -35258 44876 -35101
rect 44816 -35264 44878 -35258
rect 44816 -35324 44818 -35264
rect 44816 -35330 44878 -35324
rect 44816 -35359 44876 -35330
rect 44606 -35365 45094 -35359
rect 44606 -35399 44618 -35365
rect 45082 -35399 45094 -35365
rect 44606 -35405 45094 -35399
rect 44310 -35526 44324 -35458
rect 42570 -36093 43058 -36087
rect 42570 -36127 42582 -36093
rect 43046 -36127 43058 -36093
rect 42570 -36133 43058 -36127
rect 42268 -36248 42274 -36188
rect 42334 -36248 42340 -36188
rect 41744 -36388 41804 -36382
rect 42776 -36318 42836 -36133
rect 42776 -36384 42836 -36378
rect 40534 -36790 40540 -36726
rect 40604 -36790 40610 -36726
rect 40540 -36848 40604 -36790
rect 41260 -36820 41320 -36590
rect 43290 -36430 43350 -36034
rect 44318 -36034 44324 -35526
rect 44358 -35526 44370 -35458
rect 45328 -35458 45388 -35002
rect 46346 -35002 46360 -34926
rect 46394 -34926 46400 -34426
rect 47372 -34426 47418 -34414
rect 46394 -35002 46406 -34926
rect 47372 -34976 47378 -34426
rect 45624 -35061 46112 -35055
rect 45624 -35095 45636 -35061
rect 46100 -35095 46112 -35061
rect 45624 -35101 46112 -35095
rect 45838 -35258 45898 -35101
rect 46346 -35154 46406 -35002
rect 47362 -35002 47378 -34976
rect 47412 -34976 47418 -34426
rect 47412 -35002 47422 -34976
rect 46642 -35061 47130 -35055
rect 46642 -35095 46654 -35061
rect 47118 -35095 47130 -35061
rect 46642 -35101 47130 -35095
rect 46868 -35154 46928 -35101
rect 47362 -35154 47422 -35002
rect 46346 -35156 47422 -35154
rect 46340 -35216 46346 -35156
rect 46406 -35214 47422 -35156
rect 46406 -35216 46412 -35214
rect 45838 -35264 45900 -35258
rect 45838 -35324 45840 -35264
rect 45838 -35330 45900 -35324
rect 45838 -35359 45898 -35330
rect 45624 -35365 46112 -35359
rect 45624 -35399 45636 -35365
rect 46100 -35399 46112 -35365
rect 45624 -35405 46112 -35399
rect 46642 -35365 47130 -35359
rect 46642 -35399 46654 -35365
rect 47118 -35399 47130 -35365
rect 46642 -35405 47130 -35399
rect 44358 -36034 44364 -35526
rect 44318 -36046 44364 -36034
rect 45328 -36034 45342 -35458
rect 45376 -36034 45388 -35458
rect 46354 -35458 46400 -35446
rect 46354 -35958 46360 -35458
rect 43792 -36087 43852 -36084
rect 43588 -36093 44076 -36087
rect 43588 -36127 43600 -36093
rect 44064 -36127 44076 -36093
rect 43588 -36133 44076 -36127
rect 44606 -36093 45094 -36087
rect 44606 -36127 44618 -36093
rect 45082 -36127 45094 -36093
rect 44606 -36133 45094 -36127
rect 43792 -36322 43852 -36133
rect 43792 -36388 43852 -36382
rect 44820 -36322 44880 -36133
rect 44820 -36388 44880 -36382
rect 45328 -36430 45388 -36034
rect 46342 -36034 46360 -35958
rect 46394 -35958 46400 -35458
rect 47372 -35458 47418 -35446
rect 46394 -36034 46402 -35958
rect 47372 -35962 47378 -35458
rect 45840 -36087 45900 -36084
rect 45624 -36093 46112 -36087
rect 45624 -36127 45636 -36093
rect 46100 -36127 46112 -36093
rect 45624 -36133 46112 -36127
rect 45840 -36322 45900 -36133
rect 46342 -36184 46402 -36034
rect 47362 -36034 47378 -35962
rect 47412 -35962 47418 -35458
rect 47412 -36034 47422 -35962
rect 46642 -36093 47130 -36087
rect 46642 -36127 46654 -36093
rect 47118 -36127 47130 -36093
rect 46642 -36133 47130 -36127
rect 46830 -36184 46890 -36133
rect 47362 -36184 47422 -36034
rect 47504 -36184 47564 -34280
rect 46340 -36188 47564 -36184
rect 46336 -36248 46342 -36188
rect 46402 -36244 47564 -36188
rect 46402 -36248 46408 -36244
rect 48292 -36380 48298 -36320
rect 48358 -36380 48364 -36320
rect 45840 -36388 45900 -36382
rect 43290 -36490 45388 -36430
rect 43290 -36820 43350 -36490
rect 47152 -36606 47158 -36546
rect 47218 -36606 47224 -36546
rect 44598 -36790 44604 -36726
rect 44668 -36790 44674 -36726
rect 45622 -36790 45628 -36726
rect 45692 -36790 45698 -36726
rect 46634 -36790 46640 -36726
rect 46704 -36790 46710 -36726
rect 40536 -36912 40542 -36848
rect 40606 -36912 40612 -36848
rect 41260 -36880 43654 -36820
rect 44604 -36844 44668 -36790
rect 40540 -36963 40604 -36912
rect 41572 -36963 41632 -36880
rect 40326 -36969 40814 -36963
rect 40326 -37003 40338 -36969
rect 40802 -37003 40814 -36969
rect 40326 -37009 40814 -37003
rect 41344 -36969 41832 -36963
rect 41344 -37003 41356 -36969
rect 41820 -37003 41832 -36969
rect 41344 -37009 41832 -37003
rect 39060 -37638 39072 -37614
rect 38290 -37697 38778 -37691
rect 38290 -37731 38302 -37697
rect 38766 -37731 38778 -37697
rect 38290 -37737 38778 -37731
rect 38506 -37792 38566 -37737
rect 39012 -37792 39072 -37638
rect 40032 -37638 40044 -37062
rect 40078 -37638 40092 -37062
rect 41056 -37062 41102 -37050
rect 41056 -37560 41062 -37062
rect 39308 -37697 39796 -37691
rect 39308 -37731 39320 -37697
rect 39784 -37731 39796 -37697
rect 39308 -37737 39796 -37731
rect 39516 -37792 39576 -37737
rect 34940 -37992 35000 -37856
rect 35448 -37910 36514 -37850
rect 36970 -37856 36976 -37796
rect 37036 -37856 37042 -37796
rect 37312 -37854 37318 -37794
rect 37378 -37854 37384 -37794
rect 37486 -37852 39576 -37792
rect 40032 -37794 40092 -37638
rect 41050 -37638 41062 -37560
rect 41096 -37560 41102 -37062
rect 42066 -37062 42126 -36880
rect 42594 -36963 42654 -36880
rect 42362 -36969 42850 -36963
rect 42362 -37003 42374 -36969
rect 42838 -37003 42850 -36969
rect 42362 -37009 42850 -37003
rect 42594 -37010 42654 -37009
rect 41096 -37638 41110 -37560
rect 40326 -37697 40814 -37691
rect 40326 -37731 40338 -37697
rect 40802 -37731 40814 -37697
rect 40326 -37737 40814 -37731
rect 34934 -38052 34940 -37992
rect 35000 -38052 35006 -37992
rect 35448 -38098 35508 -37910
rect 35954 -38050 35960 -37990
rect 36020 -38050 36026 -37990
rect 33920 -38162 33926 -38102
rect 33986 -38162 33992 -38102
rect 34410 -38158 35508 -38098
rect 35960 -38102 36020 -38050
rect 33200 -38225 33688 -38219
rect 33200 -38259 33212 -38225
rect 33676 -38259 33688 -38225
rect 33200 -38265 33688 -38259
rect 32912 -38318 32958 -38306
rect 32912 -38858 32918 -38318
rect 32908 -38894 32918 -38858
rect 32952 -38858 32958 -38318
rect 33926 -38318 33986 -38162
rect 34410 -38219 34470 -38158
rect 35448 -38219 35508 -38158
rect 35954 -38162 35960 -38102
rect 36020 -38162 36026 -38102
rect 34218 -38225 34706 -38219
rect 34218 -38259 34230 -38225
rect 34694 -38259 34706 -38225
rect 34218 -38265 34706 -38259
rect 35236 -38225 35724 -38219
rect 35236 -38259 35248 -38225
rect 35712 -38259 35724 -38225
rect 35236 -38265 35724 -38259
rect 33926 -38344 33936 -38318
rect 32952 -38894 32968 -38858
rect 33930 -38870 33936 -38344
rect 32908 -39052 32968 -38894
rect 33924 -38894 33936 -38870
rect 33970 -38344 33986 -38318
rect 34948 -38318 34994 -38306
rect 33970 -38870 33976 -38344
rect 34948 -38868 34954 -38318
rect 33970 -38894 33984 -38870
rect 33200 -38953 33688 -38947
rect 33200 -38987 33212 -38953
rect 33676 -38987 33688 -38953
rect 33200 -38993 33688 -38987
rect 33422 -39052 33482 -38993
rect 33924 -39052 33984 -38894
rect 34942 -38894 34954 -38868
rect 34988 -38868 34994 -38318
rect 35960 -38318 36020 -38162
rect 36454 -38219 36514 -37910
rect 37318 -38108 37378 -37854
rect 36976 -38168 37378 -38108
rect 36254 -38225 36742 -38219
rect 36254 -38259 36266 -38225
rect 36730 -38259 36742 -38225
rect 36254 -38265 36742 -38259
rect 35960 -38340 35972 -38318
rect 34988 -38894 35002 -38868
rect 34404 -38947 34464 -38946
rect 34218 -38953 34706 -38947
rect 34218 -38987 34230 -38953
rect 34694 -38987 34706 -38953
rect 34218 -38993 34706 -38987
rect 32908 -39112 33984 -39052
rect 32908 -39266 32968 -39112
rect 32902 -39326 32908 -39266
rect 32968 -39326 32974 -39266
rect 32906 -39436 33982 -39376
rect 32906 -39574 32966 -39436
rect 33420 -39475 33480 -39436
rect 33200 -39481 33688 -39475
rect 33200 -39515 33212 -39481
rect 33676 -39515 33688 -39481
rect 33200 -39521 33688 -39515
rect 32906 -39608 32918 -39574
rect 32912 -40150 32918 -39608
rect 32952 -39608 32966 -39574
rect 33922 -39574 33982 -39436
rect 34404 -39475 34464 -38993
rect 34942 -39156 35002 -38894
rect 35966 -38894 35972 -38340
rect 36006 -38340 36020 -38318
rect 36976 -38318 37036 -38168
rect 37272 -38225 37760 -38219
rect 37272 -38259 37284 -38225
rect 37748 -38259 37760 -38225
rect 37272 -38265 37760 -38259
rect 36006 -38894 36012 -38340
rect 36976 -38376 36990 -38318
rect 36984 -38864 36990 -38376
rect 35966 -38906 36012 -38894
rect 36978 -38894 36990 -38864
rect 37024 -38376 37036 -38318
rect 37992 -38318 38052 -37852
rect 40026 -37854 40032 -37794
rect 40092 -37854 40098 -37794
rect 41050 -37990 41110 -37638
rect 42066 -37638 42080 -37062
rect 42114 -37638 42126 -37062
rect 41344 -37697 41832 -37691
rect 41344 -37731 41356 -37697
rect 41820 -37731 41832 -37697
rect 41344 -37737 41832 -37731
rect 41560 -37792 41620 -37737
rect 42066 -37792 42126 -37638
rect 43082 -37062 43142 -36880
rect 43594 -36963 43654 -36880
rect 44098 -36908 44104 -36848
rect 44164 -36908 44170 -36848
rect 43380 -36969 43868 -36963
rect 43380 -37003 43392 -36969
rect 43856 -37003 43868 -36969
rect 43380 -37009 43868 -37003
rect 43594 -37016 43654 -37009
rect 43082 -37638 43098 -37062
rect 43132 -37638 43142 -37062
rect 44104 -37062 44164 -36908
rect 44604 -36963 44668 -36908
rect 45628 -36963 45692 -36790
rect 46132 -36908 46138 -36848
rect 46198 -36908 46204 -36848
rect 44398 -36969 44886 -36963
rect 44398 -37003 44410 -36969
rect 44874 -37003 44886 -36969
rect 44398 -37009 44886 -37003
rect 45416 -36969 45904 -36963
rect 45416 -37003 45428 -36969
rect 45892 -37003 45904 -36969
rect 45416 -37009 45904 -37003
rect 44104 -37090 44116 -37062
rect 42362 -37697 42850 -37691
rect 42362 -37731 42374 -37697
rect 42838 -37731 42850 -37697
rect 42362 -37737 42850 -37731
rect 42586 -37792 42646 -37737
rect 43082 -37792 43142 -37638
rect 44110 -37638 44116 -37090
rect 44150 -37090 44164 -37062
rect 45128 -37062 45174 -37050
rect 44150 -37638 44156 -37090
rect 45128 -37614 45134 -37062
rect 44110 -37650 44156 -37638
rect 45120 -37638 45134 -37614
rect 45168 -37614 45174 -37062
rect 46138 -37062 46198 -36908
rect 46640 -36963 46704 -36790
rect 47158 -36844 47218 -36606
rect 47158 -36904 48234 -36844
rect 46434 -36969 46922 -36963
rect 46434 -37003 46446 -36969
rect 46910 -37003 46922 -36969
rect 46434 -37009 46922 -37003
rect 46138 -37086 46152 -37062
rect 45168 -37638 45180 -37614
rect 43380 -37697 43868 -37691
rect 43380 -37731 43392 -37697
rect 43856 -37731 43868 -37697
rect 43380 -37737 43868 -37731
rect 44398 -37697 44886 -37691
rect 44398 -37731 44410 -37697
rect 44874 -37731 44886 -37697
rect 44398 -37737 44886 -37731
rect 43598 -37792 43658 -37737
rect 41560 -37852 43658 -37792
rect 41044 -38050 41050 -37990
rect 41110 -38050 41116 -37990
rect 39010 -38164 39016 -38104
rect 39076 -38164 39082 -38104
rect 41044 -38164 41050 -38104
rect 41110 -38164 41116 -38104
rect 38290 -38225 38778 -38219
rect 38290 -38259 38302 -38225
rect 38766 -38259 38778 -38225
rect 38290 -38265 38778 -38259
rect 37992 -38362 38008 -38318
rect 37024 -38864 37030 -38376
rect 38002 -38864 38008 -38362
rect 37024 -38894 37038 -38864
rect 35442 -38947 35502 -38946
rect 36448 -38947 36508 -38946
rect 35236 -38953 35724 -38947
rect 35236 -38987 35248 -38953
rect 35712 -38987 35724 -38953
rect 35236 -38993 35724 -38987
rect 36254 -38953 36742 -38947
rect 36254 -38987 36266 -38953
rect 36730 -38987 36742 -38953
rect 36254 -38993 36742 -38987
rect 34942 -39222 35002 -39216
rect 34936 -39420 34942 -39360
rect 35002 -39420 35008 -39360
rect 34218 -39481 34706 -39475
rect 34218 -39515 34230 -39481
rect 34694 -39515 34706 -39481
rect 34218 -39521 34706 -39515
rect 33922 -39596 33936 -39574
rect 32952 -40150 32958 -39608
rect 33930 -40122 33936 -39596
rect 32912 -40162 32958 -40150
rect 33924 -40150 33936 -40122
rect 33970 -39596 33982 -39574
rect 34942 -39574 35002 -39420
rect 35442 -39475 35502 -38993
rect 36448 -39475 36508 -38993
rect 36978 -39156 37038 -38894
rect 37994 -38894 38008 -38864
rect 38042 -38362 38052 -38318
rect 39016 -38318 39076 -38164
rect 39308 -38225 39796 -38219
rect 39308 -38259 39320 -38225
rect 39784 -38259 39796 -38225
rect 39308 -38265 39796 -38259
rect 40326 -38225 40814 -38219
rect 40326 -38259 40338 -38225
rect 40802 -38259 40814 -38225
rect 40326 -38265 40814 -38259
rect 39016 -38346 39026 -38318
rect 38042 -38864 38048 -38362
rect 38042 -38894 38054 -38864
rect 37272 -38953 37760 -38947
rect 37272 -38987 37284 -38953
rect 37748 -38987 37760 -38953
rect 37272 -38993 37760 -38987
rect 37498 -39048 37558 -38993
rect 37994 -39048 38054 -38894
rect 39020 -38894 39026 -38346
rect 39060 -38346 39076 -38318
rect 40038 -38318 40084 -38306
rect 39060 -38894 39066 -38346
rect 40038 -38870 40044 -38318
rect 39020 -38906 39066 -38894
rect 40032 -38894 40044 -38870
rect 40078 -38870 40084 -38318
rect 41050 -38318 41110 -38164
rect 41344 -38225 41832 -38219
rect 41344 -38259 41356 -38225
rect 41820 -38259 41832 -38225
rect 41344 -38265 41832 -38259
rect 42362 -38225 42850 -38219
rect 42362 -38259 42374 -38225
rect 42838 -38259 42850 -38225
rect 42362 -38265 42850 -38259
rect 41050 -38348 41062 -38318
rect 41056 -38866 41062 -38348
rect 40078 -38894 40092 -38870
rect 38290 -38953 38778 -38947
rect 38290 -38987 38302 -38953
rect 38766 -38987 38778 -38953
rect 38290 -38993 38778 -38987
rect 39308 -38953 39796 -38947
rect 39308 -38987 39320 -38953
rect 39784 -38987 39796 -38953
rect 39308 -38993 39796 -38987
rect 38510 -39048 38570 -38993
rect 37498 -39108 38570 -39048
rect 36972 -39216 36978 -39156
rect 37038 -39216 37044 -39156
rect 36970 -39318 36976 -39258
rect 37036 -39318 37042 -39258
rect 36976 -39360 37036 -39318
rect 36970 -39420 36976 -39360
rect 37036 -39420 37042 -39360
rect 35236 -39481 35724 -39475
rect 35236 -39515 35248 -39481
rect 35712 -39515 35724 -39481
rect 35236 -39521 35724 -39515
rect 36254 -39481 36742 -39475
rect 36254 -39515 36266 -39481
rect 36730 -39515 36742 -39481
rect 36254 -39521 36742 -39515
rect 33970 -40122 33976 -39596
rect 34942 -39598 34954 -39574
rect 33970 -40150 33984 -40122
rect 33200 -40209 33688 -40203
rect 33200 -40243 33212 -40209
rect 33676 -40243 33688 -40209
rect 33200 -40249 33688 -40243
rect 33924 -40308 33984 -40150
rect 34948 -40150 34954 -39598
rect 34988 -39598 35002 -39574
rect 35966 -39574 36012 -39562
rect 34988 -40150 34994 -39598
rect 35966 -40126 35972 -39574
rect 34948 -40162 34994 -40150
rect 35960 -40150 35972 -40126
rect 36006 -40126 36012 -39574
rect 36976 -39574 37036 -39420
rect 37272 -39481 37760 -39475
rect 37272 -39515 37284 -39481
rect 37748 -39515 37760 -39481
rect 37272 -39521 37760 -39515
rect 36976 -39602 36990 -39574
rect 36006 -40150 36020 -40126
rect 36984 -40131 36990 -39602
rect 34416 -40203 34476 -40196
rect 35454 -40203 35514 -40196
rect 34218 -40209 34706 -40203
rect 34218 -40243 34230 -40209
rect 34694 -40243 34706 -40209
rect 34218 -40249 34706 -40243
rect 35236 -40209 35724 -40203
rect 35236 -40243 35248 -40209
rect 35712 -40243 35724 -40209
rect 35236 -40249 35724 -40243
rect 33918 -40368 33924 -40308
rect 33984 -40368 33990 -40308
rect 32750 -40576 32756 -40516
rect 32816 -40576 32822 -40516
rect 32906 -40674 33982 -40614
rect 32906 -40830 32966 -40674
rect 33420 -40731 33480 -40674
rect 33200 -40737 33688 -40731
rect 33200 -40771 33212 -40737
rect 33676 -40771 33688 -40737
rect 33200 -40777 33688 -40771
rect 32906 -40868 32918 -40830
rect 32912 -41406 32918 -40868
rect 32952 -40868 32966 -40830
rect 33922 -40830 33982 -40674
rect 34416 -40731 34476 -40249
rect 34932 -40678 34938 -40618
rect 34998 -40678 35004 -40618
rect 34218 -40737 34706 -40731
rect 34218 -40771 34230 -40737
rect 34694 -40771 34706 -40737
rect 34218 -40777 34706 -40771
rect 33922 -40856 33936 -40830
rect 32952 -41406 32958 -40868
rect 33930 -41380 33936 -40856
rect 32912 -41418 32958 -41406
rect 33920 -41406 33936 -41380
rect 33970 -40856 33982 -40830
rect 34938 -40830 34998 -40678
rect 35454 -40731 35514 -40249
rect 35960 -40308 36020 -40150
rect 36978 -40150 36990 -40131
rect 37024 -39602 37036 -39574
rect 37994 -39574 38054 -39108
rect 39006 -39112 39012 -39052
rect 39072 -39112 39078 -39052
rect 38290 -39481 38778 -39475
rect 38290 -39515 38302 -39481
rect 38766 -39515 38778 -39481
rect 38290 -39521 38778 -39515
rect 37024 -40131 37030 -39602
rect 37994 -39612 38008 -39574
rect 38002 -40116 38008 -39612
rect 37024 -40150 37038 -40131
rect 36460 -40203 36520 -40196
rect 36254 -40209 36742 -40203
rect 36254 -40243 36266 -40209
rect 36730 -40243 36742 -40209
rect 36254 -40249 36742 -40243
rect 35954 -40368 35960 -40308
rect 36020 -40368 36026 -40308
rect 35960 -40416 36020 -40368
rect 35954 -40476 35960 -40416
rect 36020 -40476 36026 -40416
rect 36460 -40466 36520 -40249
rect 36978 -40300 37038 -40150
rect 37992 -40150 38008 -40116
rect 38042 -39612 38054 -39574
rect 39012 -39574 39072 -39112
rect 39514 -39214 39574 -38993
rect 40032 -39052 40092 -38894
rect 41050 -38894 41062 -38866
rect 41096 -38348 41110 -38318
rect 42074 -38318 42120 -38306
rect 41096 -38866 41102 -38348
rect 42074 -38866 42080 -38318
rect 41096 -38894 41110 -38866
rect 40544 -38947 40604 -38940
rect 40326 -38953 40814 -38947
rect 40326 -38987 40338 -38953
rect 40802 -38987 40814 -38953
rect 40326 -38993 40814 -38987
rect 40026 -39112 40032 -39052
rect 40092 -39112 40098 -39052
rect 40544 -39214 40604 -38993
rect 39514 -39274 40604 -39214
rect 39514 -39475 39574 -39274
rect 40026 -39418 40032 -39358
rect 40092 -39418 40098 -39358
rect 39308 -39481 39796 -39475
rect 39308 -39515 39320 -39481
rect 39784 -39515 39796 -39481
rect 39308 -39521 39796 -39515
rect 39514 -39526 39574 -39521
rect 39012 -39598 39026 -39574
rect 38042 -40116 38048 -39612
rect 38042 -40150 38052 -40116
rect 39020 -40120 39026 -39598
rect 37272 -40209 37760 -40203
rect 37272 -40243 37284 -40209
rect 37748 -40243 37760 -40209
rect 37272 -40249 37760 -40243
rect 37496 -40300 37556 -40249
rect 37992 -40300 38052 -40150
rect 39014 -40150 39026 -40120
rect 39060 -39598 39072 -39574
rect 40032 -39574 40092 -39418
rect 40544 -39475 40604 -39274
rect 41050 -39358 41110 -38894
rect 42068 -38894 42080 -38866
rect 42114 -38866 42120 -38318
rect 43082 -38318 43142 -37852
rect 44100 -38164 44106 -38104
rect 44166 -38164 44172 -38104
rect 43380 -38225 43868 -38219
rect 43380 -38259 43392 -38225
rect 43856 -38259 43868 -38225
rect 43380 -38265 43868 -38259
rect 43082 -38338 43098 -38318
rect 43092 -38866 43098 -38338
rect 42114 -38894 42128 -38866
rect 41556 -38947 41616 -38940
rect 41344 -38953 41832 -38947
rect 41344 -38987 41356 -38953
rect 41820 -38987 41832 -38953
rect 41344 -38993 41832 -38987
rect 41044 -39418 41050 -39358
rect 41110 -39418 41116 -39358
rect 41556 -39475 41616 -38993
rect 42068 -39052 42128 -38894
rect 43082 -38894 43098 -38866
rect 43132 -38338 43142 -38318
rect 44106 -38318 44166 -38164
rect 44606 -38219 44666 -37737
rect 45120 -37796 45180 -37638
rect 46146 -37638 46152 -37086
rect 46186 -37086 46198 -37062
rect 47158 -37062 47218 -36904
rect 47672 -36963 47732 -36904
rect 47452 -36969 47940 -36963
rect 47452 -37003 47464 -36969
rect 47928 -37003 47940 -36969
rect 47452 -37009 47940 -37003
rect 46186 -37638 46192 -37086
rect 47158 -37098 47170 -37062
rect 47164 -37610 47170 -37098
rect 46146 -37650 46192 -37638
rect 47156 -37638 47170 -37610
rect 47204 -37098 47218 -37062
rect 48174 -37062 48234 -36904
rect 48174 -37086 48188 -37062
rect 47204 -37610 47210 -37098
rect 47204 -37638 47216 -37610
rect 46636 -37691 46696 -37685
rect 45416 -37697 45904 -37691
rect 45416 -37731 45428 -37697
rect 45892 -37731 45904 -37697
rect 45416 -37737 45904 -37731
rect 46434 -37697 46922 -37691
rect 46434 -37731 46446 -37697
rect 46910 -37731 46922 -37697
rect 46434 -37737 46922 -37731
rect 45114 -37856 45120 -37796
rect 45180 -37856 45186 -37796
rect 45630 -38219 45690 -37737
rect 46134 -38164 46140 -38104
rect 46200 -38164 46206 -38104
rect 44398 -38225 44886 -38219
rect 44398 -38259 44410 -38225
rect 44874 -38259 44886 -38225
rect 44398 -38265 44886 -38259
rect 45416 -38225 45904 -38219
rect 45416 -38259 45428 -38225
rect 45892 -38259 45904 -38225
rect 45416 -38265 45904 -38259
rect 43132 -38866 43138 -38338
rect 44106 -38346 44116 -38318
rect 43132 -38894 43142 -38866
rect 42362 -38953 42850 -38947
rect 42362 -38987 42374 -38953
rect 42838 -38987 42850 -38953
rect 42362 -38993 42850 -38987
rect 42586 -39050 42646 -38993
rect 43082 -39050 43142 -38894
rect 44110 -38894 44116 -38346
rect 44150 -38346 44166 -38318
rect 45128 -38318 45174 -38306
rect 44150 -38894 44156 -38346
rect 45128 -38858 45134 -38318
rect 44110 -38906 44156 -38894
rect 45118 -38894 45134 -38858
rect 45168 -38858 45174 -38318
rect 46140 -38318 46200 -38164
rect 46636 -38219 46696 -37737
rect 47156 -37796 47216 -37638
rect 48182 -37638 48188 -37086
rect 48222 -37086 48234 -37062
rect 48222 -37638 48228 -37086
rect 48182 -37650 48228 -37638
rect 47452 -37697 47940 -37691
rect 47452 -37731 47464 -37697
rect 47928 -37731 47940 -37697
rect 47452 -37737 47940 -37731
rect 47150 -37856 47156 -37796
rect 47216 -37856 47222 -37796
rect 47158 -38158 48234 -38098
rect 46434 -38225 46922 -38219
rect 46434 -38259 46446 -38225
rect 46910 -38259 46922 -38225
rect 46434 -38265 46922 -38259
rect 46140 -38342 46152 -38318
rect 45168 -38894 45178 -38858
rect 46146 -38866 46152 -38342
rect 44600 -38947 44660 -38946
rect 43380 -38953 43868 -38947
rect 43380 -38987 43392 -38953
rect 43856 -38987 43868 -38953
rect 43380 -38993 43868 -38987
rect 44398 -38953 44886 -38947
rect 44398 -38987 44410 -38953
rect 44874 -38987 44886 -38953
rect 44398 -38993 44886 -38987
rect 43598 -39050 43658 -38993
rect 42062 -39112 42068 -39052
rect 42128 -39112 42134 -39052
rect 42586 -39110 43658 -39050
rect 42060 -39418 42066 -39358
rect 42126 -39418 42132 -39358
rect 40326 -39481 40814 -39475
rect 40326 -39515 40338 -39481
rect 40802 -39515 40814 -39481
rect 40326 -39521 40814 -39515
rect 41344 -39481 41832 -39475
rect 41344 -39515 41356 -39481
rect 41820 -39515 41832 -39481
rect 41344 -39521 41832 -39515
rect 40032 -39596 40044 -39574
rect 39060 -40120 39066 -39598
rect 39060 -40150 39074 -40120
rect 38290 -40209 38778 -40203
rect 38290 -40243 38302 -40209
rect 38766 -40243 38778 -40209
rect 38290 -40249 38778 -40243
rect 38508 -40300 38568 -40249
rect 36972 -40360 36978 -40300
rect 37038 -40360 37044 -40300
rect 37496 -40360 38568 -40300
rect 38774 -40360 38780 -40300
rect 38840 -40360 38846 -40300
rect 39014 -40306 39074 -40150
rect 40038 -40150 40044 -39596
rect 40078 -39596 40092 -39574
rect 41056 -39574 41102 -39562
rect 40078 -40150 40084 -39596
rect 41056 -40124 41062 -39574
rect 40038 -40162 40084 -40150
rect 41050 -40150 41062 -40124
rect 41096 -40124 41102 -39574
rect 42066 -39574 42126 -39418
rect 42362 -39481 42850 -39475
rect 42362 -39515 42374 -39481
rect 42838 -39515 42850 -39481
rect 42362 -39521 42850 -39515
rect 42066 -39600 42080 -39574
rect 41096 -40150 41110 -40124
rect 39308 -40209 39796 -40203
rect 39308 -40243 39320 -40209
rect 39784 -40243 39796 -40209
rect 39308 -40249 39796 -40243
rect 40326 -40209 40814 -40203
rect 40326 -40243 40338 -40209
rect 40802 -40243 40814 -40209
rect 40326 -40249 40814 -40243
rect 36460 -40526 37236 -40466
rect 36460 -40731 36520 -40526
rect 36966 -40678 36972 -40618
rect 37032 -40678 37038 -40618
rect 37176 -40630 37236 -40526
rect 35236 -40737 35724 -40731
rect 35236 -40771 35248 -40737
rect 35712 -40771 35724 -40737
rect 35236 -40777 35724 -40771
rect 36254 -40737 36742 -40731
rect 36254 -40771 36266 -40737
rect 36730 -40771 36742 -40737
rect 36254 -40777 36742 -40771
rect 34938 -40856 34954 -40830
rect 33970 -41380 33976 -40856
rect 33970 -41406 33980 -41380
rect 33200 -41465 33688 -41459
rect 33200 -41499 33212 -41465
rect 33676 -41499 33688 -41465
rect 33200 -41505 33688 -41499
rect 33920 -41566 33980 -41406
rect 34948 -41406 34954 -40856
rect 34988 -40856 34998 -40830
rect 35966 -40830 36012 -40818
rect 34988 -41406 34994 -40856
rect 35966 -41384 35972 -40830
rect 34948 -41418 34994 -41406
rect 35956 -41406 35972 -41384
rect 36006 -41384 36012 -40830
rect 36972 -40830 37032 -40678
rect 37170 -40690 37176 -40630
rect 37236 -40690 37242 -40630
rect 37272 -40737 37760 -40731
rect 37272 -40771 37284 -40737
rect 37748 -40771 37760 -40737
rect 37272 -40777 37760 -40771
rect 36972 -40860 36990 -40830
rect 36984 -41370 36990 -40860
rect 36006 -41406 36016 -41384
rect 34218 -41465 34706 -41459
rect 34218 -41499 34230 -41465
rect 34694 -41499 34706 -41465
rect 34218 -41505 34706 -41499
rect 35236 -41465 35724 -41459
rect 35236 -41499 35248 -41465
rect 35712 -41499 35724 -41465
rect 35236 -41505 35724 -41499
rect 33914 -41626 33920 -41566
rect 33980 -41626 33986 -41566
rect 34428 -41680 34488 -41505
rect 35452 -41680 35512 -41505
rect 35956 -41566 36016 -41406
rect 36978 -41406 36990 -41370
rect 37024 -40860 37032 -40830
rect 37992 -40830 38052 -40360
rect 38780 -40570 38840 -40360
rect 39008 -40366 39014 -40306
rect 39074 -40366 39080 -40306
rect 39510 -40428 39570 -40249
rect 40538 -40428 40598 -40249
rect 41050 -40306 41110 -40150
rect 42074 -40150 42080 -39600
rect 42114 -39600 42126 -39574
rect 43082 -39574 43142 -39110
rect 44096 -39216 44102 -39156
rect 44162 -39216 44168 -39156
rect 43380 -39481 43868 -39475
rect 43380 -39515 43392 -39481
rect 43856 -39515 43868 -39481
rect 43380 -39521 43868 -39515
rect 42114 -40150 42120 -39600
rect 43082 -39604 43098 -39574
rect 43092 -40118 43098 -39604
rect 42074 -40162 42120 -40150
rect 43080 -40150 43098 -40118
rect 43132 -39604 43142 -39574
rect 44102 -39574 44162 -39216
rect 44600 -39475 44660 -38993
rect 44964 -39098 44970 -39038
rect 45030 -39098 45036 -39038
rect 44970 -39358 45030 -39098
rect 45118 -39148 45178 -38894
rect 46138 -38894 46152 -38866
rect 46186 -38342 46200 -38318
rect 47158 -38318 47218 -38158
rect 47672 -38219 47732 -38158
rect 47452 -38225 47940 -38219
rect 47452 -38259 47464 -38225
rect 47928 -38259 47940 -38225
rect 47452 -38265 47940 -38259
rect 46186 -38866 46192 -38342
rect 47158 -38352 47170 -38318
rect 47164 -38854 47170 -38352
rect 46186 -38894 46198 -38866
rect 45624 -38947 45684 -38946
rect 45416 -38953 45904 -38947
rect 45416 -38987 45428 -38953
rect 45892 -38987 45904 -38953
rect 45416 -38993 45904 -38987
rect 45112 -39208 45118 -39148
rect 45178 -39208 45184 -39148
rect 44964 -39418 44970 -39358
rect 45030 -39418 45036 -39358
rect 45116 -39416 45122 -39356
rect 45182 -39416 45188 -39356
rect 44398 -39481 44886 -39475
rect 44398 -39515 44410 -39481
rect 44874 -39515 44886 -39481
rect 44398 -39521 44886 -39515
rect 43132 -40118 43138 -39604
rect 44102 -39606 44116 -39574
rect 44110 -40118 44116 -39606
rect 43132 -40150 43140 -40118
rect 41344 -40209 41832 -40203
rect 41344 -40243 41356 -40209
rect 41820 -40243 41832 -40209
rect 41344 -40249 41832 -40243
rect 42362 -40209 42850 -40203
rect 42362 -40243 42374 -40209
rect 42838 -40243 42850 -40209
rect 42362 -40249 42850 -40243
rect 41044 -40366 41050 -40306
rect 41110 -40366 41116 -40306
rect 39510 -40488 40598 -40428
rect 41042 -40476 41048 -40416
rect 41108 -40476 41114 -40416
rect 38780 -40630 40088 -40570
rect 38290 -40737 38778 -40731
rect 38290 -40771 38302 -40737
rect 38766 -40771 38778 -40737
rect 38290 -40777 38778 -40771
rect 39308 -40737 39796 -40731
rect 39308 -40771 39320 -40737
rect 39784 -40771 39796 -40737
rect 39308 -40777 39796 -40771
rect 37024 -41370 37030 -40860
rect 37992 -40888 38008 -40830
rect 37024 -41406 37038 -41370
rect 38002 -41374 38008 -40888
rect 36254 -41465 36742 -41459
rect 36254 -41499 36266 -41465
rect 36730 -41499 36742 -41465
rect 36254 -41505 36742 -41499
rect 35950 -41626 35956 -41566
rect 36016 -41626 36022 -41566
rect 36458 -41680 36518 -41505
rect 32618 -41756 32624 -41696
rect 32684 -41756 32690 -41696
rect 34428 -41740 36518 -41680
rect 30192 -41882 32302 -41824
rect 27840 -41884 32302 -41882
rect 27780 -41890 27840 -41884
rect 30132 -41888 30192 -41884
rect 27660 -41942 27720 -41936
rect 32624 -41942 32684 -41756
rect 27720 -42002 32684 -41942
rect 27660 -42008 27720 -42002
rect 27214 -42060 27274 -42054
rect 34428 -42060 34488 -41740
rect 36458 -41950 36518 -41740
rect 36978 -41836 37038 -41406
rect 37992 -41406 38008 -41374
rect 38042 -40888 38052 -40830
rect 39020 -40830 39066 -40818
rect 38042 -41374 38048 -40888
rect 39020 -41362 39026 -40830
rect 38042 -41406 38052 -41374
rect 37272 -41465 37760 -41459
rect 37272 -41499 37284 -41465
rect 37748 -41499 37760 -41465
rect 37272 -41505 37760 -41499
rect 37496 -41560 37556 -41505
rect 37992 -41560 38052 -41406
rect 39014 -41406 39026 -41362
rect 39060 -41362 39066 -40830
rect 40028 -40830 40088 -40630
rect 40538 -40630 40598 -40488
rect 40538 -40731 40598 -40690
rect 40326 -40737 40814 -40731
rect 40326 -40771 40338 -40737
rect 40802 -40771 40814 -40737
rect 40326 -40777 40814 -40771
rect 40028 -40882 40044 -40830
rect 39060 -41406 39074 -41362
rect 38290 -41465 38778 -41459
rect 38290 -41499 38302 -41465
rect 38766 -41499 38778 -41465
rect 38290 -41505 38778 -41499
rect 38508 -41560 38568 -41505
rect 39014 -41560 39074 -41406
rect 40038 -41406 40044 -40882
rect 40078 -40882 40088 -40830
rect 41048 -40830 41108 -40476
rect 41554 -40630 41614 -40249
rect 42584 -40302 42644 -40249
rect 43080 -40302 43140 -40150
rect 44104 -40150 44116 -40118
rect 44150 -39606 44162 -39574
rect 45122 -39574 45182 -39416
rect 45624 -39475 45684 -38993
rect 46138 -39258 46198 -38894
rect 47158 -38894 47170 -38854
rect 47204 -38352 47218 -38318
rect 48174 -38318 48234 -38158
rect 48174 -38340 48188 -38318
rect 47204 -38854 47210 -38352
rect 47204 -38894 47218 -38854
rect 46630 -38947 46690 -38940
rect 46434 -38953 46922 -38947
rect 46434 -38987 46446 -38953
rect 46910 -38987 46922 -38953
rect 46434 -38993 46922 -38987
rect 46132 -39318 46138 -39258
rect 46198 -39318 46204 -39258
rect 46630 -39475 46690 -38993
rect 47158 -39148 47218 -38894
rect 48182 -38894 48188 -38340
rect 48222 -38340 48234 -38318
rect 48222 -38894 48228 -38340
rect 48182 -38906 48228 -38894
rect 47452 -38953 47940 -38947
rect 47452 -38987 47464 -38953
rect 47928 -38987 47940 -38953
rect 47452 -38993 47940 -38987
rect 48298 -39148 48358 -36380
rect 48440 -36548 48500 -33832
rect 48728 -36248 48734 -36188
rect 48794 -36248 48800 -36188
rect 48440 -36614 48500 -36608
rect 48576 -36908 48582 -36848
rect 48642 -36908 48648 -36848
rect 48416 -38050 48422 -37990
rect 48482 -38050 48488 -37990
rect 47152 -39208 47158 -39148
rect 47218 -39208 47224 -39148
rect 48292 -39208 48298 -39148
rect 48358 -39208 48364 -39148
rect 47150 -39416 47156 -39356
rect 47216 -39416 47222 -39356
rect 45416 -39481 45904 -39475
rect 45416 -39515 45428 -39481
rect 45892 -39515 45904 -39481
rect 45416 -39521 45904 -39515
rect 46434 -39481 46922 -39475
rect 46434 -39515 46446 -39481
rect 46910 -39515 46922 -39481
rect 46434 -39521 46922 -39515
rect 45122 -39594 45134 -39574
rect 44150 -40118 44156 -39606
rect 44150 -40150 44164 -40118
rect 43380 -40209 43868 -40203
rect 43380 -40243 43392 -40209
rect 43856 -40243 43868 -40209
rect 43380 -40249 43868 -40243
rect 43596 -40302 43656 -40249
rect 42584 -40362 43656 -40302
rect 44104 -40304 44164 -40150
rect 45128 -40150 45134 -39594
rect 45168 -39594 45182 -39574
rect 46146 -39574 46192 -39562
rect 45168 -40150 45174 -39594
rect 46146 -40122 46152 -39574
rect 45128 -40162 45174 -40150
rect 46140 -40150 46152 -40122
rect 46186 -40122 46192 -39574
rect 47156 -39574 47216 -39416
rect 47452 -39481 47940 -39475
rect 47452 -39515 47464 -39481
rect 47928 -39515 47940 -39481
rect 47452 -39521 47940 -39515
rect 47156 -39598 47170 -39574
rect 47164 -40114 47170 -39598
rect 46186 -40150 46200 -40122
rect 44612 -40203 44672 -40196
rect 45636 -40203 45696 -40196
rect 44398 -40209 44886 -40203
rect 44398 -40243 44410 -40209
rect 44874 -40243 44886 -40209
rect 44398 -40249 44886 -40243
rect 45416 -40209 45904 -40203
rect 45416 -40243 45428 -40209
rect 45892 -40243 45904 -40209
rect 45416 -40249 45904 -40243
rect 41554 -40696 41614 -40690
rect 41344 -40737 41832 -40731
rect 41344 -40771 41356 -40737
rect 41820 -40771 41832 -40737
rect 41344 -40777 41832 -40771
rect 42362 -40737 42850 -40731
rect 42362 -40771 42374 -40737
rect 42838 -40771 42850 -40737
rect 42362 -40777 42850 -40771
rect 40078 -41406 40084 -40882
rect 41048 -40894 41062 -40830
rect 40038 -41418 40084 -41406
rect 41056 -41406 41062 -40894
rect 41096 -40894 41108 -40830
rect 42074 -40830 42120 -40818
rect 41096 -41406 41102 -40894
rect 42074 -41378 42080 -40830
rect 41056 -41418 41102 -41406
rect 42066 -41406 42080 -41378
rect 42114 -41378 42120 -40830
rect 43080 -40830 43140 -40362
rect 44098 -40364 44104 -40304
rect 44164 -40364 44170 -40304
rect 44612 -40624 44672 -40249
rect 44612 -40630 44674 -40624
rect 44612 -40690 44614 -40630
rect 45120 -40678 45126 -40618
rect 45186 -40678 45192 -40618
rect 44612 -40696 44674 -40690
rect 44612 -40731 44672 -40696
rect 43380 -40737 43868 -40731
rect 43380 -40771 43392 -40737
rect 43856 -40771 43868 -40737
rect 43380 -40777 43868 -40771
rect 44398 -40737 44886 -40731
rect 44398 -40771 44410 -40737
rect 44874 -40771 44886 -40737
rect 44398 -40777 44886 -40771
rect 43080 -40868 43098 -40830
rect 43092 -41376 43098 -40868
rect 42114 -41406 42126 -41378
rect 39308 -41465 39796 -41459
rect 39308 -41499 39320 -41465
rect 39784 -41499 39796 -41465
rect 39308 -41505 39796 -41499
rect 40326 -41465 40814 -41459
rect 40326 -41499 40338 -41465
rect 40802 -41499 40814 -41465
rect 40326 -41505 40814 -41499
rect 41344 -41465 41832 -41459
rect 41344 -41499 41356 -41465
rect 41820 -41499 41832 -41465
rect 41344 -41505 41832 -41499
rect 39524 -41560 39584 -41505
rect 41550 -41560 41610 -41505
rect 42066 -41560 42126 -41406
rect 43080 -41406 43098 -41376
rect 43132 -40868 43140 -40830
rect 44110 -40830 44156 -40818
rect 43132 -41376 43138 -40868
rect 43132 -41406 43140 -41376
rect 44110 -41380 44116 -40830
rect 42362 -41465 42850 -41459
rect 42362 -41499 42374 -41465
rect 42838 -41499 42850 -41465
rect 42362 -41505 42850 -41499
rect 42584 -41560 42644 -41505
rect 43080 -41560 43140 -41406
rect 44108 -41406 44116 -41380
rect 44150 -41380 44156 -40830
rect 45126 -40830 45186 -40678
rect 45636 -40731 45696 -40249
rect 46140 -40304 46200 -40150
rect 47156 -40150 47170 -40114
rect 47204 -39598 47216 -39574
rect 48182 -39574 48228 -39562
rect 47204 -40114 47210 -39598
rect 47204 -40150 47216 -40114
rect 48182 -40126 48188 -39574
rect 46642 -40203 46702 -40190
rect 46434 -40209 46922 -40203
rect 46434 -40243 46446 -40209
rect 46910 -40243 46922 -40209
rect 46434 -40249 46922 -40243
rect 46134 -40364 46140 -40304
rect 46200 -40364 46206 -40304
rect 46642 -40731 46702 -40249
rect 47156 -40308 47216 -40150
rect 48172 -40150 48188 -40126
rect 48222 -40126 48228 -39574
rect 48222 -40150 48232 -40126
rect 47452 -40209 47940 -40203
rect 47452 -40243 47464 -40209
rect 47928 -40243 47940 -40209
rect 47452 -40249 47940 -40243
rect 47670 -40308 47730 -40249
rect 48172 -40308 48232 -40150
rect 47156 -40368 48232 -40308
rect 48298 -40416 48358 -39208
rect 48422 -39356 48482 -38050
rect 48416 -39416 48422 -39356
rect 48482 -39416 48488 -39356
rect 48292 -40476 48298 -40416
rect 48358 -40476 48364 -40416
rect 47154 -40678 47160 -40618
rect 47220 -40678 47226 -40618
rect 45416 -40737 45904 -40731
rect 45416 -40771 45428 -40737
rect 45892 -40771 45904 -40737
rect 45416 -40777 45904 -40771
rect 46434 -40737 46922 -40731
rect 46434 -40771 46446 -40737
rect 46910 -40771 46922 -40737
rect 46434 -40777 46922 -40771
rect 45126 -40856 45134 -40830
rect 44150 -41406 44168 -41380
rect 43380 -41465 43868 -41459
rect 43380 -41499 43392 -41465
rect 43856 -41499 43868 -41465
rect 43380 -41505 43868 -41499
rect 43596 -41560 43656 -41505
rect 37496 -41620 43656 -41560
rect 44108 -41566 44168 -41406
rect 45128 -41406 45134 -40856
rect 45168 -40856 45186 -40830
rect 46146 -40830 46192 -40818
rect 45168 -41406 45174 -40856
rect 46146 -41384 46152 -40830
rect 45128 -41418 45174 -41406
rect 46144 -41406 46152 -41384
rect 46186 -41384 46192 -40830
rect 47160 -40830 47220 -40678
rect 47452 -40737 47940 -40731
rect 47452 -40771 47464 -40737
rect 47928 -40771 47940 -40737
rect 47452 -40777 47940 -40771
rect 47160 -40860 47170 -40830
rect 47164 -41368 47170 -40860
rect 46186 -41406 46204 -41384
rect 44616 -41459 44676 -41452
rect 44398 -41465 44886 -41459
rect 44398 -41499 44410 -41465
rect 44874 -41499 44886 -41465
rect 44398 -41505 44886 -41499
rect 45416 -41465 45904 -41459
rect 45416 -41499 45428 -41465
rect 45892 -41499 45904 -41465
rect 45416 -41505 45904 -41499
rect 44102 -41626 44108 -41566
rect 44168 -41626 44174 -41566
rect 44616 -41678 44676 -41505
rect 45636 -41678 45696 -41505
rect 46144 -41566 46204 -41406
rect 47158 -41406 47170 -41368
rect 47204 -40860 47220 -40830
rect 48182 -40830 48228 -40818
rect 47204 -41368 47210 -40860
rect 47204 -41406 47218 -41368
rect 48182 -41380 48188 -40830
rect 46434 -41465 46922 -41459
rect 46434 -41499 46446 -41465
rect 46910 -41499 46922 -41465
rect 46434 -41505 46922 -41499
rect 46138 -41626 46144 -41566
rect 46204 -41626 46210 -41566
rect 46638 -41678 46698 -41505
rect 47158 -41562 47218 -41406
rect 48174 -41406 48188 -41380
rect 48222 -41380 48228 -40830
rect 48222 -41406 48234 -41380
rect 47452 -41465 47940 -41459
rect 47452 -41499 47464 -41465
rect 47928 -41499 47940 -41465
rect 47452 -41505 47940 -41499
rect 47672 -41562 47732 -41505
rect 48174 -41562 48234 -41406
rect 47158 -41622 48234 -41562
rect 44616 -41738 46698 -41678
rect 36972 -41896 36978 -41836
rect 37038 -41896 37044 -41836
rect 44616 -41950 44676 -41738
rect 48582 -41836 48642 -36908
rect 48734 -38104 48794 -36248
rect 48728 -38164 48734 -38104
rect 48794 -38164 48800 -38104
rect 50160 -41706 50166 -28276
rect 50266 -41706 50272 -28276
rect 48576 -41896 48582 -41836
rect 48642 -41896 48648 -41836
rect 36458 -42010 44676 -41950
rect 27274 -42120 34488 -42060
rect 27214 -42126 27274 -42120
rect 50160 -42220 50272 -41706
rect 25816 -42226 50272 -42220
rect 25816 -42326 25922 -42226
rect 50166 -42326 50272 -42226
rect 25816 -42332 50272 -42326
rect 52150 -38980 55526 -38974
rect 52150 -39080 52256 -38980
rect 55420 -39080 55526 -38980
rect 52150 -39086 55526 -39080
rect 52150 -39217 52262 -39086
rect 52150 -42087 52156 -39217
rect 52256 -39386 52262 -39217
rect 55130 -39386 55148 -39086
rect 52256 -39406 55148 -39386
rect 55414 -39217 55526 -39086
rect 52256 -42087 52262 -39406
rect 52312 -40260 52372 -39406
rect 52584 -39599 52792 -39593
rect 52584 -39633 52596 -39599
rect 52780 -39633 52792 -39599
rect 52584 -39639 52792 -39633
rect 53042 -39599 53250 -39593
rect 53042 -39633 53054 -39599
rect 53238 -39633 53250 -39599
rect 53042 -39639 53250 -39633
rect 52436 -39692 52482 -39680
rect 52436 -39848 52442 -39692
rect 52430 -39868 52442 -39848
rect 52476 -39848 52482 -39692
rect 52894 -39692 52940 -39680
rect 52894 -39826 52900 -39692
rect 52476 -39868 52490 -39848
rect 52430 -40134 52490 -39868
rect 52888 -39868 52900 -39826
rect 52934 -39826 52940 -39692
rect 53344 -39692 53404 -39406
rect 53500 -39599 53708 -39593
rect 53500 -39633 53512 -39599
rect 53696 -39633 53708 -39599
rect 53500 -39639 53708 -39633
rect 53958 -39599 54166 -39593
rect 53958 -39633 53970 -39599
rect 54154 -39633 54166 -39599
rect 53958 -39639 54166 -39633
rect 53344 -39728 53358 -39692
rect 52934 -39868 52948 -39826
rect 52584 -39927 52792 -39921
rect 52584 -39961 52596 -39927
rect 52780 -39961 52792 -39927
rect 52584 -39967 52792 -39961
rect 52658 -40134 52718 -39967
rect 52888 -40134 52948 -39868
rect 53352 -39868 53358 -39728
rect 53392 -39728 53404 -39692
rect 53810 -39692 53856 -39680
rect 53392 -39868 53398 -39728
rect 53810 -39834 53816 -39692
rect 53352 -39880 53398 -39868
rect 53802 -39868 53816 -39834
rect 53850 -39834 53856 -39692
rect 54258 -39692 54318 -39406
rect 54416 -39599 54624 -39593
rect 54416 -39633 54428 -39599
rect 54612 -39633 54624 -39599
rect 54416 -39639 54624 -39633
rect 54874 -39599 55082 -39593
rect 54874 -39633 54886 -39599
rect 55070 -39633 55082 -39599
rect 54874 -39639 55082 -39633
rect 54258 -39720 54274 -39692
rect 53850 -39868 53862 -39834
rect 53042 -39927 53250 -39921
rect 53042 -39961 53054 -39927
rect 53238 -39961 53250 -39927
rect 53042 -39967 53250 -39961
rect 53500 -39927 53708 -39921
rect 53500 -39961 53512 -39927
rect 53696 -39961 53708 -39927
rect 53500 -39967 53708 -39961
rect 53114 -40017 53174 -39967
rect 53570 -40017 53630 -39967
rect 53802 -40017 53862 -39868
rect 54268 -39868 54274 -39720
rect 54308 -39720 54318 -39692
rect 54726 -39692 54772 -39680
rect 54308 -39868 54314 -39720
rect 54726 -39833 54732 -39692
rect 54268 -39880 54314 -39868
rect 54716 -39868 54732 -39833
rect 54766 -39833 54772 -39692
rect 55184 -39692 55230 -39680
rect 55184 -39830 55190 -39692
rect 54766 -39868 54776 -39833
rect 53958 -39927 54166 -39921
rect 53958 -39961 53970 -39927
rect 54154 -39961 54166 -39927
rect 53958 -39967 54166 -39961
rect 54416 -39927 54624 -39921
rect 54416 -39961 54428 -39927
rect 54612 -39961 54624 -39927
rect 54416 -39967 54624 -39961
rect 54028 -40017 54088 -39967
rect 54492 -40017 54552 -39967
rect 53108 -40077 53114 -40017
rect 53174 -40077 54552 -40017
rect 54716 -40134 54776 -39868
rect 55174 -39868 55190 -39830
rect 55224 -39830 55230 -39692
rect 55224 -39868 55234 -39830
rect 54874 -39927 55082 -39921
rect 54874 -39961 54886 -39927
rect 55070 -39961 55082 -39927
rect 54874 -39967 55082 -39961
rect 54948 -40134 55008 -39967
rect 55174 -40134 55234 -39868
rect 52430 -40194 55234 -40134
rect 52312 -40320 52676 -40260
rect 52374 -40434 52380 -40374
rect 52440 -40434 52446 -40374
rect 52380 -41962 52440 -40434
rect 52488 -40575 52548 -40320
rect 52616 -40476 52676 -40320
rect 52593 -40482 52701 -40476
rect 52593 -40516 52605 -40482
rect 52689 -40516 52701 -40482
rect 52593 -40522 52701 -40516
rect 52851 -40482 52959 -40476
rect 52851 -40516 52863 -40482
rect 52947 -40516 52959 -40482
rect 52851 -40522 52959 -40516
rect 52488 -40592 52501 -40575
rect 52495 -40920 52501 -40592
rect 52492 -40951 52501 -40920
rect 52535 -40592 52548 -40575
rect 52753 -40575 52799 -40563
rect 52535 -40920 52541 -40592
rect 52535 -40951 52552 -40920
rect 52753 -40932 52759 -40575
rect 52492 -41162 52552 -40951
rect 52748 -40951 52759 -40932
rect 52793 -40932 52799 -40575
rect 53002 -40575 53062 -40194
rect 53258 -40316 53264 -40256
rect 53324 -40316 53330 -40256
rect 53128 -40434 53134 -40374
rect 53194 -40434 53200 -40374
rect 53134 -40476 53194 -40434
rect 53109 -40482 53217 -40476
rect 53109 -40516 53121 -40482
rect 53205 -40516 53217 -40482
rect 53109 -40522 53217 -40516
rect 52793 -40951 52808 -40932
rect 52593 -41010 52701 -41004
rect 52593 -41044 52605 -41010
rect 52689 -41044 52701 -41010
rect 52593 -41050 52701 -41044
rect 52616 -41162 52676 -41050
rect 52492 -41222 52676 -41162
rect 52492 -41435 52552 -41222
rect 52616 -41336 52676 -41222
rect 52748 -41226 52808 -40951
rect 53002 -40951 53017 -40575
rect 53051 -40951 53062 -40575
rect 53264 -40575 53324 -40316
rect 53386 -40434 53392 -40374
rect 53452 -40434 53458 -40374
rect 53392 -40476 53452 -40434
rect 53367 -40482 53475 -40476
rect 53367 -40516 53379 -40482
rect 53463 -40516 53475 -40482
rect 53367 -40522 53475 -40516
rect 53264 -40634 53275 -40575
rect 52851 -41010 52959 -41004
rect 52851 -41044 52863 -41010
rect 52947 -41044 52959 -41010
rect 52851 -41050 52959 -41044
rect 52878 -41106 52938 -41050
rect 52872 -41166 52878 -41106
rect 52938 -41166 52944 -41106
rect 52742 -41286 52748 -41226
rect 52808 -41286 52814 -41226
rect 52593 -41342 52701 -41336
rect 52593 -41376 52605 -41342
rect 52689 -41376 52701 -41342
rect 52593 -41382 52701 -41376
rect 52851 -41342 52959 -41336
rect 52851 -41376 52863 -41342
rect 52947 -41376 52959 -41342
rect 52851 -41382 52959 -41376
rect 52492 -41470 52501 -41435
rect 52495 -41762 52501 -41470
rect 52488 -41811 52501 -41762
rect 52535 -41470 52552 -41435
rect 52753 -41435 52799 -41423
rect 52535 -41762 52541 -41470
rect 52535 -41811 52548 -41762
rect 52753 -41780 52759 -41435
rect 52488 -41958 52548 -41811
rect 52748 -41811 52759 -41780
rect 52793 -41780 52799 -41435
rect 53002 -41435 53062 -40951
rect 53269 -40951 53275 -40634
rect 53309 -40634 53324 -40575
rect 53520 -40575 53580 -40194
rect 53625 -40482 53733 -40476
rect 53625 -40516 53637 -40482
rect 53721 -40516 53733 -40482
rect 53625 -40522 53733 -40516
rect 53883 -40482 53991 -40476
rect 53883 -40516 53895 -40482
rect 53979 -40516 53991 -40482
rect 53883 -40522 53991 -40516
rect 53309 -40951 53315 -40634
rect 53269 -40963 53315 -40951
rect 53520 -40951 53533 -40575
rect 53567 -40951 53580 -40575
rect 53785 -40575 53831 -40563
rect 53785 -40910 53791 -40575
rect 53109 -41010 53217 -41004
rect 53109 -41044 53121 -41010
rect 53205 -41044 53217 -41010
rect 53109 -41050 53217 -41044
rect 53367 -41010 53475 -41004
rect 53367 -41044 53379 -41010
rect 53463 -41044 53475 -41010
rect 53367 -41050 53475 -41044
rect 53126 -41166 53132 -41106
rect 53192 -41166 53198 -41106
rect 53386 -41166 53392 -41106
rect 53452 -41166 53458 -41106
rect 53132 -41336 53192 -41166
rect 53256 -41286 53262 -41226
rect 53322 -41286 53328 -41226
rect 53109 -41342 53217 -41336
rect 53109 -41376 53121 -41342
rect 53205 -41376 53217 -41342
rect 53109 -41382 53217 -41376
rect 53002 -41498 53017 -41435
rect 52793 -41811 52808 -41780
rect 52593 -41870 52701 -41864
rect 52593 -41904 52605 -41870
rect 52689 -41904 52701 -41870
rect 52593 -41910 52701 -41904
rect 52618 -41958 52678 -41910
rect 52374 -42022 52380 -41962
rect 52440 -42022 52446 -41962
rect 52488 -42018 52678 -41958
rect 52748 -41996 52808 -41811
rect 53011 -41811 53017 -41498
rect 53051 -41498 53062 -41435
rect 53262 -41435 53322 -41286
rect 53392 -41336 53452 -41166
rect 53367 -41342 53475 -41336
rect 53367 -41376 53379 -41342
rect 53463 -41376 53475 -41342
rect 53367 -41382 53475 -41376
rect 53262 -41472 53275 -41435
rect 53051 -41811 53057 -41498
rect 53011 -41823 53057 -41811
rect 53269 -41811 53275 -41472
rect 53309 -41472 53322 -41435
rect 53520 -41435 53580 -40951
rect 53778 -40951 53791 -40910
rect 53825 -40910 53831 -40575
rect 54036 -40575 54096 -40194
rect 54288 -40316 54294 -40256
rect 54354 -40316 54360 -40256
rect 54160 -40434 54166 -40374
rect 54226 -40434 54232 -40374
rect 54166 -40476 54226 -40434
rect 54141 -40482 54249 -40476
rect 54141 -40516 54153 -40482
rect 54237 -40516 54249 -40482
rect 54141 -40522 54249 -40516
rect 53825 -40951 53838 -40910
rect 53625 -41010 53733 -41004
rect 53625 -41044 53637 -41010
rect 53721 -41044 53733 -41010
rect 53625 -41050 53733 -41044
rect 53650 -41106 53710 -41050
rect 53644 -41166 53650 -41106
rect 53710 -41166 53716 -41106
rect 53778 -41226 53838 -40951
rect 54036 -40951 54049 -40575
rect 54083 -40951 54096 -40575
rect 54294 -40575 54354 -40316
rect 54420 -40434 54426 -40374
rect 54486 -40434 54492 -40374
rect 54426 -40476 54486 -40434
rect 54399 -40482 54507 -40476
rect 54399 -40516 54411 -40482
rect 54495 -40516 54507 -40482
rect 54399 -40522 54507 -40516
rect 54294 -40606 54307 -40575
rect 53883 -41010 53991 -41004
rect 53883 -41044 53895 -41010
rect 53979 -41044 53991 -41010
rect 53883 -41050 53991 -41044
rect 53908 -41106 53968 -41050
rect 53902 -41166 53908 -41106
rect 53968 -41166 53974 -41106
rect 53772 -41286 53778 -41226
rect 53838 -41286 53844 -41226
rect 53625 -41342 53733 -41336
rect 53625 -41376 53637 -41342
rect 53721 -41376 53733 -41342
rect 53625 -41382 53733 -41376
rect 53883 -41342 53991 -41336
rect 53883 -41376 53895 -41342
rect 53979 -41376 53991 -41342
rect 53883 -41382 53991 -41376
rect 53309 -41811 53315 -41472
rect 53520 -41486 53533 -41435
rect 53269 -41823 53315 -41811
rect 53527 -41811 53533 -41486
rect 53567 -41486 53580 -41435
rect 53785 -41435 53831 -41423
rect 53567 -41811 53573 -41486
rect 53785 -41762 53791 -41435
rect 53527 -41823 53573 -41811
rect 53778 -41811 53791 -41762
rect 53825 -41762 53831 -41435
rect 54036 -41435 54096 -40951
rect 54301 -40951 54307 -40606
rect 54341 -40606 54354 -40575
rect 54550 -40575 54610 -40194
rect 55180 -40316 55186 -40256
rect 55246 -40316 55252 -40256
rect 54940 -40434 55004 -40374
rect 55064 -40434 55128 -40374
rect 54940 -40476 55000 -40434
rect 54657 -40482 54765 -40476
rect 54657 -40516 54669 -40482
rect 54753 -40516 54765 -40482
rect 54657 -40522 54765 -40516
rect 54915 -40482 55023 -40476
rect 54915 -40516 54927 -40482
rect 55011 -40516 55023 -40482
rect 54915 -40522 55023 -40516
rect 54341 -40951 54347 -40606
rect 54301 -40963 54347 -40951
rect 54550 -40951 54565 -40575
rect 54599 -40951 54610 -40575
rect 54817 -40575 54863 -40563
rect 54817 -40886 54823 -40575
rect 54141 -41010 54249 -41004
rect 54141 -41044 54153 -41010
rect 54237 -41044 54249 -41010
rect 54141 -41050 54249 -41044
rect 54399 -41010 54507 -41004
rect 54399 -41044 54411 -41010
rect 54495 -41044 54507 -41010
rect 54399 -41050 54507 -41044
rect 54160 -41166 54166 -41106
rect 54226 -41166 54232 -41106
rect 54418 -41166 54424 -41106
rect 54484 -41166 54490 -41106
rect 54166 -41336 54226 -41166
rect 54288 -41286 54294 -41226
rect 54354 -41286 54360 -41226
rect 54141 -41342 54249 -41336
rect 54141 -41376 54153 -41342
rect 54237 -41376 54249 -41342
rect 54141 -41382 54249 -41376
rect 54036 -41496 54049 -41435
rect 53825 -41811 53838 -41762
rect 52851 -41870 52959 -41864
rect 52851 -41904 52863 -41870
rect 52947 -41904 52959 -41870
rect 52851 -41910 52959 -41904
rect 53109 -41870 53217 -41864
rect 53109 -41904 53121 -41870
rect 53205 -41904 53217 -41870
rect 53109 -41910 53217 -41904
rect 53367 -41870 53475 -41864
rect 53367 -41904 53379 -41870
rect 53463 -41904 53475 -41870
rect 53367 -41910 53475 -41904
rect 53625 -41870 53733 -41864
rect 53625 -41904 53637 -41870
rect 53721 -41904 53733 -41870
rect 53625 -41910 53733 -41904
rect 52874 -41962 52934 -41910
rect 53650 -41962 53710 -41910
rect 52746 -42078 52808 -41996
rect 52868 -42022 52874 -41962
rect 52934 -42022 52940 -41962
rect 53644 -42022 53650 -41962
rect 53710 -42022 53716 -41962
rect 52150 -42218 52262 -42087
rect 52740 -42138 52746 -42078
rect 52806 -42138 52812 -42078
rect 53778 -42080 53838 -41811
rect 54043 -41811 54049 -41496
rect 54083 -41496 54096 -41435
rect 54294 -41435 54354 -41286
rect 54424 -41336 54484 -41166
rect 54399 -41342 54507 -41336
rect 54399 -41376 54411 -41342
rect 54495 -41376 54507 -41342
rect 54399 -41382 54507 -41376
rect 54294 -41486 54307 -41435
rect 54083 -41811 54089 -41496
rect 54043 -41823 54089 -41811
rect 54301 -41811 54307 -41486
rect 54341 -41486 54354 -41435
rect 54550 -41435 54610 -40951
rect 54806 -40951 54823 -40886
rect 54857 -40886 54863 -40575
rect 55068 -40575 55128 -40434
rect 55068 -40618 55081 -40575
rect 54857 -40951 54866 -40886
rect 55075 -40906 55081 -40618
rect 54657 -41010 54765 -41004
rect 54657 -41044 54669 -41010
rect 54753 -41044 54765 -41010
rect 54657 -41050 54765 -41044
rect 54682 -41106 54742 -41050
rect 54676 -41166 54682 -41106
rect 54742 -41166 54748 -41106
rect 54806 -41226 54866 -40951
rect 55068 -40951 55081 -40906
rect 55115 -40618 55128 -40575
rect 55115 -40906 55121 -40618
rect 55115 -40951 55128 -40906
rect 54915 -41010 55023 -41004
rect 54915 -41044 54927 -41010
rect 55011 -41044 55023 -41010
rect 54915 -41050 55023 -41044
rect 54940 -41168 55000 -41050
rect 55068 -41168 55128 -40951
rect 54800 -41286 54806 -41226
rect 54866 -41286 54872 -41226
rect 54940 -41228 55128 -41168
rect 54940 -41336 55000 -41228
rect 54657 -41342 54765 -41336
rect 54657 -41376 54669 -41342
rect 54753 -41376 54765 -41342
rect 54657 -41382 54765 -41376
rect 54915 -41342 55023 -41336
rect 54915 -41376 54927 -41342
rect 55011 -41376 55023 -41342
rect 54915 -41382 55023 -41376
rect 54341 -41811 54347 -41486
rect 54550 -41496 54565 -41435
rect 54301 -41823 54347 -41811
rect 54559 -41811 54565 -41496
rect 54599 -41496 54610 -41435
rect 54817 -41435 54863 -41423
rect 54599 -41811 54605 -41496
rect 54817 -41768 54823 -41435
rect 54559 -41823 54605 -41811
rect 54808 -41811 54823 -41768
rect 54857 -41768 54863 -41435
rect 55068 -41435 55128 -41228
rect 55068 -41474 55081 -41435
rect 54857 -41811 54868 -41768
rect 55075 -41770 55081 -41474
rect 53883 -41870 53991 -41864
rect 53883 -41904 53895 -41870
rect 53979 -41904 53991 -41870
rect 53883 -41910 53991 -41904
rect 54141 -41870 54249 -41864
rect 54141 -41904 54153 -41870
rect 54237 -41904 54249 -41870
rect 54141 -41910 54249 -41904
rect 54399 -41870 54507 -41864
rect 54399 -41904 54411 -41870
rect 54495 -41904 54507 -41870
rect 54399 -41910 54507 -41904
rect 54657 -41870 54765 -41864
rect 54657 -41904 54669 -41870
rect 54753 -41904 54765 -41870
rect 54657 -41910 54765 -41904
rect 53906 -41962 53966 -41910
rect 54678 -41962 54738 -41910
rect 53900 -42022 53906 -41962
rect 53966 -42022 53972 -41962
rect 54672 -42022 54678 -41962
rect 54738 -42022 54744 -41962
rect 53778 -42146 53838 -42140
rect 54808 -42080 54868 -41811
rect 55066 -41811 55081 -41770
rect 55115 -41474 55128 -41435
rect 55115 -41770 55121 -41474
rect 55115 -41811 55126 -41770
rect 54915 -41870 55023 -41864
rect 54915 -41904 54927 -41870
rect 55011 -41904 55023 -41870
rect 54915 -41910 55023 -41904
rect 54940 -41960 55000 -41910
rect 55066 -41960 55126 -41811
rect 54940 -42020 55126 -41960
rect 54808 -42146 54868 -42140
rect 55186 -42080 55246 -40316
rect 55186 -42146 55246 -42140
rect 55414 -42087 55420 -39217
rect 55520 -42087 55526 -39217
rect 55852 -38980 58268 -38974
rect 55852 -39080 55958 -38980
rect 58162 -39080 58268 -38980
rect 55852 -39086 58268 -39080
rect 55852 -39172 55964 -39086
rect 55726 -40604 55732 -40544
rect 55792 -40604 55798 -40544
rect 55580 -41286 55586 -41226
rect 55646 -41286 55652 -41226
rect 55414 -42218 55526 -42087
rect 52150 -42224 55526 -42218
rect 52150 -42324 52256 -42224
rect 55420 -42324 55526 -42224
rect 52150 -42330 55526 -42324
rect 11452 -42648 11814 -42356
rect 22578 -42648 22722 -42356
rect 53908 -42428 53914 -42368
rect 53974 -42428 53980 -42368
rect 54090 -42384 55526 -42330
rect 54090 -42418 54200 -42384
rect 55424 -42418 55526 -42384
rect 11452 -42956 22722 -42648
rect 11452 -43150 23804 -42956
rect 53914 -43046 53974 -42428
rect 54090 -42432 55526 -42418
rect 54090 -42454 54148 -42432
rect 54090 -42922 54104 -42454
rect 54138 -42922 54148 -42454
rect 54200 -42476 54272 -42470
rect 54194 -42548 54200 -42476
rect 54260 -42482 54272 -42476
rect 54266 -42542 54272 -42482
rect 54260 -42548 54272 -42542
rect 54200 -42554 54272 -42548
rect 55283 -42471 55365 -42465
rect 55283 -42477 55295 -42471
rect 55283 -42547 55289 -42477
rect 55283 -42553 55295 -42547
rect 55365 -42553 55371 -42471
rect 55468 -42476 55526 -42432
rect 55283 -42559 55365 -42553
rect 54212 -42606 54258 -42594
rect 54212 -42756 54218 -42606
rect 54202 -42782 54218 -42756
rect 54252 -42756 54258 -42606
rect 54340 -42606 54386 -42594
rect 54340 -42736 54346 -42606
rect 54380 -42736 54386 -42606
rect 54468 -42606 54514 -42594
rect 54468 -42702 54474 -42606
rect 54252 -42782 54275 -42756
rect 54202 -42827 54275 -42782
rect 54326 -42796 54332 -42736
rect 54392 -42796 54398 -42736
rect 54462 -42782 54474 -42702
rect 54508 -42702 54514 -42606
rect 54596 -42606 54642 -42594
rect 54508 -42782 54522 -42702
rect 54596 -42726 54602 -42606
rect 54636 -42726 54642 -42606
rect 54724 -42606 54770 -42594
rect 54189 -42833 54286 -42827
rect 54189 -42906 54201 -42833
rect 54274 -42906 54286 -42833
rect 54462 -42844 54522 -42782
rect 54582 -42786 54588 -42726
rect 54648 -42786 54654 -42726
rect 54724 -42758 54730 -42606
rect 54716 -42782 54730 -42758
rect 54764 -42758 54770 -42606
rect 54852 -42606 54898 -42594
rect 54852 -42716 54858 -42606
rect 54892 -42716 54898 -42606
rect 54980 -42606 55026 -42594
rect 54764 -42782 54776 -42758
rect 54840 -42776 54846 -42716
rect 54906 -42776 54912 -42716
rect 54980 -42744 54986 -42606
rect 54596 -42794 54642 -42786
rect 54716 -42844 54776 -42782
rect 54852 -42782 54858 -42776
rect 54892 -42782 54898 -42776
rect 54852 -42794 54898 -42782
rect 54972 -42782 54986 -42744
rect 55020 -42744 55026 -42606
rect 55108 -42606 55154 -42594
rect 55108 -42718 55114 -42606
rect 55148 -42718 55154 -42606
rect 55236 -42606 55282 -42594
rect 55236 -42716 55242 -42606
rect 55276 -42716 55282 -42606
rect 55364 -42606 55410 -42594
rect 55020 -42782 55032 -42744
rect 55092 -42778 55098 -42718
rect 55158 -42778 55164 -42718
rect 55226 -42776 55232 -42716
rect 55292 -42776 55298 -42716
rect 55364 -42729 55370 -42606
rect 54972 -42844 55032 -42782
rect 55108 -42782 55114 -42778
rect 55148 -42782 55154 -42778
rect 55108 -42794 55154 -42782
rect 55228 -42782 55242 -42776
rect 55276 -42782 55288 -42776
rect 55228 -42844 55288 -42782
rect 55349 -42782 55370 -42729
rect 55404 -42729 55410 -42606
rect 55404 -42782 55424 -42729
rect 55349 -42826 55424 -42782
rect 54462 -42904 55288 -42844
rect 55336 -42832 55435 -42826
rect 54189 -42912 54286 -42906
rect 55336 -42907 55348 -42832
rect 55423 -42907 55435 -42832
rect 54090 -42949 54148 -42922
rect 54202 -42949 54275 -42912
rect 55336 -42913 55435 -42907
rect 55349 -42949 55424 -42913
rect 55468 -42922 55484 -42476
rect 55518 -42922 55526 -42476
rect 55468 -42949 55526 -42922
rect 54090 -42966 55526 -42949
rect 54090 -43000 54198 -42966
rect 55422 -43000 55526 -42966
rect 54090 -43008 55526 -43000
rect 55098 -43046 55158 -43040
rect 53914 -43048 54588 -43046
rect 53914 -43106 54332 -43048
rect 54326 -43108 54332 -43106
rect 54392 -43106 54588 -43048
rect 54648 -43106 54846 -43046
rect 54906 -43106 55098 -43046
rect 54392 -43108 54398 -43106
rect 55098 -43112 55158 -43106
rect 55586 -43066 55646 -41286
rect 55732 -41866 55792 -40604
rect 55852 -41338 55858 -39172
rect 55958 -41338 55964 -39172
rect 56516 -39386 56534 -39086
rect 58154 -39172 58268 -39086
rect 58154 -39386 58166 -39172
rect 56516 -39406 58166 -39386
rect 56568 -39556 56628 -39406
rect 56056 -39616 56628 -39556
rect 56056 -39892 56116 -39616
rect 56186 -39793 56246 -39616
rect 56312 -39726 56318 -39666
rect 56378 -39726 56384 -39666
rect 56162 -39799 56270 -39793
rect 56162 -39833 56174 -39799
rect 56258 -39833 56270 -39799
rect 56162 -39839 56270 -39833
rect 56056 -39946 56070 -39892
rect 56064 -40120 56070 -39946
rect 55852 -41424 55964 -41338
rect 56052 -40268 56070 -40120
rect 56104 -39946 56116 -39892
rect 56318 -39892 56378 -39726
rect 56420 -39799 56528 -39793
rect 56420 -39833 56432 -39799
rect 56516 -39833 56528 -39799
rect 56420 -39839 56528 -39833
rect 56318 -39932 56328 -39892
rect 56104 -40120 56110 -39946
rect 56104 -40268 56112 -40120
rect 56052 -40478 56112 -40268
rect 56322 -40268 56328 -39932
rect 56362 -39932 56378 -39892
rect 56568 -39892 56628 -39616
rect 56698 -39726 56704 -39666
rect 56764 -39726 56770 -39666
rect 56956 -39726 56962 -39666
rect 57022 -39726 57028 -39666
rect 56704 -39793 56764 -39726
rect 56962 -39793 57022 -39726
rect 56678 -39799 56786 -39793
rect 56678 -39833 56690 -39799
rect 56774 -39833 56786 -39799
rect 56678 -39839 56786 -39833
rect 56936 -39799 57044 -39793
rect 56936 -39833 56948 -39799
rect 57032 -39833 57044 -39799
rect 56936 -39839 57044 -39833
rect 56362 -40268 56368 -39932
rect 56322 -40280 56368 -40268
rect 56568 -40268 56586 -39892
rect 56620 -40268 56628 -39892
rect 56838 -39892 56884 -39880
rect 56838 -40224 56844 -39892
rect 56162 -40327 56270 -40321
rect 56162 -40361 56174 -40327
rect 56258 -40361 56270 -40327
rect 56162 -40367 56270 -40361
rect 56420 -40327 56528 -40321
rect 56420 -40361 56432 -40327
rect 56516 -40361 56528 -40327
rect 56420 -40367 56528 -40361
rect 56186 -40478 56246 -40367
rect 56052 -40538 56246 -40478
rect 56052 -40752 56112 -40538
rect 56186 -40653 56246 -40538
rect 56442 -40544 56502 -40367
rect 56312 -40604 56318 -40544
rect 56378 -40604 56384 -40544
rect 56436 -40604 56442 -40544
rect 56502 -40604 56508 -40544
rect 56162 -40659 56270 -40653
rect 56162 -40693 56174 -40659
rect 56258 -40693 56270 -40659
rect 56162 -40699 56270 -40693
rect 56052 -41128 56070 -40752
rect 56104 -41128 56112 -40752
rect 56318 -40752 56378 -40604
rect 56420 -40659 56528 -40653
rect 56420 -40693 56432 -40659
rect 56516 -40693 56528 -40659
rect 56420 -40699 56528 -40693
rect 56318 -40906 56328 -40752
rect 56052 -41282 56112 -41128
rect 56322 -41128 56328 -40906
rect 56362 -40906 56378 -40752
rect 56568 -40752 56628 -40268
rect 56832 -40268 56844 -40224
rect 56878 -40224 56884 -39892
rect 57084 -39892 57144 -39406
rect 57340 -39726 57346 -39666
rect 57406 -39726 57412 -39666
rect 57194 -39799 57302 -39793
rect 57194 -39833 57206 -39799
rect 57290 -39833 57302 -39799
rect 57194 -39839 57302 -39833
rect 56878 -40268 56892 -40224
rect 56678 -40327 56786 -40321
rect 56678 -40361 56690 -40327
rect 56774 -40361 56786 -40327
rect 56678 -40367 56786 -40361
rect 56832 -40544 56892 -40268
rect 57084 -40268 57102 -39892
rect 57136 -40268 57144 -39892
rect 57346 -39892 57406 -39726
rect 57452 -39799 57560 -39793
rect 57452 -39833 57464 -39799
rect 57548 -39833 57560 -39799
rect 57452 -39839 57560 -39833
rect 57346 -39924 57360 -39892
rect 56936 -40327 57044 -40321
rect 56936 -40361 56948 -40327
rect 57032 -40361 57044 -40327
rect 56936 -40367 57044 -40361
rect 56698 -40604 56704 -40544
rect 56764 -40604 56770 -40544
rect 56826 -40604 56832 -40544
rect 56892 -40604 56898 -40544
rect 56952 -40604 56958 -40544
rect 57018 -40604 57024 -40544
rect 56704 -40653 56764 -40604
rect 56958 -40653 57018 -40604
rect 56678 -40659 56786 -40653
rect 56678 -40693 56690 -40659
rect 56774 -40693 56786 -40659
rect 56678 -40699 56786 -40693
rect 56936 -40659 57044 -40653
rect 56936 -40693 56948 -40659
rect 57032 -40693 57044 -40659
rect 56936 -40699 57044 -40693
rect 56568 -40820 56586 -40752
rect 56362 -41128 56368 -40906
rect 56322 -41140 56368 -41128
rect 56580 -41128 56586 -40820
rect 56620 -40820 56628 -40752
rect 56838 -40752 56884 -40740
rect 56620 -41128 56626 -40820
rect 56838 -41082 56844 -40752
rect 56580 -41140 56626 -41128
rect 56828 -41128 56844 -41082
rect 56878 -41082 56884 -40752
rect 57084 -40752 57144 -40268
rect 57354 -40268 57360 -39924
rect 57394 -39924 57406 -39892
rect 57602 -39892 57662 -39406
rect 57710 -39799 57818 -39793
rect 57710 -39833 57722 -39799
rect 57806 -39833 57818 -39799
rect 57710 -39839 57818 -39833
rect 57394 -40268 57400 -39924
rect 57354 -40280 57400 -40268
rect 57602 -40268 57618 -39892
rect 57652 -40268 57662 -39892
rect 57194 -40327 57302 -40321
rect 57194 -40361 57206 -40327
rect 57290 -40361 57302 -40327
rect 57194 -40367 57302 -40361
rect 57452 -40327 57560 -40321
rect 57452 -40361 57464 -40327
rect 57548 -40361 57560 -40327
rect 57452 -40367 57560 -40361
rect 57216 -40544 57276 -40367
rect 57474 -40476 57534 -40367
rect 57602 -40472 57662 -40268
rect 57864 -39892 57924 -39406
rect 57980 -39726 57986 -39666
rect 58046 -39726 58052 -39666
rect 57864 -40268 57876 -39892
rect 57910 -40268 57924 -39892
rect 57710 -40327 57818 -40321
rect 57710 -40361 57722 -40327
rect 57806 -40361 57818 -40327
rect 57710 -40367 57818 -40361
rect 57738 -40472 57798 -40367
rect 57864 -40472 57924 -40268
rect 57468 -40536 57474 -40476
rect 57534 -40536 57540 -40476
rect 57602 -40532 57924 -40472
rect 57210 -40604 57216 -40544
rect 57276 -40604 57282 -40544
rect 57340 -40604 57346 -40544
rect 57406 -40604 57412 -40544
rect 57194 -40659 57302 -40653
rect 57194 -40693 57206 -40659
rect 57290 -40693 57302 -40659
rect 57194 -40699 57302 -40693
rect 57084 -40816 57102 -40752
rect 56878 -41128 56888 -41082
rect 56162 -41187 56270 -41181
rect 56162 -41221 56174 -41187
rect 56258 -41221 56270 -41187
rect 56162 -41227 56270 -41221
rect 56420 -41187 56528 -41181
rect 56420 -41221 56432 -41187
rect 56516 -41221 56528 -41187
rect 56420 -41227 56528 -41221
rect 56678 -41187 56786 -41181
rect 56678 -41221 56690 -41187
rect 56774 -41221 56786 -41187
rect 56678 -41227 56786 -41221
rect 56190 -41282 56250 -41227
rect 56052 -41342 56250 -41282
rect 56438 -41298 56498 -41227
rect 56828 -41298 56888 -41128
rect 57096 -41128 57102 -40816
rect 57136 -40816 57144 -40752
rect 57346 -40752 57406 -40604
rect 57474 -40653 57534 -40536
rect 57452 -40659 57560 -40653
rect 57452 -40693 57464 -40659
rect 57548 -40693 57560 -40659
rect 57452 -40699 57560 -40693
rect 57346 -40798 57360 -40752
rect 57136 -41128 57142 -40816
rect 57096 -41140 57142 -41128
rect 57354 -41128 57360 -40798
rect 57394 -40798 57406 -40752
rect 57602 -40752 57662 -40532
rect 57738 -40653 57798 -40532
rect 57710 -40659 57818 -40653
rect 57710 -40693 57722 -40659
rect 57806 -40693 57818 -40659
rect 57710 -40699 57818 -40693
rect 57602 -40798 57618 -40752
rect 57394 -41128 57400 -40798
rect 57354 -41140 57400 -41128
rect 57612 -41128 57618 -40798
rect 57652 -40798 57662 -40752
rect 57864 -40752 57924 -40532
rect 57864 -40794 57876 -40752
rect 57652 -41128 57658 -40798
rect 57612 -41140 57658 -41128
rect 57870 -41128 57876 -40794
rect 57910 -40794 57924 -40752
rect 57910 -41128 57916 -40794
rect 57870 -41140 57916 -41128
rect 56936 -41187 57044 -41181
rect 56936 -41221 56948 -41187
rect 57032 -41221 57044 -41187
rect 56936 -41227 57044 -41221
rect 57194 -41187 57302 -41181
rect 57194 -41221 57206 -41187
rect 57290 -41221 57302 -41187
rect 57194 -41227 57302 -41221
rect 57452 -41187 57560 -41181
rect 57452 -41221 57464 -41187
rect 57548 -41221 57560 -41187
rect 57452 -41227 57560 -41221
rect 57710 -41187 57818 -41181
rect 57710 -41221 57722 -41187
rect 57806 -41221 57818 -41187
rect 57710 -41227 57818 -41221
rect 57216 -41298 57276 -41227
rect 57986 -41298 58046 -39726
rect 56432 -41358 56438 -41298
rect 56498 -41358 56504 -41298
rect 56822 -41358 56828 -41298
rect 56888 -41358 56894 -41298
rect 57210 -41358 57216 -41298
rect 57276 -41358 57282 -41298
rect 57980 -41358 57986 -41298
rect 58046 -41358 58052 -41298
rect 58156 -41338 58162 -39406
rect 58262 -41338 58268 -39172
rect 58156 -41424 58268 -41338
rect 55852 -41430 58268 -41424
rect 55852 -41530 55958 -41430
rect 58162 -41530 58268 -41430
rect 55852 -41536 58268 -41530
rect 56104 -41574 57948 -41536
rect 56104 -41575 56958 -41574
rect 56104 -41609 56133 -41575
rect 56167 -41609 56225 -41575
rect 56259 -41609 56317 -41575
rect 56351 -41609 56409 -41575
rect 56443 -41609 56501 -41575
rect 56535 -41609 56593 -41575
rect 56627 -41609 56685 -41575
rect 56719 -41609 56777 -41575
rect 56811 -41609 56869 -41575
rect 56903 -41608 56958 -41575
rect 56992 -41608 57050 -41574
rect 57084 -41575 57948 -41574
rect 57084 -41608 57147 -41575
rect 56903 -41609 57147 -41608
rect 57181 -41609 57239 -41575
rect 57273 -41609 57331 -41575
rect 57365 -41609 57423 -41575
rect 57457 -41609 57515 -41575
rect 57549 -41609 57607 -41575
rect 57641 -41609 57699 -41575
rect 57733 -41609 57791 -41575
rect 57825 -41609 57883 -41575
rect 57917 -41609 57948 -41575
rect 56104 -41622 57948 -41609
rect 56104 -41640 57946 -41622
rect 58250 -41650 58256 -41590
rect 58316 -41650 58322 -41590
rect 56276 -41866 56336 -41860
rect 56436 -41866 56496 -41860
rect 55732 -41872 56230 -41866
rect 55732 -41920 56170 -41872
rect 56218 -41920 56230 -41872
rect 55732 -41926 56230 -41920
rect 56276 -41872 56496 -41866
rect 56276 -41920 56282 -41872
rect 56330 -41920 56442 -41872
rect 56490 -41920 56496 -41872
rect 56276 -41926 56496 -41920
rect 56538 -41872 56742 -41866
rect 56538 -41920 56550 -41872
rect 56598 -41920 56682 -41872
rect 56730 -41920 56742 -41872
rect 56538 -41926 56742 -41920
rect 56844 -41872 57090 -41866
rect 56844 -41920 56856 -41872
rect 56904 -41920 57090 -41872
rect 57324 -41868 57384 -41862
rect 57438 -41868 57498 -41862
rect 57554 -41866 57614 -41860
rect 57714 -41866 57774 -41860
rect 57324 -41874 57506 -41868
rect 56844 -41926 57090 -41920
rect 55732 -42958 55792 -41926
rect 56276 -41932 56336 -41926
rect 56436 -41932 56496 -41926
rect 56856 -41984 56916 -41978
rect 57030 -41984 57090 -41926
rect 57130 -41934 57136 -41874
rect 57196 -41934 57202 -41874
rect 57324 -41922 57330 -41874
rect 57378 -41922 57444 -41874
rect 57492 -41922 57506 -41874
rect 57324 -41928 57506 -41922
rect 57554 -41872 57774 -41866
rect 57554 -41920 57560 -41872
rect 57608 -41920 57720 -41872
rect 57768 -41920 57774 -41872
rect 57554 -41926 57774 -41920
rect 57324 -41934 57384 -41928
rect 57438 -41934 57498 -41928
rect 57554 -41932 57614 -41926
rect 57714 -41932 57774 -41926
rect 57826 -41866 57886 -41860
rect 58256 -41866 58316 -41650
rect 57826 -41872 58316 -41866
rect 57826 -41920 57832 -41872
rect 57880 -41920 58316 -41872
rect 57826 -41926 58316 -41920
rect 57826 -41932 57886 -41926
rect 57134 -41984 57196 -41978
rect 56850 -42044 56856 -41984
rect 56916 -42044 56922 -41984
rect 57030 -42044 57134 -41984
rect 57194 -42044 57196 -41984
rect 56856 -42050 56916 -42044
rect 57134 -42050 57196 -42044
rect 56104 -42118 57946 -42088
rect 56104 -42119 57050 -42118
rect 56104 -42153 56133 -42119
rect 56167 -42153 56225 -42119
rect 56259 -42153 56317 -42119
rect 56351 -42153 56409 -42119
rect 56443 -42153 56501 -42119
rect 56535 -42153 56593 -42119
rect 56627 -42153 56685 -42119
rect 56719 -42153 56777 -42119
rect 56811 -42153 56869 -42119
rect 56903 -42120 57050 -42119
rect 56903 -42153 56958 -42120
rect 56104 -42154 56958 -42153
rect 56992 -42152 57050 -42120
rect 57084 -42119 57946 -42118
rect 57084 -42152 57147 -42119
rect 56992 -42153 57147 -42152
rect 57181 -42153 57239 -42119
rect 57273 -42153 57331 -42119
rect 57365 -42153 57423 -42119
rect 57457 -42153 57515 -42119
rect 57549 -42153 57607 -42119
rect 57641 -42153 57699 -42119
rect 57733 -42153 57791 -42119
rect 57825 -42153 57883 -42119
rect 57917 -42153 57946 -42119
rect 56992 -42154 57946 -42153
rect 56104 -42184 57946 -42154
rect 56364 -42346 57734 -42184
rect 56364 -42446 56470 -42346
rect 57628 -42446 57734 -42346
rect 56364 -42452 57734 -42446
rect 56364 -42487 56476 -42452
rect 55890 -42624 55950 -42610
rect 55890 -42918 55902 -42624
rect 55936 -42918 55950 -42624
rect 56036 -42672 56042 -42572
rect 56142 -42672 56148 -42572
rect 56234 -42624 56298 -42612
rect 56010 -42714 56056 -42702
rect 56128 -42704 56174 -42702
rect 56010 -42734 56016 -42714
rect 55726 -43018 55732 -42958
rect 55792 -43018 55798 -42958
rect 55586 -43132 55646 -43126
rect 11452 -43156 50372 -43150
rect 11452 -43256 13222 -43156
rect 50266 -43256 50372 -43156
rect 55890 -43252 55950 -42918
rect 56004 -42890 56016 -42734
rect 56050 -42734 56056 -42714
rect 56120 -42714 56180 -42704
rect 56050 -42890 56064 -42734
rect 56004 -42958 56064 -42890
rect 56120 -42890 56134 -42714
rect 56168 -42764 56180 -42714
rect 56168 -42890 56182 -42764
rect 56120 -42896 56182 -42890
rect 56120 -42958 56180 -42896
rect 56234 -42918 56248 -42624
rect 56282 -42918 56298 -42624
rect 55998 -43018 56004 -42958
rect 56064 -43018 56070 -42958
rect 56114 -43018 56120 -42958
rect 56180 -43018 56186 -42958
rect 56234 -43252 56298 -42918
rect 56364 -43252 56370 -42487
rect 11452 -43262 50372 -43256
rect 11452 -43278 23802 -43262
rect 13116 -44048 13228 -43278
rect 27332 -43336 27392 -43330
rect 27654 -43386 27660 -43326
rect 27720 -43386 27726 -43326
rect 27780 -43334 27840 -43328
rect 26720 -43532 26726 -43472
rect 26786 -43532 26792 -43472
rect 26840 -43530 26846 -43470
rect 26906 -43530 26912 -43470
rect 26980 -43512 26986 -43452
rect 27046 -43512 27052 -43452
rect 27208 -43496 27214 -43436
rect 27274 -43496 27280 -43436
rect 26588 -43660 26594 -43600
rect 26654 -43660 26660 -43600
rect 10528 -56672 11876 -56612
rect 9350 -56724 9452 -56700
rect 9350 -57518 9372 -56724
rect 9436 -56726 10454 -56724
rect 10528 -56726 10588 -56672
rect 9436 -56738 10588 -56726
rect 9436 -56772 10342 -56738
rect 10562 -56772 10588 -56738
rect 9436 -56784 10588 -56772
rect 9436 -57094 9452 -56784
rect 10284 -56786 10588 -56784
rect 10284 -56836 10344 -56786
rect 10284 -57094 10294 -56836
rect 9436 -57154 10294 -57094
rect 9436 -57458 9452 -57154
rect 10284 -57408 10294 -57154
rect 10332 -57094 10344 -56836
rect 10394 -56934 10454 -56786
rect 10528 -56835 10588 -56786
rect 10784 -56720 10844 -56719
rect 11560 -56720 11620 -56714
rect 10784 -56780 11560 -56720
rect 10784 -56835 10844 -56780
rect 11042 -56835 11102 -56780
rect 11300 -56835 11360 -56780
rect 11560 -56835 11620 -56780
rect 11816 -56722 11876 -56672
rect 11816 -56738 12118 -56722
rect 11816 -56772 11834 -56738
rect 12036 -56772 12118 -56738
rect 11816 -56786 12118 -56772
rect 11816 -56835 11876 -56786
rect 10502 -56841 10610 -56835
rect 10502 -56875 10514 -56841
rect 10598 -56875 10610 -56841
rect 10502 -56881 10610 -56875
rect 10760 -56841 10868 -56835
rect 10760 -56875 10772 -56841
rect 10856 -56875 10868 -56841
rect 10760 -56881 10868 -56875
rect 11018 -56841 11126 -56835
rect 11018 -56875 11030 -56841
rect 11114 -56875 11126 -56841
rect 11018 -56881 11126 -56875
rect 11276 -56841 11384 -56835
rect 11276 -56875 11288 -56841
rect 11372 -56875 11384 -56841
rect 11276 -56881 11384 -56875
rect 11534 -56841 11642 -56835
rect 11534 -56875 11546 -56841
rect 11630 -56875 11642 -56841
rect 11534 -56881 11642 -56875
rect 11792 -56841 11900 -56835
rect 11792 -56875 11804 -56841
rect 11888 -56875 11900 -56841
rect 11792 -56881 11900 -56875
rect 10394 -57094 10410 -56934
rect 10332 -57154 10410 -57094
rect 10332 -57408 10344 -57154
rect 10404 -57276 10410 -57154
rect 10284 -57458 10344 -57408
rect 10396 -57310 10410 -57276
rect 10444 -57154 10454 -56934
rect 10662 -56934 10708 -56922
rect 10444 -57276 10450 -57154
rect 10662 -57265 10668 -56934
rect 10444 -57310 10456 -57276
rect 10396 -57458 10456 -57310
rect 10654 -57310 10668 -57265
rect 10702 -57265 10708 -56934
rect 10920 -56934 10966 -56922
rect 10702 -57310 10714 -57265
rect 10920 -57290 10926 -56934
rect 10502 -57369 10610 -57363
rect 10502 -57403 10514 -57369
rect 10598 -57403 10610 -57369
rect 10502 -57409 10610 -57403
rect 10524 -57458 10584 -57409
rect 9436 -57472 10584 -57458
rect 9436 -57506 10342 -57472
rect 10562 -57506 10584 -57472
rect 9436 -57518 10584 -57506
rect 9350 -57536 9452 -57518
rect 10654 -57635 10714 -57310
rect 10912 -57310 10926 -57290
rect 10960 -57290 10966 -56934
rect 11178 -56934 11224 -56922
rect 11178 -57267 11184 -56934
rect 10960 -57310 10972 -57290
rect 10760 -57369 10868 -57363
rect 10760 -57403 10772 -57369
rect 10856 -57403 10868 -57369
rect 10760 -57409 10868 -57403
rect 10912 -57486 10972 -57310
rect 11170 -57310 11184 -57267
rect 11218 -57267 11224 -56934
rect 11436 -56934 11482 -56922
rect 11218 -57310 11230 -57267
rect 11436 -57272 11442 -56934
rect 11018 -57369 11126 -57363
rect 11018 -57403 11030 -57369
rect 11114 -57403 11126 -57369
rect 11018 -57409 11126 -57403
rect 10906 -57546 10912 -57486
rect 10972 -57546 10978 -57486
rect 10282 -57670 10586 -57660
rect 10282 -57708 10366 -57670
rect 10574 -57708 10586 -57670
rect 10648 -57695 10654 -57635
rect 10714 -57695 10720 -57635
rect 10282 -57720 10586 -57708
rect 10282 -57768 10342 -57720
rect 10282 -58124 10294 -57768
rect 10330 -58124 10342 -57768
rect 10396 -57858 10456 -57720
rect 10526 -57768 10586 -57720
rect 10502 -57774 10610 -57768
rect 10502 -57808 10514 -57774
rect 10598 -57808 10610 -57774
rect 10502 -57814 10610 -57808
rect 10396 -57908 10410 -57858
rect 10404 -57995 10410 -57908
rect 10282 -58173 10342 -58124
rect 10398 -58034 10410 -57995
rect 10444 -57908 10456 -57858
rect 10654 -57858 10714 -57695
rect 10760 -57774 10868 -57768
rect 10760 -57808 10772 -57774
rect 10856 -57808 10868 -57774
rect 10760 -57814 10868 -57808
rect 10654 -57895 10668 -57858
rect 10444 -57995 10450 -57908
rect 10444 -58034 10458 -57995
rect 10398 -58173 10458 -58034
rect 10662 -58034 10668 -57895
rect 10702 -57895 10714 -57858
rect 10912 -57828 10972 -57546
rect 11170 -57635 11230 -57310
rect 11430 -57310 11442 -57272
rect 11476 -57272 11482 -56934
rect 11694 -56934 11740 -56922
rect 11694 -57267 11700 -56934
rect 11476 -57310 11490 -57272
rect 11276 -57369 11384 -57363
rect 11276 -57403 11288 -57369
rect 11372 -57403 11384 -57369
rect 11276 -57409 11384 -57403
rect 11430 -57486 11490 -57310
rect 11688 -57310 11700 -57267
rect 11734 -57267 11740 -56934
rect 11944 -56934 12004 -56786
rect 11944 -57152 11958 -56934
rect 11734 -57310 11748 -57267
rect 11952 -57280 11958 -57152
rect 11534 -57369 11642 -57363
rect 11534 -57403 11546 -57369
rect 11630 -57403 11642 -57369
rect 11534 -57409 11642 -57403
rect 11424 -57546 11430 -57486
rect 11490 -57546 11496 -57486
rect 11164 -57695 11170 -57635
rect 11230 -57695 11236 -57635
rect 11018 -57774 11126 -57768
rect 11018 -57808 11030 -57774
rect 11114 -57808 11126 -57774
rect 11018 -57814 11126 -57808
rect 10912 -57858 10974 -57828
rect 10912 -57894 10926 -57858
rect 10702 -58034 10708 -57895
rect 10662 -58046 10708 -58034
rect 10914 -58034 10926 -57894
rect 10960 -58034 10974 -57858
rect 11170 -57858 11230 -57695
rect 11276 -57774 11384 -57768
rect 11276 -57808 11288 -57774
rect 11372 -57808 11384 -57774
rect 11276 -57814 11384 -57808
rect 11170 -58014 11184 -57858
rect 10914 -58074 10974 -58034
rect 11178 -58034 11184 -58014
rect 11218 -58014 11230 -57858
rect 11430 -57858 11490 -57546
rect 11688 -57635 11748 -57310
rect 11946 -57310 11958 -57280
rect 11992 -57092 12004 -56934
rect 12058 -56834 12118 -56786
rect 12058 -57092 12070 -56834
rect 11992 -57152 12070 -57092
rect 11992 -57280 11998 -57152
rect 11992 -57310 12006 -57280
rect 11792 -57369 11900 -57363
rect 11792 -57403 11804 -57369
rect 11888 -57403 11900 -57369
rect 11792 -57409 11900 -57403
rect 11812 -57458 11872 -57409
rect 11946 -57458 12006 -57310
rect 12058 -57410 12070 -57152
rect 12106 -57210 12118 -56834
rect 12106 -57241 12456 -57210
rect 12106 -57275 12209 -57241
rect 12243 -57275 12301 -57241
rect 12335 -57275 12393 -57241
rect 12427 -57275 12456 -57241
rect 12106 -57306 12456 -57275
rect 12106 -57410 12118 -57306
rect 12058 -57458 12118 -57410
rect 11812 -57470 12118 -57458
rect 11812 -57504 11834 -57470
rect 12036 -57504 12118 -57470
rect 11812 -57518 12118 -57504
rect 12176 -57532 12236 -57526
rect 12524 -57532 12584 -57526
rect 12236 -57538 12298 -57532
rect 12236 -57586 12238 -57538
rect 12286 -57586 12298 -57538
rect 12236 -57592 12298 -57586
rect 12330 -57538 12524 -57532
rect 12330 -57586 12342 -57538
rect 12390 -57586 12524 -57538
rect 12330 -57592 12524 -57586
rect 12176 -57598 12236 -57592
rect 12524 -57598 12584 -57592
rect 11534 -57774 11642 -57768
rect 11534 -57808 11546 -57774
rect 11630 -57808 11642 -57774
rect 11534 -57814 11642 -57808
rect 11218 -58034 11224 -58014
rect 11178 -58046 11224 -58034
rect 11430 -58034 11442 -57858
rect 11476 -58034 11490 -57858
rect 11688 -57858 11748 -57695
rect 11818 -57668 12120 -57658
rect 11818 -57706 11838 -57668
rect 12036 -57706 12120 -57668
rect 11818 -57718 12120 -57706
rect 11818 -57768 11878 -57718
rect 11792 -57774 11900 -57768
rect 11792 -57808 11804 -57774
rect 11888 -57808 11900 -57774
rect 11792 -57814 11900 -57808
rect 11688 -57897 11700 -57858
rect 11430 -58074 11490 -58034
rect 11694 -58034 11700 -57897
rect 11734 -57897 11748 -57858
rect 11946 -57858 12006 -57718
rect 11734 -58034 11740 -57897
rect 11946 -57904 11958 -57858
rect 11952 -58001 11958 -57904
rect 11694 -58046 11740 -58034
rect 11944 -58034 11958 -58001
rect 11992 -57904 12006 -57858
rect 12060 -57754 12120 -57718
rect 13116 -57754 13122 -44048
rect 12060 -57768 13122 -57754
rect 11992 -58001 11998 -57904
rect 11992 -58034 12004 -58001
rect 10502 -58084 10610 -58078
rect 10502 -58118 10514 -58084
rect 10598 -58118 10610 -58084
rect 10502 -58124 10610 -58118
rect 10760 -58084 10868 -58078
rect 10760 -58118 10772 -58084
rect 10856 -58118 10868 -58084
rect 10760 -58124 10868 -58118
rect 10526 -58173 10586 -58124
rect 10282 -58184 10586 -58173
rect 10282 -58220 10364 -58184
rect 10572 -58220 10586 -58184
rect 10282 -58233 10586 -58220
rect 10282 -58390 10342 -58233
rect 10398 -58390 10458 -58233
rect 10526 -58390 10586 -58233
rect 10784 -58183 10844 -58124
rect 10908 -58134 10914 -58074
rect 10974 -58134 10980 -58074
rect 11018 -58084 11126 -58078
rect 11018 -58118 11030 -58084
rect 11114 -58118 11126 -58084
rect 11018 -58124 11126 -58118
rect 11276 -58084 11384 -58078
rect 11276 -58118 11288 -58084
rect 11372 -58118 11384 -58084
rect 11276 -58124 11384 -58118
rect 11044 -58183 11104 -58124
rect 11302 -58183 11362 -58124
rect 11424 -58134 11430 -58074
rect 11490 -58134 11496 -58074
rect 11534 -58084 11642 -58078
rect 11534 -58118 11546 -58084
rect 11630 -58118 11642 -58084
rect 11534 -58124 11642 -58118
rect 11792 -58084 11900 -58078
rect 11792 -58118 11804 -58084
rect 11888 -58118 11900 -58084
rect 11792 -58124 11900 -58118
rect 11558 -58183 11618 -58124
rect 11816 -58173 11876 -58124
rect 11944 -58173 12004 -58034
rect 12060 -58124 12070 -57768
rect 12108 -57785 13122 -57768
rect 12108 -57819 12209 -57785
rect 12243 -57819 12301 -57785
rect 12335 -57819 12393 -57785
rect 12427 -57819 13122 -57785
rect 12108 -57850 13122 -57819
rect 12108 -58124 12120 -57850
rect 12060 -58173 12120 -58124
rect 10784 -58243 11558 -58183
rect 11618 -58243 11624 -58183
rect 11816 -58186 12120 -58173
rect 11816 -58222 11836 -58186
rect 12038 -58222 12120 -58186
rect 11816 -58233 12120 -58222
rect 11816 -58390 11876 -58233
rect 11944 -58390 12004 -58233
rect 12060 -58390 12120 -58233
rect 13116 -58308 13122 -57850
rect 13222 -58308 13228 -44048
rect 23876 -44258 23882 -44198
rect 23942 -44258 23948 -44198
rect 23882 -44302 23942 -44258
rect 16248 -44362 23942 -44302
rect 16248 -44502 16308 -44362
rect 16758 -44412 16818 -44362
rect 16542 -44418 17030 -44412
rect 16542 -44452 16554 -44418
rect 17018 -44452 17030 -44418
rect 16542 -44458 17030 -44452
rect 16248 -44532 16260 -44502
rect 16254 -45060 16260 -44532
rect 16244 -45078 16260 -45060
rect 16294 -44532 16308 -44502
rect 17264 -44502 17324 -44362
rect 17766 -44412 17826 -44362
rect 18794 -44412 18854 -44362
rect 17560 -44418 18048 -44412
rect 17560 -44452 17572 -44418
rect 18036 -44452 18048 -44418
rect 17560 -44458 18048 -44452
rect 18578 -44418 19066 -44412
rect 18578 -44452 18590 -44418
rect 19054 -44452 19066 -44418
rect 18578 -44458 19066 -44452
rect 17264 -44526 17278 -44502
rect 16294 -45060 16300 -44532
rect 17272 -45056 17278 -44526
rect 16294 -45078 16304 -45060
rect 16244 -45320 16304 -45078
rect 17264 -45078 17278 -45056
rect 17312 -44526 17324 -44502
rect 18290 -44502 18336 -44490
rect 17312 -45056 17318 -44526
rect 18290 -45054 18296 -44502
rect 17312 -45078 17324 -45056
rect 16542 -45128 17030 -45122
rect 16542 -45162 16554 -45128
rect 17018 -45162 17030 -45128
rect 16542 -45168 17030 -45162
rect 16758 -45230 16818 -45168
rect 16542 -45236 17030 -45230
rect 16542 -45270 16554 -45236
rect 17018 -45270 17030 -45236
rect 16542 -45276 17030 -45270
rect 16244 -45350 16260 -45320
rect 16254 -45874 16260 -45350
rect 16246 -45896 16260 -45874
rect 16294 -45350 16304 -45320
rect 17264 -45320 17324 -45078
rect 18284 -45078 18296 -45054
rect 18330 -45054 18336 -44502
rect 19302 -44502 19362 -44362
rect 19808 -44412 19868 -44362
rect 20822 -44412 20882 -44362
rect 19596 -44418 20084 -44412
rect 19596 -44452 19608 -44418
rect 20072 -44452 20084 -44418
rect 19596 -44458 20084 -44452
rect 20614 -44418 21102 -44412
rect 20614 -44452 20626 -44418
rect 21090 -44452 21102 -44418
rect 20614 -44458 21102 -44452
rect 19302 -44540 19314 -44502
rect 18330 -45078 18344 -45054
rect 19308 -45058 19314 -44540
rect 17560 -45128 18048 -45122
rect 17560 -45162 17572 -45128
rect 18036 -45162 18048 -45128
rect 17560 -45168 18048 -45162
rect 17762 -45230 17822 -45168
rect 17560 -45236 18048 -45230
rect 17560 -45270 17572 -45236
rect 18036 -45270 18048 -45236
rect 17560 -45276 18048 -45270
rect 17264 -45346 17278 -45320
rect 16294 -45874 16300 -45350
rect 17272 -45870 17278 -45346
rect 16294 -45896 16306 -45874
rect 16246 -46138 16306 -45896
rect 17266 -45896 17278 -45870
rect 17312 -45346 17324 -45320
rect 18284 -45320 18344 -45078
rect 19302 -45078 19314 -45058
rect 19348 -44540 19362 -44502
rect 20326 -44502 20372 -44490
rect 21338 -44502 21398 -44362
rect 21854 -44412 21914 -44362
rect 22860 -44412 22920 -44362
rect 21632 -44418 22120 -44412
rect 21632 -44452 21644 -44418
rect 22108 -44452 22120 -44418
rect 21632 -44458 22120 -44452
rect 22650 -44418 23138 -44412
rect 22650 -44452 22662 -44418
rect 23126 -44452 23138 -44418
rect 22650 -44458 23138 -44452
rect 19348 -45058 19354 -44540
rect 20326 -45050 20332 -44502
rect 19348 -45078 19362 -45058
rect 18578 -45128 19066 -45122
rect 18578 -45162 18590 -45128
rect 19054 -45162 19066 -45128
rect 18578 -45168 19066 -45162
rect 18792 -45230 18852 -45168
rect 18578 -45236 19066 -45230
rect 18578 -45270 18590 -45236
rect 19054 -45270 19066 -45236
rect 18578 -45276 19066 -45270
rect 18284 -45344 18296 -45320
rect 17312 -45870 17318 -45346
rect 18290 -45868 18296 -45344
rect 17312 -45896 17326 -45870
rect 16542 -45946 17030 -45940
rect 16542 -45980 16554 -45946
rect 17018 -45980 17030 -45946
rect 16542 -45986 17030 -45980
rect 16758 -46048 16818 -45986
rect 16542 -46054 17030 -46048
rect 16542 -46088 16554 -46054
rect 17018 -46088 17030 -46054
rect 16542 -46094 17030 -46088
rect 16246 -46164 16260 -46138
rect 16254 -46702 16260 -46164
rect 16246 -46714 16260 -46702
rect 16294 -46164 16306 -46138
rect 17266 -46138 17326 -45896
rect 18286 -45896 18296 -45868
rect 18330 -45344 18344 -45320
rect 19302 -45320 19362 -45078
rect 20322 -45078 20332 -45050
rect 20366 -45050 20372 -44502
rect 21336 -44536 21350 -44502
rect 21338 -44548 21350 -44536
rect 20366 -45078 20382 -45050
rect 21344 -45058 21350 -44548
rect 19596 -45128 20084 -45122
rect 19596 -45162 19608 -45128
rect 20072 -45162 20084 -45128
rect 19596 -45168 20084 -45162
rect 19794 -45230 19854 -45168
rect 19596 -45236 20084 -45230
rect 19596 -45270 19608 -45236
rect 20072 -45270 20084 -45236
rect 19596 -45276 20084 -45270
rect 18330 -45868 18336 -45344
rect 19302 -45348 19314 -45320
rect 18330 -45896 18346 -45868
rect 19308 -45872 19314 -45348
rect 17560 -45946 18048 -45940
rect 17560 -45980 17572 -45946
rect 18036 -45980 18048 -45946
rect 17560 -45986 18048 -45980
rect 17774 -46048 17834 -45986
rect 17560 -46054 18048 -46048
rect 17560 -46088 17572 -46054
rect 18036 -46088 18048 -46054
rect 17560 -46094 18048 -46088
rect 17266 -46160 17278 -46138
rect 16294 -46702 16300 -46164
rect 17272 -46698 17278 -46160
rect 16294 -46714 16306 -46702
rect 16246 -46956 16306 -46714
rect 17266 -46714 17278 -46698
rect 17312 -46160 17326 -46138
rect 18286 -46138 18346 -45896
rect 19304 -45896 19314 -45872
rect 19348 -45348 19362 -45320
rect 20322 -45320 20382 -45078
rect 21334 -45078 21350 -45058
rect 21384 -44548 21398 -44502
rect 22362 -44502 22408 -44490
rect 21384 -45058 21390 -44548
rect 22362 -45058 22368 -44502
rect 21384 -45078 21394 -45058
rect 20614 -45128 21102 -45122
rect 20614 -45162 20626 -45128
rect 21090 -45162 21102 -45128
rect 20614 -45168 21102 -45162
rect 20824 -45230 20884 -45168
rect 20614 -45236 21102 -45230
rect 20614 -45270 20626 -45236
rect 21090 -45270 21102 -45236
rect 20614 -45276 21102 -45270
rect 20322 -45340 20332 -45320
rect 19348 -45872 19354 -45348
rect 20326 -45864 20332 -45340
rect 19348 -45896 19364 -45872
rect 18578 -45946 19066 -45940
rect 18578 -45980 18590 -45946
rect 19054 -45980 19066 -45946
rect 18578 -45986 19066 -45980
rect 18792 -46048 18852 -45986
rect 18578 -46054 19066 -46048
rect 18578 -46088 18590 -46054
rect 19054 -46088 19066 -46054
rect 18578 -46094 19066 -46088
rect 18286 -46158 18296 -46138
rect 17312 -46698 17318 -46160
rect 18290 -46696 18296 -46158
rect 17312 -46714 17326 -46698
rect 16542 -46764 17030 -46758
rect 16542 -46798 16554 -46764
rect 17018 -46798 17030 -46764
rect 16542 -46804 17030 -46798
rect 16752 -46866 16812 -46804
rect 16542 -46872 17030 -46866
rect 16542 -46906 16554 -46872
rect 17018 -46906 17030 -46872
rect 16542 -46912 17030 -46906
rect 16246 -46992 16260 -46956
rect 16254 -47514 16260 -46992
rect 16246 -47532 16260 -47514
rect 16294 -46992 16306 -46956
rect 17266 -46956 17326 -46714
rect 18286 -46714 18296 -46696
rect 18330 -46158 18346 -46138
rect 19304 -46138 19364 -45896
rect 20324 -45896 20332 -45864
rect 20366 -45340 20382 -45320
rect 21334 -45320 21394 -45078
rect 22356 -45078 22368 -45058
rect 22402 -45058 22408 -44502
rect 23372 -44502 23432 -44362
rect 23882 -44412 23942 -44362
rect 25402 -44392 25408 -44332
rect 25468 -44392 25474 -44332
rect 23668 -44418 24156 -44412
rect 23668 -44452 23680 -44418
rect 24144 -44452 24156 -44418
rect 23668 -44458 24156 -44452
rect 24686 -44418 25174 -44412
rect 24686 -44452 24698 -44418
rect 25162 -44452 25174 -44418
rect 24686 -44458 25174 -44452
rect 23372 -44538 23386 -44502
rect 23380 -45058 23386 -44538
rect 22402 -45078 22416 -45058
rect 21632 -45128 22120 -45122
rect 21632 -45162 21644 -45128
rect 22108 -45162 22120 -45128
rect 21632 -45168 22120 -45162
rect 21840 -45230 21900 -45168
rect 21632 -45236 22120 -45230
rect 21632 -45270 21644 -45236
rect 22108 -45270 22120 -45236
rect 21632 -45276 22120 -45270
rect 20366 -45864 20372 -45340
rect 21334 -45348 21350 -45320
rect 20366 -45896 20384 -45864
rect 21344 -45872 21350 -45348
rect 19596 -45946 20084 -45940
rect 19596 -45980 19608 -45946
rect 20072 -45980 20084 -45946
rect 19596 -45986 20084 -45980
rect 19794 -46048 19854 -45986
rect 19596 -46054 20084 -46048
rect 19596 -46088 19608 -46054
rect 20072 -46088 20084 -46054
rect 19596 -46094 20084 -46088
rect 18330 -46696 18336 -46158
rect 19304 -46162 19314 -46138
rect 18330 -46714 18346 -46696
rect 19308 -46700 19314 -46162
rect 17560 -46764 18048 -46758
rect 17560 -46798 17572 -46764
rect 18036 -46798 18048 -46764
rect 17560 -46804 18048 -46798
rect 17774 -46866 17834 -46804
rect 17560 -46872 18048 -46866
rect 17560 -46906 17572 -46872
rect 18036 -46906 18048 -46872
rect 17560 -46912 18048 -46906
rect 17266 -46988 17278 -46956
rect 16294 -47514 16300 -46992
rect 17272 -47510 17278 -46988
rect 16294 -47532 16306 -47514
rect 16246 -47774 16306 -47532
rect 17266 -47532 17278 -47510
rect 17312 -46988 17326 -46956
rect 18286 -46956 18346 -46714
rect 19304 -46714 19314 -46700
rect 19348 -46162 19364 -46138
rect 20324 -46138 20384 -45896
rect 21336 -45896 21350 -45872
rect 21384 -45348 21394 -45320
rect 22356 -45320 22416 -45078
rect 23376 -45078 23386 -45058
rect 23420 -44538 23432 -44502
rect 24398 -44502 24444 -44490
rect 23420 -45058 23426 -44538
rect 24398 -45054 24404 -44502
rect 23420 -45078 23436 -45058
rect 22650 -45128 23138 -45122
rect 22650 -45162 22662 -45128
rect 23126 -45162 23138 -45128
rect 22650 -45168 23138 -45162
rect 22862 -45230 22922 -45168
rect 22650 -45236 23138 -45230
rect 22650 -45270 22662 -45236
rect 23126 -45270 23138 -45236
rect 22650 -45276 23138 -45270
rect 22356 -45348 22368 -45320
rect 21384 -45872 21390 -45348
rect 22362 -45872 22368 -45348
rect 21384 -45896 21396 -45872
rect 20614 -45946 21102 -45940
rect 20614 -45980 20626 -45946
rect 21090 -45980 21102 -45946
rect 20614 -45986 21102 -45980
rect 20824 -46048 20884 -45986
rect 20614 -46054 21102 -46048
rect 20614 -46088 20626 -46054
rect 21090 -46088 21102 -46054
rect 20614 -46094 21102 -46088
rect 20324 -46154 20332 -46138
rect 19348 -46700 19354 -46162
rect 20326 -46692 20332 -46154
rect 19348 -46714 19364 -46700
rect 18578 -46764 19066 -46758
rect 18578 -46798 18590 -46764
rect 19054 -46798 19066 -46764
rect 18578 -46804 19066 -46798
rect 18786 -46866 18846 -46804
rect 18578 -46872 19066 -46866
rect 18578 -46906 18590 -46872
rect 19054 -46906 19066 -46872
rect 18578 -46912 19066 -46906
rect 18286 -46986 18296 -46956
rect 17312 -47510 17318 -46988
rect 18290 -47508 18296 -46986
rect 17312 -47532 17326 -47510
rect 16542 -47582 17030 -47576
rect 16542 -47616 16554 -47582
rect 17018 -47616 17030 -47582
rect 16542 -47622 17030 -47616
rect 16750 -47684 16810 -47622
rect 16542 -47690 17030 -47684
rect 16542 -47724 16554 -47690
rect 17018 -47724 17030 -47690
rect 16542 -47730 17030 -47724
rect 16246 -47804 16260 -47774
rect 16254 -48334 16260 -47804
rect 16246 -48350 16260 -48334
rect 16294 -47804 16306 -47774
rect 17266 -47774 17326 -47532
rect 18286 -47532 18296 -47508
rect 18330 -46986 18346 -46956
rect 19304 -46956 19364 -46714
rect 20324 -46714 20332 -46692
rect 20366 -46154 20384 -46138
rect 21336 -46138 21396 -45896
rect 22358 -45896 22368 -45872
rect 22402 -45348 22416 -45320
rect 23376 -45320 23436 -45078
rect 24392 -45078 24404 -45054
rect 24438 -45054 24444 -44502
rect 25408 -44502 25468 -44392
rect 25408 -44538 25422 -44502
rect 24438 -45078 24452 -45054
rect 25416 -45058 25422 -44538
rect 23668 -45128 24156 -45122
rect 23668 -45162 23680 -45128
rect 24144 -45162 24156 -45128
rect 23668 -45168 24156 -45162
rect 23874 -45230 23934 -45168
rect 23668 -45236 24156 -45230
rect 23668 -45270 23680 -45236
rect 24144 -45270 24156 -45236
rect 23668 -45276 24156 -45270
rect 23376 -45348 23386 -45320
rect 22402 -45872 22408 -45348
rect 23380 -45872 23386 -45348
rect 22402 -45896 22418 -45872
rect 21632 -45946 22120 -45940
rect 21632 -45980 21644 -45946
rect 22108 -45980 22120 -45946
rect 21632 -45986 22120 -45980
rect 21840 -46048 21900 -45986
rect 21632 -46054 22120 -46048
rect 21632 -46088 21644 -46054
rect 22108 -46088 22120 -46054
rect 21632 -46094 22120 -46088
rect 20366 -46692 20372 -46154
rect 21336 -46162 21350 -46138
rect 20366 -46714 20384 -46692
rect 21344 -46700 21350 -46162
rect 19596 -46764 20084 -46758
rect 19596 -46798 19608 -46764
rect 20072 -46798 20084 -46764
rect 19596 -46804 20084 -46798
rect 19788 -46866 19848 -46804
rect 19596 -46872 20084 -46866
rect 19596 -46906 19608 -46872
rect 20072 -46906 20084 -46872
rect 19596 -46912 20084 -46906
rect 18330 -47508 18336 -46986
rect 19304 -46990 19314 -46956
rect 18330 -47532 18346 -47508
rect 19308 -47512 19314 -46990
rect 17560 -47582 18048 -47576
rect 17560 -47616 17572 -47582
rect 18036 -47616 18048 -47582
rect 17560 -47622 18048 -47616
rect 17768 -47684 17828 -47622
rect 17560 -47690 18048 -47684
rect 17560 -47724 17572 -47690
rect 18036 -47724 18048 -47690
rect 17560 -47730 18048 -47724
rect 17266 -47800 17278 -47774
rect 16294 -48334 16300 -47804
rect 17272 -48330 17278 -47800
rect 16294 -48350 16306 -48334
rect 16246 -48592 16306 -48350
rect 17266 -48350 17278 -48330
rect 17312 -47800 17326 -47774
rect 18286 -47774 18346 -47532
rect 19304 -47532 19314 -47512
rect 19348 -46990 19364 -46956
rect 20324 -46956 20384 -46714
rect 21336 -46714 21350 -46700
rect 21384 -46162 21396 -46138
rect 22358 -46138 22418 -45896
rect 23378 -45896 23386 -45872
rect 23420 -45348 23436 -45320
rect 24392 -45320 24452 -45078
rect 25414 -45078 25422 -45058
rect 25456 -44538 25468 -44502
rect 25456 -45058 25462 -44538
rect 25456 -45078 25474 -45058
rect 24686 -45128 25174 -45122
rect 24686 -45162 24698 -45128
rect 25162 -45162 25174 -45128
rect 24686 -45168 25174 -45162
rect 24894 -45230 24954 -45168
rect 24686 -45236 25174 -45230
rect 24686 -45270 24698 -45236
rect 25162 -45270 25174 -45236
rect 24686 -45276 25174 -45270
rect 24392 -45344 24404 -45320
rect 23420 -45872 23426 -45348
rect 24398 -45868 24404 -45344
rect 23420 -45896 23438 -45872
rect 22650 -45946 23138 -45940
rect 22650 -45980 22662 -45946
rect 23126 -45980 23138 -45946
rect 22650 -45986 23138 -45980
rect 22862 -46048 22922 -45986
rect 22650 -46054 23138 -46048
rect 22650 -46088 22662 -46054
rect 23126 -46088 23138 -46054
rect 22650 -46094 23138 -46088
rect 22358 -46162 22368 -46138
rect 21384 -46700 21390 -46162
rect 22362 -46700 22368 -46162
rect 21384 -46714 21396 -46700
rect 20614 -46764 21102 -46758
rect 20614 -46798 20626 -46764
rect 21090 -46798 21102 -46764
rect 20614 -46804 21102 -46798
rect 20818 -46866 20878 -46804
rect 20614 -46872 21102 -46866
rect 20614 -46906 20626 -46872
rect 21090 -46906 21102 -46872
rect 20614 -46912 21102 -46906
rect 20324 -46982 20332 -46956
rect 19348 -47512 19354 -46990
rect 20326 -47504 20332 -46982
rect 19348 -47532 19364 -47512
rect 18578 -47582 19066 -47576
rect 18578 -47616 18590 -47582
rect 19054 -47616 19066 -47582
rect 18578 -47622 19066 -47616
rect 18784 -47684 18844 -47622
rect 18578 -47690 19066 -47684
rect 18578 -47724 18590 -47690
rect 19054 -47724 19066 -47690
rect 18578 -47730 19066 -47724
rect 18286 -47798 18296 -47774
rect 17312 -48330 17318 -47800
rect 18290 -48328 18296 -47798
rect 17312 -48350 17326 -48330
rect 16542 -48400 17030 -48394
rect 16542 -48434 16554 -48400
rect 17018 -48434 17030 -48400
rect 16542 -48440 17030 -48434
rect 16752 -48502 16812 -48440
rect 16542 -48508 17030 -48502
rect 16542 -48542 16554 -48508
rect 17018 -48542 17030 -48508
rect 16542 -48548 17030 -48542
rect 16246 -48624 16260 -48592
rect 16254 -49146 16260 -48624
rect 16246 -49168 16260 -49146
rect 16294 -48624 16306 -48592
rect 17266 -48592 17326 -48350
rect 18286 -48350 18296 -48328
rect 18330 -47798 18346 -47774
rect 19304 -47774 19364 -47532
rect 20324 -47532 20332 -47504
rect 20366 -46982 20384 -46956
rect 21336 -46956 21396 -46714
rect 22358 -46714 22368 -46700
rect 22402 -46162 22418 -46138
rect 23378 -46138 23438 -45896
rect 24394 -45896 24404 -45868
rect 24438 -45344 24452 -45320
rect 25414 -45320 25474 -45078
rect 24438 -45868 24444 -45344
rect 25414 -45348 25422 -45320
rect 24438 -45896 24454 -45868
rect 23668 -45946 24156 -45940
rect 23668 -45980 23680 -45946
rect 24144 -45980 24156 -45946
rect 23668 -45986 24156 -45980
rect 23874 -46048 23934 -45986
rect 23668 -46054 24156 -46048
rect 23668 -46088 23680 -46054
rect 24144 -46088 24156 -46054
rect 23668 -46094 24156 -46088
rect 23378 -46162 23386 -46138
rect 22402 -46700 22408 -46162
rect 23380 -46700 23386 -46162
rect 22402 -46714 22418 -46700
rect 21632 -46764 22120 -46758
rect 21632 -46798 21644 -46764
rect 22108 -46798 22120 -46764
rect 21632 -46804 22120 -46798
rect 21834 -46866 21894 -46804
rect 21632 -46872 22120 -46866
rect 21632 -46906 21644 -46872
rect 22108 -46906 22120 -46872
rect 21632 -46912 22120 -46906
rect 20366 -47504 20372 -46982
rect 21336 -46990 21350 -46956
rect 20366 -47532 20384 -47504
rect 21344 -47512 21350 -46990
rect 19596 -47582 20084 -47576
rect 19596 -47616 19608 -47582
rect 20072 -47616 20084 -47582
rect 19596 -47622 20084 -47616
rect 19786 -47684 19846 -47622
rect 19596 -47690 20084 -47684
rect 19596 -47724 19608 -47690
rect 20072 -47724 20084 -47690
rect 19596 -47730 20084 -47724
rect 18330 -48328 18336 -47798
rect 19304 -47802 19314 -47774
rect 18330 -48350 18346 -48328
rect 19308 -48332 19314 -47802
rect 17560 -48400 18048 -48394
rect 17560 -48434 17572 -48400
rect 18036 -48434 18048 -48400
rect 17560 -48440 18048 -48434
rect 17766 -48502 17826 -48440
rect 17560 -48508 18048 -48502
rect 17560 -48542 17572 -48508
rect 18036 -48542 18048 -48508
rect 17560 -48548 18048 -48542
rect 17266 -48620 17278 -48592
rect 16294 -49146 16300 -48624
rect 17272 -49142 17278 -48620
rect 16294 -49168 16306 -49146
rect 16246 -49410 16306 -49168
rect 17266 -49168 17278 -49142
rect 17312 -48620 17326 -48592
rect 18286 -48592 18346 -48350
rect 19304 -48350 19314 -48332
rect 19348 -47802 19364 -47774
rect 20324 -47774 20384 -47532
rect 21336 -47532 21350 -47512
rect 21384 -46990 21396 -46956
rect 22358 -46956 22418 -46714
rect 23378 -46714 23386 -46700
rect 23420 -46162 23438 -46138
rect 24394 -46138 24454 -45896
rect 25416 -45896 25422 -45348
rect 25456 -45348 25474 -45320
rect 25456 -45872 25462 -45348
rect 25456 -45896 25476 -45872
rect 24686 -45946 25174 -45940
rect 24686 -45980 24698 -45946
rect 25162 -45980 25174 -45946
rect 24686 -45986 25174 -45980
rect 24894 -46048 24954 -45986
rect 24686 -46054 25174 -46048
rect 24686 -46088 24698 -46054
rect 25162 -46088 25174 -46054
rect 24686 -46094 25174 -46088
rect 24394 -46158 24404 -46138
rect 23420 -46700 23426 -46162
rect 24398 -46696 24404 -46158
rect 23420 -46714 23438 -46700
rect 22650 -46764 23138 -46758
rect 22650 -46798 22662 -46764
rect 23126 -46798 23138 -46764
rect 22650 -46804 23138 -46798
rect 22856 -46866 22916 -46804
rect 22650 -46872 23138 -46866
rect 22650 -46906 22662 -46872
rect 23126 -46906 23138 -46872
rect 22650 -46912 23138 -46906
rect 22358 -46990 22368 -46956
rect 21384 -47512 21390 -46990
rect 22362 -47512 22368 -46990
rect 21384 -47532 21396 -47512
rect 20614 -47582 21102 -47576
rect 20614 -47616 20626 -47582
rect 21090 -47616 21102 -47582
rect 20614 -47622 21102 -47616
rect 20816 -47684 20876 -47622
rect 20614 -47690 21102 -47684
rect 20614 -47724 20626 -47690
rect 21090 -47724 21102 -47690
rect 20614 -47730 21102 -47724
rect 20324 -47794 20332 -47774
rect 19348 -48332 19354 -47802
rect 20326 -48324 20332 -47794
rect 19348 -48350 19364 -48332
rect 18578 -48400 19066 -48394
rect 18578 -48434 18590 -48400
rect 19054 -48434 19066 -48400
rect 18578 -48440 19066 -48434
rect 18786 -48502 18846 -48440
rect 18578 -48508 19066 -48502
rect 18578 -48542 18590 -48508
rect 19054 -48542 19066 -48508
rect 18578 -48548 19066 -48542
rect 18286 -48618 18296 -48592
rect 17312 -49142 17318 -48620
rect 18290 -49140 18296 -48618
rect 17312 -49168 17326 -49142
rect 16542 -49218 17030 -49212
rect 16542 -49252 16554 -49218
rect 17018 -49252 17030 -49218
rect 16542 -49258 17030 -49252
rect 16754 -49320 16814 -49258
rect 16542 -49326 17030 -49320
rect 16542 -49360 16554 -49326
rect 17018 -49360 17030 -49326
rect 16542 -49366 17030 -49360
rect 16246 -49436 16260 -49410
rect 16254 -49964 16260 -49436
rect 16246 -49986 16260 -49964
rect 16294 -49436 16306 -49410
rect 17266 -49410 17326 -49168
rect 18286 -49168 18296 -49140
rect 18330 -48618 18346 -48592
rect 19304 -48592 19364 -48350
rect 20324 -48350 20332 -48324
rect 20366 -47794 20384 -47774
rect 21336 -47774 21396 -47532
rect 22358 -47532 22368 -47512
rect 22402 -46990 22418 -46956
rect 23378 -46956 23438 -46714
rect 24394 -46714 24404 -46696
rect 24438 -46158 24454 -46138
rect 25416 -46138 25476 -45896
rect 24438 -46696 24444 -46158
rect 24438 -46714 24454 -46696
rect 23668 -46764 24156 -46758
rect 23668 -46798 23680 -46764
rect 24144 -46798 24156 -46764
rect 23668 -46804 24156 -46798
rect 23868 -46866 23928 -46804
rect 23668 -46872 24156 -46866
rect 23668 -46906 23680 -46872
rect 24144 -46906 24156 -46872
rect 23668 -46912 24156 -46906
rect 23378 -46990 23386 -46956
rect 22402 -47512 22408 -46990
rect 23380 -47512 23386 -46990
rect 22402 -47532 22418 -47512
rect 21632 -47582 22120 -47576
rect 21632 -47616 21644 -47582
rect 22108 -47616 22120 -47582
rect 21632 -47622 22120 -47616
rect 21832 -47684 21892 -47622
rect 21632 -47690 22120 -47684
rect 21632 -47724 21644 -47690
rect 22108 -47724 22120 -47690
rect 21632 -47730 22120 -47724
rect 20366 -48324 20372 -47794
rect 21336 -47802 21350 -47774
rect 20366 -48350 20384 -48324
rect 21344 -48332 21350 -47802
rect 19596 -48400 20084 -48394
rect 19596 -48434 19608 -48400
rect 20072 -48434 20084 -48400
rect 19596 -48440 20084 -48434
rect 19788 -48502 19848 -48440
rect 19596 -48508 20084 -48502
rect 19596 -48542 19608 -48508
rect 20072 -48542 20084 -48508
rect 19596 -48548 20084 -48542
rect 18330 -49140 18336 -48618
rect 19304 -48622 19314 -48592
rect 18330 -49168 18346 -49140
rect 19308 -49144 19314 -48622
rect 17560 -49218 18048 -49212
rect 17560 -49252 17572 -49218
rect 18036 -49252 18048 -49218
rect 17560 -49258 18048 -49252
rect 17768 -49320 17828 -49258
rect 17560 -49326 18048 -49320
rect 17560 -49360 17572 -49326
rect 18036 -49360 18048 -49326
rect 17560 -49366 18048 -49360
rect 17266 -49432 17278 -49410
rect 16294 -49964 16300 -49436
rect 17272 -49960 17278 -49432
rect 16294 -49986 16306 -49964
rect 16246 -50228 16306 -49986
rect 17266 -49986 17278 -49960
rect 17312 -49432 17326 -49410
rect 18286 -49410 18346 -49168
rect 19304 -49168 19314 -49144
rect 19348 -48622 19364 -48592
rect 20324 -48592 20384 -48350
rect 21336 -48350 21350 -48332
rect 21384 -47802 21396 -47774
rect 22358 -47774 22418 -47532
rect 23378 -47532 23386 -47512
rect 23420 -46990 23438 -46956
rect 24394 -46956 24454 -46714
rect 25416 -46714 25422 -46138
rect 25456 -46162 25476 -46138
rect 25456 -46700 25462 -46162
rect 25456 -46714 25476 -46700
rect 24686 -46764 25174 -46758
rect 24686 -46798 24698 -46764
rect 25162 -46798 25174 -46764
rect 24686 -46804 25174 -46798
rect 24888 -46866 24948 -46804
rect 24686 -46872 25174 -46866
rect 24686 -46906 24698 -46872
rect 25162 -46906 25174 -46872
rect 24686 -46912 25174 -46906
rect 24394 -46986 24404 -46956
rect 23420 -47512 23426 -46990
rect 24398 -47508 24404 -46986
rect 23420 -47532 23438 -47512
rect 22650 -47582 23138 -47576
rect 22650 -47616 22662 -47582
rect 23126 -47616 23138 -47582
rect 22650 -47622 23138 -47616
rect 22854 -47684 22914 -47622
rect 22650 -47690 23138 -47684
rect 22650 -47724 22662 -47690
rect 23126 -47724 23138 -47690
rect 22650 -47730 23138 -47724
rect 22358 -47802 22368 -47774
rect 21384 -48332 21390 -47802
rect 22362 -48332 22368 -47802
rect 21384 -48350 21396 -48332
rect 20614 -48400 21102 -48394
rect 20614 -48434 20626 -48400
rect 21090 -48434 21102 -48400
rect 20614 -48440 21102 -48434
rect 20818 -48502 20878 -48440
rect 20614 -48508 21102 -48502
rect 20614 -48542 20626 -48508
rect 21090 -48542 21102 -48508
rect 20614 -48548 21102 -48542
rect 20324 -48614 20332 -48592
rect 19348 -49144 19354 -48622
rect 20326 -49136 20332 -48614
rect 19348 -49168 19364 -49144
rect 18578 -49218 19066 -49212
rect 18578 -49252 18590 -49218
rect 19054 -49252 19066 -49218
rect 18578 -49258 19066 -49252
rect 18788 -49320 18848 -49258
rect 18578 -49326 19066 -49320
rect 18578 -49360 18590 -49326
rect 19054 -49360 19066 -49326
rect 18578 -49366 19066 -49360
rect 18286 -49430 18296 -49410
rect 17312 -49960 17318 -49432
rect 18290 -49958 18296 -49430
rect 17312 -49986 17326 -49960
rect 16542 -50036 17030 -50030
rect 16542 -50070 16554 -50036
rect 17018 -50070 17030 -50036
rect 16542 -50076 17030 -50070
rect 16756 -50138 16816 -50076
rect 16542 -50144 17030 -50138
rect 16542 -50178 16554 -50144
rect 17018 -50178 17030 -50144
rect 16542 -50184 17030 -50178
rect 16246 -50254 16260 -50228
rect 16254 -50804 16260 -50254
rect 16294 -50254 16306 -50228
rect 17266 -50228 17326 -49986
rect 18286 -49986 18296 -49958
rect 18330 -49430 18346 -49410
rect 19304 -49410 19364 -49168
rect 20324 -49168 20332 -49136
rect 20366 -48614 20384 -48592
rect 21336 -48592 21396 -48350
rect 22358 -48350 22368 -48332
rect 22402 -47802 22418 -47774
rect 23378 -47774 23438 -47532
rect 24394 -47532 24404 -47508
rect 24438 -46986 24454 -46956
rect 25416 -46956 25476 -46714
rect 24438 -47508 24444 -46986
rect 24438 -47532 24454 -47508
rect 23668 -47582 24156 -47576
rect 23668 -47616 23680 -47582
rect 24144 -47616 24156 -47582
rect 23668 -47622 24156 -47616
rect 23866 -47684 23926 -47622
rect 23668 -47690 24156 -47684
rect 23668 -47724 23680 -47690
rect 24144 -47724 24156 -47690
rect 23668 -47730 24156 -47724
rect 23378 -47802 23386 -47774
rect 22402 -48332 22408 -47802
rect 23380 -48332 23386 -47802
rect 22402 -48350 22418 -48332
rect 21632 -48400 22120 -48394
rect 21632 -48434 21644 -48400
rect 22108 -48434 22120 -48400
rect 21632 -48440 22120 -48434
rect 21834 -48502 21894 -48440
rect 21632 -48508 22120 -48502
rect 21632 -48542 21644 -48508
rect 22108 -48542 22120 -48508
rect 21632 -48548 22120 -48542
rect 20366 -49136 20372 -48614
rect 21336 -48622 21350 -48592
rect 20366 -49168 20384 -49136
rect 21344 -49144 21350 -48622
rect 19596 -49218 20084 -49212
rect 19596 -49252 19608 -49218
rect 20072 -49252 20084 -49218
rect 19596 -49258 20084 -49252
rect 19790 -49320 19850 -49258
rect 19596 -49326 20084 -49320
rect 19596 -49360 19608 -49326
rect 20072 -49360 20084 -49326
rect 19596 -49366 20084 -49360
rect 18330 -49958 18336 -49430
rect 19304 -49434 19314 -49410
rect 18330 -49986 18346 -49958
rect 19308 -49962 19314 -49434
rect 17560 -50036 18048 -50030
rect 17560 -50070 17572 -50036
rect 18036 -50070 18048 -50036
rect 17560 -50076 18048 -50070
rect 17770 -50138 17830 -50076
rect 17560 -50144 18048 -50138
rect 17560 -50178 17572 -50144
rect 18036 -50178 18048 -50144
rect 17560 -50184 18048 -50178
rect 17266 -50250 17278 -50228
rect 16294 -50804 16300 -50254
rect 16254 -50816 16300 -50804
rect 17272 -50804 17278 -50250
rect 17312 -50250 17326 -50228
rect 18286 -50228 18346 -49986
rect 19304 -49986 19314 -49962
rect 19348 -49434 19364 -49410
rect 20324 -49410 20384 -49168
rect 21336 -49168 21350 -49144
rect 21384 -48622 21396 -48592
rect 22358 -48592 22418 -48350
rect 23378 -48350 23386 -48332
rect 23420 -47802 23438 -47774
rect 24394 -47774 24454 -47532
rect 25416 -47532 25422 -46956
rect 25456 -46990 25476 -46956
rect 25456 -47512 25462 -46990
rect 25456 -47532 25476 -47512
rect 24686 -47582 25174 -47576
rect 24686 -47616 24698 -47582
rect 25162 -47616 25174 -47582
rect 24686 -47622 25174 -47616
rect 24886 -47684 24946 -47622
rect 24686 -47690 25174 -47684
rect 24686 -47724 24698 -47690
rect 25162 -47724 25174 -47690
rect 24686 -47730 25174 -47724
rect 24394 -47798 24404 -47774
rect 23420 -48332 23426 -47802
rect 24398 -48328 24404 -47798
rect 23420 -48350 23438 -48332
rect 22650 -48400 23138 -48394
rect 22650 -48434 22662 -48400
rect 23126 -48434 23138 -48400
rect 22650 -48440 23138 -48434
rect 22856 -48502 22916 -48440
rect 22650 -48508 23138 -48502
rect 22650 -48542 22662 -48508
rect 23126 -48542 23138 -48508
rect 22650 -48548 23138 -48542
rect 22358 -48622 22368 -48592
rect 21384 -49144 21390 -48622
rect 22362 -49144 22368 -48622
rect 21384 -49168 21396 -49144
rect 20614 -49218 21102 -49212
rect 20614 -49252 20626 -49218
rect 21090 -49252 21102 -49218
rect 20614 -49258 21102 -49252
rect 20820 -49320 20880 -49258
rect 20614 -49326 21102 -49320
rect 20614 -49360 20626 -49326
rect 21090 -49360 21102 -49326
rect 20614 -49366 21102 -49360
rect 20324 -49426 20332 -49410
rect 19348 -49962 19354 -49434
rect 20326 -49954 20332 -49426
rect 19348 -49986 19364 -49962
rect 18578 -50036 19066 -50030
rect 18578 -50070 18590 -50036
rect 19054 -50070 19066 -50036
rect 18578 -50076 19066 -50070
rect 18790 -50138 18850 -50076
rect 18578 -50144 19066 -50138
rect 18578 -50178 18590 -50144
rect 19054 -50178 19066 -50144
rect 18578 -50184 19066 -50178
rect 18286 -50248 18296 -50228
rect 17312 -50804 17318 -50250
rect 18290 -50758 18296 -50248
rect 17272 -50816 17318 -50804
rect 18280 -50804 18296 -50758
rect 18330 -50248 18346 -50228
rect 19304 -50228 19364 -49986
rect 20324 -49986 20332 -49954
rect 20366 -49426 20384 -49410
rect 21336 -49410 21396 -49168
rect 22358 -49168 22368 -49144
rect 22402 -48622 22418 -48592
rect 23378 -48592 23438 -48350
rect 24394 -48350 24404 -48328
rect 24438 -47798 24454 -47774
rect 25416 -47774 25476 -47532
rect 24438 -48328 24444 -47798
rect 24438 -48350 24454 -48328
rect 23668 -48400 24156 -48394
rect 23668 -48434 23680 -48400
rect 24144 -48434 24156 -48400
rect 23668 -48440 24156 -48434
rect 23868 -48502 23928 -48440
rect 23668 -48508 24156 -48502
rect 23668 -48542 23680 -48508
rect 24144 -48542 24156 -48508
rect 23668 -48548 24156 -48542
rect 23378 -48622 23386 -48592
rect 22402 -49144 22408 -48622
rect 23380 -49144 23386 -48622
rect 22402 -49168 22418 -49144
rect 21632 -49218 22120 -49212
rect 21632 -49252 21644 -49218
rect 22108 -49252 22120 -49218
rect 21632 -49258 22120 -49252
rect 21836 -49320 21896 -49258
rect 21632 -49326 22120 -49320
rect 21632 -49360 21644 -49326
rect 22108 -49360 22120 -49326
rect 21632 -49366 22120 -49360
rect 20366 -49954 20372 -49426
rect 21336 -49434 21350 -49410
rect 20366 -49986 20384 -49954
rect 21344 -49962 21350 -49434
rect 19596 -50036 20084 -50030
rect 19596 -50070 19608 -50036
rect 20072 -50070 20084 -50036
rect 19596 -50076 20084 -50070
rect 19792 -50138 19852 -50076
rect 19596 -50144 20084 -50138
rect 19596 -50178 19608 -50144
rect 20072 -50178 20084 -50144
rect 19596 -50184 20084 -50178
rect 18330 -50758 18336 -50248
rect 19304 -50252 19314 -50228
rect 18330 -50804 18340 -50758
rect 16542 -50854 17030 -50848
rect 16542 -50888 16554 -50854
rect 17018 -50888 17030 -50854
rect 16542 -50894 17030 -50888
rect 17560 -50854 18048 -50848
rect 17560 -50888 17572 -50854
rect 18036 -50888 18048 -50854
rect 17560 -50894 18048 -50888
rect 18280 -50978 18340 -50804
rect 19308 -50804 19314 -50252
rect 19348 -50252 19364 -50228
rect 20324 -50228 20384 -49986
rect 21336 -49986 21350 -49962
rect 21384 -49434 21396 -49410
rect 22358 -49410 22418 -49168
rect 23378 -49168 23386 -49144
rect 23420 -48622 23438 -48592
rect 24394 -48592 24454 -48350
rect 25416 -48350 25422 -47774
rect 25456 -47802 25476 -47774
rect 25456 -48332 25462 -47802
rect 25456 -48350 25476 -48332
rect 24686 -48400 25174 -48394
rect 24686 -48434 24698 -48400
rect 25162 -48434 25174 -48400
rect 24686 -48440 25174 -48434
rect 24888 -48502 24948 -48440
rect 24686 -48508 25174 -48502
rect 24686 -48542 24698 -48508
rect 25162 -48542 25174 -48508
rect 24686 -48548 25174 -48542
rect 24394 -48618 24404 -48592
rect 23420 -49144 23426 -48622
rect 24398 -49140 24404 -48618
rect 23420 -49168 23438 -49144
rect 22650 -49218 23138 -49212
rect 22650 -49252 22662 -49218
rect 23126 -49252 23138 -49218
rect 22650 -49258 23138 -49252
rect 22858 -49320 22918 -49258
rect 22650 -49326 23138 -49320
rect 22650 -49360 22662 -49326
rect 23126 -49360 23138 -49326
rect 22650 -49366 23138 -49360
rect 22358 -49434 22368 -49410
rect 21384 -49962 21390 -49434
rect 22362 -49962 22368 -49434
rect 21384 -49986 21396 -49962
rect 20614 -50036 21102 -50030
rect 20614 -50070 20626 -50036
rect 21090 -50070 21102 -50036
rect 20614 -50076 21102 -50070
rect 20822 -50138 20882 -50076
rect 20614 -50144 21102 -50138
rect 20614 -50178 20626 -50144
rect 21090 -50178 21102 -50144
rect 20614 -50184 21102 -50178
rect 20324 -50244 20332 -50228
rect 19348 -50804 19354 -50252
rect 20326 -50756 20332 -50244
rect 19308 -50816 19354 -50804
rect 20318 -50804 20332 -50756
rect 20366 -50244 20384 -50228
rect 21336 -50228 21396 -49986
rect 22358 -49986 22368 -49962
rect 22402 -49434 22418 -49410
rect 23378 -49410 23438 -49168
rect 24394 -49168 24404 -49140
rect 24438 -48618 24454 -48592
rect 25416 -48592 25476 -48350
rect 24438 -49140 24444 -48618
rect 24438 -49168 24454 -49140
rect 23668 -49218 24156 -49212
rect 23668 -49252 23680 -49218
rect 24144 -49252 24156 -49218
rect 23668 -49258 24156 -49252
rect 23870 -49320 23930 -49258
rect 23668 -49326 24156 -49320
rect 23668 -49360 23680 -49326
rect 24144 -49360 24156 -49326
rect 23668 -49366 24156 -49360
rect 23378 -49434 23386 -49410
rect 22402 -49962 22408 -49434
rect 23380 -49962 23386 -49434
rect 22402 -49986 22418 -49962
rect 21632 -50036 22120 -50030
rect 21632 -50070 21644 -50036
rect 22108 -50070 22120 -50036
rect 21632 -50076 22120 -50070
rect 21838 -50138 21898 -50076
rect 21632 -50144 22120 -50138
rect 21632 -50178 21644 -50144
rect 22108 -50178 22120 -50144
rect 21632 -50184 22120 -50178
rect 20366 -50756 20372 -50244
rect 21336 -50252 21350 -50228
rect 20366 -50804 20378 -50756
rect 18578 -50854 19066 -50848
rect 18578 -50888 18590 -50854
rect 19054 -50888 19066 -50854
rect 18578 -50894 19066 -50888
rect 19596 -50854 20084 -50848
rect 19596 -50888 19608 -50854
rect 20072 -50888 20084 -50854
rect 19596 -50894 20084 -50888
rect 20318 -50978 20378 -50804
rect 21344 -50804 21350 -50252
rect 21384 -50252 21396 -50228
rect 22358 -50228 22418 -49986
rect 23378 -49986 23386 -49962
rect 23420 -49434 23438 -49410
rect 24394 -49410 24454 -49168
rect 25416 -49168 25422 -48592
rect 25456 -48622 25476 -48592
rect 25456 -49144 25462 -48622
rect 25456 -49168 25476 -49144
rect 24686 -49218 25174 -49212
rect 24686 -49252 24698 -49218
rect 25162 -49252 25174 -49218
rect 24686 -49258 25174 -49252
rect 24890 -49320 24950 -49258
rect 24686 -49326 25174 -49320
rect 24686 -49360 24698 -49326
rect 25162 -49360 25174 -49326
rect 24686 -49366 25174 -49360
rect 24394 -49430 24404 -49410
rect 23420 -49962 23426 -49434
rect 24398 -49958 24404 -49430
rect 23420 -49986 23438 -49962
rect 22650 -50036 23138 -50030
rect 22650 -50070 22662 -50036
rect 23126 -50070 23138 -50036
rect 22650 -50076 23138 -50070
rect 22860 -50138 22920 -50076
rect 22650 -50144 23138 -50138
rect 22650 -50178 22662 -50144
rect 23126 -50178 23138 -50144
rect 22650 -50184 23138 -50178
rect 22358 -50252 22368 -50228
rect 21384 -50804 21390 -50252
rect 22362 -50760 22368 -50252
rect 21344 -50816 21390 -50804
rect 22354 -50804 22368 -50760
rect 22402 -50252 22418 -50228
rect 23378 -50228 23438 -49986
rect 24394 -49986 24404 -49958
rect 24438 -49430 24454 -49410
rect 25416 -49410 25476 -49168
rect 24438 -49958 24444 -49430
rect 24438 -49986 24454 -49958
rect 23668 -50036 24156 -50030
rect 23668 -50070 23680 -50036
rect 24144 -50070 24156 -50036
rect 23668 -50076 24156 -50070
rect 23872 -50138 23932 -50076
rect 23668 -50144 24156 -50138
rect 23668 -50178 23680 -50144
rect 24144 -50178 24156 -50144
rect 23668 -50184 24156 -50178
rect 23378 -50252 23386 -50228
rect 22402 -50760 22408 -50252
rect 22402 -50804 22414 -50760
rect 20614 -50854 21102 -50848
rect 20614 -50888 20626 -50854
rect 21090 -50888 21102 -50854
rect 20614 -50894 21102 -50888
rect 21632 -50854 22120 -50848
rect 21632 -50888 21644 -50854
rect 22108 -50888 22120 -50854
rect 21632 -50894 22120 -50888
rect 22354 -50978 22414 -50804
rect 23380 -50804 23386 -50252
rect 23420 -50252 23438 -50228
rect 24394 -50228 24454 -49986
rect 25416 -49986 25422 -49410
rect 25456 -49434 25476 -49410
rect 25456 -49962 25462 -49434
rect 25456 -49986 25476 -49962
rect 24686 -50036 25174 -50030
rect 24686 -50070 24698 -50036
rect 25162 -50070 25174 -50036
rect 24686 -50076 25174 -50070
rect 24892 -50138 24952 -50076
rect 24686 -50144 25174 -50138
rect 24686 -50178 24698 -50144
rect 25162 -50178 25174 -50144
rect 24686 -50184 25174 -50178
rect 24394 -50248 24404 -50228
rect 23420 -50804 23426 -50252
rect 24398 -50762 24404 -50248
rect 23380 -50816 23426 -50804
rect 24390 -50804 24404 -50762
rect 24438 -50248 24454 -50228
rect 25416 -50228 25476 -49986
rect 24438 -50762 24444 -50248
rect 25416 -50750 25422 -50228
rect 24438 -50804 24450 -50762
rect 22650 -50854 23138 -50848
rect 22650 -50888 22662 -50854
rect 23126 -50888 23138 -50854
rect 22650 -50894 23138 -50888
rect 23668 -50854 24156 -50848
rect 23668 -50888 23680 -50854
rect 24144 -50888 24156 -50854
rect 23668 -50894 24156 -50888
rect 24390 -50978 24450 -50804
rect 25410 -50804 25422 -50750
rect 25456 -50252 25476 -50228
rect 25456 -50750 25462 -50252
rect 25456 -50804 25470 -50750
rect 26594 -50800 26654 -43660
rect 24686 -50854 25174 -50848
rect 24686 -50888 24698 -50854
rect 25162 -50888 25174 -50854
rect 24686 -50894 25174 -50888
rect 24904 -50978 24964 -50894
rect 25410 -50978 25470 -50804
rect 26588 -50860 26594 -50800
rect 26654 -50860 26660 -50800
rect 18280 -51038 26574 -50978
rect 22040 -51786 22046 -51726
rect 22106 -51786 22112 -51726
rect 15936 -51872 15996 -51866
rect 20010 -51932 20016 -51872
rect 20076 -51932 20082 -51872
rect 14776 -52060 14782 -52000
rect 14842 -52060 14848 -52000
rect 14782 -52942 14842 -52060
rect 15936 -52064 15996 -51932
rect 17454 -52060 17460 -52000
rect 17520 -52060 17526 -52000
rect 18486 -52060 18492 -52000
rect 18552 -52060 18558 -52000
rect 14920 -52124 15996 -52064
rect 14920 -52252 14980 -52124
rect 15428 -52162 15488 -52124
rect 15218 -52168 15706 -52162
rect 15218 -52202 15230 -52168
rect 15694 -52202 15706 -52168
rect 15218 -52208 15706 -52202
rect 14920 -52298 14936 -52252
rect 14930 -52828 14936 -52298
rect 14970 -52298 14980 -52252
rect 15936 -52252 15996 -52124
rect 17460 -52162 17520 -52060
rect 18492 -52162 18552 -52060
rect 16236 -52168 16724 -52162
rect 16236 -52202 16248 -52168
rect 16712 -52202 16724 -52168
rect 16236 -52208 16724 -52202
rect 17254 -52168 17742 -52162
rect 17254 -52202 17266 -52168
rect 17730 -52202 17742 -52168
rect 17254 -52208 17742 -52202
rect 18272 -52168 18760 -52162
rect 18272 -52202 18284 -52168
rect 18748 -52202 18760 -52168
rect 18272 -52208 18760 -52202
rect 19290 -52168 19778 -52162
rect 19290 -52202 19302 -52168
rect 19766 -52202 19778 -52168
rect 19290 -52208 19778 -52202
rect 15936 -52292 15954 -52252
rect 14970 -52828 14976 -52298
rect 14930 -52840 14976 -52828
rect 15948 -52828 15954 -52292
rect 15988 -52292 15996 -52252
rect 16966 -52252 17012 -52240
rect 15988 -52828 15994 -52292
rect 16966 -52764 16972 -52252
rect 15948 -52840 15994 -52828
rect 16958 -52828 16972 -52764
rect 17006 -52764 17012 -52252
rect 17984 -52252 18030 -52240
rect 17006 -52828 17018 -52764
rect 17984 -52782 17990 -52252
rect 15218 -52878 15706 -52872
rect 15218 -52912 15230 -52878
rect 15694 -52912 15706 -52878
rect 15218 -52918 15706 -52912
rect 16236 -52878 16724 -52872
rect 16236 -52912 16248 -52878
rect 16712 -52912 16724 -52878
rect 16236 -52918 16724 -52912
rect 14762 -52948 14862 -52942
rect 16440 -52962 16500 -52918
rect 16434 -53022 16440 -52962
rect 16500 -53022 16506 -52962
rect 14762 -53054 14862 -53048
rect 14782 -53936 14842 -53054
rect 15934 -53126 15940 -53066
rect 16000 -53126 16006 -53066
rect 15940 -53168 16000 -53126
rect 14920 -53228 16000 -53168
rect 14920 -53364 14980 -53228
rect 15424 -53274 15484 -53228
rect 15218 -53280 15706 -53274
rect 15218 -53314 15230 -53280
rect 15694 -53314 15706 -53280
rect 15218 -53320 15706 -53314
rect 14920 -53410 14936 -53364
rect 14764 -53942 14864 -53936
rect 14930 -53940 14936 -53410
rect 14970 -53410 14980 -53364
rect 15940 -53364 16000 -53228
rect 16958 -53170 17018 -52828
rect 17976 -52828 17990 -52782
rect 18024 -52782 18030 -52252
rect 19002 -52252 19048 -52240
rect 19002 -52766 19008 -52252
rect 18024 -52828 18036 -52782
rect 17254 -52878 17742 -52872
rect 17254 -52912 17266 -52878
rect 17730 -52912 17742 -52878
rect 17254 -52918 17742 -52912
rect 17458 -53022 17464 -52962
rect 17524 -53022 17530 -52962
rect 16236 -53280 16724 -53274
rect 16236 -53314 16248 -53280
rect 16712 -53314 16724 -53280
rect 16236 -53320 16724 -53314
rect 14970 -53940 14976 -53410
rect 14930 -53952 14976 -53940
rect 15940 -53940 15954 -53364
rect 15988 -53940 16000 -53364
rect 15218 -53990 15706 -53984
rect 15218 -54024 15230 -53990
rect 15694 -54024 15706 -53990
rect 15218 -54030 15706 -54024
rect 14764 -54048 14864 -54042
rect 14782 -54232 14842 -54048
rect 14776 -54292 14782 -54232
rect 14842 -54292 14848 -54232
rect 14782 -54942 14842 -54292
rect 15218 -54392 15706 -54386
rect 15218 -54426 15230 -54392
rect 15694 -54426 15706 -54392
rect 15218 -54432 15706 -54426
rect 14930 -54476 14976 -54464
rect 14764 -54948 14864 -54942
rect 14930 -55018 14936 -54476
rect 14764 -55054 14864 -55048
rect 14924 -55052 14936 -55018
rect 14970 -55018 14976 -54476
rect 15940 -54476 16000 -53940
rect 16958 -53364 17018 -53230
rect 17464 -53274 17524 -53022
rect 17976 -53066 18036 -52828
rect 18994 -52828 19008 -52766
rect 19042 -52766 19048 -52252
rect 20016 -52252 20076 -51932
rect 21546 -52060 21552 -52000
rect 21612 -52060 21618 -52000
rect 21552 -52162 21612 -52060
rect 20308 -52168 20796 -52162
rect 20308 -52202 20320 -52168
rect 20784 -52202 20796 -52168
rect 20308 -52208 20796 -52202
rect 21326 -52168 21814 -52162
rect 21326 -52202 21338 -52168
rect 21802 -52202 21814 -52168
rect 21326 -52208 21814 -52202
rect 20016 -52316 20026 -52252
rect 19042 -52828 19054 -52766
rect 18272 -52878 18760 -52872
rect 18272 -52912 18284 -52878
rect 18748 -52912 18760 -52878
rect 18272 -52918 18760 -52912
rect 18490 -53022 18496 -52962
rect 18556 -53022 18562 -52962
rect 17970 -53126 17976 -53066
rect 18036 -53126 18042 -53066
rect 18496 -53274 18556 -53022
rect 18994 -53170 19054 -52828
rect 20020 -52828 20026 -52316
rect 20060 -52316 20076 -52252
rect 21038 -52252 21084 -52240
rect 20060 -52828 20066 -52316
rect 21038 -52756 21044 -52252
rect 20020 -52840 20066 -52828
rect 21026 -52828 21044 -52756
rect 21078 -52756 21084 -52252
rect 22046 -52252 22106 -51786
rect 24070 -51932 24076 -51872
rect 24136 -51932 24142 -51872
rect 26254 -51932 26260 -51872
rect 26320 -51932 26326 -51872
rect 22542 -52060 22548 -52000
rect 22608 -52060 22614 -52000
rect 22548 -52162 22608 -52060
rect 22344 -52168 22832 -52162
rect 22344 -52202 22356 -52168
rect 22820 -52202 22832 -52168
rect 22344 -52208 22832 -52202
rect 23362 -52168 23850 -52162
rect 23362 -52202 23374 -52168
rect 23838 -52202 23850 -52168
rect 23362 -52208 23850 -52202
rect 22548 -52210 22608 -52208
rect 24076 -52240 24136 -51932
rect 24380 -52168 24868 -52162
rect 24380 -52202 24392 -52168
rect 24856 -52202 24868 -52168
rect 24380 -52208 24868 -52202
rect 25398 -52168 25886 -52162
rect 25398 -52202 25410 -52168
rect 25874 -52202 25886 -52168
rect 25398 -52208 25886 -52202
rect 21078 -52828 21086 -52756
rect 19290 -52878 19778 -52872
rect 19290 -52912 19302 -52878
rect 19766 -52912 19778 -52878
rect 19290 -52918 19778 -52912
rect 20308 -52878 20796 -52872
rect 20308 -52912 20320 -52878
rect 20784 -52912 20796 -52878
rect 20308 -52918 20796 -52912
rect 19496 -52962 19556 -52918
rect 20516 -52962 20576 -52918
rect 19490 -53022 19496 -52962
rect 19556 -53022 19562 -52962
rect 20510 -53022 20516 -52962
rect 20576 -53022 20582 -52962
rect 20006 -53126 20012 -53066
rect 20072 -53126 20078 -53066
rect 17254 -53280 17742 -53274
rect 17254 -53314 17266 -53280
rect 17730 -53314 17742 -53280
rect 17254 -53320 17742 -53314
rect 18272 -53280 18760 -53274
rect 18272 -53314 18284 -53280
rect 18748 -53314 18760 -53280
rect 18272 -53320 18760 -53314
rect 16958 -53940 16972 -53364
rect 17006 -53940 17018 -53364
rect 17984 -53364 18030 -53352
rect 17984 -53902 17990 -53364
rect 16236 -53990 16724 -53984
rect 16236 -54024 16248 -53990
rect 16712 -54024 16724 -53990
rect 16236 -54030 16724 -54024
rect 16432 -54232 16492 -54030
rect 16426 -54292 16432 -54232
rect 16492 -54292 16498 -54232
rect 16432 -54386 16492 -54292
rect 16236 -54392 16724 -54386
rect 16236 -54426 16248 -54392
rect 16712 -54426 16724 -54392
rect 16236 -54432 16724 -54426
rect 15940 -54548 15954 -54476
rect 14970 -55052 14984 -55018
rect 15948 -55022 15954 -54548
rect 14782 -56358 14842 -55054
rect 14924 -55184 14984 -55052
rect 15944 -55052 15954 -55022
rect 15988 -54548 16000 -54476
rect 16958 -54476 17018 -53940
rect 17970 -53940 17990 -53902
rect 18024 -53940 18030 -53364
rect 17254 -53990 17742 -53984
rect 17254 -54024 17266 -53990
rect 17730 -54024 17742 -53990
rect 17254 -54030 17742 -54024
rect 17970 -54112 18030 -53940
rect 18994 -53364 19054 -53230
rect 19290 -53280 19778 -53274
rect 19290 -53314 19302 -53280
rect 19766 -53314 19778 -53280
rect 19290 -53320 19778 -53314
rect 18994 -53940 19008 -53364
rect 19042 -53940 19054 -53364
rect 18272 -53990 18760 -53984
rect 18272 -54024 18284 -53990
rect 18748 -54024 18760 -53990
rect 18272 -54030 18760 -54024
rect 17964 -54172 17970 -54112
rect 18030 -54172 18036 -54112
rect 17254 -54392 17742 -54386
rect 17254 -54426 17266 -54392
rect 17730 -54426 17742 -54392
rect 17254 -54432 17742 -54426
rect 15988 -55022 15994 -54548
rect 15988 -55052 16004 -55022
rect 15218 -55102 15706 -55096
rect 15218 -55136 15230 -55102
rect 15694 -55136 15706 -55102
rect 15218 -55142 15706 -55136
rect 15416 -55184 15476 -55142
rect 15944 -55184 16004 -55052
rect 16958 -55052 16972 -54476
rect 17006 -55052 17018 -54476
rect 17970 -54476 18030 -54172
rect 18272 -54392 18760 -54386
rect 18272 -54426 18284 -54392
rect 18748 -54426 18760 -54392
rect 18272 -54432 18760 -54426
rect 17970 -54546 17990 -54476
rect 16236 -55102 16724 -55096
rect 16236 -55136 16248 -55102
rect 16712 -55136 16724 -55102
rect 16236 -55142 16724 -55136
rect 14924 -55244 16004 -55184
rect 15944 -55284 16004 -55244
rect 16958 -55176 17018 -55052
rect 17984 -55052 17990 -54546
rect 18024 -55052 18030 -54476
rect 17984 -55064 18030 -55052
rect 18994 -54476 19054 -53940
rect 20012 -53364 20072 -53126
rect 21026 -53170 21086 -52828
rect 22046 -52828 22062 -52252
rect 22096 -52828 22106 -52252
rect 23074 -52252 23120 -52240
rect 23074 -52766 23080 -52252
rect 21326 -52878 21814 -52872
rect 21326 -52912 21338 -52878
rect 21802 -52912 21814 -52878
rect 21326 -52918 21814 -52912
rect 21530 -53022 21536 -52962
rect 21596 -53022 21602 -52962
rect 21020 -53230 21026 -53170
rect 21086 -53230 21092 -53170
rect 20308 -53280 20796 -53274
rect 20308 -53314 20320 -53280
rect 20784 -53314 20796 -53280
rect 20308 -53320 20796 -53314
rect 20012 -53940 20026 -53364
rect 20060 -53940 20072 -53364
rect 19290 -53990 19778 -53984
rect 19290 -54024 19302 -53990
rect 19766 -54024 19778 -53990
rect 19290 -54030 19778 -54024
rect 19502 -54232 19562 -54030
rect 19496 -54292 19502 -54232
rect 19562 -54292 19568 -54232
rect 19502 -54386 19562 -54292
rect 19290 -54392 19778 -54386
rect 19290 -54426 19302 -54392
rect 19766 -54426 19778 -54392
rect 19290 -54432 19778 -54426
rect 18994 -55052 19008 -54476
rect 19042 -55052 19054 -54476
rect 20012 -54476 20072 -53940
rect 21026 -53364 21086 -53230
rect 21536 -53274 21596 -53022
rect 22046 -53066 22106 -52828
rect 23060 -52828 23080 -52766
rect 23114 -52828 23120 -52252
rect 24076 -52252 24138 -52240
rect 24076 -52284 24098 -52252
rect 22344 -52878 22832 -52872
rect 22344 -52912 22356 -52878
rect 22820 -52912 22832 -52878
rect 22344 -52918 22832 -52912
rect 22546 -52962 22606 -52956
rect 22040 -53126 22046 -53066
rect 22106 -53126 22112 -53066
rect 22546 -53274 22606 -53022
rect 23060 -53170 23120 -52828
rect 24092 -52828 24098 -52284
rect 24132 -52828 24138 -52252
rect 25110 -52252 25156 -52240
rect 25110 -52794 25116 -52252
rect 24092 -52840 24138 -52828
rect 25104 -52828 25116 -52794
rect 25150 -52794 25156 -52252
rect 26128 -52252 26174 -52240
rect 26128 -52774 26134 -52252
rect 25150 -52828 25164 -52794
rect 23362 -52878 23850 -52872
rect 23362 -52912 23374 -52878
rect 23838 -52912 23850 -52878
rect 23362 -52918 23850 -52912
rect 24380 -52878 24868 -52872
rect 24380 -52912 24392 -52878
rect 24856 -52912 24868 -52878
rect 24380 -52918 24868 -52912
rect 23560 -52962 23620 -52918
rect 24578 -52962 24638 -52918
rect 23554 -53022 23560 -52962
rect 23620 -53022 23626 -52962
rect 24578 -53028 24638 -53022
rect 25104 -53056 25164 -52828
rect 26120 -52828 26134 -52774
rect 26168 -52774 26174 -52252
rect 26168 -52828 26180 -52774
rect 25398 -52878 25886 -52872
rect 25398 -52912 25410 -52878
rect 25874 -52912 25886 -52878
rect 25398 -52918 25886 -52912
rect 25608 -53056 25668 -52918
rect 26120 -53056 26180 -52828
rect 24076 -53126 24082 -53066
rect 24142 -53126 24148 -53066
rect 25104 -53116 26180 -53056
rect 21326 -53280 21814 -53274
rect 21326 -53314 21338 -53280
rect 21802 -53314 21814 -53280
rect 21326 -53320 21814 -53314
rect 22344 -53280 22832 -53274
rect 22344 -53314 22356 -53280
rect 22820 -53314 22832 -53280
rect 22344 -53320 22832 -53314
rect 21026 -53940 21044 -53364
rect 21078 -53940 21086 -53364
rect 22056 -53364 22102 -53352
rect 22056 -53884 22062 -53364
rect 20308 -53990 20796 -53984
rect 20308 -54024 20320 -53990
rect 20784 -54024 20796 -53990
rect 20308 -54030 20796 -54024
rect 20510 -54232 20570 -54030
rect 20504 -54292 20510 -54232
rect 20570 -54292 20576 -54232
rect 20510 -54386 20570 -54292
rect 20308 -54392 20796 -54386
rect 20308 -54426 20320 -54392
rect 20784 -54426 20796 -54392
rect 20308 -54432 20796 -54426
rect 20012 -54582 20026 -54476
rect 20020 -54990 20026 -54582
rect 17254 -55102 17742 -55096
rect 17254 -55136 17266 -55102
rect 17730 -55136 17742 -55102
rect 17254 -55142 17742 -55136
rect 18272 -55102 18760 -55096
rect 18272 -55136 18284 -55102
rect 18748 -55136 18760 -55102
rect 18272 -55142 18760 -55136
rect 15938 -55344 15944 -55284
rect 16004 -55344 16010 -55284
rect 16432 -55456 16438 -55396
rect 16498 -55456 16504 -55396
rect 16438 -55498 16498 -55456
rect 15218 -55504 15706 -55498
rect 15218 -55538 15230 -55504
rect 15694 -55538 15706 -55504
rect 15218 -55544 15706 -55538
rect 16236 -55504 16724 -55498
rect 16236 -55538 16248 -55504
rect 16712 -55538 16724 -55504
rect 16236 -55544 16724 -55538
rect 14930 -55588 14976 -55576
rect 14930 -56122 14936 -55588
rect 14920 -56164 14936 -56122
rect 14970 -56122 14976 -55588
rect 15948 -55588 15994 -55576
rect 14970 -56164 14980 -56122
rect 15948 -56128 15954 -55588
rect 14920 -56308 14980 -56164
rect 15938 -56164 15954 -56128
rect 15988 -56128 15994 -55588
rect 16958 -55588 17018 -55236
rect 17462 -55396 17522 -55142
rect 17974 -55344 17980 -55284
rect 18040 -55344 18046 -55284
rect 17456 -55456 17462 -55396
rect 17522 -55456 17528 -55396
rect 17254 -55504 17742 -55498
rect 17254 -55538 17266 -55504
rect 17730 -55538 17742 -55504
rect 17254 -55544 17742 -55538
rect 16958 -55690 16972 -55588
rect 15988 -56164 15998 -56128
rect 15218 -56214 15706 -56208
rect 15218 -56248 15230 -56214
rect 15694 -56248 15706 -56214
rect 15218 -56254 15706 -56248
rect 15424 -56308 15484 -56254
rect 15938 -56308 15998 -56164
rect 16966 -56164 16972 -55690
rect 17006 -55690 17018 -55588
rect 17980 -55588 18040 -55344
rect 18494 -55396 18554 -55142
rect 18994 -55176 19054 -55052
rect 20016 -55052 20026 -54990
rect 20060 -54582 20072 -54476
rect 21026 -54476 21086 -53940
rect 22046 -53940 22062 -53884
rect 22096 -53884 22102 -53364
rect 23060 -53364 23120 -53230
rect 23362 -53280 23850 -53274
rect 23362 -53314 23374 -53280
rect 23838 -53314 23850 -53280
rect 23362 -53320 23850 -53314
rect 22096 -53940 22106 -53884
rect 21326 -53990 21814 -53984
rect 21326 -54024 21338 -53990
rect 21802 -54024 21814 -53990
rect 21326 -54030 21814 -54024
rect 22046 -54112 22106 -53940
rect 23060 -53940 23080 -53364
rect 23114 -53940 23120 -53364
rect 22344 -53990 22832 -53984
rect 22344 -54024 22356 -53990
rect 22820 -54024 22832 -53990
rect 22344 -54030 22832 -54024
rect 22040 -54172 22046 -54112
rect 22106 -54172 22112 -54112
rect 21326 -54392 21814 -54386
rect 21326 -54426 21338 -54392
rect 21802 -54426 21814 -54392
rect 21326 -54432 21814 -54426
rect 20060 -54990 20066 -54582
rect 20060 -55052 20076 -54990
rect 19290 -55102 19778 -55096
rect 19290 -55136 19302 -55102
rect 19766 -55136 19778 -55102
rect 19290 -55142 19778 -55136
rect 18488 -55456 18494 -55396
rect 18554 -55456 18560 -55396
rect 18272 -55504 18760 -55498
rect 18272 -55538 18284 -55504
rect 18748 -55538 18760 -55504
rect 18272 -55544 18760 -55538
rect 17980 -55628 17990 -55588
rect 17006 -56164 17012 -55690
rect 16966 -56176 17012 -56164
rect 17984 -56164 17990 -55628
rect 18024 -55628 18040 -55588
rect 18994 -55588 19054 -55236
rect 20016 -55284 20076 -55052
rect 21026 -55052 21044 -54476
rect 21078 -55052 21086 -54476
rect 22046 -54476 22106 -54172
rect 22344 -54392 22832 -54386
rect 22344 -54426 22356 -54392
rect 22820 -54426 22832 -54392
rect 22344 -54432 22832 -54426
rect 22046 -54518 22062 -54476
rect 20308 -55102 20796 -55096
rect 20308 -55136 20320 -55102
rect 20784 -55136 20796 -55102
rect 20308 -55142 20796 -55136
rect 21026 -55176 21086 -55052
rect 22056 -55052 22062 -54518
rect 22096 -54518 22106 -54476
rect 23060 -54476 23120 -53940
rect 24082 -53364 24142 -53126
rect 25104 -53170 25164 -53116
rect 24380 -53280 24868 -53274
rect 24380 -53314 24392 -53280
rect 24856 -53314 24868 -53280
rect 24380 -53320 24868 -53314
rect 24082 -53940 24098 -53364
rect 24132 -53940 24142 -53364
rect 23362 -53990 23850 -53984
rect 23362 -54024 23374 -53990
rect 23838 -54024 23850 -53990
rect 23362 -54030 23850 -54024
rect 23572 -54232 23632 -54030
rect 23566 -54292 23572 -54232
rect 23632 -54292 23638 -54232
rect 23572 -54386 23632 -54292
rect 23362 -54392 23850 -54386
rect 23362 -54426 23374 -54392
rect 23838 -54426 23850 -54392
rect 23362 -54432 23850 -54426
rect 22096 -55052 22102 -54518
rect 22056 -55064 22102 -55052
rect 23060 -55052 23080 -54476
rect 23114 -55052 23120 -54476
rect 24082 -54476 24142 -53940
rect 25104 -53364 25164 -53230
rect 25608 -53274 25668 -53116
rect 25398 -53280 25886 -53274
rect 25398 -53314 25410 -53280
rect 25874 -53314 25886 -53280
rect 25398 -53320 25886 -53314
rect 25104 -53940 25116 -53364
rect 25150 -53940 25164 -53364
rect 24380 -53990 24868 -53984
rect 24380 -54024 24392 -53990
rect 24856 -54024 24868 -53990
rect 24380 -54030 24868 -54024
rect 24598 -54232 24658 -54030
rect 25104 -54176 25164 -53940
rect 26120 -53364 26180 -53116
rect 26120 -53940 26134 -53364
rect 26168 -53940 26180 -53364
rect 25398 -53990 25886 -53984
rect 25398 -54024 25410 -53990
rect 25874 -54024 25886 -53990
rect 25398 -54030 25886 -54024
rect 25604 -54176 25664 -54030
rect 26120 -54176 26180 -53940
rect 26260 -54112 26320 -51932
rect 26374 -53022 26380 -52962
rect 26440 -53022 26446 -52962
rect 26380 -53564 26440 -53022
rect 26374 -53624 26380 -53564
rect 26440 -53624 26446 -53564
rect 26254 -54172 26260 -54112
rect 26320 -54172 26326 -54112
rect 24592 -54292 24598 -54232
rect 24658 -54292 24664 -54232
rect 25104 -54236 26180 -54176
rect 24598 -54386 24658 -54292
rect 24380 -54392 24868 -54386
rect 24380 -54426 24392 -54392
rect 24856 -54426 24868 -54392
rect 24380 -54432 24868 -54426
rect 24082 -54532 24098 -54476
rect 24092 -55006 24098 -54532
rect 21326 -55102 21814 -55096
rect 21326 -55136 21338 -55102
rect 21802 -55136 21814 -55102
rect 21326 -55142 21814 -55136
rect 22344 -55102 22832 -55096
rect 22344 -55136 22356 -55102
rect 22820 -55136 22832 -55102
rect 22344 -55142 22832 -55136
rect 20010 -55344 20016 -55284
rect 20076 -55344 20082 -55284
rect 19488 -55456 19494 -55396
rect 19554 -55456 19560 -55396
rect 20508 -55456 20514 -55396
rect 20574 -55456 20580 -55396
rect 19494 -55498 19554 -55456
rect 20514 -55498 20574 -55456
rect 19290 -55504 19778 -55498
rect 19290 -55538 19302 -55504
rect 19766 -55538 19778 -55504
rect 19290 -55544 19778 -55538
rect 20308 -55504 20796 -55498
rect 20308 -55538 20320 -55504
rect 20784 -55538 20796 -55504
rect 20308 -55544 20796 -55538
rect 18994 -55626 19008 -55588
rect 18024 -56164 18030 -55628
rect 17984 -56176 18030 -56164
rect 19002 -56164 19008 -55626
rect 19042 -55626 19054 -55588
rect 20020 -55588 20066 -55576
rect 19042 -56164 19048 -55626
rect 20020 -56104 20026 -55588
rect 19002 -56176 19048 -56164
rect 20018 -56164 20026 -56104
rect 20060 -56104 20066 -55588
rect 21026 -55588 21086 -55236
rect 21534 -55396 21594 -55142
rect 22044 -55344 22050 -55284
rect 22110 -55344 22116 -55284
rect 21528 -55456 21534 -55396
rect 21594 -55456 21600 -55396
rect 21326 -55504 21814 -55498
rect 21326 -55538 21338 -55504
rect 21802 -55538 21814 -55504
rect 21326 -55544 21814 -55538
rect 21026 -55648 21044 -55588
rect 20060 -56164 20078 -56104
rect 16236 -56214 16724 -56208
rect 16236 -56248 16248 -56214
rect 16712 -56248 16724 -56214
rect 16236 -56254 16724 -56248
rect 17254 -56214 17742 -56208
rect 17254 -56248 17266 -56214
rect 17730 -56248 17742 -56214
rect 17254 -56254 17742 -56248
rect 18272 -56214 18760 -56208
rect 18272 -56248 18284 -56214
rect 18748 -56248 18760 -56214
rect 18272 -56254 18760 -56248
rect 19290 -56214 19778 -56208
rect 19290 -56248 19302 -56214
rect 19766 -56248 19778 -56214
rect 19290 -56254 19778 -56248
rect 14776 -56418 14782 -56358
rect 14842 -56418 14848 -56358
rect 14920 -56368 15998 -56308
rect 17452 -56358 17512 -56254
rect 18484 -56358 18544 -56254
rect 15938 -56488 15998 -56368
rect 17446 -56418 17452 -56358
rect 17512 -56418 17518 -56358
rect 18478 -56418 18484 -56358
rect 18544 -56418 18550 -56358
rect 20018 -56488 20078 -56164
rect 21038 -56164 21044 -55648
rect 21078 -55648 21086 -55588
rect 22050 -55588 22110 -55344
rect 22544 -55396 22604 -55142
rect 22544 -55462 22604 -55456
rect 23060 -55176 23120 -55052
rect 24086 -55052 24098 -55006
rect 24132 -54532 24142 -54476
rect 25104 -54476 25164 -54236
rect 25604 -54386 25664 -54236
rect 25398 -54392 25886 -54386
rect 25398 -54426 25410 -54392
rect 25874 -54426 25886 -54392
rect 25398 -54432 25886 -54426
rect 24132 -55006 24138 -54532
rect 24132 -55052 24146 -55006
rect 23362 -55102 23850 -55096
rect 23362 -55136 23374 -55102
rect 23838 -55136 23850 -55102
rect 23362 -55142 23850 -55136
rect 22344 -55504 22832 -55498
rect 22344 -55538 22356 -55504
rect 22820 -55538 22832 -55504
rect 22344 -55544 22832 -55538
rect 22050 -55634 22062 -55588
rect 21078 -56164 21084 -55648
rect 21038 -56176 21084 -56164
rect 22056 -56164 22062 -55634
rect 22096 -55634 22110 -55588
rect 23060 -55588 23120 -55236
rect 24086 -55284 24146 -55052
rect 25104 -55052 25116 -54476
rect 25150 -55052 25164 -54476
rect 24380 -55102 24868 -55096
rect 24380 -55136 24392 -55102
rect 24856 -55136 24868 -55102
rect 24380 -55142 24868 -55136
rect 25104 -55176 25164 -55052
rect 26120 -54476 26180 -54236
rect 26120 -55052 26134 -54476
rect 26168 -55052 26180 -54476
rect 25398 -55102 25886 -55096
rect 25398 -55136 25410 -55102
rect 25874 -55136 25886 -55102
rect 25398 -55142 25886 -55136
rect 25098 -55236 25104 -55176
rect 25164 -55236 25170 -55176
rect 24080 -55344 24086 -55284
rect 24146 -55344 24152 -55284
rect 25104 -55288 25164 -55236
rect 25612 -55288 25672 -55142
rect 26120 -55288 26180 -55052
rect 25104 -55348 26180 -55288
rect 24576 -55396 24636 -55390
rect 23552 -55456 23558 -55396
rect 23618 -55456 23624 -55396
rect 23558 -55498 23618 -55456
rect 24576 -55498 24636 -55456
rect 23362 -55504 23850 -55498
rect 23362 -55538 23374 -55504
rect 23838 -55538 23850 -55504
rect 23362 -55544 23850 -55538
rect 24380 -55504 24868 -55498
rect 24380 -55538 24392 -55504
rect 24856 -55538 24868 -55504
rect 24380 -55544 24868 -55538
rect 23060 -55630 23080 -55588
rect 22096 -56164 22102 -55634
rect 22056 -56176 22102 -56164
rect 23074 -56164 23080 -55630
rect 23114 -56164 23120 -55588
rect 24092 -55588 24138 -55576
rect 24092 -56136 24098 -55588
rect 23074 -56176 23120 -56164
rect 24078 -56164 24098 -56136
rect 24132 -56164 24138 -55588
rect 25104 -55588 25164 -55348
rect 25612 -55498 25672 -55348
rect 25398 -55504 25886 -55498
rect 25398 -55538 25410 -55504
rect 25874 -55538 25886 -55504
rect 25398 -55544 25886 -55538
rect 25104 -55652 25116 -55588
rect 20308 -56214 20796 -56208
rect 20308 -56248 20320 -56214
rect 20784 -56248 20796 -56214
rect 20308 -56254 20796 -56248
rect 21326 -56214 21814 -56208
rect 21326 -56248 21338 -56214
rect 21802 -56248 21814 -56214
rect 21326 -56254 21814 -56248
rect 22344 -56214 22832 -56208
rect 22344 -56248 22356 -56214
rect 22820 -56248 22832 -56214
rect 22344 -56254 22832 -56248
rect 23362 -56214 23850 -56208
rect 23362 -56248 23374 -56214
rect 23838 -56248 23850 -56214
rect 23362 -56254 23850 -56248
rect 21544 -56358 21604 -56254
rect 22540 -56358 22600 -56254
rect 21538 -56418 21544 -56358
rect 21604 -56418 21610 -56358
rect 22534 -56418 22540 -56358
rect 22600 -56418 22606 -56358
rect 24078 -56488 24138 -56164
rect 25110 -56164 25116 -55652
rect 25150 -55652 25164 -55588
rect 26120 -55588 26180 -55348
rect 26120 -55630 26134 -55588
rect 25150 -56164 25156 -55652
rect 25110 -56176 25156 -56164
rect 26128 -56164 26134 -55630
rect 26168 -55630 26180 -55588
rect 26168 -56164 26174 -55630
rect 26128 -56176 26174 -56164
rect 24380 -56214 24868 -56208
rect 24380 -56248 24392 -56214
rect 24856 -56248 24868 -56214
rect 24380 -56254 24868 -56248
rect 25398 -56214 25886 -56208
rect 25398 -56248 25410 -56214
rect 25874 -56248 25886 -56214
rect 25398 -56254 25886 -56248
rect 26260 -56488 26320 -54172
rect 26380 -55396 26440 -53624
rect 26374 -55456 26380 -55396
rect 26440 -55456 26446 -55396
rect 20012 -56548 20018 -56488
rect 20078 -56548 20084 -56488
rect 24072 -56548 24078 -56488
rect 24138 -56548 24144 -56488
rect 26254 -56548 26260 -56488
rect 26320 -56548 26326 -56488
rect 15938 -56554 15998 -56548
rect 15194 -56954 25616 -56894
rect 15380 -57130 15440 -56954
rect 15880 -57040 15940 -56954
rect 15676 -57046 16164 -57040
rect 15676 -57080 15688 -57046
rect 16152 -57080 16164 -57046
rect 15676 -57086 16164 -57080
rect 15380 -57164 15394 -57130
rect 15388 -57706 15394 -57164
rect 15428 -57164 15440 -57130
rect 16402 -57130 16462 -56954
rect 16900 -57040 16960 -56954
rect 17934 -57040 17994 -56954
rect 18956 -57040 19016 -56954
rect 19946 -57040 20006 -56954
rect 16694 -57046 17182 -57040
rect 16694 -57080 16706 -57046
rect 17170 -57080 17182 -57046
rect 16694 -57086 17182 -57080
rect 17712 -57046 18200 -57040
rect 17712 -57080 17724 -57046
rect 18188 -57080 18200 -57046
rect 17712 -57086 18200 -57080
rect 18730 -57046 19218 -57040
rect 18730 -57080 18742 -57046
rect 19206 -57080 19218 -57046
rect 18730 -57086 19218 -57080
rect 19748 -57046 20236 -57040
rect 19748 -57080 19760 -57046
rect 20224 -57080 20236 -57046
rect 19748 -57086 20236 -57080
rect 15428 -57706 15434 -57164
rect 16402 -57174 16412 -57130
rect 15388 -57718 15434 -57706
rect 16406 -57706 16412 -57174
rect 16446 -57174 16462 -57130
rect 17424 -57130 17470 -57118
rect 16446 -57706 16452 -57174
rect 17424 -57648 17430 -57130
rect 16406 -57718 16452 -57706
rect 17416 -57706 17430 -57648
rect 17464 -57648 17470 -57130
rect 18442 -57130 18488 -57118
rect 17464 -57706 17476 -57648
rect 18442 -57672 18448 -57130
rect 15676 -57756 16164 -57750
rect 15676 -57790 15688 -57756
rect 16152 -57790 16164 -57756
rect 15676 -57796 16164 -57790
rect 16694 -57756 17182 -57750
rect 16694 -57790 16706 -57756
rect 17170 -57790 17182 -57756
rect 16694 -57796 17182 -57790
rect 17416 -57854 17476 -57706
rect 18434 -57706 18448 -57672
rect 18482 -57672 18488 -57130
rect 19460 -57130 19506 -57118
rect 19460 -57660 19466 -57130
rect 18482 -57706 18494 -57672
rect 17712 -57756 18200 -57750
rect 17712 -57790 17724 -57756
rect 18188 -57790 18200 -57756
rect 17712 -57796 18200 -57790
rect 17410 -57914 17416 -57854
rect 17476 -57914 17482 -57854
rect 10276 -58408 12130 -58390
rect 10276 -58514 10294 -58408
rect 12110 -58514 12130 -58408
rect 10276 -58528 12130 -58514
rect 13116 -59094 13228 -58308
rect 17416 -58408 17476 -57914
rect 18434 -57966 18494 -57706
rect 19454 -57706 19466 -57660
rect 19500 -57660 19506 -57130
rect 20470 -57130 20530 -56954
rect 20980 -57040 21040 -56954
rect 21970 -57040 22030 -56954
rect 23002 -57040 23062 -56954
rect 24006 -57040 24066 -56954
rect 20766 -57046 21254 -57040
rect 20766 -57080 20778 -57046
rect 21242 -57080 21254 -57046
rect 20766 -57086 21254 -57080
rect 21784 -57046 22272 -57040
rect 21784 -57080 21796 -57046
rect 22260 -57080 22272 -57046
rect 21784 -57086 22272 -57080
rect 22802 -57046 23290 -57040
rect 22802 -57080 22814 -57046
rect 23278 -57080 23290 -57046
rect 22802 -57086 23290 -57080
rect 23820 -57046 24308 -57040
rect 23820 -57080 23832 -57046
rect 24296 -57080 24308 -57046
rect 23820 -57086 24308 -57080
rect 20980 -57088 21040 -57086
rect 23002 -57088 23062 -57086
rect 20470 -57172 20484 -57130
rect 19500 -57706 19514 -57660
rect 18730 -57756 19218 -57750
rect 18730 -57790 18742 -57756
rect 19206 -57790 19218 -57756
rect 18730 -57796 19218 -57790
rect 19454 -57854 19514 -57706
rect 20478 -57706 20484 -57172
rect 20518 -57172 20530 -57130
rect 21496 -57130 21542 -57118
rect 20518 -57706 20524 -57172
rect 21496 -57660 21502 -57130
rect 20478 -57718 20524 -57706
rect 21490 -57706 21502 -57660
rect 21536 -57660 21542 -57130
rect 22514 -57130 22560 -57118
rect 21536 -57706 21550 -57660
rect 22514 -57668 22520 -57130
rect 19748 -57756 20236 -57750
rect 19748 -57790 19760 -57756
rect 20224 -57790 20236 -57756
rect 19748 -57796 20236 -57790
rect 20766 -57756 21254 -57750
rect 20766 -57790 20778 -57756
rect 21242 -57790 21254 -57756
rect 20766 -57796 21254 -57790
rect 21490 -57854 21550 -57706
rect 22508 -57706 22520 -57668
rect 22554 -57668 22560 -57130
rect 23532 -57130 23578 -57118
rect 22554 -57706 22568 -57668
rect 23532 -57674 23538 -57130
rect 21784 -57756 22272 -57750
rect 21784 -57790 21796 -57756
rect 22260 -57790 22272 -57756
rect 21784 -57796 22272 -57790
rect 19448 -57914 19454 -57854
rect 19514 -57914 19520 -57854
rect 21484 -57914 21490 -57854
rect 21550 -57914 21556 -57854
rect 18428 -58026 18434 -57966
rect 18494 -58026 18500 -57966
rect 19454 -58408 19514 -57914
rect 21490 -58408 21550 -57914
rect 22508 -57966 22568 -57706
rect 23526 -57706 23538 -57674
rect 23572 -57674 23578 -57130
rect 24546 -57130 24606 -56954
rect 25026 -57040 25086 -56954
rect 24838 -57046 25326 -57040
rect 24838 -57080 24850 -57046
rect 25314 -57080 25326 -57046
rect 24838 -57086 25326 -57080
rect 24546 -57198 24556 -57130
rect 23572 -57706 23586 -57674
rect 22802 -57756 23290 -57750
rect 22802 -57790 22814 -57756
rect 23278 -57790 23290 -57756
rect 22802 -57796 23290 -57790
rect 23526 -57854 23586 -57706
rect 24550 -57706 24556 -57198
rect 24590 -57198 24606 -57130
rect 25556 -57130 25616 -56954
rect 25556 -57170 25574 -57130
rect 24590 -57706 24596 -57198
rect 24550 -57718 24596 -57706
rect 25568 -57706 25574 -57170
rect 25608 -57170 25616 -57130
rect 25608 -57706 25614 -57170
rect 25568 -57718 25614 -57706
rect 23820 -57756 24308 -57750
rect 23820 -57790 23832 -57756
rect 24296 -57790 24308 -57756
rect 23820 -57796 24308 -57790
rect 24838 -57756 25326 -57750
rect 24838 -57790 24850 -57756
rect 25314 -57790 25326 -57756
rect 24838 -57796 25326 -57790
rect 23520 -57914 23526 -57854
rect 23586 -57914 23592 -57854
rect 22502 -58026 22508 -57966
rect 22568 -58026 22574 -57966
rect 23526 -58408 23586 -57914
rect 26514 -57966 26574 -51038
rect 26726 -51872 26786 -43532
rect 26720 -51932 26726 -51872
rect 26786 -51932 26792 -51872
rect 26846 -52000 26906 -43530
rect 26986 -45104 27046 -43512
rect 27098 -43650 27104 -43590
rect 27164 -43650 27170 -43590
rect 26980 -45164 26986 -45104
rect 27046 -45164 27052 -45104
rect 26986 -46860 27046 -45164
rect 26980 -46920 26986 -46860
rect 27046 -46920 27052 -46860
rect 26986 -48374 27046 -46920
rect 26980 -48434 26986 -48374
rect 27046 -48434 27052 -48374
rect 26986 -49616 27046 -48434
rect 26976 -49676 26982 -49616
rect 27042 -49676 27048 -49616
rect 26986 -50852 27046 -49676
rect 27104 -49718 27164 -43650
rect 27214 -44332 27274 -43496
rect 27208 -44392 27214 -44332
rect 27274 -44392 27280 -44332
rect 27332 -47252 27392 -43396
rect 27660 -44198 27720 -43386
rect 27654 -44258 27660 -44198
rect 27720 -44258 27726 -44198
rect 27780 -45104 27840 -43394
rect 27886 -43470 27946 -43464
rect 27774 -45164 27780 -45104
rect 27840 -45164 27846 -45104
rect 27450 -45616 27456 -45556
rect 27516 -45616 27522 -45556
rect 27330 -47258 27392 -47252
rect 27390 -47318 27392 -47258
rect 27330 -47324 27392 -47318
rect 27098 -49778 27104 -49718
rect 27164 -49778 27170 -49718
rect 26980 -50912 26986 -50852
rect 27046 -50912 27052 -50852
rect 26840 -52060 26846 -52000
rect 26906 -52060 26912 -52000
rect 26986 -52962 27046 -50912
rect 26980 -53022 26986 -52962
rect 27046 -53022 27052 -52962
rect 27332 -53320 27392 -47324
rect 27456 -48252 27516 -45616
rect 27662 -45952 27668 -45892
rect 27728 -45952 27734 -45892
rect 27558 -47212 27564 -47152
rect 27624 -47212 27630 -47152
rect 27450 -48312 27456 -48252
rect 27516 -48312 27522 -48252
rect 27564 -53170 27624 -47212
rect 27668 -48488 27728 -45952
rect 27780 -46860 27840 -45164
rect 27886 -46014 27946 -43530
rect 38692 -43826 38698 -43820
rect 28012 -43880 38698 -43826
rect 38758 -43826 38764 -43820
rect 43796 -43826 43802 -43820
rect 38758 -43880 43802 -43826
rect 43862 -43826 43868 -43820
rect 47862 -43826 47922 -43820
rect 43862 -43880 47862 -43826
rect 28012 -43886 47862 -43880
rect 47922 -43886 48434 -43826
rect 28012 -44026 28072 -43886
rect 28534 -43936 28594 -43886
rect 29544 -43936 29604 -43886
rect 28308 -43942 28796 -43936
rect 28308 -43976 28320 -43942
rect 28784 -43976 28796 -43942
rect 28308 -43982 28796 -43976
rect 29326 -43942 29814 -43936
rect 29326 -43976 29338 -43942
rect 29802 -43976 29814 -43942
rect 29326 -43982 29814 -43976
rect 29544 -43988 29604 -43982
rect 28012 -44602 28026 -44026
rect 28060 -44602 28072 -44026
rect 29038 -44026 29084 -44014
rect 29038 -44568 29044 -44026
rect 28012 -44844 28072 -44602
rect 29030 -44602 29044 -44568
rect 29078 -44568 29084 -44026
rect 30050 -44026 30110 -43886
rect 30574 -43936 30634 -43886
rect 31586 -43936 31646 -43886
rect 30344 -43942 30832 -43936
rect 30344 -43976 30356 -43942
rect 30820 -43976 30832 -43942
rect 30344 -43982 30832 -43976
rect 31362 -43942 31850 -43936
rect 31362 -43976 31374 -43942
rect 31838 -43976 31850 -43942
rect 31362 -43982 31850 -43976
rect 31586 -43988 31646 -43982
rect 29078 -44602 29090 -44568
rect 28308 -44652 28796 -44646
rect 28308 -44686 28320 -44652
rect 28784 -44686 28796 -44652
rect 28308 -44692 28796 -44686
rect 28524 -44754 28584 -44692
rect 28308 -44760 28796 -44754
rect 28308 -44794 28320 -44760
rect 28784 -44794 28796 -44760
rect 28308 -44800 28796 -44794
rect 28524 -44806 28584 -44800
rect 28012 -45420 28026 -44844
rect 28060 -45420 28072 -44844
rect 28012 -45892 28072 -45420
rect 29030 -44844 29090 -44602
rect 30050 -44602 30062 -44026
rect 30096 -44602 30110 -44026
rect 31074 -44026 31120 -44014
rect 31074 -44556 31080 -44026
rect 29530 -44646 29590 -44644
rect 29326 -44652 29814 -44646
rect 29326 -44686 29338 -44652
rect 29802 -44686 29814 -44652
rect 29326 -44692 29814 -44686
rect 29530 -44754 29590 -44692
rect 29326 -44760 29814 -44754
rect 29326 -44794 29338 -44760
rect 29802 -44794 29814 -44760
rect 29326 -44800 29814 -44794
rect 29030 -45420 29044 -44844
rect 29078 -45420 29090 -44844
rect 30050 -44844 30110 -44602
rect 31064 -44602 31080 -44556
rect 31114 -44556 31120 -44026
rect 32082 -44026 32142 -43886
rect 32598 -43936 32658 -43886
rect 33598 -43936 33658 -43886
rect 32380 -43942 32868 -43936
rect 32380 -43976 32392 -43942
rect 32856 -43976 32868 -43942
rect 32380 -43982 32868 -43976
rect 33398 -43942 33886 -43936
rect 33398 -43976 33410 -43942
rect 33874 -43976 33886 -43942
rect 33398 -43982 33886 -43976
rect 31114 -44602 31124 -44556
rect 30542 -44646 30602 -44638
rect 30344 -44652 30832 -44646
rect 30344 -44686 30356 -44652
rect 30820 -44686 30832 -44652
rect 30344 -44692 30832 -44686
rect 30542 -44754 30602 -44692
rect 30344 -44760 30832 -44754
rect 30344 -44794 30356 -44760
rect 30820 -44794 30832 -44760
rect 30344 -44800 30832 -44794
rect 30050 -44902 30062 -44844
rect 28308 -45470 28796 -45464
rect 28308 -45504 28320 -45470
rect 28784 -45504 28796 -45470
rect 28308 -45510 28796 -45504
rect 29030 -45556 29090 -45420
rect 30056 -45420 30062 -44902
rect 30096 -44902 30110 -44844
rect 31064 -44844 31124 -44602
rect 32082 -44602 32098 -44026
rect 32132 -44602 32142 -44026
rect 33110 -44026 33156 -44014
rect 33110 -44562 33116 -44026
rect 31362 -44652 31850 -44646
rect 31362 -44686 31374 -44652
rect 31838 -44686 31850 -44652
rect 31362 -44692 31850 -44686
rect 31564 -44754 31624 -44692
rect 31362 -44760 31850 -44754
rect 31362 -44794 31374 -44760
rect 31838 -44794 31850 -44760
rect 31362 -44800 31850 -44794
rect 31564 -44806 31624 -44800
rect 30096 -45420 30102 -44902
rect 30056 -45432 30102 -45420
rect 31064 -45420 31080 -44844
rect 31114 -45420 31124 -44844
rect 32082 -44844 32142 -44602
rect 33100 -44602 33116 -44562
rect 33150 -44562 33156 -44026
rect 34120 -44026 34180 -43886
rect 34632 -43936 34692 -43886
rect 35644 -43936 35704 -43886
rect 34416 -43942 34904 -43936
rect 34416 -43976 34428 -43942
rect 34892 -43976 34904 -43942
rect 34416 -43982 34904 -43976
rect 35434 -43942 35922 -43936
rect 35434 -43976 35446 -43942
rect 35910 -43976 35922 -43942
rect 35434 -43982 35922 -43976
rect 33150 -44602 33160 -44562
rect 32380 -44652 32868 -44646
rect 32380 -44686 32392 -44652
rect 32856 -44686 32868 -44652
rect 32380 -44692 32868 -44686
rect 32576 -44754 32636 -44692
rect 32380 -44760 32868 -44754
rect 32380 -44794 32392 -44760
rect 32856 -44794 32868 -44760
rect 32380 -44800 32868 -44794
rect 32576 -44806 32636 -44800
rect 32082 -44906 32098 -44844
rect 29326 -45470 29814 -45464
rect 29326 -45504 29338 -45470
rect 29802 -45504 29814 -45470
rect 29326 -45510 29814 -45504
rect 30344 -45470 30832 -45464
rect 30344 -45504 30356 -45470
rect 30820 -45504 30832 -45470
rect 30344 -45510 30832 -45504
rect 31064 -45558 31124 -45420
rect 32092 -45420 32098 -44906
rect 32132 -44906 32142 -44844
rect 33100 -44844 33160 -44602
rect 34120 -44602 34134 -44026
rect 34168 -44602 34180 -44026
rect 35146 -44026 35192 -44014
rect 35146 -44562 35152 -44026
rect 33398 -44652 33886 -44646
rect 33398 -44686 33410 -44652
rect 33874 -44686 33886 -44652
rect 33398 -44692 33886 -44686
rect 33606 -44754 33666 -44692
rect 33398 -44760 33886 -44754
rect 33398 -44794 33410 -44760
rect 33874 -44794 33886 -44760
rect 33398 -44800 33886 -44794
rect 33606 -44806 33666 -44800
rect 32132 -45420 32138 -44906
rect 32092 -45432 32138 -45420
rect 33100 -45420 33116 -44844
rect 33150 -45420 33160 -44844
rect 34120 -44844 34180 -44602
rect 35138 -44602 35152 -44562
rect 35186 -44562 35192 -44026
rect 36156 -44026 36216 -43886
rect 36668 -43936 36728 -43886
rect 37680 -43936 37740 -43886
rect 36452 -43942 36940 -43936
rect 36452 -43976 36464 -43942
rect 36928 -43976 36940 -43942
rect 36452 -43982 36940 -43976
rect 37470 -43942 37958 -43936
rect 37470 -43976 37482 -43942
rect 37946 -43976 37958 -43942
rect 37470 -43982 37958 -43976
rect 35186 -44602 35198 -44562
rect 34612 -44646 34672 -44644
rect 34416 -44652 34904 -44646
rect 34416 -44686 34428 -44652
rect 34892 -44686 34904 -44652
rect 34416 -44692 34904 -44686
rect 34612 -44754 34672 -44692
rect 34416 -44760 34904 -44754
rect 34416 -44794 34428 -44760
rect 34892 -44794 34904 -44760
rect 34416 -44800 34904 -44794
rect 34120 -44886 34134 -44844
rect 31362 -45470 31850 -45464
rect 31362 -45504 31374 -45470
rect 31838 -45504 31850 -45470
rect 31362 -45510 31850 -45504
rect 32380 -45470 32868 -45464
rect 32380 -45504 32392 -45470
rect 32856 -45504 32868 -45470
rect 32380 -45510 32868 -45504
rect 33100 -45558 33160 -45420
rect 34128 -45420 34134 -44886
rect 34168 -44886 34180 -44844
rect 35138 -44844 35198 -44602
rect 36156 -44602 36170 -44026
rect 36204 -44602 36216 -44026
rect 37182 -44026 37228 -44014
rect 37182 -44556 37188 -44026
rect 35634 -44646 35694 -44644
rect 35434 -44652 35922 -44646
rect 35434 -44686 35446 -44652
rect 35910 -44686 35922 -44652
rect 35434 -44692 35922 -44686
rect 35634 -44754 35694 -44692
rect 35434 -44760 35922 -44754
rect 35434 -44794 35446 -44760
rect 35910 -44794 35922 -44760
rect 35434 -44800 35922 -44794
rect 34168 -45420 34174 -44886
rect 34128 -45432 34174 -45420
rect 35138 -45420 35152 -44844
rect 35186 -45420 35198 -44844
rect 36156 -44844 36216 -44602
rect 37176 -44602 37188 -44556
rect 37222 -44556 37228 -44026
rect 38188 -44026 38248 -43886
rect 38702 -43936 38762 -43886
rect 39714 -43936 39774 -43886
rect 38488 -43942 38976 -43936
rect 38488 -43976 38500 -43942
rect 38964 -43976 38976 -43942
rect 38488 -43982 38976 -43976
rect 39506 -43942 39994 -43936
rect 39506 -43976 39518 -43942
rect 39982 -43976 39994 -43942
rect 39506 -43982 39994 -43976
rect 39714 -43988 39774 -43982
rect 37222 -44602 37236 -44556
rect 36452 -44652 36940 -44646
rect 36452 -44686 36464 -44652
rect 36928 -44686 36940 -44652
rect 36452 -44692 36940 -44686
rect 36658 -44754 36718 -44692
rect 36452 -44760 36940 -44754
rect 36452 -44794 36464 -44760
rect 36928 -44794 36940 -44760
rect 36452 -44800 36940 -44794
rect 36658 -44806 36718 -44800
rect 36156 -44894 36170 -44844
rect 33398 -45470 33886 -45464
rect 33398 -45504 33410 -45470
rect 33874 -45504 33886 -45470
rect 33398 -45510 33886 -45504
rect 34416 -45470 34904 -45464
rect 34416 -45504 34428 -45470
rect 34892 -45504 34904 -45470
rect 34416 -45510 34904 -45504
rect 35138 -45558 35198 -45420
rect 36164 -45420 36170 -44894
rect 36204 -44894 36216 -44844
rect 37176 -44844 37236 -44602
rect 38188 -44602 38206 -44026
rect 38240 -44602 38248 -44026
rect 39218 -44026 39264 -44014
rect 39218 -44556 39224 -44026
rect 37664 -44646 37724 -44644
rect 37470 -44652 37958 -44646
rect 37470 -44686 37482 -44652
rect 37946 -44686 37958 -44652
rect 37470 -44692 37958 -44686
rect 37664 -44754 37724 -44692
rect 37470 -44760 37958 -44754
rect 37470 -44794 37482 -44760
rect 37946 -44794 37958 -44760
rect 37470 -44800 37958 -44794
rect 36204 -45420 36210 -44894
rect 36164 -45432 36210 -45420
rect 37176 -45420 37188 -44844
rect 37222 -45420 37236 -44844
rect 38188 -44844 38248 -44602
rect 39210 -44602 39224 -44556
rect 39258 -44556 39264 -44026
rect 40226 -44026 40286 -43886
rect 40738 -43936 40798 -43886
rect 41756 -43936 41816 -43886
rect 40524 -43942 41012 -43936
rect 40524 -43976 40536 -43942
rect 41000 -43976 41012 -43942
rect 40524 -43982 41012 -43976
rect 41542 -43942 42030 -43936
rect 41542 -43976 41554 -43942
rect 42018 -43976 42030 -43942
rect 41542 -43982 42030 -43976
rect 40738 -43988 40798 -43982
rect 39258 -44602 39270 -44556
rect 38688 -44646 38748 -44638
rect 38488 -44652 38976 -44646
rect 38488 -44686 38500 -44652
rect 38964 -44686 38976 -44652
rect 38488 -44692 38976 -44686
rect 38688 -44754 38748 -44692
rect 38488 -44760 38976 -44754
rect 38488 -44794 38500 -44760
rect 38964 -44794 38976 -44760
rect 38488 -44800 38976 -44794
rect 38188 -44892 38206 -44844
rect 35434 -45470 35922 -45464
rect 35434 -45504 35446 -45470
rect 35910 -45504 35922 -45470
rect 35434 -45510 35922 -45504
rect 36452 -45470 36940 -45464
rect 36452 -45504 36464 -45470
rect 36928 -45504 36940 -45470
rect 36452 -45510 36940 -45504
rect 37176 -45558 37236 -45420
rect 38200 -45420 38206 -44892
rect 38240 -44892 38248 -44844
rect 39210 -44844 39270 -44602
rect 40226 -44602 40242 -44026
rect 40276 -44602 40286 -44026
rect 41254 -44026 41300 -44014
rect 41254 -44556 41260 -44026
rect 39710 -44646 39770 -44644
rect 39506 -44652 39994 -44646
rect 39506 -44686 39518 -44652
rect 39982 -44686 39994 -44652
rect 39506 -44692 39994 -44686
rect 39710 -44754 39770 -44692
rect 39506 -44760 39994 -44754
rect 39506 -44794 39518 -44760
rect 39982 -44794 39994 -44760
rect 39506 -44800 39994 -44794
rect 38240 -45420 38246 -44892
rect 38200 -45432 38246 -45420
rect 39210 -45420 39224 -44844
rect 39258 -45420 39270 -44844
rect 40226 -44844 40286 -44602
rect 41246 -44602 41260 -44556
rect 41294 -44556 41300 -44026
rect 42262 -44026 42322 -43886
rect 42778 -43936 42838 -43886
rect 43802 -43936 43862 -43886
rect 42560 -43942 43048 -43936
rect 42560 -43976 42572 -43942
rect 43036 -43976 43048 -43942
rect 42560 -43982 43048 -43976
rect 43578 -43942 44066 -43936
rect 43578 -43976 43590 -43942
rect 44054 -43976 44066 -43942
rect 43578 -43982 44066 -43976
rect 41294 -44602 41306 -44556
rect 40722 -44646 40782 -44644
rect 40524 -44652 41012 -44646
rect 40524 -44686 40536 -44652
rect 41000 -44686 41012 -44652
rect 40524 -44692 41012 -44686
rect 40722 -44754 40782 -44692
rect 40524 -44760 41012 -44754
rect 40524 -44794 40536 -44760
rect 41000 -44794 41012 -44760
rect 40524 -44800 41012 -44794
rect 40226 -44894 40242 -44844
rect 37470 -45470 37958 -45464
rect 37470 -45504 37482 -45470
rect 37946 -45504 37958 -45470
rect 37470 -45510 37958 -45504
rect 38488 -45470 38976 -45464
rect 38488 -45504 38500 -45470
rect 38964 -45504 38976 -45470
rect 38488 -45510 38976 -45504
rect 39210 -45558 39270 -45420
rect 40236 -45420 40242 -44894
rect 40276 -44894 40286 -44844
rect 41246 -44844 41306 -44602
rect 42262 -44602 42278 -44026
rect 42312 -44602 42322 -44026
rect 43290 -44026 43336 -44014
rect 43290 -44532 43296 -44026
rect 41542 -44652 42030 -44646
rect 41542 -44686 41554 -44652
rect 42018 -44686 42030 -44652
rect 41542 -44692 42030 -44686
rect 41734 -44754 41794 -44692
rect 41542 -44760 42030 -44754
rect 41542 -44794 41554 -44760
rect 42018 -44794 42030 -44760
rect 41542 -44800 42030 -44794
rect 41734 -44806 41794 -44800
rect 40276 -45420 40282 -44894
rect 40236 -45432 40282 -45420
rect 41246 -45420 41260 -44844
rect 41294 -45420 41306 -44844
rect 42262 -44844 42322 -44602
rect 43284 -44602 43296 -44532
rect 43330 -44532 43336 -44026
rect 44298 -44026 44358 -43886
rect 44820 -43936 44880 -43886
rect 45832 -43936 45892 -43886
rect 44596 -43942 45084 -43936
rect 44596 -43976 44608 -43942
rect 45072 -43976 45084 -43942
rect 44596 -43982 45084 -43976
rect 45614 -43942 46102 -43936
rect 45614 -43976 45626 -43942
rect 46090 -43976 46102 -43942
rect 45614 -43982 46102 -43976
rect 43330 -44602 43344 -44532
rect 42758 -44646 42818 -44638
rect 42560 -44652 43048 -44646
rect 42560 -44686 42572 -44652
rect 43036 -44686 43048 -44652
rect 42560 -44692 43048 -44686
rect 42758 -44754 42818 -44692
rect 42560 -44760 43048 -44754
rect 42560 -44794 42572 -44760
rect 43036 -44794 43048 -44760
rect 42560 -44800 43048 -44794
rect 42262 -44868 42278 -44844
rect 39506 -45470 39994 -45464
rect 39506 -45504 39518 -45470
rect 39982 -45504 39994 -45470
rect 39506 -45510 39994 -45504
rect 40524 -45470 41012 -45464
rect 40524 -45504 40536 -45470
rect 41000 -45504 41012 -45470
rect 40524 -45510 41012 -45504
rect 41246 -45558 41306 -45420
rect 42272 -45420 42278 -44868
rect 42312 -44868 42322 -44844
rect 43284 -44844 43344 -44602
rect 44298 -44602 44314 -44026
rect 44348 -44602 44358 -44026
rect 45326 -44026 45372 -44014
rect 45326 -44492 45332 -44026
rect 43578 -44652 44066 -44646
rect 43578 -44686 43590 -44652
rect 44054 -44686 44066 -44652
rect 43578 -44692 44066 -44686
rect 43780 -44754 43840 -44692
rect 43578 -44760 44066 -44754
rect 43578 -44794 43590 -44760
rect 44054 -44794 44066 -44760
rect 43578 -44800 44066 -44794
rect 43780 -44812 43840 -44800
rect 42312 -45420 42318 -44868
rect 42272 -45432 42318 -45420
rect 43284 -45420 43296 -44844
rect 43330 -45420 43344 -44844
rect 44298 -44844 44358 -44602
rect 45318 -44602 45332 -44492
rect 45366 -44492 45372 -44026
rect 46336 -44026 46396 -43886
rect 46842 -43936 46902 -43886
rect 47860 -43892 47922 -43886
rect 47860 -43936 47920 -43892
rect 46632 -43942 47120 -43936
rect 46632 -43976 46644 -43942
rect 47108 -43976 47120 -43942
rect 46632 -43982 47120 -43976
rect 47650 -43942 48138 -43936
rect 47650 -43976 47662 -43942
rect 48126 -43976 48138 -43942
rect 47650 -43982 48138 -43976
rect 45366 -44602 45378 -44492
rect 44798 -44646 44858 -44644
rect 44596 -44652 45084 -44646
rect 44596 -44686 44608 -44652
rect 45072 -44686 45084 -44652
rect 44596 -44692 45084 -44686
rect 44798 -44754 44858 -44692
rect 44596 -44760 45084 -44754
rect 44596 -44794 44608 -44760
rect 45072 -44794 45084 -44760
rect 44596 -44800 45084 -44794
rect 44298 -44886 44314 -44844
rect 41542 -45470 42030 -45464
rect 41542 -45504 41554 -45470
rect 42018 -45504 42030 -45470
rect 41542 -45510 42030 -45504
rect 42560 -45470 43048 -45464
rect 42560 -45504 42572 -45470
rect 43036 -45504 43048 -45470
rect 42560 -45510 43048 -45504
rect 43284 -45558 43344 -45420
rect 44308 -45420 44314 -44886
rect 44348 -44886 44358 -44844
rect 45318 -44844 45378 -44602
rect 46336 -44602 46350 -44026
rect 46384 -44602 46396 -44026
rect 47362 -44026 47408 -44014
rect 47362 -44542 47368 -44026
rect 45828 -44646 45888 -44632
rect 45614 -44652 46102 -44646
rect 45614 -44686 45626 -44652
rect 46090 -44686 46102 -44652
rect 45614 -44692 46102 -44686
rect 45828 -44754 45888 -44692
rect 45614 -44760 46102 -44754
rect 45614 -44794 45626 -44760
rect 46090 -44794 46102 -44760
rect 45614 -44800 46102 -44794
rect 44348 -45420 44354 -44886
rect 44308 -45432 44354 -45420
rect 45318 -45420 45332 -44844
rect 45366 -45420 45378 -44844
rect 46336 -44844 46396 -44602
rect 47354 -44602 47368 -44542
rect 47402 -44542 47408 -44026
rect 48374 -44026 48434 -43886
rect 47402 -44602 47414 -44542
rect 46840 -44646 46900 -44632
rect 46632 -44652 47120 -44646
rect 46632 -44686 46644 -44652
rect 47108 -44686 47120 -44652
rect 46632 -44692 47120 -44686
rect 46840 -44754 46900 -44692
rect 46632 -44760 47120 -44754
rect 46632 -44794 46644 -44760
rect 47108 -44794 47120 -44760
rect 46632 -44800 47120 -44794
rect 46336 -44886 46350 -44844
rect 43578 -45470 44066 -45464
rect 43578 -45504 43590 -45470
rect 44054 -45504 44066 -45470
rect 43578 -45510 44066 -45504
rect 44596 -45470 45084 -45464
rect 44596 -45504 44608 -45470
rect 45072 -45504 45084 -45470
rect 44596 -45510 45084 -45504
rect 45318 -45558 45378 -45420
rect 46344 -45420 46350 -44886
rect 46384 -44886 46396 -44844
rect 47354 -44844 47414 -44602
rect 48374 -44602 48386 -44026
rect 48420 -44602 48434 -44026
rect 47650 -44652 48138 -44646
rect 47650 -44686 47662 -44652
rect 48126 -44686 48138 -44652
rect 47650 -44692 48138 -44686
rect 47840 -44754 47900 -44692
rect 48374 -44694 48434 -44602
rect 50260 -44048 50372 -43262
rect 55800 -43278 56370 -43252
rect 56470 -43250 56476 -42487
rect 57622 -42486 57734 -42452
rect 56608 -42502 56668 -42496
rect 56720 -42502 56792 -42490
rect 57310 -42502 57382 -42490
rect 56668 -42562 56726 -42502
rect 56786 -42562 57316 -42502
rect 57376 -42562 57382 -42502
rect 56608 -42568 56668 -42562
rect 56720 -42574 56792 -42562
rect 56556 -42628 56602 -42616
rect 56556 -42784 56562 -42628
rect 56548 -42804 56562 -42784
rect 56596 -42784 56602 -42628
rect 56674 -42628 56720 -42616
rect 56674 -42784 56680 -42628
rect 56596 -42804 56608 -42784
rect 56548 -42854 56608 -42804
rect 56666 -42804 56680 -42784
rect 56714 -42784 56720 -42628
rect 56792 -42628 56838 -42616
rect 56792 -42778 56798 -42628
rect 56714 -42804 56726 -42784
rect 56542 -42866 56614 -42854
rect 56542 -42926 56548 -42866
rect 56608 -42926 56614 -42866
rect 56542 -42938 56614 -42926
rect 56548 -43250 56608 -42938
rect 56666 -43068 56726 -42804
rect 56788 -42804 56798 -42778
rect 56832 -42778 56838 -42628
rect 56902 -42628 56962 -42562
rect 56902 -42650 56916 -42628
rect 56832 -42804 56848 -42778
rect 56660 -43128 56666 -43068
rect 56726 -43128 56732 -43068
rect 56788 -43250 56848 -42804
rect 56910 -42804 56916 -42650
rect 56950 -42650 56962 -42628
rect 57028 -42628 57074 -42616
rect 56950 -42804 56956 -42650
rect 57028 -42792 57034 -42628
rect 56910 -42816 56956 -42804
rect 57020 -42804 57034 -42792
rect 57068 -42792 57074 -42628
rect 57140 -42628 57200 -42562
rect 57310 -42574 57382 -42562
rect 57140 -42642 57152 -42628
rect 57068 -42804 57080 -42792
rect 56918 -42868 56978 -42862
rect 56912 -42928 56918 -42868
rect 56978 -42928 56984 -42868
rect 56918 -42934 56978 -42928
rect 57020 -43250 57080 -42804
rect 57146 -42804 57152 -42642
rect 57186 -42642 57200 -42628
rect 57264 -42628 57310 -42616
rect 57186 -42804 57192 -42642
rect 57264 -42780 57270 -42628
rect 57146 -42816 57192 -42804
rect 57256 -42804 57270 -42780
rect 57304 -42780 57310 -42628
rect 57382 -42628 57428 -42616
rect 57382 -42780 57388 -42628
rect 57304 -42804 57316 -42780
rect 57138 -42868 57198 -42862
rect 57132 -42928 57138 -42868
rect 57198 -42928 57204 -42868
rect 57138 -42934 57198 -42928
rect 57256 -43250 57316 -42804
rect 57374 -42804 57388 -42780
rect 57422 -42780 57428 -42628
rect 57500 -42628 57546 -42616
rect 57500 -42762 57506 -42628
rect 57422 -42804 57434 -42780
rect 57374 -43068 57434 -42804
rect 57496 -42804 57506 -42762
rect 57540 -42762 57546 -42628
rect 57540 -42804 57556 -42762
rect 57496 -42854 57556 -42804
rect 57490 -42866 57562 -42854
rect 57490 -42926 57496 -42866
rect 57556 -42926 57562 -42866
rect 57490 -42938 57562 -42926
rect 57368 -43128 57374 -43068
rect 57434 -43128 57440 -43068
rect 57496 -43250 57556 -42938
rect 57622 -43250 57628 -42486
rect 56470 -43278 57628 -43250
rect 57728 -43250 57734 -42486
rect 57794 -42624 57854 -42612
rect 57794 -42918 57806 -42624
rect 57840 -42918 57854 -42624
rect 57940 -42674 57946 -42574
rect 58046 -42674 58052 -42574
rect 58140 -42624 58200 -42614
rect 57914 -42714 57960 -42702
rect 57914 -42854 57920 -42714
rect 57794 -43250 57854 -42918
rect 57904 -42890 57920 -42854
rect 57954 -42854 57960 -42714
rect 58032 -42714 58078 -42702
rect 58032 -42848 58038 -42714
rect 57954 -42890 57964 -42854
rect 57904 -43068 57964 -42890
rect 58024 -42890 58038 -42848
rect 58072 -42848 58078 -42714
rect 58072 -42890 58084 -42848
rect 58024 -42968 58084 -42890
rect 58140 -42918 58152 -42624
rect 58186 -42918 58200 -42624
rect 58018 -43028 58024 -42968
rect 58084 -43028 58090 -42968
rect 57898 -43128 57904 -43068
rect 57964 -43128 57970 -43068
rect 58140 -43250 58200 -42918
rect 58256 -42968 58316 -41926
rect 58250 -43028 58256 -42968
rect 58316 -43028 58322 -42968
rect 57728 -43278 58288 -43250
rect 55800 -43584 55824 -43278
rect 58268 -43584 58288 -43278
rect 55800 -43602 58288 -43584
rect 56364 -43604 57734 -43602
rect 56364 -43704 56470 -43604
rect 57628 -43704 57734 -43604
rect 56364 -43710 57734 -43704
rect 48374 -44754 49154 -44694
rect 47650 -44760 48138 -44754
rect 47650 -44794 47662 -44760
rect 48126 -44794 48138 -44760
rect 47650 -44800 48138 -44794
rect 47840 -44806 47900 -44800
rect 46384 -45420 46390 -44886
rect 46344 -45432 46390 -45420
rect 47354 -45420 47368 -44844
rect 47402 -45420 47414 -44844
rect 48374 -44844 48434 -44754
rect 48374 -44894 48386 -44844
rect 45614 -45470 46102 -45464
rect 45614 -45504 45626 -45470
rect 46090 -45504 46102 -45470
rect 45614 -45510 46102 -45504
rect 46632 -45470 47120 -45464
rect 46632 -45504 46644 -45470
rect 47108 -45504 47120 -45470
rect 46632 -45510 47120 -45504
rect 47354 -45558 47414 -45420
rect 48380 -45420 48386 -44894
rect 48420 -44894 48434 -44844
rect 48420 -45420 48426 -44894
rect 48380 -45432 48426 -45420
rect 47650 -45470 48138 -45464
rect 47650 -45504 47662 -45470
rect 48126 -45504 48138 -45470
rect 47650 -45510 48138 -45504
rect 29090 -45616 49032 -45558
rect 29030 -45618 49032 -45616
rect 29030 -45622 29090 -45618
rect 30038 -45832 30044 -45772
rect 30104 -45832 30110 -45772
rect 32078 -45832 32084 -45772
rect 32144 -45832 32150 -45772
rect 34118 -45832 34124 -45772
rect 34184 -45832 34190 -45772
rect 36148 -45832 36154 -45772
rect 36214 -45832 36220 -45772
rect 38188 -45832 38194 -45772
rect 38254 -45832 38260 -45772
rect 40220 -45832 40226 -45772
rect 40286 -45832 40292 -45772
rect 42260 -45832 42266 -45772
rect 42326 -45832 42332 -45772
rect 44296 -45832 44302 -45772
rect 44362 -45832 44368 -45772
rect 46330 -45832 46336 -45772
rect 46396 -45832 46402 -45772
rect 28006 -45952 28012 -45892
rect 28072 -45952 28078 -45892
rect 29530 -45958 29536 -45898
rect 29596 -45958 29602 -45898
rect 27880 -46074 27886 -46014
rect 27946 -46074 27952 -46014
rect 27774 -46920 27780 -46860
rect 27840 -46920 27846 -46860
rect 27780 -48374 27840 -46920
rect 27886 -48148 27946 -46074
rect 29536 -46132 29596 -45958
rect 28308 -46138 28796 -46132
rect 28308 -46172 28320 -46138
rect 28784 -46172 28796 -46138
rect 28308 -46178 28796 -46172
rect 29326 -46138 29814 -46132
rect 29326 -46172 29338 -46138
rect 29802 -46172 29814 -46138
rect 29326 -46178 29814 -46172
rect 28020 -46222 28066 -46210
rect 29038 -46222 29084 -46210
rect 30044 -46222 30104 -45832
rect 30550 -45898 30610 -45892
rect 30550 -46132 30610 -45958
rect 31572 -45898 31632 -45892
rect 31572 -46132 31632 -45958
rect 30344 -46138 30832 -46132
rect 30344 -46172 30356 -46138
rect 30820 -46172 30832 -46138
rect 30344 -46178 30832 -46172
rect 31362 -46138 31850 -46132
rect 31362 -46172 31374 -46138
rect 31838 -46172 31850 -46138
rect 31362 -46178 31850 -46172
rect 31074 -46222 31120 -46210
rect 28012 -46256 28026 -46222
rect 28020 -46748 28026 -46256
rect 28012 -46798 28026 -46748
rect 28060 -46256 28072 -46222
rect 28060 -46748 28066 -46256
rect 29030 -46270 29044 -46222
rect 28060 -46798 28072 -46748
rect 29038 -46762 29044 -46270
rect 28012 -46936 28072 -46798
rect 29030 -46798 29044 -46762
rect 29078 -46270 29090 -46222
rect 29078 -46762 29084 -46270
rect 30044 -46290 30062 -46222
rect 30056 -46734 30062 -46290
rect 29078 -46798 29090 -46762
rect 28308 -46848 28796 -46842
rect 28308 -46882 28320 -46848
rect 28784 -46882 28796 -46848
rect 28308 -46888 28796 -46882
rect 28514 -46936 28574 -46888
rect 29030 -46936 29090 -46798
rect 30048 -46798 30062 -46734
rect 30096 -46254 30108 -46222
rect 30096 -46290 30104 -46254
rect 30096 -46734 30102 -46290
rect 30096 -46798 30108 -46734
rect 31074 -46752 31080 -46222
rect 31070 -46770 31080 -46752
rect 31068 -46798 31080 -46770
rect 31114 -46752 31120 -46222
rect 32084 -46222 32144 -45832
rect 32586 -45898 32646 -45892
rect 32584 -45958 32586 -45952
rect 33612 -45898 33672 -45892
rect 32584 -45964 32646 -45958
rect 33610 -45958 33612 -45952
rect 33610 -45964 33672 -45958
rect 32584 -46132 32644 -45964
rect 33094 -46074 33100 -46014
rect 33160 -46074 33166 -46014
rect 32380 -46138 32868 -46132
rect 32380 -46172 32392 -46138
rect 32856 -46172 32868 -46138
rect 32380 -46178 32868 -46172
rect 32084 -46276 32098 -46222
rect 32092 -46726 32098 -46276
rect 32088 -46750 32098 -46726
rect 31114 -46798 31130 -46752
rect 32086 -46798 32098 -46750
rect 32132 -46276 32144 -46222
rect 33100 -46222 33160 -46074
rect 33610 -46132 33670 -45964
rect 33398 -46138 33886 -46132
rect 33398 -46172 33410 -46138
rect 33874 -46172 33886 -46138
rect 33398 -46178 33886 -46172
rect 33100 -46264 33116 -46222
rect 32132 -46726 32138 -46276
rect 33110 -46722 33116 -46264
rect 32132 -46798 32148 -46726
rect 33100 -46798 33116 -46722
rect 33150 -46264 33160 -46222
rect 34124 -46222 34184 -45832
rect 34624 -45898 34684 -45892
rect 34624 -46132 34684 -45958
rect 35660 -45898 35720 -45892
rect 35660 -46132 35720 -45958
rect 34416 -46138 34904 -46132
rect 34416 -46172 34428 -46138
rect 34892 -46172 34904 -46138
rect 34416 -46178 34904 -46172
rect 35434 -46138 35922 -46132
rect 35434 -46172 35446 -46138
rect 35910 -46172 35922 -46138
rect 35434 -46178 35922 -46172
rect 35146 -46222 35192 -46210
rect 36154 -46222 36214 -45832
rect 36666 -45898 36726 -45892
rect 37674 -45958 37680 -45898
rect 37740 -45958 37746 -45898
rect 36666 -46132 36726 -45958
rect 37680 -46132 37740 -45958
rect 36452 -46138 36940 -46132
rect 36452 -46172 36464 -46138
rect 36928 -46172 36940 -46138
rect 36452 -46178 36940 -46172
rect 37470 -46138 37958 -46132
rect 37470 -46172 37482 -46138
rect 37946 -46172 37958 -46138
rect 37470 -46178 37958 -46172
rect 33150 -46722 33156 -46264
rect 34124 -46296 34134 -46222
rect 33150 -46738 33160 -46722
rect 33150 -46798 33164 -46738
rect 34128 -46742 34134 -46296
rect 34120 -46798 34134 -46742
rect 34168 -46296 34184 -46222
rect 35140 -46272 35152 -46222
rect 34168 -46742 34174 -46296
rect 35146 -46734 35152 -46272
rect 34168 -46798 34180 -46742
rect 35140 -46762 35152 -46734
rect 35138 -46798 35152 -46762
rect 35186 -46272 35200 -46222
rect 35186 -46734 35192 -46272
rect 36154 -46290 36170 -46222
rect 36164 -46722 36170 -46290
rect 35186 -46798 35200 -46734
rect 29326 -46848 29814 -46842
rect 29326 -46882 29338 -46848
rect 29802 -46882 29814 -46848
rect 29326 -46888 29814 -46882
rect 28012 -46996 29090 -46936
rect 29030 -47152 29090 -46996
rect 29540 -47046 29600 -46888
rect 30048 -46936 30108 -46798
rect 30344 -46848 30832 -46842
rect 30344 -46882 30356 -46848
rect 30820 -46882 30832 -46848
rect 30344 -46888 30832 -46882
rect 30042 -46996 30048 -46936
rect 30108 -46996 30114 -46936
rect 29534 -47106 29540 -47046
rect 29600 -47106 29606 -47046
rect 29024 -47212 29030 -47152
rect 29090 -47212 29096 -47152
rect 28010 -47318 28016 -47258
rect 28076 -47318 28082 -47258
rect 28508 -47318 28514 -47258
rect 28574 -47318 28580 -47258
rect 29020 -47318 29026 -47258
rect 29086 -47318 29092 -47258
rect 28016 -47454 28076 -47318
rect 28514 -47364 28574 -47318
rect 28308 -47370 28796 -47364
rect 28308 -47404 28320 -47370
rect 28784 -47404 28796 -47370
rect 28308 -47410 28796 -47404
rect 28016 -47494 28026 -47454
rect 28020 -48030 28026 -47494
rect 28060 -47494 28076 -47454
rect 29026 -47454 29086 -47318
rect 29540 -47364 29600 -47106
rect 29326 -47370 29814 -47364
rect 29326 -47404 29338 -47370
rect 29802 -47404 29814 -47370
rect 29326 -47410 29814 -47404
rect 28060 -48030 28066 -47494
rect 29026 -47500 29044 -47454
rect 28020 -48042 28066 -48030
rect 29038 -48030 29044 -47500
rect 29078 -47500 29086 -47454
rect 30048 -47454 30108 -46996
rect 30562 -47046 30622 -46888
rect 30556 -47106 30562 -47046
rect 30622 -47106 30628 -47046
rect 30562 -47364 30622 -47106
rect 31070 -47152 31130 -46798
rect 31362 -46848 31850 -46842
rect 31362 -46882 31374 -46848
rect 31838 -46882 31850 -46848
rect 31362 -46888 31850 -46882
rect 31576 -47046 31636 -46888
rect 32088 -46936 32148 -46798
rect 33110 -46810 33156 -46798
rect 32380 -46848 32868 -46842
rect 32380 -46882 32392 -46848
rect 32856 -46882 32868 -46848
rect 32380 -46888 32868 -46882
rect 33398 -46848 33886 -46842
rect 33398 -46882 33410 -46848
rect 33874 -46882 33886 -46848
rect 33398 -46888 33886 -46882
rect 32082 -46996 32088 -46936
rect 32148 -46996 32154 -46936
rect 31570 -47106 31576 -47046
rect 31636 -47106 31642 -47046
rect 31064 -47212 31070 -47152
rect 31130 -47212 31136 -47152
rect 31576 -47364 31636 -47106
rect 30344 -47370 30832 -47364
rect 30344 -47404 30356 -47370
rect 30820 -47404 30832 -47370
rect 30344 -47410 30832 -47404
rect 31362 -47370 31850 -47364
rect 31362 -47404 31374 -47370
rect 31838 -47404 31850 -47370
rect 31362 -47410 31850 -47404
rect 31074 -47454 31120 -47442
rect 32088 -47454 32148 -46996
rect 32590 -47046 32650 -46888
rect 33608 -47046 33668 -46888
rect 34120 -46936 34180 -46798
rect 34416 -46848 34904 -46842
rect 34416 -46882 34428 -46848
rect 34892 -46882 34904 -46848
rect 34416 -46888 34904 -46882
rect 34114 -46996 34120 -46936
rect 34180 -46996 34186 -46936
rect 32584 -47106 32590 -47046
rect 32650 -47106 32656 -47046
rect 33602 -47106 33608 -47046
rect 33668 -47106 33674 -47046
rect 32590 -47364 32650 -47106
rect 33094 -47212 33100 -47152
rect 33160 -47212 33166 -47152
rect 32380 -47370 32868 -47364
rect 32380 -47404 32392 -47370
rect 32856 -47404 32868 -47370
rect 32380 -47410 32868 -47404
rect 30048 -47492 30062 -47454
rect 29078 -48030 29084 -47500
rect 30056 -47972 30062 -47492
rect 29038 -48042 29084 -48030
rect 30042 -48030 30062 -47972
rect 30096 -47492 30108 -47454
rect 30096 -48030 30102 -47492
rect 31068 -47506 31080 -47454
rect 31074 -48010 31080 -47506
rect 28308 -48080 28796 -48074
rect 28308 -48114 28320 -48080
rect 28784 -48114 28796 -48080
rect 28308 -48120 28796 -48114
rect 29326 -48080 29814 -48074
rect 29326 -48114 29338 -48080
rect 29802 -48114 29814 -48080
rect 29326 -48120 29814 -48114
rect 27880 -48208 27886 -48148
rect 27946 -48208 27952 -48148
rect 30042 -48252 30102 -48030
rect 31064 -48030 31080 -48010
rect 31114 -47506 31128 -47454
rect 31114 -48010 31120 -47506
rect 32086 -47518 32098 -47454
rect 32092 -47966 32098 -47518
rect 31114 -48030 31124 -48010
rect 30344 -48080 30832 -48074
rect 30344 -48114 30356 -48080
rect 30820 -48114 30832 -48080
rect 30344 -48120 30832 -48114
rect 28004 -48312 28010 -48252
rect 28070 -48312 28076 -48252
rect 29524 -48312 29530 -48252
rect 29590 -48312 29596 -48252
rect 30036 -48312 30042 -48252
rect 30102 -48312 30108 -48252
rect 27774 -48434 27780 -48374
rect 27840 -48434 27846 -48374
rect 27662 -48548 27668 -48488
rect 27728 -48548 27734 -48488
rect 27780 -49616 27840 -48434
rect 28010 -48688 28070 -48312
rect 28510 -48548 28516 -48488
rect 28576 -48548 28582 -48488
rect 28516 -48598 28576 -48548
rect 29530 -48598 29590 -48312
rect 30042 -48546 30048 -48486
rect 30108 -48546 30114 -48486
rect 28306 -48604 28794 -48598
rect 28306 -48638 28318 -48604
rect 28782 -48638 28794 -48604
rect 28306 -48644 28794 -48638
rect 29324 -48604 29812 -48598
rect 29324 -48638 29336 -48604
rect 29800 -48638 29812 -48604
rect 29324 -48644 29812 -48638
rect 29036 -48688 29082 -48676
rect 30048 -48688 30108 -48546
rect 30546 -48598 30606 -48120
rect 31064 -48148 31124 -48030
rect 32078 -48030 32098 -47966
rect 32132 -47488 32148 -47454
rect 33100 -47454 33160 -47212
rect 33608 -47364 33668 -47106
rect 33398 -47370 33886 -47364
rect 33398 -47404 33410 -47370
rect 33874 -47404 33886 -47370
rect 33398 -47410 33886 -47404
rect 34120 -47454 34180 -46996
rect 34634 -47046 34694 -46888
rect 35140 -47006 35200 -46798
rect 36152 -46798 36170 -46722
rect 36204 -46290 36214 -46222
rect 37182 -46222 37228 -46210
rect 36204 -46722 36210 -46290
rect 36204 -46798 36212 -46722
rect 37182 -46736 37188 -46222
rect 37176 -46738 37188 -46736
rect 35434 -46848 35922 -46842
rect 35434 -46882 35446 -46848
rect 35910 -46882 35922 -46848
rect 35434 -46888 35922 -46882
rect 34628 -47106 34634 -47046
rect 34694 -47106 34700 -47046
rect 35140 -47066 35366 -47006
rect 35654 -47046 35714 -46888
rect 36152 -46936 36212 -46798
rect 37174 -46798 37188 -46738
rect 37222 -46736 37228 -46222
rect 38194 -46222 38254 -45832
rect 38696 -45898 38756 -45892
rect 38696 -46132 38756 -45958
rect 39704 -45898 39764 -45892
rect 39764 -45958 39766 -45952
rect 39704 -45964 39766 -45958
rect 39706 -46132 39766 -45964
rect 38488 -46138 38976 -46132
rect 38488 -46172 38500 -46138
rect 38964 -46172 38976 -46138
rect 38488 -46178 38976 -46172
rect 39506 -46138 39994 -46132
rect 39506 -46172 39518 -46138
rect 39982 -46172 39994 -46138
rect 39506 -46178 39994 -46172
rect 39218 -46222 39264 -46210
rect 40226 -46222 40286 -45832
rect 40720 -45898 40780 -45892
rect 41744 -45898 41804 -45892
rect 40780 -45958 40782 -45952
rect 40720 -45964 40782 -45958
rect 40722 -46132 40782 -45964
rect 41744 -46132 41804 -45958
rect 40524 -46138 41012 -46132
rect 40524 -46172 40536 -46138
rect 41000 -46172 41012 -46138
rect 40524 -46178 41012 -46172
rect 41542 -46138 42030 -46132
rect 41542 -46172 41554 -46138
rect 42018 -46172 42030 -46138
rect 41542 -46178 42030 -46172
rect 41254 -46222 41300 -46210
rect 42266 -46222 42326 -45832
rect 42766 -45898 42826 -45892
rect 43788 -45898 43848 -45892
rect 42766 -46132 42826 -45958
rect 43786 -45958 43788 -45952
rect 43786 -45964 43848 -45958
rect 43282 -46074 43288 -46014
rect 43348 -46074 43354 -46014
rect 42560 -46138 43048 -46132
rect 42560 -46172 42572 -46138
rect 43036 -46172 43048 -46138
rect 42560 -46178 43048 -46172
rect 38194 -46290 38206 -46222
rect 38200 -46732 38206 -46290
rect 37222 -46798 37236 -46736
rect 38188 -46798 38206 -46732
rect 38240 -46290 38254 -46222
rect 39208 -46256 39224 -46222
rect 38240 -46732 38246 -46290
rect 38240 -46798 38248 -46732
rect 39218 -46750 39224 -46256
rect 36452 -46848 36940 -46842
rect 36452 -46882 36464 -46848
rect 36928 -46882 36940 -46848
rect 36452 -46888 36940 -46882
rect 36146 -46996 36152 -46936
rect 36212 -46996 36218 -46936
rect 34634 -47364 34694 -47106
rect 35134 -47212 35140 -47152
rect 35200 -47212 35206 -47152
rect 34416 -47370 34904 -47364
rect 34416 -47404 34428 -47370
rect 34892 -47404 34904 -47370
rect 34416 -47410 34904 -47404
rect 35140 -47454 35200 -47212
rect 35306 -47258 35366 -47066
rect 35648 -47106 35654 -47046
rect 35714 -47106 35720 -47046
rect 35300 -47318 35306 -47258
rect 35366 -47318 35372 -47258
rect 35654 -47364 35714 -47106
rect 35434 -47370 35922 -47364
rect 35434 -47404 35446 -47370
rect 35910 -47404 35922 -47370
rect 35434 -47410 35922 -47404
rect 32132 -47518 32146 -47488
rect 33100 -47498 33116 -47454
rect 32132 -48030 32138 -47518
rect 31362 -48080 31850 -48074
rect 31362 -48114 31374 -48080
rect 31838 -48114 31850 -48080
rect 31362 -48120 31850 -48114
rect 31058 -48208 31064 -48148
rect 31124 -48208 31130 -48148
rect 31060 -48312 31066 -48252
rect 31126 -48312 31132 -48252
rect 30342 -48604 30830 -48598
rect 30342 -48638 30354 -48604
rect 30818 -48638 30830 -48604
rect 30342 -48644 30830 -48638
rect 28010 -48744 28024 -48688
rect 28018 -49264 28024 -48744
rect 28058 -48744 28070 -48688
rect 29030 -48720 29042 -48688
rect 28058 -49264 28064 -48744
rect 29036 -49220 29042 -48720
rect 28018 -49276 28064 -49264
rect 29030 -49264 29042 -49220
rect 29076 -48720 29090 -48688
rect 30048 -48714 30060 -48688
rect 29076 -49220 29082 -48720
rect 29076 -49264 29090 -49220
rect 28306 -49314 28794 -49308
rect 28306 -49348 28318 -49314
rect 28782 -49348 28794 -49314
rect 28306 -49354 28794 -49348
rect 29030 -49416 29090 -49264
rect 30054 -49264 30060 -48714
rect 30094 -48714 30108 -48688
rect 31066 -48688 31126 -48312
rect 31566 -48598 31626 -48120
rect 32078 -48252 32138 -48030
rect 33110 -48030 33116 -47498
rect 33150 -47488 33162 -47454
rect 33150 -47498 33160 -47488
rect 34120 -47496 34134 -47454
rect 33150 -48030 33156 -47498
rect 34128 -47988 34134 -47496
rect 34120 -48030 34134 -47988
rect 34168 -47496 34180 -47454
rect 34168 -47988 34174 -47496
rect 35136 -47516 35152 -47454
rect 34168 -48030 34180 -47988
rect 35146 -48030 35152 -47516
rect 35186 -47494 35200 -47454
rect 36152 -47454 36212 -46996
rect 36674 -47046 36734 -46888
rect 36668 -47106 36674 -47046
rect 36734 -47106 36740 -47046
rect 36674 -47364 36734 -47106
rect 37174 -47152 37234 -46798
rect 37470 -46848 37958 -46842
rect 37470 -46882 37482 -46848
rect 37946 -46882 37958 -46848
rect 37470 -46888 37958 -46882
rect 37676 -47046 37736 -46888
rect 38188 -46936 38248 -46798
rect 39210 -46798 39224 -46750
rect 39258 -46256 39268 -46222
rect 39258 -46750 39264 -46256
rect 40226 -46276 40242 -46222
rect 40236 -46738 40242 -46276
rect 39258 -46798 39270 -46750
rect 38488 -46848 38976 -46842
rect 38488 -46882 38500 -46848
rect 38964 -46882 38976 -46848
rect 38488 -46888 38976 -46882
rect 38182 -46996 38188 -46936
rect 38248 -46996 38254 -46936
rect 37670 -47106 37676 -47046
rect 37736 -47106 37742 -47046
rect 37168 -47212 37174 -47152
rect 37234 -47212 37240 -47152
rect 37168 -47318 37174 -47258
rect 37234 -47318 37240 -47258
rect 36452 -47370 36940 -47364
rect 36452 -47404 36464 -47370
rect 36928 -47404 36940 -47370
rect 36452 -47410 36940 -47404
rect 37174 -47454 37234 -47318
rect 37676 -47364 37736 -47106
rect 37470 -47370 37958 -47364
rect 37470 -47404 37482 -47370
rect 37946 -47404 37958 -47370
rect 37470 -47410 37958 -47404
rect 38188 -47454 38248 -46996
rect 38702 -47046 38762 -46888
rect 38696 -47106 38702 -47046
rect 38762 -47106 38768 -47046
rect 38702 -47364 38762 -47106
rect 39210 -47152 39270 -46798
rect 40224 -46798 40242 -46738
rect 40276 -46276 40286 -46222
rect 41246 -46262 41260 -46222
rect 40276 -46738 40282 -46276
rect 41254 -46732 41260 -46262
rect 40276 -46798 40284 -46738
rect 41250 -46758 41260 -46732
rect 39506 -46848 39994 -46842
rect 39506 -46882 39518 -46848
rect 39982 -46882 39994 -46848
rect 39506 -46888 39994 -46882
rect 39720 -47046 39780 -46888
rect 40224 -46936 40284 -46798
rect 41248 -46798 41260 -46758
rect 41294 -46262 41306 -46222
rect 41294 -46732 41300 -46262
rect 42266 -46276 42278 -46222
rect 41294 -46798 41310 -46732
rect 42272 -46748 42278 -46276
rect 42262 -46798 42278 -46748
rect 42312 -46276 42326 -46222
rect 43288 -46222 43348 -46074
rect 43786 -46132 43846 -45964
rect 43578 -46138 44066 -46132
rect 43578 -46172 43590 -46138
rect 44054 -46172 44066 -46138
rect 43578 -46178 44066 -46172
rect 42312 -46748 42318 -46276
rect 43288 -46286 43296 -46222
rect 43290 -46742 43296 -46286
rect 42312 -46798 42322 -46748
rect 43282 -46798 43296 -46742
rect 43330 -46286 43348 -46222
rect 44302 -46222 44362 -45832
rect 44806 -45898 44866 -45892
rect 45820 -45898 45880 -45892
rect 44866 -45958 44868 -45952
rect 44806 -45964 44868 -45958
rect 45880 -45958 45882 -45952
rect 45820 -45964 45882 -45958
rect 44808 -46132 44868 -45964
rect 45822 -46132 45882 -45964
rect 44596 -46138 45084 -46132
rect 44596 -46172 44608 -46138
rect 45072 -46172 45084 -46138
rect 44596 -46178 45084 -46172
rect 45614 -46138 46102 -46132
rect 45614 -46172 45626 -46138
rect 46090 -46172 46102 -46138
rect 45614 -46178 46102 -46172
rect 45326 -46222 45372 -46210
rect 46336 -46222 46396 -45832
rect 46844 -45898 46904 -45892
rect 46842 -45958 46844 -45952
rect 46842 -45964 46904 -45958
rect 46842 -46132 46902 -45964
rect 47354 -46074 47360 -46014
rect 47420 -46074 47426 -46014
rect 48486 -46074 48492 -46014
rect 48552 -46074 48558 -46014
rect 46632 -46138 47120 -46132
rect 46632 -46172 46644 -46138
rect 47108 -46172 47120 -46138
rect 46632 -46178 47120 -46172
rect 47360 -46222 47420 -46074
rect 47650 -46138 48138 -46132
rect 47650 -46172 47662 -46138
rect 48126 -46172 48138 -46138
rect 47650 -46178 48138 -46172
rect 44302 -46282 44314 -46222
rect 43330 -46742 43336 -46286
rect 43330 -46744 43342 -46742
rect 43330 -46798 43344 -46744
rect 44308 -46762 44314 -46282
rect 44300 -46798 44314 -46762
rect 44348 -46282 44362 -46222
rect 45318 -46262 45332 -46222
rect 44348 -46762 44354 -46282
rect 45326 -46742 45332 -46262
rect 44348 -46798 44360 -46762
rect 40524 -46848 41012 -46842
rect 40524 -46882 40536 -46848
rect 41000 -46882 41012 -46848
rect 40524 -46888 41012 -46882
rect 40218 -46996 40224 -46936
rect 40284 -46996 40290 -46936
rect 39714 -47106 39720 -47046
rect 39780 -47106 39786 -47046
rect 39204 -47212 39210 -47152
rect 39270 -47212 39276 -47152
rect 39206 -47318 39212 -47258
rect 39272 -47318 39278 -47258
rect 38488 -47370 38976 -47364
rect 38488 -47404 38500 -47370
rect 38964 -47404 38976 -47370
rect 38488 -47410 38976 -47404
rect 39212 -47454 39272 -47318
rect 39720 -47364 39780 -47106
rect 39506 -47370 39994 -47364
rect 39506 -47404 39518 -47370
rect 39982 -47404 39994 -47370
rect 39506 -47410 39994 -47404
rect 40224 -47454 40284 -46996
rect 40728 -47046 40788 -46888
rect 41248 -47014 41308 -46798
rect 41740 -46842 41800 -46840
rect 41542 -46848 42030 -46842
rect 41542 -46882 41554 -46848
rect 42018 -46882 42030 -46848
rect 41542 -46888 42030 -46882
rect 40722 -47106 40728 -47046
rect 40788 -47106 40794 -47046
rect 41092 -47074 41308 -47014
rect 41740 -47046 41800 -46888
rect 42262 -46936 42322 -46798
rect 43290 -46810 43336 -46798
rect 42772 -46842 42832 -46840
rect 42560 -46848 43048 -46842
rect 42560 -46882 42572 -46848
rect 43036 -46882 43048 -46848
rect 42560 -46888 43048 -46882
rect 43578 -46848 44066 -46842
rect 43578 -46882 43590 -46848
rect 44054 -46882 44066 -46848
rect 43578 -46888 44066 -46882
rect 42256 -46996 42262 -46936
rect 42322 -46996 42328 -46936
rect 40728 -47364 40788 -47106
rect 41092 -47258 41152 -47074
rect 41734 -47106 41740 -47046
rect 41800 -47106 41806 -47046
rect 41240 -47212 41246 -47152
rect 41306 -47212 41312 -47152
rect 41086 -47318 41092 -47258
rect 41152 -47318 41158 -47258
rect 40524 -47370 41012 -47364
rect 40524 -47404 40536 -47370
rect 41000 -47404 41012 -47370
rect 40524 -47410 41012 -47404
rect 35186 -47516 35196 -47494
rect 36152 -47510 36170 -47454
rect 35186 -48030 35192 -47516
rect 36164 -47988 36170 -47510
rect 33110 -48042 33156 -48030
rect 34128 -48042 34174 -48030
rect 35146 -48042 35192 -48030
rect 36156 -48030 36170 -47988
rect 36204 -47510 36212 -47454
rect 37172 -47506 37188 -47454
rect 36204 -47988 36210 -47510
rect 36204 -48030 36216 -47988
rect 32380 -48080 32868 -48074
rect 32380 -48114 32392 -48080
rect 32856 -48114 32868 -48080
rect 32380 -48120 32868 -48114
rect 33398 -48080 33886 -48074
rect 33398 -48114 33410 -48080
rect 33874 -48114 33886 -48080
rect 33398 -48120 33886 -48114
rect 34416 -48080 34904 -48074
rect 34416 -48114 34428 -48080
rect 34892 -48114 34904 -48080
rect 34416 -48120 34904 -48114
rect 35434 -48080 35922 -48074
rect 35434 -48114 35446 -48080
rect 35910 -48114 35922 -48080
rect 35434 -48120 35922 -48114
rect 32072 -48312 32078 -48252
rect 32138 -48312 32144 -48252
rect 32078 -48546 32084 -48486
rect 32144 -48546 32150 -48486
rect 31360 -48604 31848 -48598
rect 31360 -48638 31372 -48604
rect 31836 -48638 31848 -48604
rect 31360 -48644 31848 -48638
rect 30094 -49264 30100 -48714
rect 31066 -48720 31078 -48688
rect 31072 -49224 31078 -48720
rect 30054 -49276 30100 -49264
rect 31064 -49264 31078 -49224
rect 31112 -48720 31126 -48688
rect 32084 -48688 32144 -48546
rect 32578 -48598 32638 -48120
rect 33092 -48312 33098 -48252
rect 33158 -48312 33164 -48252
rect 32378 -48604 32866 -48598
rect 32378 -48638 32390 -48604
rect 32854 -48638 32866 -48604
rect 32378 -48644 32866 -48638
rect 32084 -48718 32096 -48688
rect 31112 -49224 31118 -48720
rect 31112 -49264 31124 -49224
rect 29324 -49314 29812 -49308
rect 29324 -49348 29336 -49314
rect 29800 -49348 29812 -49314
rect 29324 -49354 29812 -49348
rect 30342 -49314 30830 -49308
rect 30342 -49348 30354 -49314
rect 30818 -49348 30830 -49314
rect 30342 -49354 30830 -49348
rect 27886 -49476 27892 -49416
rect 27952 -49476 27958 -49416
rect 29024 -49476 29030 -49416
rect 29090 -49476 29096 -49416
rect 27774 -49676 27780 -49616
rect 27840 -49676 27846 -49616
rect 27668 -49778 27674 -49718
rect 27734 -49778 27740 -49718
rect 27558 -53230 27564 -53170
rect 27624 -53230 27630 -53170
rect 27674 -53208 27734 -49778
rect 27780 -50852 27840 -49676
rect 27774 -50912 27780 -50852
rect 27840 -50912 27846 -50852
rect 27780 -52962 27840 -50912
rect 27892 -52190 27952 -49476
rect 29022 -49676 29028 -49616
rect 29088 -49676 29094 -49616
rect 29028 -49720 29088 -49676
rect 28012 -49780 29088 -49720
rect 28012 -49782 28576 -49780
rect 28012 -49922 28072 -49782
rect 28516 -49832 28576 -49782
rect 28306 -49838 28794 -49832
rect 28306 -49872 28318 -49838
rect 28782 -49872 28794 -49838
rect 28306 -49878 28794 -49872
rect 28012 -49954 28024 -49922
rect 28018 -50498 28024 -49954
rect 28058 -49954 28072 -49922
rect 29028 -49922 29088 -49780
rect 29532 -49832 29592 -49354
rect 30040 -49556 30046 -49496
rect 30106 -49556 30112 -49496
rect 29324 -49838 29812 -49832
rect 29324 -49872 29336 -49838
rect 29800 -49872 29812 -49838
rect 29324 -49878 29812 -49872
rect 28058 -50498 28064 -49954
rect 29028 -49958 29042 -49922
rect 28018 -50510 28064 -50498
rect 29036 -50498 29042 -49958
rect 29076 -49958 29088 -49922
rect 30046 -49922 30106 -49556
rect 30560 -49610 30620 -49354
rect 31064 -49392 31124 -49264
rect 32090 -49264 32096 -48718
rect 32130 -48718 32144 -48688
rect 33098 -48688 33158 -48312
rect 33604 -48598 33664 -48120
rect 34114 -48208 34120 -48148
rect 34180 -48208 34186 -48148
rect 33396 -48604 33884 -48598
rect 33396 -48638 33408 -48604
rect 33872 -48638 33884 -48604
rect 33396 -48644 33884 -48638
rect 32130 -49264 32136 -48718
rect 33098 -48732 33114 -48688
rect 33108 -49214 33114 -48732
rect 32090 -49276 32136 -49264
rect 33100 -49264 33114 -49214
rect 33148 -48732 33158 -48688
rect 34120 -48688 34180 -48208
rect 36156 -48252 36216 -48030
rect 37182 -48030 37188 -47506
rect 37222 -47498 37236 -47454
rect 37222 -47506 37232 -47498
rect 38188 -47502 38206 -47454
rect 37222 -48030 37228 -47506
rect 38200 -47982 38206 -47502
rect 37182 -48042 37228 -48030
rect 38194 -48030 38206 -47982
rect 38240 -47502 38248 -47454
rect 39208 -47494 39224 -47454
rect 38240 -47982 38246 -47502
rect 38240 -48030 38254 -47982
rect 36452 -48080 36940 -48074
rect 36452 -48114 36464 -48080
rect 36928 -48114 36940 -48080
rect 36452 -48120 36940 -48114
rect 37470 -48080 37958 -48074
rect 37470 -48114 37482 -48080
rect 37946 -48114 37958 -48080
rect 37470 -48120 37958 -48114
rect 38194 -48252 38254 -48030
rect 39218 -48030 39224 -47494
rect 39258 -47492 39274 -47454
rect 39258 -47494 39272 -47492
rect 39258 -48030 39264 -47494
rect 40224 -47500 40242 -47454
rect 40236 -47976 40242 -47500
rect 40224 -48030 40242 -47976
rect 40276 -47500 40284 -47454
rect 41246 -47454 41306 -47212
rect 41740 -47364 41800 -47106
rect 41542 -47370 42030 -47364
rect 41542 -47404 41554 -47370
rect 42018 -47404 42030 -47370
rect 41542 -47410 42030 -47404
rect 42262 -47454 42322 -46996
rect 42772 -47046 42832 -46888
rect 43786 -47046 43846 -46888
rect 44300 -46936 44360 -46798
rect 45316 -46798 45332 -46742
rect 45366 -46262 45378 -46222
rect 45366 -46742 45372 -46262
rect 45366 -46798 45376 -46742
rect 44596 -46848 45084 -46842
rect 44596 -46882 44608 -46848
rect 45072 -46882 45084 -46848
rect 44596 -46888 45084 -46882
rect 44294 -46996 44300 -46936
rect 44360 -46996 44366 -46936
rect 42766 -47106 42772 -47046
rect 42832 -47106 42838 -47046
rect 43780 -47106 43786 -47046
rect 43846 -47106 43852 -47046
rect 42772 -47364 42832 -47106
rect 43280 -47212 43286 -47152
rect 43346 -47212 43352 -47152
rect 42560 -47370 43048 -47364
rect 42560 -47404 42572 -47370
rect 43036 -47404 43048 -47370
rect 42560 -47410 43048 -47404
rect 43286 -47454 43346 -47212
rect 43786 -47364 43846 -47106
rect 43578 -47370 44066 -47364
rect 43578 -47404 43590 -47370
rect 44054 -47404 44066 -47370
rect 43578 -47410 44066 -47404
rect 40276 -47976 40282 -47500
rect 41246 -47506 41260 -47454
rect 40276 -48030 40284 -47976
rect 41254 -48030 41260 -47506
rect 41294 -47496 41310 -47454
rect 41294 -47506 41306 -47496
rect 41294 -48030 41300 -47506
rect 39218 -48042 39264 -48030
rect 40236 -48042 40282 -48030
rect 41254 -48042 41300 -48030
rect 42262 -48030 42278 -47454
rect 42312 -48030 42322 -47454
rect 43282 -47496 43296 -47454
rect 43286 -47516 43296 -47496
rect 38488 -48080 38976 -48074
rect 38488 -48114 38500 -48080
rect 38964 -48114 38976 -48080
rect 38488 -48120 38976 -48114
rect 39506 -48080 39994 -48074
rect 39506 -48114 39518 -48080
rect 39982 -48114 39994 -48080
rect 39506 -48120 39994 -48114
rect 40524 -48080 41012 -48074
rect 40524 -48114 40536 -48080
rect 41000 -48114 41012 -48080
rect 40524 -48120 41012 -48114
rect 41542 -48080 42030 -48074
rect 41542 -48114 41554 -48080
rect 42018 -48114 42030 -48080
rect 41542 -48120 42030 -48114
rect 40220 -48208 40226 -48148
rect 40286 -48208 40292 -48148
rect 36150 -48312 36156 -48252
rect 36216 -48312 36222 -48252
rect 38188 -48312 38194 -48252
rect 38254 -48312 38260 -48252
rect 35134 -48434 35140 -48374
rect 35200 -48434 35206 -48374
rect 37168 -48434 37174 -48374
rect 37234 -48434 37240 -48374
rect 39198 -48434 39204 -48374
rect 39264 -48434 39270 -48374
rect 34414 -48604 34902 -48598
rect 34414 -48638 34426 -48604
rect 34890 -48638 34902 -48604
rect 34414 -48644 34902 -48638
rect 33148 -49214 33154 -48732
rect 34120 -48750 34132 -48688
rect 33148 -49264 33160 -49214
rect 34126 -49228 34132 -48750
rect 31360 -49314 31848 -49308
rect 31360 -49348 31372 -49314
rect 31836 -49348 31848 -49314
rect 31360 -49354 31848 -49348
rect 32378 -49314 32866 -49308
rect 32378 -49348 32390 -49314
rect 32854 -49348 32866 -49314
rect 32378 -49354 32866 -49348
rect 31058 -49452 31064 -49392
rect 31124 -49452 31130 -49392
rect 30554 -49670 30560 -49610
rect 30620 -49670 30626 -49610
rect 30560 -49832 30620 -49670
rect 30342 -49838 30830 -49832
rect 30342 -49872 30354 -49838
rect 30818 -49872 30830 -49838
rect 30342 -49878 30830 -49872
rect 29076 -50498 29082 -49958
rect 30046 -49964 30060 -49922
rect 30054 -50440 30060 -49964
rect 29036 -50510 29082 -50498
rect 30048 -50498 30060 -50440
rect 30094 -49964 30106 -49922
rect 31064 -49922 31124 -49452
rect 31562 -49604 31622 -49354
rect 32080 -49556 32086 -49496
rect 32146 -49556 32152 -49496
rect 31562 -49610 31624 -49604
rect 31562 -49670 31564 -49610
rect 31562 -49676 31624 -49670
rect 31562 -49832 31622 -49676
rect 31360 -49838 31848 -49832
rect 31360 -49872 31372 -49838
rect 31836 -49872 31848 -49838
rect 31360 -49878 31848 -49872
rect 30094 -50440 30100 -49964
rect 31064 -49966 31078 -49922
rect 30094 -50498 30108 -50440
rect 31072 -50450 31078 -49966
rect 28306 -50548 28794 -50542
rect 28306 -50582 28318 -50548
rect 28782 -50582 28794 -50548
rect 28306 -50588 28794 -50582
rect 29324 -50548 29812 -50542
rect 29324 -50582 29336 -50548
rect 29800 -50582 29812 -50548
rect 29324 -50588 29812 -50582
rect 29022 -50708 29028 -50648
rect 29088 -50708 29094 -50648
rect 28306 -51070 28794 -51064
rect 28306 -51104 28318 -51070
rect 28782 -51104 28794 -51070
rect 28306 -51110 28794 -51104
rect 28018 -51154 28064 -51142
rect 28018 -51684 28024 -51154
rect 28008 -51730 28024 -51684
rect 28058 -51684 28064 -51154
rect 29028 -51154 29088 -50708
rect 29534 -50750 29594 -50588
rect 29528 -50810 29534 -50750
rect 29594 -50810 29600 -50750
rect 30048 -50952 30108 -50498
rect 31066 -50498 31078 -50450
rect 31112 -49966 31124 -49922
rect 32086 -49922 32146 -49556
rect 32578 -49604 32638 -49354
rect 33100 -49392 33160 -49264
rect 34118 -49264 34132 -49228
rect 34166 -48750 34180 -48688
rect 35140 -48688 35200 -48434
rect 35432 -48604 35920 -48598
rect 35432 -48638 35444 -48604
rect 35908 -48638 35920 -48604
rect 35432 -48644 35920 -48638
rect 36450 -48604 36938 -48598
rect 36450 -48638 36462 -48604
rect 36926 -48638 36938 -48604
rect 36450 -48644 36938 -48638
rect 35140 -48744 35150 -48688
rect 34166 -49228 34172 -48750
rect 34166 -49264 34178 -49228
rect 33396 -49314 33884 -49308
rect 33396 -49348 33408 -49314
rect 33872 -49348 33884 -49314
rect 33396 -49354 33884 -49348
rect 33094 -49452 33100 -49392
rect 33160 -49452 33166 -49392
rect 32576 -49610 32638 -49604
rect 32636 -49670 32638 -49610
rect 32576 -49676 32638 -49670
rect 32578 -49832 32638 -49676
rect 32378 -49838 32866 -49832
rect 32378 -49872 32390 -49838
rect 32854 -49872 32866 -49838
rect 32378 -49878 32866 -49872
rect 32086 -49964 32096 -49922
rect 31112 -50450 31118 -49966
rect 31112 -50498 31126 -50450
rect 30342 -50548 30830 -50542
rect 30342 -50582 30354 -50548
rect 30818 -50582 30830 -50548
rect 30342 -50588 30830 -50582
rect 31066 -50648 31126 -50498
rect 32090 -50498 32096 -49964
rect 32130 -49964 32146 -49922
rect 33100 -49922 33160 -49452
rect 33596 -49610 33656 -49354
rect 34118 -49496 34178 -49264
rect 35144 -49264 35150 -48744
rect 35184 -48744 35200 -48688
rect 36162 -48688 36208 -48676
rect 35184 -49264 35190 -48744
rect 36162 -49234 36168 -48688
rect 35144 -49276 35190 -49264
rect 36152 -49264 36168 -49234
rect 36202 -49234 36208 -48688
rect 37174 -48688 37234 -48434
rect 37468 -48604 37956 -48598
rect 37468 -48638 37480 -48604
rect 37944 -48638 37956 -48604
rect 37468 -48644 37956 -48638
rect 38486 -48604 38974 -48598
rect 38486 -48638 38498 -48604
rect 38962 -48638 38974 -48604
rect 38486 -48644 38974 -48638
rect 37174 -48738 37186 -48688
rect 36202 -49264 36212 -49234
rect 34414 -49314 34902 -49308
rect 34414 -49348 34426 -49314
rect 34890 -49348 34902 -49314
rect 34414 -49354 34902 -49348
rect 35432 -49314 35920 -49308
rect 35432 -49348 35444 -49314
rect 35908 -49348 35920 -49314
rect 35432 -49354 35920 -49348
rect 34112 -49556 34118 -49496
rect 34178 -49556 34184 -49496
rect 34608 -49552 34668 -49354
rect 35650 -49552 35710 -49354
rect 36152 -49496 36212 -49264
rect 37180 -49264 37186 -48738
rect 37220 -48738 37234 -48688
rect 38198 -48688 38244 -48676
rect 37220 -49264 37226 -48738
rect 38198 -49222 38204 -48688
rect 37180 -49276 37226 -49264
rect 38192 -49264 38204 -49222
rect 38238 -49222 38244 -48688
rect 39204 -48688 39264 -48434
rect 39504 -48604 39992 -48598
rect 39504 -48638 39516 -48604
rect 39980 -48638 39992 -48604
rect 39504 -48644 39992 -48638
rect 39204 -48732 39222 -48688
rect 38238 -49264 38252 -49222
rect 36450 -49314 36938 -49308
rect 36450 -49348 36462 -49314
rect 36926 -49348 36938 -49314
rect 36450 -49354 36938 -49348
rect 37468 -49314 37956 -49308
rect 37468 -49348 37480 -49314
rect 37944 -49348 37956 -49314
rect 37468 -49354 37956 -49348
rect 34112 -49668 34118 -49608
rect 34178 -49668 34184 -49608
rect 34608 -49612 35710 -49552
rect 36146 -49556 36152 -49496
rect 36212 -49556 36218 -49496
rect 33596 -49832 33656 -49670
rect 33396 -49838 33884 -49832
rect 33396 -49872 33408 -49838
rect 33872 -49872 33884 -49838
rect 33396 -49878 33884 -49872
rect 32130 -50498 32136 -49964
rect 33100 -49970 33114 -49922
rect 33108 -50448 33114 -49970
rect 32090 -50510 32136 -50498
rect 33102 -50498 33114 -50448
rect 33148 -49970 33160 -49922
rect 34118 -49922 34178 -49668
rect 34608 -49832 34668 -49612
rect 35130 -49778 35136 -49718
rect 35196 -49778 35202 -49718
rect 34414 -49838 34902 -49832
rect 34414 -49872 34426 -49838
rect 34890 -49872 34902 -49838
rect 34414 -49878 34902 -49872
rect 33148 -50448 33154 -49970
rect 34118 -49980 34132 -49922
rect 33148 -50498 33162 -50448
rect 31360 -50548 31848 -50542
rect 31360 -50582 31372 -50548
rect 31836 -50582 31848 -50548
rect 31360 -50588 31848 -50582
rect 32378 -50548 32866 -50542
rect 32378 -50582 32390 -50548
rect 32854 -50582 32866 -50548
rect 32378 -50588 32866 -50582
rect 31060 -50708 31066 -50648
rect 31126 -50708 31132 -50648
rect 31058 -50912 31064 -50852
rect 31124 -50912 31130 -50852
rect 31572 -50858 31632 -50588
rect 32594 -50858 32654 -50588
rect 33102 -50648 33162 -50498
rect 34126 -50498 34132 -49980
rect 34166 -49980 34178 -49922
rect 35136 -49922 35196 -49778
rect 35650 -49832 35710 -49612
rect 36148 -49668 36154 -49608
rect 36214 -49668 36220 -49608
rect 35432 -49838 35920 -49832
rect 35432 -49872 35444 -49838
rect 35908 -49872 35920 -49838
rect 35432 -49878 35920 -49872
rect 35136 -49968 35150 -49922
rect 34166 -50498 34172 -49980
rect 34126 -50510 34172 -50498
rect 35144 -50498 35150 -49968
rect 35184 -49968 35196 -49922
rect 36154 -49922 36214 -49668
rect 36650 -49832 36710 -49354
rect 37164 -49778 37170 -49718
rect 37230 -49778 37236 -49718
rect 36450 -49838 36938 -49832
rect 36450 -49872 36462 -49838
rect 36926 -49872 36938 -49838
rect 36450 -49878 36938 -49872
rect 35184 -50498 35190 -49968
rect 36154 -49990 36168 -49922
rect 35144 -50510 35190 -50498
rect 36162 -50498 36168 -49990
rect 36202 -49990 36214 -49922
rect 37170 -49922 37230 -49778
rect 37684 -49832 37744 -49354
rect 38192 -49496 38252 -49264
rect 39216 -49264 39222 -48732
rect 39256 -48732 39264 -48688
rect 40226 -48688 40286 -48208
rect 40748 -48598 40808 -48120
rect 41238 -48312 41244 -48252
rect 41304 -48312 41310 -48252
rect 40522 -48604 41010 -48598
rect 40522 -48638 40534 -48604
rect 40998 -48638 41010 -48604
rect 40522 -48644 41010 -48638
rect 39256 -49264 39262 -48732
rect 40226 -48740 40240 -48688
rect 40234 -49212 40240 -48740
rect 39216 -49276 39262 -49264
rect 40226 -49264 40240 -49212
rect 40274 -48740 40286 -48688
rect 41244 -48688 41304 -48312
rect 41750 -48598 41810 -48120
rect 42262 -48252 42322 -48030
rect 43290 -48030 43296 -47516
rect 43330 -47516 43346 -47454
rect 44300 -47454 44360 -46996
rect 44804 -47046 44864 -46888
rect 44798 -47106 44804 -47046
rect 44864 -47106 44870 -47046
rect 44804 -47364 44864 -47106
rect 45316 -47152 45376 -46798
rect 46336 -46798 46350 -46222
rect 46384 -46254 46398 -46222
rect 47356 -46250 47368 -46222
rect 46384 -46798 46396 -46254
rect 47360 -46286 47368 -46250
rect 47362 -46738 47368 -46286
rect 45614 -46848 46102 -46842
rect 45614 -46882 45626 -46848
rect 46090 -46882 46102 -46848
rect 45614 -46888 46102 -46882
rect 45828 -47046 45888 -46888
rect 46336 -46936 46396 -46798
rect 47356 -46798 47368 -46738
rect 47402 -46286 47420 -46222
rect 48380 -46222 48426 -46210
rect 47402 -46738 47408 -46286
rect 47402 -46798 47416 -46738
rect 48380 -46750 48386 -46222
rect 46632 -46848 47120 -46842
rect 46632 -46882 46644 -46848
rect 47108 -46882 47120 -46848
rect 46632 -46888 47120 -46882
rect 46330 -46996 46336 -46936
rect 46396 -46996 46402 -46936
rect 45822 -47106 45828 -47046
rect 45888 -47106 45894 -47046
rect 45310 -47212 45316 -47152
rect 45376 -47212 45382 -47152
rect 45310 -47316 45316 -47256
rect 45376 -47316 45382 -47256
rect 44596 -47370 45084 -47364
rect 44596 -47404 44608 -47370
rect 45072 -47404 45084 -47370
rect 44596 -47410 45084 -47404
rect 44796 -47422 44856 -47410
rect 45316 -47454 45376 -47316
rect 45828 -47364 45888 -47106
rect 45614 -47370 46102 -47364
rect 45614 -47404 45626 -47370
rect 46090 -47404 46102 -47370
rect 45614 -47410 46102 -47404
rect 44300 -47512 44314 -47454
rect 43330 -48030 43336 -47516
rect 44308 -47982 44314 -47512
rect 43290 -48042 43336 -48030
rect 44298 -48030 44314 -47982
rect 44348 -47512 44360 -47454
rect 45314 -47500 45332 -47454
rect 44348 -47982 44354 -47512
rect 45316 -47528 45332 -47500
rect 45326 -47976 45332 -47528
rect 44348 -48030 44358 -47982
rect 42560 -48080 43048 -48074
rect 42560 -48114 42572 -48080
rect 43036 -48114 43048 -48080
rect 42560 -48120 43048 -48114
rect 43578 -48080 44066 -48074
rect 43578 -48114 43590 -48080
rect 44054 -48114 44066 -48080
rect 43578 -48120 44066 -48114
rect 42256 -48312 42262 -48252
rect 42322 -48312 42328 -48252
rect 42762 -48598 42822 -48120
rect 43276 -48312 43282 -48252
rect 43342 -48312 43348 -48252
rect 41540 -48604 42028 -48598
rect 41540 -48638 41552 -48604
rect 42016 -48638 42028 -48604
rect 41540 -48644 42028 -48638
rect 42558 -48604 43046 -48598
rect 42558 -48638 42570 -48604
rect 43034 -48638 43046 -48604
rect 42558 -48644 43046 -48638
rect 41244 -48736 41258 -48688
rect 40274 -49212 40280 -48740
rect 40274 -49264 40286 -49212
rect 41252 -49232 41258 -48736
rect 38486 -49314 38974 -49308
rect 38486 -49348 38498 -49314
rect 38962 -49348 38974 -49314
rect 38486 -49354 38974 -49348
rect 39504 -49314 39992 -49308
rect 39504 -49348 39516 -49314
rect 39980 -49348 39992 -49314
rect 39504 -49354 39992 -49348
rect 38186 -49556 38192 -49496
rect 38252 -49556 38258 -49496
rect 38706 -49552 38766 -49354
rect 39714 -49552 39774 -49354
rect 40226 -49496 40286 -49264
rect 41244 -49264 41258 -49232
rect 41292 -48736 41304 -48688
rect 42270 -48688 42316 -48676
rect 41292 -49232 41298 -48736
rect 42270 -49228 42276 -48688
rect 41292 -49264 41304 -49232
rect 40522 -49314 41010 -49308
rect 40522 -49348 40534 -49314
rect 40998 -49348 41010 -49314
rect 40522 -49354 41010 -49348
rect 38184 -49668 38190 -49608
rect 38250 -49668 38256 -49608
rect 38706 -49612 39774 -49552
rect 40220 -49556 40226 -49496
rect 40286 -49556 40292 -49496
rect 40416 -49560 40422 -49500
rect 40482 -49560 40488 -49500
rect 37468 -49838 37956 -49832
rect 37468 -49872 37480 -49838
rect 37944 -49872 37956 -49838
rect 37468 -49878 37956 -49872
rect 37170 -49970 37186 -49922
rect 36202 -50498 36208 -49990
rect 36162 -50510 36208 -50498
rect 37180 -50498 37186 -49970
rect 37220 -49970 37230 -49922
rect 38190 -49922 38250 -49668
rect 38706 -49832 38766 -49612
rect 39204 -49778 39210 -49718
rect 39270 -49778 39276 -49718
rect 38486 -49838 38974 -49832
rect 38486 -49872 38498 -49838
rect 38962 -49872 38974 -49838
rect 38486 -49878 38974 -49872
rect 37220 -50498 37226 -49970
rect 38190 -49972 38204 -49922
rect 37180 -50510 37226 -50498
rect 38198 -50498 38204 -49972
rect 38238 -49972 38250 -49922
rect 39210 -49922 39270 -49778
rect 39714 -49832 39774 -49612
rect 40220 -49668 40226 -49608
rect 40286 -49668 40292 -49608
rect 39504 -49838 39992 -49832
rect 39504 -49872 39516 -49838
rect 39980 -49872 39992 -49838
rect 39504 -49878 39992 -49872
rect 39210 -49960 39222 -49922
rect 38238 -50498 38244 -49972
rect 39216 -50452 39222 -49960
rect 38198 -50510 38244 -50498
rect 39210 -50498 39222 -50452
rect 39256 -49960 39270 -49922
rect 40226 -49922 40286 -49668
rect 40422 -49718 40482 -49560
rect 40716 -49716 40776 -49354
rect 41244 -49392 41304 -49264
rect 42260 -49264 42276 -49228
rect 42310 -49228 42316 -48688
rect 43282 -48688 43342 -48312
rect 43796 -48598 43856 -48120
rect 44298 -48252 44358 -48030
rect 45320 -48030 45332 -47976
rect 45366 -47528 45376 -47454
rect 46336 -47454 46396 -46996
rect 46848 -47046 46908 -46888
rect 47356 -46946 47416 -46798
rect 48372 -46798 48386 -46750
rect 48420 -46750 48426 -46222
rect 48420 -46798 48432 -46750
rect 47650 -46848 48138 -46842
rect 47650 -46882 47662 -46848
rect 48126 -46882 48138 -46848
rect 47650 -46888 48138 -46882
rect 47866 -46946 47926 -46888
rect 48372 -46946 48432 -46798
rect 48492 -46946 48552 -46074
rect 47356 -47006 48552 -46946
rect 46842 -47106 46848 -47046
rect 46908 -47106 46914 -47046
rect 46848 -47364 46908 -47106
rect 47350 -47212 47356 -47152
rect 47416 -47212 47422 -47152
rect 47356 -47254 47416 -47212
rect 47356 -47314 48434 -47254
rect 48492 -47256 48552 -47006
rect 46632 -47370 47120 -47364
rect 46632 -47404 46644 -47370
rect 47108 -47404 47120 -47370
rect 46632 -47410 47120 -47404
rect 46336 -47480 46350 -47454
rect 45366 -47976 45372 -47528
rect 46344 -47972 46350 -47480
rect 45366 -48030 45380 -47976
rect 44596 -48080 45084 -48074
rect 44596 -48114 44608 -48080
rect 45072 -48114 45084 -48080
rect 44596 -48120 45084 -48114
rect 45320 -48148 45380 -48030
rect 46334 -48030 46350 -47972
rect 46384 -47480 46396 -47454
rect 47356 -47454 47416 -47314
rect 47842 -47364 47902 -47314
rect 47650 -47370 48138 -47364
rect 47650 -47404 47662 -47370
rect 48126 -47404 48138 -47370
rect 47650 -47410 48138 -47404
rect 48374 -47454 48434 -47314
rect 48486 -47316 48492 -47256
rect 48552 -47316 48558 -47256
rect 46384 -47972 46390 -47480
rect 47356 -47510 47368 -47454
rect 46384 -48030 46394 -47972
rect 45614 -48080 46102 -48074
rect 45614 -48114 45626 -48080
rect 46090 -48114 46102 -48080
rect 45614 -48120 46102 -48114
rect 45314 -48208 45320 -48148
rect 45380 -48208 45386 -48148
rect 46334 -48252 46394 -48030
rect 47362 -48030 47368 -47510
rect 47402 -47510 47416 -47454
rect 48370 -47490 48386 -47454
rect 48374 -47496 48386 -47490
rect 47402 -48030 47408 -47510
rect 48380 -47986 48386 -47496
rect 47362 -48042 47408 -48030
rect 48376 -48030 48386 -47986
rect 48420 -47496 48434 -47454
rect 48420 -47986 48426 -47496
rect 48420 -48030 48436 -47986
rect 46632 -48080 47120 -48074
rect 46632 -48114 46644 -48080
rect 47108 -48114 47120 -48080
rect 46632 -48120 47120 -48114
rect 47650 -48080 48138 -48074
rect 47650 -48114 47662 -48080
rect 48126 -48114 48138 -48080
rect 47650 -48120 48138 -48114
rect 44292 -48312 44298 -48252
rect 44358 -48312 44364 -48252
rect 46328 -48312 46334 -48252
rect 46394 -48312 46400 -48252
rect 46824 -48598 46884 -48120
rect 48376 -48156 48436 -48030
rect 48376 -48216 48666 -48156
rect 47862 -48522 48430 -48462
rect 47862 -48598 47922 -48522
rect 43576 -48604 44064 -48598
rect 43576 -48638 43588 -48604
rect 44052 -48638 44064 -48604
rect 43576 -48644 44064 -48638
rect 44594 -48604 45082 -48598
rect 44594 -48638 44606 -48604
rect 45070 -48638 45082 -48604
rect 44594 -48644 45082 -48638
rect 45612 -48604 46100 -48598
rect 45612 -48638 45624 -48604
rect 46088 -48638 46100 -48604
rect 45612 -48644 46100 -48638
rect 46630 -48604 47118 -48598
rect 46630 -48638 46642 -48604
rect 47106 -48638 47118 -48604
rect 46630 -48644 47118 -48638
rect 47648 -48604 48136 -48598
rect 47648 -48638 47660 -48604
rect 48124 -48638 48136 -48604
rect 47648 -48644 48136 -48638
rect 43282 -48746 43294 -48688
rect 43288 -49218 43294 -48746
rect 42310 -49264 42320 -49228
rect 41540 -49314 42028 -49308
rect 41540 -49348 41552 -49314
rect 42016 -49348 42028 -49314
rect 41540 -49354 42028 -49348
rect 41238 -49452 41244 -49392
rect 41304 -49452 41310 -49392
rect 40416 -49778 40422 -49718
rect 40482 -49778 40488 -49718
rect 40710 -49776 40716 -49716
rect 40776 -49776 40782 -49716
rect 40716 -49832 40776 -49776
rect 40522 -49838 41010 -49832
rect 40522 -49872 40534 -49838
rect 40998 -49872 41010 -49838
rect 40522 -49878 41010 -49872
rect 39256 -50452 39262 -49960
rect 40226 -49966 40240 -49922
rect 39256 -50498 39270 -50452
rect 33396 -50548 33884 -50542
rect 33396 -50582 33408 -50548
rect 33872 -50582 33884 -50548
rect 33396 -50588 33884 -50582
rect 34414 -50548 34902 -50542
rect 34414 -50582 34426 -50548
rect 34890 -50582 34902 -50548
rect 34414 -50588 34902 -50582
rect 35432 -50548 35920 -50542
rect 35432 -50582 35444 -50548
rect 35908 -50582 35920 -50548
rect 35432 -50588 35920 -50582
rect 36450 -50548 36938 -50542
rect 36450 -50582 36462 -50548
rect 36926 -50582 36938 -50548
rect 36450 -50588 36938 -50582
rect 37468 -50548 37956 -50542
rect 37468 -50582 37480 -50548
rect 37944 -50582 37956 -50548
rect 37468 -50588 37956 -50582
rect 38486 -50548 38974 -50542
rect 38486 -50582 38498 -50548
rect 38962 -50582 38974 -50548
rect 38486 -50588 38974 -50582
rect 33096 -50708 33102 -50648
rect 33162 -50708 33168 -50648
rect 30042 -51012 30048 -50952
rect 30108 -51012 30114 -50952
rect 29324 -51070 29812 -51064
rect 29324 -51104 29336 -51070
rect 29800 -51104 29812 -51070
rect 29324 -51110 29812 -51104
rect 29028 -51192 29042 -51154
rect 28058 -51730 28068 -51684
rect 29036 -51688 29042 -51192
rect 28008 -51892 28068 -51730
rect 29026 -51730 29042 -51688
rect 29076 -51192 29088 -51154
rect 30048 -51154 30108 -51012
rect 30342 -51070 30830 -51064
rect 30342 -51104 30354 -51070
rect 30818 -51104 30830 -51070
rect 30342 -51110 30830 -51104
rect 29076 -51688 29082 -51192
rect 30048 -51194 30060 -51154
rect 29076 -51730 29086 -51688
rect 28306 -51780 28794 -51774
rect 28306 -51814 28318 -51780
rect 28782 -51814 28794 -51780
rect 28306 -51820 28794 -51814
rect 28520 -51892 28580 -51820
rect 29026 -51892 29086 -51730
rect 30054 -51730 30060 -51194
rect 30094 -51194 30108 -51154
rect 31064 -51154 31124 -50912
rect 31566 -50918 31572 -50858
rect 31632 -50918 31638 -50858
rect 32588 -50918 32594 -50858
rect 32654 -50918 32660 -50858
rect 32076 -51012 32082 -50952
rect 32142 -51012 32148 -50952
rect 31360 -51070 31848 -51064
rect 31360 -51104 31372 -51070
rect 31836 -51104 31848 -51070
rect 31360 -51110 31848 -51104
rect 30094 -51730 30100 -51194
rect 31064 -51206 31078 -51154
rect 30054 -51742 30100 -51730
rect 31072 -51730 31078 -51206
rect 31112 -51206 31124 -51154
rect 32082 -51154 32142 -51012
rect 32594 -51064 32654 -50918
rect 32378 -51070 32866 -51064
rect 32378 -51104 32390 -51070
rect 32854 -51104 32866 -51070
rect 32378 -51110 32866 -51104
rect 32082 -51198 32096 -51154
rect 31112 -51730 31118 -51206
rect 32090 -51694 32096 -51198
rect 31072 -51742 31118 -51730
rect 32082 -51730 32096 -51694
rect 32130 -51198 32142 -51154
rect 33102 -51154 33162 -50708
rect 33608 -50858 33668 -50588
rect 34626 -50750 34686 -50588
rect 35646 -50638 35706 -50588
rect 36646 -50638 36706 -50588
rect 37684 -50638 37744 -50588
rect 38712 -50638 38772 -50588
rect 35128 -50708 35134 -50648
rect 35194 -50708 35200 -50648
rect 35646 -50698 38772 -50638
rect 34620 -50810 34626 -50750
rect 34686 -50810 34692 -50750
rect 33602 -50918 33608 -50858
rect 33668 -50918 33674 -50858
rect 34620 -50918 34626 -50858
rect 34686 -50918 34692 -50858
rect 33608 -51064 33668 -50918
rect 34112 -51012 34118 -50952
rect 34178 -51012 34184 -50952
rect 33396 -51070 33884 -51064
rect 33396 -51104 33408 -51070
rect 33872 -51104 33884 -51070
rect 33396 -51110 33884 -51104
rect 32130 -51694 32136 -51198
rect 32130 -51730 32142 -51694
rect 29324 -51780 29812 -51774
rect 29324 -51814 29336 -51780
rect 29800 -51814 29812 -51780
rect 29324 -51820 29812 -51814
rect 30342 -51780 30830 -51774
rect 30342 -51814 30354 -51780
rect 30818 -51814 30830 -51780
rect 30342 -51820 30830 -51814
rect 31360 -51780 31848 -51774
rect 31360 -51814 31372 -51780
rect 31836 -51814 31848 -51780
rect 31360 -51820 31848 -51814
rect 29530 -51876 29590 -51820
rect 28008 -51952 29086 -51892
rect 29524 -51936 29530 -51876
rect 29590 -51936 29596 -51876
rect 30434 -51936 30440 -51876
rect 30500 -51936 30506 -51876
rect 29524 -52152 29530 -52092
rect 29590 -52152 29596 -52092
rect 29530 -52158 29592 -52152
rect 27892 -52196 27954 -52190
rect 27892 -52256 27894 -52196
rect 27892 -52262 27954 -52256
rect 27776 -53022 27782 -52962
rect 27842 -53022 27848 -52962
rect 27326 -53380 27332 -53320
rect 27392 -53380 27398 -53320
rect 27564 -56906 27624 -53230
rect 27668 -53268 27674 -53208
rect 27734 -53268 27740 -53208
rect 27674 -55698 27734 -53268
rect 27780 -53564 27840 -53022
rect 27774 -53624 27780 -53564
rect 27840 -53624 27846 -53564
rect 27780 -55396 27840 -53624
rect 27892 -54440 27952 -52262
rect 29532 -52298 29592 -52158
rect 30440 -52298 30500 -51936
rect 30568 -52092 30628 -51820
rect 31436 -51936 31442 -51876
rect 31502 -51936 31508 -51876
rect 30568 -52158 30628 -52152
rect 31442 -52298 31502 -51936
rect 31582 -52092 31642 -51820
rect 32082 -51978 32142 -51730
rect 33102 -51730 33114 -51154
rect 33148 -51730 33162 -51154
rect 34118 -51154 34178 -51012
rect 34626 -51064 34686 -50918
rect 34414 -51070 34902 -51064
rect 34414 -51104 34426 -51070
rect 34890 -51104 34902 -51070
rect 34414 -51110 34902 -51104
rect 34118 -51190 34132 -51154
rect 32378 -51780 32866 -51774
rect 32378 -51814 32390 -51780
rect 32854 -51814 32866 -51780
rect 32378 -51820 32866 -51814
rect 32594 -51876 32654 -51820
rect 32588 -51936 32594 -51876
rect 32654 -51936 32660 -51876
rect 32076 -52038 32082 -51978
rect 32142 -52038 32148 -51978
rect 31576 -52152 31582 -52092
rect 31642 -52152 31648 -52092
rect 32594 -52298 32654 -51936
rect 28306 -52304 28794 -52298
rect 28306 -52338 28318 -52304
rect 28782 -52338 28794 -52304
rect 28306 -52344 28794 -52338
rect 29324 -52304 29812 -52298
rect 29324 -52338 29336 -52304
rect 29800 -52338 29812 -52304
rect 29324 -52344 29812 -52338
rect 30342 -52304 30830 -52298
rect 30342 -52338 30354 -52304
rect 30818 -52338 30830 -52304
rect 30342 -52344 30830 -52338
rect 31360 -52304 31848 -52298
rect 31360 -52338 31372 -52304
rect 31836 -52338 31848 -52304
rect 31360 -52344 31848 -52338
rect 32378 -52304 32866 -52298
rect 32378 -52338 32390 -52304
rect 32854 -52338 32866 -52304
rect 32378 -52344 32866 -52338
rect 28018 -52388 28064 -52376
rect 28018 -52926 28024 -52388
rect 28012 -52964 28024 -52926
rect 28058 -52926 28064 -52388
rect 29036 -52388 29082 -52376
rect 29036 -52926 29042 -52388
rect 28058 -52964 28072 -52926
rect 28012 -53094 28072 -52964
rect 29030 -52964 29042 -52926
rect 29076 -52926 29082 -52388
rect 30054 -52388 30100 -52376
rect 30054 -52914 30060 -52388
rect 29076 -52964 29090 -52926
rect 28306 -53014 28794 -53008
rect 28306 -53048 28318 -53014
rect 28782 -53048 28794 -53014
rect 28306 -53054 28794 -53048
rect 28510 -53094 28570 -53054
rect 29030 -53094 29090 -52964
rect 30046 -52964 30060 -52914
rect 30094 -52914 30100 -52388
rect 31072 -52388 31118 -52376
rect 31072 -52906 31078 -52388
rect 30094 -52964 30106 -52914
rect 29324 -53014 29812 -53008
rect 29324 -53048 29336 -53014
rect 29800 -53048 29812 -53014
rect 29324 -53054 29812 -53048
rect 28012 -53154 29090 -53094
rect 29030 -53208 29090 -53154
rect 29522 -53164 29528 -53104
rect 29588 -53164 29594 -53104
rect 29024 -53268 29030 -53208
rect 29090 -53268 29096 -53208
rect 29020 -53478 29026 -53418
rect 29086 -53478 29092 -53418
rect 28306 -53538 28794 -53532
rect 28306 -53572 28318 -53538
rect 28782 -53572 28794 -53538
rect 28306 -53578 28794 -53572
rect 28018 -53622 28064 -53610
rect 28018 -54164 28024 -53622
rect 28008 -54198 28024 -54164
rect 28058 -54164 28064 -53622
rect 29026 -53622 29086 -53478
rect 29528 -53532 29588 -53164
rect 30046 -53320 30106 -52964
rect 31064 -52964 31078 -52906
rect 31112 -52906 31118 -52388
rect 32090 -52388 32136 -52376
rect 31112 -52964 31124 -52906
rect 32090 -52918 32096 -52388
rect 30342 -53014 30830 -53008
rect 30342 -53048 30354 -53014
rect 30818 -53048 30830 -53014
rect 30342 -53054 30830 -53048
rect 30536 -53104 30596 -53054
rect 30530 -53164 30536 -53104
rect 30596 -53164 30602 -53104
rect 30040 -53380 30046 -53320
rect 30106 -53380 30112 -53320
rect 31064 -53418 31124 -52964
rect 32084 -52964 32096 -52918
rect 32130 -52918 32136 -52388
rect 33102 -52388 33162 -51730
rect 34126 -51730 34132 -51190
rect 34166 -51190 34178 -51154
rect 35134 -51154 35194 -50708
rect 35640 -50918 35646 -50858
rect 35706 -50918 35712 -50858
rect 38712 -50874 38772 -50698
rect 39210 -50764 39270 -50498
rect 40234 -50498 40240 -49966
rect 40274 -49966 40286 -49922
rect 41244 -49922 41304 -49452
rect 41746 -49710 41806 -49354
rect 42260 -49608 42320 -49264
rect 43280 -49264 43294 -49218
rect 43328 -48746 43342 -48688
rect 44306 -48688 44352 -48676
rect 43328 -49218 43334 -48746
rect 44306 -49208 44312 -48688
rect 43328 -49264 43340 -49218
rect 42558 -49314 43046 -49308
rect 42558 -49348 42570 -49314
rect 43034 -49348 43046 -49314
rect 42558 -49354 43046 -49348
rect 42254 -49668 42260 -49608
rect 42320 -49668 42326 -49608
rect 41744 -49716 41806 -49710
rect 41804 -49776 41806 -49716
rect 41744 -49782 41806 -49776
rect 42256 -49782 42262 -49722
rect 42322 -49782 42328 -49722
rect 41746 -49832 41806 -49782
rect 41540 -49838 42028 -49832
rect 41540 -49872 41552 -49838
rect 42016 -49872 42028 -49838
rect 41540 -49878 42028 -49872
rect 41244 -49966 41258 -49922
rect 40274 -50498 40280 -49966
rect 40234 -50510 40280 -50498
rect 41252 -50498 41258 -49966
rect 41292 -49966 41304 -49922
rect 42262 -49922 42322 -49782
rect 42770 -49832 42830 -49354
rect 43280 -49392 43340 -49264
rect 44298 -49264 44312 -49208
rect 44346 -49208 44352 -48688
rect 45324 -48688 45370 -48676
rect 44346 -49264 44358 -49208
rect 45324 -49220 45330 -48688
rect 43576 -49314 44064 -49308
rect 43576 -49348 43588 -49314
rect 44052 -49348 44064 -49314
rect 43576 -49354 44064 -49348
rect 43274 -49452 43280 -49392
rect 43340 -49452 43346 -49392
rect 42558 -49838 43046 -49832
rect 42558 -49872 42570 -49838
rect 43034 -49872 43046 -49838
rect 42558 -49878 43046 -49872
rect 42262 -49952 42276 -49922
rect 41292 -50498 41298 -49966
rect 42270 -50458 42276 -49952
rect 41252 -50510 41298 -50498
rect 42262 -50498 42276 -50458
rect 42310 -49952 42322 -49922
rect 43280 -49922 43340 -49452
rect 43796 -49832 43856 -49354
rect 44298 -49608 44358 -49264
rect 45314 -49264 45330 -49220
rect 45364 -49220 45370 -48688
rect 46342 -48688 46388 -48676
rect 46342 -49220 46348 -48688
rect 45364 -49264 45374 -49220
rect 44594 -49314 45082 -49308
rect 44594 -49348 44606 -49314
rect 45070 -49348 45082 -49314
rect 44594 -49354 45082 -49348
rect 44292 -49668 44298 -49608
rect 44358 -49668 44364 -49608
rect 44804 -49658 44864 -49354
rect 45314 -49500 45374 -49264
rect 46338 -49264 46348 -49220
rect 46382 -49220 46388 -48688
rect 47360 -48688 47406 -48676
rect 47360 -49214 47366 -48688
rect 46382 -49264 46398 -49220
rect 45612 -49314 46100 -49308
rect 45612 -49348 45624 -49314
rect 46088 -49348 46100 -49314
rect 45612 -49354 46100 -49348
rect 45820 -49498 45880 -49354
rect 45308 -49560 45314 -49500
rect 45374 -49560 45380 -49500
rect 45818 -49504 45880 -49498
rect 45878 -49564 45880 -49504
rect 45818 -49570 45880 -49564
rect 45820 -49658 45880 -49570
rect 46338 -49608 46398 -49264
rect 47354 -49264 47366 -49214
rect 47400 -49214 47406 -48688
rect 48370 -48688 48430 -48522
rect 48472 -48546 48478 -48486
rect 48538 -48546 48544 -48486
rect 48606 -48504 48666 -48216
rect 48370 -48716 48384 -48688
rect 48378 -49206 48384 -48716
rect 47400 -49264 47414 -49214
rect 46630 -49314 47118 -49308
rect 46630 -49348 46642 -49314
rect 47106 -49348 47118 -49314
rect 46630 -49354 47118 -49348
rect 44804 -49718 45880 -49658
rect 46332 -49668 46338 -49608
rect 46398 -49668 46404 -49608
rect 44292 -49782 44298 -49722
rect 44358 -49782 44364 -49722
rect 43576 -49838 44064 -49832
rect 43576 -49872 43588 -49838
rect 44052 -49872 44064 -49838
rect 43576 -49878 44064 -49872
rect 42310 -50458 42316 -49952
rect 43280 -49962 43294 -49922
rect 42310 -50498 42322 -50458
rect 43288 -50464 43294 -49962
rect 39504 -50548 39992 -50542
rect 39504 -50582 39516 -50548
rect 39980 -50582 39992 -50548
rect 39504 -50588 39992 -50582
rect 40522 -50548 41010 -50542
rect 40522 -50582 40534 -50548
rect 40998 -50582 41010 -50548
rect 40522 -50588 41010 -50582
rect 41540 -50548 42028 -50542
rect 41540 -50582 41552 -50548
rect 42016 -50582 42028 -50548
rect 41540 -50588 42028 -50582
rect 39716 -50636 39776 -50588
rect 39204 -50824 39210 -50764
rect 39270 -50824 39276 -50764
rect 39716 -50874 39776 -50696
rect 35646 -51064 35706 -50918
rect 38712 -50934 39776 -50874
rect 41240 -51022 41246 -50962
rect 41306 -51022 41312 -50962
rect 35432 -51070 35920 -51064
rect 35432 -51104 35444 -51070
rect 35908 -51104 35920 -51070
rect 35432 -51110 35920 -51104
rect 36450 -51070 36938 -51064
rect 36450 -51104 36462 -51070
rect 36926 -51104 36938 -51070
rect 36450 -51110 36938 -51104
rect 37468 -51070 37956 -51064
rect 37468 -51104 37480 -51070
rect 37944 -51104 37956 -51070
rect 37468 -51110 37956 -51104
rect 38486 -51070 38974 -51064
rect 38486 -51104 38498 -51070
rect 38962 -51104 38974 -51070
rect 38486 -51110 38974 -51104
rect 39504 -51070 39992 -51064
rect 39504 -51104 39516 -51070
rect 39980 -51104 39992 -51070
rect 39504 -51110 39992 -51104
rect 40522 -51070 41010 -51064
rect 40522 -51104 40534 -51070
rect 40998 -51104 41010 -51070
rect 40522 -51110 41010 -51104
rect 34166 -51730 34172 -51190
rect 35134 -51192 35150 -51154
rect 34126 -51742 34172 -51730
rect 35144 -51730 35150 -51192
rect 35184 -51192 35194 -51154
rect 36162 -51154 36208 -51142
rect 35184 -51730 35190 -51192
rect 36162 -51688 36168 -51154
rect 35144 -51742 35190 -51730
rect 36154 -51730 36168 -51688
rect 36202 -51688 36208 -51154
rect 37180 -51154 37226 -51142
rect 36202 -51730 36214 -51688
rect 37180 -51692 37186 -51154
rect 33396 -51780 33884 -51774
rect 33396 -51814 33408 -51780
rect 33872 -51814 33884 -51780
rect 33396 -51820 33884 -51814
rect 34414 -51780 34902 -51774
rect 34414 -51814 34426 -51780
rect 34890 -51814 34902 -51780
rect 34414 -51820 34902 -51814
rect 35432 -51780 35920 -51774
rect 35432 -51814 35444 -51780
rect 35908 -51814 35920 -51780
rect 35432 -51820 35920 -51814
rect 33604 -51876 33664 -51820
rect 34610 -51876 34670 -51820
rect 35654 -51876 35714 -51820
rect 36154 -51870 36214 -51730
rect 37174 -51730 37186 -51692
rect 37220 -51692 37226 -51154
rect 38198 -51154 38244 -51142
rect 37220 -51730 37234 -51692
rect 38198 -51698 38204 -51154
rect 36450 -51780 36938 -51774
rect 36450 -51814 36462 -51780
rect 36926 -51814 36938 -51780
rect 36450 -51820 36938 -51814
rect 33598 -51936 33604 -51876
rect 33664 -51936 33670 -51876
rect 34604 -51936 34610 -51876
rect 34670 -51936 34676 -51876
rect 35648 -51936 35654 -51876
rect 35714 -51936 35720 -51876
rect 36148 -51930 36154 -51870
rect 36214 -51930 36220 -51870
rect 33604 -52298 33664 -51936
rect 34602 -52152 34608 -52092
rect 34668 -52152 34674 -52092
rect 35642 -52152 35648 -52092
rect 35708 -52152 35714 -52092
rect 34608 -52298 34668 -52152
rect 35126 -52256 35132 -52196
rect 35192 -52256 35198 -52196
rect 33396 -52304 33884 -52298
rect 33396 -52338 33408 -52304
rect 33872 -52338 33884 -52304
rect 33396 -52344 33884 -52338
rect 34414 -52304 34902 -52298
rect 34414 -52338 34426 -52304
rect 34890 -52338 34902 -52304
rect 34414 -52344 34902 -52338
rect 33102 -52470 33114 -52388
rect 33108 -52918 33114 -52470
rect 32130 -52964 32144 -52918
rect 31360 -53014 31848 -53008
rect 31360 -53048 31372 -53014
rect 31836 -53048 31848 -53014
rect 31360 -53054 31848 -53048
rect 31550 -53104 31610 -53054
rect 31544 -53164 31550 -53104
rect 31610 -53164 31616 -53104
rect 32084 -53320 32144 -52964
rect 33104 -52964 33114 -52918
rect 33148 -52470 33162 -52388
rect 34126 -52388 34172 -52376
rect 33148 -52918 33154 -52470
rect 33148 -52964 33164 -52918
rect 34126 -52920 34132 -52388
rect 32378 -53014 32866 -53008
rect 32378 -53048 32390 -53014
rect 32854 -53048 32866 -53014
rect 32378 -53054 32866 -53048
rect 32588 -53104 32648 -53054
rect 32582 -53164 32588 -53104
rect 32648 -53164 32654 -53104
rect 32078 -53380 32084 -53320
rect 32144 -53380 32150 -53320
rect 31058 -53478 31064 -53418
rect 31124 -53478 31130 -53418
rect 32588 -53532 32648 -53164
rect 33104 -53418 33164 -52964
rect 34122 -52964 34132 -52920
rect 34166 -52920 34172 -52388
rect 35132 -52388 35192 -52256
rect 35648 -52298 35708 -52152
rect 35432 -52304 35920 -52298
rect 35432 -52338 35444 -52304
rect 35908 -52338 35920 -52304
rect 35432 -52344 35920 -52338
rect 35132 -52452 35150 -52388
rect 34166 -52964 34182 -52920
rect 33396 -53014 33884 -53008
rect 33396 -53048 33408 -53014
rect 33872 -53048 33884 -53014
rect 33396 -53054 33884 -53048
rect 33606 -53104 33666 -53054
rect 34122 -53098 34182 -52964
rect 35144 -52964 35150 -52452
rect 35184 -52452 35192 -52388
rect 36154 -52388 36214 -51930
rect 36662 -52092 36722 -51820
rect 36656 -52152 36662 -52092
rect 36722 -52152 36728 -52092
rect 36662 -52298 36722 -52152
rect 37174 -52196 37234 -51730
rect 38190 -51730 38204 -51698
rect 38238 -51698 38244 -51154
rect 39216 -51154 39262 -51142
rect 39216 -51696 39222 -51154
rect 38238 -51730 38250 -51698
rect 37468 -51780 37956 -51774
rect 37468 -51814 37480 -51780
rect 37944 -51814 37956 -51780
rect 37468 -51820 37956 -51814
rect 37670 -52092 37730 -51820
rect 38190 -51870 38250 -51730
rect 39212 -51730 39222 -51696
rect 39256 -51696 39262 -51154
rect 40234 -51154 40280 -51142
rect 39256 -51730 39272 -51696
rect 40234 -51698 40240 -51154
rect 38486 -51780 38974 -51774
rect 38486 -51814 38498 -51780
rect 38962 -51814 38974 -51780
rect 38486 -51820 38974 -51814
rect 38184 -51930 38190 -51870
rect 38250 -51930 38256 -51870
rect 38714 -52092 38774 -51820
rect 37664 -52152 37670 -52092
rect 37730 -52152 37736 -52092
rect 38708 -52152 38714 -52092
rect 38774 -52152 38780 -52092
rect 37168 -52256 37174 -52196
rect 37234 -52256 37240 -52196
rect 36450 -52304 36938 -52298
rect 36450 -52338 36462 -52304
rect 36926 -52338 36938 -52304
rect 36450 -52344 36938 -52338
rect 36154 -52424 36168 -52388
rect 35184 -52964 35190 -52452
rect 36162 -52906 36168 -52424
rect 35144 -52976 35190 -52964
rect 36158 -52964 36168 -52906
rect 36202 -52424 36214 -52388
rect 37174 -52388 37234 -52256
rect 37670 -52298 37730 -52152
rect 38714 -52298 38774 -52152
rect 39212 -52196 39272 -51730
rect 40226 -51730 40240 -51698
rect 40274 -51698 40280 -51154
rect 41246 -51154 41306 -51022
rect 41540 -51070 42028 -51064
rect 41540 -51104 41552 -51070
rect 42016 -51104 42028 -51070
rect 41540 -51110 42028 -51104
rect 40274 -51730 40286 -51698
rect 39504 -51780 39992 -51774
rect 39504 -51814 39516 -51780
rect 39980 -51814 39992 -51780
rect 39504 -51820 39992 -51814
rect 39704 -52092 39764 -51820
rect 40226 -51870 40286 -51730
rect 41246 -51730 41258 -51154
rect 41292 -51730 41306 -51154
rect 42262 -51154 42322 -50498
rect 43282 -50498 43294 -50464
rect 43328 -49962 43340 -49922
rect 44298 -49922 44358 -49782
rect 44804 -49832 44864 -49718
rect 45820 -49832 45880 -49718
rect 46330 -49782 46336 -49722
rect 46396 -49782 46402 -49722
rect 44594 -49838 45082 -49832
rect 44594 -49872 44606 -49838
rect 45070 -49872 45082 -49838
rect 44594 -49878 45082 -49872
rect 45612 -49838 46100 -49832
rect 45612 -49872 45624 -49838
rect 46088 -49872 46100 -49838
rect 45612 -49878 46100 -49872
rect 43328 -50464 43334 -49962
rect 44298 -49964 44312 -49922
rect 43328 -50498 43342 -50464
rect 42558 -50548 43046 -50542
rect 42558 -50582 42570 -50548
rect 43034 -50582 43046 -50548
rect 42558 -50588 43046 -50582
rect 42758 -50858 42818 -50588
rect 42752 -50918 42758 -50858
rect 42818 -50918 42824 -50858
rect 42758 -51064 42818 -50918
rect 42558 -51070 43046 -51064
rect 42558 -51104 42570 -51070
rect 43034 -51104 43046 -51070
rect 42558 -51110 43046 -51104
rect 42262 -51194 42276 -51154
rect 42270 -51698 42276 -51194
rect 40522 -51780 41010 -51774
rect 40522 -51814 40534 -51780
rect 40998 -51814 41010 -51780
rect 40522 -51820 41010 -51814
rect 40220 -51930 40226 -51870
rect 40286 -51930 40292 -51870
rect 40722 -52092 40782 -51820
rect 39698 -52152 39704 -52092
rect 39764 -52152 39770 -52092
rect 40716 -52152 40722 -52092
rect 40782 -52152 40788 -52092
rect 39206 -52256 39212 -52196
rect 39272 -52256 39278 -52196
rect 37468 -52304 37956 -52298
rect 37468 -52338 37480 -52304
rect 37944 -52338 37956 -52304
rect 37468 -52344 37956 -52338
rect 38486 -52304 38974 -52298
rect 38486 -52338 38498 -52304
rect 38962 -52338 38974 -52304
rect 38486 -52344 38974 -52338
rect 36202 -52906 36208 -52424
rect 37174 -52426 37186 -52388
rect 36202 -52964 36218 -52906
rect 34414 -53014 34902 -53008
rect 34414 -53048 34426 -53014
rect 34890 -53048 34902 -53014
rect 34414 -53054 34902 -53048
rect 35432 -53014 35920 -53008
rect 35432 -53048 35444 -53014
rect 35908 -53048 35920 -53014
rect 35432 -53054 35920 -53048
rect 36158 -53098 36218 -52964
rect 37180 -52964 37186 -52426
rect 37220 -52426 37234 -52388
rect 38198 -52388 38244 -52376
rect 37220 -52964 37226 -52426
rect 38198 -52914 38204 -52388
rect 37180 -52976 37226 -52964
rect 38190 -52964 38204 -52914
rect 38238 -52914 38244 -52388
rect 39212 -52388 39272 -52256
rect 39704 -52298 39764 -52152
rect 41246 -52196 41306 -51730
rect 42264 -51730 42276 -51698
rect 42310 -51194 42322 -51154
rect 43282 -51154 43342 -50498
rect 44306 -50498 44312 -49964
rect 44346 -49964 44358 -49922
rect 45324 -49922 45370 -49910
rect 44346 -50498 44352 -49964
rect 45324 -50440 45330 -49922
rect 44306 -50510 44352 -50498
rect 45316 -50498 45330 -50440
rect 45364 -50440 45370 -49922
rect 46336 -49922 46396 -49782
rect 46838 -49832 46898 -49354
rect 47354 -49392 47414 -49264
rect 48372 -49264 48384 -49206
rect 48418 -48716 48430 -48688
rect 48418 -49206 48424 -48716
rect 48418 -49264 48432 -49206
rect 47648 -49314 48136 -49308
rect 47648 -49348 47660 -49314
rect 48124 -49348 48136 -49314
rect 47648 -49354 48136 -49348
rect 48372 -49374 48432 -49264
rect 47348 -49452 47354 -49392
rect 47414 -49452 47420 -49392
rect 48366 -49434 48372 -49374
rect 48432 -49434 48438 -49374
rect 47354 -49670 47414 -49452
rect 47354 -49730 48428 -49670
rect 48478 -49722 48538 -48546
rect 48600 -48564 48606 -48504
rect 48666 -48564 48672 -48504
rect 48972 -49504 49032 -45618
rect 48966 -49564 48972 -49504
rect 49032 -49564 49038 -49504
rect 48716 -49668 48722 -49608
rect 48782 -49668 48788 -49608
rect 46630 -49838 47118 -49832
rect 46630 -49872 46642 -49838
rect 47106 -49872 47118 -49838
rect 46630 -49878 47118 -49872
rect 46336 -49964 46348 -49922
rect 45364 -50498 45376 -50440
rect 43788 -50542 43848 -50540
rect 43576 -50548 44064 -50542
rect 43576 -50582 43588 -50548
rect 44052 -50582 44064 -50548
rect 43576 -50588 44064 -50582
rect 44594 -50548 45082 -50542
rect 44594 -50582 44606 -50548
rect 45070 -50582 45082 -50548
rect 44594 -50588 45082 -50582
rect 43788 -50858 43848 -50588
rect 44810 -50636 44870 -50588
rect 44804 -50696 44810 -50636
rect 44870 -50696 44876 -50636
rect 44942 -50692 44948 -50632
rect 45008 -50692 45014 -50632
rect 44948 -50858 45008 -50692
rect 45316 -50858 45376 -50498
rect 46342 -50498 46348 -49964
rect 46382 -49964 46396 -49922
rect 47354 -49922 47414 -49730
rect 47858 -49832 47918 -49730
rect 47648 -49838 48136 -49832
rect 47648 -49872 47660 -49838
rect 48124 -49872 48136 -49838
rect 47648 -49878 48136 -49872
rect 47354 -49956 47366 -49922
rect 46382 -50498 46388 -49964
rect 47360 -50458 47366 -49956
rect 46342 -50510 46388 -50498
rect 47354 -50498 47366 -50458
rect 47400 -49956 47414 -49922
rect 48368 -49922 48428 -49730
rect 48472 -49782 48478 -49722
rect 48538 -49782 48544 -49722
rect 48368 -49946 48384 -49922
rect 47400 -50458 47406 -49956
rect 47400 -50498 47414 -50458
rect 45612 -50548 46100 -50542
rect 45612 -50582 45624 -50548
rect 46088 -50582 46100 -50548
rect 45612 -50588 46100 -50582
rect 46630 -50548 47118 -50542
rect 46630 -50582 46642 -50548
rect 47106 -50582 47118 -50548
rect 46630 -50588 47118 -50582
rect 46836 -50632 46896 -50588
rect 45824 -50692 45830 -50632
rect 45890 -50692 45896 -50632
rect 46830 -50692 46836 -50632
rect 46896 -50692 46902 -50632
rect 47354 -50636 47414 -50498
rect 48378 -50498 48384 -49946
rect 48418 -49946 48428 -49922
rect 48418 -50498 48424 -49946
rect 48378 -50510 48424 -50498
rect 47648 -50548 48136 -50542
rect 47648 -50582 47660 -50548
rect 48124 -50582 48136 -50548
rect 47648 -50588 48136 -50582
rect 43782 -50918 43788 -50858
rect 43848 -50918 43854 -50858
rect 44942 -50918 44948 -50858
rect 45008 -50918 45014 -50858
rect 45310 -50918 45316 -50858
rect 45376 -50918 45382 -50858
rect 43788 -51064 43848 -50918
rect 44948 -51064 45008 -50918
rect 45316 -50962 45376 -50918
rect 45310 -51022 45316 -50962
rect 45376 -51022 45382 -50962
rect 45830 -51064 45890 -50692
rect 47348 -50696 47354 -50636
rect 47414 -50696 47420 -50636
rect 47348 -50824 47354 -50764
rect 47414 -50824 47420 -50764
rect 46326 -51020 46332 -50960
rect 46392 -51020 46398 -50960
rect 43576 -51070 44064 -51064
rect 43576 -51104 43588 -51070
rect 44052 -51104 44064 -51070
rect 43576 -51110 44064 -51104
rect 44594 -51070 45082 -51064
rect 44594 -51104 44606 -51070
rect 45070 -51104 45082 -51070
rect 44594 -51110 45082 -51104
rect 45612 -51070 46100 -51064
rect 45612 -51104 45624 -51070
rect 46088 -51104 46100 -51070
rect 45612 -51110 46100 -51104
rect 45830 -51112 45890 -51110
rect 42310 -51698 42316 -51194
rect 43282 -51200 43294 -51154
rect 43288 -51686 43294 -51200
rect 42310 -51730 42324 -51698
rect 41540 -51780 42028 -51774
rect 41540 -51814 41552 -51780
rect 42016 -51814 42028 -51780
rect 41540 -51820 42028 -51814
rect 41756 -52092 41816 -51820
rect 42264 -51870 42324 -51730
rect 43280 -51730 43294 -51686
rect 43328 -51200 43342 -51154
rect 44306 -51154 44352 -51142
rect 43328 -51686 43334 -51200
rect 43328 -51730 43340 -51686
rect 44306 -51690 44312 -51154
rect 42558 -51780 43046 -51774
rect 42558 -51814 42570 -51780
rect 43034 -51814 43046 -51780
rect 42558 -51820 43046 -51814
rect 42258 -51930 42264 -51870
rect 42324 -51930 42330 -51870
rect 42250 -52038 42256 -51978
rect 42316 -52038 42322 -51978
rect 41750 -52152 41756 -52092
rect 41816 -52152 41822 -52092
rect 41240 -52256 41246 -52196
rect 41306 -52256 41312 -52196
rect 41752 -52260 41758 -52200
rect 41818 -52260 41824 -52200
rect 41758 -52298 41818 -52260
rect 39504 -52304 39992 -52298
rect 39504 -52338 39516 -52304
rect 39980 -52338 39992 -52304
rect 39504 -52344 39992 -52338
rect 40522 -52304 41010 -52298
rect 40522 -52338 40534 -52304
rect 40998 -52338 41010 -52304
rect 40522 -52344 41010 -52338
rect 41540 -52304 42028 -52298
rect 41540 -52338 41552 -52304
rect 42016 -52338 42028 -52304
rect 41540 -52344 42028 -52338
rect 39212 -52424 39222 -52388
rect 38238 -52964 38250 -52914
rect 36450 -53014 36938 -53008
rect 36450 -53048 36462 -53014
rect 36926 -53048 36938 -53014
rect 36450 -53054 36938 -53048
rect 37468 -53014 37956 -53008
rect 37468 -53048 37480 -53014
rect 37944 -53048 37956 -53014
rect 37468 -53054 37956 -53048
rect 38190 -53098 38250 -52964
rect 39216 -52964 39222 -52424
rect 39256 -52424 39272 -52388
rect 40234 -52388 40280 -52376
rect 39256 -52964 39262 -52424
rect 40234 -52902 40240 -52388
rect 39216 -52976 39262 -52964
rect 40224 -52964 40240 -52902
rect 40274 -52902 40280 -52388
rect 41252 -52388 41298 -52376
rect 40274 -52964 40284 -52902
rect 41252 -52922 41258 -52388
rect 38486 -53014 38974 -53008
rect 38486 -53048 38498 -53014
rect 38962 -53048 38974 -53014
rect 38486 -53054 38974 -53048
rect 39504 -53014 39992 -53008
rect 39504 -53048 39516 -53014
rect 39980 -53048 39992 -53014
rect 39504 -53054 39992 -53048
rect 40224 -53098 40284 -52964
rect 41246 -52964 41258 -52922
rect 41292 -52922 41298 -52388
rect 42256 -52388 42316 -52038
rect 42780 -52200 42840 -51820
rect 43280 -52194 43340 -51730
rect 44300 -51730 44312 -51690
rect 44346 -51690 44352 -51154
rect 45324 -51154 45370 -51142
rect 45324 -51686 45330 -51154
rect 44346 -51730 44360 -51690
rect 43576 -51780 44064 -51774
rect 43576 -51814 43588 -51780
rect 44052 -51814 44064 -51780
rect 43576 -51820 44064 -51814
rect 42774 -52260 42780 -52200
rect 42840 -52260 42846 -52200
rect 43274 -52254 43280 -52194
rect 43340 -52254 43346 -52194
rect 42780 -52298 42840 -52260
rect 42558 -52304 43046 -52298
rect 42558 -52338 42570 -52304
rect 43034 -52338 43046 -52304
rect 42558 -52344 43046 -52338
rect 42256 -52424 42276 -52388
rect 41292 -52964 41306 -52922
rect 40522 -53014 41010 -53008
rect 40522 -53048 40534 -53014
rect 40998 -53048 41010 -53014
rect 40522 -53054 41010 -53048
rect 33600 -53164 33606 -53104
rect 33666 -53164 33672 -53104
rect 34116 -53158 34122 -53098
rect 34182 -53158 34188 -53098
rect 38184 -53158 38190 -53098
rect 38250 -53158 38256 -53098
rect 40218 -53158 40224 -53098
rect 40284 -53158 40290 -53098
rect 33098 -53478 33104 -53418
rect 33164 -53478 33170 -53418
rect 29324 -53538 29812 -53532
rect 29324 -53572 29336 -53538
rect 29800 -53572 29812 -53538
rect 29324 -53578 29812 -53572
rect 30342 -53538 30830 -53532
rect 30342 -53572 30354 -53538
rect 30818 -53572 30830 -53538
rect 30342 -53578 30830 -53572
rect 31360 -53538 31848 -53532
rect 31360 -53572 31372 -53538
rect 31836 -53572 31848 -53538
rect 31360 -53578 31848 -53572
rect 32378 -53538 32866 -53532
rect 32378 -53572 32390 -53538
rect 32854 -53572 32866 -53538
rect 32378 -53578 32866 -53572
rect 29026 -53676 29042 -53622
rect 28058 -54198 28068 -54164
rect 29036 -54168 29042 -53676
rect 28008 -54330 28068 -54198
rect 29032 -54198 29042 -54168
rect 29076 -53676 29086 -53622
rect 30054 -53622 30100 -53610
rect 29076 -54168 29082 -53676
rect 30054 -54152 30060 -53622
rect 29076 -54198 29092 -54168
rect 28306 -54248 28794 -54242
rect 28306 -54282 28318 -54248
rect 28782 -54282 28794 -54248
rect 28306 -54288 28794 -54282
rect 28528 -54330 28588 -54288
rect 29032 -54330 29092 -54198
rect 30046 -54198 30060 -54152
rect 30094 -54152 30100 -53622
rect 31072 -53622 31118 -53610
rect 30094 -54198 30106 -54152
rect 31072 -54168 31078 -53622
rect 29324 -54248 29812 -54242
rect 29324 -54282 29336 -54248
rect 29800 -54282 29812 -54248
rect 29324 -54288 29812 -54282
rect 28008 -54390 29092 -54330
rect 27886 -54500 27892 -54440
rect 27952 -54500 27958 -54440
rect 29032 -54536 29092 -54390
rect 28008 -54596 29092 -54536
rect 28008 -54854 28068 -54596
rect 28520 -54764 28580 -54596
rect 29032 -54656 29092 -54596
rect 29026 -54716 29032 -54656
rect 29092 -54716 29098 -54656
rect 28306 -54770 28794 -54764
rect 28306 -54804 28318 -54770
rect 28782 -54804 28794 -54770
rect 28306 -54810 28794 -54804
rect 28008 -54890 28024 -54854
rect 27774 -55456 27780 -55396
rect 27840 -55456 27846 -55396
rect 28018 -55430 28024 -54890
rect 28058 -54890 28068 -54854
rect 29032 -54854 29092 -54716
rect 29524 -54764 29584 -54288
rect 30046 -54342 30106 -54198
rect 31064 -54198 31078 -54168
rect 31112 -54168 31118 -53622
rect 32090 -53622 32136 -53610
rect 32090 -54156 32096 -53622
rect 31112 -54198 31124 -54168
rect 30342 -54248 30830 -54242
rect 30342 -54282 30354 -54248
rect 30818 -54282 30830 -54248
rect 30342 -54288 30830 -54282
rect 30040 -54402 30046 -54342
rect 30106 -54402 30112 -54342
rect 30044 -54596 30050 -54536
rect 30110 -54596 30116 -54536
rect 29324 -54770 29812 -54764
rect 29324 -54804 29336 -54770
rect 29800 -54804 29812 -54770
rect 29324 -54810 29812 -54804
rect 28058 -55430 28064 -54890
rect 29032 -54894 29042 -54854
rect 28018 -55442 28064 -55430
rect 29036 -55430 29042 -54894
rect 29076 -54894 29092 -54854
rect 30050 -54854 30110 -54596
rect 30544 -54600 30604 -54288
rect 31064 -54440 31124 -54198
rect 32082 -54198 32096 -54156
rect 32130 -54156 32136 -53622
rect 33104 -53622 33164 -53478
rect 33606 -53532 33666 -53164
rect 33396 -53538 33884 -53532
rect 33396 -53572 33408 -53538
rect 33872 -53572 33884 -53538
rect 33396 -53578 33884 -53572
rect 33104 -53652 33114 -53622
rect 33108 -54134 33114 -53652
rect 32130 -54198 32142 -54156
rect 31360 -54248 31848 -54242
rect 31360 -54282 31372 -54248
rect 31836 -54282 31848 -54248
rect 31360 -54288 31848 -54282
rect 31058 -54500 31064 -54440
rect 31124 -54500 31130 -54440
rect 31578 -54600 31638 -54288
rect 32082 -54342 32142 -54198
rect 33100 -54198 33114 -54134
rect 33148 -53652 33164 -53622
rect 34122 -53622 34182 -53158
rect 36158 -53164 36218 -53158
rect 37168 -53268 37174 -53208
rect 37234 -53268 37240 -53208
rect 39204 -53268 39210 -53208
rect 39270 -53268 39276 -53208
rect 36150 -53380 36156 -53320
rect 36216 -53380 36222 -53320
rect 35134 -53478 35140 -53418
rect 35200 -53478 35206 -53418
rect 34414 -53538 34902 -53532
rect 34414 -53572 34426 -53538
rect 34890 -53572 34902 -53538
rect 34414 -53578 34902 -53572
rect 33148 -54134 33154 -53652
rect 34122 -53664 34132 -53622
rect 33148 -54198 33160 -54134
rect 34126 -54158 34132 -53664
rect 32378 -54248 32866 -54242
rect 32378 -54282 32390 -54248
rect 32854 -54282 32866 -54248
rect 32378 -54288 32866 -54282
rect 32076 -54402 32082 -54342
rect 32142 -54402 32148 -54342
rect 32588 -54440 32648 -54288
rect 32582 -54500 32588 -54440
rect 32648 -54500 32654 -54440
rect 32080 -54596 32086 -54536
rect 32146 -54596 32152 -54536
rect 30544 -54660 31638 -54600
rect 30544 -54764 30604 -54660
rect 31578 -54764 31638 -54660
rect 30342 -54770 30830 -54764
rect 30342 -54804 30354 -54770
rect 30818 -54804 30830 -54770
rect 30342 -54810 30830 -54804
rect 31360 -54770 31848 -54764
rect 31360 -54804 31372 -54770
rect 31836 -54804 31848 -54770
rect 31360 -54810 31848 -54804
rect 29076 -55430 29082 -54894
rect 30050 -54898 30060 -54854
rect 29036 -55442 29082 -55430
rect 30054 -55430 30060 -54898
rect 30094 -54898 30110 -54854
rect 31072 -54854 31118 -54842
rect 30094 -55430 30100 -54898
rect 31072 -55388 31078 -54854
rect 30054 -55442 30100 -55430
rect 31064 -55430 31078 -55388
rect 31112 -55388 31118 -54854
rect 32086 -54854 32146 -54596
rect 32588 -54764 32648 -54500
rect 33100 -54656 33160 -54198
rect 34120 -54198 34132 -54158
rect 34166 -53664 34182 -53622
rect 35140 -53622 35200 -53478
rect 35432 -53538 35920 -53532
rect 35432 -53572 35444 -53538
rect 35908 -53572 35920 -53538
rect 35432 -53578 35920 -53572
rect 35140 -53658 35150 -53622
rect 34166 -54158 34172 -53664
rect 34166 -54198 34180 -54158
rect 35144 -54164 35150 -53658
rect 33396 -54248 33884 -54242
rect 33396 -54282 33408 -54248
rect 33872 -54282 33884 -54248
rect 33396 -54288 33884 -54282
rect 33610 -54440 33670 -54288
rect 34120 -54342 34180 -54198
rect 35134 -54198 35150 -54164
rect 35184 -53658 35200 -53622
rect 36156 -53622 36216 -53380
rect 36450 -53538 36938 -53532
rect 36450 -53572 36462 -53538
rect 36926 -53572 36938 -53538
rect 36450 -53578 36938 -53572
rect 36156 -53648 36168 -53622
rect 35184 -54164 35190 -53658
rect 36162 -54142 36168 -53648
rect 35184 -54198 35194 -54164
rect 34414 -54248 34902 -54242
rect 34414 -54282 34426 -54248
rect 34890 -54282 34902 -54248
rect 34414 -54288 34902 -54282
rect 34114 -54402 34120 -54342
rect 34180 -54402 34186 -54342
rect 34634 -54434 34694 -54288
rect 33094 -54716 33100 -54656
rect 33160 -54716 33166 -54656
rect 32378 -54770 32866 -54764
rect 32378 -54804 32390 -54770
rect 32854 -54804 32866 -54770
rect 32378 -54810 32866 -54804
rect 32086 -54906 32096 -54854
rect 31112 -55430 31124 -55388
rect 27780 -55572 27840 -55456
rect 28306 -55480 28794 -55474
rect 28306 -55514 28318 -55480
rect 28782 -55514 28794 -55480
rect 28306 -55520 28794 -55514
rect 29324 -55480 29812 -55474
rect 29324 -55514 29336 -55480
rect 29800 -55514 29812 -55480
rect 29324 -55520 29812 -55514
rect 30342 -55480 30830 -55474
rect 30342 -55514 30354 -55480
rect 30818 -55514 30830 -55480
rect 30342 -55520 30830 -55514
rect 27774 -55632 27780 -55572
rect 27840 -55632 27846 -55572
rect 27668 -55758 27674 -55698
rect 27734 -55758 27740 -55698
rect 28008 -55938 29088 -55878
rect 28008 -56088 28068 -55938
rect 28516 -55998 28576 -55938
rect 28306 -56004 28794 -55998
rect 28306 -56038 28318 -56004
rect 28782 -56038 28794 -56004
rect 28306 -56044 28794 -56038
rect 28008 -56144 28024 -56088
rect 28018 -56664 28024 -56144
rect 28058 -56144 28068 -56088
rect 29028 -56088 29088 -55938
rect 29526 -55998 29586 -55520
rect 31064 -55698 31124 -55430
rect 32090 -55430 32096 -54906
rect 32130 -54906 32146 -54854
rect 33100 -54854 33160 -54716
rect 33610 -54764 33670 -54500
rect 34632 -54440 34694 -54434
rect 34692 -54500 34694 -54440
rect 34632 -54506 34694 -54500
rect 34108 -54596 34114 -54536
rect 34174 -54596 34180 -54536
rect 33396 -54770 33884 -54764
rect 33396 -54804 33408 -54770
rect 33872 -54804 33884 -54770
rect 33396 -54810 33884 -54804
rect 33100 -54894 33114 -54854
rect 32130 -55430 32136 -54906
rect 33108 -55376 33114 -54894
rect 32090 -55442 32136 -55430
rect 33102 -55430 33114 -55376
rect 33148 -54894 33160 -54854
rect 34114 -54854 34174 -54596
rect 34634 -54764 34694 -54506
rect 35134 -54656 35194 -54198
rect 36152 -54198 36168 -54142
rect 36202 -53648 36216 -53622
rect 37174 -53622 37234 -53268
rect 37468 -53538 37956 -53532
rect 37468 -53572 37480 -53538
rect 37944 -53572 37956 -53538
rect 37468 -53578 37956 -53572
rect 38486 -53538 38974 -53532
rect 38486 -53572 38498 -53538
rect 38962 -53572 38974 -53538
rect 38486 -53578 38974 -53572
rect 36202 -54142 36208 -53648
rect 37174 -53654 37186 -53622
rect 36202 -54198 36212 -54142
rect 35432 -54248 35920 -54242
rect 35432 -54282 35444 -54248
rect 35908 -54282 35920 -54248
rect 35432 -54288 35920 -54282
rect 35636 -54440 35696 -54288
rect 35982 -54322 36042 -54316
rect 36152 -54322 36212 -54198
rect 37180 -54198 37186 -53654
rect 37220 -53654 37234 -53622
rect 38198 -53622 38244 -53610
rect 37220 -54198 37226 -53654
rect 38198 -54128 38204 -53622
rect 37180 -54210 37226 -54198
rect 38194 -54198 38204 -54128
rect 38238 -54128 38244 -53622
rect 39210 -53622 39270 -53268
rect 40752 -53306 40812 -53054
rect 41246 -53096 41306 -52964
rect 42270 -52964 42276 -52424
rect 42310 -52964 42316 -52388
rect 43280 -52388 43340 -52254
rect 43758 -52298 43818 -51820
rect 44300 -51870 44360 -51730
rect 45314 -51730 45330 -51686
rect 45364 -51686 45370 -51154
rect 46332 -51154 46392 -51020
rect 46630 -51070 47118 -51064
rect 46630 -51104 46642 -51070
rect 47106 -51104 47118 -51070
rect 46630 -51110 47118 -51104
rect 46332 -51204 46348 -51154
rect 45364 -51730 45374 -51686
rect 46342 -51702 46348 -51204
rect 44594 -51780 45082 -51774
rect 44594 -51814 44606 -51780
rect 45070 -51814 45082 -51780
rect 44594 -51820 45082 -51814
rect 44294 -51930 44300 -51870
rect 44360 -51930 44366 -51870
rect 44290 -52038 44296 -51978
rect 44356 -52038 44362 -51978
rect 43576 -52304 44064 -52298
rect 43576 -52338 43588 -52304
rect 44052 -52338 44064 -52304
rect 43576 -52344 44064 -52338
rect 43280 -52482 43294 -52388
rect 43288 -52922 43294 -52482
rect 42270 -52976 42316 -52964
rect 43280 -52964 43294 -52922
rect 43328 -52482 43340 -52388
rect 44296 -52388 44356 -52038
rect 44782 -52152 44788 -52092
rect 44848 -52152 44854 -52092
rect 44788 -52298 44848 -52152
rect 45314 -52194 45374 -51730
rect 46338 -51730 46348 -51702
rect 46382 -51204 46392 -51154
rect 47354 -51154 47414 -50824
rect 47648 -51070 48136 -51064
rect 47648 -51104 47660 -51070
rect 48124 -51104 48136 -51070
rect 47648 -51110 48136 -51104
rect 46382 -51702 46388 -51204
rect 47354 -51206 47366 -51154
rect 47360 -51702 47366 -51206
rect 46382 -51730 46398 -51702
rect 45612 -51780 46100 -51774
rect 45612 -51814 45624 -51780
rect 46088 -51814 46100 -51780
rect 45612 -51820 46100 -51814
rect 46338 -51870 46398 -51730
rect 47354 -51730 47366 -51702
rect 47400 -51206 47414 -51154
rect 48378 -51154 48424 -51142
rect 47400 -51702 47406 -51206
rect 48378 -51696 48384 -51154
rect 47400 -51730 47414 -51702
rect 46630 -51780 47118 -51774
rect 46630 -51814 46642 -51780
rect 47106 -51814 47118 -51780
rect 46630 -51820 47118 -51814
rect 46332 -51930 46338 -51870
rect 46398 -51930 46404 -51870
rect 46328 -52038 46334 -51978
rect 46394 -52038 46400 -51978
rect 45820 -52152 45826 -52092
rect 45886 -52152 45892 -52092
rect 45308 -52254 45314 -52194
rect 45374 -52254 45380 -52194
rect 45826 -52298 45886 -52152
rect 44594 -52304 45082 -52298
rect 44594 -52338 44606 -52304
rect 45070 -52338 45082 -52304
rect 44594 -52344 45082 -52338
rect 45612 -52304 46100 -52298
rect 45612 -52338 45624 -52304
rect 46088 -52338 46100 -52304
rect 45612 -52344 46100 -52338
rect 44296 -52454 44312 -52388
rect 43328 -52922 43334 -52482
rect 43328 -52964 43340 -52922
rect 41540 -53014 42028 -53008
rect 41540 -53048 41552 -53014
rect 42016 -53048 42028 -53014
rect 41540 -53054 42028 -53048
rect 42558 -53014 43046 -53008
rect 42558 -53048 42570 -53014
rect 43034 -53048 43046 -53014
rect 42558 -53054 43046 -53048
rect 41240 -53156 41246 -53096
rect 41306 -53156 41312 -53096
rect 41594 -53156 41600 -53096
rect 41660 -53156 41666 -53096
rect 41236 -53268 41242 -53208
rect 41302 -53268 41308 -53208
rect 40746 -53366 40752 -53306
rect 40812 -53366 40818 -53306
rect 39504 -53538 39992 -53532
rect 39504 -53572 39516 -53538
rect 39980 -53572 39992 -53538
rect 39504 -53578 39992 -53572
rect 40522 -53538 41010 -53532
rect 40522 -53572 40534 -53538
rect 40998 -53572 41010 -53538
rect 40522 -53578 41010 -53572
rect 39210 -53660 39222 -53622
rect 38238 -54198 38254 -54128
rect 36450 -54248 36938 -54242
rect 36450 -54282 36462 -54248
rect 36926 -54282 36938 -54248
rect 36450 -54288 36938 -54282
rect 37468 -54248 37956 -54242
rect 37468 -54282 37480 -54248
rect 37944 -54282 37956 -54248
rect 37468 -54288 37956 -54282
rect 36146 -54382 36152 -54322
rect 36212 -54382 36218 -54322
rect 35630 -54500 35636 -54440
rect 35696 -54500 35702 -54440
rect 35128 -54716 35134 -54656
rect 35194 -54716 35200 -54656
rect 34414 -54770 34902 -54764
rect 34414 -54804 34426 -54770
rect 34890 -54804 34902 -54770
rect 34414 -54810 34902 -54804
rect 33148 -55376 33154 -54894
rect 34114 -54914 34132 -54854
rect 33148 -55430 33162 -55376
rect 31360 -55480 31848 -55474
rect 31360 -55514 31372 -55480
rect 31836 -55514 31848 -55480
rect 31360 -55520 31848 -55514
rect 32378 -55480 32866 -55474
rect 32378 -55514 32390 -55480
rect 32854 -55514 32866 -55480
rect 32378 -55520 32866 -55514
rect 31584 -55686 31644 -55520
rect 31058 -55758 31064 -55698
rect 31124 -55758 31130 -55698
rect 31578 -55746 31584 -55686
rect 31644 -55746 31650 -55686
rect 30040 -55860 30046 -55800
rect 30106 -55860 30112 -55800
rect 32076 -55860 32082 -55800
rect 32142 -55860 32148 -55800
rect 29324 -56004 29812 -55998
rect 29324 -56038 29336 -56004
rect 29800 -56038 29812 -56004
rect 29324 -56044 29812 -56038
rect 28058 -56664 28064 -56144
rect 28018 -56676 28064 -56664
rect 29028 -56664 29042 -56088
rect 29076 -56664 29088 -56088
rect 30046 -56088 30106 -55860
rect 31058 -55964 31064 -55904
rect 31124 -55964 31130 -55904
rect 30342 -56004 30830 -55998
rect 30342 -56038 30354 -56004
rect 30818 -56038 30830 -56004
rect 30342 -56044 30830 -56038
rect 30046 -56148 30060 -56088
rect 30054 -56628 30060 -56148
rect 28306 -56714 28794 -56708
rect 28306 -56748 28318 -56714
rect 28782 -56748 28794 -56714
rect 28306 -56754 28794 -56748
rect 27886 -56862 27892 -56802
rect 27952 -56862 27958 -56802
rect 27558 -56966 27564 -56906
rect 27624 -56966 27630 -56906
rect 27892 -57132 27952 -56862
rect 29028 -56906 29088 -56664
rect 30048 -56664 30060 -56628
rect 30094 -56148 30106 -56088
rect 31064 -56088 31124 -55964
rect 31360 -56004 31848 -55998
rect 31360 -56038 31372 -56004
rect 31836 -56038 31848 -56004
rect 31360 -56044 31848 -56038
rect 31064 -56142 31078 -56088
rect 30094 -56628 30100 -56148
rect 31072 -56624 31078 -56142
rect 30094 -56664 30108 -56628
rect 29324 -56714 29812 -56708
rect 29324 -56748 29336 -56714
rect 29800 -56748 29812 -56714
rect 29324 -56754 29812 -56748
rect 29022 -56966 29028 -56906
rect 29088 -56966 29094 -56906
rect 29536 -57012 29596 -56754
rect 29530 -57072 29536 -57012
rect 29596 -57072 29602 -57012
rect 27892 -57192 29092 -57132
rect 26508 -58026 26514 -57966
rect 26574 -58026 26580 -57966
rect 27892 -58044 27952 -57192
rect 28012 -57320 28072 -57192
rect 28498 -57230 28558 -57192
rect 28306 -57236 28794 -57230
rect 28306 -57270 28318 -57236
rect 28782 -57270 28794 -57236
rect 28306 -57276 28794 -57270
rect 28012 -57392 28024 -57320
rect 28018 -57896 28024 -57392
rect 28058 -57392 28072 -57320
rect 29032 -57320 29092 -57192
rect 29536 -57230 29596 -57072
rect 30048 -57122 30108 -56664
rect 31062 -56664 31078 -56624
rect 31112 -56142 31124 -56088
rect 32082 -56088 32142 -55860
rect 32584 -55998 32644 -55520
rect 33102 -55800 33162 -55430
rect 34126 -55430 34132 -54914
rect 34166 -54914 34174 -54854
rect 35134 -54854 35194 -54716
rect 35636 -54764 35696 -54500
rect 35982 -54536 36042 -54382
rect 35976 -54596 35982 -54536
rect 36042 -54596 36048 -54536
rect 36152 -54590 36158 -54530
rect 36218 -54590 36224 -54530
rect 35432 -54770 35920 -54764
rect 35432 -54804 35444 -54770
rect 35908 -54804 35920 -54770
rect 35432 -54810 35920 -54804
rect 35134 -54894 35150 -54854
rect 34166 -55430 34172 -54914
rect 35144 -55364 35150 -54894
rect 34126 -55442 34172 -55430
rect 35138 -55430 35150 -55364
rect 35184 -54894 35194 -54854
rect 36158 -54854 36218 -54590
rect 36674 -54592 36734 -54288
rect 37688 -54428 37748 -54288
rect 38194 -54322 38254 -54198
rect 39216 -54198 39222 -53660
rect 39256 -53660 39270 -53622
rect 40234 -53622 40280 -53610
rect 39256 -54198 39262 -53660
rect 40234 -54128 40240 -53622
rect 39216 -54210 39262 -54198
rect 40226 -54198 40240 -54128
rect 40274 -54128 40280 -53622
rect 41242 -53622 41302 -53268
rect 41600 -53414 41660 -53156
rect 41790 -53306 41850 -53054
rect 42766 -53306 42826 -53054
rect 41784 -53366 41790 -53306
rect 41850 -53366 41856 -53306
rect 42760 -53366 42766 -53306
rect 42826 -53366 42832 -53306
rect 43280 -53418 43340 -52964
rect 44306 -52964 44312 -52454
rect 44346 -52454 44356 -52388
rect 45324 -52388 45370 -52376
rect 44346 -52964 44352 -52454
rect 45324 -52920 45330 -52388
rect 44306 -52976 44352 -52964
rect 45318 -52964 45330 -52920
rect 45364 -52920 45370 -52388
rect 46334 -52388 46394 -52038
rect 46852 -52092 46912 -51820
rect 47354 -51912 47414 -51730
rect 48368 -51730 48384 -51696
rect 48418 -51696 48424 -51154
rect 48418 -51730 48428 -51696
rect 47648 -51780 48136 -51774
rect 47648 -51814 47660 -51780
rect 48124 -51814 48136 -51780
rect 47648 -51820 48136 -51814
rect 47862 -51912 47922 -51820
rect 48368 -51912 48428 -51730
rect 47354 -51972 48428 -51912
rect 46846 -52152 46852 -52092
rect 46912 -52152 46918 -52092
rect 47350 -52254 47356 -52194
rect 47416 -52254 47422 -52194
rect 46630 -52304 47118 -52298
rect 46630 -52338 46642 -52304
rect 47106 -52338 47118 -52304
rect 46630 -52344 47118 -52338
rect 46334 -52440 46348 -52388
rect 46342 -52914 46348 -52440
rect 45364 -52964 45378 -52920
rect 43576 -53014 44064 -53008
rect 43576 -53048 43588 -53014
rect 44052 -53048 44064 -53014
rect 43576 -53054 44064 -53048
rect 44594 -53014 45082 -53008
rect 44594 -53048 44606 -53014
rect 45070 -53048 45082 -53014
rect 44594 -53054 45082 -53048
rect 43782 -53306 43842 -53054
rect 45318 -53096 45378 -52964
rect 46336 -52964 46348 -52914
rect 46382 -52440 46394 -52388
rect 47356 -52388 47416 -52254
rect 47648 -52304 48136 -52298
rect 47648 -52338 47660 -52304
rect 48124 -52338 48136 -52304
rect 47648 -52344 48136 -52338
rect 47356 -52422 47366 -52388
rect 46382 -52914 46388 -52440
rect 46382 -52964 46396 -52914
rect 47360 -52920 47366 -52422
rect 45612 -53014 46100 -53008
rect 45612 -53048 45624 -53014
rect 46088 -53048 46100 -53014
rect 45612 -53054 46100 -53048
rect 45312 -53156 45318 -53096
rect 45378 -53156 45384 -53096
rect 43776 -53366 43782 -53306
rect 43842 -53366 43848 -53306
rect 45802 -53366 45808 -53306
rect 45868 -53366 45874 -53306
rect 41600 -53480 41660 -53474
rect 43274 -53478 43280 -53418
rect 43340 -53478 43346 -53418
rect 45310 -53478 45316 -53418
rect 45376 -53478 45382 -53418
rect 41540 -53538 42028 -53532
rect 41540 -53572 41552 -53538
rect 42016 -53572 42028 -53538
rect 41540 -53578 42028 -53572
rect 42558 -53538 43046 -53532
rect 42558 -53572 42570 -53538
rect 43034 -53572 43046 -53538
rect 42558 -53578 43046 -53572
rect 41242 -53664 41258 -53622
rect 40274 -54198 40286 -54128
rect 38486 -54248 38974 -54242
rect 38486 -54282 38498 -54248
rect 38962 -54282 38974 -54248
rect 38486 -54288 38974 -54282
rect 39504 -54248 39992 -54242
rect 39504 -54282 39516 -54248
rect 39980 -54282 39992 -54248
rect 39504 -54288 39992 -54282
rect 38188 -54382 38194 -54322
rect 38254 -54382 38260 -54322
rect 38710 -54428 38770 -54288
rect 39724 -54428 39784 -54288
rect 40226 -54322 40286 -54198
rect 41252 -54198 41258 -53664
rect 41292 -53664 41302 -53622
rect 42270 -53622 42316 -53610
rect 41292 -54198 41298 -53664
rect 42270 -54162 42276 -53622
rect 41252 -54210 41298 -54198
rect 42266 -54198 42276 -54162
rect 42310 -54162 42316 -53622
rect 43280 -53622 43340 -53478
rect 43576 -53538 44064 -53532
rect 43576 -53572 43588 -53538
rect 44052 -53572 44064 -53538
rect 43576 -53578 44064 -53572
rect 44594 -53538 45082 -53532
rect 44594 -53572 44606 -53538
rect 45070 -53572 45082 -53538
rect 44594 -53578 45082 -53572
rect 43280 -53660 43294 -53622
rect 43288 -54146 43294 -53660
rect 42310 -54198 42326 -54162
rect 40522 -54248 41010 -54242
rect 40522 -54282 40534 -54248
rect 40998 -54282 41010 -54248
rect 40522 -54288 41010 -54282
rect 41540 -54248 42028 -54242
rect 41540 -54282 41552 -54248
rect 42016 -54282 42028 -54248
rect 41540 -54288 42028 -54282
rect 40220 -54382 40226 -54322
rect 40286 -54382 40292 -54322
rect 40726 -54328 40786 -54288
rect 41752 -54328 41812 -54288
rect 42266 -54322 42326 -54198
rect 43284 -54198 43294 -54146
rect 43328 -53660 43340 -53622
rect 44306 -53622 44352 -53610
rect 43328 -54146 43334 -53660
rect 43328 -54198 43344 -54146
rect 44306 -54154 44312 -53622
rect 42558 -54248 43046 -54242
rect 42558 -54282 42570 -54248
rect 43034 -54282 43046 -54248
rect 42558 -54288 43046 -54282
rect 40726 -54388 41812 -54328
rect 42260 -54382 42266 -54322
rect 42326 -54382 42332 -54322
rect 40726 -54428 40786 -54388
rect 37688 -54488 40786 -54428
rect 41238 -54480 41244 -54420
rect 41304 -54480 41310 -54420
rect 37688 -54592 37748 -54488
rect 38180 -54590 38186 -54530
rect 38246 -54590 38252 -54530
rect 36674 -54652 37748 -54592
rect 36674 -54764 36734 -54652
rect 37688 -54764 37748 -54652
rect 36450 -54770 36938 -54764
rect 36450 -54804 36462 -54770
rect 36926 -54804 36938 -54770
rect 36450 -54810 36938 -54804
rect 37468 -54770 37956 -54764
rect 37468 -54804 37480 -54770
rect 37944 -54804 37956 -54770
rect 37468 -54810 37956 -54804
rect 35184 -55364 35190 -54894
rect 36158 -54898 36168 -54854
rect 35184 -55430 35198 -55364
rect 36162 -55372 36168 -54898
rect 33396 -55480 33884 -55474
rect 33396 -55514 33408 -55480
rect 33872 -55514 33884 -55480
rect 33396 -55520 33884 -55514
rect 34414 -55480 34902 -55474
rect 34414 -55514 34426 -55480
rect 34890 -55514 34902 -55480
rect 34414 -55520 34902 -55514
rect 33096 -55860 33102 -55800
rect 33162 -55860 33168 -55800
rect 33606 -55998 33666 -55520
rect 34112 -55860 34118 -55800
rect 34178 -55860 34184 -55800
rect 32378 -56004 32866 -55998
rect 32378 -56038 32390 -56004
rect 32854 -56038 32866 -56004
rect 32378 -56044 32866 -56038
rect 33396 -56004 33884 -55998
rect 33396 -56038 33408 -56004
rect 33872 -56038 33884 -56004
rect 33396 -56044 33884 -56038
rect 32082 -56138 32096 -56088
rect 31112 -56624 31118 -56142
rect 31112 -56664 31122 -56624
rect 32090 -56640 32096 -56138
rect 30342 -56714 30830 -56708
rect 30342 -56748 30354 -56714
rect 30818 -56748 30830 -56714
rect 30342 -56754 30830 -56748
rect 30556 -57012 30616 -56754
rect 31062 -56802 31122 -56664
rect 32084 -56664 32096 -56640
rect 32130 -56138 32142 -56088
rect 33108 -56088 33154 -56076
rect 32130 -56640 32136 -56138
rect 32130 -56664 32144 -56640
rect 33108 -56650 33114 -56088
rect 31360 -56714 31848 -56708
rect 31360 -56748 31372 -56714
rect 31836 -56748 31848 -56714
rect 31360 -56754 31848 -56748
rect 31056 -56862 31062 -56802
rect 31122 -56862 31128 -56802
rect 31062 -56966 31068 -56906
rect 31128 -56966 31134 -56906
rect 30550 -57072 30556 -57012
rect 30616 -57072 30622 -57012
rect 30042 -57182 30048 -57122
rect 30108 -57182 30114 -57122
rect 29324 -57236 29812 -57230
rect 29324 -57270 29336 -57236
rect 29800 -57270 29812 -57236
rect 29324 -57276 29812 -57270
rect 28058 -57896 28064 -57392
rect 29032 -57396 29042 -57320
rect 29036 -57848 29042 -57396
rect 28018 -57908 28064 -57896
rect 29028 -57896 29042 -57848
rect 29076 -57396 29092 -57320
rect 30048 -57320 30108 -57182
rect 30556 -57230 30616 -57072
rect 30342 -57236 30830 -57230
rect 30342 -57270 30354 -57236
rect 30818 -57270 30830 -57236
rect 30342 -57276 30830 -57270
rect 29076 -57848 29082 -57396
rect 29076 -57896 29088 -57848
rect 28306 -57946 28794 -57940
rect 28306 -57980 28318 -57946
rect 28782 -57980 28794 -57946
rect 28306 -57986 28794 -57980
rect 29028 -58044 29088 -57896
rect 30048 -57896 30060 -57320
rect 30094 -57896 30108 -57320
rect 31068 -57320 31128 -56966
rect 31580 -57012 31640 -56754
rect 31574 -57072 31580 -57012
rect 31640 -57072 31646 -57012
rect 31580 -57230 31640 -57072
rect 32084 -57122 32144 -56664
rect 33098 -56664 33114 -56650
rect 33148 -56650 33154 -56088
rect 34118 -56088 34178 -55860
rect 34618 -55998 34678 -55520
rect 35138 -55800 35198 -55430
rect 36150 -55430 36168 -55372
rect 36202 -54898 36218 -54854
rect 37180 -54854 37226 -54842
rect 36202 -55372 36208 -54898
rect 36202 -55430 36210 -55372
rect 37180 -55378 37186 -54854
rect 35432 -55480 35920 -55474
rect 35432 -55514 35444 -55480
rect 35908 -55514 35920 -55480
rect 35432 -55520 35920 -55514
rect 35132 -55860 35138 -55800
rect 35198 -55860 35204 -55800
rect 35648 -55998 35708 -55520
rect 36150 -55632 36210 -55430
rect 37168 -55430 37186 -55378
rect 37220 -55378 37226 -54854
rect 38186 -54854 38246 -54590
rect 38710 -54764 38770 -54488
rect 39724 -54764 39784 -54488
rect 40224 -54590 40230 -54530
rect 40290 -54590 40296 -54530
rect 38486 -54770 38974 -54764
rect 38486 -54804 38498 -54770
rect 38962 -54804 38974 -54770
rect 38486 -54810 38974 -54804
rect 39504 -54770 39992 -54764
rect 39504 -54804 39516 -54770
rect 39980 -54804 39992 -54770
rect 39504 -54810 39992 -54804
rect 38186 -54898 38204 -54854
rect 37220 -55430 37228 -55378
rect 36450 -55480 36938 -55474
rect 36450 -55514 36462 -55480
rect 36926 -55514 36938 -55480
rect 36450 -55520 36938 -55514
rect 36000 -55692 36210 -55632
rect 36664 -55686 36724 -55520
rect 37168 -55572 37228 -55430
rect 38198 -55430 38204 -54898
rect 38238 -54898 38246 -54854
rect 39216 -54854 39262 -54842
rect 38238 -55430 38244 -54898
rect 39216 -55378 39222 -54854
rect 38198 -55442 38244 -55430
rect 39210 -55430 39222 -55378
rect 39256 -55378 39262 -54854
rect 40230 -54854 40290 -54590
rect 40726 -54764 40786 -54488
rect 40522 -54770 41010 -54764
rect 40522 -54804 40534 -54770
rect 40998 -54804 41010 -54770
rect 40522 -54810 41010 -54804
rect 40230 -54902 40240 -54854
rect 39256 -55430 39270 -55378
rect 37468 -55480 37956 -55474
rect 37468 -55514 37480 -55480
rect 37944 -55514 37956 -55480
rect 37468 -55520 37956 -55514
rect 38486 -55480 38974 -55474
rect 38486 -55514 38498 -55480
rect 38962 -55514 38974 -55480
rect 38486 -55520 38974 -55514
rect 39210 -55572 39270 -55430
rect 40234 -55430 40240 -54902
rect 40274 -54902 40290 -54854
rect 41244 -54854 41304 -54480
rect 41752 -54764 41812 -54388
rect 42252 -54590 42258 -54530
rect 42318 -54590 42324 -54530
rect 41540 -54770 42028 -54764
rect 41540 -54804 41552 -54770
rect 42016 -54804 42028 -54770
rect 41540 -54810 42028 -54804
rect 41244 -54890 41258 -54854
rect 40274 -55430 40280 -54902
rect 41252 -55386 41258 -54890
rect 40234 -55442 40280 -55430
rect 41246 -55430 41258 -55386
rect 41292 -54890 41304 -54854
rect 42258 -54854 42318 -54590
rect 42772 -54764 42832 -54288
rect 43284 -54656 43344 -54198
rect 44296 -54198 44312 -54154
rect 44346 -54154 44352 -53622
rect 45316 -53622 45376 -53478
rect 45808 -53532 45868 -53366
rect 45612 -53538 46100 -53532
rect 45612 -53572 45624 -53538
rect 46088 -53572 46100 -53538
rect 45612 -53578 46100 -53572
rect 45316 -53680 45330 -53622
rect 44346 -54198 44356 -54154
rect 45324 -54158 45330 -53680
rect 43576 -54248 44064 -54242
rect 43576 -54282 43588 -54248
rect 44052 -54282 44064 -54248
rect 43576 -54288 44064 -54282
rect 43278 -54716 43284 -54656
rect 43344 -54716 43350 -54656
rect 42558 -54770 43046 -54764
rect 42558 -54804 42570 -54770
rect 43034 -54804 43046 -54770
rect 42558 -54810 43046 -54804
rect 41292 -55386 41298 -54890
rect 42258 -54902 42276 -54854
rect 41292 -55430 41306 -55386
rect 42270 -55390 42276 -54902
rect 39504 -55480 39992 -55474
rect 39504 -55514 39516 -55480
rect 39980 -55514 39992 -55480
rect 39504 -55520 39992 -55514
rect 40522 -55480 41010 -55474
rect 40522 -55514 40534 -55480
rect 40998 -55514 41010 -55480
rect 40522 -55520 41010 -55514
rect 41246 -55572 41306 -55430
rect 42260 -55430 42276 -55390
rect 42310 -54902 42318 -54854
rect 43284 -54854 43344 -54716
rect 43788 -54764 43848 -54288
rect 44296 -54530 44356 -54198
rect 45314 -54198 45330 -54158
rect 45364 -53680 45376 -53622
rect 46336 -53622 46396 -52964
rect 47352 -52964 47366 -52920
rect 47400 -52422 47416 -52388
rect 48378 -52388 48424 -52376
rect 47400 -52920 47406 -52422
rect 47400 -52964 47412 -52920
rect 48378 -52934 48384 -52388
rect 46630 -53014 47118 -53008
rect 46630 -53048 46642 -53014
rect 47106 -53048 47118 -53014
rect 46630 -53054 47118 -53048
rect 46838 -53306 46898 -53054
rect 47352 -53146 47412 -52964
rect 48368 -52964 48384 -52934
rect 48418 -52934 48424 -52388
rect 48418 -52964 48428 -52934
rect 47648 -53014 48136 -53008
rect 47648 -53048 47660 -53014
rect 48124 -53048 48136 -53014
rect 47648 -53054 48136 -53048
rect 47858 -53146 47918 -53054
rect 48368 -53146 48428 -52964
rect 47352 -53206 48428 -53146
rect 46832 -53366 46838 -53306
rect 46898 -53366 46904 -53306
rect 47352 -53418 47412 -53206
rect 47346 -53478 47352 -53418
rect 47412 -53478 47418 -53418
rect 46630 -53538 47118 -53532
rect 46630 -53572 46642 -53538
rect 47106 -53572 47118 -53538
rect 46630 -53578 47118 -53572
rect 47648 -53538 48136 -53532
rect 47648 -53572 47660 -53538
rect 48124 -53572 48136 -53538
rect 47648 -53578 48136 -53572
rect 46336 -53664 46348 -53622
rect 45364 -54158 45370 -53680
rect 46342 -54144 46348 -53664
rect 45364 -54198 45374 -54158
rect 44594 -54248 45082 -54242
rect 44594 -54282 44606 -54248
rect 45070 -54282 45082 -54248
rect 44594 -54288 45082 -54282
rect 44290 -54590 44296 -54530
rect 44356 -54590 44362 -54530
rect 44822 -54764 44882 -54288
rect 45314 -54656 45374 -54198
rect 46336 -54198 46348 -54144
rect 46382 -53664 46396 -53622
rect 47360 -53622 47406 -53610
rect 46382 -54144 46388 -53664
rect 46382 -54198 46396 -54144
rect 47360 -54152 47366 -53622
rect 45612 -54248 46100 -54242
rect 45612 -54282 45624 -54248
rect 46088 -54282 46100 -54248
rect 45612 -54288 46100 -54282
rect 45840 -54654 45900 -54288
rect 46336 -54530 46396 -54198
rect 47350 -54198 47366 -54152
rect 47400 -54152 47406 -53622
rect 48378 -53622 48424 -53610
rect 47400 -54198 47410 -54152
rect 48378 -54170 48384 -53622
rect 46630 -54248 47118 -54242
rect 46630 -54282 46642 -54248
rect 47106 -54282 47118 -54248
rect 46630 -54288 47118 -54282
rect 46854 -54526 46914 -54288
rect 47350 -54324 47410 -54198
rect 48370 -54198 48384 -54170
rect 48418 -54170 48424 -53622
rect 48418 -54198 48430 -54170
rect 47648 -54248 48136 -54242
rect 47648 -54282 47660 -54248
rect 48124 -54282 48136 -54248
rect 47648 -54288 48136 -54282
rect 47856 -54322 47916 -54288
rect 48370 -54322 48430 -54198
rect 47856 -54324 48430 -54322
rect 47350 -54384 48430 -54324
rect 47350 -54420 47410 -54384
rect 47344 -54480 47350 -54420
rect 47410 -54480 47416 -54420
rect 46330 -54590 46336 -54530
rect 46396 -54590 46402 -54530
rect 46848 -54586 46854 -54526
rect 46914 -54586 46920 -54526
rect 48360 -54586 48366 -54526
rect 48426 -54586 48432 -54526
rect 45308 -54716 45314 -54656
rect 45374 -54716 45380 -54656
rect 43576 -54770 44064 -54764
rect 43576 -54804 43588 -54770
rect 44052 -54804 44064 -54770
rect 43576 -54810 44064 -54804
rect 44594 -54770 45082 -54764
rect 44594 -54804 44606 -54770
rect 45070 -54804 45082 -54770
rect 44594 -54810 45082 -54804
rect 43284 -54900 43294 -54854
rect 42310 -55390 42316 -54902
rect 43288 -55370 43294 -54900
rect 42310 -55430 42320 -55390
rect 41540 -55480 42028 -55474
rect 41540 -55514 41552 -55480
rect 42016 -55514 42028 -55480
rect 41540 -55520 42028 -55514
rect 37162 -55632 37168 -55572
rect 37228 -55632 37234 -55572
rect 39204 -55632 39210 -55572
rect 39270 -55632 39276 -55572
rect 41240 -55632 41246 -55572
rect 41306 -55632 41312 -55572
rect 41752 -55682 41812 -55520
rect 42260 -55580 42320 -55430
rect 43282 -55430 43294 -55370
rect 43328 -54900 43344 -54854
rect 44306 -54854 44352 -54842
rect 43328 -55370 43334 -54900
rect 43328 -55430 43342 -55370
rect 44306 -55386 44312 -54854
rect 42558 -55480 43046 -55474
rect 42558 -55514 42570 -55480
rect 43034 -55514 43046 -55480
rect 42558 -55520 43046 -55514
rect 42260 -55640 42466 -55580
rect 36000 -55904 36060 -55692
rect 36658 -55746 36664 -55686
rect 36724 -55746 36730 -55686
rect 41746 -55742 41752 -55682
rect 41812 -55742 41818 -55682
rect 36150 -55860 36156 -55800
rect 36216 -55860 36222 -55800
rect 38180 -55860 38186 -55800
rect 38246 -55860 38252 -55800
rect 40218 -55860 40224 -55800
rect 40284 -55860 40290 -55800
rect 42254 -55860 42260 -55800
rect 42320 -55860 42326 -55800
rect 35994 -55964 36000 -55904
rect 36060 -55964 36066 -55904
rect 34414 -56004 34902 -55998
rect 34414 -56038 34426 -56004
rect 34890 -56038 34902 -56004
rect 34414 -56044 34902 -56038
rect 35432 -56004 35920 -55998
rect 35432 -56038 35444 -56004
rect 35908 -56038 35920 -56004
rect 35432 -56044 35920 -56038
rect 34118 -56570 34132 -56088
rect 34126 -56644 34132 -56570
rect 33148 -56664 33158 -56650
rect 32378 -56714 32866 -56708
rect 32378 -56748 32390 -56714
rect 32854 -56748 32866 -56714
rect 32378 -56754 32866 -56748
rect 32598 -57012 32658 -56754
rect 33098 -56906 33158 -56664
rect 34122 -56664 34132 -56644
rect 34166 -56570 34178 -56088
rect 35144 -56088 35190 -56076
rect 34166 -56644 34172 -56570
rect 35144 -56638 35150 -56088
rect 34166 -56664 34182 -56644
rect 33396 -56714 33884 -56708
rect 33396 -56748 33408 -56714
rect 33872 -56748 33884 -56714
rect 33396 -56754 33884 -56748
rect 33092 -56966 33098 -56906
rect 33158 -56966 33164 -56906
rect 33612 -57012 33672 -56754
rect 32592 -57072 32598 -57012
rect 32658 -57072 32664 -57012
rect 33606 -57072 33612 -57012
rect 33672 -57072 33678 -57012
rect 32078 -57182 32084 -57122
rect 32144 -57182 32150 -57122
rect 31360 -57236 31848 -57230
rect 31360 -57270 31372 -57236
rect 31836 -57270 31848 -57236
rect 31360 -57276 31848 -57270
rect 31068 -57334 31078 -57320
rect 29324 -57946 29812 -57940
rect 29324 -57980 29336 -57946
rect 29800 -57980 29812 -57946
rect 29324 -57986 29812 -57980
rect 27886 -58104 27892 -58044
rect 27952 -58104 27958 -58044
rect 29022 -58104 29028 -58044
rect 29088 -58104 29094 -58044
rect 29540 -58152 29600 -57986
rect 29534 -58212 29540 -58152
rect 29600 -58212 29606 -58152
rect 30048 -58408 30108 -57896
rect 31072 -57896 31078 -57334
rect 31112 -57334 31128 -57320
rect 32084 -57320 32144 -57182
rect 32598 -57230 32658 -57072
rect 33612 -57230 33672 -57072
rect 34122 -57122 34182 -56664
rect 35138 -56664 35150 -56638
rect 35184 -56638 35190 -56088
rect 36156 -56088 36216 -55860
rect 36450 -56004 36938 -55998
rect 36450 -56038 36462 -56004
rect 36926 -56038 36938 -56004
rect 36450 -56044 36938 -56038
rect 37468 -56004 37956 -55998
rect 37468 -56038 37480 -56004
rect 37944 -56038 37956 -56004
rect 37468 -56044 37956 -56038
rect 37180 -56088 37226 -56076
rect 38186 -56088 38246 -55860
rect 38486 -56004 38974 -55998
rect 38486 -56038 38498 -56004
rect 38962 -56038 38974 -56004
rect 38486 -56044 38974 -56038
rect 39504 -56004 39992 -55998
rect 39504 -56038 39516 -56004
rect 39980 -56038 39992 -56004
rect 39504 -56044 39992 -56038
rect 39216 -56088 39262 -56076
rect 40224 -56088 40284 -55860
rect 40522 -56004 41010 -55998
rect 40522 -56038 40534 -56004
rect 40998 -56038 41010 -56004
rect 40522 -56044 41010 -56038
rect 41540 -56004 42028 -55998
rect 41540 -56038 41552 -56004
rect 42016 -56038 42028 -56004
rect 41540 -56044 42028 -56038
rect 36156 -56144 36168 -56088
rect 35184 -56664 35198 -56638
rect 36162 -56640 36168 -56144
rect 34414 -56714 34902 -56708
rect 34414 -56748 34426 -56714
rect 34890 -56748 34902 -56714
rect 34414 -56754 34902 -56748
rect 34644 -57012 34704 -56754
rect 35138 -56906 35198 -56664
rect 36160 -56664 36168 -56640
rect 36202 -56144 36216 -56088
rect 37174 -56124 37186 -56088
rect 36202 -56640 36208 -56144
rect 37180 -56612 37186 -56124
rect 36202 -56664 36220 -56640
rect 35432 -56714 35920 -56708
rect 35432 -56748 35444 -56714
rect 35908 -56748 35920 -56714
rect 35432 -56754 35920 -56748
rect 35286 -56860 35292 -56800
rect 35352 -56860 35358 -56800
rect 35132 -56966 35138 -56906
rect 35198 -56966 35204 -56906
rect 34638 -57072 34644 -57012
rect 34704 -57072 34710 -57012
rect 35292 -57044 35352 -56860
rect 35656 -57012 35716 -56754
rect 34116 -57182 34122 -57122
rect 34182 -57182 34188 -57122
rect 32378 -57236 32866 -57230
rect 32378 -57270 32390 -57236
rect 32854 -57270 32866 -57236
rect 32378 -57276 32866 -57270
rect 33396 -57236 33884 -57230
rect 33396 -57270 33408 -57236
rect 33872 -57270 33884 -57236
rect 33396 -57276 33884 -57270
rect 31112 -57896 31118 -57334
rect 31072 -57908 31118 -57896
rect 32084 -57896 32096 -57320
rect 32130 -57896 32144 -57320
rect 33108 -57320 33154 -57308
rect 33108 -57854 33114 -57320
rect 30342 -57946 30830 -57940
rect 30342 -57980 30354 -57946
rect 30818 -57980 30830 -57946
rect 30342 -57986 30830 -57980
rect 31360 -57946 31848 -57940
rect 31360 -57980 31372 -57946
rect 31836 -57980 31848 -57946
rect 31360 -57986 31848 -57980
rect 30554 -58152 30614 -57986
rect 30554 -58218 30614 -58212
rect 31576 -58152 31636 -57986
rect 31576 -58218 31636 -58212
rect 32084 -58408 32144 -57896
rect 33098 -57896 33114 -57854
rect 33148 -57854 33154 -57320
rect 34122 -57320 34182 -57182
rect 34644 -57230 34704 -57072
rect 35136 -57104 35352 -57044
rect 35650 -57072 35656 -57012
rect 35716 -57072 35722 -57012
rect 34414 -57236 34902 -57230
rect 34414 -57270 34426 -57236
rect 34890 -57270 34902 -57236
rect 34414 -57276 34902 -57270
rect 33148 -57896 33158 -57854
rect 32378 -57946 32866 -57940
rect 32378 -57980 32390 -57946
rect 32854 -57980 32866 -57946
rect 32378 -57986 32866 -57980
rect 32588 -58146 32648 -57986
rect 33098 -58044 33158 -57896
rect 34122 -57896 34132 -57320
rect 34166 -57896 34182 -57320
rect 35136 -57320 35196 -57104
rect 35656 -57230 35716 -57072
rect 36160 -57122 36220 -56664
rect 37170 -56664 37186 -56612
rect 37220 -56124 37234 -56088
rect 37220 -56612 37226 -56124
rect 38186 -56138 38204 -56088
rect 37220 -56664 37230 -56612
rect 38198 -56634 38204 -56138
rect 36450 -56714 36938 -56708
rect 36450 -56748 36462 -56714
rect 36926 -56748 36938 -56714
rect 36450 -56754 36938 -56748
rect 36664 -57012 36724 -56754
rect 37170 -56800 37230 -56664
rect 38196 -56664 38204 -56634
rect 38238 -56138 38246 -56088
rect 39210 -56120 39222 -56088
rect 38238 -56634 38244 -56138
rect 39216 -56624 39222 -56120
rect 38238 -56664 38256 -56634
rect 37468 -56714 37956 -56708
rect 37468 -56748 37480 -56714
rect 37944 -56748 37956 -56714
rect 37468 -56754 37956 -56748
rect 37164 -56860 37170 -56800
rect 37230 -56860 37236 -56800
rect 37168 -56966 37174 -56906
rect 37234 -56966 37240 -56906
rect 36658 -57072 36664 -57012
rect 36724 -57072 36730 -57012
rect 36154 -57182 36160 -57122
rect 36220 -57182 36226 -57122
rect 35432 -57236 35920 -57230
rect 35432 -57270 35444 -57236
rect 35908 -57270 35920 -57236
rect 35432 -57276 35920 -57270
rect 35136 -57346 35150 -57320
rect 33396 -57946 33884 -57940
rect 33396 -57980 33408 -57946
rect 33872 -57980 33884 -57946
rect 33396 -57986 33884 -57980
rect 33092 -58104 33098 -58044
rect 33158 -58104 33164 -58044
rect 33614 -58146 33674 -57986
rect 32588 -58152 32650 -58146
rect 32588 -58158 32590 -58152
rect 33614 -58152 33676 -58146
rect 33614 -58158 33616 -58152
rect 32590 -58218 32650 -58212
rect 33616 -58218 33676 -58212
rect 34122 -58408 34182 -57896
rect 35144 -57896 35150 -57346
rect 35184 -57346 35196 -57320
rect 36160 -57320 36220 -57182
rect 36664 -57230 36724 -57072
rect 36450 -57236 36938 -57230
rect 36450 -57270 36462 -57236
rect 36926 -57270 36938 -57236
rect 36450 -57276 36938 -57270
rect 35184 -57896 35190 -57346
rect 35144 -57908 35190 -57896
rect 36160 -57896 36168 -57320
rect 36202 -57896 36220 -57320
rect 37174 -57320 37234 -56966
rect 37682 -57012 37742 -56754
rect 37676 -57072 37682 -57012
rect 37742 -57072 37748 -57012
rect 37682 -57230 37742 -57072
rect 38196 -57122 38256 -56664
rect 39208 -56664 39222 -56624
rect 39256 -56120 39270 -56088
rect 39256 -56624 39262 -56120
rect 40224 -56132 40240 -56088
rect 39256 -56664 39268 -56624
rect 40234 -56640 40240 -56132
rect 38486 -56714 38974 -56708
rect 38486 -56748 38498 -56714
rect 38962 -56748 38974 -56714
rect 38486 -56754 38974 -56748
rect 38708 -57012 38768 -56754
rect 39208 -56800 39268 -56664
rect 40232 -56664 40240 -56640
rect 40274 -56132 40284 -56088
rect 41252 -56088 41298 -56076
rect 40274 -56640 40280 -56132
rect 41252 -56618 41258 -56088
rect 40274 -56664 40292 -56640
rect 39504 -56714 39992 -56708
rect 39504 -56748 39516 -56714
rect 39980 -56748 39992 -56714
rect 39504 -56754 39992 -56748
rect 39202 -56860 39208 -56800
rect 39268 -56860 39274 -56800
rect 39204 -56966 39210 -56906
rect 39270 -56966 39276 -56906
rect 38702 -57072 38708 -57012
rect 38768 -57072 38774 -57012
rect 38190 -57182 38196 -57122
rect 38256 -57182 38262 -57122
rect 37468 -57236 37956 -57230
rect 37468 -57270 37480 -57236
rect 37944 -57270 37956 -57236
rect 37468 -57276 37956 -57270
rect 37174 -57346 37186 -57320
rect 34414 -57946 34902 -57940
rect 34414 -57980 34426 -57946
rect 34890 -57980 34902 -57946
rect 34414 -57986 34902 -57980
rect 35432 -57946 35920 -57940
rect 35432 -57980 35444 -57946
rect 35908 -57980 35920 -57946
rect 35432 -57986 35920 -57980
rect 34628 -58152 34688 -57986
rect 34628 -58218 34688 -58212
rect 35664 -58152 35724 -57986
rect 35664 -58218 35724 -58212
rect 36160 -58408 36220 -57896
rect 37180 -57896 37186 -57346
rect 37220 -57346 37234 -57320
rect 38196 -57320 38256 -57182
rect 38708 -57230 38768 -57072
rect 38486 -57236 38974 -57230
rect 38486 -57270 38498 -57236
rect 38962 -57270 38974 -57236
rect 38486 -57276 38974 -57270
rect 37220 -57896 37226 -57346
rect 37180 -57908 37226 -57896
rect 38196 -57896 38204 -57320
rect 38238 -57896 38256 -57320
rect 39210 -57320 39270 -56966
rect 39710 -57012 39770 -56754
rect 39704 -57072 39710 -57012
rect 39770 -57072 39776 -57012
rect 39710 -57230 39770 -57072
rect 40232 -57122 40292 -56664
rect 41244 -56664 41258 -56618
rect 41292 -56618 41298 -56088
rect 42260 -56088 42320 -55860
rect 42406 -55904 42466 -55640
rect 42400 -55964 42406 -55904
rect 42466 -55964 42472 -55904
rect 42770 -55998 42830 -55520
rect 43282 -55800 43342 -55430
rect 44300 -55430 44312 -55386
rect 44346 -55386 44352 -54854
rect 45314 -54854 45374 -54716
rect 45840 -54764 45900 -54714
rect 46854 -54764 46914 -54586
rect 47348 -54714 47354 -54654
rect 47414 -54714 47420 -54654
rect 45612 -54770 46100 -54764
rect 45612 -54804 45624 -54770
rect 46088 -54804 46100 -54770
rect 45612 -54810 46100 -54804
rect 46630 -54770 47118 -54764
rect 46630 -54804 46642 -54770
rect 47106 -54804 47118 -54770
rect 46630 -54810 47118 -54804
rect 45314 -54900 45330 -54854
rect 45324 -55382 45330 -54900
rect 44346 -55430 44360 -55386
rect 43576 -55480 44064 -55474
rect 43576 -55514 43588 -55480
rect 44052 -55514 44064 -55480
rect 43576 -55520 44064 -55514
rect 43276 -55860 43282 -55800
rect 43342 -55860 43348 -55800
rect 43790 -55998 43850 -55520
rect 44300 -55572 44360 -55430
rect 45316 -55430 45330 -55382
rect 45364 -54900 45374 -54854
rect 46342 -54854 46388 -54842
rect 47354 -54854 47414 -54714
rect 47648 -54770 48136 -54764
rect 47648 -54804 47660 -54770
rect 48124 -54804 48136 -54770
rect 47648 -54810 48136 -54804
rect 45364 -55382 45370 -54900
rect 45364 -55430 45376 -55382
rect 46342 -55386 46348 -54854
rect 44594 -55480 45082 -55474
rect 44594 -55514 44606 -55480
rect 45070 -55514 45082 -55480
rect 44594 -55520 45082 -55514
rect 44294 -55632 44300 -55572
rect 44360 -55632 44366 -55572
rect 44296 -55860 44302 -55800
rect 44362 -55860 44368 -55800
rect 42558 -56004 43046 -55998
rect 42558 -56038 42570 -56004
rect 43034 -56038 43046 -56004
rect 42558 -56044 43046 -56038
rect 43576 -56004 44064 -55998
rect 43576 -56038 43588 -56004
rect 44052 -56038 44064 -56004
rect 43576 -56044 44064 -56038
rect 42260 -56132 42276 -56088
rect 41292 -56664 41304 -56618
rect 42270 -56638 42276 -56132
rect 40522 -56714 41010 -56708
rect 40522 -56748 40534 -56714
rect 40998 -56748 41010 -56714
rect 40522 -56754 41010 -56748
rect 40730 -57012 40790 -56754
rect 41072 -56860 41078 -56800
rect 41138 -56860 41144 -56800
rect 40724 -57072 40730 -57012
rect 40790 -57072 40796 -57012
rect 41078 -57052 41138 -56860
rect 41244 -56906 41304 -56664
rect 42264 -56664 42276 -56638
rect 42310 -56132 42320 -56088
rect 43288 -56088 43334 -56076
rect 42310 -56638 42316 -56132
rect 43288 -56624 43294 -56088
rect 42310 -56664 42324 -56638
rect 41540 -56714 42028 -56708
rect 41540 -56748 41552 -56714
rect 42016 -56748 42028 -56714
rect 41540 -56754 42028 -56748
rect 41238 -56966 41244 -56906
rect 41304 -56966 41310 -56906
rect 41750 -57012 41810 -56754
rect 40226 -57182 40232 -57122
rect 40292 -57182 40298 -57122
rect 39504 -57236 39992 -57230
rect 39504 -57270 39516 -57236
rect 39980 -57270 39992 -57236
rect 39504 -57276 39992 -57270
rect 39210 -57356 39222 -57320
rect 36450 -57946 36938 -57940
rect 36450 -57980 36462 -57946
rect 36926 -57980 36938 -57946
rect 36450 -57986 36938 -57980
rect 37468 -57946 37956 -57940
rect 37468 -57980 37480 -57946
rect 37944 -57980 37956 -57946
rect 37468 -57986 37956 -57980
rect 36670 -58152 36730 -57986
rect 37684 -58152 37744 -57986
rect 37678 -58212 37684 -58152
rect 37744 -58212 37750 -58152
rect 36670 -58218 36730 -58212
rect 38196 -58408 38256 -57896
rect 39216 -57896 39222 -57356
rect 39256 -57356 39270 -57320
rect 40232 -57320 40292 -57182
rect 40730 -57230 40790 -57072
rect 41078 -57112 41304 -57052
rect 41744 -57072 41750 -57012
rect 41810 -57072 41816 -57012
rect 40522 -57236 41010 -57230
rect 40522 -57270 40534 -57236
rect 40998 -57270 41010 -57236
rect 40522 -57276 41010 -57270
rect 39256 -57896 39262 -57356
rect 39216 -57908 39262 -57896
rect 40232 -57896 40240 -57320
rect 40274 -57896 40292 -57320
rect 41244 -57320 41304 -57112
rect 41750 -57230 41810 -57072
rect 42264 -57122 42324 -56664
rect 43284 -56664 43294 -56624
rect 43328 -56624 43334 -56088
rect 44302 -56088 44362 -55860
rect 44804 -55998 44864 -55520
rect 45316 -55800 45376 -55430
rect 46332 -55430 46348 -55386
rect 46382 -55386 46388 -54854
rect 47352 -54888 47366 -54854
rect 47354 -54898 47366 -54888
rect 46382 -55430 46392 -55386
rect 45612 -55480 46100 -55474
rect 45612 -55514 45624 -55480
rect 46088 -55514 46100 -55480
rect 45612 -55520 46100 -55514
rect 45310 -55860 45316 -55800
rect 45376 -55860 45382 -55800
rect 45310 -55964 45316 -55904
rect 45376 -55964 45382 -55904
rect 44594 -56004 45082 -55998
rect 44594 -56038 44606 -56004
rect 45070 -56038 45082 -56004
rect 44594 -56044 45082 -56038
rect 44812 -56048 44872 -56044
rect 44302 -56154 44312 -56088
rect 44306 -56618 44312 -56154
rect 43328 -56664 43344 -56624
rect 42558 -56714 43046 -56708
rect 42558 -56748 42570 -56714
rect 43034 -56748 43046 -56714
rect 42558 -56754 43046 -56748
rect 42776 -57012 42836 -56754
rect 43284 -56906 43344 -56664
rect 44296 -56664 44312 -56618
rect 44346 -56154 44362 -56088
rect 45316 -56088 45376 -55964
rect 45840 -55998 45900 -55520
rect 46332 -55572 46392 -55430
rect 47360 -55430 47366 -54898
rect 47400 -54898 47414 -54854
rect 48366 -54854 48426 -54586
rect 47400 -55430 47406 -54898
rect 48366 -54908 48384 -54854
rect 47360 -55442 47406 -55430
rect 48378 -55430 48384 -54908
rect 48418 -54892 48430 -54854
rect 48418 -54908 48426 -54892
rect 48418 -55430 48424 -54908
rect 48378 -55442 48424 -55430
rect 46630 -55480 47118 -55474
rect 46630 -55514 46642 -55480
rect 47106 -55514 47118 -55480
rect 46630 -55520 47118 -55514
rect 47648 -55480 48136 -55474
rect 47648 -55514 47660 -55480
rect 48124 -55514 48136 -55480
rect 47648 -55520 48136 -55514
rect 46326 -55632 46332 -55572
rect 46392 -55632 46398 -55572
rect 46852 -55682 46912 -55520
rect 47860 -55682 47920 -55520
rect 48478 -55572 48538 -49782
rect 48600 -50696 48606 -50636
rect 48666 -50696 48672 -50636
rect 48606 -52194 48666 -50696
rect 48722 -50960 48782 -49668
rect 48838 -50918 48844 -50858
rect 48904 -50918 48910 -50858
rect 48716 -51020 48722 -50960
rect 48782 -51020 48788 -50960
rect 48600 -52254 48606 -52194
rect 48666 -52254 48672 -52194
rect 48596 -53156 48602 -53096
rect 48662 -53156 48668 -53096
rect 48602 -54420 48662 -53156
rect 48722 -54322 48782 -51020
rect 48716 -54382 48722 -54322
rect 48782 -54382 48788 -54322
rect 48596 -54480 48602 -54420
rect 48662 -54480 48668 -54420
rect 48472 -55632 48478 -55572
rect 48538 -55632 48544 -55572
rect 46846 -55742 46852 -55682
rect 46912 -55742 46918 -55682
rect 47854 -55742 47860 -55682
rect 47920 -55742 47926 -55682
rect 48722 -55798 48782 -54382
rect 48844 -54654 48904 -50918
rect 48972 -52086 49032 -49564
rect 48970 -52092 49032 -52086
rect 49030 -52152 49032 -52092
rect 48970 -52158 49032 -52152
rect 48972 -54526 49032 -52158
rect 48966 -54586 48972 -54526
rect 49032 -54586 49038 -54526
rect 48838 -54714 48844 -54654
rect 48904 -54714 48910 -54654
rect 49094 -55682 49154 -44754
rect 49200 -48564 49206 -48504
rect 49266 -48564 49272 -48504
rect 49088 -55742 49094 -55682
rect 49154 -55742 49160 -55682
rect 46332 -55860 46338 -55800
rect 46398 -55860 46404 -55800
rect 47354 -55858 48782 -55798
rect 45612 -56004 46100 -55998
rect 45612 -56038 45624 -56004
rect 46088 -56038 46100 -56004
rect 45612 -56044 46100 -56038
rect 45316 -56134 45330 -56088
rect 44346 -56618 44352 -56154
rect 44346 -56664 44356 -56618
rect 43576 -56714 44064 -56708
rect 43576 -56748 43588 -56714
rect 44052 -56748 44064 -56714
rect 43576 -56754 44064 -56748
rect 43278 -56966 43284 -56906
rect 43344 -56966 43350 -56906
rect 43794 -57012 43854 -56754
rect 42770 -57072 42776 -57012
rect 42836 -57072 42842 -57012
rect 43788 -57072 43794 -57012
rect 43854 -57072 43860 -57012
rect 42258 -57182 42264 -57122
rect 42324 -57182 42330 -57122
rect 41540 -57236 42028 -57230
rect 41540 -57270 41552 -57236
rect 42016 -57270 42028 -57236
rect 41540 -57276 42028 -57270
rect 41244 -57356 41258 -57320
rect 38486 -57946 38974 -57940
rect 38486 -57980 38498 -57946
rect 38962 -57980 38974 -57946
rect 38486 -57986 38974 -57980
rect 39504 -57946 39992 -57940
rect 39504 -57980 39516 -57946
rect 39980 -57980 39992 -57946
rect 39504 -57986 39992 -57980
rect 38700 -58152 38760 -57986
rect 39710 -58146 39770 -57986
rect 38700 -58218 38760 -58212
rect 39708 -58152 39770 -58146
rect 39768 -58158 39770 -58152
rect 39708 -58218 39768 -58212
rect 40232 -58408 40292 -57896
rect 41252 -57896 41258 -57356
rect 41292 -57356 41304 -57320
rect 42264 -57320 42324 -57182
rect 42776 -57230 42836 -57072
rect 43794 -57230 43854 -57072
rect 44296 -57122 44356 -56664
rect 45324 -56664 45330 -56134
rect 45364 -56134 45376 -56088
rect 46338 -56088 46398 -55860
rect 46630 -56004 47118 -55998
rect 46630 -56038 46642 -56004
rect 47106 -56038 47118 -56004
rect 46630 -56044 47118 -56038
rect 45364 -56664 45370 -56134
rect 46338 -56148 46348 -56088
rect 46342 -56640 46348 -56148
rect 45324 -56676 45370 -56664
rect 46336 -56664 46348 -56640
rect 46382 -56148 46398 -56088
rect 47354 -56088 47414 -55858
rect 47852 -55998 47912 -55858
rect 47648 -56004 48136 -55998
rect 47648 -56038 47660 -56004
rect 48124 -56038 48136 -56004
rect 47648 -56044 48136 -56038
rect 46382 -56640 46388 -56148
rect 46382 -56664 46396 -56640
rect 44594 -56714 45082 -56708
rect 44594 -56748 44606 -56714
rect 45070 -56748 45082 -56714
rect 44594 -56754 45082 -56748
rect 45612 -56714 46100 -56708
rect 45612 -56748 45624 -56714
rect 46088 -56748 46100 -56714
rect 45612 -56754 46100 -56748
rect 44808 -57012 44868 -56754
rect 45308 -56966 45314 -56906
rect 45374 -56966 45380 -56906
rect 44802 -57072 44808 -57012
rect 44868 -57072 44874 -57012
rect 44290 -57182 44296 -57122
rect 44356 -57182 44362 -57122
rect 42558 -57236 43046 -57230
rect 42558 -57270 42570 -57236
rect 43034 -57270 43046 -57236
rect 42558 -57276 43046 -57270
rect 43576 -57236 44064 -57230
rect 43576 -57270 43588 -57236
rect 44052 -57270 44064 -57236
rect 43576 -57276 44064 -57270
rect 41292 -57896 41298 -57356
rect 41252 -57908 41298 -57896
rect 42264 -57896 42276 -57320
rect 42310 -57896 42324 -57320
rect 43288 -57320 43334 -57308
rect 43288 -57844 43294 -57320
rect 41748 -57940 41808 -57938
rect 40522 -57946 41010 -57940
rect 40522 -57980 40534 -57946
rect 40998 -57980 41010 -57946
rect 40522 -57986 41010 -57980
rect 41540 -57946 42028 -57940
rect 41540 -57980 41552 -57946
rect 42016 -57980 42028 -57946
rect 41540 -57986 42028 -57980
rect 40726 -58146 40786 -57986
rect 40724 -58152 40786 -58146
rect 40784 -58158 40786 -58152
rect 41748 -58152 41808 -57986
rect 40724 -58218 40784 -58212
rect 41748 -58218 41808 -58212
rect 42264 -58408 42324 -57896
rect 43278 -57896 43294 -57844
rect 43328 -57844 43334 -57320
rect 44296 -57320 44356 -57182
rect 44808 -57230 44868 -57072
rect 44594 -57236 45082 -57230
rect 44594 -57270 44606 -57236
rect 45070 -57270 45082 -57236
rect 44594 -57276 45082 -57270
rect 43328 -57896 43338 -57844
rect 42558 -57946 43046 -57940
rect 42558 -57980 42570 -57946
rect 43034 -57980 43046 -57946
rect 42558 -57986 43046 -57980
rect 42770 -58152 42830 -57986
rect 43278 -58044 43338 -57896
rect 44296 -57896 44312 -57320
rect 44346 -57896 44356 -57320
rect 45314 -57320 45374 -56966
rect 45822 -57012 45882 -56754
rect 45816 -57072 45822 -57012
rect 45882 -57072 45888 -57012
rect 45822 -57230 45882 -57072
rect 46336 -57122 46396 -56664
rect 47354 -56664 47366 -56088
rect 47400 -56664 47414 -56088
rect 48368 -56088 48428 -55858
rect 48492 -55964 48498 -55904
rect 48558 -55964 48564 -55904
rect 48368 -56142 48384 -56088
rect 46630 -56714 47118 -56708
rect 46630 -56748 46642 -56714
rect 47106 -56748 47118 -56714
rect 46630 -56754 47118 -56748
rect 46844 -57012 46904 -56754
rect 47354 -56800 47414 -56664
rect 48378 -56664 48384 -56142
rect 48418 -56142 48428 -56088
rect 48418 -56664 48424 -56142
rect 48378 -56676 48424 -56664
rect 47648 -56714 48136 -56708
rect 47648 -56748 47660 -56714
rect 48124 -56748 48136 -56714
rect 47648 -56754 48136 -56748
rect 47348 -56860 47354 -56800
rect 47414 -56860 47420 -56800
rect 47348 -56966 47354 -56906
rect 47414 -56966 47420 -56906
rect 46838 -57072 46844 -57012
rect 46904 -57072 46910 -57012
rect 46330 -57182 46336 -57122
rect 46396 -57182 46402 -57122
rect 45612 -57236 46100 -57230
rect 45612 -57270 45624 -57236
rect 46088 -57270 46100 -57236
rect 45612 -57276 46100 -57270
rect 45314 -57364 45330 -57320
rect 43576 -57946 44064 -57940
rect 43576 -57980 43588 -57946
rect 44052 -57980 44064 -57946
rect 43576 -57986 44064 -57980
rect 43272 -58104 43278 -58044
rect 43338 -58104 43344 -58044
rect 43790 -58146 43850 -57986
rect 43790 -58152 43852 -58146
rect 43790 -58158 43792 -58152
rect 42770 -58218 42830 -58212
rect 43792 -58218 43852 -58212
rect 44296 -58408 44356 -57896
rect 45324 -57896 45330 -57364
rect 45364 -57364 45374 -57320
rect 46336 -57320 46396 -57182
rect 46844 -57230 46904 -57072
rect 47354 -57122 47414 -56966
rect 47354 -57182 48432 -57122
rect 46630 -57236 47118 -57230
rect 46630 -57270 46642 -57236
rect 47106 -57270 47118 -57236
rect 46630 -57276 47118 -57270
rect 45364 -57896 45370 -57364
rect 45324 -57908 45370 -57896
rect 46336 -57896 46348 -57320
rect 46382 -57896 46396 -57320
rect 47354 -57320 47414 -57182
rect 47870 -57230 47930 -57182
rect 47648 -57236 48136 -57230
rect 47648 -57270 47660 -57236
rect 48124 -57270 48136 -57236
rect 47648 -57276 48136 -57270
rect 47354 -57328 47366 -57320
rect 44812 -57940 44872 -57938
rect 44594 -57946 45082 -57940
rect 44594 -57980 44606 -57946
rect 45070 -57980 45082 -57946
rect 44594 -57986 45082 -57980
rect 45612 -57946 46100 -57940
rect 45612 -57980 45624 -57946
rect 46088 -57980 46100 -57946
rect 45612 -57986 46100 -57980
rect 44812 -58146 44872 -57986
rect 45826 -58146 45886 -57986
rect 44810 -58152 44872 -58146
rect 44870 -58158 44872 -58152
rect 45824 -58152 45886 -58146
rect 44810 -58218 44870 -58212
rect 45884 -58158 45886 -58152
rect 45824 -58218 45884 -58212
rect 46336 -58408 46396 -57896
rect 47360 -57896 47366 -57328
rect 47400 -57328 47414 -57320
rect 48372 -57320 48432 -57182
rect 47400 -57896 47406 -57328
rect 48372 -57338 48384 -57320
rect 47360 -57908 47406 -57896
rect 48378 -57896 48384 -57338
rect 48418 -57338 48432 -57320
rect 48418 -57896 48424 -57338
rect 48378 -57908 48424 -57896
rect 46846 -57940 46906 -57938
rect 46630 -57946 47118 -57940
rect 46630 -57980 46642 -57946
rect 47106 -57980 47118 -57946
rect 46630 -57986 47118 -57980
rect 47648 -57946 48136 -57940
rect 47648 -57980 47660 -57946
rect 48124 -57980 48136 -57946
rect 47648 -57986 48136 -57980
rect 46846 -58146 46906 -57986
rect 48498 -58044 48558 -55964
rect 49206 -56906 49266 -48564
rect 49200 -56966 49206 -56906
rect 49266 -56966 49272 -56906
rect 48492 -58104 48498 -58044
rect 48558 -58104 48564 -58044
rect 46846 -58152 46908 -58146
rect 46846 -58158 46848 -58152
rect 46848 -58218 46908 -58212
rect 50260 -58308 50266 -44048
rect 50366 -58308 50372 -44048
rect 17326 -58454 17476 -58408
rect 17522 -58454 20696 -58408
rect 20756 -58454 27148 -58408
rect 27208 -58454 49250 -58408
rect 49310 -58454 49412 -58408
rect 17326 -58608 17372 -58454
rect 49372 -58608 49412 -58454
rect 17326 -58654 49412 -58608
rect 13828 -59094 13838 -58794
rect 49650 -59094 49660 -58794
rect 50260 -59094 50372 -58308
rect 13116 -59100 50372 -59094
rect 13116 -59200 13222 -59100
rect 50266 -59200 50372 -59100
rect 13116 -59206 50372 -59200
rect -27690 -64426 -25354 -64420
rect -27690 -64526 -27584 -64426
rect -25460 -64526 -25354 -64426
rect -27690 -64532 -25354 -64526
rect -27690 -64666 -27578 -64532
rect -27690 -67234 -27684 -64666
rect -28072 -67265 -27684 -67234
rect -28072 -67299 -28043 -67265
rect -28009 -67299 -27951 -67265
rect -27917 -67299 -27859 -67265
rect -27825 -67290 -27684 -67265
rect -27584 -67290 -27578 -64666
rect -26978 -64832 -26968 -64532
rect -26076 -64832 -26066 -64532
rect -25466 -64666 -25354 -64532
rect -27422 -65036 -25520 -65006
rect -27422 -65100 -27388 -65036
rect -25564 -65100 -25520 -65036
rect -27422 -65130 -25520 -65100
rect -27348 -65394 -27288 -65130
rect -27218 -65394 -27158 -65130
rect -26840 -65274 -26834 -65214
rect -26774 -65274 -26768 -65214
rect -26322 -65274 -26316 -65214
rect -26256 -65274 -26250 -65214
rect -27502 -65506 -27496 -65446
rect -27436 -65506 -27430 -65446
rect -27348 -65454 -27158 -65394
rect -27496 -66040 -27436 -65506
rect -27348 -65637 -27288 -65454
rect -27218 -65538 -27158 -65454
rect -27245 -65544 -27137 -65538
rect -27245 -65578 -27233 -65544
rect -27149 -65578 -27137 -65544
rect -27245 -65584 -27137 -65578
rect -26987 -65544 -26879 -65538
rect -26987 -65578 -26975 -65544
rect -26891 -65578 -26879 -65544
rect -26987 -65584 -26879 -65578
rect -27348 -65670 -27337 -65637
rect -27343 -65970 -27337 -65670
rect -27496 -67020 -27436 -66100
rect -27348 -66013 -27337 -65970
rect -27303 -65670 -27288 -65637
rect -27085 -65637 -27039 -65625
rect -27303 -65970 -27297 -65670
rect -27303 -66013 -27288 -65970
rect -27085 -65988 -27079 -65637
rect -27348 -66236 -27288 -66013
rect -27092 -66013 -27079 -65988
rect -27045 -65988 -27039 -65637
rect -26834 -65637 -26774 -65274
rect -26584 -65386 -26578 -65326
rect -26518 -65386 -26512 -65326
rect -26712 -65506 -26706 -65446
rect -26646 -65506 -26640 -65446
rect -26706 -65538 -26646 -65506
rect -26729 -65544 -26621 -65538
rect -26729 -65578 -26717 -65544
rect -26633 -65578 -26621 -65544
rect -26729 -65584 -26621 -65578
rect -27045 -66013 -27032 -65988
rect -27245 -66072 -27137 -66066
rect -27245 -66106 -27233 -66072
rect -27149 -66106 -27137 -66072
rect -27245 -66112 -27137 -66106
rect -27218 -66236 -27158 -66112
rect -27348 -66296 -27158 -66236
rect -27092 -66284 -27032 -66013
rect -26834 -66013 -26821 -65637
rect -26787 -66013 -26774 -65637
rect -26578 -65637 -26518 -65386
rect -26456 -65506 -26450 -65446
rect -26390 -65506 -26384 -65446
rect -26450 -65538 -26390 -65506
rect -26471 -65544 -26363 -65538
rect -26471 -65578 -26459 -65544
rect -26375 -65578 -26363 -65544
rect -26471 -65584 -26363 -65578
rect -26578 -65670 -26563 -65637
rect -26987 -66072 -26879 -66066
rect -26987 -66106 -26975 -66072
rect -26891 -66106 -26879 -66072
rect -26987 -66112 -26879 -66106
rect -26962 -66170 -26902 -66112
rect -26968 -66230 -26962 -66170
rect -26902 -66230 -26896 -66170
rect -27348 -66497 -27288 -66296
rect -27218 -66398 -27158 -66296
rect -27098 -66344 -27092 -66284
rect -27032 -66344 -27026 -66284
rect -27245 -66404 -27137 -66398
rect -27245 -66438 -27233 -66404
rect -27149 -66438 -27137 -66404
rect -27245 -66444 -27137 -66438
rect -26987 -66404 -26879 -66398
rect -26987 -66438 -26975 -66404
rect -26891 -66438 -26879 -66404
rect -26987 -66444 -26879 -66438
rect -27348 -66550 -27337 -66497
rect -27343 -66873 -27337 -66550
rect -27303 -66550 -27288 -66497
rect -27085 -66497 -27039 -66485
rect -27303 -66873 -27297 -66550
rect -27085 -66828 -27079 -66497
rect -27343 -66885 -27297 -66873
rect -27094 -66873 -27079 -66828
rect -27045 -66828 -27039 -66497
rect -26834 -66497 -26774 -66013
rect -26569 -66013 -26563 -65670
rect -26529 -65670 -26518 -65637
rect -26316 -65637 -26256 -65274
rect -25928 -65406 -25868 -65130
rect -25800 -65406 -25740 -65130
rect -25654 -65386 -25648 -65326
rect -25588 -65386 -25582 -65326
rect -25928 -65466 -25740 -65406
rect -25928 -65538 -25868 -65466
rect -26213 -65544 -26105 -65538
rect -26213 -65578 -26201 -65544
rect -26117 -65578 -26105 -65544
rect -26213 -65584 -26105 -65578
rect -25955 -65544 -25847 -65538
rect -25955 -65578 -25943 -65544
rect -25859 -65578 -25847 -65544
rect -25955 -65584 -25847 -65578
rect -26529 -66013 -26523 -65670
rect -26316 -65698 -26305 -65637
rect -26311 -65956 -26305 -65698
rect -26569 -66025 -26523 -66013
rect -26322 -66013 -26305 -65956
rect -26271 -65698 -26256 -65637
rect -26053 -65637 -26007 -65625
rect -26271 -65956 -26265 -65698
rect -26271 -66013 -26262 -65956
rect -26053 -65964 -26047 -65637
rect -26729 -66072 -26621 -66066
rect -26729 -66106 -26717 -66072
rect -26633 -66106 -26621 -66072
rect -26729 -66112 -26621 -66106
rect -26471 -66072 -26363 -66066
rect -26471 -66106 -26459 -66072
rect -26375 -66106 -26363 -66072
rect -26471 -66112 -26363 -66106
rect -26710 -66230 -26704 -66170
rect -26644 -66230 -26638 -66170
rect -26452 -66230 -26446 -66170
rect -26386 -66230 -26380 -66170
rect -26704 -66398 -26644 -66230
rect -26580 -66344 -26574 -66284
rect -26514 -66344 -26508 -66284
rect -26729 -66404 -26621 -66398
rect -26729 -66438 -26717 -66404
rect -26633 -66438 -26621 -66404
rect -26729 -66444 -26621 -66438
rect -27045 -66873 -27034 -66828
rect -26834 -66836 -26821 -66497
rect -27245 -66932 -27137 -66926
rect -27245 -66966 -27233 -66932
rect -27149 -66966 -27137 -66932
rect -27245 -66972 -27137 -66966
rect -27496 -67080 -27246 -67020
rect -27186 -67080 -27180 -67020
rect -27094 -67132 -27034 -66873
rect -26827 -66873 -26821 -66836
rect -26787 -66836 -26774 -66497
rect -26574 -66497 -26514 -66344
rect -26446 -66398 -26386 -66230
rect -26471 -66404 -26363 -66398
rect -26471 -66438 -26459 -66404
rect -26375 -66438 -26363 -66404
rect -26471 -66444 -26363 -66438
rect -26574 -66530 -26563 -66497
rect -26569 -66834 -26563 -66530
rect -26787 -66873 -26781 -66836
rect -26827 -66885 -26781 -66873
rect -26578 -66873 -26563 -66834
rect -26529 -66530 -26514 -66497
rect -26322 -66497 -26262 -66013
rect -26058 -66013 -26047 -65964
rect -26013 -65964 -26007 -65637
rect -25800 -65637 -25740 -65466
rect -26013 -66013 -25998 -65964
rect -26213 -66072 -26105 -66066
rect -26213 -66106 -26201 -66072
rect -26117 -66106 -26105 -66072
rect -26213 -66112 -26105 -66106
rect -26188 -66170 -26128 -66112
rect -26194 -66230 -26188 -66170
rect -26128 -66230 -26122 -66170
rect -26058 -66284 -25998 -66013
rect -25800 -66013 -25789 -65637
rect -25755 -66013 -25740 -65637
rect -25955 -66072 -25847 -66066
rect -25955 -66106 -25943 -66072
rect -25859 -66106 -25847 -66072
rect -25955 -66112 -25847 -66106
rect -25800 -66228 -25740 -66013
rect -26064 -66344 -26058 -66284
rect -25998 -66344 -25992 -66284
rect -25932 -66288 -25740 -66228
rect -25932 -66398 -25872 -66288
rect -26213 -66404 -26105 -66398
rect -26213 -66438 -26201 -66404
rect -26117 -66438 -26105 -66404
rect -26213 -66444 -26105 -66438
rect -25955 -66404 -25847 -66398
rect -25955 -66438 -25943 -66404
rect -25859 -66438 -25847 -66404
rect -25955 -66444 -25847 -66438
rect -26529 -66834 -26523 -66530
rect -26322 -66542 -26305 -66497
rect -26311 -66820 -26305 -66542
rect -26529 -66873 -26518 -66834
rect -26987 -66932 -26879 -66926
rect -26987 -66966 -26975 -66932
rect -26891 -66966 -26879 -66932
rect -26987 -66972 -26879 -66966
rect -26729 -66932 -26621 -66926
rect -26729 -66966 -26717 -66932
rect -26633 -66966 -26621 -66932
rect -26729 -66972 -26621 -66966
rect -26962 -67020 -26902 -66972
rect -26968 -67080 -26962 -67020
rect -26902 -67080 -26896 -67020
rect -27100 -67192 -27094 -67132
rect -27034 -67192 -27028 -67132
rect -26578 -67280 -26518 -66873
rect -26320 -66873 -26305 -66820
rect -26271 -66542 -26262 -66497
rect -26053 -66497 -26007 -66485
rect -26271 -66820 -26265 -66542
rect -26053 -66796 -26047 -66497
rect -26271 -66873 -26260 -66820
rect -26471 -66932 -26363 -66926
rect -26471 -66966 -26459 -66932
rect -26375 -66966 -26363 -66932
rect -26471 -66972 -26363 -66966
rect -26450 -67026 -26390 -66972
rect -26320 -67240 -26260 -66873
rect -26058 -66873 -26047 -66796
rect -26013 -66796 -26007 -66497
rect -25800 -66497 -25740 -66288
rect -26013 -66873 -25998 -66796
rect -26213 -66932 -26105 -66926
rect -26213 -66966 -26201 -66932
rect -26117 -66966 -26105 -66932
rect -26213 -66972 -26105 -66966
rect -26186 -67020 -26126 -66972
rect -26192 -67080 -26186 -67020
rect -26126 -67080 -26120 -67020
rect -26058 -67132 -25998 -66873
rect -25800 -66873 -25789 -66497
rect -25755 -66873 -25740 -66497
rect -25955 -66932 -25847 -66926
rect -25955 -66966 -25943 -66932
rect -25859 -66966 -25847 -66932
rect -25955 -66972 -25847 -66966
rect -25934 -67018 -25874 -66972
rect -25800 -67018 -25740 -66873
rect -25934 -67078 -25740 -67018
rect -26064 -67192 -26058 -67132
rect -25998 -67192 -25992 -67132
rect -27825 -67299 -27578 -67290
rect -28072 -67330 -27578 -67299
rect -27690 -67424 -27578 -67330
rect -26584 -67340 -26578 -67280
rect -26518 -67340 -26512 -67280
rect -26326 -67300 -26320 -67240
rect -26260 -67300 -26254 -67240
rect -25934 -67424 -25874 -67078
rect -25800 -67424 -25740 -67078
rect -25648 -67132 -25588 -65386
rect -25654 -67192 -25648 -67132
rect -25588 -67192 -25582 -67132
rect -25466 -67290 -25460 -64666
rect -25360 -67290 -25354 -64666
rect -23690 -64426 -21354 -64420
rect -23690 -64526 -23584 -64426
rect -21460 -64526 -21354 -64426
rect -23690 -64532 -21354 -64526
rect -23690 -64666 -23578 -64532
rect -23690 -67234 -23684 -64666
rect -25466 -67424 -25354 -67290
rect -24072 -67265 -23684 -67234
rect -24072 -67299 -24043 -67265
rect -24009 -67299 -23951 -67265
rect -23917 -67299 -23859 -67265
rect -23825 -67290 -23684 -67265
rect -23584 -67290 -23578 -64666
rect -22978 -64832 -22968 -64532
rect -22076 -64832 -22066 -64532
rect -21466 -64666 -21354 -64532
rect -23422 -65036 -21520 -65006
rect -23422 -65100 -23388 -65036
rect -21564 -65100 -21520 -65036
rect -23422 -65130 -21520 -65100
rect -23348 -65394 -23288 -65130
rect -23218 -65394 -23158 -65130
rect -22840 -65274 -22834 -65214
rect -22774 -65274 -22768 -65214
rect -22322 -65274 -22316 -65214
rect -22256 -65274 -22250 -65214
rect -23502 -65506 -23496 -65446
rect -23436 -65506 -23430 -65446
rect -23348 -65454 -23158 -65394
rect -23496 -66040 -23436 -65506
rect -23348 -65637 -23288 -65454
rect -23218 -65538 -23158 -65454
rect -23245 -65544 -23137 -65538
rect -23245 -65578 -23233 -65544
rect -23149 -65578 -23137 -65544
rect -23245 -65584 -23137 -65578
rect -22987 -65544 -22879 -65538
rect -22987 -65578 -22975 -65544
rect -22891 -65578 -22879 -65544
rect -22987 -65584 -22879 -65578
rect -23348 -65670 -23337 -65637
rect -23343 -65970 -23337 -65670
rect -23496 -67020 -23436 -66100
rect -23348 -66013 -23337 -65970
rect -23303 -65670 -23288 -65637
rect -23085 -65637 -23039 -65625
rect -23303 -65970 -23297 -65670
rect -23303 -66013 -23288 -65970
rect -23085 -65988 -23079 -65637
rect -23348 -66236 -23288 -66013
rect -23092 -66013 -23079 -65988
rect -23045 -65988 -23039 -65637
rect -22834 -65637 -22774 -65274
rect -22584 -65386 -22578 -65326
rect -22518 -65386 -22512 -65326
rect -22712 -65506 -22706 -65446
rect -22646 -65506 -22640 -65446
rect -22706 -65538 -22646 -65506
rect -22729 -65544 -22621 -65538
rect -22729 -65578 -22717 -65544
rect -22633 -65578 -22621 -65544
rect -22729 -65584 -22621 -65578
rect -23045 -66013 -23032 -65988
rect -23245 -66072 -23137 -66066
rect -23245 -66106 -23233 -66072
rect -23149 -66106 -23137 -66072
rect -23245 -66112 -23137 -66106
rect -23218 -66236 -23158 -66112
rect -23348 -66296 -23158 -66236
rect -23092 -66284 -23032 -66013
rect -22834 -66013 -22821 -65637
rect -22787 -66013 -22774 -65637
rect -22578 -65637 -22518 -65386
rect -22456 -65506 -22450 -65446
rect -22390 -65506 -22384 -65446
rect -22450 -65538 -22390 -65506
rect -22471 -65544 -22363 -65538
rect -22471 -65578 -22459 -65544
rect -22375 -65578 -22363 -65544
rect -22471 -65584 -22363 -65578
rect -22578 -65670 -22563 -65637
rect -22987 -66072 -22879 -66066
rect -22987 -66106 -22975 -66072
rect -22891 -66106 -22879 -66072
rect -22987 -66112 -22879 -66106
rect -22962 -66170 -22902 -66112
rect -22968 -66230 -22962 -66170
rect -22902 -66230 -22896 -66170
rect -23348 -66497 -23288 -66296
rect -23218 -66398 -23158 -66296
rect -23098 -66344 -23092 -66284
rect -23032 -66344 -23026 -66284
rect -23245 -66404 -23137 -66398
rect -23245 -66438 -23233 -66404
rect -23149 -66438 -23137 -66404
rect -23245 -66444 -23137 -66438
rect -22987 -66404 -22879 -66398
rect -22987 -66438 -22975 -66404
rect -22891 -66438 -22879 -66404
rect -22987 -66444 -22879 -66438
rect -23348 -66550 -23337 -66497
rect -23343 -66873 -23337 -66550
rect -23303 -66550 -23288 -66497
rect -23085 -66497 -23039 -66485
rect -23303 -66873 -23297 -66550
rect -23085 -66828 -23079 -66497
rect -23343 -66885 -23297 -66873
rect -23094 -66873 -23079 -66828
rect -23045 -66828 -23039 -66497
rect -22834 -66497 -22774 -66013
rect -22569 -66013 -22563 -65670
rect -22529 -65670 -22518 -65637
rect -22316 -65637 -22256 -65274
rect -21928 -65406 -21868 -65130
rect -21800 -65406 -21740 -65130
rect -21654 -65386 -21648 -65326
rect -21588 -65386 -21582 -65326
rect -21928 -65466 -21740 -65406
rect -21928 -65538 -21868 -65466
rect -22213 -65544 -22105 -65538
rect -22213 -65578 -22201 -65544
rect -22117 -65578 -22105 -65544
rect -22213 -65584 -22105 -65578
rect -21955 -65544 -21847 -65538
rect -21955 -65578 -21943 -65544
rect -21859 -65578 -21847 -65544
rect -21955 -65584 -21847 -65578
rect -22529 -66013 -22523 -65670
rect -22316 -65698 -22305 -65637
rect -22311 -65956 -22305 -65698
rect -22569 -66025 -22523 -66013
rect -22322 -66013 -22305 -65956
rect -22271 -65698 -22256 -65637
rect -22053 -65637 -22007 -65625
rect -22271 -65956 -22265 -65698
rect -22271 -66013 -22262 -65956
rect -22053 -65964 -22047 -65637
rect -22729 -66072 -22621 -66066
rect -22729 -66106 -22717 -66072
rect -22633 -66106 -22621 -66072
rect -22729 -66112 -22621 -66106
rect -22471 -66072 -22363 -66066
rect -22471 -66106 -22459 -66072
rect -22375 -66106 -22363 -66072
rect -22471 -66112 -22363 -66106
rect -22710 -66230 -22704 -66170
rect -22644 -66230 -22638 -66170
rect -22452 -66230 -22446 -66170
rect -22386 -66230 -22380 -66170
rect -22704 -66398 -22644 -66230
rect -22580 -66344 -22574 -66284
rect -22514 -66344 -22508 -66284
rect -22729 -66404 -22621 -66398
rect -22729 -66438 -22717 -66404
rect -22633 -66438 -22621 -66404
rect -22729 -66444 -22621 -66438
rect -23045 -66873 -23034 -66828
rect -22834 -66836 -22821 -66497
rect -23245 -66932 -23137 -66926
rect -23245 -66966 -23233 -66932
rect -23149 -66966 -23137 -66932
rect -23245 -66972 -23137 -66966
rect -23496 -67080 -23246 -67020
rect -23186 -67080 -23180 -67020
rect -23094 -67132 -23034 -66873
rect -22827 -66873 -22821 -66836
rect -22787 -66836 -22774 -66497
rect -22574 -66497 -22514 -66344
rect -22446 -66398 -22386 -66230
rect -22471 -66404 -22363 -66398
rect -22471 -66438 -22459 -66404
rect -22375 -66438 -22363 -66404
rect -22471 -66444 -22363 -66438
rect -22574 -66530 -22563 -66497
rect -22569 -66834 -22563 -66530
rect -22787 -66873 -22781 -66836
rect -22827 -66885 -22781 -66873
rect -22578 -66873 -22563 -66834
rect -22529 -66530 -22514 -66497
rect -22322 -66497 -22262 -66013
rect -22058 -66013 -22047 -65964
rect -22013 -65964 -22007 -65637
rect -21800 -65637 -21740 -65466
rect -22013 -66013 -21998 -65964
rect -22213 -66072 -22105 -66066
rect -22213 -66106 -22201 -66072
rect -22117 -66106 -22105 -66072
rect -22213 -66112 -22105 -66106
rect -22188 -66170 -22128 -66112
rect -22194 -66230 -22188 -66170
rect -22128 -66230 -22122 -66170
rect -22058 -66284 -21998 -66013
rect -21800 -66013 -21789 -65637
rect -21755 -66013 -21740 -65637
rect -21955 -66072 -21847 -66066
rect -21955 -66106 -21943 -66072
rect -21859 -66106 -21847 -66072
rect -21955 -66112 -21847 -66106
rect -21800 -66228 -21740 -66013
rect -22064 -66344 -22058 -66284
rect -21998 -66344 -21992 -66284
rect -21932 -66288 -21740 -66228
rect -21932 -66398 -21872 -66288
rect -22213 -66404 -22105 -66398
rect -22213 -66438 -22201 -66404
rect -22117 -66438 -22105 -66404
rect -22213 -66444 -22105 -66438
rect -21955 -66404 -21847 -66398
rect -21955 -66438 -21943 -66404
rect -21859 -66438 -21847 -66404
rect -21955 -66444 -21847 -66438
rect -22529 -66834 -22523 -66530
rect -22322 -66542 -22305 -66497
rect -22311 -66820 -22305 -66542
rect -22529 -66873 -22518 -66834
rect -22987 -66932 -22879 -66926
rect -22987 -66966 -22975 -66932
rect -22891 -66966 -22879 -66932
rect -22987 -66972 -22879 -66966
rect -22729 -66932 -22621 -66926
rect -22729 -66966 -22717 -66932
rect -22633 -66966 -22621 -66932
rect -22729 -66972 -22621 -66966
rect -22962 -67020 -22902 -66972
rect -22968 -67080 -22962 -67020
rect -22902 -67080 -22896 -67020
rect -23100 -67192 -23094 -67132
rect -23034 -67192 -23028 -67132
rect -22578 -67280 -22518 -66873
rect -22320 -66873 -22305 -66820
rect -22271 -66542 -22262 -66497
rect -22053 -66497 -22007 -66485
rect -22271 -66820 -22265 -66542
rect -22053 -66796 -22047 -66497
rect -22271 -66873 -22260 -66820
rect -22471 -66932 -22363 -66926
rect -22471 -66966 -22459 -66932
rect -22375 -66966 -22363 -66932
rect -22471 -66972 -22363 -66966
rect -22450 -67026 -22390 -66972
rect -22320 -67240 -22260 -66873
rect -22058 -66873 -22047 -66796
rect -22013 -66796 -22007 -66497
rect -21800 -66497 -21740 -66288
rect -22013 -66873 -21998 -66796
rect -22213 -66932 -22105 -66926
rect -22213 -66966 -22201 -66932
rect -22117 -66966 -22105 -66932
rect -22213 -66972 -22105 -66966
rect -22186 -67020 -22126 -66972
rect -22192 -67080 -22186 -67020
rect -22126 -67080 -22120 -67020
rect -22058 -67132 -21998 -66873
rect -21800 -66873 -21789 -66497
rect -21755 -66873 -21740 -66497
rect -21955 -66932 -21847 -66926
rect -21955 -66966 -21943 -66932
rect -21859 -66966 -21847 -66932
rect -21955 -66972 -21847 -66966
rect -21934 -67018 -21874 -66972
rect -21800 -67018 -21740 -66873
rect -21934 -67078 -21740 -67018
rect -22064 -67192 -22058 -67132
rect -21998 -67192 -21992 -67132
rect -23825 -67299 -23578 -67290
rect -24072 -67330 -23578 -67299
rect -27690 -67430 -25354 -67424
rect -27690 -67530 -27584 -67430
rect -25460 -67530 -25354 -67430
rect -27690 -67536 -25354 -67530
rect -23690 -67424 -23578 -67330
rect -22584 -67340 -22578 -67280
rect -22518 -67340 -22512 -67280
rect -22326 -67300 -22320 -67240
rect -22260 -67300 -22254 -67240
rect -21934 -67424 -21874 -67078
rect -21800 -67424 -21740 -67078
rect -21648 -67132 -21588 -65386
rect -21654 -67192 -21648 -67132
rect -21588 -67192 -21582 -67132
rect -21466 -67290 -21460 -64666
rect -21360 -67290 -21354 -64666
rect -19690 -64426 -17354 -64420
rect -19690 -64526 -19584 -64426
rect -17460 -64526 -17354 -64426
rect -19690 -64532 -17354 -64526
rect -19690 -64666 -19578 -64532
rect -19690 -67234 -19684 -64666
rect -21466 -67424 -21354 -67290
rect -20072 -67265 -19684 -67234
rect -20072 -67299 -20043 -67265
rect -20009 -67299 -19951 -67265
rect -19917 -67299 -19859 -67265
rect -19825 -67290 -19684 -67265
rect -19584 -67290 -19578 -64666
rect -18978 -64832 -18968 -64532
rect -18076 -64832 -18066 -64532
rect -17466 -64666 -17354 -64532
rect -19422 -65036 -17520 -65006
rect -19422 -65100 -19388 -65036
rect -17564 -65100 -17520 -65036
rect -19422 -65130 -17520 -65100
rect -19348 -65394 -19288 -65130
rect -19218 -65394 -19158 -65130
rect -18840 -65274 -18834 -65214
rect -18774 -65274 -18768 -65214
rect -18322 -65274 -18316 -65214
rect -18256 -65274 -18250 -65214
rect -19502 -65506 -19496 -65446
rect -19436 -65506 -19430 -65446
rect -19348 -65454 -19158 -65394
rect -19496 -66040 -19436 -65506
rect -19348 -65637 -19288 -65454
rect -19218 -65538 -19158 -65454
rect -19245 -65544 -19137 -65538
rect -19245 -65578 -19233 -65544
rect -19149 -65578 -19137 -65544
rect -19245 -65584 -19137 -65578
rect -18987 -65544 -18879 -65538
rect -18987 -65578 -18975 -65544
rect -18891 -65578 -18879 -65544
rect -18987 -65584 -18879 -65578
rect -19348 -65670 -19337 -65637
rect -19343 -65970 -19337 -65670
rect -19496 -67020 -19436 -66100
rect -19348 -66013 -19337 -65970
rect -19303 -65670 -19288 -65637
rect -19085 -65637 -19039 -65625
rect -19303 -65970 -19297 -65670
rect -19303 -66013 -19288 -65970
rect -19085 -65988 -19079 -65637
rect -19348 -66236 -19288 -66013
rect -19092 -66013 -19079 -65988
rect -19045 -65988 -19039 -65637
rect -18834 -65637 -18774 -65274
rect -18584 -65386 -18578 -65326
rect -18518 -65386 -18512 -65326
rect -18712 -65506 -18706 -65446
rect -18646 -65506 -18640 -65446
rect -18706 -65538 -18646 -65506
rect -18729 -65544 -18621 -65538
rect -18729 -65578 -18717 -65544
rect -18633 -65578 -18621 -65544
rect -18729 -65584 -18621 -65578
rect -19045 -66013 -19032 -65988
rect -19245 -66072 -19137 -66066
rect -19245 -66106 -19233 -66072
rect -19149 -66106 -19137 -66072
rect -19245 -66112 -19137 -66106
rect -19218 -66236 -19158 -66112
rect -19348 -66296 -19158 -66236
rect -19092 -66284 -19032 -66013
rect -18834 -66013 -18821 -65637
rect -18787 -66013 -18774 -65637
rect -18578 -65637 -18518 -65386
rect -18456 -65506 -18450 -65446
rect -18390 -65506 -18384 -65446
rect -18450 -65538 -18390 -65506
rect -18471 -65544 -18363 -65538
rect -18471 -65578 -18459 -65544
rect -18375 -65578 -18363 -65544
rect -18471 -65584 -18363 -65578
rect -18578 -65670 -18563 -65637
rect -18987 -66072 -18879 -66066
rect -18987 -66106 -18975 -66072
rect -18891 -66106 -18879 -66072
rect -18987 -66112 -18879 -66106
rect -18962 -66170 -18902 -66112
rect -18968 -66230 -18962 -66170
rect -18902 -66230 -18896 -66170
rect -19348 -66497 -19288 -66296
rect -19218 -66398 -19158 -66296
rect -19098 -66344 -19092 -66284
rect -19032 -66344 -19026 -66284
rect -19245 -66404 -19137 -66398
rect -19245 -66438 -19233 -66404
rect -19149 -66438 -19137 -66404
rect -19245 -66444 -19137 -66438
rect -18987 -66404 -18879 -66398
rect -18987 -66438 -18975 -66404
rect -18891 -66438 -18879 -66404
rect -18987 -66444 -18879 -66438
rect -19348 -66550 -19337 -66497
rect -19343 -66873 -19337 -66550
rect -19303 -66550 -19288 -66497
rect -19085 -66497 -19039 -66485
rect -19303 -66873 -19297 -66550
rect -19085 -66828 -19079 -66497
rect -19343 -66885 -19297 -66873
rect -19094 -66873 -19079 -66828
rect -19045 -66828 -19039 -66497
rect -18834 -66497 -18774 -66013
rect -18569 -66013 -18563 -65670
rect -18529 -65670 -18518 -65637
rect -18316 -65637 -18256 -65274
rect -17928 -65406 -17868 -65130
rect -17800 -65406 -17740 -65130
rect -17654 -65386 -17648 -65326
rect -17588 -65386 -17582 -65326
rect -17928 -65466 -17740 -65406
rect -17928 -65538 -17868 -65466
rect -18213 -65544 -18105 -65538
rect -18213 -65578 -18201 -65544
rect -18117 -65578 -18105 -65544
rect -18213 -65584 -18105 -65578
rect -17955 -65544 -17847 -65538
rect -17955 -65578 -17943 -65544
rect -17859 -65578 -17847 -65544
rect -17955 -65584 -17847 -65578
rect -18529 -66013 -18523 -65670
rect -18316 -65698 -18305 -65637
rect -18311 -65956 -18305 -65698
rect -18569 -66025 -18523 -66013
rect -18322 -66013 -18305 -65956
rect -18271 -65698 -18256 -65637
rect -18053 -65637 -18007 -65625
rect -18271 -65956 -18265 -65698
rect -18271 -66013 -18262 -65956
rect -18053 -65964 -18047 -65637
rect -18729 -66072 -18621 -66066
rect -18729 -66106 -18717 -66072
rect -18633 -66106 -18621 -66072
rect -18729 -66112 -18621 -66106
rect -18471 -66072 -18363 -66066
rect -18471 -66106 -18459 -66072
rect -18375 -66106 -18363 -66072
rect -18471 -66112 -18363 -66106
rect -18710 -66230 -18704 -66170
rect -18644 -66230 -18638 -66170
rect -18452 -66230 -18446 -66170
rect -18386 -66230 -18380 -66170
rect -18704 -66398 -18644 -66230
rect -18580 -66344 -18574 -66284
rect -18514 -66344 -18508 -66284
rect -18729 -66404 -18621 -66398
rect -18729 -66438 -18717 -66404
rect -18633 -66438 -18621 -66404
rect -18729 -66444 -18621 -66438
rect -19045 -66873 -19034 -66828
rect -18834 -66836 -18821 -66497
rect -19245 -66932 -19137 -66926
rect -19245 -66966 -19233 -66932
rect -19149 -66966 -19137 -66932
rect -19245 -66972 -19137 -66966
rect -19496 -67080 -19246 -67020
rect -19186 -67080 -19180 -67020
rect -19094 -67132 -19034 -66873
rect -18827 -66873 -18821 -66836
rect -18787 -66836 -18774 -66497
rect -18574 -66497 -18514 -66344
rect -18446 -66398 -18386 -66230
rect -18471 -66404 -18363 -66398
rect -18471 -66438 -18459 -66404
rect -18375 -66438 -18363 -66404
rect -18471 -66444 -18363 -66438
rect -18574 -66530 -18563 -66497
rect -18569 -66834 -18563 -66530
rect -18787 -66873 -18781 -66836
rect -18827 -66885 -18781 -66873
rect -18578 -66873 -18563 -66834
rect -18529 -66530 -18514 -66497
rect -18322 -66497 -18262 -66013
rect -18058 -66013 -18047 -65964
rect -18013 -65964 -18007 -65637
rect -17800 -65637 -17740 -65466
rect -18013 -66013 -17998 -65964
rect -18213 -66072 -18105 -66066
rect -18213 -66106 -18201 -66072
rect -18117 -66106 -18105 -66072
rect -18213 -66112 -18105 -66106
rect -18188 -66170 -18128 -66112
rect -18194 -66230 -18188 -66170
rect -18128 -66230 -18122 -66170
rect -18058 -66284 -17998 -66013
rect -17800 -66013 -17789 -65637
rect -17755 -66013 -17740 -65637
rect -17955 -66072 -17847 -66066
rect -17955 -66106 -17943 -66072
rect -17859 -66106 -17847 -66072
rect -17955 -66112 -17847 -66106
rect -17800 -66228 -17740 -66013
rect -18064 -66344 -18058 -66284
rect -17998 -66344 -17992 -66284
rect -17932 -66288 -17740 -66228
rect -17932 -66398 -17872 -66288
rect -18213 -66404 -18105 -66398
rect -18213 -66438 -18201 -66404
rect -18117 -66438 -18105 -66404
rect -18213 -66444 -18105 -66438
rect -17955 -66404 -17847 -66398
rect -17955 -66438 -17943 -66404
rect -17859 -66438 -17847 -66404
rect -17955 -66444 -17847 -66438
rect -18529 -66834 -18523 -66530
rect -18322 -66542 -18305 -66497
rect -18311 -66820 -18305 -66542
rect -18529 -66873 -18518 -66834
rect -18987 -66932 -18879 -66926
rect -18987 -66966 -18975 -66932
rect -18891 -66966 -18879 -66932
rect -18987 -66972 -18879 -66966
rect -18729 -66932 -18621 -66926
rect -18729 -66966 -18717 -66932
rect -18633 -66966 -18621 -66932
rect -18729 -66972 -18621 -66966
rect -18962 -67020 -18902 -66972
rect -18968 -67080 -18962 -67020
rect -18902 -67080 -18896 -67020
rect -19100 -67192 -19094 -67132
rect -19034 -67192 -19028 -67132
rect -18578 -67280 -18518 -66873
rect -18320 -66873 -18305 -66820
rect -18271 -66542 -18262 -66497
rect -18053 -66497 -18007 -66485
rect -18271 -66820 -18265 -66542
rect -18053 -66796 -18047 -66497
rect -18271 -66873 -18260 -66820
rect -18471 -66932 -18363 -66926
rect -18471 -66966 -18459 -66932
rect -18375 -66966 -18363 -66932
rect -18471 -66972 -18363 -66966
rect -18450 -67026 -18390 -66972
rect -18320 -67240 -18260 -66873
rect -18058 -66873 -18047 -66796
rect -18013 -66796 -18007 -66497
rect -17800 -66497 -17740 -66288
rect -18013 -66873 -17998 -66796
rect -18213 -66932 -18105 -66926
rect -18213 -66966 -18201 -66932
rect -18117 -66966 -18105 -66932
rect -18213 -66972 -18105 -66966
rect -18186 -67020 -18126 -66972
rect -18192 -67080 -18186 -67020
rect -18126 -67080 -18120 -67020
rect -18058 -67132 -17998 -66873
rect -17800 -66873 -17789 -66497
rect -17755 -66873 -17740 -66497
rect -17955 -66932 -17847 -66926
rect -17955 -66966 -17943 -66932
rect -17859 -66966 -17847 -66932
rect -17955 -66972 -17847 -66966
rect -17934 -67018 -17874 -66972
rect -17800 -67018 -17740 -66873
rect -17934 -67078 -17740 -67018
rect -18064 -67192 -18058 -67132
rect -17998 -67192 -17992 -67132
rect -19825 -67299 -19578 -67290
rect -20072 -67330 -19578 -67299
rect -23690 -67430 -21354 -67424
rect -23690 -67530 -23584 -67430
rect -21460 -67530 -21354 -67430
rect -23690 -67536 -21354 -67530
rect -19690 -67424 -19578 -67330
rect -18584 -67340 -18578 -67280
rect -18518 -67340 -18512 -67280
rect -18326 -67300 -18320 -67240
rect -18260 -67300 -18254 -67240
rect -17934 -67424 -17874 -67078
rect -17800 -67424 -17740 -67078
rect -17648 -67132 -17588 -65386
rect -17654 -67192 -17648 -67132
rect -17588 -67192 -17582 -67132
rect -17466 -67290 -17460 -64666
rect -17360 -67290 -17354 -64666
rect -15690 -64426 -13354 -64420
rect -15690 -64526 -15584 -64426
rect -13460 -64526 -13354 -64426
rect -15690 -64532 -13354 -64526
rect -15690 -64666 -15578 -64532
rect -15690 -67234 -15684 -64666
rect -17466 -67424 -17354 -67290
rect -16072 -67265 -15684 -67234
rect -16072 -67299 -16043 -67265
rect -16009 -67299 -15951 -67265
rect -15917 -67299 -15859 -67265
rect -15825 -67290 -15684 -67265
rect -15584 -67290 -15578 -64666
rect -14978 -64832 -14968 -64532
rect -14076 -64832 -14066 -64532
rect -13466 -64666 -13354 -64532
rect -15422 -65036 -13520 -65006
rect -15422 -65100 -15388 -65036
rect -13564 -65100 -13520 -65036
rect -15422 -65130 -13520 -65100
rect -15348 -65394 -15288 -65130
rect -15218 -65394 -15158 -65130
rect -14840 -65274 -14834 -65214
rect -14774 -65274 -14768 -65214
rect -14322 -65274 -14316 -65214
rect -14256 -65274 -14250 -65214
rect -15502 -65506 -15496 -65446
rect -15436 -65506 -15430 -65446
rect -15348 -65454 -15158 -65394
rect -15496 -66040 -15436 -65506
rect -15348 -65637 -15288 -65454
rect -15218 -65538 -15158 -65454
rect -15245 -65544 -15137 -65538
rect -15245 -65578 -15233 -65544
rect -15149 -65578 -15137 -65544
rect -15245 -65584 -15137 -65578
rect -14987 -65544 -14879 -65538
rect -14987 -65578 -14975 -65544
rect -14891 -65578 -14879 -65544
rect -14987 -65584 -14879 -65578
rect -15348 -65670 -15337 -65637
rect -15343 -65970 -15337 -65670
rect -15496 -67020 -15436 -66100
rect -15348 -66013 -15337 -65970
rect -15303 -65670 -15288 -65637
rect -15085 -65637 -15039 -65625
rect -15303 -65970 -15297 -65670
rect -15303 -66013 -15288 -65970
rect -15085 -65988 -15079 -65637
rect -15348 -66236 -15288 -66013
rect -15092 -66013 -15079 -65988
rect -15045 -65988 -15039 -65637
rect -14834 -65637 -14774 -65274
rect -14584 -65386 -14578 -65326
rect -14518 -65386 -14512 -65326
rect -14712 -65506 -14706 -65446
rect -14646 -65506 -14640 -65446
rect -14706 -65538 -14646 -65506
rect -14729 -65544 -14621 -65538
rect -14729 -65578 -14717 -65544
rect -14633 -65578 -14621 -65544
rect -14729 -65584 -14621 -65578
rect -15045 -66013 -15032 -65988
rect -15245 -66072 -15137 -66066
rect -15245 -66106 -15233 -66072
rect -15149 -66106 -15137 -66072
rect -15245 -66112 -15137 -66106
rect -15218 -66236 -15158 -66112
rect -15348 -66296 -15158 -66236
rect -15092 -66284 -15032 -66013
rect -14834 -66013 -14821 -65637
rect -14787 -66013 -14774 -65637
rect -14578 -65637 -14518 -65386
rect -14456 -65506 -14450 -65446
rect -14390 -65506 -14384 -65446
rect -14450 -65538 -14390 -65506
rect -14471 -65544 -14363 -65538
rect -14471 -65578 -14459 -65544
rect -14375 -65578 -14363 -65544
rect -14471 -65584 -14363 -65578
rect -14578 -65670 -14563 -65637
rect -14987 -66072 -14879 -66066
rect -14987 -66106 -14975 -66072
rect -14891 -66106 -14879 -66072
rect -14987 -66112 -14879 -66106
rect -14962 -66170 -14902 -66112
rect -14968 -66230 -14962 -66170
rect -14902 -66230 -14896 -66170
rect -15348 -66497 -15288 -66296
rect -15218 -66398 -15158 -66296
rect -15098 -66344 -15092 -66284
rect -15032 -66344 -15026 -66284
rect -15245 -66404 -15137 -66398
rect -15245 -66438 -15233 -66404
rect -15149 -66438 -15137 -66404
rect -15245 -66444 -15137 -66438
rect -14987 -66404 -14879 -66398
rect -14987 -66438 -14975 -66404
rect -14891 -66438 -14879 -66404
rect -14987 -66444 -14879 -66438
rect -15348 -66550 -15337 -66497
rect -15343 -66873 -15337 -66550
rect -15303 -66550 -15288 -66497
rect -15085 -66497 -15039 -66485
rect -15303 -66873 -15297 -66550
rect -15085 -66828 -15079 -66497
rect -15343 -66885 -15297 -66873
rect -15094 -66873 -15079 -66828
rect -15045 -66828 -15039 -66497
rect -14834 -66497 -14774 -66013
rect -14569 -66013 -14563 -65670
rect -14529 -65670 -14518 -65637
rect -14316 -65637 -14256 -65274
rect -13928 -65406 -13868 -65130
rect -13800 -65406 -13740 -65130
rect -13654 -65386 -13648 -65326
rect -13588 -65386 -13582 -65326
rect -13928 -65466 -13740 -65406
rect -13928 -65538 -13868 -65466
rect -14213 -65544 -14105 -65538
rect -14213 -65578 -14201 -65544
rect -14117 -65578 -14105 -65544
rect -14213 -65584 -14105 -65578
rect -13955 -65544 -13847 -65538
rect -13955 -65578 -13943 -65544
rect -13859 -65578 -13847 -65544
rect -13955 -65584 -13847 -65578
rect -14529 -66013 -14523 -65670
rect -14316 -65698 -14305 -65637
rect -14311 -65956 -14305 -65698
rect -14569 -66025 -14523 -66013
rect -14322 -66013 -14305 -65956
rect -14271 -65698 -14256 -65637
rect -14053 -65637 -14007 -65625
rect -14271 -65956 -14265 -65698
rect -14271 -66013 -14262 -65956
rect -14053 -65964 -14047 -65637
rect -14729 -66072 -14621 -66066
rect -14729 -66106 -14717 -66072
rect -14633 -66106 -14621 -66072
rect -14729 -66112 -14621 -66106
rect -14471 -66072 -14363 -66066
rect -14471 -66106 -14459 -66072
rect -14375 -66106 -14363 -66072
rect -14471 -66112 -14363 -66106
rect -14710 -66230 -14704 -66170
rect -14644 -66230 -14638 -66170
rect -14452 -66230 -14446 -66170
rect -14386 -66230 -14380 -66170
rect -14704 -66398 -14644 -66230
rect -14580 -66344 -14574 -66284
rect -14514 -66344 -14508 -66284
rect -14729 -66404 -14621 -66398
rect -14729 -66438 -14717 -66404
rect -14633 -66438 -14621 -66404
rect -14729 -66444 -14621 -66438
rect -15045 -66873 -15034 -66828
rect -14834 -66836 -14821 -66497
rect -15245 -66932 -15137 -66926
rect -15245 -66966 -15233 -66932
rect -15149 -66966 -15137 -66932
rect -15245 -66972 -15137 -66966
rect -15496 -67080 -15246 -67020
rect -15186 -67080 -15180 -67020
rect -15094 -67132 -15034 -66873
rect -14827 -66873 -14821 -66836
rect -14787 -66836 -14774 -66497
rect -14574 -66497 -14514 -66344
rect -14446 -66398 -14386 -66230
rect -14471 -66404 -14363 -66398
rect -14471 -66438 -14459 -66404
rect -14375 -66438 -14363 -66404
rect -14471 -66444 -14363 -66438
rect -14574 -66530 -14563 -66497
rect -14569 -66834 -14563 -66530
rect -14787 -66873 -14781 -66836
rect -14827 -66885 -14781 -66873
rect -14578 -66873 -14563 -66834
rect -14529 -66530 -14514 -66497
rect -14322 -66497 -14262 -66013
rect -14058 -66013 -14047 -65964
rect -14013 -65964 -14007 -65637
rect -13800 -65637 -13740 -65466
rect -14013 -66013 -13998 -65964
rect -14213 -66072 -14105 -66066
rect -14213 -66106 -14201 -66072
rect -14117 -66106 -14105 -66072
rect -14213 -66112 -14105 -66106
rect -14188 -66170 -14128 -66112
rect -14194 -66230 -14188 -66170
rect -14128 -66230 -14122 -66170
rect -14058 -66284 -13998 -66013
rect -13800 -66013 -13789 -65637
rect -13755 -66013 -13740 -65637
rect -13955 -66072 -13847 -66066
rect -13955 -66106 -13943 -66072
rect -13859 -66106 -13847 -66072
rect -13955 -66112 -13847 -66106
rect -13800 -66228 -13740 -66013
rect -14064 -66344 -14058 -66284
rect -13998 -66344 -13992 -66284
rect -13932 -66288 -13740 -66228
rect -13932 -66398 -13872 -66288
rect -14213 -66404 -14105 -66398
rect -14213 -66438 -14201 -66404
rect -14117 -66438 -14105 -66404
rect -14213 -66444 -14105 -66438
rect -13955 -66404 -13847 -66398
rect -13955 -66438 -13943 -66404
rect -13859 -66438 -13847 -66404
rect -13955 -66444 -13847 -66438
rect -14529 -66834 -14523 -66530
rect -14322 -66542 -14305 -66497
rect -14311 -66820 -14305 -66542
rect -14529 -66873 -14518 -66834
rect -14987 -66932 -14879 -66926
rect -14987 -66966 -14975 -66932
rect -14891 -66966 -14879 -66932
rect -14987 -66972 -14879 -66966
rect -14729 -66932 -14621 -66926
rect -14729 -66966 -14717 -66932
rect -14633 -66966 -14621 -66932
rect -14729 -66972 -14621 -66966
rect -14962 -67020 -14902 -66972
rect -14968 -67080 -14962 -67020
rect -14902 -67080 -14896 -67020
rect -15100 -67192 -15094 -67132
rect -15034 -67192 -15028 -67132
rect -14578 -67280 -14518 -66873
rect -14320 -66873 -14305 -66820
rect -14271 -66542 -14262 -66497
rect -14053 -66497 -14007 -66485
rect -14271 -66820 -14265 -66542
rect -14053 -66796 -14047 -66497
rect -14271 -66873 -14260 -66820
rect -14471 -66932 -14363 -66926
rect -14471 -66966 -14459 -66932
rect -14375 -66966 -14363 -66932
rect -14471 -66972 -14363 -66966
rect -14450 -67026 -14390 -66972
rect -14320 -67240 -14260 -66873
rect -14058 -66873 -14047 -66796
rect -14013 -66796 -14007 -66497
rect -13800 -66497 -13740 -66288
rect -14013 -66873 -13998 -66796
rect -14213 -66932 -14105 -66926
rect -14213 -66966 -14201 -66932
rect -14117 -66966 -14105 -66932
rect -14213 -66972 -14105 -66966
rect -14186 -67020 -14126 -66972
rect -14192 -67080 -14186 -67020
rect -14126 -67080 -14120 -67020
rect -14058 -67132 -13998 -66873
rect -13800 -66873 -13789 -66497
rect -13755 -66873 -13740 -66497
rect -13955 -66932 -13847 -66926
rect -13955 -66966 -13943 -66932
rect -13859 -66966 -13847 -66932
rect -13955 -66972 -13847 -66966
rect -13934 -67018 -13874 -66972
rect -13800 -67018 -13740 -66873
rect -13934 -67078 -13740 -67018
rect -14064 -67192 -14058 -67132
rect -13998 -67192 -13992 -67132
rect -15825 -67299 -15578 -67290
rect -16072 -67330 -15578 -67299
rect -19690 -67430 -17354 -67424
rect -19690 -67530 -19584 -67430
rect -17460 -67530 -17354 -67430
rect -19690 -67536 -17354 -67530
rect -15690 -67424 -15578 -67330
rect -14584 -67340 -14578 -67280
rect -14518 -67340 -14512 -67280
rect -14326 -67300 -14320 -67240
rect -14260 -67300 -14254 -67240
rect -13934 -67424 -13874 -67078
rect -13800 -67424 -13740 -67078
rect -13648 -67132 -13588 -65386
rect -13654 -67192 -13648 -67132
rect -13588 -67192 -13582 -67132
rect -13466 -67290 -13460 -64666
rect -13360 -67290 -13354 -64666
rect -11690 -64426 -9354 -64420
rect -11690 -64526 -11584 -64426
rect -9460 -64526 -9354 -64426
rect -11690 -64532 -9354 -64526
rect -11690 -64666 -11578 -64532
rect -11690 -67234 -11684 -64666
rect -13466 -67424 -13354 -67290
rect -12072 -67265 -11684 -67234
rect -12072 -67299 -12043 -67265
rect -12009 -67299 -11951 -67265
rect -11917 -67299 -11859 -67265
rect -11825 -67290 -11684 -67265
rect -11584 -67290 -11578 -64666
rect -10978 -64832 -10968 -64532
rect -10076 -64832 -10066 -64532
rect -9466 -64666 -9354 -64532
rect -11422 -65036 -9520 -65006
rect -11422 -65100 -11388 -65036
rect -9564 -65100 -9520 -65036
rect -11422 -65130 -9520 -65100
rect -11348 -65394 -11288 -65130
rect -11218 -65394 -11158 -65130
rect -10840 -65274 -10834 -65214
rect -10774 -65274 -10768 -65214
rect -10322 -65274 -10316 -65214
rect -10256 -65274 -10250 -65214
rect -11502 -65506 -11496 -65446
rect -11436 -65506 -11430 -65446
rect -11348 -65454 -11158 -65394
rect -11496 -66040 -11436 -65506
rect -11348 -65637 -11288 -65454
rect -11218 -65538 -11158 -65454
rect -11245 -65544 -11137 -65538
rect -11245 -65578 -11233 -65544
rect -11149 -65578 -11137 -65544
rect -11245 -65584 -11137 -65578
rect -10987 -65544 -10879 -65538
rect -10987 -65578 -10975 -65544
rect -10891 -65578 -10879 -65544
rect -10987 -65584 -10879 -65578
rect -11348 -65670 -11337 -65637
rect -11343 -65970 -11337 -65670
rect -11496 -67020 -11436 -66100
rect -11348 -66013 -11337 -65970
rect -11303 -65670 -11288 -65637
rect -11085 -65637 -11039 -65625
rect -11303 -65970 -11297 -65670
rect -11303 -66013 -11288 -65970
rect -11085 -65988 -11079 -65637
rect -11348 -66236 -11288 -66013
rect -11092 -66013 -11079 -65988
rect -11045 -65988 -11039 -65637
rect -10834 -65637 -10774 -65274
rect -10584 -65386 -10578 -65326
rect -10518 -65386 -10512 -65326
rect -10712 -65506 -10706 -65446
rect -10646 -65506 -10640 -65446
rect -10706 -65538 -10646 -65506
rect -10729 -65544 -10621 -65538
rect -10729 -65578 -10717 -65544
rect -10633 -65578 -10621 -65544
rect -10729 -65584 -10621 -65578
rect -11045 -66013 -11032 -65988
rect -11245 -66072 -11137 -66066
rect -11245 -66106 -11233 -66072
rect -11149 -66106 -11137 -66072
rect -11245 -66112 -11137 -66106
rect -11218 -66236 -11158 -66112
rect -11348 -66296 -11158 -66236
rect -11092 -66284 -11032 -66013
rect -10834 -66013 -10821 -65637
rect -10787 -66013 -10774 -65637
rect -10578 -65637 -10518 -65386
rect -10456 -65506 -10450 -65446
rect -10390 -65506 -10384 -65446
rect -10450 -65538 -10390 -65506
rect -10471 -65544 -10363 -65538
rect -10471 -65578 -10459 -65544
rect -10375 -65578 -10363 -65544
rect -10471 -65584 -10363 -65578
rect -10578 -65670 -10563 -65637
rect -10987 -66072 -10879 -66066
rect -10987 -66106 -10975 -66072
rect -10891 -66106 -10879 -66072
rect -10987 -66112 -10879 -66106
rect -10962 -66170 -10902 -66112
rect -10968 -66230 -10962 -66170
rect -10902 -66230 -10896 -66170
rect -11348 -66497 -11288 -66296
rect -11218 -66398 -11158 -66296
rect -11098 -66344 -11092 -66284
rect -11032 -66344 -11026 -66284
rect -11245 -66404 -11137 -66398
rect -11245 -66438 -11233 -66404
rect -11149 -66438 -11137 -66404
rect -11245 -66444 -11137 -66438
rect -10987 -66404 -10879 -66398
rect -10987 -66438 -10975 -66404
rect -10891 -66438 -10879 -66404
rect -10987 -66444 -10879 -66438
rect -11348 -66550 -11337 -66497
rect -11343 -66873 -11337 -66550
rect -11303 -66550 -11288 -66497
rect -11085 -66497 -11039 -66485
rect -11303 -66873 -11297 -66550
rect -11085 -66828 -11079 -66497
rect -11343 -66885 -11297 -66873
rect -11094 -66873 -11079 -66828
rect -11045 -66828 -11039 -66497
rect -10834 -66497 -10774 -66013
rect -10569 -66013 -10563 -65670
rect -10529 -65670 -10518 -65637
rect -10316 -65637 -10256 -65274
rect -9928 -65406 -9868 -65130
rect -9800 -65406 -9740 -65130
rect -9654 -65386 -9648 -65326
rect -9588 -65386 -9582 -65326
rect -9928 -65466 -9740 -65406
rect -9928 -65538 -9868 -65466
rect -10213 -65544 -10105 -65538
rect -10213 -65578 -10201 -65544
rect -10117 -65578 -10105 -65544
rect -10213 -65584 -10105 -65578
rect -9955 -65544 -9847 -65538
rect -9955 -65578 -9943 -65544
rect -9859 -65578 -9847 -65544
rect -9955 -65584 -9847 -65578
rect -10529 -66013 -10523 -65670
rect -10316 -65698 -10305 -65637
rect -10311 -65956 -10305 -65698
rect -10569 -66025 -10523 -66013
rect -10322 -66013 -10305 -65956
rect -10271 -65698 -10256 -65637
rect -10053 -65637 -10007 -65625
rect -10271 -65956 -10265 -65698
rect -10271 -66013 -10262 -65956
rect -10053 -65964 -10047 -65637
rect -10729 -66072 -10621 -66066
rect -10729 -66106 -10717 -66072
rect -10633 -66106 -10621 -66072
rect -10729 -66112 -10621 -66106
rect -10471 -66072 -10363 -66066
rect -10471 -66106 -10459 -66072
rect -10375 -66106 -10363 -66072
rect -10471 -66112 -10363 -66106
rect -10710 -66230 -10704 -66170
rect -10644 -66230 -10638 -66170
rect -10452 -66230 -10446 -66170
rect -10386 -66230 -10380 -66170
rect -10704 -66398 -10644 -66230
rect -10580 -66344 -10574 -66284
rect -10514 -66344 -10508 -66284
rect -10729 -66404 -10621 -66398
rect -10729 -66438 -10717 -66404
rect -10633 -66438 -10621 -66404
rect -10729 -66444 -10621 -66438
rect -11045 -66873 -11034 -66828
rect -10834 -66836 -10821 -66497
rect -11245 -66932 -11137 -66926
rect -11245 -66966 -11233 -66932
rect -11149 -66966 -11137 -66932
rect -11245 -66972 -11137 -66966
rect -11496 -67080 -11246 -67020
rect -11186 -67080 -11180 -67020
rect -11094 -67132 -11034 -66873
rect -10827 -66873 -10821 -66836
rect -10787 -66836 -10774 -66497
rect -10574 -66497 -10514 -66344
rect -10446 -66398 -10386 -66230
rect -10471 -66404 -10363 -66398
rect -10471 -66438 -10459 -66404
rect -10375 -66438 -10363 -66404
rect -10471 -66444 -10363 -66438
rect -10574 -66530 -10563 -66497
rect -10569 -66834 -10563 -66530
rect -10787 -66873 -10781 -66836
rect -10827 -66885 -10781 -66873
rect -10578 -66873 -10563 -66834
rect -10529 -66530 -10514 -66497
rect -10322 -66497 -10262 -66013
rect -10058 -66013 -10047 -65964
rect -10013 -65964 -10007 -65637
rect -9800 -65637 -9740 -65466
rect -10013 -66013 -9998 -65964
rect -10213 -66072 -10105 -66066
rect -10213 -66106 -10201 -66072
rect -10117 -66106 -10105 -66072
rect -10213 -66112 -10105 -66106
rect -10188 -66170 -10128 -66112
rect -10194 -66230 -10188 -66170
rect -10128 -66230 -10122 -66170
rect -10058 -66284 -9998 -66013
rect -9800 -66013 -9789 -65637
rect -9755 -66013 -9740 -65637
rect -9955 -66072 -9847 -66066
rect -9955 -66106 -9943 -66072
rect -9859 -66106 -9847 -66072
rect -9955 -66112 -9847 -66106
rect -9800 -66228 -9740 -66013
rect -10064 -66344 -10058 -66284
rect -9998 -66344 -9992 -66284
rect -9932 -66288 -9740 -66228
rect -9932 -66398 -9872 -66288
rect -10213 -66404 -10105 -66398
rect -10213 -66438 -10201 -66404
rect -10117 -66438 -10105 -66404
rect -10213 -66444 -10105 -66438
rect -9955 -66404 -9847 -66398
rect -9955 -66438 -9943 -66404
rect -9859 -66438 -9847 -66404
rect -9955 -66444 -9847 -66438
rect -10529 -66834 -10523 -66530
rect -10322 -66542 -10305 -66497
rect -10311 -66820 -10305 -66542
rect -10529 -66873 -10518 -66834
rect -10987 -66932 -10879 -66926
rect -10987 -66966 -10975 -66932
rect -10891 -66966 -10879 -66932
rect -10987 -66972 -10879 -66966
rect -10729 -66932 -10621 -66926
rect -10729 -66966 -10717 -66932
rect -10633 -66966 -10621 -66932
rect -10729 -66972 -10621 -66966
rect -10962 -67020 -10902 -66972
rect -10968 -67080 -10962 -67020
rect -10902 -67080 -10896 -67020
rect -11100 -67192 -11094 -67132
rect -11034 -67192 -11028 -67132
rect -10578 -67280 -10518 -66873
rect -10320 -66873 -10305 -66820
rect -10271 -66542 -10262 -66497
rect -10053 -66497 -10007 -66485
rect -10271 -66820 -10265 -66542
rect -10053 -66796 -10047 -66497
rect -10271 -66873 -10260 -66820
rect -10471 -66932 -10363 -66926
rect -10471 -66966 -10459 -66932
rect -10375 -66966 -10363 -66932
rect -10471 -66972 -10363 -66966
rect -10450 -67026 -10390 -66972
rect -10320 -67240 -10260 -66873
rect -10058 -66873 -10047 -66796
rect -10013 -66796 -10007 -66497
rect -9800 -66497 -9740 -66288
rect -10013 -66873 -9998 -66796
rect -10213 -66932 -10105 -66926
rect -10213 -66966 -10201 -66932
rect -10117 -66966 -10105 -66932
rect -10213 -66972 -10105 -66966
rect -10186 -67020 -10126 -66972
rect -10192 -67080 -10186 -67020
rect -10126 -67080 -10120 -67020
rect -10058 -67132 -9998 -66873
rect -9800 -66873 -9789 -66497
rect -9755 -66873 -9740 -66497
rect -9955 -66932 -9847 -66926
rect -9955 -66966 -9943 -66932
rect -9859 -66966 -9847 -66932
rect -9955 -66972 -9847 -66966
rect -9934 -67018 -9874 -66972
rect -9800 -67018 -9740 -66873
rect -9934 -67078 -9740 -67018
rect -10064 -67192 -10058 -67132
rect -9998 -67192 -9992 -67132
rect -11825 -67299 -11578 -67290
rect -12072 -67330 -11578 -67299
rect -15690 -67430 -13354 -67424
rect -15690 -67530 -15584 -67430
rect -13460 -67530 -13354 -67430
rect -15690 -67536 -13354 -67530
rect -11690 -67424 -11578 -67330
rect -10584 -67340 -10578 -67280
rect -10518 -67340 -10512 -67280
rect -10326 -67300 -10320 -67240
rect -10260 -67300 -10254 -67240
rect -9934 -67424 -9874 -67078
rect -9800 -67424 -9740 -67078
rect -9648 -67132 -9588 -65386
rect -9654 -67192 -9648 -67132
rect -9588 -67192 -9582 -67132
rect -9466 -67290 -9460 -64666
rect -9360 -67290 -9354 -64666
rect -7690 -64426 -5354 -64420
rect -7690 -64526 -7584 -64426
rect -5460 -64526 -5354 -64426
rect -7690 -64532 -5354 -64526
rect -7690 -64666 -7578 -64532
rect -7690 -67234 -7684 -64666
rect -9466 -67424 -9354 -67290
rect -8072 -67265 -7684 -67234
rect -8072 -67299 -8043 -67265
rect -8009 -67299 -7951 -67265
rect -7917 -67299 -7859 -67265
rect -7825 -67290 -7684 -67265
rect -7584 -67290 -7578 -64666
rect -6978 -64832 -6968 -64532
rect -6076 -64832 -6066 -64532
rect -5466 -64666 -5354 -64532
rect -7422 -65036 -5520 -65006
rect -7422 -65100 -7388 -65036
rect -5564 -65100 -5520 -65036
rect -7422 -65130 -5520 -65100
rect -7348 -65394 -7288 -65130
rect -7218 -65394 -7158 -65130
rect -6840 -65274 -6834 -65214
rect -6774 -65274 -6768 -65214
rect -6322 -65274 -6316 -65214
rect -6256 -65274 -6250 -65214
rect -7502 -65506 -7496 -65446
rect -7436 -65506 -7430 -65446
rect -7348 -65454 -7158 -65394
rect -7496 -66040 -7436 -65506
rect -7348 -65637 -7288 -65454
rect -7218 -65538 -7158 -65454
rect -7245 -65544 -7137 -65538
rect -7245 -65578 -7233 -65544
rect -7149 -65578 -7137 -65544
rect -7245 -65584 -7137 -65578
rect -6987 -65544 -6879 -65538
rect -6987 -65578 -6975 -65544
rect -6891 -65578 -6879 -65544
rect -6987 -65584 -6879 -65578
rect -7348 -65670 -7337 -65637
rect -7343 -65970 -7337 -65670
rect -7496 -67020 -7436 -66100
rect -7348 -66013 -7337 -65970
rect -7303 -65670 -7288 -65637
rect -7085 -65637 -7039 -65625
rect -7303 -65970 -7297 -65670
rect -7303 -66013 -7288 -65970
rect -7085 -65988 -7079 -65637
rect -7348 -66236 -7288 -66013
rect -7092 -66013 -7079 -65988
rect -7045 -65988 -7039 -65637
rect -6834 -65637 -6774 -65274
rect -6584 -65386 -6578 -65326
rect -6518 -65386 -6512 -65326
rect -6712 -65506 -6706 -65446
rect -6646 -65506 -6640 -65446
rect -6706 -65538 -6646 -65506
rect -6729 -65544 -6621 -65538
rect -6729 -65578 -6717 -65544
rect -6633 -65578 -6621 -65544
rect -6729 -65584 -6621 -65578
rect -7045 -66013 -7032 -65988
rect -7245 -66072 -7137 -66066
rect -7245 -66106 -7233 -66072
rect -7149 -66106 -7137 -66072
rect -7245 -66112 -7137 -66106
rect -7218 -66236 -7158 -66112
rect -7348 -66296 -7158 -66236
rect -7092 -66284 -7032 -66013
rect -6834 -66013 -6821 -65637
rect -6787 -66013 -6774 -65637
rect -6578 -65637 -6518 -65386
rect -6456 -65506 -6450 -65446
rect -6390 -65506 -6384 -65446
rect -6450 -65538 -6390 -65506
rect -6471 -65544 -6363 -65538
rect -6471 -65578 -6459 -65544
rect -6375 -65578 -6363 -65544
rect -6471 -65584 -6363 -65578
rect -6578 -65670 -6563 -65637
rect -6987 -66072 -6879 -66066
rect -6987 -66106 -6975 -66072
rect -6891 -66106 -6879 -66072
rect -6987 -66112 -6879 -66106
rect -6962 -66170 -6902 -66112
rect -6968 -66230 -6962 -66170
rect -6902 -66230 -6896 -66170
rect -7348 -66497 -7288 -66296
rect -7218 -66398 -7158 -66296
rect -7098 -66344 -7092 -66284
rect -7032 -66344 -7026 -66284
rect -7245 -66404 -7137 -66398
rect -7245 -66438 -7233 -66404
rect -7149 -66438 -7137 -66404
rect -7245 -66444 -7137 -66438
rect -6987 -66404 -6879 -66398
rect -6987 -66438 -6975 -66404
rect -6891 -66438 -6879 -66404
rect -6987 -66444 -6879 -66438
rect -7348 -66550 -7337 -66497
rect -7343 -66873 -7337 -66550
rect -7303 -66550 -7288 -66497
rect -7085 -66497 -7039 -66485
rect -7303 -66873 -7297 -66550
rect -7085 -66828 -7079 -66497
rect -7343 -66885 -7297 -66873
rect -7094 -66873 -7079 -66828
rect -7045 -66828 -7039 -66497
rect -6834 -66497 -6774 -66013
rect -6569 -66013 -6563 -65670
rect -6529 -65670 -6518 -65637
rect -6316 -65637 -6256 -65274
rect -5928 -65406 -5868 -65130
rect -5800 -65406 -5740 -65130
rect -5654 -65386 -5648 -65326
rect -5588 -65386 -5582 -65326
rect -5928 -65466 -5740 -65406
rect -5928 -65538 -5868 -65466
rect -6213 -65544 -6105 -65538
rect -6213 -65578 -6201 -65544
rect -6117 -65578 -6105 -65544
rect -6213 -65584 -6105 -65578
rect -5955 -65544 -5847 -65538
rect -5955 -65578 -5943 -65544
rect -5859 -65578 -5847 -65544
rect -5955 -65584 -5847 -65578
rect -6529 -66013 -6523 -65670
rect -6316 -65698 -6305 -65637
rect -6311 -65956 -6305 -65698
rect -6569 -66025 -6523 -66013
rect -6322 -66013 -6305 -65956
rect -6271 -65698 -6256 -65637
rect -6053 -65637 -6007 -65625
rect -6271 -65956 -6265 -65698
rect -6271 -66013 -6262 -65956
rect -6053 -65964 -6047 -65637
rect -6729 -66072 -6621 -66066
rect -6729 -66106 -6717 -66072
rect -6633 -66106 -6621 -66072
rect -6729 -66112 -6621 -66106
rect -6471 -66072 -6363 -66066
rect -6471 -66106 -6459 -66072
rect -6375 -66106 -6363 -66072
rect -6471 -66112 -6363 -66106
rect -6710 -66230 -6704 -66170
rect -6644 -66230 -6638 -66170
rect -6452 -66230 -6446 -66170
rect -6386 -66230 -6380 -66170
rect -6704 -66398 -6644 -66230
rect -6580 -66344 -6574 -66284
rect -6514 -66344 -6508 -66284
rect -6729 -66404 -6621 -66398
rect -6729 -66438 -6717 -66404
rect -6633 -66438 -6621 -66404
rect -6729 -66444 -6621 -66438
rect -7045 -66873 -7034 -66828
rect -6834 -66836 -6821 -66497
rect -7245 -66932 -7137 -66926
rect -7245 -66966 -7233 -66932
rect -7149 -66966 -7137 -66932
rect -7245 -66972 -7137 -66966
rect -7496 -67080 -7246 -67020
rect -7186 -67080 -7180 -67020
rect -7094 -67132 -7034 -66873
rect -6827 -66873 -6821 -66836
rect -6787 -66836 -6774 -66497
rect -6574 -66497 -6514 -66344
rect -6446 -66398 -6386 -66230
rect -6471 -66404 -6363 -66398
rect -6471 -66438 -6459 -66404
rect -6375 -66438 -6363 -66404
rect -6471 -66444 -6363 -66438
rect -6574 -66530 -6563 -66497
rect -6569 -66834 -6563 -66530
rect -6787 -66873 -6781 -66836
rect -6827 -66885 -6781 -66873
rect -6578 -66873 -6563 -66834
rect -6529 -66530 -6514 -66497
rect -6322 -66497 -6262 -66013
rect -6058 -66013 -6047 -65964
rect -6013 -65964 -6007 -65637
rect -5800 -65637 -5740 -65466
rect -6013 -66013 -5998 -65964
rect -6213 -66072 -6105 -66066
rect -6213 -66106 -6201 -66072
rect -6117 -66106 -6105 -66072
rect -6213 -66112 -6105 -66106
rect -6188 -66170 -6128 -66112
rect -6194 -66230 -6188 -66170
rect -6128 -66230 -6122 -66170
rect -6058 -66284 -5998 -66013
rect -5800 -66013 -5789 -65637
rect -5755 -66013 -5740 -65637
rect -5955 -66072 -5847 -66066
rect -5955 -66106 -5943 -66072
rect -5859 -66106 -5847 -66072
rect -5955 -66112 -5847 -66106
rect -5800 -66228 -5740 -66013
rect -6064 -66344 -6058 -66284
rect -5998 -66344 -5992 -66284
rect -5932 -66288 -5740 -66228
rect -5932 -66398 -5872 -66288
rect -6213 -66404 -6105 -66398
rect -6213 -66438 -6201 -66404
rect -6117 -66438 -6105 -66404
rect -6213 -66444 -6105 -66438
rect -5955 -66404 -5847 -66398
rect -5955 -66438 -5943 -66404
rect -5859 -66438 -5847 -66404
rect -5955 -66444 -5847 -66438
rect -6529 -66834 -6523 -66530
rect -6322 -66542 -6305 -66497
rect -6311 -66820 -6305 -66542
rect -6529 -66873 -6518 -66834
rect -6987 -66932 -6879 -66926
rect -6987 -66966 -6975 -66932
rect -6891 -66966 -6879 -66932
rect -6987 -66972 -6879 -66966
rect -6729 -66932 -6621 -66926
rect -6729 -66966 -6717 -66932
rect -6633 -66966 -6621 -66932
rect -6729 -66972 -6621 -66966
rect -6962 -67020 -6902 -66972
rect -6968 -67080 -6962 -67020
rect -6902 -67080 -6896 -67020
rect -7100 -67192 -7094 -67132
rect -7034 -67192 -7028 -67132
rect -6578 -67280 -6518 -66873
rect -6320 -66873 -6305 -66820
rect -6271 -66542 -6262 -66497
rect -6053 -66497 -6007 -66485
rect -6271 -66820 -6265 -66542
rect -6053 -66796 -6047 -66497
rect -6271 -66873 -6260 -66820
rect -6471 -66932 -6363 -66926
rect -6471 -66966 -6459 -66932
rect -6375 -66966 -6363 -66932
rect -6471 -66972 -6363 -66966
rect -6450 -67026 -6390 -66972
rect -6320 -67240 -6260 -66873
rect -6058 -66873 -6047 -66796
rect -6013 -66796 -6007 -66497
rect -5800 -66497 -5740 -66288
rect -6013 -66873 -5998 -66796
rect -6213 -66932 -6105 -66926
rect -6213 -66966 -6201 -66932
rect -6117 -66966 -6105 -66932
rect -6213 -66972 -6105 -66966
rect -6186 -67020 -6126 -66972
rect -6192 -67080 -6186 -67020
rect -6126 -67080 -6120 -67020
rect -6058 -67132 -5998 -66873
rect -5800 -66873 -5789 -66497
rect -5755 -66873 -5740 -66497
rect -5955 -66932 -5847 -66926
rect -5955 -66966 -5943 -66932
rect -5859 -66966 -5847 -66932
rect -5955 -66972 -5847 -66966
rect -5934 -67018 -5874 -66972
rect -5800 -67018 -5740 -66873
rect -5934 -67078 -5740 -67018
rect -6064 -67192 -6058 -67132
rect -5998 -67192 -5992 -67132
rect -7825 -67299 -7578 -67290
rect -8072 -67330 -7578 -67299
rect -11690 -67430 -9354 -67424
rect -11690 -67530 -11584 -67430
rect -9460 -67530 -9354 -67430
rect -11690 -67536 -9354 -67530
rect -7690 -67424 -7578 -67330
rect -6584 -67340 -6578 -67280
rect -6518 -67340 -6512 -67280
rect -6326 -67300 -6320 -67240
rect -6260 -67300 -6254 -67240
rect -5934 -67424 -5874 -67078
rect -5800 -67424 -5740 -67078
rect -5648 -67132 -5588 -65386
rect -5654 -67192 -5648 -67132
rect -5588 -67192 -5582 -67132
rect -5466 -67290 -5460 -64666
rect -5360 -67290 -5354 -64666
rect -3690 -64426 -1354 -64420
rect -3690 -64526 -3584 -64426
rect -1460 -64526 -1354 -64426
rect -3690 -64532 -1354 -64526
rect -3690 -64666 -3578 -64532
rect -3690 -67234 -3684 -64666
rect -5466 -67424 -5354 -67290
rect -4072 -67265 -3684 -67234
rect -4072 -67299 -4043 -67265
rect -4009 -67299 -3951 -67265
rect -3917 -67299 -3859 -67265
rect -3825 -67290 -3684 -67265
rect -3584 -67290 -3578 -64666
rect -2978 -64832 -2968 -64532
rect -2076 -64832 -2066 -64532
rect -1466 -64666 -1354 -64532
rect -3422 -65036 -1520 -65006
rect -3422 -65100 -3388 -65036
rect -1564 -65100 -1520 -65036
rect -3422 -65130 -1520 -65100
rect -3348 -65394 -3288 -65130
rect -3218 -65394 -3158 -65130
rect -2840 -65274 -2834 -65214
rect -2774 -65274 -2768 -65214
rect -2322 -65274 -2316 -65214
rect -2256 -65274 -2250 -65214
rect -3502 -65506 -3496 -65446
rect -3436 -65506 -3430 -65446
rect -3348 -65454 -3158 -65394
rect -3496 -66040 -3436 -65506
rect -3348 -65637 -3288 -65454
rect -3218 -65538 -3158 -65454
rect -3245 -65544 -3137 -65538
rect -3245 -65578 -3233 -65544
rect -3149 -65578 -3137 -65544
rect -3245 -65584 -3137 -65578
rect -2987 -65544 -2879 -65538
rect -2987 -65578 -2975 -65544
rect -2891 -65578 -2879 -65544
rect -2987 -65584 -2879 -65578
rect -3348 -65670 -3337 -65637
rect -3343 -65970 -3337 -65670
rect -3496 -67020 -3436 -66100
rect -3348 -66013 -3337 -65970
rect -3303 -65670 -3288 -65637
rect -3085 -65637 -3039 -65625
rect -3303 -65970 -3297 -65670
rect -3303 -66013 -3288 -65970
rect -3085 -65988 -3079 -65637
rect -3348 -66236 -3288 -66013
rect -3092 -66013 -3079 -65988
rect -3045 -65988 -3039 -65637
rect -2834 -65637 -2774 -65274
rect -2584 -65386 -2578 -65326
rect -2518 -65386 -2512 -65326
rect -2712 -65506 -2706 -65446
rect -2646 -65506 -2640 -65446
rect -2706 -65538 -2646 -65506
rect -2729 -65544 -2621 -65538
rect -2729 -65578 -2717 -65544
rect -2633 -65578 -2621 -65544
rect -2729 -65584 -2621 -65578
rect -3045 -66013 -3032 -65988
rect -3245 -66072 -3137 -66066
rect -3245 -66106 -3233 -66072
rect -3149 -66106 -3137 -66072
rect -3245 -66112 -3137 -66106
rect -3218 -66236 -3158 -66112
rect -3348 -66296 -3158 -66236
rect -3092 -66284 -3032 -66013
rect -2834 -66013 -2821 -65637
rect -2787 -66013 -2774 -65637
rect -2578 -65637 -2518 -65386
rect -2456 -65506 -2450 -65446
rect -2390 -65506 -2384 -65446
rect -2450 -65538 -2390 -65506
rect -2471 -65544 -2363 -65538
rect -2471 -65578 -2459 -65544
rect -2375 -65578 -2363 -65544
rect -2471 -65584 -2363 -65578
rect -2578 -65670 -2563 -65637
rect -2987 -66072 -2879 -66066
rect -2987 -66106 -2975 -66072
rect -2891 -66106 -2879 -66072
rect -2987 -66112 -2879 -66106
rect -2962 -66170 -2902 -66112
rect -2968 -66230 -2962 -66170
rect -2902 -66230 -2896 -66170
rect -3348 -66497 -3288 -66296
rect -3218 -66398 -3158 -66296
rect -3098 -66344 -3092 -66284
rect -3032 -66344 -3026 -66284
rect -3245 -66404 -3137 -66398
rect -3245 -66438 -3233 -66404
rect -3149 -66438 -3137 -66404
rect -3245 -66444 -3137 -66438
rect -2987 -66404 -2879 -66398
rect -2987 -66438 -2975 -66404
rect -2891 -66438 -2879 -66404
rect -2987 -66444 -2879 -66438
rect -3348 -66550 -3337 -66497
rect -3343 -66873 -3337 -66550
rect -3303 -66550 -3288 -66497
rect -3085 -66497 -3039 -66485
rect -3303 -66873 -3297 -66550
rect -3085 -66828 -3079 -66497
rect -3343 -66885 -3297 -66873
rect -3094 -66873 -3079 -66828
rect -3045 -66828 -3039 -66497
rect -2834 -66497 -2774 -66013
rect -2569 -66013 -2563 -65670
rect -2529 -65670 -2518 -65637
rect -2316 -65637 -2256 -65274
rect -1928 -65406 -1868 -65130
rect -1800 -65406 -1740 -65130
rect -1654 -65386 -1648 -65326
rect -1588 -65386 -1582 -65326
rect -1928 -65466 -1740 -65406
rect -1928 -65538 -1868 -65466
rect -2213 -65544 -2105 -65538
rect -2213 -65578 -2201 -65544
rect -2117 -65578 -2105 -65544
rect -2213 -65584 -2105 -65578
rect -1955 -65544 -1847 -65538
rect -1955 -65578 -1943 -65544
rect -1859 -65578 -1847 -65544
rect -1955 -65584 -1847 -65578
rect -2529 -66013 -2523 -65670
rect -2316 -65698 -2305 -65637
rect -2311 -65956 -2305 -65698
rect -2569 -66025 -2523 -66013
rect -2322 -66013 -2305 -65956
rect -2271 -65698 -2256 -65637
rect -2053 -65637 -2007 -65625
rect -2271 -65956 -2265 -65698
rect -2271 -66013 -2262 -65956
rect -2053 -65964 -2047 -65637
rect -2729 -66072 -2621 -66066
rect -2729 -66106 -2717 -66072
rect -2633 -66106 -2621 -66072
rect -2729 -66112 -2621 -66106
rect -2471 -66072 -2363 -66066
rect -2471 -66106 -2459 -66072
rect -2375 -66106 -2363 -66072
rect -2471 -66112 -2363 -66106
rect -2710 -66230 -2704 -66170
rect -2644 -66230 -2638 -66170
rect -2452 -66230 -2446 -66170
rect -2386 -66230 -2380 -66170
rect -2704 -66398 -2644 -66230
rect -2580 -66344 -2574 -66284
rect -2514 -66344 -2508 -66284
rect -2729 -66404 -2621 -66398
rect -2729 -66438 -2717 -66404
rect -2633 -66438 -2621 -66404
rect -2729 -66444 -2621 -66438
rect -3045 -66873 -3034 -66828
rect -2834 -66836 -2821 -66497
rect -3245 -66932 -3137 -66926
rect -3245 -66966 -3233 -66932
rect -3149 -66966 -3137 -66932
rect -3245 -66972 -3137 -66966
rect -3496 -67080 -3246 -67020
rect -3186 -67080 -3180 -67020
rect -3094 -67132 -3034 -66873
rect -2827 -66873 -2821 -66836
rect -2787 -66836 -2774 -66497
rect -2574 -66497 -2514 -66344
rect -2446 -66398 -2386 -66230
rect -2471 -66404 -2363 -66398
rect -2471 -66438 -2459 -66404
rect -2375 -66438 -2363 -66404
rect -2471 -66444 -2363 -66438
rect -2574 -66530 -2563 -66497
rect -2569 -66834 -2563 -66530
rect -2787 -66873 -2781 -66836
rect -2827 -66885 -2781 -66873
rect -2578 -66873 -2563 -66834
rect -2529 -66530 -2514 -66497
rect -2322 -66497 -2262 -66013
rect -2058 -66013 -2047 -65964
rect -2013 -65964 -2007 -65637
rect -1800 -65637 -1740 -65466
rect -2013 -66013 -1998 -65964
rect -2213 -66072 -2105 -66066
rect -2213 -66106 -2201 -66072
rect -2117 -66106 -2105 -66072
rect -2213 -66112 -2105 -66106
rect -2188 -66170 -2128 -66112
rect -2194 -66230 -2188 -66170
rect -2128 -66230 -2122 -66170
rect -2058 -66284 -1998 -66013
rect -1800 -66013 -1789 -65637
rect -1755 -66013 -1740 -65637
rect -1955 -66072 -1847 -66066
rect -1955 -66106 -1943 -66072
rect -1859 -66106 -1847 -66072
rect -1955 -66112 -1847 -66106
rect -1800 -66228 -1740 -66013
rect -2064 -66344 -2058 -66284
rect -1998 -66344 -1992 -66284
rect -1932 -66288 -1740 -66228
rect -1932 -66398 -1872 -66288
rect -2213 -66404 -2105 -66398
rect -2213 -66438 -2201 -66404
rect -2117 -66438 -2105 -66404
rect -2213 -66444 -2105 -66438
rect -1955 -66404 -1847 -66398
rect -1955 -66438 -1943 -66404
rect -1859 -66438 -1847 -66404
rect -1955 -66444 -1847 -66438
rect -2529 -66834 -2523 -66530
rect -2322 -66542 -2305 -66497
rect -2311 -66820 -2305 -66542
rect -2529 -66873 -2518 -66834
rect -2987 -66932 -2879 -66926
rect -2987 -66966 -2975 -66932
rect -2891 -66966 -2879 -66932
rect -2987 -66972 -2879 -66966
rect -2729 -66932 -2621 -66926
rect -2729 -66966 -2717 -66932
rect -2633 -66966 -2621 -66932
rect -2729 -66972 -2621 -66966
rect -2962 -67020 -2902 -66972
rect -2968 -67080 -2962 -67020
rect -2902 -67080 -2896 -67020
rect -3100 -67192 -3094 -67132
rect -3034 -67192 -3028 -67132
rect -2578 -67280 -2518 -66873
rect -2320 -66873 -2305 -66820
rect -2271 -66542 -2262 -66497
rect -2053 -66497 -2007 -66485
rect -2271 -66820 -2265 -66542
rect -2053 -66796 -2047 -66497
rect -2271 -66873 -2260 -66820
rect -2471 -66932 -2363 -66926
rect -2471 -66966 -2459 -66932
rect -2375 -66966 -2363 -66932
rect -2471 -66972 -2363 -66966
rect -2450 -67026 -2390 -66972
rect -2320 -67240 -2260 -66873
rect -2058 -66873 -2047 -66796
rect -2013 -66796 -2007 -66497
rect -1800 -66497 -1740 -66288
rect -2013 -66873 -1998 -66796
rect -2213 -66932 -2105 -66926
rect -2213 -66966 -2201 -66932
rect -2117 -66966 -2105 -66932
rect -2213 -66972 -2105 -66966
rect -2186 -67020 -2126 -66972
rect -2192 -67080 -2186 -67020
rect -2126 -67080 -2120 -67020
rect -2058 -67132 -1998 -66873
rect -1800 -66873 -1789 -66497
rect -1755 -66873 -1740 -66497
rect -1955 -66932 -1847 -66926
rect -1955 -66966 -1943 -66932
rect -1859 -66966 -1847 -66932
rect -1955 -66972 -1847 -66966
rect -1934 -67018 -1874 -66972
rect -1800 -67018 -1740 -66873
rect -1934 -67078 -1740 -67018
rect -2064 -67192 -2058 -67132
rect -1998 -67192 -1992 -67132
rect -3825 -67299 -3578 -67290
rect -4072 -67330 -3578 -67299
rect -7690 -67430 -5354 -67424
rect -7690 -67530 -7584 -67430
rect -5460 -67530 -5354 -67430
rect -7690 -67536 -5354 -67530
rect -3690 -67424 -3578 -67330
rect -2584 -67340 -2578 -67280
rect -2518 -67340 -2512 -67280
rect -2326 -67300 -2320 -67240
rect -2260 -67300 -2254 -67240
rect -1934 -67424 -1874 -67078
rect -1800 -67424 -1740 -67078
rect -1648 -67132 -1588 -65386
rect -1654 -67192 -1648 -67132
rect -1588 -67192 -1582 -67132
rect -1466 -67290 -1460 -64666
rect -1360 -67290 -1354 -64666
rect 310 -64426 2646 -64420
rect 310 -64526 416 -64426
rect 2540 -64526 2646 -64426
rect 310 -64532 2646 -64526
rect 310 -64666 422 -64532
rect 310 -67234 316 -64666
rect -1466 -67424 -1354 -67290
rect -72 -67265 316 -67234
rect -72 -67299 -43 -67265
rect -9 -67299 49 -67265
rect 83 -67299 141 -67265
rect 175 -67290 316 -67265
rect 416 -67290 422 -64666
rect 1022 -64832 1032 -64532
rect 1924 -64832 1934 -64532
rect 2534 -64666 2646 -64532
rect 578 -65036 2480 -65006
rect 578 -65100 612 -65036
rect 2436 -65100 2480 -65036
rect 578 -65130 2480 -65100
rect 652 -65394 712 -65130
rect 782 -65394 842 -65130
rect 1160 -65274 1166 -65214
rect 1226 -65274 1232 -65214
rect 1678 -65274 1684 -65214
rect 1744 -65274 1750 -65214
rect 498 -65506 504 -65446
rect 564 -65506 570 -65446
rect 652 -65454 842 -65394
rect 504 -66040 564 -65506
rect 652 -65637 712 -65454
rect 782 -65538 842 -65454
rect 755 -65544 863 -65538
rect 755 -65578 767 -65544
rect 851 -65578 863 -65544
rect 755 -65584 863 -65578
rect 1013 -65544 1121 -65538
rect 1013 -65578 1025 -65544
rect 1109 -65578 1121 -65544
rect 1013 -65584 1121 -65578
rect 652 -65670 663 -65637
rect 657 -65970 663 -65670
rect 504 -67020 564 -66100
rect 652 -66013 663 -65970
rect 697 -65670 712 -65637
rect 915 -65637 961 -65625
rect 697 -65970 703 -65670
rect 697 -66013 712 -65970
rect 915 -65988 921 -65637
rect 652 -66236 712 -66013
rect 908 -66013 921 -65988
rect 955 -65988 961 -65637
rect 1166 -65637 1226 -65274
rect 1416 -65386 1422 -65326
rect 1482 -65386 1488 -65326
rect 1288 -65506 1294 -65446
rect 1354 -65506 1360 -65446
rect 1294 -65538 1354 -65506
rect 1271 -65544 1379 -65538
rect 1271 -65578 1283 -65544
rect 1367 -65578 1379 -65544
rect 1271 -65584 1379 -65578
rect 955 -66013 968 -65988
rect 755 -66072 863 -66066
rect 755 -66106 767 -66072
rect 851 -66106 863 -66072
rect 755 -66112 863 -66106
rect 782 -66236 842 -66112
rect 652 -66296 842 -66236
rect 908 -66284 968 -66013
rect 1166 -66013 1179 -65637
rect 1213 -66013 1226 -65637
rect 1422 -65637 1482 -65386
rect 1544 -65506 1550 -65446
rect 1610 -65506 1616 -65446
rect 1550 -65538 1610 -65506
rect 1529 -65544 1637 -65538
rect 1529 -65578 1541 -65544
rect 1625 -65578 1637 -65544
rect 1529 -65584 1637 -65578
rect 1422 -65670 1437 -65637
rect 1013 -66072 1121 -66066
rect 1013 -66106 1025 -66072
rect 1109 -66106 1121 -66072
rect 1013 -66112 1121 -66106
rect 1038 -66170 1098 -66112
rect 1032 -66230 1038 -66170
rect 1098 -66230 1104 -66170
rect 652 -66497 712 -66296
rect 782 -66398 842 -66296
rect 902 -66344 908 -66284
rect 968 -66344 974 -66284
rect 755 -66404 863 -66398
rect 755 -66438 767 -66404
rect 851 -66438 863 -66404
rect 755 -66444 863 -66438
rect 1013 -66404 1121 -66398
rect 1013 -66438 1025 -66404
rect 1109 -66438 1121 -66404
rect 1013 -66444 1121 -66438
rect 652 -66550 663 -66497
rect 657 -66873 663 -66550
rect 697 -66550 712 -66497
rect 915 -66497 961 -66485
rect 697 -66873 703 -66550
rect 915 -66828 921 -66497
rect 657 -66885 703 -66873
rect 906 -66873 921 -66828
rect 955 -66828 961 -66497
rect 1166 -66497 1226 -66013
rect 1431 -66013 1437 -65670
rect 1471 -65670 1482 -65637
rect 1684 -65637 1744 -65274
rect 2072 -65406 2132 -65130
rect 2200 -65406 2260 -65130
rect 2346 -65386 2352 -65326
rect 2412 -65386 2418 -65326
rect 2072 -65466 2260 -65406
rect 2072 -65538 2132 -65466
rect 1787 -65544 1895 -65538
rect 1787 -65578 1799 -65544
rect 1883 -65578 1895 -65544
rect 1787 -65584 1895 -65578
rect 2045 -65544 2153 -65538
rect 2045 -65578 2057 -65544
rect 2141 -65578 2153 -65544
rect 2045 -65584 2153 -65578
rect 1471 -66013 1477 -65670
rect 1684 -65698 1695 -65637
rect 1689 -65956 1695 -65698
rect 1431 -66025 1477 -66013
rect 1678 -66013 1695 -65956
rect 1729 -65698 1744 -65637
rect 1947 -65637 1993 -65625
rect 1729 -65956 1735 -65698
rect 1729 -66013 1738 -65956
rect 1947 -65964 1953 -65637
rect 1271 -66072 1379 -66066
rect 1271 -66106 1283 -66072
rect 1367 -66106 1379 -66072
rect 1271 -66112 1379 -66106
rect 1529 -66072 1637 -66066
rect 1529 -66106 1541 -66072
rect 1625 -66106 1637 -66072
rect 1529 -66112 1637 -66106
rect 1290 -66230 1296 -66170
rect 1356 -66230 1362 -66170
rect 1548 -66230 1554 -66170
rect 1614 -66230 1620 -66170
rect 1296 -66398 1356 -66230
rect 1420 -66344 1426 -66284
rect 1486 -66344 1492 -66284
rect 1271 -66404 1379 -66398
rect 1271 -66438 1283 -66404
rect 1367 -66438 1379 -66404
rect 1271 -66444 1379 -66438
rect 955 -66873 966 -66828
rect 1166 -66836 1179 -66497
rect 755 -66932 863 -66926
rect 755 -66966 767 -66932
rect 851 -66966 863 -66932
rect 755 -66972 863 -66966
rect 504 -67080 754 -67020
rect 814 -67080 820 -67020
rect 906 -67132 966 -66873
rect 1173 -66873 1179 -66836
rect 1213 -66836 1226 -66497
rect 1426 -66497 1486 -66344
rect 1554 -66398 1614 -66230
rect 1529 -66404 1637 -66398
rect 1529 -66438 1541 -66404
rect 1625 -66438 1637 -66404
rect 1529 -66444 1637 -66438
rect 1426 -66530 1437 -66497
rect 1431 -66834 1437 -66530
rect 1213 -66873 1219 -66836
rect 1173 -66885 1219 -66873
rect 1422 -66873 1437 -66834
rect 1471 -66530 1486 -66497
rect 1678 -66497 1738 -66013
rect 1942 -66013 1953 -65964
rect 1987 -65964 1993 -65637
rect 2200 -65637 2260 -65466
rect 1987 -66013 2002 -65964
rect 1787 -66072 1895 -66066
rect 1787 -66106 1799 -66072
rect 1883 -66106 1895 -66072
rect 1787 -66112 1895 -66106
rect 1812 -66170 1872 -66112
rect 1806 -66230 1812 -66170
rect 1872 -66230 1878 -66170
rect 1942 -66284 2002 -66013
rect 2200 -66013 2211 -65637
rect 2245 -66013 2260 -65637
rect 2045 -66072 2153 -66066
rect 2045 -66106 2057 -66072
rect 2141 -66106 2153 -66072
rect 2045 -66112 2153 -66106
rect 2200 -66228 2260 -66013
rect 1936 -66344 1942 -66284
rect 2002 -66344 2008 -66284
rect 2068 -66288 2260 -66228
rect 2068 -66398 2128 -66288
rect 1787 -66404 1895 -66398
rect 1787 -66438 1799 -66404
rect 1883 -66438 1895 -66404
rect 1787 -66444 1895 -66438
rect 2045 -66404 2153 -66398
rect 2045 -66438 2057 -66404
rect 2141 -66438 2153 -66404
rect 2045 -66444 2153 -66438
rect 1471 -66834 1477 -66530
rect 1678 -66542 1695 -66497
rect 1689 -66820 1695 -66542
rect 1471 -66873 1482 -66834
rect 1013 -66932 1121 -66926
rect 1013 -66966 1025 -66932
rect 1109 -66966 1121 -66932
rect 1013 -66972 1121 -66966
rect 1271 -66932 1379 -66926
rect 1271 -66966 1283 -66932
rect 1367 -66966 1379 -66932
rect 1271 -66972 1379 -66966
rect 1038 -67020 1098 -66972
rect 1032 -67080 1038 -67020
rect 1098 -67080 1104 -67020
rect 900 -67192 906 -67132
rect 966 -67192 972 -67132
rect 1422 -67280 1482 -66873
rect 1680 -66873 1695 -66820
rect 1729 -66542 1738 -66497
rect 1947 -66497 1993 -66485
rect 1729 -66820 1735 -66542
rect 1947 -66796 1953 -66497
rect 1729 -66873 1740 -66820
rect 1529 -66932 1637 -66926
rect 1529 -66966 1541 -66932
rect 1625 -66966 1637 -66932
rect 1529 -66972 1637 -66966
rect 1550 -67026 1610 -66972
rect 1680 -67240 1740 -66873
rect 1942 -66873 1953 -66796
rect 1987 -66796 1993 -66497
rect 2200 -66497 2260 -66288
rect 1987 -66873 2002 -66796
rect 1787 -66932 1895 -66926
rect 1787 -66966 1799 -66932
rect 1883 -66966 1895 -66932
rect 1787 -66972 1895 -66966
rect 1814 -67020 1874 -66972
rect 1808 -67080 1814 -67020
rect 1874 -67080 1880 -67020
rect 1942 -67132 2002 -66873
rect 2200 -66873 2211 -66497
rect 2245 -66873 2260 -66497
rect 2045 -66932 2153 -66926
rect 2045 -66966 2057 -66932
rect 2141 -66966 2153 -66932
rect 2045 -66972 2153 -66966
rect 2066 -67018 2126 -66972
rect 2200 -67018 2260 -66873
rect 2066 -67078 2260 -67018
rect 1936 -67192 1942 -67132
rect 2002 -67192 2008 -67132
rect 175 -67299 422 -67290
rect -72 -67330 422 -67299
rect -3690 -67430 -1354 -67424
rect -3690 -67530 -3584 -67430
rect -1460 -67530 -1354 -67430
rect -3690 -67536 -1354 -67530
rect 310 -67424 422 -67330
rect 1416 -67340 1422 -67280
rect 1482 -67340 1488 -67280
rect 1674 -67300 1680 -67240
rect 1740 -67300 1746 -67240
rect 2066 -67424 2126 -67078
rect 2200 -67424 2260 -67078
rect 2352 -67132 2412 -65386
rect 2346 -67192 2352 -67132
rect 2412 -67192 2418 -67132
rect 2534 -67290 2540 -64666
rect 2640 -67290 2646 -64666
rect 4310 -64426 6646 -64420
rect 4310 -64526 4416 -64426
rect 6540 -64526 6646 -64426
rect 4310 -64532 6646 -64526
rect 4310 -64666 4422 -64532
rect 4310 -67234 4316 -64666
rect 2534 -67424 2646 -67290
rect 3928 -67265 4316 -67234
rect 3928 -67299 3957 -67265
rect 3991 -67299 4049 -67265
rect 4083 -67299 4141 -67265
rect 4175 -67290 4316 -67265
rect 4416 -67290 4422 -64666
rect 5022 -64832 5032 -64532
rect 5924 -64832 5934 -64532
rect 6534 -64666 6646 -64532
rect 4578 -65036 6480 -65006
rect 4578 -65100 4612 -65036
rect 6436 -65100 6480 -65036
rect 4578 -65130 6480 -65100
rect 4652 -65394 4712 -65130
rect 4782 -65394 4842 -65130
rect 5160 -65274 5166 -65214
rect 5226 -65274 5232 -65214
rect 5678 -65274 5684 -65214
rect 5744 -65274 5750 -65214
rect 4498 -65506 4504 -65446
rect 4564 -65506 4570 -65446
rect 4652 -65454 4842 -65394
rect 4504 -66040 4564 -65506
rect 4652 -65637 4712 -65454
rect 4782 -65538 4842 -65454
rect 4755 -65544 4863 -65538
rect 4755 -65578 4767 -65544
rect 4851 -65578 4863 -65544
rect 4755 -65584 4863 -65578
rect 5013 -65544 5121 -65538
rect 5013 -65578 5025 -65544
rect 5109 -65578 5121 -65544
rect 5013 -65584 5121 -65578
rect 4652 -65670 4663 -65637
rect 4657 -65970 4663 -65670
rect 4504 -67020 4564 -66100
rect 4652 -66013 4663 -65970
rect 4697 -65670 4712 -65637
rect 4915 -65637 4961 -65625
rect 4697 -65970 4703 -65670
rect 4697 -66013 4712 -65970
rect 4915 -65988 4921 -65637
rect 4652 -66236 4712 -66013
rect 4908 -66013 4921 -65988
rect 4955 -65988 4961 -65637
rect 5166 -65637 5226 -65274
rect 5416 -65386 5422 -65326
rect 5482 -65386 5488 -65326
rect 5288 -65506 5294 -65446
rect 5354 -65506 5360 -65446
rect 5294 -65538 5354 -65506
rect 5271 -65544 5379 -65538
rect 5271 -65578 5283 -65544
rect 5367 -65578 5379 -65544
rect 5271 -65584 5379 -65578
rect 4955 -66013 4968 -65988
rect 4755 -66072 4863 -66066
rect 4755 -66106 4767 -66072
rect 4851 -66106 4863 -66072
rect 4755 -66112 4863 -66106
rect 4782 -66236 4842 -66112
rect 4652 -66296 4842 -66236
rect 4908 -66284 4968 -66013
rect 5166 -66013 5179 -65637
rect 5213 -66013 5226 -65637
rect 5422 -65637 5482 -65386
rect 5544 -65506 5550 -65446
rect 5610 -65506 5616 -65446
rect 5550 -65538 5610 -65506
rect 5529 -65544 5637 -65538
rect 5529 -65578 5541 -65544
rect 5625 -65578 5637 -65544
rect 5529 -65584 5637 -65578
rect 5422 -65670 5437 -65637
rect 5013 -66072 5121 -66066
rect 5013 -66106 5025 -66072
rect 5109 -66106 5121 -66072
rect 5013 -66112 5121 -66106
rect 5038 -66170 5098 -66112
rect 5032 -66230 5038 -66170
rect 5098 -66230 5104 -66170
rect 4652 -66497 4712 -66296
rect 4782 -66398 4842 -66296
rect 4902 -66344 4908 -66284
rect 4968 -66344 4974 -66284
rect 4755 -66404 4863 -66398
rect 4755 -66438 4767 -66404
rect 4851 -66438 4863 -66404
rect 4755 -66444 4863 -66438
rect 5013 -66404 5121 -66398
rect 5013 -66438 5025 -66404
rect 5109 -66438 5121 -66404
rect 5013 -66444 5121 -66438
rect 4652 -66550 4663 -66497
rect 4657 -66873 4663 -66550
rect 4697 -66550 4712 -66497
rect 4915 -66497 4961 -66485
rect 4697 -66873 4703 -66550
rect 4915 -66828 4921 -66497
rect 4657 -66885 4703 -66873
rect 4906 -66873 4921 -66828
rect 4955 -66828 4961 -66497
rect 5166 -66497 5226 -66013
rect 5431 -66013 5437 -65670
rect 5471 -65670 5482 -65637
rect 5684 -65637 5744 -65274
rect 6072 -65406 6132 -65130
rect 6200 -65406 6260 -65130
rect 6346 -65386 6352 -65326
rect 6412 -65386 6418 -65326
rect 6072 -65466 6260 -65406
rect 6072 -65538 6132 -65466
rect 5787 -65544 5895 -65538
rect 5787 -65578 5799 -65544
rect 5883 -65578 5895 -65544
rect 5787 -65584 5895 -65578
rect 6045 -65544 6153 -65538
rect 6045 -65578 6057 -65544
rect 6141 -65578 6153 -65544
rect 6045 -65584 6153 -65578
rect 5471 -66013 5477 -65670
rect 5684 -65698 5695 -65637
rect 5689 -65956 5695 -65698
rect 5431 -66025 5477 -66013
rect 5678 -66013 5695 -65956
rect 5729 -65698 5744 -65637
rect 5947 -65637 5993 -65625
rect 5729 -65956 5735 -65698
rect 5729 -66013 5738 -65956
rect 5947 -65964 5953 -65637
rect 5271 -66072 5379 -66066
rect 5271 -66106 5283 -66072
rect 5367 -66106 5379 -66072
rect 5271 -66112 5379 -66106
rect 5529 -66072 5637 -66066
rect 5529 -66106 5541 -66072
rect 5625 -66106 5637 -66072
rect 5529 -66112 5637 -66106
rect 5290 -66230 5296 -66170
rect 5356 -66230 5362 -66170
rect 5548 -66230 5554 -66170
rect 5614 -66230 5620 -66170
rect 5296 -66398 5356 -66230
rect 5420 -66344 5426 -66284
rect 5486 -66344 5492 -66284
rect 5271 -66404 5379 -66398
rect 5271 -66438 5283 -66404
rect 5367 -66438 5379 -66404
rect 5271 -66444 5379 -66438
rect 4955 -66873 4966 -66828
rect 5166 -66836 5179 -66497
rect 4755 -66932 4863 -66926
rect 4755 -66966 4767 -66932
rect 4851 -66966 4863 -66932
rect 4755 -66972 4863 -66966
rect 4504 -67080 4754 -67020
rect 4814 -67080 4820 -67020
rect 4906 -67132 4966 -66873
rect 5173 -66873 5179 -66836
rect 5213 -66836 5226 -66497
rect 5426 -66497 5486 -66344
rect 5554 -66398 5614 -66230
rect 5529 -66404 5637 -66398
rect 5529 -66438 5541 -66404
rect 5625 -66438 5637 -66404
rect 5529 -66444 5637 -66438
rect 5426 -66530 5437 -66497
rect 5431 -66834 5437 -66530
rect 5213 -66873 5219 -66836
rect 5173 -66885 5219 -66873
rect 5422 -66873 5437 -66834
rect 5471 -66530 5486 -66497
rect 5678 -66497 5738 -66013
rect 5942 -66013 5953 -65964
rect 5987 -65964 5993 -65637
rect 6200 -65637 6260 -65466
rect 5987 -66013 6002 -65964
rect 5787 -66072 5895 -66066
rect 5787 -66106 5799 -66072
rect 5883 -66106 5895 -66072
rect 5787 -66112 5895 -66106
rect 5812 -66170 5872 -66112
rect 5806 -66230 5812 -66170
rect 5872 -66230 5878 -66170
rect 5942 -66284 6002 -66013
rect 6200 -66013 6211 -65637
rect 6245 -66013 6260 -65637
rect 6045 -66072 6153 -66066
rect 6045 -66106 6057 -66072
rect 6141 -66106 6153 -66072
rect 6045 -66112 6153 -66106
rect 6200 -66228 6260 -66013
rect 5936 -66344 5942 -66284
rect 6002 -66344 6008 -66284
rect 6068 -66288 6260 -66228
rect 6068 -66398 6128 -66288
rect 5787 -66404 5895 -66398
rect 5787 -66438 5799 -66404
rect 5883 -66438 5895 -66404
rect 5787 -66444 5895 -66438
rect 6045 -66404 6153 -66398
rect 6045 -66438 6057 -66404
rect 6141 -66438 6153 -66404
rect 6045 -66444 6153 -66438
rect 5471 -66834 5477 -66530
rect 5678 -66542 5695 -66497
rect 5689 -66820 5695 -66542
rect 5471 -66873 5482 -66834
rect 5013 -66932 5121 -66926
rect 5013 -66966 5025 -66932
rect 5109 -66966 5121 -66932
rect 5013 -66972 5121 -66966
rect 5271 -66932 5379 -66926
rect 5271 -66966 5283 -66932
rect 5367 -66966 5379 -66932
rect 5271 -66972 5379 -66966
rect 5038 -67020 5098 -66972
rect 5032 -67080 5038 -67020
rect 5098 -67080 5104 -67020
rect 4900 -67192 4906 -67132
rect 4966 -67192 4972 -67132
rect 5422 -67280 5482 -66873
rect 5680 -66873 5695 -66820
rect 5729 -66542 5738 -66497
rect 5947 -66497 5993 -66485
rect 5729 -66820 5735 -66542
rect 5947 -66796 5953 -66497
rect 5729 -66873 5740 -66820
rect 5529 -66932 5637 -66926
rect 5529 -66966 5541 -66932
rect 5625 -66966 5637 -66932
rect 5529 -66972 5637 -66966
rect 5550 -67026 5610 -66972
rect 5680 -67240 5740 -66873
rect 5942 -66873 5953 -66796
rect 5987 -66796 5993 -66497
rect 6200 -66497 6260 -66288
rect 5987 -66873 6002 -66796
rect 5787 -66932 5895 -66926
rect 5787 -66966 5799 -66932
rect 5883 -66966 5895 -66932
rect 5787 -66972 5895 -66966
rect 5814 -67020 5874 -66972
rect 5808 -67080 5814 -67020
rect 5874 -67080 5880 -67020
rect 5942 -67132 6002 -66873
rect 6200 -66873 6211 -66497
rect 6245 -66873 6260 -66497
rect 6045 -66932 6153 -66926
rect 6045 -66966 6057 -66932
rect 6141 -66966 6153 -66932
rect 6045 -66972 6153 -66966
rect 6066 -67018 6126 -66972
rect 6200 -67018 6260 -66873
rect 6066 -67078 6260 -67018
rect 5936 -67192 5942 -67132
rect 6002 -67192 6008 -67132
rect 4175 -67299 4422 -67290
rect 3928 -67330 4422 -67299
rect 310 -67430 2646 -67424
rect 310 -67530 416 -67430
rect 2540 -67530 2646 -67430
rect 310 -67536 2646 -67530
rect 4310 -67424 4422 -67330
rect 5416 -67340 5422 -67280
rect 5482 -67340 5488 -67280
rect 5674 -67300 5680 -67240
rect 5740 -67300 5746 -67240
rect 6066 -67424 6126 -67078
rect 6200 -67424 6260 -67078
rect 6352 -67132 6412 -65386
rect 6346 -67192 6352 -67132
rect 6412 -67192 6418 -67132
rect 6534 -67290 6540 -64666
rect 6640 -67290 6646 -64666
rect 6534 -67424 6646 -67290
rect 4310 -67430 6646 -67424
rect 4310 -67530 4416 -67430
rect 6540 -67530 6646 -67430
rect 4310 -67536 6646 -67530
rect -28230 -67556 -28170 -67550
rect -24230 -67556 -24170 -67550
rect -20230 -67556 -20170 -67550
rect -16230 -67556 -16170 -67550
rect -12230 -67556 -12170 -67550
rect -8230 -67556 -8170 -67550
rect -4230 -67556 -4170 -67550
rect -230 -67556 -170 -67550
rect 3770 -67556 3830 -67550
rect -28170 -67562 -27944 -67556
rect -28170 -67610 -28004 -67562
rect -27956 -67610 -27944 -67562
rect -28170 -67616 -27944 -67610
rect -27908 -67614 -27848 -67608
rect -28230 -67622 -28170 -67616
rect -27914 -67674 -27908 -67614
rect -27848 -67674 -27842 -67614
rect -24170 -67562 -23944 -67556
rect -24170 -67610 -24004 -67562
rect -23956 -67610 -23944 -67562
rect -24170 -67616 -23944 -67610
rect -23908 -67614 -23848 -67608
rect -24230 -67622 -24170 -67616
rect -23914 -67674 -23908 -67614
rect -23848 -67674 -23842 -67614
rect -20170 -67562 -19944 -67556
rect -20170 -67610 -20004 -67562
rect -19956 -67610 -19944 -67562
rect -20170 -67616 -19944 -67610
rect -19908 -67614 -19848 -67608
rect -20230 -67622 -20170 -67616
rect -19914 -67674 -19908 -67614
rect -19848 -67674 -19842 -67614
rect -16170 -67562 -15944 -67556
rect -16170 -67610 -16004 -67562
rect -15956 -67610 -15944 -67562
rect -16170 -67616 -15944 -67610
rect -15908 -67614 -15848 -67608
rect -16230 -67622 -16170 -67616
rect -15914 -67674 -15908 -67614
rect -15848 -67674 -15842 -67614
rect -12170 -67562 -11944 -67556
rect -12170 -67610 -12004 -67562
rect -11956 -67610 -11944 -67562
rect -12170 -67616 -11944 -67610
rect -11908 -67614 -11848 -67608
rect -12230 -67622 -12170 -67616
rect -11914 -67674 -11908 -67614
rect -11848 -67674 -11842 -67614
rect -8170 -67562 -7944 -67556
rect -8170 -67610 -8004 -67562
rect -7956 -67610 -7944 -67562
rect -8170 -67616 -7944 -67610
rect -7908 -67614 -7848 -67608
rect -8230 -67622 -8170 -67616
rect -7914 -67674 -7908 -67614
rect -7848 -67674 -7842 -67614
rect -4170 -67562 -3944 -67556
rect -4170 -67610 -4004 -67562
rect -3956 -67610 -3944 -67562
rect -4170 -67616 -3944 -67610
rect -3908 -67614 -3848 -67608
rect -4230 -67622 -4170 -67616
rect -3914 -67674 -3908 -67614
rect -3848 -67674 -3842 -67614
rect -170 -67562 56 -67556
rect -170 -67610 -4 -67562
rect 44 -67610 56 -67562
rect -170 -67616 56 -67610
rect 92 -67614 152 -67608
rect -230 -67622 -170 -67616
rect 86 -67674 92 -67614
rect 152 -67674 158 -67614
rect 3830 -67562 4056 -67556
rect 3830 -67610 3996 -67562
rect 4044 -67610 4056 -67562
rect 3830 -67616 4056 -67610
rect 4092 -67614 4152 -67608
rect 3770 -67622 3830 -67616
rect 4086 -67674 4092 -67614
rect 4152 -67674 4158 -67614
rect -27908 -67680 -27848 -67674
rect -23908 -67680 -23848 -67674
rect -19908 -67680 -19848 -67674
rect -15908 -67680 -15848 -67674
rect -11908 -67680 -11848 -67674
rect -7908 -67680 -7848 -67674
rect -3908 -67680 -3848 -67674
rect 92 -67680 152 -67674
rect 4092 -67680 4152 -67674
rect -27690 -67766 -25354 -67760
rect -27690 -67778 -27584 -67766
rect -28072 -67809 -27584 -67778
rect -28072 -67843 -28043 -67809
rect -28009 -67843 -27951 -67809
rect -27917 -67843 -27859 -67809
rect -27825 -67843 -27584 -67809
rect -28072 -67866 -27584 -67843
rect -25460 -67866 -25354 -67766
rect -23690 -67766 -21354 -67760
rect -23690 -67778 -23584 -67766
rect -28072 -67872 -25354 -67866
rect -28072 -67874 -27578 -67872
rect -27690 -67958 -27578 -67874
rect -27690 -69618 -27684 -67958
rect -27584 -69618 -27578 -67958
rect -26578 -67920 -26518 -67914
rect -27100 -68046 -27094 -67986
rect -27034 -68046 -27028 -67986
rect -27250 -68246 -27142 -68240
rect -27250 -68280 -27238 -68246
rect -27154 -68280 -27142 -68246
rect -27250 -68286 -27142 -68280
rect -27348 -68330 -27302 -68318
rect -27348 -68652 -27342 -68330
rect -27356 -68706 -27342 -68652
rect -27308 -68652 -27302 -68330
rect -27094 -68330 -27034 -68046
rect -26846 -68090 -26840 -68030
rect -26780 -68090 -26774 -68030
rect -26992 -68246 -26884 -68240
rect -26992 -68280 -26980 -68246
rect -26896 -68280 -26884 -68246
rect -26992 -68286 -26884 -68280
rect -27094 -68400 -27084 -68330
rect -27308 -68706 -27296 -68652
rect -27090 -68670 -27084 -68400
rect -27356 -68826 -27296 -68706
rect -27100 -68706 -27084 -68670
rect -27050 -68400 -27034 -68330
rect -26840 -68330 -26780 -68090
rect -26714 -68202 -26708 -68142
rect -26648 -68202 -26642 -68142
rect -26708 -68240 -26648 -68202
rect -26734 -68246 -26626 -68240
rect -26734 -68280 -26722 -68246
rect -26638 -68280 -26626 -68246
rect -26734 -68286 -26626 -68280
rect -26840 -68366 -26826 -68330
rect -27050 -68670 -27044 -68400
rect -27050 -68706 -27040 -68670
rect -27250 -68756 -27142 -68750
rect -27250 -68790 -27238 -68756
rect -27154 -68790 -27142 -68756
rect -27250 -68796 -27142 -68790
rect -27226 -68826 -27166 -68796
rect -27356 -68886 -27166 -68826
rect -27356 -69122 -27296 -68886
rect -27226 -69122 -27166 -68886
rect -27100 -68952 -27040 -68706
rect -26832 -68706 -26826 -68366
rect -26792 -68366 -26780 -68330
rect -26578 -68330 -26518 -67980
rect -25466 -67958 -25354 -67872
rect -24072 -67809 -23584 -67778
rect -24072 -67843 -24043 -67809
rect -24009 -67843 -23951 -67809
rect -23917 -67843 -23859 -67809
rect -23825 -67843 -23584 -67809
rect -24072 -67866 -23584 -67843
rect -21460 -67866 -21354 -67766
rect -19690 -67766 -17354 -67760
rect -19690 -67778 -19584 -67766
rect -24072 -67872 -21354 -67866
rect -24072 -67874 -23578 -67872
rect -26326 -68090 -26320 -68030
rect -26260 -68090 -26254 -68030
rect -26458 -68202 -26452 -68142
rect -26392 -68202 -26386 -68142
rect -26452 -68240 -26392 -68202
rect -26476 -68246 -26368 -68240
rect -26476 -68280 -26464 -68246
rect -26380 -68280 -26368 -68246
rect -26476 -68286 -26368 -68280
rect -26578 -68362 -26568 -68330
rect -26792 -68706 -26786 -68366
rect -26832 -68718 -26786 -68706
rect -26574 -68706 -26568 -68362
rect -26534 -68362 -26518 -68330
rect -26320 -68330 -26260 -68090
rect -26218 -68246 -26110 -68240
rect -26218 -68280 -26206 -68246
rect -26122 -68280 -26110 -68246
rect -26218 -68286 -26110 -68280
rect -25960 -68246 -25852 -68240
rect -25960 -68280 -25948 -68246
rect -25864 -68280 -25852 -68246
rect -25960 -68286 -25852 -68280
rect -26534 -68706 -26528 -68362
rect -26320 -68372 -26310 -68330
rect -26574 -68718 -26528 -68706
rect -26316 -68706 -26310 -68372
rect -26276 -68372 -26260 -68330
rect -26058 -68330 -26012 -68318
rect -26276 -68706 -26270 -68372
rect -26058 -68652 -26052 -68330
rect -26316 -68718 -26270 -68706
rect -26064 -68706 -26052 -68652
rect -26018 -68652 -26012 -68330
rect -25800 -68330 -25754 -68318
rect -26018 -68706 -26004 -68652
rect -25800 -68660 -25794 -68330
rect -26992 -68756 -26884 -68750
rect -26992 -68790 -26980 -68756
rect -26896 -68790 -26884 -68756
rect -26992 -68796 -26884 -68790
rect -26734 -68756 -26626 -68750
rect -26734 -68790 -26722 -68756
rect -26638 -68790 -26626 -68756
rect -26734 -68796 -26626 -68790
rect -26476 -68756 -26368 -68750
rect -26476 -68790 -26464 -68756
rect -26380 -68790 -26368 -68756
rect -26476 -68796 -26368 -68790
rect -26218 -68756 -26110 -68750
rect -26218 -68790 -26206 -68756
rect -26122 -68790 -26110 -68756
rect -26218 -68796 -26110 -68790
rect -26966 -68838 -26906 -68796
rect -26192 -68838 -26132 -68796
rect -26972 -68898 -26966 -68838
rect -26906 -68898 -26900 -68838
rect -26198 -68898 -26192 -68838
rect -26132 -68898 -26126 -68838
rect -26064 -68952 -26004 -68706
rect -25808 -68706 -25794 -68660
rect -25760 -68660 -25754 -68330
rect -25760 -68706 -25748 -68660
rect -25960 -68756 -25852 -68750
rect -25960 -68790 -25948 -68756
rect -25864 -68790 -25852 -68756
rect -25960 -68796 -25852 -68790
rect -25936 -68832 -25876 -68796
rect -25808 -68832 -25748 -68706
rect -25936 -68892 -25748 -68832
rect -27106 -69012 -27100 -68952
rect -27040 -69012 -27034 -68952
rect -26070 -69012 -26064 -68952
rect -26004 -69012 -25998 -68952
rect -25936 -69122 -25876 -68892
rect -25808 -69122 -25748 -68892
rect -27466 -69154 -25688 -69122
rect -27466 -69222 -27430 -69154
rect -25722 -69222 -25688 -69154
rect -27466 -69252 -25688 -69222
rect -27690 -69704 -27578 -69618
rect -26978 -69704 -26968 -69404
rect -26076 -69704 -26066 -69404
rect -25466 -69618 -25460 -67958
rect -25360 -69618 -25354 -67958
rect -25466 -69704 -25354 -69618
rect -27690 -69710 -25354 -69704
rect -27690 -69810 -27584 -69710
rect -25460 -69810 -25354 -69710
rect -27690 -69816 -25354 -69810
rect -23690 -67958 -23578 -67874
rect -23690 -69618 -23684 -67958
rect -23584 -69618 -23578 -67958
rect -22578 -67920 -22518 -67914
rect -23100 -68046 -23094 -67986
rect -23034 -68046 -23028 -67986
rect -23250 -68246 -23142 -68240
rect -23250 -68280 -23238 -68246
rect -23154 -68280 -23142 -68246
rect -23250 -68286 -23142 -68280
rect -23348 -68330 -23302 -68318
rect -23348 -68652 -23342 -68330
rect -23356 -68706 -23342 -68652
rect -23308 -68652 -23302 -68330
rect -23094 -68330 -23034 -68046
rect -22846 -68090 -22840 -68030
rect -22780 -68090 -22774 -68030
rect -22992 -68246 -22884 -68240
rect -22992 -68280 -22980 -68246
rect -22896 -68280 -22884 -68246
rect -22992 -68286 -22884 -68280
rect -23094 -68400 -23084 -68330
rect -23308 -68706 -23296 -68652
rect -23090 -68670 -23084 -68400
rect -23356 -68826 -23296 -68706
rect -23100 -68706 -23084 -68670
rect -23050 -68400 -23034 -68330
rect -22840 -68330 -22780 -68090
rect -22714 -68202 -22708 -68142
rect -22648 -68202 -22642 -68142
rect -22708 -68240 -22648 -68202
rect -22734 -68246 -22626 -68240
rect -22734 -68280 -22722 -68246
rect -22638 -68280 -22626 -68246
rect -22734 -68286 -22626 -68280
rect -22840 -68366 -22826 -68330
rect -23050 -68670 -23044 -68400
rect -23050 -68706 -23040 -68670
rect -23250 -68756 -23142 -68750
rect -23250 -68790 -23238 -68756
rect -23154 -68790 -23142 -68756
rect -23250 -68796 -23142 -68790
rect -23226 -68826 -23166 -68796
rect -23356 -68886 -23166 -68826
rect -23356 -69122 -23296 -68886
rect -23226 -69122 -23166 -68886
rect -23100 -68952 -23040 -68706
rect -22832 -68706 -22826 -68366
rect -22792 -68366 -22780 -68330
rect -22578 -68330 -22518 -67980
rect -21466 -67958 -21354 -67872
rect -20072 -67809 -19584 -67778
rect -20072 -67843 -20043 -67809
rect -20009 -67843 -19951 -67809
rect -19917 -67843 -19859 -67809
rect -19825 -67843 -19584 -67809
rect -20072 -67866 -19584 -67843
rect -17460 -67866 -17354 -67766
rect -15690 -67766 -13354 -67760
rect -15690 -67778 -15584 -67766
rect -20072 -67872 -17354 -67866
rect -20072 -67874 -19578 -67872
rect -22326 -68090 -22320 -68030
rect -22260 -68090 -22254 -68030
rect -22458 -68202 -22452 -68142
rect -22392 -68202 -22386 -68142
rect -22452 -68240 -22392 -68202
rect -22476 -68246 -22368 -68240
rect -22476 -68280 -22464 -68246
rect -22380 -68280 -22368 -68246
rect -22476 -68286 -22368 -68280
rect -22578 -68362 -22568 -68330
rect -22792 -68706 -22786 -68366
rect -22832 -68718 -22786 -68706
rect -22574 -68706 -22568 -68362
rect -22534 -68362 -22518 -68330
rect -22320 -68330 -22260 -68090
rect -22218 -68246 -22110 -68240
rect -22218 -68280 -22206 -68246
rect -22122 -68280 -22110 -68246
rect -22218 -68286 -22110 -68280
rect -21960 -68246 -21852 -68240
rect -21960 -68280 -21948 -68246
rect -21864 -68280 -21852 -68246
rect -21960 -68286 -21852 -68280
rect -22534 -68706 -22528 -68362
rect -22320 -68372 -22310 -68330
rect -22574 -68718 -22528 -68706
rect -22316 -68706 -22310 -68372
rect -22276 -68372 -22260 -68330
rect -22058 -68330 -22012 -68318
rect -22276 -68706 -22270 -68372
rect -22058 -68652 -22052 -68330
rect -22316 -68718 -22270 -68706
rect -22064 -68706 -22052 -68652
rect -22018 -68652 -22012 -68330
rect -21800 -68330 -21754 -68318
rect -22018 -68706 -22004 -68652
rect -21800 -68660 -21794 -68330
rect -22992 -68756 -22884 -68750
rect -22992 -68790 -22980 -68756
rect -22896 -68790 -22884 -68756
rect -22992 -68796 -22884 -68790
rect -22734 -68756 -22626 -68750
rect -22734 -68790 -22722 -68756
rect -22638 -68790 -22626 -68756
rect -22734 -68796 -22626 -68790
rect -22476 -68756 -22368 -68750
rect -22476 -68790 -22464 -68756
rect -22380 -68790 -22368 -68756
rect -22476 -68796 -22368 -68790
rect -22218 -68756 -22110 -68750
rect -22218 -68790 -22206 -68756
rect -22122 -68790 -22110 -68756
rect -22218 -68796 -22110 -68790
rect -22966 -68838 -22906 -68796
rect -22192 -68838 -22132 -68796
rect -22972 -68898 -22966 -68838
rect -22906 -68898 -22900 -68838
rect -22198 -68898 -22192 -68838
rect -22132 -68898 -22126 -68838
rect -22064 -68952 -22004 -68706
rect -21808 -68706 -21794 -68660
rect -21760 -68660 -21754 -68330
rect -21760 -68706 -21748 -68660
rect -21960 -68756 -21852 -68750
rect -21960 -68790 -21948 -68756
rect -21864 -68790 -21852 -68756
rect -21960 -68796 -21852 -68790
rect -21936 -68832 -21876 -68796
rect -21808 -68832 -21748 -68706
rect -21936 -68892 -21748 -68832
rect -23106 -69012 -23100 -68952
rect -23040 -69012 -23034 -68952
rect -22070 -69012 -22064 -68952
rect -22004 -69012 -21998 -68952
rect -21936 -69122 -21876 -68892
rect -21808 -69122 -21748 -68892
rect -23466 -69154 -21688 -69122
rect -23466 -69222 -23430 -69154
rect -21722 -69222 -21688 -69154
rect -23466 -69252 -21688 -69222
rect -23690 -69704 -23578 -69618
rect -22978 -69704 -22968 -69404
rect -22076 -69704 -22066 -69404
rect -21466 -69618 -21460 -67958
rect -21360 -69618 -21354 -67958
rect -21466 -69704 -21354 -69618
rect -23690 -69710 -21354 -69704
rect -23690 -69810 -23584 -69710
rect -21460 -69810 -21354 -69710
rect -23690 -69816 -21354 -69810
rect -19690 -67958 -19578 -67874
rect -19690 -69618 -19684 -67958
rect -19584 -69618 -19578 -67958
rect -18578 -67920 -18518 -67914
rect -19100 -68046 -19094 -67986
rect -19034 -68046 -19028 -67986
rect -19250 -68246 -19142 -68240
rect -19250 -68280 -19238 -68246
rect -19154 -68280 -19142 -68246
rect -19250 -68286 -19142 -68280
rect -19348 -68330 -19302 -68318
rect -19348 -68652 -19342 -68330
rect -19356 -68706 -19342 -68652
rect -19308 -68652 -19302 -68330
rect -19094 -68330 -19034 -68046
rect -18846 -68090 -18840 -68030
rect -18780 -68090 -18774 -68030
rect -18992 -68246 -18884 -68240
rect -18992 -68280 -18980 -68246
rect -18896 -68280 -18884 -68246
rect -18992 -68286 -18884 -68280
rect -19094 -68400 -19084 -68330
rect -19308 -68706 -19296 -68652
rect -19090 -68670 -19084 -68400
rect -19356 -68826 -19296 -68706
rect -19100 -68706 -19084 -68670
rect -19050 -68400 -19034 -68330
rect -18840 -68330 -18780 -68090
rect -18714 -68202 -18708 -68142
rect -18648 -68202 -18642 -68142
rect -18708 -68240 -18648 -68202
rect -18734 -68246 -18626 -68240
rect -18734 -68280 -18722 -68246
rect -18638 -68280 -18626 -68246
rect -18734 -68286 -18626 -68280
rect -18840 -68366 -18826 -68330
rect -19050 -68670 -19044 -68400
rect -19050 -68706 -19040 -68670
rect -19250 -68756 -19142 -68750
rect -19250 -68790 -19238 -68756
rect -19154 -68790 -19142 -68756
rect -19250 -68796 -19142 -68790
rect -19226 -68826 -19166 -68796
rect -19356 -68886 -19166 -68826
rect -19356 -69122 -19296 -68886
rect -19226 -69122 -19166 -68886
rect -19100 -68952 -19040 -68706
rect -18832 -68706 -18826 -68366
rect -18792 -68366 -18780 -68330
rect -18578 -68330 -18518 -67980
rect -17466 -67958 -17354 -67872
rect -16072 -67809 -15584 -67778
rect -16072 -67843 -16043 -67809
rect -16009 -67843 -15951 -67809
rect -15917 -67843 -15859 -67809
rect -15825 -67843 -15584 -67809
rect -16072 -67866 -15584 -67843
rect -13460 -67866 -13354 -67766
rect -11690 -67766 -9354 -67760
rect -11690 -67778 -11584 -67766
rect -16072 -67872 -13354 -67866
rect -16072 -67874 -15578 -67872
rect -18326 -68090 -18320 -68030
rect -18260 -68090 -18254 -68030
rect -18458 -68202 -18452 -68142
rect -18392 -68202 -18386 -68142
rect -18452 -68240 -18392 -68202
rect -18476 -68246 -18368 -68240
rect -18476 -68280 -18464 -68246
rect -18380 -68280 -18368 -68246
rect -18476 -68286 -18368 -68280
rect -18578 -68362 -18568 -68330
rect -18792 -68706 -18786 -68366
rect -18832 -68718 -18786 -68706
rect -18574 -68706 -18568 -68362
rect -18534 -68362 -18518 -68330
rect -18320 -68330 -18260 -68090
rect -18218 -68246 -18110 -68240
rect -18218 -68280 -18206 -68246
rect -18122 -68280 -18110 -68246
rect -18218 -68286 -18110 -68280
rect -17960 -68246 -17852 -68240
rect -17960 -68280 -17948 -68246
rect -17864 -68280 -17852 -68246
rect -17960 -68286 -17852 -68280
rect -18534 -68706 -18528 -68362
rect -18320 -68372 -18310 -68330
rect -18574 -68718 -18528 -68706
rect -18316 -68706 -18310 -68372
rect -18276 -68372 -18260 -68330
rect -18058 -68330 -18012 -68318
rect -18276 -68706 -18270 -68372
rect -18058 -68652 -18052 -68330
rect -18316 -68718 -18270 -68706
rect -18064 -68706 -18052 -68652
rect -18018 -68652 -18012 -68330
rect -17800 -68330 -17754 -68318
rect -18018 -68706 -18004 -68652
rect -17800 -68660 -17794 -68330
rect -18992 -68756 -18884 -68750
rect -18992 -68790 -18980 -68756
rect -18896 -68790 -18884 -68756
rect -18992 -68796 -18884 -68790
rect -18734 -68756 -18626 -68750
rect -18734 -68790 -18722 -68756
rect -18638 -68790 -18626 -68756
rect -18734 -68796 -18626 -68790
rect -18476 -68756 -18368 -68750
rect -18476 -68790 -18464 -68756
rect -18380 -68790 -18368 -68756
rect -18476 -68796 -18368 -68790
rect -18218 -68756 -18110 -68750
rect -18218 -68790 -18206 -68756
rect -18122 -68790 -18110 -68756
rect -18218 -68796 -18110 -68790
rect -18966 -68838 -18906 -68796
rect -18192 -68838 -18132 -68796
rect -18972 -68898 -18966 -68838
rect -18906 -68898 -18900 -68838
rect -18198 -68898 -18192 -68838
rect -18132 -68898 -18126 -68838
rect -18064 -68952 -18004 -68706
rect -17808 -68706 -17794 -68660
rect -17760 -68660 -17754 -68330
rect -17760 -68706 -17748 -68660
rect -17960 -68756 -17852 -68750
rect -17960 -68790 -17948 -68756
rect -17864 -68790 -17852 -68756
rect -17960 -68796 -17852 -68790
rect -17936 -68832 -17876 -68796
rect -17808 -68832 -17748 -68706
rect -17936 -68892 -17748 -68832
rect -19106 -69012 -19100 -68952
rect -19040 -69012 -19034 -68952
rect -18070 -69012 -18064 -68952
rect -18004 -69012 -17998 -68952
rect -17936 -69122 -17876 -68892
rect -17808 -69122 -17748 -68892
rect -19466 -69154 -17688 -69122
rect -19466 -69222 -19430 -69154
rect -17722 -69222 -17688 -69154
rect -19466 -69252 -17688 -69222
rect -19690 -69704 -19578 -69618
rect -18978 -69704 -18968 -69404
rect -18076 -69704 -18066 -69404
rect -17466 -69618 -17460 -67958
rect -17360 -69618 -17354 -67958
rect -17466 -69704 -17354 -69618
rect -19690 -69710 -17354 -69704
rect -19690 -69810 -19584 -69710
rect -17460 -69810 -17354 -69710
rect -19690 -69816 -17354 -69810
rect -15690 -67958 -15578 -67874
rect -15690 -69618 -15684 -67958
rect -15584 -69618 -15578 -67958
rect -14578 -67920 -14518 -67914
rect -15100 -68046 -15094 -67986
rect -15034 -68046 -15028 -67986
rect -15250 -68246 -15142 -68240
rect -15250 -68280 -15238 -68246
rect -15154 -68280 -15142 -68246
rect -15250 -68286 -15142 -68280
rect -15348 -68330 -15302 -68318
rect -15348 -68652 -15342 -68330
rect -15356 -68706 -15342 -68652
rect -15308 -68652 -15302 -68330
rect -15094 -68330 -15034 -68046
rect -14846 -68090 -14840 -68030
rect -14780 -68090 -14774 -68030
rect -14992 -68246 -14884 -68240
rect -14992 -68280 -14980 -68246
rect -14896 -68280 -14884 -68246
rect -14992 -68286 -14884 -68280
rect -15094 -68400 -15084 -68330
rect -15308 -68706 -15296 -68652
rect -15090 -68670 -15084 -68400
rect -15356 -68826 -15296 -68706
rect -15100 -68706 -15084 -68670
rect -15050 -68400 -15034 -68330
rect -14840 -68330 -14780 -68090
rect -14714 -68202 -14708 -68142
rect -14648 -68202 -14642 -68142
rect -14708 -68240 -14648 -68202
rect -14734 -68246 -14626 -68240
rect -14734 -68280 -14722 -68246
rect -14638 -68280 -14626 -68246
rect -14734 -68286 -14626 -68280
rect -14840 -68366 -14826 -68330
rect -15050 -68670 -15044 -68400
rect -15050 -68706 -15040 -68670
rect -15250 -68756 -15142 -68750
rect -15250 -68790 -15238 -68756
rect -15154 -68790 -15142 -68756
rect -15250 -68796 -15142 -68790
rect -15226 -68826 -15166 -68796
rect -15356 -68886 -15166 -68826
rect -15356 -69122 -15296 -68886
rect -15226 -69122 -15166 -68886
rect -15100 -68952 -15040 -68706
rect -14832 -68706 -14826 -68366
rect -14792 -68366 -14780 -68330
rect -14578 -68330 -14518 -67980
rect -13466 -67958 -13354 -67872
rect -12072 -67809 -11584 -67778
rect -12072 -67843 -12043 -67809
rect -12009 -67843 -11951 -67809
rect -11917 -67843 -11859 -67809
rect -11825 -67843 -11584 -67809
rect -12072 -67866 -11584 -67843
rect -9460 -67866 -9354 -67766
rect -7690 -67766 -5354 -67760
rect -7690 -67778 -7584 -67766
rect -12072 -67872 -9354 -67866
rect -12072 -67874 -11578 -67872
rect -14326 -68090 -14320 -68030
rect -14260 -68090 -14254 -68030
rect -14458 -68202 -14452 -68142
rect -14392 -68202 -14386 -68142
rect -14452 -68240 -14392 -68202
rect -14476 -68246 -14368 -68240
rect -14476 -68280 -14464 -68246
rect -14380 -68280 -14368 -68246
rect -14476 -68286 -14368 -68280
rect -14578 -68362 -14568 -68330
rect -14792 -68706 -14786 -68366
rect -14832 -68718 -14786 -68706
rect -14574 -68706 -14568 -68362
rect -14534 -68362 -14518 -68330
rect -14320 -68330 -14260 -68090
rect -14218 -68246 -14110 -68240
rect -14218 -68280 -14206 -68246
rect -14122 -68280 -14110 -68246
rect -14218 -68286 -14110 -68280
rect -13960 -68246 -13852 -68240
rect -13960 -68280 -13948 -68246
rect -13864 -68280 -13852 -68246
rect -13960 -68286 -13852 -68280
rect -14534 -68706 -14528 -68362
rect -14320 -68372 -14310 -68330
rect -14574 -68718 -14528 -68706
rect -14316 -68706 -14310 -68372
rect -14276 -68372 -14260 -68330
rect -14058 -68330 -14012 -68318
rect -14276 -68706 -14270 -68372
rect -14058 -68652 -14052 -68330
rect -14316 -68718 -14270 -68706
rect -14064 -68706 -14052 -68652
rect -14018 -68652 -14012 -68330
rect -13800 -68330 -13754 -68318
rect -14018 -68706 -14004 -68652
rect -13800 -68660 -13794 -68330
rect -14992 -68756 -14884 -68750
rect -14992 -68790 -14980 -68756
rect -14896 -68790 -14884 -68756
rect -14992 -68796 -14884 -68790
rect -14734 -68756 -14626 -68750
rect -14734 -68790 -14722 -68756
rect -14638 -68790 -14626 -68756
rect -14734 -68796 -14626 -68790
rect -14476 -68756 -14368 -68750
rect -14476 -68790 -14464 -68756
rect -14380 -68790 -14368 -68756
rect -14476 -68796 -14368 -68790
rect -14218 -68756 -14110 -68750
rect -14218 -68790 -14206 -68756
rect -14122 -68790 -14110 -68756
rect -14218 -68796 -14110 -68790
rect -14966 -68838 -14906 -68796
rect -14192 -68838 -14132 -68796
rect -14972 -68898 -14966 -68838
rect -14906 -68898 -14900 -68838
rect -14198 -68898 -14192 -68838
rect -14132 -68898 -14126 -68838
rect -14064 -68952 -14004 -68706
rect -13808 -68706 -13794 -68660
rect -13760 -68660 -13754 -68330
rect -13760 -68706 -13748 -68660
rect -13960 -68756 -13852 -68750
rect -13960 -68790 -13948 -68756
rect -13864 -68790 -13852 -68756
rect -13960 -68796 -13852 -68790
rect -13936 -68832 -13876 -68796
rect -13808 -68832 -13748 -68706
rect -13936 -68892 -13748 -68832
rect -15106 -69012 -15100 -68952
rect -15040 -69012 -15034 -68952
rect -14070 -69012 -14064 -68952
rect -14004 -69012 -13998 -68952
rect -13936 -69122 -13876 -68892
rect -13808 -69122 -13748 -68892
rect -15466 -69154 -13688 -69122
rect -15466 -69222 -15430 -69154
rect -13722 -69222 -13688 -69154
rect -15466 -69252 -13688 -69222
rect -15690 -69704 -15578 -69618
rect -14978 -69704 -14968 -69404
rect -14076 -69704 -14066 -69404
rect -13466 -69618 -13460 -67958
rect -13360 -69618 -13354 -67958
rect -13466 -69704 -13354 -69618
rect -15690 -69710 -13354 -69704
rect -15690 -69810 -15584 -69710
rect -13460 -69810 -13354 -69710
rect -15690 -69816 -13354 -69810
rect -11690 -67958 -11578 -67874
rect -11690 -69618 -11684 -67958
rect -11584 -69618 -11578 -67958
rect -10578 -67920 -10518 -67914
rect -11100 -68046 -11094 -67986
rect -11034 -68046 -11028 -67986
rect -11250 -68246 -11142 -68240
rect -11250 -68280 -11238 -68246
rect -11154 -68280 -11142 -68246
rect -11250 -68286 -11142 -68280
rect -11348 -68330 -11302 -68318
rect -11348 -68652 -11342 -68330
rect -11356 -68706 -11342 -68652
rect -11308 -68652 -11302 -68330
rect -11094 -68330 -11034 -68046
rect -10846 -68090 -10840 -68030
rect -10780 -68090 -10774 -68030
rect -10992 -68246 -10884 -68240
rect -10992 -68280 -10980 -68246
rect -10896 -68280 -10884 -68246
rect -10992 -68286 -10884 -68280
rect -11094 -68400 -11084 -68330
rect -11308 -68706 -11296 -68652
rect -11090 -68670 -11084 -68400
rect -11356 -68826 -11296 -68706
rect -11100 -68706 -11084 -68670
rect -11050 -68400 -11034 -68330
rect -10840 -68330 -10780 -68090
rect -10714 -68202 -10708 -68142
rect -10648 -68202 -10642 -68142
rect -10708 -68240 -10648 -68202
rect -10734 -68246 -10626 -68240
rect -10734 -68280 -10722 -68246
rect -10638 -68280 -10626 -68246
rect -10734 -68286 -10626 -68280
rect -10840 -68366 -10826 -68330
rect -11050 -68670 -11044 -68400
rect -11050 -68706 -11040 -68670
rect -11250 -68756 -11142 -68750
rect -11250 -68790 -11238 -68756
rect -11154 -68790 -11142 -68756
rect -11250 -68796 -11142 -68790
rect -11226 -68826 -11166 -68796
rect -11356 -68886 -11166 -68826
rect -11356 -69122 -11296 -68886
rect -11226 -69122 -11166 -68886
rect -11100 -68952 -11040 -68706
rect -10832 -68706 -10826 -68366
rect -10792 -68366 -10780 -68330
rect -10578 -68330 -10518 -67980
rect -9466 -67958 -9354 -67872
rect -8072 -67809 -7584 -67778
rect -8072 -67843 -8043 -67809
rect -8009 -67843 -7951 -67809
rect -7917 -67843 -7859 -67809
rect -7825 -67843 -7584 -67809
rect -8072 -67866 -7584 -67843
rect -5460 -67866 -5354 -67766
rect -3690 -67766 -1354 -67760
rect -3690 -67778 -3584 -67766
rect -8072 -67872 -5354 -67866
rect -8072 -67874 -7578 -67872
rect -10326 -68090 -10320 -68030
rect -10260 -68090 -10254 -68030
rect -10458 -68202 -10452 -68142
rect -10392 -68202 -10386 -68142
rect -10452 -68240 -10392 -68202
rect -10476 -68246 -10368 -68240
rect -10476 -68280 -10464 -68246
rect -10380 -68280 -10368 -68246
rect -10476 -68286 -10368 -68280
rect -10578 -68362 -10568 -68330
rect -10792 -68706 -10786 -68366
rect -10832 -68718 -10786 -68706
rect -10574 -68706 -10568 -68362
rect -10534 -68362 -10518 -68330
rect -10320 -68330 -10260 -68090
rect -10218 -68246 -10110 -68240
rect -10218 -68280 -10206 -68246
rect -10122 -68280 -10110 -68246
rect -10218 -68286 -10110 -68280
rect -9960 -68246 -9852 -68240
rect -9960 -68280 -9948 -68246
rect -9864 -68280 -9852 -68246
rect -9960 -68286 -9852 -68280
rect -10534 -68706 -10528 -68362
rect -10320 -68372 -10310 -68330
rect -10574 -68718 -10528 -68706
rect -10316 -68706 -10310 -68372
rect -10276 -68372 -10260 -68330
rect -10058 -68330 -10012 -68318
rect -10276 -68706 -10270 -68372
rect -10058 -68652 -10052 -68330
rect -10316 -68718 -10270 -68706
rect -10064 -68706 -10052 -68652
rect -10018 -68652 -10012 -68330
rect -9800 -68330 -9754 -68318
rect -10018 -68706 -10004 -68652
rect -9800 -68660 -9794 -68330
rect -10992 -68756 -10884 -68750
rect -10992 -68790 -10980 -68756
rect -10896 -68790 -10884 -68756
rect -10992 -68796 -10884 -68790
rect -10734 -68756 -10626 -68750
rect -10734 -68790 -10722 -68756
rect -10638 -68790 -10626 -68756
rect -10734 -68796 -10626 -68790
rect -10476 -68756 -10368 -68750
rect -10476 -68790 -10464 -68756
rect -10380 -68790 -10368 -68756
rect -10476 -68796 -10368 -68790
rect -10218 -68756 -10110 -68750
rect -10218 -68790 -10206 -68756
rect -10122 -68790 -10110 -68756
rect -10218 -68796 -10110 -68790
rect -10966 -68838 -10906 -68796
rect -10192 -68838 -10132 -68796
rect -10972 -68898 -10966 -68838
rect -10906 -68898 -10900 -68838
rect -10198 -68898 -10192 -68838
rect -10132 -68898 -10126 -68838
rect -10064 -68952 -10004 -68706
rect -9808 -68706 -9794 -68660
rect -9760 -68660 -9754 -68330
rect -9760 -68706 -9748 -68660
rect -9960 -68756 -9852 -68750
rect -9960 -68790 -9948 -68756
rect -9864 -68790 -9852 -68756
rect -9960 -68796 -9852 -68790
rect -9936 -68832 -9876 -68796
rect -9808 -68832 -9748 -68706
rect -9936 -68892 -9748 -68832
rect -11106 -69012 -11100 -68952
rect -11040 -69012 -11034 -68952
rect -10070 -69012 -10064 -68952
rect -10004 -69012 -9998 -68952
rect -9936 -69122 -9876 -68892
rect -9808 -69122 -9748 -68892
rect -11466 -69154 -9688 -69122
rect -11466 -69222 -11430 -69154
rect -9722 -69222 -9688 -69154
rect -11466 -69252 -9688 -69222
rect -11690 -69704 -11578 -69618
rect -10978 -69704 -10968 -69404
rect -10076 -69704 -10066 -69404
rect -9466 -69618 -9460 -67958
rect -9360 -69618 -9354 -67958
rect -9466 -69704 -9354 -69618
rect -11690 -69710 -9354 -69704
rect -11690 -69810 -11584 -69710
rect -9460 -69810 -9354 -69710
rect -11690 -69816 -9354 -69810
rect -7690 -67958 -7578 -67874
rect -7690 -69618 -7684 -67958
rect -7584 -69618 -7578 -67958
rect -6578 -67920 -6518 -67914
rect -7100 -68046 -7094 -67986
rect -7034 -68046 -7028 -67986
rect -7250 -68246 -7142 -68240
rect -7250 -68280 -7238 -68246
rect -7154 -68280 -7142 -68246
rect -7250 -68286 -7142 -68280
rect -7348 -68330 -7302 -68318
rect -7348 -68652 -7342 -68330
rect -7356 -68706 -7342 -68652
rect -7308 -68652 -7302 -68330
rect -7094 -68330 -7034 -68046
rect -6846 -68090 -6840 -68030
rect -6780 -68090 -6774 -68030
rect -6992 -68246 -6884 -68240
rect -6992 -68280 -6980 -68246
rect -6896 -68280 -6884 -68246
rect -6992 -68286 -6884 -68280
rect -7094 -68400 -7084 -68330
rect -7308 -68706 -7296 -68652
rect -7090 -68670 -7084 -68400
rect -7356 -68826 -7296 -68706
rect -7100 -68706 -7084 -68670
rect -7050 -68400 -7034 -68330
rect -6840 -68330 -6780 -68090
rect -6714 -68202 -6708 -68142
rect -6648 -68202 -6642 -68142
rect -6708 -68240 -6648 -68202
rect -6734 -68246 -6626 -68240
rect -6734 -68280 -6722 -68246
rect -6638 -68280 -6626 -68246
rect -6734 -68286 -6626 -68280
rect -6840 -68366 -6826 -68330
rect -7050 -68670 -7044 -68400
rect -7050 -68706 -7040 -68670
rect -7250 -68756 -7142 -68750
rect -7250 -68790 -7238 -68756
rect -7154 -68790 -7142 -68756
rect -7250 -68796 -7142 -68790
rect -7226 -68826 -7166 -68796
rect -7356 -68886 -7166 -68826
rect -7356 -69122 -7296 -68886
rect -7226 -69122 -7166 -68886
rect -7100 -68952 -7040 -68706
rect -6832 -68706 -6826 -68366
rect -6792 -68366 -6780 -68330
rect -6578 -68330 -6518 -67980
rect -5466 -67958 -5354 -67872
rect -4072 -67809 -3584 -67778
rect -4072 -67843 -4043 -67809
rect -4009 -67843 -3951 -67809
rect -3917 -67843 -3859 -67809
rect -3825 -67843 -3584 -67809
rect -4072 -67866 -3584 -67843
rect -1460 -67866 -1354 -67766
rect 310 -67766 2646 -67760
rect 310 -67778 416 -67766
rect -4072 -67872 -1354 -67866
rect -4072 -67874 -3578 -67872
rect -6326 -68090 -6320 -68030
rect -6260 -68090 -6254 -68030
rect -6458 -68202 -6452 -68142
rect -6392 -68202 -6386 -68142
rect -6452 -68240 -6392 -68202
rect -6476 -68246 -6368 -68240
rect -6476 -68280 -6464 -68246
rect -6380 -68280 -6368 -68246
rect -6476 -68286 -6368 -68280
rect -6578 -68362 -6568 -68330
rect -6792 -68706 -6786 -68366
rect -6832 -68718 -6786 -68706
rect -6574 -68706 -6568 -68362
rect -6534 -68362 -6518 -68330
rect -6320 -68330 -6260 -68090
rect -6218 -68246 -6110 -68240
rect -6218 -68280 -6206 -68246
rect -6122 -68280 -6110 -68246
rect -6218 -68286 -6110 -68280
rect -5960 -68246 -5852 -68240
rect -5960 -68280 -5948 -68246
rect -5864 -68280 -5852 -68246
rect -5960 -68286 -5852 -68280
rect -6534 -68706 -6528 -68362
rect -6320 -68372 -6310 -68330
rect -6574 -68718 -6528 -68706
rect -6316 -68706 -6310 -68372
rect -6276 -68372 -6260 -68330
rect -6058 -68330 -6012 -68318
rect -6276 -68706 -6270 -68372
rect -6058 -68652 -6052 -68330
rect -6316 -68718 -6270 -68706
rect -6064 -68706 -6052 -68652
rect -6018 -68652 -6012 -68330
rect -5800 -68330 -5754 -68318
rect -6018 -68706 -6004 -68652
rect -5800 -68660 -5794 -68330
rect -6992 -68756 -6884 -68750
rect -6992 -68790 -6980 -68756
rect -6896 -68790 -6884 -68756
rect -6992 -68796 -6884 -68790
rect -6734 -68756 -6626 -68750
rect -6734 -68790 -6722 -68756
rect -6638 -68790 -6626 -68756
rect -6734 -68796 -6626 -68790
rect -6476 -68756 -6368 -68750
rect -6476 -68790 -6464 -68756
rect -6380 -68790 -6368 -68756
rect -6476 -68796 -6368 -68790
rect -6218 -68756 -6110 -68750
rect -6218 -68790 -6206 -68756
rect -6122 -68790 -6110 -68756
rect -6218 -68796 -6110 -68790
rect -6966 -68838 -6906 -68796
rect -6192 -68838 -6132 -68796
rect -6972 -68898 -6966 -68838
rect -6906 -68898 -6900 -68838
rect -6198 -68898 -6192 -68838
rect -6132 -68898 -6126 -68838
rect -6064 -68952 -6004 -68706
rect -5808 -68706 -5794 -68660
rect -5760 -68660 -5754 -68330
rect -5760 -68706 -5748 -68660
rect -5960 -68756 -5852 -68750
rect -5960 -68790 -5948 -68756
rect -5864 -68790 -5852 -68756
rect -5960 -68796 -5852 -68790
rect -5936 -68832 -5876 -68796
rect -5808 -68832 -5748 -68706
rect -5936 -68892 -5748 -68832
rect -7106 -69012 -7100 -68952
rect -7040 -69012 -7034 -68952
rect -6070 -69012 -6064 -68952
rect -6004 -69012 -5998 -68952
rect -5936 -69122 -5876 -68892
rect -5808 -69122 -5748 -68892
rect -7466 -69154 -5688 -69122
rect -7466 -69222 -7430 -69154
rect -5722 -69222 -5688 -69154
rect -7466 -69252 -5688 -69222
rect -7690 -69704 -7578 -69618
rect -6978 -69704 -6968 -69404
rect -6076 -69704 -6066 -69404
rect -5466 -69618 -5460 -67958
rect -5360 -69618 -5354 -67958
rect -5466 -69704 -5354 -69618
rect -7690 -69710 -5354 -69704
rect -7690 -69810 -7584 -69710
rect -5460 -69810 -5354 -69710
rect -7690 -69816 -5354 -69810
rect -3690 -67958 -3578 -67874
rect -3690 -69618 -3684 -67958
rect -3584 -69618 -3578 -67958
rect -2578 -67920 -2518 -67914
rect -3100 -68046 -3094 -67986
rect -3034 -68046 -3028 -67986
rect -3250 -68246 -3142 -68240
rect -3250 -68280 -3238 -68246
rect -3154 -68280 -3142 -68246
rect -3250 -68286 -3142 -68280
rect -3348 -68330 -3302 -68318
rect -3348 -68652 -3342 -68330
rect -3356 -68706 -3342 -68652
rect -3308 -68652 -3302 -68330
rect -3094 -68330 -3034 -68046
rect -2846 -68090 -2840 -68030
rect -2780 -68090 -2774 -68030
rect -2992 -68246 -2884 -68240
rect -2992 -68280 -2980 -68246
rect -2896 -68280 -2884 -68246
rect -2992 -68286 -2884 -68280
rect -3094 -68400 -3084 -68330
rect -3308 -68706 -3296 -68652
rect -3090 -68670 -3084 -68400
rect -3356 -68826 -3296 -68706
rect -3100 -68706 -3084 -68670
rect -3050 -68400 -3034 -68330
rect -2840 -68330 -2780 -68090
rect -2714 -68202 -2708 -68142
rect -2648 -68202 -2642 -68142
rect -2708 -68240 -2648 -68202
rect -2734 -68246 -2626 -68240
rect -2734 -68280 -2722 -68246
rect -2638 -68280 -2626 -68246
rect -2734 -68286 -2626 -68280
rect -2840 -68366 -2826 -68330
rect -3050 -68670 -3044 -68400
rect -3050 -68706 -3040 -68670
rect -3250 -68756 -3142 -68750
rect -3250 -68790 -3238 -68756
rect -3154 -68790 -3142 -68756
rect -3250 -68796 -3142 -68790
rect -3226 -68826 -3166 -68796
rect -3356 -68886 -3166 -68826
rect -3356 -69122 -3296 -68886
rect -3226 -69122 -3166 -68886
rect -3100 -68952 -3040 -68706
rect -2832 -68706 -2826 -68366
rect -2792 -68366 -2780 -68330
rect -2578 -68330 -2518 -67980
rect -1466 -67958 -1354 -67872
rect -72 -67809 416 -67778
rect -72 -67843 -43 -67809
rect -9 -67843 49 -67809
rect 83 -67843 141 -67809
rect 175 -67843 416 -67809
rect -72 -67866 416 -67843
rect 2540 -67866 2646 -67766
rect 4310 -67766 6646 -67760
rect 4310 -67778 4416 -67766
rect -72 -67872 2646 -67866
rect -72 -67874 422 -67872
rect -2326 -68090 -2320 -68030
rect -2260 -68090 -2254 -68030
rect -2458 -68202 -2452 -68142
rect -2392 -68202 -2386 -68142
rect -2452 -68240 -2392 -68202
rect -2476 -68246 -2368 -68240
rect -2476 -68280 -2464 -68246
rect -2380 -68280 -2368 -68246
rect -2476 -68286 -2368 -68280
rect -2578 -68362 -2568 -68330
rect -2792 -68706 -2786 -68366
rect -2832 -68718 -2786 -68706
rect -2574 -68706 -2568 -68362
rect -2534 -68362 -2518 -68330
rect -2320 -68330 -2260 -68090
rect -2218 -68246 -2110 -68240
rect -2218 -68280 -2206 -68246
rect -2122 -68280 -2110 -68246
rect -2218 -68286 -2110 -68280
rect -1960 -68246 -1852 -68240
rect -1960 -68280 -1948 -68246
rect -1864 -68280 -1852 -68246
rect -1960 -68286 -1852 -68280
rect -2534 -68706 -2528 -68362
rect -2320 -68372 -2310 -68330
rect -2574 -68718 -2528 -68706
rect -2316 -68706 -2310 -68372
rect -2276 -68372 -2260 -68330
rect -2058 -68330 -2012 -68318
rect -2276 -68706 -2270 -68372
rect -2058 -68652 -2052 -68330
rect -2316 -68718 -2270 -68706
rect -2064 -68706 -2052 -68652
rect -2018 -68652 -2012 -68330
rect -1800 -68330 -1754 -68318
rect -2018 -68706 -2004 -68652
rect -1800 -68660 -1794 -68330
rect -2992 -68756 -2884 -68750
rect -2992 -68790 -2980 -68756
rect -2896 -68790 -2884 -68756
rect -2992 -68796 -2884 -68790
rect -2734 -68756 -2626 -68750
rect -2734 -68790 -2722 -68756
rect -2638 -68790 -2626 -68756
rect -2734 -68796 -2626 -68790
rect -2476 -68756 -2368 -68750
rect -2476 -68790 -2464 -68756
rect -2380 -68790 -2368 -68756
rect -2476 -68796 -2368 -68790
rect -2218 -68756 -2110 -68750
rect -2218 -68790 -2206 -68756
rect -2122 -68790 -2110 -68756
rect -2218 -68796 -2110 -68790
rect -2966 -68838 -2906 -68796
rect -2192 -68838 -2132 -68796
rect -2972 -68898 -2966 -68838
rect -2906 -68898 -2900 -68838
rect -2198 -68898 -2192 -68838
rect -2132 -68898 -2126 -68838
rect -2064 -68952 -2004 -68706
rect -1808 -68706 -1794 -68660
rect -1760 -68660 -1754 -68330
rect -1760 -68706 -1748 -68660
rect -1960 -68756 -1852 -68750
rect -1960 -68790 -1948 -68756
rect -1864 -68790 -1852 -68756
rect -1960 -68796 -1852 -68790
rect -1936 -68832 -1876 -68796
rect -1808 -68832 -1748 -68706
rect -1936 -68892 -1748 -68832
rect -3106 -69012 -3100 -68952
rect -3040 -69012 -3034 -68952
rect -2070 -69012 -2064 -68952
rect -2004 -69012 -1998 -68952
rect -1936 -69122 -1876 -68892
rect -1808 -69122 -1748 -68892
rect -3466 -69154 -1688 -69122
rect -3466 -69222 -3430 -69154
rect -1722 -69222 -1688 -69154
rect -3466 -69252 -1688 -69222
rect -3690 -69704 -3578 -69618
rect -2978 -69704 -2968 -69404
rect -2076 -69704 -2066 -69404
rect -1466 -69618 -1460 -67958
rect -1360 -69618 -1354 -67958
rect -1466 -69704 -1354 -69618
rect -3690 -69710 -1354 -69704
rect -3690 -69810 -3584 -69710
rect -1460 -69810 -1354 -69710
rect -3690 -69816 -1354 -69810
rect 310 -67958 422 -67874
rect 310 -69618 316 -67958
rect 416 -69618 422 -67958
rect 1422 -67920 1482 -67914
rect 900 -68046 906 -67986
rect 966 -68046 972 -67986
rect 750 -68246 858 -68240
rect 750 -68280 762 -68246
rect 846 -68280 858 -68246
rect 750 -68286 858 -68280
rect 652 -68330 698 -68318
rect 652 -68652 658 -68330
rect 644 -68706 658 -68652
rect 692 -68652 698 -68330
rect 906 -68330 966 -68046
rect 1154 -68090 1160 -68030
rect 1220 -68090 1226 -68030
rect 1008 -68246 1116 -68240
rect 1008 -68280 1020 -68246
rect 1104 -68280 1116 -68246
rect 1008 -68286 1116 -68280
rect 906 -68400 916 -68330
rect 692 -68706 704 -68652
rect 910 -68670 916 -68400
rect 644 -68826 704 -68706
rect 900 -68706 916 -68670
rect 950 -68400 966 -68330
rect 1160 -68330 1220 -68090
rect 1286 -68202 1292 -68142
rect 1352 -68202 1358 -68142
rect 1292 -68240 1352 -68202
rect 1266 -68246 1374 -68240
rect 1266 -68280 1278 -68246
rect 1362 -68280 1374 -68246
rect 1266 -68286 1374 -68280
rect 1160 -68366 1174 -68330
rect 950 -68670 956 -68400
rect 950 -68706 960 -68670
rect 750 -68756 858 -68750
rect 750 -68790 762 -68756
rect 846 -68790 858 -68756
rect 750 -68796 858 -68790
rect 774 -68826 834 -68796
rect 644 -68886 834 -68826
rect 644 -69122 704 -68886
rect 774 -69122 834 -68886
rect 900 -68952 960 -68706
rect 1168 -68706 1174 -68366
rect 1208 -68366 1220 -68330
rect 1422 -68330 1482 -67980
rect 2534 -67958 2646 -67872
rect 3928 -67809 4416 -67778
rect 3928 -67843 3957 -67809
rect 3991 -67843 4049 -67809
rect 4083 -67843 4141 -67809
rect 4175 -67843 4416 -67809
rect 3928 -67866 4416 -67843
rect 6540 -67866 6646 -67766
rect 3928 -67872 6646 -67866
rect 3928 -67874 4422 -67872
rect 1674 -68090 1680 -68030
rect 1740 -68090 1746 -68030
rect 1542 -68202 1548 -68142
rect 1608 -68202 1614 -68142
rect 1548 -68240 1608 -68202
rect 1524 -68246 1632 -68240
rect 1524 -68280 1536 -68246
rect 1620 -68280 1632 -68246
rect 1524 -68286 1632 -68280
rect 1422 -68362 1432 -68330
rect 1208 -68706 1214 -68366
rect 1168 -68718 1214 -68706
rect 1426 -68706 1432 -68362
rect 1466 -68362 1482 -68330
rect 1680 -68330 1740 -68090
rect 1782 -68246 1890 -68240
rect 1782 -68280 1794 -68246
rect 1878 -68280 1890 -68246
rect 1782 -68286 1890 -68280
rect 2040 -68246 2148 -68240
rect 2040 -68280 2052 -68246
rect 2136 -68280 2148 -68246
rect 2040 -68286 2148 -68280
rect 1466 -68706 1472 -68362
rect 1680 -68372 1690 -68330
rect 1426 -68718 1472 -68706
rect 1684 -68706 1690 -68372
rect 1724 -68372 1740 -68330
rect 1942 -68330 1988 -68318
rect 1724 -68706 1730 -68372
rect 1942 -68652 1948 -68330
rect 1684 -68718 1730 -68706
rect 1936 -68706 1948 -68652
rect 1982 -68652 1988 -68330
rect 2200 -68330 2246 -68318
rect 1982 -68706 1996 -68652
rect 2200 -68660 2206 -68330
rect 1008 -68756 1116 -68750
rect 1008 -68790 1020 -68756
rect 1104 -68790 1116 -68756
rect 1008 -68796 1116 -68790
rect 1266 -68756 1374 -68750
rect 1266 -68790 1278 -68756
rect 1362 -68790 1374 -68756
rect 1266 -68796 1374 -68790
rect 1524 -68756 1632 -68750
rect 1524 -68790 1536 -68756
rect 1620 -68790 1632 -68756
rect 1524 -68796 1632 -68790
rect 1782 -68756 1890 -68750
rect 1782 -68790 1794 -68756
rect 1878 -68790 1890 -68756
rect 1782 -68796 1890 -68790
rect 1034 -68838 1094 -68796
rect 1808 -68838 1868 -68796
rect 1028 -68898 1034 -68838
rect 1094 -68898 1100 -68838
rect 1802 -68898 1808 -68838
rect 1868 -68898 1874 -68838
rect 1936 -68952 1996 -68706
rect 2192 -68706 2206 -68660
rect 2240 -68660 2246 -68330
rect 2240 -68706 2252 -68660
rect 2040 -68756 2148 -68750
rect 2040 -68790 2052 -68756
rect 2136 -68790 2148 -68756
rect 2040 -68796 2148 -68790
rect 2064 -68832 2124 -68796
rect 2192 -68832 2252 -68706
rect 2064 -68892 2252 -68832
rect 894 -69012 900 -68952
rect 960 -69012 966 -68952
rect 1930 -69012 1936 -68952
rect 1996 -69012 2002 -68952
rect 2064 -69122 2124 -68892
rect 2192 -69122 2252 -68892
rect 534 -69154 2312 -69122
rect 534 -69222 570 -69154
rect 2278 -69222 2312 -69154
rect 534 -69252 2312 -69222
rect 310 -69704 422 -69618
rect 1022 -69704 1032 -69404
rect 1924 -69704 1934 -69404
rect 2534 -69618 2540 -67958
rect 2640 -69618 2646 -67958
rect 2534 -69704 2646 -69618
rect 310 -69710 2646 -69704
rect 310 -69810 416 -69710
rect 2540 -69810 2646 -69710
rect 310 -69816 2646 -69810
rect 4310 -67958 4422 -67874
rect 4310 -69618 4316 -67958
rect 4416 -69618 4422 -67958
rect 5422 -67920 5482 -67914
rect 4900 -68046 4906 -67986
rect 4966 -68046 4972 -67986
rect 4750 -68246 4858 -68240
rect 4750 -68280 4762 -68246
rect 4846 -68280 4858 -68246
rect 4750 -68286 4858 -68280
rect 4652 -68330 4698 -68318
rect 4652 -68652 4658 -68330
rect 4644 -68706 4658 -68652
rect 4692 -68652 4698 -68330
rect 4906 -68330 4966 -68046
rect 5154 -68090 5160 -68030
rect 5220 -68090 5226 -68030
rect 5008 -68246 5116 -68240
rect 5008 -68280 5020 -68246
rect 5104 -68280 5116 -68246
rect 5008 -68286 5116 -68280
rect 4906 -68400 4916 -68330
rect 4692 -68706 4704 -68652
rect 4910 -68670 4916 -68400
rect 4644 -68826 4704 -68706
rect 4900 -68706 4916 -68670
rect 4950 -68400 4966 -68330
rect 5160 -68330 5220 -68090
rect 5286 -68202 5292 -68142
rect 5352 -68202 5358 -68142
rect 5292 -68240 5352 -68202
rect 5266 -68246 5374 -68240
rect 5266 -68280 5278 -68246
rect 5362 -68280 5374 -68246
rect 5266 -68286 5374 -68280
rect 5160 -68366 5174 -68330
rect 4950 -68670 4956 -68400
rect 4950 -68706 4960 -68670
rect 4750 -68756 4858 -68750
rect 4750 -68790 4762 -68756
rect 4846 -68790 4858 -68756
rect 4750 -68796 4858 -68790
rect 4774 -68826 4834 -68796
rect 4644 -68886 4834 -68826
rect 4644 -69122 4704 -68886
rect 4774 -69122 4834 -68886
rect 4900 -68952 4960 -68706
rect 5168 -68706 5174 -68366
rect 5208 -68366 5220 -68330
rect 5422 -68330 5482 -67980
rect 6534 -67958 6646 -67872
rect 5674 -68090 5680 -68030
rect 5740 -68090 5746 -68030
rect 5542 -68202 5548 -68142
rect 5608 -68202 5614 -68142
rect 5548 -68240 5608 -68202
rect 5524 -68246 5632 -68240
rect 5524 -68280 5536 -68246
rect 5620 -68280 5632 -68246
rect 5524 -68286 5632 -68280
rect 5422 -68362 5432 -68330
rect 5208 -68706 5214 -68366
rect 5168 -68718 5214 -68706
rect 5426 -68706 5432 -68362
rect 5466 -68362 5482 -68330
rect 5680 -68330 5740 -68090
rect 5782 -68246 5890 -68240
rect 5782 -68280 5794 -68246
rect 5878 -68280 5890 -68246
rect 5782 -68286 5890 -68280
rect 6040 -68246 6148 -68240
rect 6040 -68280 6052 -68246
rect 6136 -68280 6148 -68246
rect 6040 -68286 6148 -68280
rect 5466 -68706 5472 -68362
rect 5680 -68372 5690 -68330
rect 5426 -68718 5472 -68706
rect 5684 -68706 5690 -68372
rect 5724 -68372 5740 -68330
rect 5942 -68330 5988 -68318
rect 5724 -68706 5730 -68372
rect 5942 -68652 5948 -68330
rect 5684 -68718 5730 -68706
rect 5936 -68706 5948 -68652
rect 5982 -68652 5988 -68330
rect 6200 -68330 6246 -68318
rect 5982 -68706 5996 -68652
rect 6200 -68660 6206 -68330
rect 5008 -68756 5116 -68750
rect 5008 -68790 5020 -68756
rect 5104 -68790 5116 -68756
rect 5008 -68796 5116 -68790
rect 5266 -68756 5374 -68750
rect 5266 -68790 5278 -68756
rect 5362 -68790 5374 -68756
rect 5266 -68796 5374 -68790
rect 5524 -68756 5632 -68750
rect 5524 -68790 5536 -68756
rect 5620 -68790 5632 -68756
rect 5524 -68796 5632 -68790
rect 5782 -68756 5890 -68750
rect 5782 -68790 5794 -68756
rect 5878 -68790 5890 -68756
rect 5782 -68796 5890 -68790
rect 5034 -68838 5094 -68796
rect 5808 -68838 5868 -68796
rect 5028 -68898 5034 -68838
rect 5094 -68898 5100 -68838
rect 5802 -68898 5808 -68838
rect 5868 -68898 5874 -68838
rect 5936 -68952 5996 -68706
rect 6192 -68706 6206 -68660
rect 6240 -68660 6246 -68330
rect 6240 -68706 6252 -68660
rect 6040 -68756 6148 -68750
rect 6040 -68790 6052 -68756
rect 6136 -68790 6148 -68756
rect 6040 -68796 6148 -68790
rect 6064 -68832 6124 -68796
rect 6192 -68832 6252 -68706
rect 6064 -68892 6252 -68832
rect 4894 -69012 4900 -68952
rect 4960 -69012 4966 -68952
rect 5930 -69012 5936 -68952
rect 5996 -69012 6002 -68952
rect 6064 -69122 6124 -68892
rect 6192 -69122 6252 -68892
rect 4534 -69154 6312 -69122
rect 4534 -69222 4570 -69154
rect 6278 -69222 6312 -69154
rect 4534 -69252 6312 -69222
rect 4310 -69704 4422 -69618
rect 5022 -69704 5032 -69404
rect 5924 -69704 5934 -69404
rect 6534 -69618 6540 -67958
rect 6640 -69618 6646 -67958
rect 6534 -69704 6646 -69618
rect 4310 -69710 6646 -69704
rect 4310 -69810 4416 -69710
rect 6540 -69810 6646 -69710
rect 4310 -69816 6646 -69810
rect -27690 -70386 -25354 -70380
rect -27690 -70486 -27584 -70386
rect -25460 -70486 -25354 -70386
rect -27690 -70492 -25354 -70486
rect -27690 -70578 -27578 -70492
rect -27690 -72238 -27684 -70578
rect -27584 -72238 -27578 -70578
rect -26978 -70792 -26968 -70492
rect -26076 -70792 -26066 -70492
rect -25466 -70578 -25354 -70492
rect -27466 -70974 -25688 -70944
rect -27466 -71042 -27430 -70974
rect -25722 -71042 -25688 -70974
rect -27466 -71074 -25688 -71042
rect -27356 -71310 -27296 -71074
rect -27226 -71310 -27166 -71074
rect -27106 -71244 -27100 -71184
rect -27040 -71244 -27034 -71184
rect -26070 -71244 -26064 -71184
rect -26004 -71244 -25998 -71184
rect -27356 -71370 -27166 -71310
rect -27356 -71490 -27296 -71370
rect -27226 -71400 -27166 -71370
rect -27250 -71406 -27142 -71400
rect -27250 -71440 -27238 -71406
rect -27154 -71440 -27142 -71406
rect -27250 -71446 -27142 -71440
rect -27356 -71544 -27342 -71490
rect -27348 -71866 -27342 -71544
rect -27308 -71544 -27296 -71490
rect -27100 -71490 -27040 -71244
rect -26972 -71358 -26966 -71298
rect -26906 -71358 -26900 -71298
rect -26198 -71358 -26192 -71298
rect -26132 -71358 -26126 -71298
rect -26966 -71400 -26906 -71358
rect -26192 -71400 -26132 -71358
rect -26992 -71406 -26884 -71400
rect -26992 -71440 -26980 -71406
rect -26896 -71440 -26884 -71406
rect -26992 -71446 -26884 -71440
rect -26734 -71406 -26626 -71400
rect -26734 -71440 -26722 -71406
rect -26638 -71440 -26626 -71406
rect -26734 -71446 -26626 -71440
rect -26476 -71406 -26368 -71400
rect -26476 -71440 -26464 -71406
rect -26380 -71440 -26368 -71406
rect -26476 -71446 -26368 -71440
rect -26218 -71406 -26110 -71400
rect -26218 -71440 -26206 -71406
rect -26122 -71440 -26110 -71406
rect -26218 -71446 -26110 -71440
rect -27100 -71526 -27084 -71490
rect -27308 -71866 -27302 -71544
rect -27090 -71796 -27084 -71526
rect -27348 -71878 -27302 -71866
rect -27094 -71866 -27084 -71796
rect -27050 -71526 -27040 -71490
rect -26832 -71490 -26786 -71478
rect -27050 -71796 -27044 -71526
rect -27050 -71866 -27034 -71796
rect -26832 -71830 -26826 -71490
rect -27250 -71916 -27142 -71910
rect -27250 -71950 -27238 -71916
rect -27154 -71950 -27142 -71916
rect -27250 -71956 -27142 -71950
rect -27094 -72150 -27034 -71866
rect -26840 -71866 -26826 -71830
rect -26792 -71830 -26786 -71490
rect -26574 -71490 -26528 -71478
rect -26792 -71866 -26780 -71830
rect -26574 -71834 -26568 -71490
rect -26992 -71916 -26884 -71910
rect -26992 -71950 -26980 -71916
rect -26896 -71950 -26884 -71916
rect -26992 -71956 -26884 -71950
rect -26840 -72106 -26780 -71866
rect -26578 -71866 -26568 -71834
rect -26534 -71834 -26528 -71490
rect -26316 -71490 -26270 -71478
rect -26316 -71824 -26310 -71490
rect -26534 -71866 -26518 -71834
rect -26734 -71916 -26626 -71910
rect -26734 -71950 -26722 -71916
rect -26638 -71950 -26626 -71916
rect -26734 -71956 -26626 -71950
rect -26708 -71994 -26648 -71956
rect -26714 -72054 -26708 -71994
rect -26648 -72054 -26642 -71994
rect -27100 -72210 -27094 -72150
rect -27034 -72210 -27028 -72150
rect -26846 -72166 -26840 -72106
rect -26780 -72166 -26774 -72106
rect -27690 -72322 -27578 -72238
rect -26578 -72216 -26518 -71866
rect -26320 -71866 -26310 -71824
rect -26276 -71824 -26270 -71490
rect -26064 -71490 -26004 -71244
rect -25936 -71304 -25876 -71074
rect -25808 -71304 -25748 -71074
rect -25936 -71364 -25748 -71304
rect -25936 -71400 -25876 -71364
rect -25960 -71406 -25852 -71400
rect -25960 -71440 -25948 -71406
rect -25864 -71440 -25852 -71406
rect -25960 -71446 -25852 -71440
rect -26064 -71544 -26052 -71490
rect -26276 -71866 -26260 -71824
rect -26476 -71916 -26368 -71910
rect -26476 -71950 -26464 -71916
rect -26380 -71950 -26368 -71916
rect -26476 -71956 -26368 -71950
rect -26452 -71994 -26392 -71956
rect -26458 -72054 -26452 -71994
rect -26392 -72054 -26386 -71994
rect -26320 -72106 -26260 -71866
rect -26058 -71866 -26052 -71544
rect -26018 -71544 -26004 -71490
rect -25808 -71490 -25748 -71364
rect -25808 -71536 -25794 -71490
rect -26018 -71866 -26012 -71544
rect -26058 -71878 -26012 -71866
rect -25800 -71866 -25794 -71536
rect -25760 -71536 -25748 -71490
rect -25760 -71866 -25754 -71536
rect -25800 -71878 -25754 -71866
rect -26218 -71916 -26110 -71910
rect -26218 -71950 -26206 -71916
rect -26122 -71950 -26110 -71916
rect -26218 -71956 -26110 -71950
rect -25960 -71916 -25852 -71910
rect -25960 -71950 -25948 -71916
rect -25864 -71950 -25852 -71916
rect -25960 -71956 -25852 -71950
rect -26326 -72166 -26320 -72106
rect -26260 -72166 -26254 -72106
rect -26578 -72282 -26518 -72276
rect -25466 -72238 -25460 -70578
rect -25360 -72238 -25354 -70578
rect -28072 -72324 -27578 -72322
rect -25466 -72324 -25354 -72238
rect -23690 -70386 -21354 -70380
rect -23690 -70486 -23584 -70386
rect -21460 -70486 -21354 -70386
rect -23690 -70492 -21354 -70486
rect -23690 -70578 -23578 -70492
rect -23690 -72238 -23684 -70578
rect -23584 -72238 -23578 -70578
rect -22978 -70792 -22968 -70492
rect -22076 -70792 -22066 -70492
rect -21466 -70578 -21354 -70492
rect -23466 -70974 -21688 -70944
rect -23466 -71042 -23430 -70974
rect -21722 -71042 -21688 -70974
rect -23466 -71074 -21688 -71042
rect -23356 -71310 -23296 -71074
rect -23226 -71310 -23166 -71074
rect -23106 -71244 -23100 -71184
rect -23040 -71244 -23034 -71184
rect -22070 -71244 -22064 -71184
rect -22004 -71244 -21998 -71184
rect -23356 -71370 -23166 -71310
rect -23356 -71490 -23296 -71370
rect -23226 -71400 -23166 -71370
rect -23250 -71406 -23142 -71400
rect -23250 -71440 -23238 -71406
rect -23154 -71440 -23142 -71406
rect -23250 -71446 -23142 -71440
rect -23356 -71544 -23342 -71490
rect -23348 -71866 -23342 -71544
rect -23308 -71544 -23296 -71490
rect -23100 -71490 -23040 -71244
rect -22972 -71358 -22966 -71298
rect -22906 -71358 -22900 -71298
rect -22198 -71358 -22192 -71298
rect -22132 -71358 -22126 -71298
rect -22966 -71400 -22906 -71358
rect -22192 -71400 -22132 -71358
rect -22992 -71406 -22884 -71400
rect -22992 -71440 -22980 -71406
rect -22896 -71440 -22884 -71406
rect -22992 -71446 -22884 -71440
rect -22734 -71406 -22626 -71400
rect -22734 -71440 -22722 -71406
rect -22638 -71440 -22626 -71406
rect -22734 -71446 -22626 -71440
rect -22476 -71406 -22368 -71400
rect -22476 -71440 -22464 -71406
rect -22380 -71440 -22368 -71406
rect -22476 -71446 -22368 -71440
rect -22218 -71406 -22110 -71400
rect -22218 -71440 -22206 -71406
rect -22122 -71440 -22110 -71406
rect -22218 -71446 -22110 -71440
rect -23100 -71526 -23084 -71490
rect -23308 -71866 -23302 -71544
rect -23090 -71796 -23084 -71526
rect -23348 -71878 -23302 -71866
rect -23094 -71866 -23084 -71796
rect -23050 -71526 -23040 -71490
rect -22832 -71490 -22786 -71478
rect -23050 -71796 -23044 -71526
rect -23050 -71866 -23034 -71796
rect -22832 -71830 -22826 -71490
rect -23250 -71916 -23142 -71910
rect -23250 -71950 -23238 -71916
rect -23154 -71950 -23142 -71916
rect -23250 -71956 -23142 -71950
rect -23094 -72150 -23034 -71866
rect -22840 -71866 -22826 -71830
rect -22792 -71830 -22786 -71490
rect -22574 -71490 -22528 -71478
rect -22792 -71866 -22780 -71830
rect -22574 -71834 -22568 -71490
rect -22992 -71916 -22884 -71910
rect -22992 -71950 -22980 -71916
rect -22896 -71950 -22884 -71916
rect -22992 -71956 -22884 -71950
rect -22840 -72106 -22780 -71866
rect -22578 -71866 -22568 -71834
rect -22534 -71834 -22528 -71490
rect -22316 -71490 -22270 -71478
rect -22316 -71824 -22310 -71490
rect -22534 -71866 -22518 -71834
rect -22734 -71916 -22626 -71910
rect -22734 -71950 -22722 -71916
rect -22638 -71950 -22626 -71916
rect -22734 -71956 -22626 -71950
rect -22708 -71994 -22648 -71956
rect -22714 -72054 -22708 -71994
rect -22648 -72054 -22642 -71994
rect -23100 -72210 -23094 -72150
rect -23034 -72210 -23028 -72150
rect -22846 -72166 -22840 -72106
rect -22780 -72166 -22774 -72106
rect -23690 -72322 -23578 -72238
rect -22578 -72216 -22518 -71866
rect -22320 -71866 -22310 -71824
rect -22276 -71824 -22270 -71490
rect -22064 -71490 -22004 -71244
rect -21936 -71304 -21876 -71074
rect -21808 -71304 -21748 -71074
rect -21936 -71364 -21748 -71304
rect -21936 -71400 -21876 -71364
rect -21960 -71406 -21852 -71400
rect -21960 -71440 -21948 -71406
rect -21864 -71440 -21852 -71406
rect -21960 -71446 -21852 -71440
rect -22064 -71544 -22052 -71490
rect -22276 -71866 -22260 -71824
rect -22476 -71916 -22368 -71910
rect -22476 -71950 -22464 -71916
rect -22380 -71950 -22368 -71916
rect -22476 -71956 -22368 -71950
rect -22452 -71994 -22392 -71956
rect -22458 -72054 -22452 -71994
rect -22392 -72054 -22386 -71994
rect -22320 -72106 -22260 -71866
rect -22058 -71866 -22052 -71544
rect -22018 -71544 -22004 -71490
rect -21808 -71490 -21748 -71364
rect -21808 -71536 -21794 -71490
rect -22018 -71866 -22012 -71544
rect -22058 -71878 -22012 -71866
rect -21800 -71866 -21794 -71536
rect -21760 -71536 -21748 -71490
rect -21760 -71866 -21754 -71536
rect -21800 -71878 -21754 -71866
rect -22218 -71916 -22110 -71910
rect -22218 -71950 -22206 -71916
rect -22122 -71950 -22110 -71916
rect -22218 -71956 -22110 -71950
rect -21960 -71916 -21852 -71910
rect -21960 -71950 -21948 -71916
rect -21864 -71950 -21852 -71916
rect -21960 -71956 -21852 -71950
rect -22326 -72166 -22320 -72106
rect -22260 -72166 -22254 -72106
rect -22578 -72282 -22518 -72276
rect -21466 -72238 -21460 -70578
rect -21360 -72238 -21354 -70578
rect -28072 -72330 -25354 -72324
rect -28072 -72353 -27584 -72330
rect -28072 -72387 -28043 -72353
rect -28009 -72387 -27951 -72353
rect -27917 -72387 -27859 -72353
rect -27825 -72387 -27584 -72353
rect -28072 -72418 -27584 -72387
rect -27690 -72430 -27584 -72418
rect -25460 -72430 -25354 -72330
rect -24072 -72324 -23578 -72322
rect -21466 -72324 -21354 -72238
rect -19690 -70386 -17354 -70380
rect -19690 -70486 -19584 -70386
rect -17460 -70486 -17354 -70386
rect -19690 -70492 -17354 -70486
rect -19690 -70578 -19578 -70492
rect -19690 -72238 -19684 -70578
rect -19584 -72238 -19578 -70578
rect -18978 -70792 -18968 -70492
rect -18076 -70792 -18066 -70492
rect -17466 -70578 -17354 -70492
rect -19466 -70974 -17688 -70944
rect -19466 -71042 -19430 -70974
rect -17722 -71042 -17688 -70974
rect -19466 -71074 -17688 -71042
rect -19356 -71310 -19296 -71074
rect -19226 -71310 -19166 -71074
rect -19106 -71244 -19100 -71184
rect -19040 -71244 -19034 -71184
rect -18070 -71244 -18064 -71184
rect -18004 -71244 -17998 -71184
rect -19356 -71370 -19166 -71310
rect -19356 -71490 -19296 -71370
rect -19226 -71400 -19166 -71370
rect -19250 -71406 -19142 -71400
rect -19250 -71440 -19238 -71406
rect -19154 -71440 -19142 -71406
rect -19250 -71446 -19142 -71440
rect -19356 -71544 -19342 -71490
rect -19348 -71866 -19342 -71544
rect -19308 -71544 -19296 -71490
rect -19100 -71490 -19040 -71244
rect -18972 -71358 -18966 -71298
rect -18906 -71358 -18900 -71298
rect -18198 -71358 -18192 -71298
rect -18132 -71358 -18126 -71298
rect -18966 -71400 -18906 -71358
rect -18192 -71400 -18132 -71358
rect -18992 -71406 -18884 -71400
rect -18992 -71440 -18980 -71406
rect -18896 -71440 -18884 -71406
rect -18992 -71446 -18884 -71440
rect -18734 -71406 -18626 -71400
rect -18734 -71440 -18722 -71406
rect -18638 -71440 -18626 -71406
rect -18734 -71446 -18626 -71440
rect -18476 -71406 -18368 -71400
rect -18476 -71440 -18464 -71406
rect -18380 -71440 -18368 -71406
rect -18476 -71446 -18368 -71440
rect -18218 -71406 -18110 -71400
rect -18218 -71440 -18206 -71406
rect -18122 -71440 -18110 -71406
rect -18218 -71446 -18110 -71440
rect -19100 -71526 -19084 -71490
rect -19308 -71866 -19302 -71544
rect -19090 -71796 -19084 -71526
rect -19348 -71878 -19302 -71866
rect -19094 -71866 -19084 -71796
rect -19050 -71526 -19040 -71490
rect -18832 -71490 -18786 -71478
rect -19050 -71796 -19044 -71526
rect -19050 -71866 -19034 -71796
rect -18832 -71830 -18826 -71490
rect -19250 -71916 -19142 -71910
rect -19250 -71950 -19238 -71916
rect -19154 -71950 -19142 -71916
rect -19250 -71956 -19142 -71950
rect -19094 -72150 -19034 -71866
rect -18840 -71866 -18826 -71830
rect -18792 -71830 -18786 -71490
rect -18574 -71490 -18528 -71478
rect -18792 -71866 -18780 -71830
rect -18574 -71834 -18568 -71490
rect -18992 -71916 -18884 -71910
rect -18992 -71950 -18980 -71916
rect -18896 -71950 -18884 -71916
rect -18992 -71956 -18884 -71950
rect -18840 -72106 -18780 -71866
rect -18578 -71866 -18568 -71834
rect -18534 -71834 -18528 -71490
rect -18316 -71490 -18270 -71478
rect -18316 -71824 -18310 -71490
rect -18534 -71866 -18518 -71834
rect -18734 -71916 -18626 -71910
rect -18734 -71950 -18722 -71916
rect -18638 -71950 -18626 -71916
rect -18734 -71956 -18626 -71950
rect -18708 -71994 -18648 -71956
rect -18714 -72054 -18708 -71994
rect -18648 -72054 -18642 -71994
rect -19100 -72210 -19094 -72150
rect -19034 -72210 -19028 -72150
rect -18846 -72166 -18840 -72106
rect -18780 -72166 -18774 -72106
rect -19690 -72322 -19578 -72238
rect -18578 -72216 -18518 -71866
rect -18320 -71866 -18310 -71824
rect -18276 -71824 -18270 -71490
rect -18064 -71490 -18004 -71244
rect -17936 -71304 -17876 -71074
rect -17808 -71304 -17748 -71074
rect -17936 -71364 -17748 -71304
rect -17936 -71400 -17876 -71364
rect -17960 -71406 -17852 -71400
rect -17960 -71440 -17948 -71406
rect -17864 -71440 -17852 -71406
rect -17960 -71446 -17852 -71440
rect -18064 -71544 -18052 -71490
rect -18276 -71866 -18260 -71824
rect -18476 -71916 -18368 -71910
rect -18476 -71950 -18464 -71916
rect -18380 -71950 -18368 -71916
rect -18476 -71956 -18368 -71950
rect -18452 -71994 -18392 -71956
rect -18458 -72054 -18452 -71994
rect -18392 -72054 -18386 -71994
rect -18320 -72106 -18260 -71866
rect -18058 -71866 -18052 -71544
rect -18018 -71544 -18004 -71490
rect -17808 -71490 -17748 -71364
rect -17808 -71536 -17794 -71490
rect -18018 -71866 -18012 -71544
rect -18058 -71878 -18012 -71866
rect -17800 -71866 -17794 -71536
rect -17760 -71536 -17748 -71490
rect -17760 -71866 -17754 -71536
rect -17800 -71878 -17754 -71866
rect -18218 -71916 -18110 -71910
rect -18218 -71950 -18206 -71916
rect -18122 -71950 -18110 -71916
rect -18218 -71956 -18110 -71950
rect -17960 -71916 -17852 -71910
rect -17960 -71950 -17948 -71916
rect -17864 -71950 -17852 -71916
rect -17960 -71956 -17852 -71950
rect -18326 -72166 -18320 -72106
rect -18260 -72166 -18254 -72106
rect -18578 -72282 -18518 -72276
rect -17466 -72238 -17460 -70578
rect -17360 -72238 -17354 -70578
rect -24072 -72330 -21354 -72324
rect -24072 -72353 -23584 -72330
rect -24072 -72387 -24043 -72353
rect -24009 -72387 -23951 -72353
rect -23917 -72387 -23859 -72353
rect -23825 -72387 -23584 -72353
rect -24072 -72418 -23584 -72387
rect -27690 -72436 -25354 -72430
rect -23690 -72430 -23584 -72418
rect -21460 -72430 -21354 -72330
rect -20072 -72324 -19578 -72322
rect -17466 -72324 -17354 -72238
rect -15690 -70386 -13354 -70380
rect -15690 -70486 -15584 -70386
rect -13460 -70486 -13354 -70386
rect -15690 -70492 -13354 -70486
rect -15690 -70578 -15578 -70492
rect -15690 -72238 -15684 -70578
rect -15584 -72238 -15578 -70578
rect -14978 -70792 -14968 -70492
rect -14076 -70792 -14066 -70492
rect -13466 -70578 -13354 -70492
rect -15466 -70974 -13688 -70944
rect -15466 -71042 -15430 -70974
rect -13722 -71042 -13688 -70974
rect -15466 -71074 -13688 -71042
rect -15356 -71310 -15296 -71074
rect -15226 -71310 -15166 -71074
rect -15106 -71244 -15100 -71184
rect -15040 -71244 -15034 -71184
rect -14070 -71244 -14064 -71184
rect -14004 -71244 -13998 -71184
rect -15356 -71370 -15166 -71310
rect -15356 -71490 -15296 -71370
rect -15226 -71400 -15166 -71370
rect -15250 -71406 -15142 -71400
rect -15250 -71440 -15238 -71406
rect -15154 -71440 -15142 -71406
rect -15250 -71446 -15142 -71440
rect -15356 -71544 -15342 -71490
rect -15348 -71866 -15342 -71544
rect -15308 -71544 -15296 -71490
rect -15100 -71490 -15040 -71244
rect -14972 -71358 -14966 -71298
rect -14906 -71358 -14900 -71298
rect -14198 -71358 -14192 -71298
rect -14132 -71358 -14126 -71298
rect -14966 -71400 -14906 -71358
rect -14192 -71400 -14132 -71358
rect -14992 -71406 -14884 -71400
rect -14992 -71440 -14980 -71406
rect -14896 -71440 -14884 -71406
rect -14992 -71446 -14884 -71440
rect -14734 -71406 -14626 -71400
rect -14734 -71440 -14722 -71406
rect -14638 -71440 -14626 -71406
rect -14734 -71446 -14626 -71440
rect -14476 -71406 -14368 -71400
rect -14476 -71440 -14464 -71406
rect -14380 -71440 -14368 -71406
rect -14476 -71446 -14368 -71440
rect -14218 -71406 -14110 -71400
rect -14218 -71440 -14206 -71406
rect -14122 -71440 -14110 -71406
rect -14218 -71446 -14110 -71440
rect -15100 -71526 -15084 -71490
rect -15308 -71866 -15302 -71544
rect -15090 -71796 -15084 -71526
rect -15348 -71878 -15302 -71866
rect -15094 -71866 -15084 -71796
rect -15050 -71526 -15040 -71490
rect -14832 -71490 -14786 -71478
rect -15050 -71796 -15044 -71526
rect -15050 -71866 -15034 -71796
rect -14832 -71830 -14826 -71490
rect -15250 -71916 -15142 -71910
rect -15250 -71950 -15238 -71916
rect -15154 -71950 -15142 -71916
rect -15250 -71956 -15142 -71950
rect -15094 -72150 -15034 -71866
rect -14840 -71866 -14826 -71830
rect -14792 -71830 -14786 -71490
rect -14574 -71490 -14528 -71478
rect -14792 -71866 -14780 -71830
rect -14574 -71834 -14568 -71490
rect -14992 -71916 -14884 -71910
rect -14992 -71950 -14980 -71916
rect -14896 -71950 -14884 -71916
rect -14992 -71956 -14884 -71950
rect -14840 -72106 -14780 -71866
rect -14578 -71866 -14568 -71834
rect -14534 -71834 -14528 -71490
rect -14316 -71490 -14270 -71478
rect -14316 -71824 -14310 -71490
rect -14534 -71866 -14518 -71834
rect -14734 -71916 -14626 -71910
rect -14734 -71950 -14722 -71916
rect -14638 -71950 -14626 -71916
rect -14734 -71956 -14626 -71950
rect -14708 -71994 -14648 -71956
rect -14714 -72054 -14708 -71994
rect -14648 -72054 -14642 -71994
rect -15100 -72210 -15094 -72150
rect -15034 -72210 -15028 -72150
rect -14846 -72166 -14840 -72106
rect -14780 -72166 -14774 -72106
rect -15690 -72322 -15578 -72238
rect -14578 -72216 -14518 -71866
rect -14320 -71866 -14310 -71824
rect -14276 -71824 -14270 -71490
rect -14064 -71490 -14004 -71244
rect -13936 -71304 -13876 -71074
rect -13808 -71304 -13748 -71074
rect -13936 -71364 -13748 -71304
rect -13936 -71400 -13876 -71364
rect -13960 -71406 -13852 -71400
rect -13960 -71440 -13948 -71406
rect -13864 -71440 -13852 -71406
rect -13960 -71446 -13852 -71440
rect -14064 -71544 -14052 -71490
rect -14276 -71866 -14260 -71824
rect -14476 -71916 -14368 -71910
rect -14476 -71950 -14464 -71916
rect -14380 -71950 -14368 -71916
rect -14476 -71956 -14368 -71950
rect -14452 -71994 -14392 -71956
rect -14458 -72054 -14452 -71994
rect -14392 -72054 -14386 -71994
rect -14320 -72106 -14260 -71866
rect -14058 -71866 -14052 -71544
rect -14018 -71544 -14004 -71490
rect -13808 -71490 -13748 -71364
rect -13808 -71536 -13794 -71490
rect -14018 -71866 -14012 -71544
rect -14058 -71878 -14012 -71866
rect -13800 -71866 -13794 -71536
rect -13760 -71536 -13748 -71490
rect -13760 -71866 -13754 -71536
rect -13800 -71878 -13754 -71866
rect -14218 -71916 -14110 -71910
rect -14218 -71950 -14206 -71916
rect -14122 -71950 -14110 -71916
rect -14218 -71956 -14110 -71950
rect -13960 -71916 -13852 -71910
rect -13960 -71950 -13948 -71916
rect -13864 -71950 -13852 -71916
rect -13960 -71956 -13852 -71950
rect -14326 -72166 -14320 -72106
rect -14260 -72166 -14254 -72106
rect -14578 -72282 -14518 -72276
rect -13466 -72238 -13460 -70578
rect -13360 -72238 -13354 -70578
rect -20072 -72330 -17354 -72324
rect -20072 -72353 -19584 -72330
rect -20072 -72387 -20043 -72353
rect -20009 -72387 -19951 -72353
rect -19917 -72387 -19859 -72353
rect -19825 -72387 -19584 -72353
rect -20072 -72418 -19584 -72387
rect -23690 -72436 -21354 -72430
rect -19690 -72430 -19584 -72418
rect -17460 -72430 -17354 -72330
rect -16072 -72324 -15578 -72322
rect -13466 -72324 -13354 -72238
rect -11690 -70386 -9354 -70380
rect -11690 -70486 -11584 -70386
rect -9460 -70486 -9354 -70386
rect -11690 -70492 -9354 -70486
rect -11690 -70578 -11578 -70492
rect -11690 -72238 -11684 -70578
rect -11584 -72238 -11578 -70578
rect -10978 -70792 -10968 -70492
rect -10076 -70792 -10066 -70492
rect -9466 -70578 -9354 -70492
rect -11466 -70974 -9688 -70944
rect -11466 -71042 -11430 -70974
rect -9722 -71042 -9688 -70974
rect -11466 -71074 -9688 -71042
rect -11356 -71310 -11296 -71074
rect -11226 -71310 -11166 -71074
rect -11106 -71244 -11100 -71184
rect -11040 -71244 -11034 -71184
rect -10070 -71244 -10064 -71184
rect -10004 -71244 -9998 -71184
rect -11356 -71370 -11166 -71310
rect -11356 -71490 -11296 -71370
rect -11226 -71400 -11166 -71370
rect -11250 -71406 -11142 -71400
rect -11250 -71440 -11238 -71406
rect -11154 -71440 -11142 -71406
rect -11250 -71446 -11142 -71440
rect -11356 -71544 -11342 -71490
rect -11348 -71866 -11342 -71544
rect -11308 -71544 -11296 -71490
rect -11100 -71490 -11040 -71244
rect -10972 -71358 -10966 -71298
rect -10906 -71358 -10900 -71298
rect -10198 -71358 -10192 -71298
rect -10132 -71358 -10126 -71298
rect -10966 -71400 -10906 -71358
rect -10192 -71400 -10132 -71358
rect -10992 -71406 -10884 -71400
rect -10992 -71440 -10980 -71406
rect -10896 -71440 -10884 -71406
rect -10992 -71446 -10884 -71440
rect -10734 -71406 -10626 -71400
rect -10734 -71440 -10722 -71406
rect -10638 -71440 -10626 -71406
rect -10734 -71446 -10626 -71440
rect -10476 -71406 -10368 -71400
rect -10476 -71440 -10464 -71406
rect -10380 -71440 -10368 -71406
rect -10476 -71446 -10368 -71440
rect -10218 -71406 -10110 -71400
rect -10218 -71440 -10206 -71406
rect -10122 -71440 -10110 -71406
rect -10218 -71446 -10110 -71440
rect -11100 -71526 -11084 -71490
rect -11308 -71866 -11302 -71544
rect -11090 -71796 -11084 -71526
rect -11348 -71878 -11302 -71866
rect -11094 -71866 -11084 -71796
rect -11050 -71526 -11040 -71490
rect -10832 -71490 -10786 -71478
rect -11050 -71796 -11044 -71526
rect -11050 -71866 -11034 -71796
rect -10832 -71830 -10826 -71490
rect -11250 -71916 -11142 -71910
rect -11250 -71950 -11238 -71916
rect -11154 -71950 -11142 -71916
rect -11250 -71956 -11142 -71950
rect -11094 -72150 -11034 -71866
rect -10840 -71866 -10826 -71830
rect -10792 -71830 -10786 -71490
rect -10574 -71490 -10528 -71478
rect -10792 -71866 -10780 -71830
rect -10574 -71834 -10568 -71490
rect -10992 -71916 -10884 -71910
rect -10992 -71950 -10980 -71916
rect -10896 -71950 -10884 -71916
rect -10992 -71956 -10884 -71950
rect -10840 -72106 -10780 -71866
rect -10578 -71866 -10568 -71834
rect -10534 -71834 -10528 -71490
rect -10316 -71490 -10270 -71478
rect -10316 -71824 -10310 -71490
rect -10534 -71866 -10518 -71834
rect -10734 -71916 -10626 -71910
rect -10734 -71950 -10722 -71916
rect -10638 -71950 -10626 -71916
rect -10734 -71956 -10626 -71950
rect -10708 -71994 -10648 -71956
rect -10714 -72054 -10708 -71994
rect -10648 -72054 -10642 -71994
rect -11100 -72210 -11094 -72150
rect -11034 -72210 -11028 -72150
rect -10846 -72166 -10840 -72106
rect -10780 -72166 -10774 -72106
rect -11690 -72322 -11578 -72238
rect -10578 -72216 -10518 -71866
rect -10320 -71866 -10310 -71824
rect -10276 -71824 -10270 -71490
rect -10064 -71490 -10004 -71244
rect -9936 -71304 -9876 -71074
rect -9808 -71304 -9748 -71074
rect -9936 -71364 -9748 -71304
rect -9936 -71400 -9876 -71364
rect -9960 -71406 -9852 -71400
rect -9960 -71440 -9948 -71406
rect -9864 -71440 -9852 -71406
rect -9960 -71446 -9852 -71440
rect -10064 -71544 -10052 -71490
rect -10276 -71866 -10260 -71824
rect -10476 -71916 -10368 -71910
rect -10476 -71950 -10464 -71916
rect -10380 -71950 -10368 -71916
rect -10476 -71956 -10368 -71950
rect -10452 -71994 -10392 -71956
rect -10458 -72054 -10452 -71994
rect -10392 -72054 -10386 -71994
rect -10320 -72106 -10260 -71866
rect -10058 -71866 -10052 -71544
rect -10018 -71544 -10004 -71490
rect -9808 -71490 -9748 -71364
rect -9808 -71536 -9794 -71490
rect -10018 -71866 -10012 -71544
rect -10058 -71878 -10012 -71866
rect -9800 -71866 -9794 -71536
rect -9760 -71536 -9748 -71490
rect -9760 -71866 -9754 -71536
rect -9800 -71878 -9754 -71866
rect -10218 -71916 -10110 -71910
rect -10218 -71950 -10206 -71916
rect -10122 -71950 -10110 -71916
rect -10218 -71956 -10110 -71950
rect -9960 -71916 -9852 -71910
rect -9960 -71950 -9948 -71916
rect -9864 -71950 -9852 -71916
rect -9960 -71956 -9852 -71950
rect -10326 -72166 -10320 -72106
rect -10260 -72166 -10254 -72106
rect -10578 -72282 -10518 -72276
rect -9466 -72238 -9460 -70578
rect -9360 -72238 -9354 -70578
rect -16072 -72330 -13354 -72324
rect -16072 -72353 -15584 -72330
rect -16072 -72387 -16043 -72353
rect -16009 -72387 -15951 -72353
rect -15917 -72387 -15859 -72353
rect -15825 -72387 -15584 -72353
rect -16072 -72418 -15584 -72387
rect -19690 -72436 -17354 -72430
rect -15690 -72430 -15584 -72418
rect -13460 -72430 -13354 -72330
rect -12072 -72324 -11578 -72322
rect -9466 -72324 -9354 -72238
rect -7690 -70386 -5354 -70380
rect -7690 -70486 -7584 -70386
rect -5460 -70486 -5354 -70386
rect -7690 -70492 -5354 -70486
rect -7690 -70578 -7578 -70492
rect -7690 -72238 -7684 -70578
rect -7584 -72238 -7578 -70578
rect -6978 -70792 -6968 -70492
rect -6076 -70792 -6066 -70492
rect -5466 -70578 -5354 -70492
rect -7466 -70974 -5688 -70944
rect -7466 -71042 -7430 -70974
rect -5722 -71042 -5688 -70974
rect -7466 -71074 -5688 -71042
rect -7356 -71310 -7296 -71074
rect -7226 -71310 -7166 -71074
rect -7106 -71244 -7100 -71184
rect -7040 -71244 -7034 -71184
rect -6070 -71244 -6064 -71184
rect -6004 -71244 -5998 -71184
rect -7356 -71370 -7166 -71310
rect -7356 -71490 -7296 -71370
rect -7226 -71400 -7166 -71370
rect -7250 -71406 -7142 -71400
rect -7250 -71440 -7238 -71406
rect -7154 -71440 -7142 -71406
rect -7250 -71446 -7142 -71440
rect -7356 -71544 -7342 -71490
rect -7348 -71866 -7342 -71544
rect -7308 -71544 -7296 -71490
rect -7100 -71490 -7040 -71244
rect -6972 -71358 -6966 -71298
rect -6906 -71358 -6900 -71298
rect -6198 -71358 -6192 -71298
rect -6132 -71358 -6126 -71298
rect -6966 -71400 -6906 -71358
rect -6192 -71400 -6132 -71358
rect -6992 -71406 -6884 -71400
rect -6992 -71440 -6980 -71406
rect -6896 -71440 -6884 -71406
rect -6992 -71446 -6884 -71440
rect -6734 -71406 -6626 -71400
rect -6734 -71440 -6722 -71406
rect -6638 -71440 -6626 -71406
rect -6734 -71446 -6626 -71440
rect -6476 -71406 -6368 -71400
rect -6476 -71440 -6464 -71406
rect -6380 -71440 -6368 -71406
rect -6476 -71446 -6368 -71440
rect -6218 -71406 -6110 -71400
rect -6218 -71440 -6206 -71406
rect -6122 -71440 -6110 -71406
rect -6218 -71446 -6110 -71440
rect -7100 -71526 -7084 -71490
rect -7308 -71866 -7302 -71544
rect -7090 -71796 -7084 -71526
rect -7348 -71878 -7302 -71866
rect -7094 -71866 -7084 -71796
rect -7050 -71526 -7040 -71490
rect -6832 -71490 -6786 -71478
rect -7050 -71796 -7044 -71526
rect -7050 -71866 -7034 -71796
rect -6832 -71830 -6826 -71490
rect -7250 -71916 -7142 -71910
rect -7250 -71950 -7238 -71916
rect -7154 -71950 -7142 -71916
rect -7250 -71956 -7142 -71950
rect -7094 -72150 -7034 -71866
rect -6840 -71866 -6826 -71830
rect -6792 -71830 -6786 -71490
rect -6574 -71490 -6528 -71478
rect -6792 -71866 -6780 -71830
rect -6574 -71834 -6568 -71490
rect -6992 -71916 -6884 -71910
rect -6992 -71950 -6980 -71916
rect -6896 -71950 -6884 -71916
rect -6992 -71956 -6884 -71950
rect -6840 -72106 -6780 -71866
rect -6578 -71866 -6568 -71834
rect -6534 -71834 -6528 -71490
rect -6316 -71490 -6270 -71478
rect -6316 -71824 -6310 -71490
rect -6534 -71866 -6518 -71834
rect -6734 -71916 -6626 -71910
rect -6734 -71950 -6722 -71916
rect -6638 -71950 -6626 -71916
rect -6734 -71956 -6626 -71950
rect -6708 -71994 -6648 -71956
rect -6714 -72054 -6708 -71994
rect -6648 -72054 -6642 -71994
rect -7100 -72210 -7094 -72150
rect -7034 -72210 -7028 -72150
rect -6846 -72166 -6840 -72106
rect -6780 -72166 -6774 -72106
rect -7690 -72322 -7578 -72238
rect -6578 -72216 -6518 -71866
rect -6320 -71866 -6310 -71824
rect -6276 -71824 -6270 -71490
rect -6064 -71490 -6004 -71244
rect -5936 -71304 -5876 -71074
rect -5808 -71304 -5748 -71074
rect -5936 -71364 -5748 -71304
rect -5936 -71400 -5876 -71364
rect -5960 -71406 -5852 -71400
rect -5960 -71440 -5948 -71406
rect -5864 -71440 -5852 -71406
rect -5960 -71446 -5852 -71440
rect -6064 -71544 -6052 -71490
rect -6276 -71866 -6260 -71824
rect -6476 -71916 -6368 -71910
rect -6476 -71950 -6464 -71916
rect -6380 -71950 -6368 -71916
rect -6476 -71956 -6368 -71950
rect -6452 -71994 -6392 -71956
rect -6458 -72054 -6452 -71994
rect -6392 -72054 -6386 -71994
rect -6320 -72106 -6260 -71866
rect -6058 -71866 -6052 -71544
rect -6018 -71544 -6004 -71490
rect -5808 -71490 -5748 -71364
rect -5808 -71536 -5794 -71490
rect -6018 -71866 -6012 -71544
rect -6058 -71878 -6012 -71866
rect -5800 -71866 -5794 -71536
rect -5760 -71536 -5748 -71490
rect -5760 -71866 -5754 -71536
rect -5800 -71878 -5754 -71866
rect -6218 -71916 -6110 -71910
rect -6218 -71950 -6206 -71916
rect -6122 -71950 -6110 -71916
rect -6218 -71956 -6110 -71950
rect -5960 -71916 -5852 -71910
rect -5960 -71950 -5948 -71916
rect -5864 -71950 -5852 -71916
rect -5960 -71956 -5852 -71950
rect -6326 -72166 -6320 -72106
rect -6260 -72166 -6254 -72106
rect -6578 -72282 -6518 -72276
rect -5466 -72238 -5460 -70578
rect -5360 -72238 -5354 -70578
rect -12072 -72330 -9354 -72324
rect -12072 -72353 -11584 -72330
rect -12072 -72387 -12043 -72353
rect -12009 -72387 -11951 -72353
rect -11917 -72387 -11859 -72353
rect -11825 -72387 -11584 -72353
rect -12072 -72418 -11584 -72387
rect -15690 -72436 -13354 -72430
rect -11690 -72430 -11584 -72418
rect -9460 -72430 -9354 -72330
rect -8072 -72324 -7578 -72322
rect -5466 -72324 -5354 -72238
rect -3690 -70386 -1354 -70380
rect -3690 -70486 -3584 -70386
rect -1460 -70486 -1354 -70386
rect -3690 -70492 -1354 -70486
rect -3690 -70578 -3578 -70492
rect -3690 -72238 -3684 -70578
rect -3584 -72238 -3578 -70578
rect -2978 -70792 -2968 -70492
rect -2076 -70792 -2066 -70492
rect -1466 -70578 -1354 -70492
rect -3466 -70974 -1688 -70944
rect -3466 -71042 -3430 -70974
rect -1722 -71042 -1688 -70974
rect -3466 -71074 -1688 -71042
rect -3356 -71310 -3296 -71074
rect -3226 -71310 -3166 -71074
rect -3106 -71244 -3100 -71184
rect -3040 -71244 -3034 -71184
rect -2070 -71244 -2064 -71184
rect -2004 -71244 -1998 -71184
rect -3356 -71370 -3166 -71310
rect -3356 -71490 -3296 -71370
rect -3226 -71400 -3166 -71370
rect -3250 -71406 -3142 -71400
rect -3250 -71440 -3238 -71406
rect -3154 -71440 -3142 -71406
rect -3250 -71446 -3142 -71440
rect -3356 -71544 -3342 -71490
rect -3348 -71866 -3342 -71544
rect -3308 -71544 -3296 -71490
rect -3100 -71490 -3040 -71244
rect -2972 -71358 -2966 -71298
rect -2906 -71358 -2900 -71298
rect -2198 -71358 -2192 -71298
rect -2132 -71358 -2126 -71298
rect -2966 -71400 -2906 -71358
rect -2192 -71400 -2132 -71358
rect -2992 -71406 -2884 -71400
rect -2992 -71440 -2980 -71406
rect -2896 -71440 -2884 -71406
rect -2992 -71446 -2884 -71440
rect -2734 -71406 -2626 -71400
rect -2734 -71440 -2722 -71406
rect -2638 -71440 -2626 -71406
rect -2734 -71446 -2626 -71440
rect -2476 -71406 -2368 -71400
rect -2476 -71440 -2464 -71406
rect -2380 -71440 -2368 -71406
rect -2476 -71446 -2368 -71440
rect -2218 -71406 -2110 -71400
rect -2218 -71440 -2206 -71406
rect -2122 -71440 -2110 -71406
rect -2218 -71446 -2110 -71440
rect -3100 -71526 -3084 -71490
rect -3308 -71866 -3302 -71544
rect -3090 -71796 -3084 -71526
rect -3348 -71878 -3302 -71866
rect -3094 -71866 -3084 -71796
rect -3050 -71526 -3040 -71490
rect -2832 -71490 -2786 -71478
rect -3050 -71796 -3044 -71526
rect -3050 -71866 -3034 -71796
rect -2832 -71830 -2826 -71490
rect -3250 -71916 -3142 -71910
rect -3250 -71950 -3238 -71916
rect -3154 -71950 -3142 -71916
rect -3250 -71956 -3142 -71950
rect -3094 -72150 -3034 -71866
rect -2840 -71866 -2826 -71830
rect -2792 -71830 -2786 -71490
rect -2574 -71490 -2528 -71478
rect -2792 -71866 -2780 -71830
rect -2574 -71834 -2568 -71490
rect -2992 -71916 -2884 -71910
rect -2992 -71950 -2980 -71916
rect -2896 -71950 -2884 -71916
rect -2992 -71956 -2884 -71950
rect -2840 -72106 -2780 -71866
rect -2578 -71866 -2568 -71834
rect -2534 -71834 -2528 -71490
rect -2316 -71490 -2270 -71478
rect -2316 -71824 -2310 -71490
rect -2534 -71866 -2518 -71834
rect -2734 -71916 -2626 -71910
rect -2734 -71950 -2722 -71916
rect -2638 -71950 -2626 -71916
rect -2734 -71956 -2626 -71950
rect -2708 -71994 -2648 -71956
rect -2714 -72054 -2708 -71994
rect -2648 -72054 -2642 -71994
rect -3100 -72210 -3094 -72150
rect -3034 -72210 -3028 -72150
rect -2846 -72166 -2840 -72106
rect -2780 -72166 -2774 -72106
rect -3690 -72322 -3578 -72238
rect -8072 -72330 -5354 -72324
rect -8072 -72353 -7584 -72330
rect -8072 -72387 -8043 -72353
rect -8009 -72387 -7951 -72353
rect -7917 -72387 -7859 -72353
rect -7825 -72387 -7584 -72353
rect -8072 -72418 -7584 -72387
rect -11690 -72436 -9354 -72430
rect -7690 -72430 -7584 -72418
rect -5460 -72430 -5354 -72330
rect -4072 -72324 -3578 -72322
rect -2708 -72324 -2648 -72054
rect -2578 -72216 -2518 -71866
rect -2320 -71866 -2310 -71824
rect -2276 -71824 -2270 -71490
rect -2064 -71490 -2004 -71244
rect -1936 -71304 -1876 -71074
rect -1808 -71304 -1748 -71074
rect -1936 -71364 -1748 -71304
rect -1936 -71400 -1876 -71364
rect -1960 -71406 -1852 -71400
rect -1960 -71440 -1948 -71406
rect -1864 -71440 -1852 -71406
rect -1960 -71446 -1852 -71440
rect -2064 -71544 -2052 -71490
rect -2276 -71866 -2260 -71824
rect -2476 -71916 -2368 -71910
rect -2476 -71950 -2464 -71916
rect -2380 -71950 -2368 -71916
rect -2476 -71956 -2368 -71950
rect -2452 -71994 -2392 -71956
rect -2458 -72054 -2452 -71994
rect -2392 -72054 -2386 -71994
rect -2578 -72282 -2518 -72276
rect -2452 -72324 -2392 -72054
rect -2320 -72106 -2260 -71866
rect -2058 -71866 -2052 -71544
rect -2018 -71544 -2004 -71490
rect -1808 -71490 -1748 -71364
rect -1808 -71536 -1794 -71490
rect -2018 -71866 -2012 -71544
rect -2058 -71878 -2012 -71866
rect -1800 -71866 -1794 -71536
rect -1760 -71536 -1748 -71490
rect -1760 -71866 -1754 -71536
rect -1800 -71878 -1754 -71866
rect -2218 -71916 -2110 -71910
rect -2218 -71950 -2206 -71916
rect -2122 -71950 -2110 -71916
rect -2218 -71956 -2110 -71950
rect -1960 -71916 -1852 -71910
rect -1960 -71950 -1948 -71916
rect -1864 -71950 -1852 -71916
rect -1960 -71956 -1852 -71950
rect -2326 -72166 -2320 -72106
rect -2260 -72166 -2254 -72106
rect -1466 -72238 -1460 -70578
rect -1360 -72238 -1354 -70578
rect -1466 -72324 -1354 -72238
rect 310 -70386 2646 -70380
rect 310 -70486 416 -70386
rect 2540 -70486 2646 -70386
rect 310 -70492 2646 -70486
rect 310 -70578 422 -70492
rect 310 -72238 316 -70578
rect 416 -72238 422 -70578
rect 1022 -70792 1032 -70492
rect 1924 -70792 1934 -70492
rect 2534 -70578 2646 -70492
rect 534 -70974 2312 -70944
rect 534 -71042 570 -70974
rect 2278 -71042 2312 -70974
rect 534 -71074 2312 -71042
rect 644 -71310 704 -71074
rect 774 -71310 834 -71074
rect 894 -71244 900 -71184
rect 960 -71244 966 -71184
rect 1930 -71244 1936 -71184
rect 1996 -71244 2002 -71184
rect 644 -71370 834 -71310
rect 644 -71490 704 -71370
rect 774 -71400 834 -71370
rect 750 -71406 858 -71400
rect 750 -71440 762 -71406
rect 846 -71440 858 -71406
rect 750 -71446 858 -71440
rect 644 -71544 658 -71490
rect 652 -71866 658 -71544
rect 692 -71544 704 -71490
rect 900 -71490 960 -71244
rect 1028 -71358 1034 -71298
rect 1094 -71358 1100 -71298
rect 1802 -71358 1808 -71298
rect 1868 -71358 1874 -71298
rect 1034 -71400 1094 -71358
rect 1808 -71400 1868 -71358
rect 1008 -71406 1116 -71400
rect 1008 -71440 1020 -71406
rect 1104 -71440 1116 -71406
rect 1008 -71446 1116 -71440
rect 1266 -71406 1374 -71400
rect 1266 -71440 1278 -71406
rect 1362 -71440 1374 -71406
rect 1266 -71446 1374 -71440
rect 1524 -71406 1632 -71400
rect 1524 -71440 1536 -71406
rect 1620 -71440 1632 -71406
rect 1524 -71446 1632 -71440
rect 1782 -71406 1890 -71400
rect 1782 -71440 1794 -71406
rect 1878 -71440 1890 -71406
rect 1782 -71446 1890 -71440
rect 900 -71526 916 -71490
rect 692 -71866 698 -71544
rect 910 -71796 916 -71526
rect 652 -71878 698 -71866
rect 906 -71866 916 -71796
rect 950 -71526 960 -71490
rect 1168 -71490 1214 -71478
rect 950 -71796 956 -71526
rect 950 -71866 966 -71796
rect 1168 -71830 1174 -71490
rect 750 -71916 858 -71910
rect 750 -71950 762 -71916
rect 846 -71950 858 -71916
rect 750 -71956 858 -71950
rect 906 -72150 966 -71866
rect 1160 -71866 1174 -71830
rect 1208 -71830 1214 -71490
rect 1426 -71490 1472 -71478
rect 1208 -71866 1220 -71830
rect 1426 -71834 1432 -71490
rect 1008 -71916 1116 -71910
rect 1008 -71950 1020 -71916
rect 1104 -71950 1116 -71916
rect 1008 -71956 1116 -71950
rect 1160 -72106 1220 -71866
rect 1422 -71866 1432 -71834
rect 1466 -71834 1472 -71490
rect 1684 -71490 1730 -71478
rect 1684 -71824 1690 -71490
rect 1466 -71866 1482 -71834
rect 1266 -71916 1374 -71910
rect 1266 -71950 1278 -71916
rect 1362 -71950 1374 -71916
rect 1266 -71956 1374 -71950
rect 1292 -71994 1352 -71956
rect 1286 -72054 1292 -71994
rect 1352 -72054 1358 -71994
rect 900 -72210 906 -72150
rect 966 -72210 972 -72150
rect 1154 -72166 1160 -72106
rect 1220 -72166 1226 -72106
rect 310 -72322 422 -72238
rect 1422 -72216 1482 -71866
rect 1680 -71866 1690 -71824
rect 1724 -71824 1730 -71490
rect 1936 -71490 1996 -71244
rect 2064 -71304 2124 -71074
rect 2192 -71304 2252 -71074
rect 2064 -71364 2252 -71304
rect 2064 -71400 2124 -71364
rect 2040 -71406 2148 -71400
rect 2040 -71440 2052 -71406
rect 2136 -71440 2148 -71406
rect 2040 -71446 2148 -71440
rect 1936 -71544 1948 -71490
rect 1724 -71866 1740 -71824
rect 1524 -71916 1632 -71910
rect 1524 -71950 1536 -71916
rect 1620 -71950 1632 -71916
rect 1524 -71956 1632 -71950
rect 1548 -71994 1608 -71956
rect 1542 -72054 1548 -71994
rect 1608 -72054 1614 -71994
rect 1680 -72106 1740 -71866
rect 1942 -71866 1948 -71544
rect 1982 -71544 1996 -71490
rect 2192 -71490 2252 -71364
rect 2192 -71536 2206 -71490
rect 1982 -71866 1988 -71544
rect 1942 -71878 1988 -71866
rect 2200 -71866 2206 -71536
rect 2240 -71536 2252 -71490
rect 2240 -71866 2246 -71536
rect 2200 -71878 2246 -71866
rect 1782 -71916 1890 -71910
rect 1782 -71950 1794 -71916
rect 1878 -71950 1890 -71916
rect 1782 -71956 1890 -71950
rect 2040 -71916 2148 -71910
rect 2040 -71950 2052 -71916
rect 2136 -71950 2148 -71916
rect 2040 -71956 2148 -71950
rect 1674 -72166 1680 -72106
rect 1740 -72166 1746 -72106
rect 1422 -72282 1482 -72276
rect 2534 -72238 2540 -70578
rect 2640 -72238 2646 -70578
rect -4072 -72330 -1354 -72324
rect -4072 -72353 -3584 -72330
rect -4072 -72387 -4043 -72353
rect -4009 -72387 -3951 -72353
rect -3917 -72387 -3859 -72353
rect -3825 -72387 -3584 -72353
rect -4072 -72418 -3584 -72387
rect -7690 -72436 -5354 -72430
rect -3690 -72430 -3584 -72418
rect -1460 -72430 -1354 -72330
rect -72 -72324 422 -72322
rect 2534 -72324 2646 -72238
rect 4310 -70386 6646 -70380
rect 4310 -70486 4416 -70386
rect 6540 -70486 6646 -70386
rect 4310 -70492 6646 -70486
rect 4310 -70578 4422 -70492
rect 4310 -72238 4316 -70578
rect 4416 -72238 4422 -70578
rect 5022 -70792 5032 -70492
rect 5924 -70792 5934 -70492
rect 6534 -70578 6646 -70492
rect 4534 -70974 6312 -70944
rect 4534 -71042 4570 -70974
rect 6278 -71042 6312 -70974
rect 4534 -71074 6312 -71042
rect 4644 -71310 4704 -71074
rect 4774 -71310 4834 -71074
rect 4894 -71244 4900 -71184
rect 4960 -71244 4966 -71184
rect 5930 -71244 5936 -71184
rect 5996 -71244 6002 -71184
rect 4644 -71370 4834 -71310
rect 4644 -71490 4704 -71370
rect 4774 -71400 4834 -71370
rect 4750 -71406 4858 -71400
rect 4750 -71440 4762 -71406
rect 4846 -71440 4858 -71406
rect 4750 -71446 4858 -71440
rect 4644 -71544 4658 -71490
rect 4652 -71866 4658 -71544
rect 4692 -71544 4704 -71490
rect 4900 -71490 4960 -71244
rect 5028 -71358 5034 -71298
rect 5094 -71358 5100 -71298
rect 5802 -71358 5808 -71298
rect 5868 -71358 5874 -71298
rect 5034 -71400 5094 -71358
rect 5808 -71400 5868 -71358
rect 5008 -71406 5116 -71400
rect 5008 -71440 5020 -71406
rect 5104 -71440 5116 -71406
rect 5008 -71446 5116 -71440
rect 5266 -71406 5374 -71400
rect 5266 -71440 5278 -71406
rect 5362 -71440 5374 -71406
rect 5266 -71446 5374 -71440
rect 5524 -71406 5632 -71400
rect 5524 -71440 5536 -71406
rect 5620 -71440 5632 -71406
rect 5524 -71446 5632 -71440
rect 5782 -71406 5890 -71400
rect 5782 -71440 5794 -71406
rect 5878 -71440 5890 -71406
rect 5782 -71446 5890 -71440
rect 4900 -71526 4916 -71490
rect 4692 -71866 4698 -71544
rect 4910 -71796 4916 -71526
rect 4652 -71878 4698 -71866
rect 4906 -71866 4916 -71796
rect 4950 -71526 4960 -71490
rect 5168 -71490 5214 -71478
rect 4950 -71796 4956 -71526
rect 4950 -71866 4966 -71796
rect 5168 -71830 5174 -71490
rect 4750 -71916 4858 -71910
rect 4750 -71950 4762 -71916
rect 4846 -71950 4858 -71916
rect 4750 -71956 4858 -71950
rect 4906 -72150 4966 -71866
rect 5160 -71866 5174 -71830
rect 5208 -71830 5214 -71490
rect 5426 -71490 5472 -71478
rect 5208 -71866 5220 -71830
rect 5426 -71834 5432 -71490
rect 5008 -71916 5116 -71910
rect 5008 -71950 5020 -71916
rect 5104 -71950 5116 -71916
rect 5008 -71956 5116 -71950
rect 5160 -72106 5220 -71866
rect 5422 -71866 5432 -71834
rect 5466 -71834 5472 -71490
rect 5684 -71490 5730 -71478
rect 5684 -71824 5690 -71490
rect 5466 -71866 5482 -71834
rect 5266 -71916 5374 -71910
rect 5266 -71950 5278 -71916
rect 5362 -71950 5374 -71916
rect 5266 -71956 5374 -71950
rect 5292 -71994 5352 -71956
rect 5286 -72054 5292 -71994
rect 5352 -72054 5358 -71994
rect 4900 -72210 4906 -72150
rect 4966 -72210 4972 -72150
rect 5154 -72166 5160 -72106
rect 5220 -72166 5226 -72106
rect 4310 -72322 4422 -72238
rect 5422 -72216 5482 -71866
rect 5680 -71866 5690 -71824
rect 5724 -71824 5730 -71490
rect 5936 -71490 5996 -71244
rect 6064 -71304 6124 -71074
rect 6192 -71304 6252 -71074
rect 6064 -71364 6252 -71304
rect 6064 -71400 6124 -71364
rect 6040 -71406 6148 -71400
rect 6040 -71440 6052 -71406
rect 6136 -71440 6148 -71406
rect 6040 -71446 6148 -71440
rect 5936 -71544 5948 -71490
rect 5724 -71866 5740 -71824
rect 5524 -71916 5632 -71910
rect 5524 -71950 5536 -71916
rect 5620 -71950 5632 -71916
rect 5524 -71956 5632 -71950
rect 5548 -71994 5608 -71956
rect 5542 -72054 5548 -71994
rect 5608 -72054 5614 -71994
rect 5680 -72106 5740 -71866
rect 5942 -71866 5948 -71544
rect 5982 -71544 5996 -71490
rect 6192 -71490 6252 -71364
rect 6192 -71536 6206 -71490
rect 5982 -71866 5988 -71544
rect 5942 -71878 5988 -71866
rect 6200 -71866 6206 -71536
rect 6240 -71536 6252 -71490
rect 6240 -71866 6246 -71536
rect 6200 -71878 6246 -71866
rect 5782 -71916 5890 -71910
rect 5782 -71950 5794 -71916
rect 5878 -71950 5890 -71916
rect 5782 -71956 5890 -71950
rect 6040 -71916 6148 -71910
rect 6040 -71950 6052 -71916
rect 6136 -71950 6148 -71916
rect 6040 -71956 6148 -71950
rect 5674 -72166 5680 -72106
rect 5740 -72166 5746 -72106
rect 5422 -72282 5482 -72276
rect 6534 -72238 6540 -70578
rect 6640 -72238 6646 -70578
rect -72 -72330 2646 -72324
rect -72 -72353 416 -72330
rect -72 -72387 -43 -72353
rect -9 -72387 49 -72353
rect 83 -72387 141 -72353
rect 175 -72387 416 -72353
rect -72 -72418 416 -72387
rect -3690 -72436 -1354 -72430
rect 310 -72430 416 -72418
rect 2540 -72430 2646 -72330
rect 3928 -72324 4422 -72322
rect 6534 -72324 6646 -72238
rect 3928 -72330 6646 -72324
rect 3928 -72353 4416 -72330
rect 3928 -72387 3957 -72353
rect 3991 -72387 4049 -72353
rect 4083 -72387 4141 -72353
rect 4175 -72387 4416 -72353
rect 3928 -72418 4416 -72387
rect 310 -72436 2646 -72430
rect 4310 -72430 4416 -72418
rect 6540 -72430 6646 -72330
rect 4310 -72436 6646 -72430
rect -27908 -72522 -27848 -72516
rect -23908 -72522 -23848 -72516
rect -19908 -72522 -19848 -72516
rect -15908 -72522 -15848 -72516
rect -11908 -72522 -11848 -72516
rect -7908 -72522 -7848 -72516
rect -3908 -72522 -3848 -72516
rect 92 -72522 152 -72516
rect 4092 -72522 4152 -72516
rect -28230 -72580 -28170 -72574
rect -28374 -72640 -28230 -72580
rect -28170 -72586 -27944 -72580
rect -27914 -72582 -27908 -72522
rect -27848 -72582 -27842 -72522
rect -24230 -72580 -24170 -72574
rect -28170 -72634 -28004 -72586
rect -27956 -72634 -27944 -72586
rect -27908 -72588 -27848 -72582
rect -28170 -72640 -27944 -72634
rect -24360 -72640 -24230 -72580
rect -24170 -72586 -23944 -72580
rect -23914 -72582 -23908 -72522
rect -23848 -72582 -23842 -72522
rect -20230 -72580 -20170 -72574
rect -24170 -72634 -24004 -72586
rect -23956 -72634 -23944 -72586
rect -23908 -72588 -23848 -72582
rect -24170 -72640 -23944 -72634
rect -20376 -72640 -20230 -72580
rect -20170 -72586 -19944 -72580
rect -19914 -72582 -19908 -72522
rect -19848 -72582 -19842 -72522
rect -16230 -72580 -16170 -72574
rect -20170 -72634 -20004 -72586
rect -19956 -72634 -19944 -72586
rect -19908 -72588 -19848 -72582
rect -20170 -72640 -19944 -72634
rect -16390 -72640 -16230 -72580
rect -16170 -72586 -15944 -72580
rect -15914 -72582 -15908 -72522
rect -15848 -72582 -15842 -72522
rect -12230 -72580 -12170 -72574
rect -16170 -72634 -16004 -72586
rect -15956 -72634 -15944 -72586
rect -15908 -72588 -15848 -72582
rect -16170 -72640 -15944 -72634
rect -12428 -72640 -12230 -72580
rect -12170 -72586 -11944 -72580
rect -11914 -72582 -11908 -72522
rect -11848 -72582 -11842 -72522
rect -8230 -72580 -8170 -72574
rect -12170 -72634 -12004 -72586
rect -11956 -72634 -11944 -72586
rect -11908 -72588 -11848 -72582
rect -12170 -72640 -11944 -72634
rect -8402 -72640 -8230 -72580
rect -8170 -72586 -7944 -72580
rect -7914 -72582 -7908 -72522
rect -7848 -72582 -7842 -72522
rect -4230 -72580 -4170 -72574
rect -8170 -72634 -8004 -72586
rect -7956 -72634 -7944 -72586
rect -7908 -72588 -7848 -72582
rect -8170 -72640 -7944 -72634
rect -4170 -72586 -3944 -72580
rect -3914 -72582 -3908 -72522
rect -3848 -72582 -3842 -72522
rect -230 -72580 -170 -72574
rect -4170 -72634 -4004 -72586
rect -3956 -72634 -3944 -72586
rect -3908 -72588 -3848 -72582
rect -4170 -72640 -3944 -72634
rect -392 -72640 -230 -72580
rect -170 -72586 56 -72580
rect 86 -72582 92 -72522
rect 152 -72582 158 -72522
rect 3770 -72580 3830 -72574
rect -170 -72634 -4 -72586
rect 44 -72634 56 -72586
rect 92 -72588 152 -72582
rect -170 -72640 56 -72634
rect 3606 -72640 3770 -72580
rect 3830 -72586 4056 -72580
rect 4086 -72582 4092 -72522
rect 4152 -72582 4158 -72522
rect 3830 -72634 3996 -72586
rect 4044 -72634 4056 -72586
rect 4092 -72588 4152 -72582
rect 3830 -72640 4056 -72634
rect -28230 -72646 -28170 -72640
rect -24230 -72646 -24170 -72640
rect -20230 -72646 -20170 -72640
rect -16230 -72646 -16170 -72640
rect -12230 -72646 -12170 -72640
rect -8230 -72646 -8170 -72640
rect -4230 -72646 -4170 -72640
rect -230 -72646 -170 -72640
rect 3770 -72646 3830 -72640
rect -27690 -72666 -25354 -72660
rect -27690 -72766 -27584 -72666
rect -25460 -72766 -25354 -72666
rect -27690 -72772 -25354 -72766
rect -27690 -72866 -27578 -72772
rect -28072 -72897 -27578 -72866
rect -28072 -72931 -28043 -72897
rect -28009 -72931 -27951 -72897
rect -27917 -72931 -27859 -72897
rect -27825 -72906 -27578 -72897
rect -27825 -72931 -27684 -72906
rect -28072 -72962 -27684 -72931
rect -27690 -75530 -27684 -72962
rect -27584 -75530 -27578 -72906
rect -26584 -72916 -26578 -72856
rect -26518 -72916 -26512 -72856
rect -27100 -73064 -27094 -73004
rect -27034 -73064 -27028 -73004
rect -27496 -73176 -27246 -73116
rect -27186 -73176 -27180 -73116
rect -27496 -74096 -27436 -73176
rect -27245 -73230 -27137 -73224
rect -27245 -73264 -27233 -73230
rect -27149 -73264 -27137 -73230
rect -27245 -73270 -27137 -73264
rect -27343 -73323 -27297 -73311
rect -27343 -73646 -27337 -73323
rect -27496 -74690 -27436 -74156
rect -27348 -73699 -27337 -73646
rect -27303 -73646 -27297 -73323
rect -27094 -73323 -27034 -73064
rect -26968 -73176 -26962 -73116
rect -26902 -73176 -26896 -73116
rect -26962 -73224 -26902 -73176
rect -26987 -73230 -26879 -73224
rect -26987 -73264 -26975 -73230
rect -26891 -73264 -26879 -73230
rect -26987 -73270 -26879 -73264
rect -26729 -73230 -26621 -73224
rect -26729 -73264 -26717 -73230
rect -26633 -73264 -26621 -73230
rect -26729 -73270 -26621 -73264
rect -27094 -73368 -27079 -73323
rect -27303 -73699 -27288 -73646
rect -27348 -73900 -27288 -73699
rect -27085 -73699 -27079 -73368
rect -27045 -73368 -27034 -73323
rect -26827 -73323 -26781 -73311
rect -26827 -73360 -26821 -73323
rect -27045 -73699 -27039 -73368
rect -27085 -73711 -27039 -73699
rect -26834 -73699 -26821 -73360
rect -26787 -73360 -26781 -73323
rect -26578 -73323 -26518 -72916
rect -26326 -72956 -26320 -72896
rect -26260 -72956 -26254 -72896
rect -26450 -73224 -26390 -73170
rect -26471 -73230 -26363 -73224
rect -26471 -73264 -26459 -73230
rect -26375 -73264 -26363 -73230
rect -26471 -73270 -26363 -73264
rect -26787 -73699 -26774 -73360
rect -26578 -73362 -26563 -73323
rect -26569 -73666 -26563 -73362
rect -27245 -73758 -27137 -73752
rect -27245 -73792 -27233 -73758
rect -27149 -73792 -27137 -73758
rect -27245 -73798 -27137 -73792
rect -26987 -73758 -26879 -73752
rect -26987 -73792 -26975 -73758
rect -26891 -73792 -26879 -73758
rect -26987 -73798 -26879 -73792
rect -27218 -73900 -27158 -73798
rect -27348 -73960 -27158 -73900
rect -27098 -73912 -27092 -73852
rect -27032 -73912 -27026 -73852
rect -27348 -74183 -27288 -73960
rect -27218 -74084 -27158 -73960
rect -27245 -74090 -27137 -74084
rect -27245 -74124 -27233 -74090
rect -27149 -74124 -27137 -74090
rect -27245 -74130 -27137 -74124
rect -27348 -74226 -27337 -74183
rect -27343 -74526 -27337 -74226
rect -27348 -74559 -27337 -74526
rect -27303 -74226 -27288 -74183
rect -27092 -74183 -27032 -73912
rect -26968 -74026 -26962 -73966
rect -26902 -74026 -26896 -73966
rect -26962 -74084 -26902 -74026
rect -26987 -74090 -26879 -74084
rect -26987 -74124 -26975 -74090
rect -26891 -74124 -26879 -74090
rect -26987 -74130 -26879 -74124
rect -27303 -74526 -27297 -74226
rect -27303 -74559 -27288 -74526
rect -27502 -74750 -27496 -74690
rect -27436 -74750 -27430 -74690
rect -27348 -74742 -27288 -74559
rect -27092 -74559 -27079 -74183
rect -27045 -74559 -27032 -74183
rect -27245 -74618 -27137 -74612
rect -27245 -74652 -27233 -74618
rect -27149 -74652 -27137 -74618
rect -27245 -74658 -27137 -74652
rect -27218 -74742 -27158 -74658
rect -27348 -74802 -27158 -74742
rect -27348 -75066 -27288 -74802
rect -27218 -75066 -27158 -74802
rect -27092 -74870 -27032 -74559
rect -26834 -74183 -26774 -73699
rect -26574 -73699 -26563 -73666
rect -26529 -73362 -26518 -73323
rect -26320 -73323 -26260 -72956
rect -26064 -73064 -26058 -73004
rect -25998 -73064 -25992 -73004
rect -26192 -73176 -26186 -73116
rect -26126 -73176 -26120 -73116
rect -26186 -73224 -26126 -73176
rect -26213 -73230 -26105 -73224
rect -26213 -73264 -26201 -73230
rect -26117 -73264 -26105 -73230
rect -26213 -73270 -26105 -73264
rect -26529 -73666 -26523 -73362
rect -26320 -73376 -26305 -73323
rect -26311 -73654 -26305 -73376
rect -26529 -73699 -26514 -73666
rect -26729 -73758 -26621 -73752
rect -26729 -73792 -26717 -73758
rect -26633 -73792 -26621 -73758
rect -26729 -73798 -26621 -73792
rect -26704 -73966 -26644 -73798
rect -26574 -73852 -26514 -73699
rect -26322 -73699 -26305 -73654
rect -26271 -73376 -26260 -73323
rect -26058 -73323 -25998 -73064
rect -25934 -73118 -25874 -72772
rect -25800 -73118 -25740 -72772
rect -25466 -72906 -25354 -72772
rect -23690 -72666 -21354 -72660
rect -23690 -72766 -23584 -72666
rect -21460 -72766 -21354 -72666
rect -23690 -72772 -21354 -72766
rect -23690 -72866 -23578 -72772
rect -25654 -73064 -25648 -73004
rect -25588 -73064 -25582 -73004
rect -25934 -73178 -25740 -73118
rect -25934 -73224 -25874 -73178
rect -25955 -73230 -25847 -73224
rect -25955 -73264 -25943 -73230
rect -25859 -73264 -25847 -73230
rect -25955 -73270 -25847 -73264
rect -26271 -73654 -26265 -73376
rect -26058 -73400 -26047 -73323
rect -26271 -73699 -26262 -73654
rect -26471 -73758 -26363 -73752
rect -26471 -73792 -26459 -73758
rect -26375 -73792 -26363 -73758
rect -26471 -73798 -26363 -73792
rect -26580 -73912 -26574 -73852
rect -26514 -73912 -26508 -73852
rect -26446 -73966 -26386 -73798
rect -26710 -74026 -26704 -73966
rect -26644 -74026 -26638 -73966
rect -26452 -74026 -26446 -73966
rect -26386 -74026 -26380 -73966
rect -26729 -74090 -26621 -74084
rect -26729 -74124 -26717 -74090
rect -26633 -74124 -26621 -74090
rect -26729 -74130 -26621 -74124
rect -26471 -74090 -26363 -74084
rect -26471 -74124 -26459 -74090
rect -26375 -74124 -26363 -74090
rect -26471 -74130 -26363 -74124
rect -26834 -74559 -26821 -74183
rect -26787 -74559 -26774 -74183
rect -26569 -74183 -26523 -74171
rect -26569 -74526 -26563 -74183
rect -26987 -74618 -26879 -74612
rect -26987 -74652 -26975 -74618
rect -26891 -74652 -26879 -74618
rect -26987 -74658 -26879 -74652
rect -27098 -74930 -27092 -74870
rect -27032 -74930 -27026 -74870
rect -26834 -74922 -26774 -74559
rect -26578 -74559 -26563 -74526
rect -26529 -74526 -26523 -74183
rect -26322 -74183 -26262 -73699
rect -26053 -73699 -26047 -73400
rect -26013 -73400 -25998 -73323
rect -25800 -73323 -25740 -73178
rect -26013 -73699 -26007 -73400
rect -26053 -73711 -26007 -73699
rect -25800 -73699 -25789 -73323
rect -25755 -73699 -25740 -73323
rect -26213 -73758 -26105 -73752
rect -26213 -73792 -26201 -73758
rect -26117 -73792 -26105 -73758
rect -26213 -73798 -26105 -73792
rect -25955 -73758 -25847 -73752
rect -25955 -73792 -25943 -73758
rect -25859 -73792 -25847 -73758
rect -25955 -73798 -25847 -73792
rect -26064 -73912 -26058 -73852
rect -25998 -73912 -25992 -73852
rect -25932 -73908 -25872 -73798
rect -25800 -73908 -25740 -73699
rect -26194 -74026 -26188 -73966
rect -26128 -74026 -26122 -73966
rect -26188 -74084 -26128 -74026
rect -26213 -74090 -26105 -74084
rect -26213 -74124 -26201 -74090
rect -26117 -74124 -26105 -74090
rect -26213 -74130 -26105 -74124
rect -26322 -74240 -26305 -74183
rect -26311 -74498 -26305 -74240
rect -26529 -74559 -26518 -74526
rect -26729 -74618 -26621 -74612
rect -26729 -74652 -26717 -74618
rect -26633 -74652 -26621 -74618
rect -26729 -74658 -26621 -74652
rect -26706 -74690 -26646 -74658
rect -26712 -74750 -26706 -74690
rect -26646 -74750 -26640 -74690
rect -26578 -74810 -26518 -74559
rect -26316 -74559 -26305 -74498
rect -26271 -74240 -26262 -74183
rect -26058 -74183 -25998 -73912
rect -25932 -73968 -25740 -73908
rect -25955 -74090 -25847 -74084
rect -25955 -74124 -25943 -74090
rect -25859 -74124 -25847 -74090
rect -25955 -74130 -25847 -74124
rect -26058 -74232 -26047 -74183
rect -26271 -74498 -26265 -74240
rect -26271 -74559 -26256 -74498
rect -26471 -74618 -26363 -74612
rect -26471 -74652 -26459 -74618
rect -26375 -74652 -26363 -74618
rect -26471 -74658 -26363 -74652
rect -26450 -74690 -26390 -74658
rect -26456 -74750 -26450 -74690
rect -26390 -74750 -26384 -74690
rect -26584 -74870 -26578 -74810
rect -26518 -74870 -26512 -74810
rect -26316 -74922 -26256 -74559
rect -26053 -74559 -26047 -74232
rect -26013 -74232 -25998 -74183
rect -25800 -74183 -25740 -73968
rect -26013 -74559 -26007 -74232
rect -26053 -74571 -26007 -74559
rect -25800 -74559 -25789 -74183
rect -25755 -74559 -25740 -74183
rect -26213 -74618 -26105 -74612
rect -26213 -74652 -26201 -74618
rect -26117 -74652 -26105 -74618
rect -26213 -74658 -26105 -74652
rect -25955 -74618 -25847 -74612
rect -25955 -74652 -25943 -74618
rect -25859 -74652 -25847 -74618
rect -25955 -74658 -25847 -74652
rect -25928 -74730 -25868 -74658
rect -25800 -74730 -25740 -74559
rect -25928 -74790 -25740 -74730
rect -26840 -74982 -26834 -74922
rect -26774 -74982 -26768 -74922
rect -26322 -74982 -26316 -74922
rect -26256 -74982 -26250 -74922
rect -25928 -75066 -25868 -74790
rect -25800 -75066 -25740 -74790
rect -25648 -74810 -25588 -73064
rect -25654 -74870 -25648 -74810
rect -25588 -74870 -25582 -74810
rect -27422 -75096 -25520 -75066
rect -27422 -75160 -27388 -75096
rect -25564 -75160 -25520 -75096
rect -27422 -75190 -25520 -75160
rect -27690 -75664 -27578 -75530
rect -26978 -75664 -26968 -75364
rect -26076 -75664 -26066 -75364
rect -25466 -75530 -25460 -72906
rect -25360 -75530 -25354 -72906
rect -24072 -72897 -23578 -72866
rect -24072 -72931 -24043 -72897
rect -24009 -72931 -23951 -72897
rect -23917 -72931 -23859 -72897
rect -23825 -72906 -23578 -72897
rect -23825 -72931 -23684 -72906
rect -24072 -72962 -23684 -72931
rect -25466 -75664 -25354 -75530
rect -27690 -75670 -25354 -75664
rect -27690 -75770 -27584 -75670
rect -25460 -75770 -25354 -75670
rect -27690 -75776 -25354 -75770
rect -23690 -75530 -23684 -72962
rect -23584 -75530 -23578 -72906
rect -22584 -72916 -22578 -72856
rect -22518 -72916 -22512 -72856
rect -23100 -73064 -23094 -73004
rect -23034 -73064 -23028 -73004
rect -23496 -73176 -23246 -73116
rect -23186 -73176 -23180 -73116
rect -23496 -74096 -23436 -73176
rect -23245 -73230 -23137 -73224
rect -23245 -73264 -23233 -73230
rect -23149 -73264 -23137 -73230
rect -23245 -73270 -23137 -73264
rect -23343 -73323 -23297 -73311
rect -23343 -73646 -23337 -73323
rect -23496 -74690 -23436 -74156
rect -23348 -73699 -23337 -73646
rect -23303 -73646 -23297 -73323
rect -23094 -73323 -23034 -73064
rect -22968 -73176 -22962 -73116
rect -22902 -73176 -22896 -73116
rect -22962 -73224 -22902 -73176
rect -22987 -73230 -22879 -73224
rect -22987 -73264 -22975 -73230
rect -22891 -73264 -22879 -73230
rect -22987 -73270 -22879 -73264
rect -22729 -73230 -22621 -73224
rect -22729 -73264 -22717 -73230
rect -22633 -73264 -22621 -73230
rect -22729 -73270 -22621 -73264
rect -23094 -73368 -23079 -73323
rect -23303 -73699 -23288 -73646
rect -23348 -73900 -23288 -73699
rect -23085 -73699 -23079 -73368
rect -23045 -73368 -23034 -73323
rect -22827 -73323 -22781 -73311
rect -22827 -73360 -22821 -73323
rect -23045 -73699 -23039 -73368
rect -23085 -73711 -23039 -73699
rect -22834 -73699 -22821 -73360
rect -22787 -73360 -22781 -73323
rect -22578 -73323 -22518 -72916
rect -22326 -72956 -22320 -72896
rect -22260 -72956 -22254 -72896
rect -22450 -73224 -22390 -73170
rect -22471 -73230 -22363 -73224
rect -22471 -73264 -22459 -73230
rect -22375 -73264 -22363 -73230
rect -22471 -73270 -22363 -73264
rect -22787 -73699 -22774 -73360
rect -22578 -73362 -22563 -73323
rect -22569 -73666 -22563 -73362
rect -23245 -73758 -23137 -73752
rect -23245 -73792 -23233 -73758
rect -23149 -73792 -23137 -73758
rect -23245 -73798 -23137 -73792
rect -22987 -73758 -22879 -73752
rect -22987 -73792 -22975 -73758
rect -22891 -73792 -22879 -73758
rect -22987 -73798 -22879 -73792
rect -23218 -73900 -23158 -73798
rect -23348 -73960 -23158 -73900
rect -23098 -73912 -23092 -73852
rect -23032 -73912 -23026 -73852
rect -23348 -74183 -23288 -73960
rect -23218 -74084 -23158 -73960
rect -23245 -74090 -23137 -74084
rect -23245 -74124 -23233 -74090
rect -23149 -74124 -23137 -74090
rect -23245 -74130 -23137 -74124
rect -23348 -74226 -23337 -74183
rect -23343 -74526 -23337 -74226
rect -23348 -74559 -23337 -74526
rect -23303 -74226 -23288 -74183
rect -23092 -74183 -23032 -73912
rect -22968 -74026 -22962 -73966
rect -22902 -74026 -22896 -73966
rect -22962 -74084 -22902 -74026
rect -22987 -74090 -22879 -74084
rect -22987 -74124 -22975 -74090
rect -22891 -74124 -22879 -74090
rect -22987 -74130 -22879 -74124
rect -23303 -74526 -23297 -74226
rect -23303 -74559 -23288 -74526
rect -23502 -74750 -23496 -74690
rect -23436 -74750 -23430 -74690
rect -23348 -74742 -23288 -74559
rect -23092 -74559 -23079 -74183
rect -23045 -74559 -23032 -74183
rect -23245 -74618 -23137 -74612
rect -23245 -74652 -23233 -74618
rect -23149 -74652 -23137 -74618
rect -23245 -74658 -23137 -74652
rect -23218 -74742 -23158 -74658
rect -23348 -74802 -23158 -74742
rect -23348 -75066 -23288 -74802
rect -23218 -75066 -23158 -74802
rect -23092 -74868 -23032 -74559
rect -22834 -74183 -22774 -73699
rect -22574 -73699 -22563 -73666
rect -22529 -73362 -22518 -73323
rect -22320 -73323 -22260 -72956
rect -22064 -73064 -22058 -73004
rect -21998 -73064 -21992 -73004
rect -22192 -73176 -22186 -73116
rect -22126 -73176 -22120 -73116
rect -22186 -73224 -22126 -73176
rect -22213 -73230 -22105 -73224
rect -22213 -73264 -22201 -73230
rect -22117 -73264 -22105 -73230
rect -22213 -73270 -22105 -73264
rect -22529 -73666 -22523 -73362
rect -22320 -73376 -22305 -73323
rect -22311 -73654 -22305 -73376
rect -22529 -73699 -22514 -73666
rect -22729 -73758 -22621 -73752
rect -22729 -73792 -22717 -73758
rect -22633 -73792 -22621 -73758
rect -22729 -73798 -22621 -73792
rect -22704 -73966 -22644 -73798
rect -22574 -73852 -22514 -73699
rect -22322 -73699 -22305 -73654
rect -22271 -73376 -22260 -73323
rect -22058 -73323 -21998 -73064
rect -21934 -73118 -21874 -72772
rect -21800 -73118 -21740 -72772
rect -21466 -72906 -21354 -72772
rect -19690 -72666 -17354 -72660
rect -19690 -72766 -19584 -72666
rect -17460 -72766 -17354 -72666
rect -19690 -72772 -17354 -72766
rect -19690 -72866 -19578 -72772
rect -21654 -73064 -21648 -73004
rect -21588 -73064 -21582 -73004
rect -21934 -73178 -21740 -73118
rect -21934 -73224 -21874 -73178
rect -21955 -73230 -21847 -73224
rect -21955 -73264 -21943 -73230
rect -21859 -73264 -21847 -73230
rect -21955 -73270 -21847 -73264
rect -22271 -73654 -22265 -73376
rect -22058 -73400 -22047 -73323
rect -22271 -73699 -22262 -73654
rect -22471 -73758 -22363 -73752
rect -22471 -73792 -22459 -73758
rect -22375 -73792 -22363 -73758
rect -22471 -73798 -22363 -73792
rect -22580 -73912 -22574 -73852
rect -22514 -73912 -22508 -73852
rect -22446 -73966 -22386 -73798
rect -22710 -74026 -22704 -73966
rect -22644 -74026 -22638 -73966
rect -22452 -74026 -22446 -73966
rect -22386 -74026 -22380 -73966
rect -22729 -74090 -22621 -74084
rect -22729 -74124 -22717 -74090
rect -22633 -74124 -22621 -74090
rect -22729 -74130 -22621 -74124
rect -22471 -74090 -22363 -74084
rect -22471 -74124 -22459 -74090
rect -22375 -74124 -22363 -74090
rect -22471 -74130 -22363 -74124
rect -22834 -74559 -22821 -74183
rect -22787 -74559 -22774 -74183
rect -22569 -74183 -22523 -74171
rect -22569 -74526 -22563 -74183
rect -22987 -74618 -22879 -74612
rect -22987 -74652 -22975 -74618
rect -22891 -74652 -22879 -74618
rect -22987 -74658 -22879 -74652
rect -23098 -74928 -23092 -74868
rect -23032 -74928 -23026 -74868
rect -22834 -74922 -22774 -74559
rect -22578 -74559 -22563 -74526
rect -22529 -74526 -22523 -74183
rect -22322 -74183 -22262 -73699
rect -22053 -73699 -22047 -73400
rect -22013 -73400 -21998 -73323
rect -21800 -73323 -21740 -73178
rect -22013 -73699 -22007 -73400
rect -22053 -73711 -22007 -73699
rect -21800 -73699 -21789 -73323
rect -21755 -73699 -21740 -73323
rect -22213 -73758 -22105 -73752
rect -22213 -73792 -22201 -73758
rect -22117 -73792 -22105 -73758
rect -22213 -73798 -22105 -73792
rect -21955 -73758 -21847 -73752
rect -21955 -73792 -21943 -73758
rect -21859 -73792 -21847 -73758
rect -21955 -73798 -21847 -73792
rect -22064 -73912 -22058 -73852
rect -21998 -73912 -21992 -73852
rect -21932 -73908 -21872 -73798
rect -21800 -73908 -21740 -73699
rect -22194 -74026 -22188 -73966
rect -22128 -74026 -22122 -73966
rect -22188 -74084 -22128 -74026
rect -22213 -74090 -22105 -74084
rect -22213 -74124 -22201 -74090
rect -22117 -74124 -22105 -74090
rect -22213 -74130 -22105 -74124
rect -22322 -74240 -22305 -74183
rect -22311 -74498 -22305 -74240
rect -22529 -74559 -22518 -74526
rect -22729 -74618 -22621 -74612
rect -22729 -74652 -22717 -74618
rect -22633 -74652 -22621 -74618
rect -22729 -74658 -22621 -74652
rect -22706 -74690 -22646 -74658
rect -22712 -74750 -22706 -74690
rect -22646 -74750 -22640 -74690
rect -22578 -74810 -22518 -74559
rect -22316 -74559 -22305 -74498
rect -22271 -74240 -22262 -74183
rect -22058 -74183 -21998 -73912
rect -21932 -73968 -21740 -73908
rect -21955 -74090 -21847 -74084
rect -21955 -74124 -21943 -74090
rect -21859 -74124 -21847 -74090
rect -21955 -74130 -21847 -74124
rect -22058 -74232 -22047 -74183
rect -22271 -74498 -22265 -74240
rect -22271 -74559 -22256 -74498
rect -22471 -74618 -22363 -74612
rect -22471 -74652 -22459 -74618
rect -22375 -74652 -22363 -74618
rect -22471 -74658 -22363 -74652
rect -22450 -74690 -22390 -74658
rect -22456 -74750 -22450 -74690
rect -22390 -74750 -22384 -74690
rect -22584 -74870 -22578 -74810
rect -22518 -74870 -22512 -74810
rect -22316 -74922 -22256 -74559
rect -22053 -74559 -22047 -74232
rect -22013 -74232 -21998 -74183
rect -21800 -74183 -21740 -73968
rect -22013 -74559 -22007 -74232
rect -22053 -74571 -22007 -74559
rect -21800 -74559 -21789 -74183
rect -21755 -74559 -21740 -74183
rect -22213 -74618 -22105 -74612
rect -22213 -74652 -22201 -74618
rect -22117 -74652 -22105 -74618
rect -22213 -74658 -22105 -74652
rect -21955 -74618 -21847 -74612
rect -21955 -74652 -21943 -74618
rect -21859 -74652 -21847 -74618
rect -21955 -74658 -21847 -74652
rect -21928 -74730 -21868 -74658
rect -21800 -74730 -21740 -74559
rect -21928 -74790 -21740 -74730
rect -22840 -74982 -22834 -74922
rect -22774 -74982 -22768 -74922
rect -22322 -74982 -22316 -74922
rect -22256 -74982 -22250 -74922
rect -21928 -75066 -21868 -74790
rect -21800 -75066 -21740 -74790
rect -21648 -74810 -21588 -73064
rect -21654 -74870 -21648 -74810
rect -21588 -74870 -21582 -74810
rect -23422 -75096 -21520 -75066
rect -23422 -75160 -23388 -75096
rect -21564 -75160 -21520 -75096
rect -23422 -75190 -21520 -75160
rect -23690 -75664 -23578 -75530
rect -22978 -75664 -22968 -75364
rect -22076 -75664 -22066 -75364
rect -21466 -75530 -21460 -72906
rect -21360 -75530 -21354 -72906
rect -20072 -72897 -19578 -72866
rect -20072 -72931 -20043 -72897
rect -20009 -72931 -19951 -72897
rect -19917 -72931 -19859 -72897
rect -19825 -72906 -19578 -72897
rect -19825 -72931 -19684 -72906
rect -20072 -72962 -19684 -72931
rect -21466 -75664 -21354 -75530
rect -23690 -75670 -21354 -75664
rect -23690 -75770 -23584 -75670
rect -21460 -75770 -21354 -75670
rect -23690 -75776 -21354 -75770
rect -19690 -75530 -19684 -72962
rect -19584 -75530 -19578 -72906
rect -18584 -72916 -18578 -72856
rect -18518 -72916 -18512 -72856
rect -19100 -73064 -19094 -73004
rect -19034 -73064 -19028 -73004
rect -19496 -73176 -19246 -73116
rect -19186 -73176 -19180 -73116
rect -19496 -74096 -19436 -73176
rect -19245 -73230 -19137 -73224
rect -19245 -73264 -19233 -73230
rect -19149 -73264 -19137 -73230
rect -19245 -73270 -19137 -73264
rect -19343 -73323 -19297 -73311
rect -19343 -73646 -19337 -73323
rect -19496 -74690 -19436 -74156
rect -19348 -73699 -19337 -73646
rect -19303 -73646 -19297 -73323
rect -19094 -73323 -19034 -73064
rect -18968 -73176 -18962 -73116
rect -18902 -73176 -18896 -73116
rect -18962 -73224 -18902 -73176
rect -18987 -73230 -18879 -73224
rect -18987 -73264 -18975 -73230
rect -18891 -73264 -18879 -73230
rect -18987 -73270 -18879 -73264
rect -18729 -73230 -18621 -73224
rect -18729 -73264 -18717 -73230
rect -18633 -73264 -18621 -73230
rect -18729 -73270 -18621 -73264
rect -19094 -73368 -19079 -73323
rect -19303 -73699 -19288 -73646
rect -19348 -73900 -19288 -73699
rect -19085 -73699 -19079 -73368
rect -19045 -73368 -19034 -73323
rect -18827 -73323 -18781 -73311
rect -18827 -73360 -18821 -73323
rect -19045 -73699 -19039 -73368
rect -19085 -73711 -19039 -73699
rect -18834 -73699 -18821 -73360
rect -18787 -73360 -18781 -73323
rect -18578 -73323 -18518 -72916
rect -18326 -72956 -18320 -72896
rect -18260 -72956 -18254 -72896
rect -18450 -73224 -18390 -73170
rect -18471 -73230 -18363 -73224
rect -18471 -73264 -18459 -73230
rect -18375 -73264 -18363 -73230
rect -18471 -73270 -18363 -73264
rect -18787 -73699 -18774 -73360
rect -18578 -73362 -18563 -73323
rect -18569 -73666 -18563 -73362
rect -19245 -73758 -19137 -73752
rect -19245 -73792 -19233 -73758
rect -19149 -73792 -19137 -73758
rect -19245 -73798 -19137 -73792
rect -18987 -73758 -18879 -73752
rect -18987 -73792 -18975 -73758
rect -18891 -73792 -18879 -73758
rect -18987 -73798 -18879 -73792
rect -19218 -73900 -19158 -73798
rect -19348 -73960 -19158 -73900
rect -19098 -73912 -19092 -73852
rect -19032 -73912 -19026 -73852
rect -19348 -74183 -19288 -73960
rect -19218 -74084 -19158 -73960
rect -19245 -74090 -19137 -74084
rect -19245 -74124 -19233 -74090
rect -19149 -74124 -19137 -74090
rect -19245 -74130 -19137 -74124
rect -19348 -74226 -19337 -74183
rect -19343 -74526 -19337 -74226
rect -19348 -74559 -19337 -74526
rect -19303 -74226 -19288 -74183
rect -19092 -74183 -19032 -73912
rect -18968 -74026 -18962 -73966
rect -18902 -74026 -18896 -73966
rect -18962 -74084 -18902 -74026
rect -18987 -74090 -18879 -74084
rect -18987 -74124 -18975 -74090
rect -18891 -74124 -18879 -74090
rect -18987 -74130 -18879 -74124
rect -19303 -74526 -19297 -74226
rect -19303 -74559 -19288 -74526
rect -19502 -74750 -19496 -74690
rect -19436 -74750 -19430 -74690
rect -19348 -74742 -19288 -74559
rect -19092 -74559 -19079 -74183
rect -19045 -74559 -19032 -74183
rect -19245 -74618 -19137 -74612
rect -19245 -74652 -19233 -74618
rect -19149 -74652 -19137 -74618
rect -19245 -74658 -19137 -74652
rect -19218 -74742 -19158 -74658
rect -19348 -74802 -19158 -74742
rect -19348 -75066 -19288 -74802
rect -19218 -75066 -19158 -74802
rect -19092 -74868 -19032 -74559
rect -18834 -74183 -18774 -73699
rect -18574 -73699 -18563 -73666
rect -18529 -73362 -18518 -73323
rect -18320 -73323 -18260 -72956
rect -18064 -73064 -18058 -73004
rect -17998 -73064 -17992 -73004
rect -18192 -73176 -18186 -73116
rect -18126 -73176 -18120 -73116
rect -18186 -73224 -18126 -73176
rect -18213 -73230 -18105 -73224
rect -18213 -73264 -18201 -73230
rect -18117 -73264 -18105 -73230
rect -18213 -73270 -18105 -73264
rect -18529 -73666 -18523 -73362
rect -18320 -73376 -18305 -73323
rect -18311 -73654 -18305 -73376
rect -18529 -73699 -18514 -73666
rect -18729 -73758 -18621 -73752
rect -18729 -73792 -18717 -73758
rect -18633 -73792 -18621 -73758
rect -18729 -73798 -18621 -73792
rect -18704 -73966 -18644 -73798
rect -18574 -73852 -18514 -73699
rect -18322 -73699 -18305 -73654
rect -18271 -73376 -18260 -73323
rect -18058 -73323 -17998 -73064
rect -17934 -73118 -17874 -72772
rect -17800 -73118 -17740 -72772
rect -17466 -72906 -17354 -72772
rect -15690 -72666 -13354 -72660
rect -15690 -72766 -15584 -72666
rect -13460 -72766 -13354 -72666
rect -15690 -72772 -13354 -72766
rect -15690 -72866 -15578 -72772
rect -17654 -73064 -17648 -73004
rect -17588 -73064 -17582 -73004
rect -17934 -73178 -17740 -73118
rect -17934 -73224 -17874 -73178
rect -17955 -73230 -17847 -73224
rect -17955 -73264 -17943 -73230
rect -17859 -73264 -17847 -73230
rect -17955 -73270 -17847 -73264
rect -18271 -73654 -18265 -73376
rect -18058 -73400 -18047 -73323
rect -18271 -73699 -18262 -73654
rect -18471 -73758 -18363 -73752
rect -18471 -73792 -18459 -73758
rect -18375 -73792 -18363 -73758
rect -18471 -73798 -18363 -73792
rect -18580 -73912 -18574 -73852
rect -18514 -73912 -18508 -73852
rect -18446 -73966 -18386 -73798
rect -18710 -74026 -18704 -73966
rect -18644 -74026 -18638 -73966
rect -18452 -74026 -18446 -73966
rect -18386 -74026 -18380 -73966
rect -18729 -74090 -18621 -74084
rect -18729 -74124 -18717 -74090
rect -18633 -74124 -18621 -74090
rect -18729 -74130 -18621 -74124
rect -18471 -74090 -18363 -74084
rect -18471 -74124 -18459 -74090
rect -18375 -74124 -18363 -74090
rect -18471 -74130 -18363 -74124
rect -18834 -74559 -18821 -74183
rect -18787 -74559 -18774 -74183
rect -18569 -74183 -18523 -74171
rect -18569 -74526 -18563 -74183
rect -18987 -74618 -18879 -74612
rect -18987 -74652 -18975 -74618
rect -18891 -74652 -18879 -74618
rect -18987 -74658 -18879 -74652
rect -19098 -74928 -19092 -74868
rect -19032 -74928 -19026 -74868
rect -18834 -74922 -18774 -74559
rect -18578 -74559 -18563 -74526
rect -18529 -74526 -18523 -74183
rect -18322 -74183 -18262 -73699
rect -18053 -73699 -18047 -73400
rect -18013 -73400 -17998 -73323
rect -17800 -73323 -17740 -73178
rect -18013 -73699 -18007 -73400
rect -18053 -73711 -18007 -73699
rect -17800 -73699 -17789 -73323
rect -17755 -73699 -17740 -73323
rect -18213 -73758 -18105 -73752
rect -18213 -73792 -18201 -73758
rect -18117 -73792 -18105 -73758
rect -18213 -73798 -18105 -73792
rect -17955 -73758 -17847 -73752
rect -17955 -73792 -17943 -73758
rect -17859 -73792 -17847 -73758
rect -17955 -73798 -17847 -73792
rect -18064 -73912 -18058 -73852
rect -17998 -73912 -17992 -73852
rect -17932 -73908 -17872 -73798
rect -17800 -73908 -17740 -73699
rect -18194 -74026 -18188 -73966
rect -18128 -74026 -18122 -73966
rect -18188 -74084 -18128 -74026
rect -18213 -74090 -18105 -74084
rect -18213 -74124 -18201 -74090
rect -18117 -74124 -18105 -74090
rect -18213 -74130 -18105 -74124
rect -18322 -74240 -18305 -74183
rect -18311 -74498 -18305 -74240
rect -18529 -74559 -18518 -74526
rect -18729 -74618 -18621 -74612
rect -18729 -74652 -18717 -74618
rect -18633 -74652 -18621 -74618
rect -18729 -74658 -18621 -74652
rect -18706 -74690 -18646 -74658
rect -18712 -74750 -18706 -74690
rect -18646 -74750 -18640 -74690
rect -18578 -74810 -18518 -74559
rect -18316 -74559 -18305 -74498
rect -18271 -74240 -18262 -74183
rect -18058 -74183 -17998 -73912
rect -17932 -73968 -17740 -73908
rect -17955 -74090 -17847 -74084
rect -17955 -74124 -17943 -74090
rect -17859 -74124 -17847 -74090
rect -17955 -74130 -17847 -74124
rect -18058 -74232 -18047 -74183
rect -18271 -74498 -18265 -74240
rect -18271 -74559 -18256 -74498
rect -18471 -74618 -18363 -74612
rect -18471 -74652 -18459 -74618
rect -18375 -74652 -18363 -74618
rect -18471 -74658 -18363 -74652
rect -18450 -74690 -18390 -74658
rect -18456 -74750 -18450 -74690
rect -18390 -74750 -18384 -74690
rect -18584 -74870 -18578 -74810
rect -18518 -74870 -18512 -74810
rect -18316 -74922 -18256 -74559
rect -18053 -74559 -18047 -74232
rect -18013 -74232 -17998 -74183
rect -17800 -74183 -17740 -73968
rect -18013 -74559 -18007 -74232
rect -18053 -74571 -18007 -74559
rect -17800 -74559 -17789 -74183
rect -17755 -74559 -17740 -74183
rect -18213 -74618 -18105 -74612
rect -18213 -74652 -18201 -74618
rect -18117 -74652 -18105 -74618
rect -18213 -74658 -18105 -74652
rect -17955 -74618 -17847 -74612
rect -17955 -74652 -17943 -74618
rect -17859 -74652 -17847 -74618
rect -17955 -74658 -17847 -74652
rect -17928 -74730 -17868 -74658
rect -17800 -74730 -17740 -74559
rect -17928 -74790 -17740 -74730
rect -18840 -74982 -18834 -74922
rect -18774 -74982 -18768 -74922
rect -18322 -74982 -18316 -74922
rect -18256 -74982 -18250 -74922
rect -17928 -75066 -17868 -74790
rect -17800 -75066 -17740 -74790
rect -17648 -74810 -17588 -73064
rect -17654 -74870 -17648 -74810
rect -17588 -74870 -17582 -74810
rect -19422 -75096 -17520 -75066
rect -19422 -75160 -19388 -75096
rect -17564 -75160 -17520 -75096
rect -19422 -75190 -17520 -75160
rect -19690 -75664 -19578 -75530
rect -18978 -75664 -18968 -75364
rect -18076 -75664 -18066 -75364
rect -17466 -75530 -17460 -72906
rect -17360 -75530 -17354 -72906
rect -16072 -72897 -15578 -72866
rect -16072 -72931 -16043 -72897
rect -16009 -72931 -15951 -72897
rect -15917 -72931 -15859 -72897
rect -15825 -72906 -15578 -72897
rect -15825 -72931 -15684 -72906
rect -16072 -72962 -15684 -72931
rect -17466 -75664 -17354 -75530
rect -19690 -75670 -17354 -75664
rect -19690 -75770 -19584 -75670
rect -17460 -75770 -17354 -75670
rect -19690 -75776 -17354 -75770
rect -15690 -75530 -15684 -72962
rect -15584 -75530 -15578 -72906
rect -14584 -72916 -14578 -72856
rect -14518 -72916 -14512 -72856
rect -15100 -73064 -15094 -73004
rect -15034 -73064 -15028 -73004
rect -15496 -73176 -15246 -73116
rect -15186 -73176 -15180 -73116
rect -15496 -74096 -15436 -73176
rect -15245 -73230 -15137 -73224
rect -15245 -73264 -15233 -73230
rect -15149 -73264 -15137 -73230
rect -15245 -73270 -15137 -73264
rect -15343 -73323 -15297 -73311
rect -15343 -73646 -15337 -73323
rect -15496 -74690 -15436 -74156
rect -15348 -73699 -15337 -73646
rect -15303 -73646 -15297 -73323
rect -15094 -73323 -15034 -73064
rect -14968 -73176 -14962 -73116
rect -14902 -73176 -14896 -73116
rect -14962 -73224 -14902 -73176
rect -14987 -73230 -14879 -73224
rect -14987 -73264 -14975 -73230
rect -14891 -73264 -14879 -73230
rect -14987 -73270 -14879 -73264
rect -14729 -73230 -14621 -73224
rect -14729 -73264 -14717 -73230
rect -14633 -73264 -14621 -73230
rect -14729 -73270 -14621 -73264
rect -15094 -73368 -15079 -73323
rect -15303 -73699 -15288 -73646
rect -15348 -73900 -15288 -73699
rect -15085 -73699 -15079 -73368
rect -15045 -73368 -15034 -73323
rect -14827 -73323 -14781 -73311
rect -14827 -73360 -14821 -73323
rect -15045 -73699 -15039 -73368
rect -15085 -73711 -15039 -73699
rect -14834 -73699 -14821 -73360
rect -14787 -73360 -14781 -73323
rect -14578 -73323 -14518 -72916
rect -14326 -72956 -14320 -72896
rect -14260 -72956 -14254 -72896
rect -14450 -73224 -14390 -73170
rect -14471 -73230 -14363 -73224
rect -14471 -73264 -14459 -73230
rect -14375 -73264 -14363 -73230
rect -14471 -73270 -14363 -73264
rect -14787 -73699 -14774 -73360
rect -14578 -73362 -14563 -73323
rect -14569 -73666 -14563 -73362
rect -15245 -73758 -15137 -73752
rect -15245 -73792 -15233 -73758
rect -15149 -73792 -15137 -73758
rect -15245 -73798 -15137 -73792
rect -14987 -73758 -14879 -73752
rect -14987 -73792 -14975 -73758
rect -14891 -73792 -14879 -73758
rect -14987 -73798 -14879 -73792
rect -15218 -73900 -15158 -73798
rect -15348 -73960 -15158 -73900
rect -15098 -73912 -15092 -73852
rect -15032 -73912 -15026 -73852
rect -15348 -74183 -15288 -73960
rect -15218 -74084 -15158 -73960
rect -15245 -74090 -15137 -74084
rect -15245 -74124 -15233 -74090
rect -15149 -74124 -15137 -74090
rect -15245 -74130 -15137 -74124
rect -15348 -74226 -15337 -74183
rect -15343 -74526 -15337 -74226
rect -15348 -74559 -15337 -74526
rect -15303 -74226 -15288 -74183
rect -15092 -74183 -15032 -73912
rect -14968 -74026 -14962 -73966
rect -14902 -74026 -14896 -73966
rect -14962 -74084 -14902 -74026
rect -14987 -74090 -14879 -74084
rect -14987 -74124 -14975 -74090
rect -14891 -74124 -14879 -74090
rect -14987 -74130 -14879 -74124
rect -15303 -74526 -15297 -74226
rect -15303 -74559 -15288 -74526
rect -15502 -74750 -15496 -74690
rect -15436 -74750 -15430 -74690
rect -15348 -74742 -15288 -74559
rect -15092 -74559 -15079 -74183
rect -15045 -74559 -15032 -74183
rect -15245 -74618 -15137 -74612
rect -15245 -74652 -15233 -74618
rect -15149 -74652 -15137 -74618
rect -15245 -74658 -15137 -74652
rect -15218 -74742 -15158 -74658
rect -15348 -74802 -15158 -74742
rect -15348 -75066 -15288 -74802
rect -15218 -75066 -15158 -74802
rect -15092 -74868 -15032 -74559
rect -14834 -74183 -14774 -73699
rect -14574 -73699 -14563 -73666
rect -14529 -73362 -14518 -73323
rect -14320 -73323 -14260 -72956
rect -14064 -73064 -14058 -73004
rect -13998 -73064 -13992 -73004
rect -14192 -73176 -14186 -73116
rect -14126 -73176 -14120 -73116
rect -14186 -73224 -14126 -73176
rect -14213 -73230 -14105 -73224
rect -14213 -73264 -14201 -73230
rect -14117 -73264 -14105 -73230
rect -14213 -73270 -14105 -73264
rect -14529 -73666 -14523 -73362
rect -14320 -73376 -14305 -73323
rect -14311 -73654 -14305 -73376
rect -14529 -73699 -14514 -73666
rect -14729 -73758 -14621 -73752
rect -14729 -73792 -14717 -73758
rect -14633 -73792 -14621 -73758
rect -14729 -73798 -14621 -73792
rect -14704 -73966 -14644 -73798
rect -14574 -73852 -14514 -73699
rect -14322 -73699 -14305 -73654
rect -14271 -73376 -14260 -73323
rect -14058 -73323 -13998 -73064
rect -13934 -73118 -13874 -72772
rect -13800 -73118 -13740 -72772
rect -13466 -72906 -13354 -72772
rect -11690 -72666 -9354 -72660
rect -11690 -72766 -11584 -72666
rect -9460 -72766 -9354 -72666
rect -11690 -72772 -9354 -72766
rect -11690 -72866 -11578 -72772
rect -13654 -73064 -13648 -73004
rect -13588 -73064 -13582 -73004
rect -13934 -73178 -13740 -73118
rect -13934 -73224 -13874 -73178
rect -13955 -73230 -13847 -73224
rect -13955 -73264 -13943 -73230
rect -13859 -73264 -13847 -73230
rect -13955 -73270 -13847 -73264
rect -14271 -73654 -14265 -73376
rect -14058 -73400 -14047 -73323
rect -14271 -73699 -14262 -73654
rect -14471 -73758 -14363 -73752
rect -14471 -73792 -14459 -73758
rect -14375 -73792 -14363 -73758
rect -14471 -73798 -14363 -73792
rect -14580 -73912 -14574 -73852
rect -14514 -73912 -14508 -73852
rect -14446 -73966 -14386 -73798
rect -14710 -74026 -14704 -73966
rect -14644 -74026 -14638 -73966
rect -14452 -74026 -14446 -73966
rect -14386 -74026 -14380 -73966
rect -14729 -74090 -14621 -74084
rect -14729 -74124 -14717 -74090
rect -14633 -74124 -14621 -74090
rect -14729 -74130 -14621 -74124
rect -14471 -74090 -14363 -74084
rect -14471 -74124 -14459 -74090
rect -14375 -74124 -14363 -74090
rect -14471 -74130 -14363 -74124
rect -14834 -74559 -14821 -74183
rect -14787 -74559 -14774 -74183
rect -14569 -74183 -14523 -74171
rect -14569 -74526 -14563 -74183
rect -14987 -74618 -14879 -74612
rect -14987 -74652 -14975 -74618
rect -14891 -74652 -14879 -74618
rect -14987 -74658 -14879 -74652
rect -15098 -74928 -15092 -74868
rect -15032 -74928 -15026 -74868
rect -14834 -74922 -14774 -74559
rect -14578 -74559 -14563 -74526
rect -14529 -74526 -14523 -74183
rect -14322 -74183 -14262 -73699
rect -14053 -73699 -14047 -73400
rect -14013 -73400 -13998 -73323
rect -13800 -73323 -13740 -73178
rect -14013 -73699 -14007 -73400
rect -14053 -73711 -14007 -73699
rect -13800 -73699 -13789 -73323
rect -13755 -73699 -13740 -73323
rect -14213 -73758 -14105 -73752
rect -14213 -73792 -14201 -73758
rect -14117 -73792 -14105 -73758
rect -14213 -73798 -14105 -73792
rect -13955 -73758 -13847 -73752
rect -13955 -73792 -13943 -73758
rect -13859 -73792 -13847 -73758
rect -13955 -73798 -13847 -73792
rect -14064 -73912 -14058 -73852
rect -13998 -73912 -13992 -73852
rect -13932 -73908 -13872 -73798
rect -13800 -73908 -13740 -73699
rect -14194 -74026 -14188 -73966
rect -14128 -74026 -14122 -73966
rect -14188 -74084 -14128 -74026
rect -14213 -74090 -14105 -74084
rect -14213 -74124 -14201 -74090
rect -14117 -74124 -14105 -74090
rect -14213 -74130 -14105 -74124
rect -14322 -74240 -14305 -74183
rect -14311 -74498 -14305 -74240
rect -14529 -74559 -14518 -74526
rect -14729 -74618 -14621 -74612
rect -14729 -74652 -14717 -74618
rect -14633 -74652 -14621 -74618
rect -14729 -74658 -14621 -74652
rect -14706 -74690 -14646 -74658
rect -14712 -74750 -14706 -74690
rect -14646 -74750 -14640 -74690
rect -14578 -74810 -14518 -74559
rect -14316 -74559 -14305 -74498
rect -14271 -74240 -14262 -74183
rect -14058 -74183 -13998 -73912
rect -13932 -73968 -13740 -73908
rect -13955 -74090 -13847 -74084
rect -13955 -74124 -13943 -74090
rect -13859 -74124 -13847 -74090
rect -13955 -74130 -13847 -74124
rect -14058 -74232 -14047 -74183
rect -14271 -74498 -14265 -74240
rect -14271 -74559 -14256 -74498
rect -14471 -74618 -14363 -74612
rect -14471 -74652 -14459 -74618
rect -14375 -74652 -14363 -74618
rect -14471 -74658 -14363 -74652
rect -14450 -74690 -14390 -74658
rect -14456 -74750 -14450 -74690
rect -14390 -74750 -14384 -74690
rect -14584 -74870 -14578 -74810
rect -14518 -74870 -14512 -74810
rect -14316 -74922 -14256 -74559
rect -14053 -74559 -14047 -74232
rect -14013 -74232 -13998 -74183
rect -13800 -74183 -13740 -73968
rect -14013 -74559 -14007 -74232
rect -14053 -74571 -14007 -74559
rect -13800 -74559 -13789 -74183
rect -13755 -74559 -13740 -74183
rect -14213 -74618 -14105 -74612
rect -14213 -74652 -14201 -74618
rect -14117 -74652 -14105 -74618
rect -14213 -74658 -14105 -74652
rect -13955 -74618 -13847 -74612
rect -13955 -74652 -13943 -74618
rect -13859 -74652 -13847 -74618
rect -13955 -74658 -13847 -74652
rect -13928 -74730 -13868 -74658
rect -13800 -74730 -13740 -74559
rect -13928 -74790 -13740 -74730
rect -14840 -74982 -14834 -74922
rect -14774 -74982 -14768 -74922
rect -14322 -74982 -14316 -74922
rect -14256 -74982 -14250 -74922
rect -13928 -75066 -13868 -74790
rect -13800 -75066 -13740 -74790
rect -13648 -74810 -13588 -73064
rect -13654 -74870 -13648 -74810
rect -13588 -74870 -13582 -74810
rect -15422 -75096 -13520 -75066
rect -15422 -75160 -15388 -75096
rect -13564 -75160 -13520 -75096
rect -15422 -75190 -13520 -75160
rect -15690 -75664 -15578 -75530
rect -14978 -75664 -14968 -75364
rect -14076 -75664 -14066 -75364
rect -13466 -75530 -13460 -72906
rect -13360 -75530 -13354 -72906
rect -12072 -72897 -11578 -72866
rect -12072 -72931 -12043 -72897
rect -12009 -72931 -11951 -72897
rect -11917 -72931 -11859 -72897
rect -11825 -72906 -11578 -72897
rect -11825 -72931 -11684 -72906
rect -12072 -72962 -11684 -72931
rect -13466 -75664 -13354 -75530
rect -15690 -75670 -13354 -75664
rect -15690 -75770 -15584 -75670
rect -13460 -75770 -13354 -75670
rect -15690 -75776 -13354 -75770
rect -11690 -75530 -11684 -72962
rect -11584 -75530 -11578 -72906
rect -10584 -72916 -10578 -72856
rect -10518 -72916 -10512 -72856
rect -11100 -73064 -11094 -73004
rect -11034 -73064 -11028 -73004
rect -11496 -73176 -11246 -73116
rect -11186 -73176 -11180 -73116
rect -11496 -74096 -11436 -73176
rect -11245 -73230 -11137 -73224
rect -11245 -73264 -11233 -73230
rect -11149 -73264 -11137 -73230
rect -11245 -73270 -11137 -73264
rect -11343 -73323 -11297 -73311
rect -11343 -73646 -11337 -73323
rect -11496 -74690 -11436 -74156
rect -11348 -73699 -11337 -73646
rect -11303 -73646 -11297 -73323
rect -11094 -73323 -11034 -73064
rect -10968 -73176 -10962 -73116
rect -10902 -73176 -10896 -73116
rect -10962 -73224 -10902 -73176
rect -10987 -73230 -10879 -73224
rect -10987 -73264 -10975 -73230
rect -10891 -73264 -10879 -73230
rect -10987 -73270 -10879 -73264
rect -10729 -73230 -10621 -73224
rect -10729 -73264 -10717 -73230
rect -10633 -73264 -10621 -73230
rect -10729 -73270 -10621 -73264
rect -11094 -73368 -11079 -73323
rect -11303 -73699 -11288 -73646
rect -11348 -73900 -11288 -73699
rect -11085 -73699 -11079 -73368
rect -11045 -73368 -11034 -73323
rect -10827 -73323 -10781 -73311
rect -10827 -73360 -10821 -73323
rect -11045 -73699 -11039 -73368
rect -11085 -73711 -11039 -73699
rect -10834 -73699 -10821 -73360
rect -10787 -73360 -10781 -73323
rect -10578 -73323 -10518 -72916
rect -10326 -72956 -10320 -72896
rect -10260 -72956 -10254 -72896
rect -10450 -73224 -10390 -73170
rect -10471 -73230 -10363 -73224
rect -10471 -73264 -10459 -73230
rect -10375 -73264 -10363 -73230
rect -10471 -73270 -10363 -73264
rect -10787 -73699 -10774 -73360
rect -10578 -73362 -10563 -73323
rect -10569 -73666 -10563 -73362
rect -11245 -73758 -11137 -73752
rect -11245 -73792 -11233 -73758
rect -11149 -73792 -11137 -73758
rect -11245 -73798 -11137 -73792
rect -10987 -73758 -10879 -73752
rect -10987 -73792 -10975 -73758
rect -10891 -73792 -10879 -73758
rect -10987 -73798 -10879 -73792
rect -11218 -73900 -11158 -73798
rect -11348 -73960 -11158 -73900
rect -11098 -73912 -11092 -73852
rect -11032 -73912 -11026 -73852
rect -11348 -74183 -11288 -73960
rect -11218 -74084 -11158 -73960
rect -11245 -74090 -11137 -74084
rect -11245 -74124 -11233 -74090
rect -11149 -74124 -11137 -74090
rect -11245 -74130 -11137 -74124
rect -11348 -74226 -11337 -74183
rect -11343 -74526 -11337 -74226
rect -11348 -74559 -11337 -74526
rect -11303 -74226 -11288 -74183
rect -11092 -74183 -11032 -73912
rect -10968 -74026 -10962 -73966
rect -10902 -74026 -10896 -73966
rect -10962 -74084 -10902 -74026
rect -10987 -74090 -10879 -74084
rect -10987 -74124 -10975 -74090
rect -10891 -74124 -10879 -74090
rect -10987 -74130 -10879 -74124
rect -11303 -74526 -11297 -74226
rect -11303 -74559 -11288 -74526
rect -11502 -74750 -11496 -74690
rect -11436 -74750 -11430 -74690
rect -11348 -74742 -11288 -74559
rect -11092 -74559 -11079 -74183
rect -11045 -74559 -11032 -74183
rect -11245 -74618 -11137 -74612
rect -11245 -74652 -11233 -74618
rect -11149 -74652 -11137 -74618
rect -11245 -74658 -11137 -74652
rect -11218 -74742 -11158 -74658
rect -11348 -74802 -11158 -74742
rect -11348 -75066 -11288 -74802
rect -11218 -75066 -11158 -74802
rect -11092 -74870 -11032 -74559
rect -10834 -74183 -10774 -73699
rect -10574 -73699 -10563 -73666
rect -10529 -73362 -10518 -73323
rect -10320 -73323 -10260 -72956
rect -10064 -73064 -10058 -73004
rect -9998 -73064 -9992 -73004
rect -10192 -73176 -10186 -73116
rect -10126 -73176 -10120 -73116
rect -10186 -73224 -10126 -73176
rect -10213 -73230 -10105 -73224
rect -10213 -73264 -10201 -73230
rect -10117 -73264 -10105 -73230
rect -10213 -73270 -10105 -73264
rect -10529 -73666 -10523 -73362
rect -10320 -73376 -10305 -73323
rect -10311 -73654 -10305 -73376
rect -10529 -73699 -10514 -73666
rect -10729 -73758 -10621 -73752
rect -10729 -73792 -10717 -73758
rect -10633 -73792 -10621 -73758
rect -10729 -73798 -10621 -73792
rect -10704 -73966 -10644 -73798
rect -10574 -73852 -10514 -73699
rect -10322 -73699 -10305 -73654
rect -10271 -73376 -10260 -73323
rect -10058 -73323 -9998 -73064
rect -9934 -73118 -9874 -72772
rect -9800 -73118 -9740 -72772
rect -9466 -72906 -9354 -72772
rect -7690 -72666 -5354 -72660
rect -7690 -72766 -7584 -72666
rect -5460 -72766 -5354 -72666
rect -7690 -72772 -5354 -72766
rect -7690 -72866 -7578 -72772
rect -9654 -73064 -9648 -73004
rect -9588 -73064 -9582 -73004
rect -9934 -73178 -9740 -73118
rect -9934 -73224 -9874 -73178
rect -9955 -73230 -9847 -73224
rect -9955 -73264 -9943 -73230
rect -9859 -73264 -9847 -73230
rect -9955 -73270 -9847 -73264
rect -10271 -73654 -10265 -73376
rect -10058 -73400 -10047 -73323
rect -10271 -73699 -10262 -73654
rect -10471 -73758 -10363 -73752
rect -10471 -73792 -10459 -73758
rect -10375 -73792 -10363 -73758
rect -10471 -73798 -10363 -73792
rect -10580 -73912 -10574 -73852
rect -10514 -73912 -10508 -73852
rect -10446 -73966 -10386 -73798
rect -10710 -74026 -10704 -73966
rect -10644 -74026 -10638 -73966
rect -10452 -74026 -10446 -73966
rect -10386 -74026 -10380 -73966
rect -10729 -74090 -10621 -74084
rect -10729 -74124 -10717 -74090
rect -10633 -74124 -10621 -74090
rect -10729 -74130 -10621 -74124
rect -10471 -74090 -10363 -74084
rect -10471 -74124 -10459 -74090
rect -10375 -74124 -10363 -74090
rect -10471 -74130 -10363 -74124
rect -10834 -74559 -10821 -74183
rect -10787 -74559 -10774 -74183
rect -10569 -74183 -10523 -74171
rect -10569 -74526 -10563 -74183
rect -10987 -74618 -10879 -74612
rect -10987 -74652 -10975 -74618
rect -10891 -74652 -10879 -74618
rect -10987 -74658 -10879 -74652
rect -11098 -74930 -11092 -74870
rect -11032 -74930 -11026 -74870
rect -10834 -74922 -10774 -74559
rect -10578 -74559 -10563 -74526
rect -10529 -74526 -10523 -74183
rect -10322 -74183 -10262 -73699
rect -10053 -73699 -10047 -73400
rect -10013 -73400 -9998 -73323
rect -9800 -73323 -9740 -73178
rect -10013 -73699 -10007 -73400
rect -10053 -73711 -10007 -73699
rect -9800 -73699 -9789 -73323
rect -9755 -73699 -9740 -73323
rect -10213 -73758 -10105 -73752
rect -10213 -73792 -10201 -73758
rect -10117 -73792 -10105 -73758
rect -10213 -73798 -10105 -73792
rect -9955 -73758 -9847 -73752
rect -9955 -73792 -9943 -73758
rect -9859 -73792 -9847 -73758
rect -9955 -73798 -9847 -73792
rect -10064 -73912 -10058 -73852
rect -9998 -73912 -9992 -73852
rect -9932 -73908 -9872 -73798
rect -9800 -73908 -9740 -73699
rect -10194 -74026 -10188 -73966
rect -10128 -74026 -10122 -73966
rect -10188 -74084 -10128 -74026
rect -10213 -74090 -10105 -74084
rect -10213 -74124 -10201 -74090
rect -10117 -74124 -10105 -74090
rect -10213 -74130 -10105 -74124
rect -10322 -74240 -10305 -74183
rect -10311 -74498 -10305 -74240
rect -10529 -74559 -10518 -74526
rect -10729 -74618 -10621 -74612
rect -10729 -74652 -10717 -74618
rect -10633 -74652 -10621 -74618
rect -10729 -74658 -10621 -74652
rect -10706 -74690 -10646 -74658
rect -10712 -74750 -10706 -74690
rect -10646 -74750 -10640 -74690
rect -10578 -74810 -10518 -74559
rect -10316 -74559 -10305 -74498
rect -10271 -74240 -10262 -74183
rect -10058 -74183 -9998 -73912
rect -9932 -73968 -9740 -73908
rect -9955 -74090 -9847 -74084
rect -9955 -74124 -9943 -74090
rect -9859 -74124 -9847 -74090
rect -9955 -74130 -9847 -74124
rect -10058 -74232 -10047 -74183
rect -10271 -74498 -10265 -74240
rect -10271 -74559 -10256 -74498
rect -10471 -74618 -10363 -74612
rect -10471 -74652 -10459 -74618
rect -10375 -74652 -10363 -74618
rect -10471 -74658 -10363 -74652
rect -10450 -74690 -10390 -74658
rect -10456 -74750 -10450 -74690
rect -10390 -74750 -10384 -74690
rect -10584 -74870 -10578 -74810
rect -10518 -74870 -10512 -74810
rect -10316 -74922 -10256 -74559
rect -10053 -74559 -10047 -74232
rect -10013 -74232 -9998 -74183
rect -9800 -74183 -9740 -73968
rect -10013 -74559 -10007 -74232
rect -10053 -74571 -10007 -74559
rect -9800 -74559 -9789 -74183
rect -9755 -74559 -9740 -74183
rect -10213 -74618 -10105 -74612
rect -10213 -74652 -10201 -74618
rect -10117 -74652 -10105 -74618
rect -10213 -74658 -10105 -74652
rect -9955 -74618 -9847 -74612
rect -9955 -74652 -9943 -74618
rect -9859 -74652 -9847 -74618
rect -9955 -74658 -9847 -74652
rect -9928 -74730 -9868 -74658
rect -9800 -74730 -9740 -74559
rect -9928 -74790 -9740 -74730
rect -10840 -74982 -10834 -74922
rect -10774 -74982 -10768 -74922
rect -10322 -74982 -10316 -74922
rect -10256 -74982 -10250 -74922
rect -9928 -75066 -9868 -74790
rect -9800 -75066 -9740 -74790
rect -9648 -74810 -9588 -73064
rect -9654 -74870 -9648 -74810
rect -9588 -74870 -9582 -74810
rect -11422 -75096 -9520 -75066
rect -11422 -75160 -11388 -75096
rect -9564 -75160 -9520 -75096
rect -11422 -75190 -9520 -75160
rect -11690 -75664 -11578 -75530
rect -10978 -75664 -10968 -75364
rect -10076 -75664 -10066 -75364
rect -9466 -75530 -9460 -72906
rect -9360 -75530 -9354 -72906
rect -8072 -72897 -7578 -72866
rect -8072 -72931 -8043 -72897
rect -8009 -72931 -7951 -72897
rect -7917 -72931 -7859 -72897
rect -7825 -72906 -7578 -72897
rect -7825 -72931 -7684 -72906
rect -8072 -72962 -7684 -72931
rect -9466 -75664 -9354 -75530
rect -11690 -75670 -9354 -75664
rect -11690 -75770 -11584 -75670
rect -9460 -75770 -9354 -75670
rect -11690 -75776 -9354 -75770
rect -7690 -75530 -7684 -72962
rect -7584 -75530 -7578 -72906
rect -6584 -72916 -6578 -72856
rect -6518 -72916 -6512 -72856
rect -7100 -73064 -7094 -73004
rect -7034 -73064 -7028 -73004
rect -7496 -73176 -7246 -73116
rect -7186 -73176 -7180 -73116
rect -7496 -74096 -7436 -73176
rect -7245 -73230 -7137 -73224
rect -7245 -73264 -7233 -73230
rect -7149 -73264 -7137 -73230
rect -7245 -73270 -7137 -73264
rect -7343 -73323 -7297 -73311
rect -7343 -73646 -7337 -73323
rect -7496 -74690 -7436 -74156
rect -7348 -73699 -7337 -73646
rect -7303 -73646 -7297 -73323
rect -7094 -73323 -7034 -73064
rect -6968 -73176 -6962 -73116
rect -6902 -73176 -6896 -73116
rect -6962 -73224 -6902 -73176
rect -6987 -73230 -6879 -73224
rect -6987 -73264 -6975 -73230
rect -6891 -73264 -6879 -73230
rect -6987 -73270 -6879 -73264
rect -6729 -73230 -6621 -73224
rect -6729 -73264 -6717 -73230
rect -6633 -73264 -6621 -73230
rect -6729 -73270 -6621 -73264
rect -7094 -73368 -7079 -73323
rect -7303 -73699 -7288 -73646
rect -7348 -73900 -7288 -73699
rect -7085 -73699 -7079 -73368
rect -7045 -73368 -7034 -73323
rect -6827 -73323 -6781 -73311
rect -6827 -73360 -6821 -73323
rect -7045 -73699 -7039 -73368
rect -7085 -73711 -7039 -73699
rect -6834 -73699 -6821 -73360
rect -6787 -73360 -6781 -73323
rect -6578 -73323 -6518 -72916
rect -6326 -72956 -6320 -72896
rect -6260 -72956 -6254 -72896
rect -6450 -73224 -6390 -73170
rect -6471 -73230 -6363 -73224
rect -6471 -73264 -6459 -73230
rect -6375 -73264 -6363 -73230
rect -6471 -73270 -6363 -73264
rect -6787 -73699 -6774 -73360
rect -6578 -73362 -6563 -73323
rect -6569 -73666 -6563 -73362
rect -7245 -73758 -7137 -73752
rect -7245 -73792 -7233 -73758
rect -7149 -73792 -7137 -73758
rect -7245 -73798 -7137 -73792
rect -6987 -73758 -6879 -73752
rect -6987 -73792 -6975 -73758
rect -6891 -73792 -6879 -73758
rect -6987 -73798 -6879 -73792
rect -7218 -73900 -7158 -73798
rect -7348 -73960 -7158 -73900
rect -7098 -73912 -7092 -73852
rect -7032 -73912 -7026 -73852
rect -7348 -74183 -7288 -73960
rect -7218 -74084 -7158 -73960
rect -7245 -74090 -7137 -74084
rect -7245 -74124 -7233 -74090
rect -7149 -74124 -7137 -74090
rect -7245 -74130 -7137 -74124
rect -7348 -74226 -7337 -74183
rect -7343 -74526 -7337 -74226
rect -7348 -74559 -7337 -74526
rect -7303 -74226 -7288 -74183
rect -7092 -74183 -7032 -73912
rect -6968 -74026 -6962 -73966
rect -6902 -74026 -6896 -73966
rect -6962 -74084 -6902 -74026
rect -6987 -74090 -6879 -74084
rect -6987 -74124 -6975 -74090
rect -6891 -74124 -6879 -74090
rect -6987 -74130 -6879 -74124
rect -7303 -74526 -7297 -74226
rect -7303 -74559 -7288 -74526
rect -7502 -74750 -7496 -74690
rect -7436 -74750 -7430 -74690
rect -7348 -74742 -7288 -74559
rect -7092 -74559 -7079 -74183
rect -7045 -74559 -7032 -74183
rect -7245 -74618 -7137 -74612
rect -7245 -74652 -7233 -74618
rect -7149 -74652 -7137 -74618
rect -7245 -74658 -7137 -74652
rect -7218 -74742 -7158 -74658
rect -7348 -74802 -7158 -74742
rect -7348 -75066 -7288 -74802
rect -7218 -75066 -7158 -74802
rect -7092 -74870 -7032 -74559
rect -6834 -74183 -6774 -73699
rect -6574 -73699 -6563 -73666
rect -6529 -73362 -6518 -73323
rect -6320 -73323 -6260 -72956
rect -6064 -73064 -6058 -73004
rect -5998 -73064 -5992 -73004
rect -6192 -73176 -6186 -73116
rect -6126 -73176 -6120 -73116
rect -6186 -73224 -6126 -73176
rect -6213 -73230 -6105 -73224
rect -6213 -73264 -6201 -73230
rect -6117 -73264 -6105 -73230
rect -6213 -73270 -6105 -73264
rect -6529 -73666 -6523 -73362
rect -6320 -73376 -6305 -73323
rect -6311 -73654 -6305 -73376
rect -6529 -73699 -6514 -73666
rect -6729 -73758 -6621 -73752
rect -6729 -73792 -6717 -73758
rect -6633 -73792 -6621 -73758
rect -6729 -73798 -6621 -73792
rect -6704 -73966 -6644 -73798
rect -6574 -73852 -6514 -73699
rect -6322 -73699 -6305 -73654
rect -6271 -73376 -6260 -73323
rect -6058 -73323 -5998 -73064
rect -5934 -73118 -5874 -72772
rect -5800 -73118 -5740 -72772
rect -5466 -72906 -5354 -72772
rect -3690 -72666 -1354 -72660
rect -3690 -72766 -3584 -72666
rect -1460 -72766 -1354 -72666
rect -3690 -72772 -1354 -72766
rect -3690 -72866 -3578 -72772
rect -5654 -73064 -5648 -73004
rect -5588 -73064 -5582 -73004
rect -5934 -73178 -5740 -73118
rect -5934 -73224 -5874 -73178
rect -5955 -73230 -5847 -73224
rect -5955 -73264 -5943 -73230
rect -5859 -73264 -5847 -73230
rect -5955 -73270 -5847 -73264
rect -6271 -73654 -6265 -73376
rect -6058 -73400 -6047 -73323
rect -6271 -73699 -6262 -73654
rect -6471 -73758 -6363 -73752
rect -6471 -73792 -6459 -73758
rect -6375 -73792 -6363 -73758
rect -6471 -73798 -6363 -73792
rect -6580 -73912 -6574 -73852
rect -6514 -73912 -6508 -73852
rect -6446 -73966 -6386 -73798
rect -6710 -74026 -6704 -73966
rect -6644 -74026 -6638 -73966
rect -6452 -74026 -6446 -73966
rect -6386 -74026 -6380 -73966
rect -6729 -74090 -6621 -74084
rect -6729 -74124 -6717 -74090
rect -6633 -74124 -6621 -74090
rect -6729 -74130 -6621 -74124
rect -6471 -74090 -6363 -74084
rect -6471 -74124 -6459 -74090
rect -6375 -74124 -6363 -74090
rect -6471 -74130 -6363 -74124
rect -6834 -74559 -6821 -74183
rect -6787 -74559 -6774 -74183
rect -6569 -74183 -6523 -74171
rect -6569 -74526 -6563 -74183
rect -6987 -74618 -6879 -74612
rect -6987 -74652 -6975 -74618
rect -6891 -74652 -6879 -74618
rect -6987 -74658 -6879 -74652
rect -7098 -74930 -7092 -74870
rect -7032 -74930 -7026 -74870
rect -6834 -74922 -6774 -74559
rect -6578 -74559 -6563 -74526
rect -6529 -74526 -6523 -74183
rect -6322 -74183 -6262 -73699
rect -6053 -73699 -6047 -73400
rect -6013 -73400 -5998 -73323
rect -5800 -73323 -5740 -73178
rect -6013 -73699 -6007 -73400
rect -6053 -73711 -6007 -73699
rect -5800 -73699 -5789 -73323
rect -5755 -73699 -5740 -73323
rect -6213 -73758 -6105 -73752
rect -6213 -73792 -6201 -73758
rect -6117 -73792 -6105 -73758
rect -6213 -73798 -6105 -73792
rect -5955 -73758 -5847 -73752
rect -5955 -73792 -5943 -73758
rect -5859 -73792 -5847 -73758
rect -5955 -73798 -5847 -73792
rect -6064 -73912 -6058 -73852
rect -5998 -73912 -5992 -73852
rect -5932 -73908 -5872 -73798
rect -5800 -73908 -5740 -73699
rect -6194 -74026 -6188 -73966
rect -6128 -74026 -6122 -73966
rect -6188 -74084 -6128 -74026
rect -6213 -74090 -6105 -74084
rect -6213 -74124 -6201 -74090
rect -6117 -74124 -6105 -74090
rect -6213 -74130 -6105 -74124
rect -6322 -74240 -6305 -74183
rect -6311 -74498 -6305 -74240
rect -6529 -74559 -6518 -74526
rect -6729 -74618 -6621 -74612
rect -6729 -74652 -6717 -74618
rect -6633 -74652 -6621 -74618
rect -6729 -74658 -6621 -74652
rect -6706 -74690 -6646 -74658
rect -6712 -74750 -6706 -74690
rect -6646 -74750 -6640 -74690
rect -6578 -74810 -6518 -74559
rect -6316 -74559 -6305 -74498
rect -6271 -74240 -6262 -74183
rect -6058 -74183 -5998 -73912
rect -5932 -73968 -5740 -73908
rect -5955 -74090 -5847 -74084
rect -5955 -74124 -5943 -74090
rect -5859 -74124 -5847 -74090
rect -5955 -74130 -5847 -74124
rect -6058 -74232 -6047 -74183
rect -6271 -74498 -6265 -74240
rect -6271 -74559 -6256 -74498
rect -6471 -74618 -6363 -74612
rect -6471 -74652 -6459 -74618
rect -6375 -74652 -6363 -74618
rect -6471 -74658 -6363 -74652
rect -6450 -74690 -6390 -74658
rect -6456 -74750 -6450 -74690
rect -6390 -74750 -6384 -74690
rect -6584 -74870 -6578 -74810
rect -6518 -74870 -6512 -74810
rect -6316 -74922 -6256 -74559
rect -6053 -74559 -6047 -74232
rect -6013 -74232 -5998 -74183
rect -5800 -74183 -5740 -73968
rect -6013 -74559 -6007 -74232
rect -6053 -74571 -6007 -74559
rect -5800 -74559 -5789 -74183
rect -5755 -74559 -5740 -74183
rect -6213 -74618 -6105 -74612
rect -6213 -74652 -6201 -74618
rect -6117 -74652 -6105 -74618
rect -6213 -74658 -6105 -74652
rect -5955 -74618 -5847 -74612
rect -5955 -74652 -5943 -74618
rect -5859 -74652 -5847 -74618
rect -5955 -74658 -5847 -74652
rect -5928 -74730 -5868 -74658
rect -5800 -74730 -5740 -74559
rect -5928 -74790 -5740 -74730
rect -6840 -74982 -6834 -74922
rect -6774 -74982 -6768 -74922
rect -6322 -74982 -6316 -74922
rect -6256 -74982 -6250 -74922
rect -5928 -75066 -5868 -74790
rect -5800 -75066 -5740 -74790
rect -5648 -74810 -5588 -73064
rect -5654 -74870 -5648 -74810
rect -5588 -74870 -5582 -74810
rect -7422 -75096 -5520 -75066
rect -7422 -75160 -7388 -75096
rect -5564 -75160 -5520 -75096
rect -7422 -75190 -5520 -75160
rect -7690 -75664 -7578 -75530
rect -6978 -75664 -6968 -75364
rect -6076 -75664 -6066 -75364
rect -5466 -75530 -5460 -72906
rect -5360 -75530 -5354 -72906
rect -4072 -72897 -3578 -72866
rect -4072 -72931 -4043 -72897
rect -4009 -72931 -3951 -72897
rect -3917 -72931 -3859 -72897
rect -3825 -72906 -3578 -72897
rect -3825 -72931 -3684 -72906
rect -4072 -72962 -3684 -72931
rect -5466 -75664 -5354 -75530
rect -7690 -75670 -5354 -75664
rect -7690 -75770 -7584 -75670
rect -5460 -75770 -5354 -75670
rect -7690 -75776 -5354 -75770
rect -3690 -75530 -3684 -72962
rect -3584 -75530 -3578 -72906
rect -2584 -72916 -2578 -72856
rect -2518 -72916 -2512 -72856
rect -3100 -73064 -3094 -73004
rect -3034 -73064 -3028 -73004
rect -3496 -73176 -3246 -73116
rect -3186 -73176 -3180 -73116
rect -3496 -74096 -3436 -73176
rect -3245 -73230 -3137 -73224
rect -3245 -73264 -3233 -73230
rect -3149 -73264 -3137 -73230
rect -3245 -73270 -3137 -73264
rect -3343 -73323 -3297 -73311
rect -3343 -73646 -3337 -73323
rect -3496 -74690 -3436 -74156
rect -3348 -73699 -3337 -73646
rect -3303 -73646 -3297 -73323
rect -3094 -73323 -3034 -73064
rect -2968 -73176 -2962 -73116
rect -2902 -73176 -2896 -73116
rect -2962 -73224 -2902 -73176
rect -2987 -73230 -2879 -73224
rect -2987 -73264 -2975 -73230
rect -2891 -73264 -2879 -73230
rect -2987 -73270 -2879 -73264
rect -2729 -73230 -2621 -73224
rect -2729 -73264 -2717 -73230
rect -2633 -73264 -2621 -73230
rect -2729 -73270 -2621 -73264
rect -3094 -73368 -3079 -73323
rect -3303 -73699 -3288 -73646
rect -3348 -73900 -3288 -73699
rect -3085 -73699 -3079 -73368
rect -3045 -73368 -3034 -73323
rect -2827 -73323 -2781 -73311
rect -2827 -73360 -2821 -73323
rect -3045 -73699 -3039 -73368
rect -3085 -73711 -3039 -73699
rect -2834 -73699 -2821 -73360
rect -2787 -73360 -2781 -73323
rect -2578 -73323 -2518 -72916
rect -2326 -72956 -2320 -72896
rect -2260 -72956 -2254 -72896
rect -2450 -73224 -2390 -73170
rect -2471 -73230 -2363 -73224
rect -2471 -73264 -2459 -73230
rect -2375 -73264 -2363 -73230
rect -2471 -73270 -2363 -73264
rect -2787 -73699 -2774 -73360
rect -2578 -73362 -2563 -73323
rect -2569 -73666 -2563 -73362
rect -3245 -73758 -3137 -73752
rect -3245 -73792 -3233 -73758
rect -3149 -73792 -3137 -73758
rect -3245 -73798 -3137 -73792
rect -2987 -73758 -2879 -73752
rect -2987 -73792 -2975 -73758
rect -2891 -73792 -2879 -73758
rect -2987 -73798 -2879 -73792
rect -3218 -73900 -3158 -73798
rect -3348 -73960 -3158 -73900
rect -3098 -73912 -3092 -73852
rect -3032 -73912 -3026 -73852
rect -3348 -74183 -3288 -73960
rect -3218 -74084 -3158 -73960
rect -3245 -74090 -3137 -74084
rect -3245 -74124 -3233 -74090
rect -3149 -74124 -3137 -74090
rect -3245 -74130 -3137 -74124
rect -3348 -74226 -3337 -74183
rect -3343 -74526 -3337 -74226
rect -3348 -74559 -3337 -74526
rect -3303 -74226 -3288 -74183
rect -3092 -74183 -3032 -73912
rect -2968 -74026 -2962 -73966
rect -2902 -74026 -2896 -73966
rect -2962 -74084 -2902 -74026
rect -2987 -74090 -2879 -74084
rect -2987 -74124 -2975 -74090
rect -2891 -74124 -2879 -74090
rect -2987 -74130 -2879 -74124
rect -3303 -74526 -3297 -74226
rect -3303 -74559 -3288 -74526
rect -3502 -74750 -3496 -74690
rect -3436 -74750 -3430 -74690
rect -3348 -74742 -3288 -74559
rect -3092 -74559 -3079 -74183
rect -3045 -74559 -3032 -74183
rect -3245 -74618 -3137 -74612
rect -3245 -74652 -3233 -74618
rect -3149 -74652 -3137 -74618
rect -3245 -74658 -3137 -74652
rect -3218 -74742 -3158 -74658
rect -3348 -74802 -3158 -74742
rect -3348 -75066 -3288 -74802
rect -3218 -75066 -3158 -74802
rect -3092 -74868 -3032 -74559
rect -2834 -74183 -2774 -73699
rect -2574 -73699 -2563 -73666
rect -2529 -73362 -2518 -73323
rect -2320 -73323 -2260 -72956
rect -2064 -73064 -2058 -73004
rect -1998 -73064 -1992 -73004
rect -2192 -73176 -2186 -73116
rect -2126 -73176 -2120 -73116
rect -2186 -73224 -2126 -73176
rect -2213 -73230 -2105 -73224
rect -2213 -73264 -2201 -73230
rect -2117 -73264 -2105 -73230
rect -2213 -73270 -2105 -73264
rect -2529 -73666 -2523 -73362
rect -2320 -73376 -2305 -73323
rect -2311 -73654 -2305 -73376
rect -2529 -73699 -2514 -73666
rect -2729 -73758 -2621 -73752
rect -2729 -73792 -2717 -73758
rect -2633 -73792 -2621 -73758
rect -2729 -73798 -2621 -73792
rect -2704 -73966 -2644 -73798
rect -2574 -73852 -2514 -73699
rect -2322 -73699 -2305 -73654
rect -2271 -73376 -2260 -73323
rect -2058 -73323 -1998 -73064
rect -1934 -73118 -1874 -72772
rect -1800 -73118 -1740 -72772
rect -1466 -72906 -1354 -72772
rect 310 -72666 2646 -72660
rect 310 -72766 416 -72666
rect 2540 -72766 2646 -72666
rect 310 -72772 2646 -72766
rect 310 -72866 422 -72772
rect -1654 -73064 -1648 -73004
rect -1588 -73064 -1582 -73004
rect -1934 -73178 -1740 -73118
rect -1934 -73224 -1874 -73178
rect -1955 -73230 -1847 -73224
rect -1955 -73264 -1943 -73230
rect -1859 -73264 -1847 -73230
rect -1955 -73270 -1847 -73264
rect -2271 -73654 -2265 -73376
rect -2058 -73400 -2047 -73323
rect -2271 -73699 -2262 -73654
rect -2471 -73758 -2363 -73752
rect -2471 -73792 -2459 -73758
rect -2375 -73792 -2363 -73758
rect -2471 -73798 -2363 -73792
rect -2580 -73912 -2574 -73852
rect -2514 -73912 -2508 -73852
rect -2446 -73966 -2386 -73798
rect -2710 -74026 -2704 -73966
rect -2644 -74026 -2638 -73966
rect -2452 -74026 -2446 -73966
rect -2386 -74026 -2380 -73966
rect -2729 -74090 -2621 -74084
rect -2729 -74124 -2717 -74090
rect -2633 -74124 -2621 -74090
rect -2729 -74130 -2621 -74124
rect -2471 -74090 -2363 -74084
rect -2471 -74124 -2459 -74090
rect -2375 -74124 -2363 -74090
rect -2471 -74130 -2363 -74124
rect -2834 -74559 -2821 -74183
rect -2787 -74559 -2774 -74183
rect -2569 -74183 -2523 -74171
rect -2569 -74526 -2563 -74183
rect -2987 -74618 -2879 -74612
rect -2987 -74652 -2975 -74618
rect -2891 -74652 -2879 -74618
rect -2987 -74658 -2879 -74652
rect -3098 -74928 -3092 -74868
rect -3032 -74928 -3026 -74868
rect -2834 -74922 -2774 -74559
rect -2578 -74559 -2563 -74526
rect -2529 -74526 -2523 -74183
rect -2322 -74183 -2262 -73699
rect -2053 -73699 -2047 -73400
rect -2013 -73400 -1998 -73323
rect -1800 -73323 -1740 -73178
rect -2013 -73699 -2007 -73400
rect -2053 -73711 -2007 -73699
rect -1800 -73699 -1789 -73323
rect -1755 -73699 -1740 -73323
rect -2213 -73758 -2105 -73752
rect -2213 -73792 -2201 -73758
rect -2117 -73792 -2105 -73758
rect -2213 -73798 -2105 -73792
rect -1955 -73758 -1847 -73752
rect -1955 -73792 -1943 -73758
rect -1859 -73792 -1847 -73758
rect -1955 -73798 -1847 -73792
rect -2064 -73912 -2058 -73852
rect -1998 -73912 -1992 -73852
rect -1932 -73908 -1872 -73798
rect -1800 -73908 -1740 -73699
rect -2194 -74026 -2188 -73966
rect -2128 -74026 -2122 -73966
rect -2188 -74084 -2128 -74026
rect -2213 -74090 -2105 -74084
rect -2213 -74124 -2201 -74090
rect -2117 -74124 -2105 -74090
rect -2213 -74130 -2105 -74124
rect -2322 -74240 -2305 -74183
rect -2311 -74498 -2305 -74240
rect -2529 -74559 -2518 -74526
rect -2729 -74618 -2621 -74612
rect -2729 -74652 -2717 -74618
rect -2633 -74652 -2621 -74618
rect -2729 -74658 -2621 -74652
rect -2706 -74690 -2646 -74658
rect -2712 -74750 -2706 -74690
rect -2646 -74750 -2640 -74690
rect -2578 -74810 -2518 -74559
rect -2316 -74559 -2305 -74498
rect -2271 -74240 -2262 -74183
rect -2058 -74183 -1998 -73912
rect -1932 -73968 -1740 -73908
rect -1955 -74090 -1847 -74084
rect -1955 -74124 -1943 -74090
rect -1859 -74124 -1847 -74090
rect -1955 -74130 -1847 -74124
rect -2058 -74232 -2047 -74183
rect -2271 -74498 -2265 -74240
rect -2271 -74559 -2256 -74498
rect -2471 -74618 -2363 -74612
rect -2471 -74652 -2459 -74618
rect -2375 -74652 -2363 -74618
rect -2471 -74658 -2363 -74652
rect -2450 -74690 -2390 -74658
rect -2456 -74750 -2450 -74690
rect -2390 -74750 -2384 -74690
rect -2584 -74870 -2578 -74810
rect -2518 -74870 -2512 -74810
rect -2316 -74922 -2256 -74559
rect -2053 -74559 -2047 -74232
rect -2013 -74232 -1998 -74183
rect -1800 -74183 -1740 -73968
rect -2013 -74559 -2007 -74232
rect -2053 -74571 -2007 -74559
rect -1800 -74559 -1789 -74183
rect -1755 -74559 -1740 -74183
rect -2213 -74618 -2105 -74612
rect -2213 -74652 -2201 -74618
rect -2117 -74652 -2105 -74618
rect -2213 -74658 -2105 -74652
rect -1955 -74618 -1847 -74612
rect -1955 -74652 -1943 -74618
rect -1859 -74652 -1847 -74618
rect -1955 -74658 -1847 -74652
rect -1928 -74730 -1868 -74658
rect -1800 -74730 -1740 -74559
rect -1928 -74790 -1740 -74730
rect -2840 -74982 -2834 -74922
rect -2774 -74982 -2768 -74922
rect -2322 -74982 -2316 -74922
rect -2256 -74982 -2250 -74922
rect -1928 -75066 -1868 -74790
rect -1800 -75066 -1740 -74790
rect -1648 -74810 -1588 -73064
rect -1654 -74870 -1648 -74810
rect -1588 -74870 -1582 -74810
rect -3422 -75096 -1520 -75066
rect -3422 -75160 -3388 -75096
rect -1564 -75160 -1520 -75096
rect -3422 -75190 -1520 -75160
rect -3690 -75664 -3578 -75530
rect -2978 -75664 -2968 -75364
rect -2076 -75664 -2066 -75364
rect -1466 -75530 -1460 -72906
rect -1360 -75530 -1354 -72906
rect -72 -72897 422 -72866
rect -72 -72931 -43 -72897
rect -9 -72931 49 -72897
rect 83 -72931 141 -72897
rect 175 -72906 422 -72897
rect 175 -72931 316 -72906
rect -72 -72962 316 -72931
rect -1466 -75664 -1354 -75530
rect -3690 -75670 -1354 -75664
rect -3690 -75770 -3584 -75670
rect -1460 -75770 -1354 -75670
rect -3690 -75776 -1354 -75770
rect 310 -75530 316 -72962
rect 416 -75530 422 -72906
rect 1416 -72916 1422 -72856
rect 1482 -72916 1488 -72856
rect 900 -73064 906 -73004
rect 966 -73064 972 -73004
rect 504 -73176 754 -73116
rect 814 -73176 820 -73116
rect 504 -74096 564 -73176
rect 755 -73230 863 -73224
rect 755 -73264 767 -73230
rect 851 -73264 863 -73230
rect 755 -73270 863 -73264
rect 657 -73323 703 -73311
rect 657 -73646 663 -73323
rect 504 -74690 564 -74156
rect 652 -73699 663 -73646
rect 697 -73646 703 -73323
rect 906 -73323 966 -73064
rect 1032 -73176 1038 -73116
rect 1098 -73176 1104 -73116
rect 1038 -73224 1098 -73176
rect 1013 -73230 1121 -73224
rect 1013 -73264 1025 -73230
rect 1109 -73264 1121 -73230
rect 1013 -73270 1121 -73264
rect 1271 -73230 1379 -73224
rect 1271 -73264 1283 -73230
rect 1367 -73264 1379 -73230
rect 1271 -73270 1379 -73264
rect 906 -73368 921 -73323
rect 697 -73699 712 -73646
rect 652 -73900 712 -73699
rect 915 -73699 921 -73368
rect 955 -73368 966 -73323
rect 1173 -73323 1219 -73311
rect 1173 -73360 1179 -73323
rect 955 -73699 961 -73368
rect 915 -73711 961 -73699
rect 1166 -73699 1179 -73360
rect 1213 -73360 1219 -73323
rect 1422 -73323 1482 -72916
rect 1674 -72956 1680 -72896
rect 1740 -72956 1746 -72896
rect 1550 -73224 1610 -73170
rect 1529 -73230 1637 -73224
rect 1529 -73264 1541 -73230
rect 1625 -73264 1637 -73230
rect 1529 -73270 1637 -73264
rect 1213 -73699 1226 -73360
rect 1422 -73362 1437 -73323
rect 1431 -73666 1437 -73362
rect 755 -73758 863 -73752
rect 755 -73792 767 -73758
rect 851 -73792 863 -73758
rect 755 -73798 863 -73792
rect 1013 -73758 1121 -73752
rect 1013 -73792 1025 -73758
rect 1109 -73792 1121 -73758
rect 1013 -73798 1121 -73792
rect 782 -73900 842 -73798
rect 652 -73960 842 -73900
rect 902 -73912 908 -73852
rect 968 -73912 974 -73852
rect 652 -74183 712 -73960
rect 782 -74084 842 -73960
rect 755 -74090 863 -74084
rect 755 -74124 767 -74090
rect 851 -74124 863 -74090
rect 755 -74130 863 -74124
rect 652 -74226 663 -74183
rect 657 -74526 663 -74226
rect 652 -74559 663 -74526
rect 697 -74226 712 -74183
rect 908 -74183 968 -73912
rect 1032 -74026 1038 -73966
rect 1098 -74026 1104 -73966
rect 1038 -74084 1098 -74026
rect 1013 -74090 1121 -74084
rect 1013 -74124 1025 -74090
rect 1109 -74124 1121 -74090
rect 1013 -74130 1121 -74124
rect 697 -74526 703 -74226
rect 697 -74559 712 -74526
rect 498 -74750 504 -74690
rect 564 -74750 570 -74690
rect 652 -74742 712 -74559
rect 908 -74559 921 -74183
rect 955 -74559 968 -74183
rect 755 -74618 863 -74612
rect 755 -74652 767 -74618
rect 851 -74652 863 -74618
rect 755 -74658 863 -74652
rect 782 -74742 842 -74658
rect 652 -74802 842 -74742
rect 652 -75066 712 -74802
rect 782 -75066 842 -74802
rect 908 -74868 968 -74559
rect 1166 -74183 1226 -73699
rect 1426 -73699 1437 -73666
rect 1471 -73362 1482 -73323
rect 1680 -73323 1740 -72956
rect 1936 -73064 1942 -73004
rect 2002 -73064 2008 -73004
rect 1808 -73176 1814 -73116
rect 1874 -73176 1880 -73116
rect 1814 -73224 1874 -73176
rect 1787 -73230 1895 -73224
rect 1787 -73264 1799 -73230
rect 1883 -73264 1895 -73230
rect 1787 -73270 1895 -73264
rect 1471 -73666 1477 -73362
rect 1680 -73376 1695 -73323
rect 1689 -73654 1695 -73376
rect 1471 -73699 1486 -73666
rect 1271 -73758 1379 -73752
rect 1271 -73792 1283 -73758
rect 1367 -73792 1379 -73758
rect 1271 -73798 1379 -73792
rect 1296 -73966 1356 -73798
rect 1426 -73852 1486 -73699
rect 1678 -73699 1695 -73654
rect 1729 -73376 1740 -73323
rect 1942 -73323 2002 -73064
rect 2066 -73118 2126 -72772
rect 2200 -73118 2260 -72772
rect 2534 -72906 2646 -72772
rect 4310 -72666 6646 -72660
rect 4310 -72766 4416 -72666
rect 6540 -72766 6646 -72666
rect 4310 -72772 6646 -72766
rect 4310 -72866 4422 -72772
rect 2346 -73064 2352 -73004
rect 2412 -73064 2418 -73004
rect 2066 -73178 2260 -73118
rect 2066 -73224 2126 -73178
rect 2045 -73230 2153 -73224
rect 2045 -73264 2057 -73230
rect 2141 -73264 2153 -73230
rect 2045 -73270 2153 -73264
rect 1729 -73654 1735 -73376
rect 1942 -73400 1953 -73323
rect 1729 -73699 1738 -73654
rect 1529 -73758 1637 -73752
rect 1529 -73792 1541 -73758
rect 1625 -73792 1637 -73758
rect 1529 -73798 1637 -73792
rect 1420 -73912 1426 -73852
rect 1486 -73912 1492 -73852
rect 1554 -73966 1614 -73798
rect 1290 -74026 1296 -73966
rect 1356 -74026 1362 -73966
rect 1548 -74026 1554 -73966
rect 1614 -74026 1620 -73966
rect 1271 -74090 1379 -74084
rect 1271 -74124 1283 -74090
rect 1367 -74124 1379 -74090
rect 1271 -74130 1379 -74124
rect 1529 -74090 1637 -74084
rect 1529 -74124 1541 -74090
rect 1625 -74124 1637 -74090
rect 1529 -74130 1637 -74124
rect 1166 -74559 1179 -74183
rect 1213 -74559 1226 -74183
rect 1431 -74183 1477 -74171
rect 1431 -74526 1437 -74183
rect 1013 -74618 1121 -74612
rect 1013 -74652 1025 -74618
rect 1109 -74652 1121 -74618
rect 1013 -74658 1121 -74652
rect 902 -74928 908 -74868
rect 968 -74928 974 -74868
rect 1166 -74922 1226 -74559
rect 1422 -74559 1437 -74526
rect 1471 -74526 1477 -74183
rect 1678 -74183 1738 -73699
rect 1947 -73699 1953 -73400
rect 1987 -73400 2002 -73323
rect 2200 -73323 2260 -73178
rect 1987 -73699 1993 -73400
rect 1947 -73711 1993 -73699
rect 2200 -73699 2211 -73323
rect 2245 -73699 2260 -73323
rect 1787 -73758 1895 -73752
rect 1787 -73792 1799 -73758
rect 1883 -73792 1895 -73758
rect 1787 -73798 1895 -73792
rect 2045 -73758 2153 -73752
rect 2045 -73792 2057 -73758
rect 2141 -73792 2153 -73758
rect 2045 -73798 2153 -73792
rect 1936 -73912 1942 -73852
rect 2002 -73912 2008 -73852
rect 2068 -73908 2128 -73798
rect 2200 -73908 2260 -73699
rect 1806 -74026 1812 -73966
rect 1872 -74026 1878 -73966
rect 1812 -74084 1872 -74026
rect 1787 -74090 1895 -74084
rect 1787 -74124 1799 -74090
rect 1883 -74124 1895 -74090
rect 1787 -74130 1895 -74124
rect 1678 -74240 1695 -74183
rect 1689 -74498 1695 -74240
rect 1471 -74559 1482 -74526
rect 1271 -74618 1379 -74612
rect 1271 -74652 1283 -74618
rect 1367 -74652 1379 -74618
rect 1271 -74658 1379 -74652
rect 1294 -74690 1354 -74658
rect 1288 -74750 1294 -74690
rect 1354 -74750 1360 -74690
rect 1422 -74810 1482 -74559
rect 1684 -74559 1695 -74498
rect 1729 -74240 1738 -74183
rect 1942 -74183 2002 -73912
rect 2068 -73968 2260 -73908
rect 2045 -74090 2153 -74084
rect 2045 -74124 2057 -74090
rect 2141 -74124 2153 -74090
rect 2045 -74130 2153 -74124
rect 1942 -74232 1953 -74183
rect 1729 -74498 1735 -74240
rect 1729 -74559 1744 -74498
rect 1529 -74618 1637 -74612
rect 1529 -74652 1541 -74618
rect 1625 -74652 1637 -74618
rect 1529 -74658 1637 -74652
rect 1550 -74690 1610 -74658
rect 1544 -74750 1550 -74690
rect 1610 -74750 1616 -74690
rect 1416 -74870 1422 -74810
rect 1482 -74870 1488 -74810
rect 1684 -74922 1744 -74559
rect 1947 -74559 1953 -74232
rect 1987 -74232 2002 -74183
rect 2200 -74183 2260 -73968
rect 1987 -74559 1993 -74232
rect 1947 -74571 1993 -74559
rect 2200 -74559 2211 -74183
rect 2245 -74559 2260 -74183
rect 1787 -74618 1895 -74612
rect 1787 -74652 1799 -74618
rect 1883 -74652 1895 -74618
rect 1787 -74658 1895 -74652
rect 2045 -74618 2153 -74612
rect 2045 -74652 2057 -74618
rect 2141 -74652 2153 -74618
rect 2045 -74658 2153 -74652
rect 2072 -74730 2132 -74658
rect 2200 -74730 2260 -74559
rect 2072 -74790 2260 -74730
rect 1160 -74982 1166 -74922
rect 1226 -74982 1232 -74922
rect 1678 -74982 1684 -74922
rect 1744 -74982 1750 -74922
rect 2072 -75066 2132 -74790
rect 2200 -75066 2260 -74790
rect 2352 -74810 2412 -73064
rect 2346 -74870 2352 -74810
rect 2412 -74870 2418 -74810
rect 578 -75096 2480 -75066
rect 578 -75160 612 -75096
rect 2436 -75160 2480 -75096
rect 578 -75190 2480 -75160
rect 310 -75664 422 -75530
rect 1022 -75664 1032 -75364
rect 1924 -75664 1934 -75364
rect 2534 -75530 2540 -72906
rect 2640 -75530 2646 -72906
rect 3928 -72897 4422 -72866
rect 3928 -72931 3957 -72897
rect 3991 -72931 4049 -72897
rect 4083 -72931 4141 -72897
rect 4175 -72906 4422 -72897
rect 4175 -72931 4316 -72906
rect 3928 -72962 4316 -72931
rect 2534 -75664 2646 -75530
rect 310 -75670 2646 -75664
rect 310 -75770 416 -75670
rect 2540 -75770 2646 -75670
rect 310 -75776 2646 -75770
rect 4310 -75530 4316 -72962
rect 4416 -75530 4422 -72906
rect 5416 -72916 5422 -72856
rect 5482 -72916 5488 -72856
rect 4900 -73064 4906 -73004
rect 4966 -73064 4972 -73004
rect 4504 -73176 4754 -73116
rect 4814 -73176 4820 -73116
rect 4504 -74096 4564 -73176
rect 4755 -73230 4863 -73224
rect 4755 -73264 4767 -73230
rect 4851 -73264 4863 -73230
rect 4755 -73270 4863 -73264
rect 4657 -73323 4703 -73311
rect 4657 -73646 4663 -73323
rect 4504 -74690 4564 -74156
rect 4652 -73699 4663 -73646
rect 4697 -73646 4703 -73323
rect 4906 -73323 4966 -73064
rect 5032 -73176 5038 -73116
rect 5098 -73176 5104 -73116
rect 5038 -73224 5098 -73176
rect 5013 -73230 5121 -73224
rect 5013 -73264 5025 -73230
rect 5109 -73264 5121 -73230
rect 5013 -73270 5121 -73264
rect 5271 -73230 5379 -73224
rect 5271 -73264 5283 -73230
rect 5367 -73264 5379 -73230
rect 5271 -73270 5379 -73264
rect 4906 -73368 4921 -73323
rect 4697 -73699 4712 -73646
rect 4652 -73900 4712 -73699
rect 4915 -73699 4921 -73368
rect 4955 -73368 4966 -73323
rect 5173 -73323 5219 -73311
rect 5173 -73360 5179 -73323
rect 4955 -73699 4961 -73368
rect 4915 -73711 4961 -73699
rect 5166 -73699 5179 -73360
rect 5213 -73360 5219 -73323
rect 5422 -73323 5482 -72916
rect 5674 -72956 5680 -72896
rect 5740 -72956 5746 -72896
rect 5550 -73224 5610 -73170
rect 5529 -73230 5637 -73224
rect 5529 -73264 5541 -73230
rect 5625 -73264 5637 -73230
rect 5529 -73270 5637 -73264
rect 5213 -73699 5226 -73360
rect 5422 -73362 5437 -73323
rect 5431 -73666 5437 -73362
rect 4755 -73758 4863 -73752
rect 4755 -73792 4767 -73758
rect 4851 -73792 4863 -73758
rect 4755 -73798 4863 -73792
rect 5013 -73758 5121 -73752
rect 5013 -73792 5025 -73758
rect 5109 -73792 5121 -73758
rect 5013 -73798 5121 -73792
rect 4782 -73900 4842 -73798
rect 4652 -73960 4842 -73900
rect 4902 -73912 4908 -73852
rect 4968 -73912 4974 -73852
rect 4652 -74183 4712 -73960
rect 4782 -74084 4842 -73960
rect 4755 -74090 4863 -74084
rect 4755 -74124 4767 -74090
rect 4851 -74124 4863 -74090
rect 4755 -74130 4863 -74124
rect 4652 -74226 4663 -74183
rect 4657 -74526 4663 -74226
rect 4652 -74559 4663 -74526
rect 4697 -74226 4712 -74183
rect 4908 -74183 4968 -73912
rect 5032 -74026 5038 -73966
rect 5098 -74026 5104 -73966
rect 5038 -74084 5098 -74026
rect 5013 -74090 5121 -74084
rect 5013 -74124 5025 -74090
rect 5109 -74124 5121 -74090
rect 5013 -74130 5121 -74124
rect 4697 -74526 4703 -74226
rect 4697 -74559 4712 -74526
rect 4498 -74750 4504 -74690
rect 4564 -74750 4570 -74690
rect 4652 -74742 4712 -74559
rect 4908 -74559 4921 -74183
rect 4955 -74559 4968 -74183
rect 4755 -74618 4863 -74612
rect 4755 -74652 4767 -74618
rect 4851 -74652 4863 -74618
rect 4755 -74658 4863 -74652
rect 4782 -74742 4842 -74658
rect 4652 -74802 4842 -74742
rect 4652 -75066 4712 -74802
rect 4782 -75066 4842 -74802
rect 4908 -74866 4968 -74559
rect 5166 -74183 5226 -73699
rect 5426 -73699 5437 -73666
rect 5471 -73362 5482 -73323
rect 5680 -73323 5740 -72956
rect 5936 -73064 5942 -73004
rect 6002 -73064 6008 -73004
rect 5808 -73176 5814 -73116
rect 5874 -73176 5880 -73116
rect 5814 -73224 5874 -73176
rect 5787 -73230 5895 -73224
rect 5787 -73264 5799 -73230
rect 5883 -73264 5895 -73230
rect 5787 -73270 5895 -73264
rect 5471 -73666 5477 -73362
rect 5680 -73376 5695 -73323
rect 5689 -73654 5695 -73376
rect 5471 -73699 5486 -73666
rect 5271 -73758 5379 -73752
rect 5271 -73792 5283 -73758
rect 5367 -73792 5379 -73758
rect 5271 -73798 5379 -73792
rect 5296 -73966 5356 -73798
rect 5426 -73852 5486 -73699
rect 5678 -73699 5695 -73654
rect 5729 -73376 5740 -73323
rect 5942 -73323 6002 -73064
rect 6066 -73118 6126 -72772
rect 6200 -73118 6260 -72772
rect 6534 -72906 6646 -72772
rect 6346 -73064 6352 -73004
rect 6412 -73064 6418 -73004
rect 6066 -73178 6260 -73118
rect 6066 -73224 6126 -73178
rect 6045 -73230 6153 -73224
rect 6045 -73264 6057 -73230
rect 6141 -73264 6153 -73230
rect 6045 -73270 6153 -73264
rect 5729 -73654 5735 -73376
rect 5942 -73400 5953 -73323
rect 5729 -73699 5738 -73654
rect 5529 -73758 5637 -73752
rect 5529 -73792 5541 -73758
rect 5625 -73792 5637 -73758
rect 5529 -73798 5637 -73792
rect 5420 -73912 5426 -73852
rect 5486 -73912 5492 -73852
rect 5554 -73966 5614 -73798
rect 5290 -74026 5296 -73966
rect 5356 -74026 5362 -73966
rect 5548 -74026 5554 -73966
rect 5614 -74026 5620 -73966
rect 5271 -74090 5379 -74084
rect 5271 -74124 5283 -74090
rect 5367 -74124 5379 -74090
rect 5271 -74130 5379 -74124
rect 5529 -74090 5637 -74084
rect 5529 -74124 5541 -74090
rect 5625 -74124 5637 -74090
rect 5529 -74130 5637 -74124
rect 5166 -74559 5179 -74183
rect 5213 -74559 5226 -74183
rect 5431 -74183 5477 -74171
rect 5431 -74526 5437 -74183
rect 5013 -74618 5121 -74612
rect 5013 -74652 5025 -74618
rect 5109 -74652 5121 -74618
rect 5013 -74658 5121 -74652
rect 4902 -74926 4908 -74866
rect 4968 -74926 4974 -74866
rect 5166 -74922 5226 -74559
rect 5422 -74559 5437 -74526
rect 5471 -74526 5477 -74183
rect 5678 -74183 5738 -73699
rect 5947 -73699 5953 -73400
rect 5987 -73400 6002 -73323
rect 6200 -73323 6260 -73178
rect 5987 -73699 5993 -73400
rect 5947 -73711 5993 -73699
rect 6200 -73699 6211 -73323
rect 6245 -73699 6260 -73323
rect 5787 -73758 5895 -73752
rect 5787 -73792 5799 -73758
rect 5883 -73792 5895 -73758
rect 5787 -73798 5895 -73792
rect 6045 -73758 6153 -73752
rect 6045 -73792 6057 -73758
rect 6141 -73792 6153 -73758
rect 6045 -73798 6153 -73792
rect 5936 -73912 5942 -73852
rect 6002 -73912 6008 -73852
rect 6068 -73908 6128 -73798
rect 6200 -73908 6260 -73699
rect 5806 -74026 5812 -73966
rect 5872 -74026 5878 -73966
rect 5812 -74084 5872 -74026
rect 5787 -74090 5895 -74084
rect 5787 -74124 5799 -74090
rect 5883 -74124 5895 -74090
rect 5787 -74130 5895 -74124
rect 5678 -74240 5695 -74183
rect 5689 -74498 5695 -74240
rect 5471 -74559 5482 -74526
rect 5271 -74618 5379 -74612
rect 5271 -74652 5283 -74618
rect 5367 -74652 5379 -74618
rect 5271 -74658 5379 -74652
rect 5294 -74690 5354 -74658
rect 5288 -74750 5294 -74690
rect 5354 -74750 5360 -74690
rect 5422 -74810 5482 -74559
rect 5684 -74559 5695 -74498
rect 5729 -74240 5738 -74183
rect 5942 -74183 6002 -73912
rect 6068 -73968 6260 -73908
rect 6045 -74090 6153 -74084
rect 6045 -74124 6057 -74090
rect 6141 -74124 6153 -74090
rect 6045 -74130 6153 -74124
rect 5942 -74232 5953 -74183
rect 5729 -74498 5735 -74240
rect 5729 -74559 5744 -74498
rect 5529 -74618 5637 -74612
rect 5529 -74652 5541 -74618
rect 5625 -74652 5637 -74618
rect 5529 -74658 5637 -74652
rect 5550 -74690 5610 -74658
rect 5544 -74750 5550 -74690
rect 5610 -74750 5616 -74690
rect 5416 -74870 5422 -74810
rect 5482 -74870 5488 -74810
rect 5684 -74922 5744 -74559
rect 5947 -74559 5953 -74232
rect 5987 -74232 6002 -74183
rect 6200 -74183 6260 -73968
rect 5987 -74559 5993 -74232
rect 5947 -74571 5993 -74559
rect 6200 -74559 6211 -74183
rect 6245 -74559 6260 -74183
rect 5787 -74618 5895 -74612
rect 5787 -74652 5799 -74618
rect 5883 -74652 5895 -74618
rect 5787 -74658 5895 -74652
rect 6045 -74618 6153 -74612
rect 6045 -74652 6057 -74618
rect 6141 -74652 6153 -74618
rect 6045 -74658 6153 -74652
rect 6072 -74730 6132 -74658
rect 6200 -74730 6260 -74559
rect 6072 -74790 6260 -74730
rect 5160 -74982 5166 -74922
rect 5226 -74982 5232 -74922
rect 5678 -74982 5684 -74922
rect 5744 -74982 5750 -74922
rect 6072 -75066 6132 -74790
rect 6200 -75066 6260 -74790
rect 6352 -74810 6412 -73064
rect 6346 -74870 6352 -74810
rect 6412 -74870 6418 -74810
rect 4578 -75096 6480 -75066
rect 4578 -75160 4612 -75096
rect 6436 -75160 6480 -75096
rect 4578 -75190 6480 -75160
rect 4310 -75664 4422 -75530
rect 5022 -75664 5032 -75364
rect 5924 -75664 5934 -75364
rect 6534 -75530 6540 -72906
rect 6640 -75530 6646 -72906
rect 6534 -75664 6646 -75530
rect 4310 -75670 6646 -75664
rect 4310 -75770 4416 -75670
rect 6540 -75770 6646 -75670
rect 4310 -75776 6646 -75770
<< via1 >>
rect 25928 -28062 26528 -27762
rect 49560 -28062 50160 -27762
rect 29505 -28358 46290 -28144
rect 33430 -30120 33490 -30060
rect 34512 -30120 34572 -30060
rect 35470 -30120 35530 -30060
rect 33956 -30366 34016 -30306
rect 35992 -30366 36052 -30306
rect 31774 -31298 31834 -31238
rect 32938 -31298 32998 -31238
rect 31644 -31502 31704 -31442
rect 29636 -33686 29696 -33626
rect 32938 -31502 32998 -31442
rect 38534 -30120 38594 -30060
rect 39552 -30120 39612 -30060
rect 38030 -30364 38090 -30304
rect 34974 -31402 35034 -31342
rect 33424 -32652 33484 -32592
rect 40576 -30120 40636 -30060
rect 41588 -30120 41648 -30060
rect 40060 -30364 40120 -30304
rect 37010 -31402 37070 -31342
rect 42102 -30362 42162 -30302
rect 39048 -31298 39108 -31238
rect 39044 -31502 39104 -31442
rect 35480 -32436 35540 -32376
rect 35990 -32436 36050 -32376
rect 34972 -32538 35036 -32474
rect 34462 -32652 34522 -32592
rect 35474 -32652 35534 -32592
rect 31774 -33972 31834 -33912
rect 32130 -36380 32190 -36320
rect 32004 -36990 32064 -36930
rect 29120 -37944 29180 -37884
rect 29228 -38056 29288 -37996
rect 27458 -38978 27518 -38918
rect 30142 -37944 30202 -37884
rect 30012 -38056 30072 -37996
rect 28618 -39088 28678 -39028
rect 30652 -38978 30712 -38918
rect 27332 -40066 27392 -40006
rect 29134 -40012 29194 -39952
rect 29240 -40112 29300 -40052
rect 31804 -39088 31864 -39028
rect 30144 -40012 30204 -39952
rect 31996 -39216 32056 -39156
rect 30026 -40112 30086 -40052
rect 26846 -41122 26906 -41062
rect 26986 -41298 27046 -41238
rect 30132 -41300 30192 -41240
rect 27886 -41472 27946 -41412
rect 32246 -36990 32306 -36930
rect 32932 -33826 32996 -33762
rect 32756 -33972 32816 -33912
rect 36848 -32538 36912 -32474
rect 43112 -30362 43172 -30302
rect 44646 -30120 44706 -30060
rect 45658 -30120 45718 -30060
rect 44134 -30362 44194 -30302
rect 41082 -31298 41142 -31238
rect 41080 -31502 41140 -31442
rect 41582 -31502 41642 -31442
rect 38024 -32436 38084 -32376
rect 36484 -32644 36544 -32584
rect 37508 -32644 37568 -32584
rect 33954 -33574 34014 -33514
rect 34970 -33688 35034 -33624
rect 38536 -32644 38596 -32584
rect 46676 -30120 46736 -30060
rect 46170 -30362 46230 -30302
rect 43116 -31402 43176 -31342
rect 42602 -31502 42662 -31442
rect 40062 -32438 40122 -32378
rect 35990 -33574 36050 -33514
rect 36512 -33574 36572 -33514
rect 37010 -33574 37070 -33514
rect 43628 -31502 43688 -31442
rect 45150 -31402 45210 -31342
rect 44134 -31506 44194 -31446
rect 44648 -31506 44708 -31446
rect 45152 -31506 45212 -31446
rect 45658 -31506 45718 -31446
rect 46178 -31506 46238 -31446
rect 41082 -32536 41142 -32476
rect 47190 -31298 47250 -31238
rect 48440 -31298 48500 -31238
rect 42098 -32438 42158 -32378
rect 42598 -32438 42658 -32378
rect 43112 -32438 43172 -32378
rect 43636 -32438 43696 -32378
rect 44134 -32438 44194 -32378
rect 44636 -32438 44696 -32378
rect 37484 -33578 37544 -33518
rect 32872 -34078 32932 -34018
rect 33434 -34078 33494 -34018
rect 34476 -34078 34536 -34018
rect 35476 -34078 35536 -34018
rect 38024 -33516 38084 -33514
rect 37992 -33574 38084 -33516
rect 38484 -33574 38544 -33514
rect 37992 -33576 38052 -33574
rect 39042 -33830 39106 -33766
rect 39528 -33572 39588 -33512
rect 38638 -34078 38698 -34018
rect 40060 -33574 40120 -33514
rect 45150 -32440 45210 -32380
rect 45658 -32440 45718 -32380
rect 46168 -32440 46228 -32380
rect 44640 -32652 44700 -32592
rect 45652 -32652 45712 -32592
rect 41572 -33572 41632 -33512
rect 41078 -33972 41142 -33908
rect 39648 -34078 39708 -34018
rect 40590 -34078 40650 -34018
rect 42098 -33518 42158 -33516
rect 42066 -33576 42158 -33518
rect 42066 -33578 42126 -33576
rect 42594 -33582 42654 -33522
rect 43082 -33520 43142 -33518
rect 43082 -33578 43176 -33520
rect 43116 -33580 43176 -33578
rect 47190 -32536 47250 -32476
rect 46654 -32652 46714 -32592
rect 43594 -33582 43654 -33522
rect 44134 -33578 44194 -33518
rect 46168 -33578 46228 -33518
rect 45150 -33688 45214 -33624
rect 48436 -33826 48500 -33762
rect 47184 -33972 47244 -33912
rect 32986 -34280 33046 -34220
rect 36164 -34280 36224 -34220
rect 34130 -35216 34190 -35156
rect 34634 -35324 34694 -35264
rect 36164 -35216 36224 -35156
rect 35656 -35324 35716 -35264
rect 36674 -35324 36734 -35264
rect 34126 -36248 34186 -36188
rect 34632 -36382 34692 -36322
rect 40232 -34280 40292 -34220
rect 38206 -35216 38266 -35156
rect 37698 -35324 37758 -35264
rect 38712 -35324 38772 -35264
rect 35646 -36386 35706 -36326
rect 36678 -36378 36738 -36318
rect 40232 -35216 40292 -35156
rect 39730 -35324 39790 -35264
rect 40740 -35324 40800 -35264
rect 38206 -36248 38266 -36188
rect 37676 -36378 37736 -36318
rect 38720 -36378 38780 -36318
rect 44308 -34280 44368 -34220
rect 42274 -35216 42334 -35156
rect 41762 -35324 41822 -35264
rect 42776 -35324 42836 -35264
rect 39724 -36382 39784 -36322
rect 40740 -36382 40800 -36322
rect 39524 -36590 39584 -36530
rect 32756 -36908 32816 -36848
rect 33922 -36908 33982 -36848
rect 32488 -37954 32548 -37894
rect 32246 -39112 32306 -39052
rect 32242 -39326 32302 -39266
rect 32130 -40368 32190 -40308
rect 26726 -41622 26786 -41562
rect 27780 -41884 27840 -41824
rect 30132 -41882 30192 -41822
rect 32624 -38052 32684 -37992
rect 32488 -41626 32548 -41566
rect 35958 -36908 36018 -36848
rect 36466 -36912 36530 -36848
rect 34940 -37856 35000 -37796
rect 47504 -34280 47564 -34220
rect 44310 -35216 44370 -35156
rect 43808 -35324 43868 -35264
rect 44818 -35324 44878 -35264
rect 42274 -36248 42334 -36188
rect 41744 -36382 41804 -36322
rect 42776 -36378 42836 -36318
rect 41260 -36590 41320 -36530
rect 40540 -36790 40604 -36726
rect 46346 -35216 46406 -35156
rect 45840 -35324 45900 -35264
rect 43792 -36382 43852 -36322
rect 44820 -36382 44880 -36322
rect 46342 -36248 46402 -36188
rect 45840 -36382 45900 -36322
rect 48298 -36380 48358 -36320
rect 47158 -36606 47218 -36546
rect 44604 -36790 44668 -36726
rect 45628 -36790 45692 -36726
rect 46640 -36790 46704 -36726
rect 40542 -36912 40606 -36848
rect 36976 -37856 37036 -37796
rect 37318 -37854 37378 -37794
rect 34940 -38052 35000 -37992
rect 35960 -38050 36020 -37990
rect 33926 -38162 33986 -38102
rect 35960 -38162 36020 -38102
rect 32908 -39326 32968 -39266
rect 40032 -37854 40092 -37794
rect 44104 -36908 44164 -36848
rect 46138 -36908 46198 -36848
rect 41050 -38050 41110 -37990
rect 39016 -38164 39076 -38104
rect 41050 -38164 41110 -38104
rect 34942 -39216 35002 -39156
rect 34942 -39420 35002 -39360
rect 36978 -39216 37038 -39156
rect 36976 -39318 37036 -39258
rect 36976 -39420 37036 -39360
rect 33924 -40368 33984 -40308
rect 32756 -40576 32816 -40516
rect 34938 -40678 34998 -40618
rect 39012 -39112 39072 -39052
rect 35960 -40368 36020 -40308
rect 35960 -40476 36020 -40416
rect 40032 -39112 40092 -39052
rect 40032 -39418 40092 -39358
rect 44106 -38164 44166 -38104
rect 41050 -39418 41110 -39358
rect 45120 -37856 45180 -37796
rect 46140 -38164 46200 -38104
rect 47156 -37856 47216 -37796
rect 42068 -39112 42128 -39052
rect 42066 -39418 42126 -39358
rect 36978 -40360 37038 -40300
rect 38780 -40360 38840 -40300
rect 36972 -40678 37032 -40618
rect 37176 -40690 37236 -40630
rect 33920 -41626 33980 -41566
rect 39014 -40366 39074 -40306
rect 44102 -39216 44162 -39156
rect 44970 -39098 45030 -39038
rect 45118 -39208 45178 -39148
rect 44970 -39418 45030 -39358
rect 45122 -39416 45182 -39356
rect 41050 -40366 41110 -40306
rect 41048 -40476 41108 -40416
rect 35956 -41626 36016 -41566
rect 32624 -41756 32684 -41696
rect 27660 -42002 27720 -41942
rect 40538 -40690 40598 -40630
rect 46138 -39318 46198 -39258
rect 48734 -36248 48794 -36188
rect 48440 -36608 48500 -36548
rect 48582 -36908 48642 -36848
rect 48422 -38050 48482 -37990
rect 47158 -39208 47218 -39148
rect 48298 -39208 48358 -39148
rect 47156 -39416 47216 -39356
rect 41554 -40690 41614 -40630
rect 44104 -40364 44164 -40304
rect 44614 -40690 44674 -40630
rect 45126 -40678 45186 -40618
rect 46140 -40364 46200 -40304
rect 48422 -39416 48482 -39356
rect 48298 -40476 48358 -40416
rect 47160 -40678 47220 -40618
rect 44108 -41626 44168 -41566
rect 46144 -41626 46204 -41566
rect 36978 -41896 37038 -41836
rect 48734 -38164 48794 -38104
rect 48582 -41896 48642 -41836
rect 27214 -42120 27274 -42060
rect 52262 -39386 55130 -39086
rect 53114 -40077 53174 -40017
rect 52380 -40434 52440 -40374
rect 53264 -40316 53324 -40256
rect 53134 -40434 53194 -40374
rect 53392 -40434 53452 -40374
rect 52878 -41166 52938 -41106
rect 52748 -41286 52808 -41226
rect 53132 -41166 53192 -41106
rect 53392 -41166 53452 -41106
rect 53262 -41286 53322 -41226
rect 52380 -42022 52440 -41962
rect 54294 -40316 54354 -40256
rect 54166 -40434 54226 -40374
rect 53650 -41166 53710 -41106
rect 54426 -40434 54486 -40374
rect 53908 -41166 53968 -41106
rect 53778 -41286 53838 -41226
rect 55186 -40316 55246 -40256
rect 55004 -40434 55064 -40374
rect 54166 -41166 54226 -41106
rect 54424 -41166 54484 -41106
rect 54294 -41286 54354 -41226
rect 52874 -42022 52934 -41962
rect 53650 -42022 53710 -41962
rect 52746 -42138 52806 -42078
rect 54682 -41166 54742 -41106
rect 54806 -41286 54866 -41226
rect 53906 -42022 53966 -41962
rect 54678 -42022 54738 -41962
rect 53778 -42140 53838 -42080
rect 54808 -42140 54868 -42080
rect 55186 -42140 55246 -42080
rect 55732 -40604 55792 -40544
rect 55586 -41286 55646 -41226
rect 11814 -42648 22578 -42356
rect 53914 -42428 53974 -42368
rect 54200 -42482 54260 -42476
rect 54200 -42542 54206 -42482
rect 54206 -42542 54260 -42482
rect 54200 -42548 54260 -42542
rect 55295 -42477 55365 -42471
rect 55295 -42547 55359 -42477
rect 55359 -42547 55365 -42477
rect 55295 -42553 55365 -42547
rect 54332 -42782 54346 -42736
rect 54346 -42782 54380 -42736
rect 54380 -42782 54392 -42736
rect 54332 -42796 54392 -42782
rect 54588 -42782 54602 -42726
rect 54602 -42782 54636 -42726
rect 54636 -42782 54648 -42726
rect 54588 -42786 54648 -42782
rect 54846 -42776 54858 -42716
rect 54858 -42776 54892 -42716
rect 54892 -42776 54906 -42716
rect 55098 -42778 55114 -42718
rect 55114 -42778 55148 -42718
rect 55148 -42778 55158 -42718
rect 55232 -42776 55242 -42716
rect 55242 -42776 55276 -42716
rect 55276 -42776 55292 -42716
rect 54332 -43108 54392 -43048
rect 54588 -43106 54648 -43046
rect 54846 -43106 54906 -43046
rect 55098 -43106 55158 -43046
rect 56534 -39386 58154 -39086
rect 56318 -39726 56378 -39666
rect 56704 -39726 56764 -39666
rect 56962 -39726 57022 -39666
rect 56318 -40604 56378 -40544
rect 56442 -40604 56502 -40544
rect 57346 -39726 57406 -39666
rect 56704 -40604 56764 -40544
rect 56832 -40604 56892 -40544
rect 56958 -40604 57018 -40544
rect 57986 -39726 58046 -39666
rect 57474 -40536 57534 -40476
rect 57216 -40604 57276 -40544
rect 57346 -40604 57406 -40544
rect 56438 -41358 56498 -41298
rect 56828 -41358 56888 -41298
rect 57216 -41358 57276 -41298
rect 57986 -41358 58046 -41298
rect 58256 -41650 58316 -41590
rect 57136 -41886 57196 -41874
rect 57136 -41920 57152 -41886
rect 57152 -41920 57186 -41886
rect 57186 -41920 57196 -41886
rect 57136 -41934 57196 -41920
rect 56856 -41990 56916 -41984
rect 56856 -42038 56862 -41990
rect 56862 -42038 56910 -41990
rect 56910 -42038 56916 -41990
rect 56856 -42044 56916 -42038
rect 57134 -41990 57194 -41984
rect 57134 -42038 57142 -41990
rect 57142 -42038 57190 -41990
rect 57190 -42038 57194 -41990
rect 57134 -42044 57194 -42038
rect 56042 -42630 56142 -42572
rect 56042 -42664 56075 -42630
rect 56075 -42664 56109 -42630
rect 56109 -42664 56142 -42630
rect 56042 -42672 56142 -42664
rect 55732 -43018 55792 -42958
rect 55586 -43126 55646 -43066
rect 56004 -43018 56064 -42958
rect 56120 -43018 56180 -42958
rect 27332 -43396 27392 -43336
rect 27660 -43386 27720 -43326
rect 26726 -43532 26786 -43472
rect 26846 -43530 26906 -43470
rect 26986 -43512 27046 -43452
rect 27214 -43496 27274 -43436
rect 26594 -43660 26654 -43600
rect 9372 -57518 9436 -56724
rect 11560 -56780 11620 -56720
rect 10912 -57546 10972 -57486
rect 10654 -57695 10714 -57635
rect 11430 -57546 11490 -57486
rect 11170 -57695 11230 -57635
rect 12176 -57592 12236 -57532
rect 12524 -57592 12584 -57532
rect 11688 -57695 11748 -57635
rect 10914 -58134 10974 -58074
rect 11430 -58134 11490 -58074
rect 11558 -58243 11618 -58183
rect 23882 -44258 23942 -44198
rect 25408 -44392 25468 -44332
rect 26594 -50860 26654 -50800
rect 22046 -51786 22106 -51726
rect 15936 -51932 15996 -51872
rect 20016 -51932 20076 -51872
rect 14782 -52060 14842 -52000
rect 17460 -52060 17520 -52000
rect 18492 -52060 18552 -52000
rect 14762 -53048 14862 -52948
rect 16440 -53022 16500 -52962
rect 15940 -53126 16000 -53066
rect 14764 -54042 14864 -53942
rect 17464 -53022 17524 -52962
rect 16958 -53230 17018 -53170
rect 14782 -54292 14842 -54232
rect 14764 -55048 14864 -54948
rect 21552 -52060 21612 -52000
rect 18496 -53022 18556 -52962
rect 17976 -53126 18036 -53066
rect 24076 -51932 24136 -51872
rect 26260 -51932 26320 -51872
rect 22548 -52060 22608 -52000
rect 19496 -53022 19556 -52962
rect 20516 -53022 20576 -52962
rect 20012 -53126 20072 -53066
rect 18994 -53230 19054 -53170
rect 16432 -54292 16492 -54232
rect 17970 -54172 18030 -54112
rect 21536 -53022 21596 -52962
rect 21026 -53230 21086 -53170
rect 19502 -54292 19562 -54232
rect 22546 -53022 22606 -52962
rect 22046 -53126 22106 -53066
rect 23560 -53022 23620 -52962
rect 24578 -53022 24638 -52962
rect 24082 -53126 24142 -53066
rect 23060 -53230 23120 -53170
rect 20510 -54292 20570 -54232
rect 16958 -55236 17018 -55176
rect 15944 -55344 16004 -55284
rect 16438 -55456 16498 -55396
rect 17980 -55344 18040 -55284
rect 17462 -55456 17522 -55396
rect 22046 -54172 22106 -54112
rect 18994 -55236 19054 -55176
rect 18494 -55456 18554 -55396
rect 25104 -53230 25164 -53170
rect 23572 -54292 23632 -54232
rect 26380 -53022 26440 -52962
rect 26380 -53624 26440 -53564
rect 26260 -54172 26320 -54112
rect 24598 -54292 24658 -54232
rect 21026 -55236 21086 -55176
rect 20016 -55344 20076 -55284
rect 19494 -55456 19554 -55396
rect 20514 -55456 20574 -55396
rect 22050 -55344 22110 -55284
rect 21534 -55456 21594 -55396
rect 14782 -56418 14842 -56358
rect 17452 -56418 17512 -56358
rect 18484 -56418 18544 -56358
rect 22544 -55456 22604 -55396
rect 23060 -55236 23120 -55176
rect 25104 -55236 25164 -55176
rect 24086 -55344 24146 -55284
rect 23558 -55456 23618 -55396
rect 24576 -55456 24636 -55396
rect 21544 -56418 21604 -56358
rect 22540 -56418 22600 -56358
rect 26380 -55456 26440 -55396
rect 15938 -56548 15998 -56488
rect 20018 -56548 20078 -56488
rect 24078 -56548 24138 -56488
rect 26260 -56548 26320 -56488
rect 17416 -57914 17476 -57854
rect 10294 -58514 12110 -58408
rect 19454 -57914 19514 -57854
rect 21490 -57914 21550 -57854
rect 18434 -58026 18494 -57966
rect 23526 -57914 23586 -57854
rect 22508 -58026 22568 -57966
rect 26726 -51932 26786 -51872
rect 27104 -43650 27164 -43590
rect 26986 -45164 27046 -45104
rect 26986 -46920 27046 -46860
rect 26986 -48434 27046 -48374
rect 26982 -49676 27042 -49616
rect 27214 -44392 27274 -44332
rect 27780 -43394 27840 -43334
rect 27660 -44258 27720 -44198
rect 27886 -43530 27946 -43470
rect 27780 -45164 27840 -45104
rect 27456 -45616 27516 -45556
rect 27330 -47318 27390 -47258
rect 27104 -49778 27164 -49718
rect 26986 -50912 27046 -50852
rect 26846 -52060 26906 -52000
rect 26986 -53022 27046 -52962
rect 27668 -45952 27728 -45892
rect 27564 -47212 27624 -47152
rect 27456 -48312 27516 -48252
rect 38698 -43880 38758 -43820
rect 43802 -43880 43862 -43820
rect 47862 -43886 47922 -43826
rect 29030 -45616 29090 -45556
rect 56608 -42562 56668 -42502
rect 56666 -43128 56726 -43068
rect 56918 -42874 56978 -42868
rect 56918 -42922 56924 -42874
rect 56924 -42922 56972 -42874
rect 56972 -42922 56978 -42874
rect 56918 -42928 56978 -42922
rect 57138 -42874 57198 -42868
rect 57138 -42922 57144 -42874
rect 57144 -42922 57192 -42874
rect 57192 -42922 57198 -42874
rect 57138 -42928 57198 -42922
rect 57374 -43128 57434 -43068
rect 57946 -42630 58046 -42574
rect 57946 -42664 57979 -42630
rect 57979 -42664 58013 -42630
rect 58013 -42664 58046 -42630
rect 57946 -42674 58046 -42664
rect 58024 -43028 58084 -42968
rect 57904 -43128 57964 -43068
rect 58256 -43028 58316 -42968
rect 55824 -43563 56370 -43278
rect 56370 -43563 56470 -43278
rect 56470 -43563 57628 -43278
rect 57628 -43563 57728 -43278
rect 57728 -43563 58268 -43278
rect 55824 -43584 58268 -43563
rect 30044 -45832 30104 -45772
rect 32084 -45832 32144 -45772
rect 34124 -45832 34184 -45772
rect 36154 -45832 36214 -45772
rect 38194 -45832 38254 -45772
rect 40226 -45832 40286 -45772
rect 42266 -45832 42326 -45772
rect 44302 -45832 44362 -45772
rect 46336 -45832 46396 -45772
rect 28012 -45952 28072 -45892
rect 29536 -45958 29596 -45898
rect 27886 -46074 27946 -46014
rect 27780 -46920 27840 -46860
rect 30550 -45958 30610 -45898
rect 31572 -45958 31632 -45898
rect 32586 -45958 32646 -45898
rect 33612 -45958 33672 -45898
rect 33100 -46074 33160 -46014
rect 34624 -45958 34684 -45898
rect 35660 -45958 35720 -45898
rect 36666 -45958 36726 -45898
rect 37680 -45958 37740 -45898
rect 30048 -46996 30108 -46936
rect 29540 -47106 29600 -47046
rect 29030 -47212 29090 -47152
rect 28016 -47318 28076 -47258
rect 28514 -47318 28574 -47258
rect 29026 -47318 29086 -47258
rect 30562 -47106 30622 -47046
rect 32088 -46996 32148 -46936
rect 31576 -47106 31636 -47046
rect 31070 -47212 31130 -47152
rect 34120 -46996 34180 -46936
rect 32590 -47106 32650 -47046
rect 33608 -47106 33668 -47046
rect 33100 -47212 33160 -47152
rect 27886 -48208 27946 -48148
rect 28010 -48312 28070 -48252
rect 29530 -48312 29590 -48252
rect 30042 -48312 30102 -48252
rect 27780 -48434 27840 -48374
rect 27668 -48548 27728 -48488
rect 28516 -48548 28576 -48488
rect 30048 -48546 30108 -48486
rect 34634 -47106 34694 -47046
rect 38696 -45958 38756 -45898
rect 39704 -45958 39764 -45898
rect 40720 -45958 40780 -45898
rect 41744 -45958 41804 -45898
rect 42766 -45958 42826 -45898
rect 43788 -45958 43848 -45898
rect 43288 -46074 43348 -46014
rect 36152 -46996 36212 -46936
rect 35140 -47212 35200 -47152
rect 35654 -47106 35714 -47046
rect 35306 -47318 35366 -47258
rect 31064 -48208 31124 -48148
rect 31066 -48312 31126 -48252
rect 36674 -47106 36734 -47046
rect 38188 -46996 38248 -46936
rect 37676 -47106 37736 -47046
rect 37174 -47212 37234 -47152
rect 37174 -47318 37234 -47258
rect 38702 -47106 38762 -47046
rect 44806 -45958 44866 -45898
rect 45820 -45958 45880 -45898
rect 46844 -45958 46904 -45898
rect 47360 -46074 47420 -46014
rect 48492 -46074 48552 -46014
rect 40224 -46996 40284 -46936
rect 39720 -47106 39780 -47046
rect 39210 -47212 39270 -47152
rect 39212 -47318 39272 -47258
rect 40728 -47106 40788 -47046
rect 42262 -46996 42322 -46936
rect 41740 -47106 41800 -47046
rect 41246 -47212 41306 -47152
rect 41092 -47318 41152 -47258
rect 32078 -48312 32138 -48252
rect 32084 -48546 32144 -48486
rect 33098 -48312 33158 -48252
rect 27892 -49476 27952 -49416
rect 29030 -49476 29090 -49416
rect 27780 -49676 27840 -49616
rect 27674 -49778 27734 -49718
rect 27564 -53230 27624 -53170
rect 27780 -50912 27840 -50852
rect 29028 -49676 29088 -49616
rect 30046 -49556 30106 -49496
rect 34120 -48208 34180 -48148
rect 44300 -46996 44360 -46936
rect 42772 -47106 42832 -47046
rect 43786 -47106 43846 -47046
rect 43286 -47212 43346 -47152
rect 40226 -48208 40286 -48148
rect 36156 -48312 36216 -48252
rect 38194 -48312 38254 -48252
rect 35140 -48434 35200 -48374
rect 37174 -48434 37234 -48374
rect 39204 -48434 39264 -48374
rect 31064 -49452 31124 -49392
rect 30560 -49670 30620 -49610
rect 32086 -49556 32146 -49496
rect 31564 -49670 31624 -49610
rect 29028 -50708 29088 -50648
rect 29534 -50810 29594 -50750
rect 33100 -49452 33160 -49392
rect 32576 -49670 32636 -49610
rect 34118 -49556 34178 -49496
rect 33596 -49670 33656 -49610
rect 34118 -49668 34178 -49608
rect 36152 -49556 36212 -49496
rect 35136 -49778 35196 -49718
rect 31066 -50708 31126 -50648
rect 31064 -50912 31124 -50852
rect 36154 -49668 36214 -49608
rect 37170 -49778 37230 -49718
rect 41244 -48312 41304 -48252
rect 44804 -47106 44864 -47046
rect 46336 -46996 46396 -46936
rect 45828 -47106 45888 -47046
rect 45316 -47212 45376 -47152
rect 45316 -47316 45376 -47256
rect 42262 -48312 42322 -48252
rect 43282 -48312 43342 -48252
rect 38192 -49556 38252 -49496
rect 38190 -49668 38250 -49608
rect 40226 -49556 40286 -49496
rect 40422 -49560 40482 -49500
rect 39210 -49778 39270 -49718
rect 40226 -49668 40286 -49608
rect 46848 -47106 46908 -47046
rect 47356 -47212 47416 -47152
rect 48492 -47316 48552 -47256
rect 45320 -48208 45380 -48148
rect 44298 -48312 44358 -48252
rect 46334 -48312 46394 -48252
rect 41244 -49452 41304 -49392
rect 40422 -49778 40482 -49718
rect 40716 -49776 40776 -49716
rect 33102 -50708 33162 -50648
rect 30048 -51012 30108 -50952
rect 31572 -50918 31632 -50858
rect 32594 -50918 32654 -50858
rect 32082 -51012 32142 -50952
rect 35134 -50708 35194 -50648
rect 34626 -50810 34686 -50750
rect 33608 -50918 33668 -50858
rect 34626 -50918 34686 -50858
rect 34118 -51012 34178 -50952
rect 29530 -51936 29590 -51876
rect 30440 -51936 30500 -51876
rect 29530 -52152 29590 -52092
rect 27894 -52256 27954 -52196
rect 27782 -53022 27842 -52962
rect 27332 -53380 27392 -53320
rect 27674 -53268 27734 -53208
rect 27780 -53624 27840 -53564
rect 31442 -51936 31502 -51876
rect 30568 -52152 30628 -52092
rect 32594 -51936 32654 -51876
rect 32082 -52038 32142 -51978
rect 31582 -52152 31642 -52092
rect 29528 -53164 29588 -53104
rect 29030 -53268 29090 -53208
rect 29026 -53478 29086 -53418
rect 30536 -53164 30596 -53104
rect 30046 -53380 30106 -53320
rect 35646 -50918 35706 -50858
rect 42260 -49668 42320 -49608
rect 41744 -49776 41804 -49716
rect 42262 -49782 42322 -49722
rect 43280 -49452 43340 -49392
rect 44298 -49668 44358 -49608
rect 45314 -49560 45374 -49500
rect 45818 -49564 45878 -49504
rect 48478 -48546 48538 -48486
rect 46338 -49668 46398 -49608
rect 44298 -49782 44358 -49722
rect 39716 -50696 39776 -50636
rect 39210 -50824 39270 -50764
rect 41246 -51022 41306 -50962
rect 33604 -51936 33664 -51876
rect 34610 -51936 34670 -51876
rect 35654 -51936 35714 -51876
rect 36154 -51930 36214 -51870
rect 34608 -52152 34668 -52092
rect 35648 -52152 35708 -52092
rect 35132 -52256 35192 -52196
rect 31550 -53164 31610 -53104
rect 32588 -53164 32648 -53104
rect 32084 -53380 32144 -53320
rect 31064 -53478 31124 -53418
rect 36662 -52152 36722 -52092
rect 38190 -51930 38250 -51870
rect 37670 -52152 37730 -52092
rect 38714 -52152 38774 -52092
rect 37174 -52256 37234 -52196
rect 46336 -49782 46396 -49722
rect 42758 -50918 42818 -50858
rect 40226 -51930 40286 -51870
rect 39704 -52152 39764 -52092
rect 40722 -52152 40782 -52092
rect 39212 -52256 39272 -52196
rect 47354 -49452 47414 -49392
rect 48372 -49434 48432 -49374
rect 48606 -48564 48666 -48504
rect 48972 -49564 49032 -49504
rect 48722 -49668 48782 -49608
rect 44810 -50696 44870 -50636
rect 44948 -50692 45008 -50632
rect 48478 -49782 48538 -49722
rect 45830 -50692 45890 -50632
rect 46836 -50692 46896 -50632
rect 43788 -50918 43848 -50858
rect 44948 -50918 45008 -50858
rect 45316 -50918 45376 -50858
rect 45316 -51022 45376 -50962
rect 47354 -50696 47414 -50636
rect 47354 -50824 47414 -50764
rect 46332 -51020 46392 -50960
rect 42264 -51930 42324 -51870
rect 42256 -52038 42316 -51978
rect 41756 -52152 41816 -52092
rect 41246 -52256 41306 -52196
rect 41758 -52260 41818 -52200
rect 42780 -52260 42840 -52200
rect 43280 -52254 43340 -52194
rect 33606 -53164 33666 -53104
rect 34122 -53158 34182 -53098
rect 36158 -53158 36218 -53098
rect 38190 -53158 38250 -53098
rect 40224 -53158 40284 -53098
rect 33104 -53478 33164 -53418
rect 27892 -54500 27952 -54440
rect 29032 -54716 29092 -54656
rect 27780 -55456 27840 -55396
rect 30046 -54402 30106 -54342
rect 30050 -54596 30110 -54536
rect 31064 -54500 31124 -54440
rect 37174 -53268 37234 -53208
rect 39210 -53268 39270 -53208
rect 36156 -53380 36216 -53320
rect 35140 -53478 35200 -53418
rect 32082 -54402 32142 -54342
rect 32588 -54500 32648 -54440
rect 32086 -54596 32146 -54536
rect 34120 -54402 34180 -54342
rect 33610 -54500 33670 -54440
rect 33100 -54716 33160 -54656
rect 27780 -55632 27840 -55572
rect 27674 -55758 27734 -55698
rect 34632 -54500 34692 -54440
rect 34114 -54596 34174 -54536
rect 44300 -51930 44360 -51870
rect 44296 -52038 44356 -51978
rect 44788 -52152 44848 -52092
rect 46338 -51930 46398 -51870
rect 46334 -52038 46394 -51978
rect 45826 -52152 45886 -52092
rect 45314 -52254 45374 -52194
rect 41246 -53156 41306 -53096
rect 41600 -53156 41660 -53096
rect 41242 -53268 41302 -53208
rect 40752 -53366 40812 -53306
rect 35982 -54382 36042 -54322
rect 36152 -54382 36212 -54322
rect 35636 -54500 35696 -54440
rect 35134 -54716 35194 -54656
rect 31064 -55758 31124 -55698
rect 31584 -55746 31644 -55686
rect 30046 -55860 30106 -55800
rect 32082 -55860 32142 -55800
rect 31064 -55964 31124 -55904
rect 27892 -56862 27952 -56802
rect 27564 -56966 27624 -56906
rect 29028 -56966 29088 -56906
rect 29536 -57072 29596 -57012
rect 26514 -58026 26574 -57966
rect 35982 -54596 36042 -54536
rect 36158 -54590 36218 -54530
rect 41790 -53366 41850 -53306
rect 42766 -53366 42826 -53306
rect 41600 -53474 41660 -53414
rect 46852 -52152 46912 -52092
rect 47356 -52254 47416 -52194
rect 45318 -53156 45378 -53096
rect 43782 -53366 43842 -53306
rect 45808 -53366 45868 -53306
rect 43280 -53478 43340 -53418
rect 45316 -53478 45376 -53418
rect 38194 -54382 38254 -54322
rect 40226 -54382 40286 -54322
rect 42266 -54382 42326 -54322
rect 41244 -54480 41304 -54420
rect 38186 -54590 38246 -54530
rect 33102 -55860 33162 -55800
rect 34118 -55860 34178 -55800
rect 31062 -56862 31122 -56802
rect 31068 -56966 31128 -56906
rect 30556 -57072 30616 -57012
rect 30048 -57182 30108 -57122
rect 31580 -57072 31640 -57012
rect 35138 -55860 35198 -55800
rect 40230 -54590 40290 -54530
rect 42258 -54590 42318 -54530
rect 43284 -54716 43344 -54656
rect 46838 -53366 46898 -53306
rect 47352 -53478 47412 -53418
rect 44296 -54590 44356 -54530
rect 47350 -54480 47410 -54420
rect 46336 -54590 46396 -54530
rect 46854 -54586 46914 -54526
rect 48366 -54586 48426 -54526
rect 45314 -54716 45374 -54656
rect 45840 -54714 45900 -54654
rect 37168 -55632 37228 -55572
rect 39210 -55632 39270 -55572
rect 41246 -55632 41306 -55572
rect 36664 -55746 36724 -55686
rect 41752 -55742 41812 -55682
rect 36156 -55860 36216 -55800
rect 38186 -55860 38246 -55800
rect 40224 -55860 40284 -55800
rect 42260 -55860 42320 -55800
rect 36000 -55964 36060 -55904
rect 33098 -56966 33158 -56906
rect 32598 -57072 32658 -57012
rect 33612 -57072 33672 -57012
rect 32084 -57182 32144 -57122
rect 27892 -58104 27952 -58044
rect 29028 -58104 29088 -58044
rect 29540 -58212 29600 -58152
rect 35292 -56860 35352 -56800
rect 35138 -56966 35198 -56906
rect 34644 -57072 34704 -57012
rect 34122 -57182 34182 -57122
rect 30554 -58212 30614 -58152
rect 31576 -58212 31636 -58152
rect 35656 -57072 35716 -57012
rect 37170 -56860 37230 -56800
rect 37174 -56966 37234 -56906
rect 36664 -57072 36724 -57012
rect 36160 -57182 36220 -57122
rect 33098 -58104 33158 -58044
rect 32590 -58212 32650 -58152
rect 33616 -58212 33676 -58152
rect 37682 -57072 37742 -57012
rect 39208 -56860 39268 -56800
rect 39210 -56966 39270 -56906
rect 38708 -57072 38768 -57012
rect 38196 -57182 38256 -57122
rect 34628 -58212 34688 -58152
rect 35664 -58212 35724 -58152
rect 39710 -57072 39770 -57012
rect 42406 -55964 42466 -55904
rect 47354 -54714 47414 -54654
rect 43282 -55860 43342 -55800
rect 44300 -55632 44360 -55572
rect 44302 -55860 44362 -55800
rect 41078 -56860 41138 -56800
rect 40730 -57072 40790 -57012
rect 41244 -56966 41304 -56906
rect 40232 -57182 40292 -57122
rect 36670 -58212 36730 -58152
rect 37684 -58212 37744 -58152
rect 41750 -57072 41810 -57012
rect 45316 -55860 45376 -55800
rect 45316 -55964 45376 -55904
rect 46332 -55632 46392 -55572
rect 48606 -50696 48666 -50636
rect 48844 -50918 48904 -50858
rect 48722 -51020 48782 -50960
rect 48606 -52254 48666 -52194
rect 48602 -53156 48662 -53096
rect 48722 -54382 48782 -54322
rect 48602 -54480 48662 -54420
rect 48478 -55632 48538 -55572
rect 46852 -55742 46912 -55682
rect 47860 -55742 47920 -55682
rect 48970 -52152 49030 -52092
rect 48972 -54586 49032 -54526
rect 48844 -54714 48904 -54654
rect 49206 -48564 49266 -48504
rect 49094 -55742 49154 -55682
rect 46338 -55860 46398 -55800
rect 43284 -56966 43344 -56906
rect 42776 -57072 42836 -57012
rect 43794 -57072 43854 -57012
rect 42264 -57182 42324 -57122
rect 38700 -58212 38760 -58152
rect 39708 -58212 39768 -58152
rect 45314 -56966 45374 -56906
rect 44808 -57072 44868 -57012
rect 44296 -57182 44356 -57122
rect 40724 -58212 40784 -58152
rect 41748 -58212 41808 -58152
rect 45822 -57072 45882 -57012
rect 48498 -55964 48558 -55904
rect 47354 -56860 47414 -56800
rect 47354 -56966 47414 -56906
rect 46844 -57072 46904 -57012
rect 46336 -57182 46396 -57122
rect 43278 -58104 43338 -58044
rect 42770 -58212 42830 -58152
rect 43792 -58212 43852 -58152
rect 44810 -58212 44870 -58152
rect 45824 -58212 45884 -58152
rect 49206 -56966 49266 -56906
rect 48498 -58104 48558 -58044
rect 46848 -58212 46908 -58152
rect 17372 -58608 49372 -58454
rect 13228 -59094 13828 -58794
rect 49660 -59094 50260 -58794
rect -27578 -64832 -26978 -64532
rect -26066 -64832 -25466 -64532
rect -27388 -65100 -25564 -65036
rect -26834 -65274 -26774 -65214
rect -26316 -65274 -26256 -65214
rect -27496 -65506 -27436 -65446
rect -27496 -66100 -27436 -66040
rect -26578 -65386 -26518 -65326
rect -26706 -65506 -26646 -65446
rect -26450 -65506 -26390 -65446
rect -26962 -66230 -26902 -66170
rect -27092 -66344 -27032 -66284
rect -25648 -65386 -25588 -65326
rect -26704 -66230 -26644 -66170
rect -26446 -66230 -26386 -66170
rect -26574 -66344 -26514 -66284
rect -27246 -67080 -27186 -67020
rect -26188 -66230 -26128 -66170
rect -26058 -66344 -25998 -66284
rect -26962 -67080 -26902 -67020
rect -27094 -67192 -27034 -67132
rect -26186 -67080 -26126 -67020
rect -26058 -67192 -25998 -67132
rect -26578 -67340 -26518 -67280
rect -26320 -67300 -26260 -67240
rect -25648 -67192 -25588 -67132
rect -23578 -64832 -22978 -64532
rect -22066 -64832 -21466 -64532
rect -23388 -65100 -21564 -65036
rect -22834 -65274 -22774 -65214
rect -22316 -65274 -22256 -65214
rect -23496 -65506 -23436 -65446
rect -23496 -66100 -23436 -66040
rect -22578 -65386 -22518 -65326
rect -22706 -65506 -22646 -65446
rect -22450 -65506 -22390 -65446
rect -22962 -66230 -22902 -66170
rect -23092 -66344 -23032 -66284
rect -21648 -65386 -21588 -65326
rect -22704 -66230 -22644 -66170
rect -22446 -66230 -22386 -66170
rect -22574 -66344 -22514 -66284
rect -23246 -67080 -23186 -67020
rect -22188 -66230 -22128 -66170
rect -22058 -66344 -21998 -66284
rect -22962 -67080 -22902 -67020
rect -23094 -67192 -23034 -67132
rect -22186 -67080 -22126 -67020
rect -22058 -67192 -21998 -67132
rect -22578 -67340 -22518 -67280
rect -22320 -67300 -22260 -67240
rect -21648 -67192 -21588 -67132
rect -19578 -64832 -18978 -64532
rect -18066 -64832 -17466 -64532
rect -19388 -65100 -17564 -65036
rect -18834 -65274 -18774 -65214
rect -18316 -65274 -18256 -65214
rect -19496 -65506 -19436 -65446
rect -19496 -66100 -19436 -66040
rect -18578 -65386 -18518 -65326
rect -18706 -65506 -18646 -65446
rect -18450 -65506 -18390 -65446
rect -18962 -66230 -18902 -66170
rect -19092 -66344 -19032 -66284
rect -17648 -65386 -17588 -65326
rect -18704 -66230 -18644 -66170
rect -18446 -66230 -18386 -66170
rect -18574 -66344 -18514 -66284
rect -19246 -67080 -19186 -67020
rect -18188 -66230 -18128 -66170
rect -18058 -66344 -17998 -66284
rect -18962 -67080 -18902 -67020
rect -19094 -67192 -19034 -67132
rect -18186 -67080 -18126 -67020
rect -18058 -67192 -17998 -67132
rect -18578 -67340 -18518 -67280
rect -18320 -67300 -18260 -67240
rect -17648 -67192 -17588 -67132
rect -15578 -64832 -14978 -64532
rect -14066 -64832 -13466 -64532
rect -15388 -65100 -13564 -65036
rect -14834 -65274 -14774 -65214
rect -14316 -65274 -14256 -65214
rect -15496 -65506 -15436 -65446
rect -15496 -66100 -15436 -66040
rect -14578 -65386 -14518 -65326
rect -14706 -65506 -14646 -65446
rect -14450 -65506 -14390 -65446
rect -14962 -66230 -14902 -66170
rect -15092 -66344 -15032 -66284
rect -13648 -65386 -13588 -65326
rect -14704 -66230 -14644 -66170
rect -14446 -66230 -14386 -66170
rect -14574 -66344 -14514 -66284
rect -15246 -67080 -15186 -67020
rect -14188 -66230 -14128 -66170
rect -14058 -66344 -13998 -66284
rect -14962 -67080 -14902 -67020
rect -15094 -67192 -15034 -67132
rect -14186 -67080 -14126 -67020
rect -14058 -67192 -13998 -67132
rect -14578 -67340 -14518 -67280
rect -14320 -67300 -14260 -67240
rect -13648 -67192 -13588 -67132
rect -11578 -64832 -10978 -64532
rect -10066 -64832 -9466 -64532
rect -11388 -65100 -9564 -65036
rect -10834 -65274 -10774 -65214
rect -10316 -65274 -10256 -65214
rect -11496 -65506 -11436 -65446
rect -11496 -66100 -11436 -66040
rect -10578 -65386 -10518 -65326
rect -10706 -65506 -10646 -65446
rect -10450 -65506 -10390 -65446
rect -10962 -66230 -10902 -66170
rect -11092 -66344 -11032 -66284
rect -9648 -65386 -9588 -65326
rect -10704 -66230 -10644 -66170
rect -10446 -66230 -10386 -66170
rect -10574 -66344 -10514 -66284
rect -11246 -67080 -11186 -67020
rect -10188 -66230 -10128 -66170
rect -10058 -66344 -9998 -66284
rect -10962 -67080 -10902 -67020
rect -11094 -67192 -11034 -67132
rect -10186 -67080 -10126 -67020
rect -10058 -67192 -9998 -67132
rect -10578 -67340 -10518 -67280
rect -10320 -67300 -10260 -67240
rect -9648 -67192 -9588 -67132
rect -7578 -64832 -6978 -64532
rect -6066 -64832 -5466 -64532
rect -7388 -65100 -5564 -65036
rect -6834 -65274 -6774 -65214
rect -6316 -65274 -6256 -65214
rect -7496 -65506 -7436 -65446
rect -7496 -66100 -7436 -66040
rect -6578 -65386 -6518 -65326
rect -6706 -65506 -6646 -65446
rect -6450 -65506 -6390 -65446
rect -6962 -66230 -6902 -66170
rect -7092 -66344 -7032 -66284
rect -5648 -65386 -5588 -65326
rect -6704 -66230 -6644 -66170
rect -6446 -66230 -6386 -66170
rect -6574 -66344 -6514 -66284
rect -7246 -67080 -7186 -67020
rect -6188 -66230 -6128 -66170
rect -6058 -66344 -5998 -66284
rect -6962 -67080 -6902 -67020
rect -7094 -67192 -7034 -67132
rect -6186 -67080 -6126 -67020
rect -6058 -67192 -5998 -67132
rect -6578 -67340 -6518 -67280
rect -6320 -67300 -6260 -67240
rect -5648 -67192 -5588 -67132
rect -3578 -64832 -2978 -64532
rect -2066 -64832 -1466 -64532
rect -3388 -65100 -1564 -65036
rect -2834 -65274 -2774 -65214
rect -2316 -65274 -2256 -65214
rect -3496 -65506 -3436 -65446
rect -3496 -66100 -3436 -66040
rect -2578 -65386 -2518 -65326
rect -2706 -65506 -2646 -65446
rect -2450 -65506 -2390 -65446
rect -2962 -66230 -2902 -66170
rect -3092 -66344 -3032 -66284
rect -1648 -65386 -1588 -65326
rect -2704 -66230 -2644 -66170
rect -2446 -66230 -2386 -66170
rect -2574 -66344 -2514 -66284
rect -3246 -67080 -3186 -67020
rect -2188 -66230 -2128 -66170
rect -2058 -66344 -1998 -66284
rect -2962 -67080 -2902 -67020
rect -3094 -67192 -3034 -67132
rect -2186 -67080 -2126 -67020
rect -2058 -67192 -1998 -67132
rect -2578 -67340 -2518 -67280
rect -2320 -67300 -2260 -67240
rect -1648 -67192 -1588 -67132
rect 422 -64832 1022 -64532
rect 1934 -64832 2534 -64532
rect 612 -65100 2436 -65036
rect 1166 -65274 1226 -65214
rect 1684 -65274 1744 -65214
rect 504 -65506 564 -65446
rect 504 -66100 564 -66040
rect 1422 -65386 1482 -65326
rect 1294 -65506 1354 -65446
rect 1550 -65506 1610 -65446
rect 1038 -66230 1098 -66170
rect 908 -66344 968 -66284
rect 2352 -65386 2412 -65326
rect 1296 -66230 1356 -66170
rect 1554 -66230 1614 -66170
rect 1426 -66344 1486 -66284
rect 754 -67080 814 -67020
rect 1812 -66230 1872 -66170
rect 1942 -66344 2002 -66284
rect 1038 -67080 1098 -67020
rect 906 -67192 966 -67132
rect 1814 -67080 1874 -67020
rect 1942 -67192 2002 -67132
rect 1422 -67340 1482 -67280
rect 1680 -67300 1740 -67240
rect 2352 -67192 2412 -67132
rect 4422 -64832 5022 -64532
rect 5934 -64832 6534 -64532
rect 4612 -65100 6436 -65036
rect 5166 -65274 5226 -65214
rect 5684 -65274 5744 -65214
rect 4504 -65506 4564 -65446
rect 4504 -66100 4564 -66040
rect 5422 -65386 5482 -65326
rect 5294 -65506 5354 -65446
rect 5550 -65506 5610 -65446
rect 5038 -66230 5098 -66170
rect 4908 -66344 4968 -66284
rect 6352 -65386 6412 -65326
rect 5296 -66230 5356 -66170
rect 5554 -66230 5614 -66170
rect 5426 -66344 5486 -66284
rect 4754 -67080 4814 -67020
rect 5812 -66230 5872 -66170
rect 5942 -66344 6002 -66284
rect 5038 -67080 5098 -67020
rect 4906 -67192 4966 -67132
rect 5814 -67080 5874 -67020
rect 5942 -67192 6002 -67132
rect 5422 -67340 5482 -67280
rect 5680 -67300 5740 -67240
rect 6352 -67192 6412 -67132
rect -28230 -67616 -28170 -67556
rect -27908 -67620 -27848 -67614
rect -27908 -67668 -27902 -67620
rect -27902 -67668 -27854 -67620
rect -27854 -67668 -27848 -67620
rect -27908 -67674 -27848 -67668
rect -24230 -67616 -24170 -67556
rect -23908 -67620 -23848 -67614
rect -23908 -67668 -23902 -67620
rect -23902 -67668 -23854 -67620
rect -23854 -67668 -23848 -67620
rect -23908 -67674 -23848 -67668
rect -20230 -67616 -20170 -67556
rect -19908 -67620 -19848 -67614
rect -19908 -67668 -19902 -67620
rect -19902 -67668 -19854 -67620
rect -19854 -67668 -19848 -67620
rect -19908 -67674 -19848 -67668
rect -16230 -67616 -16170 -67556
rect -15908 -67620 -15848 -67614
rect -15908 -67668 -15902 -67620
rect -15902 -67668 -15854 -67620
rect -15854 -67668 -15848 -67620
rect -15908 -67674 -15848 -67668
rect -12230 -67616 -12170 -67556
rect -11908 -67620 -11848 -67614
rect -11908 -67668 -11902 -67620
rect -11902 -67668 -11854 -67620
rect -11854 -67668 -11848 -67620
rect -11908 -67674 -11848 -67668
rect -8230 -67616 -8170 -67556
rect -7908 -67620 -7848 -67614
rect -7908 -67668 -7902 -67620
rect -7902 -67668 -7854 -67620
rect -7854 -67668 -7848 -67620
rect -7908 -67674 -7848 -67668
rect -4230 -67616 -4170 -67556
rect -3908 -67620 -3848 -67614
rect -3908 -67668 -3902 -67620
rect -3902 -67668 -3854 -67620
rect -3854 -67668 -3848 -67620
rect -3908 -67674 -3848 -67668
rect -230 -67616 -170 -67556
rect 92 -67620 152 -67614
rect 92 -67668 98 -67620
rect 98 -67668 146 -67620
rect 146 -67668 152 -67620
rect 92 -67674 152 -67668
rect 3770 -67616 3830 -67556
rect 4092 -67620 4152 -67614
rect 4092 -67668 4098 -67620
rect 4098 -67668 4146 -67620
rect 4146 -67668 4152 -67620
rect 4092 -67674 4152 -67668
rect -26578 -67980 -26518 -67920
rect -27094 -68046 -27034 -67986
rect -26840 -68090 -26780 -68030
rect -26708 -68202 -26648 -68142
rect -26320 -68090 -26260 -68030
rect -26452 -68202 -26392 -68142
rect -26966 -68898 -26906 -68838
rect -26192 -68898 -26132 -68838
rect -27100 -69012 -27040 -68952
rect -26064 -69012 -26004 -68952
rect -27430 -69222 -25722 -69154
rect -27578 -69704 -26978 -69404
rect -26066 -69704 -25466 -69404
rect -22578 -67980 -22518 -67920
rect -23094 -68046 -23034 -67986
rect -22840 -68090 -22780 -68030
rect -22708 -68202 -22648 -68142
rect -22320 -68090 -22260 -68030
rect -22452 -68202 -22392 -68142
rect -22966 -68898 -22906 -68838
rect -22192 -68898 -22132 -68838
rect -23100 -69012 -23040 -68952
rect -22064 -69012 -22004 -68952
rect -23430 -69222 -21722 -69154
rect -23578 -69704 -22978 -69404
rect -22066 -69704 -21466 -69404
rect -18578 -67980 -18518 -67920
rect -19094 -68046 -19034 -67986
rect -18840 -68090 -18780 -68030
rect -18708 -68202 -18648 -68142
rect -18320 -68090 -18260 -68030
rect -18452 -68202 -18392 -68142
rect -18966 -68898 -18906 -68838
rect -18192 -68898 -18132 -68838
rect -19100 -69012 -19040 -68952
rect -18064 -69012 -18004 -68952
rect -19430 -69222 -17722 -69154
rect -19578 -69704 -18978 -69404
rect -18066 -69704 -17466 -69404
rect -14578 -67980 -14518 -67920
rect -15094 -68046 -15034 -67986
rect -14840 -68090 -14780 -68030
rect -14708 -68202 -14648 -68142
rect -14320 -68090 -14260 -68030
rect -14452 -68202 -14392 -68142
rect -14966 -68898 -14906 -68838
rect -14192 -68898 -14132 -68838
rect -15100 -69012 -15040 -68952
rect -14064 -69012 -14004 -68952
rect -15430 -69222 -13722 -69154
rect -15578 -69704 -14978 -69404
rect -14066 -69704 -13466 -69404
rect -10578 -67980 -10518 -67920
rect -11094 -68046 -11034 -67986
rect -10840 -68090 -10780 -68030
rect -10708 -68202 -10648 -68142
rect -10320 -68090 -10260 -68030
rect -10452 -68202 -10392 -68142
rect -10966 -68898 -10906 -68838
rect -10192 -68898 -10132 -68838
rect -11100 -69012 -11040 -68952
rect -10064 -69012 -10004 -68952
rect -11430 -69222 -9722 -69154
rect -11578 -69704 -10978 -69404
rect -10066 -69704 -9466 -69404
rect -6578 -67980 -6518 -67920
rect -7094 -68046 -7034 -67986
rect -6840 -68090 -6780 -68030
rect -6708 -68202 -6648 -68142
rect -6320 -68090 -6260 -68030
rect -6452 -68202 -6392 -68142
rect -6966 -68898 -6906 -68838
rect -6192 -68898 -6132 -68838
rect -7100 -69012 -7040 -68952
rect -6064 -69012 -6004 -68952
rect -7430 -69222 -5722 -69154
rect -7578 -69704 -6978 -69404
rect -6066 -69704 -5466 -69404
rect -2578 -67980 -2518 -67920
rect -3094 -68046 -3034 -67986
rect -2840 -68090 -2780 -68030
rect -2708 -68202 -2648 -68142
rect -2320 -68090 -2260 -68030
rect -2452 -68202 -2392 -68142
rect -2966 -68898 -2906 -68838
rect -2192 -68898 -2132 -68838
rect -3100 -69012 -3040 -68952
rect -2064 -69012 -2004 -68952
rect -3430 -69222 -1722 -69154
rect -3578 -69704 -2978 -69404
rect -2066 -69704 -1466 -69404
rect 1422 -67980 1482 -67920
rect 906 -68046 966 -67986
rect 1160 -68090 1220 -68030
rect 1292 -68202 1352 -68142
rect 1680 -68090 1740 -68030
rect 1548 -68202 1608 -68142
rect 1034 -68898 1094 -68838
rect 1808 -68898 1868 -68838
rect 900 -69012 960 -68952
rect 1936 -69012 1996 -68952
rect 570 -69222 2278 -69154
rect 422 -69704 1022 -69404
rect 1934 -69704 2534 -69404
rect 5422 -67980 5482 -67920
rect 4906 -68046 4966 -67986
rect 5160 -68090 5220 -68030
rect 5292 -68202 5352 -68142
rect 5680 -68090 5740 -68030
rect 5548 -68202 5608 -68142
rect 5034 -68898 5094 -68838
rect 5808 -68898 5868 -68838
rect 4900 -69012 4960 -68952
rect 5936 -69012 5996 -68952
rect 4570 -69222 6278 -69154
rect 4422 -69704 5022 -69404
rect 5934 -69704 6534 -69404
rect -27578 -70792 -26978 -70492
rect -26066 -70792 -25466 -70492
rect -27430 -71042 -25722 -70974
rect -27100 -71244 -27040 -71184
rect -26064 -71244 -26004 -71184
rect -26966 -71358 -26906 -71298
rect -26192 -71358 -26132 -71298
rect -26708 -72054 -26648 -71994
rect -27094 -72210 -27034 -72150
rect -26840 -72166 -26780 -72106
rect -26452 -72054 -26392 -71994
rect -26320 -72166 -26260 -72106
rect -26578 -72276 -26518 -72216
rect -23578 -70792 -22978 -70492
rect -22066 -70792 -21466 -70492
rect -23430 -71042 -21722 -70974
rect -23100 -71244 -23040 -71184
rect -22064 -71244 -22004 -71184
rect -22966 -71358 -22906 -71298
rect -22192 -71358 -22132 -71298
rect -22708 -72054 -22648 -71994
rect -23094 -72210 -23034 -72150
rect -22840 -72166 -22780 -72106
rect -22452 -72054 -22392 -71994
rect -22320 -72166 -22260 -72106
rect -22578 -72276 -22518 -72216
rect -19578 -70792 -18978 -70492
rect -18066 -70792 -17466 -70492
rect -19430 -71042 -17722 -70974
rect -19100 -71244 -19040 -71184
rect -18064 -71244 -18004 -71184
rect -18966 -71358 -18906 -71298
rect -18192 -71358 -18132 -71298
rect -18708 -72054 -18648 -71994
rect -19094 -72210 -19034 -72150
rect -18840 -72166 -18780 -72106
rect -18452 -72054 -18392 -71994
rect -18320 -72166 -18260 -72106
rect -18578 -72276 -18518 -72216
rect -15578 -70792 -14978 -70492
rect -14066 -70792 -13466 -70492
rect -15430 -71042 -13722 -70974
rect -15100 -71244 -15040 -71184
rect -14064 -71244 -14004 -71184
rect -14966 -71358 -14906 -71298
rect -14192 -71358 -14132 -71298
rect -14708 -72054 -14648 -71994
rect -15094 -72210 -15034 -72150
rect -14840 -72166 -14780 -72106
rect -14452 -72054 -14392 -71994
rect -14320 -72166 -14260 -72106
rect -14578 -72276 -14518 -72216
rect -11578 -70792 -10978 -70492
rect -10066 -70792 -9466 -70492
rect -11430 -71042 -9722 -70974
rect -11100 -71244 -11040 -71184
rect -10064 -71244 -10004 -71184
rect -10966 -71358 -10906 -71298
rect -10192 -71358 -10132 -71298
rect -10708 -72054 -10648 -71994
rect -11094 -72210 -11034 -72150
rect -10840 -72166 -10780 -72106
rect -10452 -72054 -10392 -71994
rect -10320 -72166 -10260 -72106
rect -10578 -72276 -10518 -72216
rect -7578 -70792 -6978 -70492
rect -6066 -70792 -5466 -70492
rect -7430 -71042 -5722 -70974
rect -7100 -71244 -7040 -71184
rect -6064 -71244 -6004 -71184
rect -6966 -71358 -6906 -71298
rect -6192 -71358 -6132 -71298
rect -6708 -72054 -6648 -71994
rect -7094 -72210 -7034 -72150
rect -6840 -72166 -6780 -72106
rect -6452 -72054 -6392 -71994
rect -6320 -72166 -6260 -72106
rect -6578 -72276 -6518 -72216
rect -3578 -70792 -2978 -70492
rect -2066 -70792 -1466 -70492
rect -3430 -71042 -1722 -70974
rect -3100 -71244 -3040 -71184
rect -2064 -71244 -2004 -71184
rect -2966 -71358 -2906 -71298
rect -2192 -71358 -2132 -71298
rect -2708 -72054 -2648 -71994
rect -3094 -72210 -3034 -72150
rect -2840 -72166 -2780 -72106
rect -2452 -72054 -2392 -71994
rect -2578 -72276 -2518 -72216
rect -2320 -72166 -2260 -72106
rect 422 -70792 1022 -70492
rect 1934 -70792 2534 -70492
rect 570 -71042 2278 -70974
rect 900 -71244 960 -71184
rect 1936 -71244 1996 -71184
rect 1034 -71358 1094 -71298
rect 1808 -71358 1868 -71298
rect 1292 -72054 1352 -71994
rect 906 -72210 966 -72150
rect 1160 -72166 1220 -72106
rect 1548 -72054 1608 -71994
rect 1680 -72166 1740 -72106
rect 1422 -72276 1482 -72216
rect -3246 -72392 -3186 -72332
rect 4422 -70792 5022 -70492
rect 5934 -70792 6534 -70492
rect 4570 -71042 6278 -70974
rect 4900 -71244 4960 -71184
rect 5936 -71244 5996 -71184
rect 5034 -71358 5094 -71298
rect 5808 -71358 5868 -71298
rect 5292 -72054 5352 -71994
rect 4906 -72210 4966 -72150
rect 5160 -72166 5220 -72106
rect 5548 -72054 5608 -71994
rect 5680 -72166 5740 -72106
rect 5422 -72276 5482 -72216
rect -28230 -72640 -28170 -72580
rect -27908 -72528 -27848 -72522
rect -27908 -72576 -27902 -72528
rect -27902 -72576 -27854 -72528
rect -27854 -72576 -27848 -72528
rect -27908 -72582 -27848 -72576
rect -24230 -72640 -24170 -72580
rect -23908 -72528 -23848 -72522
rect -23908 -72576 -23902 -72528
rect -23902 -72576 -23854 -72528
rect -23854 -72576 -23848 -72528
rect -23908 -72582 -23848 -72576
rect -20230 -72640 -20170 -72580
rect -19908 -72528 -19848 -72522
rect -19908 -72576 -19902 -72528
rect -19902 -72576 -19854 -72528
rect -19854 -72576 -19848 -72528
rect -19908 -72582 -19848 -72576
rect -16230 -72640 -16170 -72580
rect -15908 -72528 -15848 -72522
rect -15908 -72576 -15902 -72528
rect -15902 -72576 -15854 -72528
rect -15854 -72576 -15848 -72528
rect -15908 -72582 -15848 -72576
rect -12230 -72640 -12170 -72580
rect -11908 -72528 -11848 -72522
rect -11908 -72576 -11902 -72528
rect -11902 -72576 -11854 -72528
rect -11854 -72576 -11848 -72528
rect -11908 -72582 -11848 -72576
rect -8230 -72640 -8170 -72580
rect -7908 -72528 -7848 -72522
rect -7908 -72576 -7902 -72528
rect -7902 -72576 -7854 -72528
rect -7854 -72576 -7848 -72528
rect -7908 -72582 -7848 -72576
rect -4230 -72640 -4170 -72580
rect -3908 -72528 -3848 -72522
rect -3908 -72576 -3902 -72528
rect -3902 -72576 -3854 -72528
rect -3854 -72576 -3848 -72528
rect -3908 -72582 -3848 -72576
rect -230 -72640 -170 -72580
rect 92 -72528 152 -72522
rect 92 -72576 98 -72528
rect 98 -72576 146 -72528
rect 146 -72576 152 -72528
rect 92 -72582 152 -72576
rect 3770 -72640 3830 -72580
rect 4092 -72528 4152 -72522
rect 4092 -72576 4098 -72528
rect 4098 -72576 4146 -72528
rect 4146 -72576 4152 -72528
rect 4092 -72582 4152 -72576
rect -26578 -72916 -26518 -72856
rect -27094 -73064 -27034 -73004
rect -27246 -73176 -27186 -73116
rect -27496 -74156 -27436 -74096
rect -26962 -73176 -26902 -73116
rect -26320 -72956 -26260 -72896
rect -27092 -73912 -27032 -73852
rect -26962 -74026 -26902 -73966
rect -27496 -74750 -27436 -74690
rect -26058 -73064 -25998 -73004
rect -26186 -73176 -26126 -73116
rect -25648 -73064 -25588 -73004
rect -26574 -73912 -26514 -73852
rect -26704 -74026 -26644 -73966
rect -26446 -74026 -26386 -73966
rect -27092 -74930 -27032 -74870
rect -26058 -73912 -25998 -73852
rect -26188 -74026 -26128 -73966
rect -26706 -74750 -26646 -74690
rect -26450 -74750 -26390 -74690
rect -26578 -74870 -26518 -74810
rect -26834 -74982 -26774 -74922
rect -26316 -74982 -26256 -74922
rect -25648 -74870 -25588 -74810
rect -27388 -75160 -25564 -75096
rect -27578 -75664 -26978 -75364
rect -26066 -75664 -25466 -75364
rect -22578 -72916 -22518 -72856
rect -23094 -73064 -23034 -73004
rect -23246 -73176 -23186 -73116
rect -23496 -74156 -23436 -74096
rect -22962 -73176 -22902 -73116
rect -22320 -72956 -22260 -72896
rect -23092 -73912 -23032 -73852
rect -22962 -74026 -22902 -73966
rect -23496 -74750 -23436 -74690
rect -22058 -73064 -21998 -73004
rect -22186 -73176 -22126 -73116
rect -21648 -73064 -21588 -73004
rect -22574 -73912 -22514 -73852
rect -22704 -74026 -22644 -73966
rect -22446 -74026 -22386 -73966
rect -23092 -74928 -23032 -74868
rect -22058 -73912 -21998 -73852
rect -22188 -74026 -22128 -73966
rect -22706 -74750 -22646 -74690
rect -22450 -74750 -22390 -74690
rect -22578 -74870 -22518 -74810
rect -22834 -74982 -22774 -74922
rect -22316 -74982 -22256 -74922
rect -21648 -74870 -21588 -74810
rect -23388 -75160 -21564 -75096
rect -23578 -75664 -22978 -75364
rect -22066 -75664 -21466 -75364
rect -18578 -72916 -18518 -72856
rect -19094 -73064 -19034 -73004
rect -19246 -73176 -19186 -73116
rect -19496 -74156 -19436 -74096
rect -18962 -73176 -18902 -73116
rect -18320 -72956 -18260 -72896
rect -19092 -73912 -19032 -73852
rect -18962 -74026 -18902 -73966
rect -19496 -74750 -19436 -74690
rect -18058 -73064 -17998 -73004
rect -18186 -73176 -18126 -73116
rect -17648 -73064 -17588 -73004
rect -18574 -73912 -18514 -73852
rect -18704 -74026 -18644 -73966
rect -18446 -74026 -18386 -73966
rect -19092 -74928 -19032 -74868
rect -18058 -73912 -17998 -73852
rect -18188 -74026 -18128 -73966
rect -18706 -74750 -18646 -74690
rect -18450 -74750 -18390 -74690
rect -18578 -74870 -18518 -74810
rect -18834 -74982 -18774 -74922
rect -18316 -74982 -18256 -74922
rect -17648 -74870 -17588 -74810
rect -19388 -75160 -17564 -75096
rect -19578 -75664 -18978 -75364
rect -18066 -75664 -17466 -75364
rect -14578 -72916 -14518 -72856
rect -15094 -73064 -15034 -73004
rect -15246 -73176 -15186 -73116
rect -15496 -74156 -15436 -74096
rect -14962 -73176 -14902 -73116
rect -14320 -72956 -14260 -72896
rect -15092 -73912 -15032 -73852
rect -14962 -74026 -14902 -73966
rect -15496 -74750 -15436 -74690
rect -14058 -73064 -13998 -73004
rect -14186 -73176 -14126 -73116
rect -13648 -73064 -13588 -73004
rect -14574 -73912 -14514 -73852
rect -14704 -74026 -14644 -73966
rect -14446 -74026 -14386 -73966
rect -15092 -74928 -15032 -74868
rect -14058 -73912 -13998 -73852
rect -14188 -74026 -14128 -73966
rect -14706 -74750 -14646 -74690
rect -14450 -74750 -14390 -74690
rect -14578 -74870 -14518 -74810
rect -14834 -74982 -14774 -74922
rect -14316 -74982 -14256 -74922
rect -13648 -74870 -13588 -74810
rect -15388 -75160 -13564 -75096
rect -15578 -75664 -14978 -75364
rect -14066 -75664 -13466 -75364
rect -10578 -72916 -10518 -72856
rect -11094 -73064 -11034 -73004
rect -11246 -73176 -11186 -73116
rect -11496 -74156 -11436 -74096
rect -10962 -73176 -10902 -73116
rect -10320 -72956 -10260 -72896
rect -11092 -73912 -11032 -73852
rect -10962 -74026 -10902 -73966
rect -11496 -74750 -11436 -74690
rect -10058 -73064 -9998 -73004
rect -10186 -73176 -10126 -73116
rect -9648 -73064 -9588 -73004
rect -10574 -73912 -10514 -73852
rect -10704 -74026 -10644 -73966
rect -10446 -74026 -10386 -73966
rect -11092 -74930 -11032 -74870
rect -10058 -73912 -9998 -73852
rect -10188 -74026 -10128 -73966
rect -10706 -74750 -10646 -74690
rect -10450 -74750 -10390 -74690
rect -10578 -74870 -10518 -74810
rect -10834 -74982 -10774 -74922
rect -10316 -74982 -10256 -74922
rect -9648 -74870 -9588 -74810
rect -11388 -75160 -9564 -75096
rect -11578 -75664 -10978 -75364
rect -10066 -75664 -9466 -75364
rect -6578 -72916 -6518 -72856
rect -7094 -73064 -7034 -73004
rect -7246 -73176 -7186 -73116
rect -7496 -74156 -7436 -74096
rect -6962 -73176 -6902 -73116
rect -6320 -72956 -6260 -72896
rect -7092 -73912 -7032 -73852
rect -6962 -74026 -6902 -73966
rect -7496 -74750 -7436 -74690
rect -6058 -73064 -5998 -73004
rect -6186 -73176 -6126 -73116
rect -5648 -73064 -5588 -73004
rect -6574 -73912 -6514 -73852
rect -6704 -74026 -6644 -73966
rect -6446 -74026 -6386 -73966
rect -7092 -74930 -7032 -74870
rect -6058 -73912 -5998 -73852
rect -6188 -74026 -6128 -73966
rect -6706 -74750 -6646 -74690
rect -6450 -74750 -6390 -74690
rect -6578 -74870 -6518 -74810
rect -6834 -74982 -6774 -74922
rect -6316 -74982 -6256 -74922
rect -5648 -74870 -5588 -74810
rect -7388 -75160 -5564 -75096
rect -7578 -75664 -6978 -75364
rect -6066 -75664 -5466 -75364
rect -2578 -72916 -2518 -72856
rect -3094 -73064 -3034 -73004
rect -3246 -73176 -3186 -73116
rect -3496 -74156 -3436 -74096
rect -2962 -73176 -2902 -73116
rect -2320 -72956 -2260 -72896
rect -3092 -73912 -3032 -73852
rect -2962 -74026 -2902 -73966
rect -3496 -74750 -3436 -74690
rect -2058 -73064 -1998 -73004
rect -2186 -73176 -2126 -73116
rect -1648 -73064 -1588 -73004
rect -2574 -73912 -2514 -73852
rect -2704 -74026 -2644 -73966
rect -2446 -74026 -2386 -73966
rect -3092 -74928 -3032 -74868
rect -2058 -73912 -1998 -73852
rect -2188 -74026 -2128 -73966
rect -2706 -74750 -2646 -74690
rect -2450 -74750 -2390 -74690
rect -2578 -74870 -2518 -74810
rect -2834 -74982 -2774 -74922
rect -2316 -74982 -2256 -74922
rect -1648 -74870 -1588 -74810
rect -3388 -75160 -1564 -75096
rect -3578 -75664 -2978 -75364
rect -2066 -75664 -1466 -75364
rect 1422 -72916 1482 -72856
rect 906 -73064 966 -73004
rect 754 -73176 814 -73116
rect 504 -74156 564 -74096
rect 1038 -73176 1098 -73116
rect 1680 -72956 1740 -72896
rect 908 -73912 968 -73852
rect 1038 -74026 1098 -73966
rect 504 -74750 564 -74690
rect 1942 -73064 2002 -73004
rect 1814 -73176 1874 -73116
rect 2352 -73064 2412 -73004
rect 1426 -73912 1486 -73852
rect 1296 -74026 1356 -73966
rect 1554 -74026 1614 -73966
rect 908 -74928 968 -74868
rect 1942 -73912 2002 -73852
rect 1812 -74026 1872 -73966
rect 1294 -74750 1354 -74690
rect 1550 -74750 1610 -74690
rect 1422 -74870 1482 -74810
rect 1166 -74982 1226 -74922
rect 1684 -74982 1744 -74922
rect 2352 -74870 2412 -74810
rect 612 -75160 2436 -75096
rect 422 -75664 1022 -75364
rect 1934 -75664 2534 -75364
rect 5422 -72916 5482 -72856
rect 4906 -73064 4966 -73004
rect 4754 -73176 4814 -73116
rect 4504 -74156 4564 -74096
rect 5038 -73176 5098 -73116
rect 5680 -72956 5740 -72896
rect 4908 -73912 4968 -73852
rect 5038 -74026 5098 -73966
rect 4504 -74750 4564 -74690
rect 5942 -73064 6002 -73004
rect 5814 -73176 5874 -73116
rect 6352 -73064 6412 -73004
rect 5426 -73912 5486 -73852
rect 5296 -74026 5356 -73966
rect 5554 -74026 5614 -73966
rect 4908 -74926 4968 -74866
rect 5942 -73912 6002 -73852
rect 5812 -74026 5872 -73966
rect 5294 -74750 5354 -74690
rect 5550 -74750 5610 -74690
rect 5422 -74870 5482 -74810
rect 5166 -74982 5226 -74922
rect 5684 -74982 5744 -74922
rect 6352 -74870 6412 -74810
rect 4612 -75160 6436 -75096
rect 4422 -75664 5022 -75364
rect 5934 -75664 6534 -75364
<< metal2 >>
rect 25928 -27762 26528 -27752
rect 25928 -28072 26528 -28062
rect 49560 -27762 50160 -27752
rect 49560 -28072 50160 -28062
rect 29442 -28144 46322 -28112
rect 29442 -28358 29505 -28144
rect 46290 -28358 46322 -28144
rect 29442 -28378 46322 -28358
rect 29442 -28380 33796 -28378
rect 33430 -30060 33490 -30054
rect 34512 -30060 34572 -30054
rect 35470 -30060 35530 -30054
rect 38534 -30060 38594 -30054
rect 39552 -30060 39612 -30054
rect 40576 -30060 40636 -30054
rect 41588 -30060 41648 -30054
rect 44646 -30060 44706 -30054
rect 45658 -30060 45718 -30054
rect 46676 -30060 46736 -30054
rect 33490 -30120 34512 -30060
rect 34572 -30120 35470 -30060
rect 35530 -30120 38534 -30060
rect 38594 -30120 39552 -30060
rect 39612 -30120 40576 -30060
rect 40636 -30120 41588 -30060
rect 41648 -30120 44646 -30060
rect 44706 -30120 45658 -30060
rect 45718 -30120 46676 -30060
rect 33430 -30126 33490 -30120
rect 34512 -30126 34572 -30120
rect 35470 -30126 35530 -30120
rect 38534 -30126 38594 -30120
rect 39552 -30126 39612 -30120
rect 40576 -30126 40636 -30120
rect 41588 -30126 41648 -30120
rect 44646 -30126 44706 -30120
rect 45658 -30126 45718 -30120
rect 46676 -30126 46736 -30120
rect 33956 -30306 34016 -30300
rect 35992 -30306 36052 -30300
rect 38030 -30304 38090 -30298
rect 40060 -30304 40120 -30298
rect 42102 -30302 42162 -30296
rect 43112 -30302 43172 -30296
rect 44134 -30302 44194 -30296
rect 46170 -30302 46230 -30296
rect 34016 -30366 35992 -30306
rect 36052 -30364 38030 -30306
rect 38090 -30364 40060 -30304
rect 40120 -30362 42102 -30304
rect 42162 -30362 43112 -30302
rect 43172 -30362 44134 -30302
rect 44194 -30362 46170 -30302
rect 40120 -30364 42300 -30362
rect 36052 -30366 38212 -30364
rect 33956 -30372 34016 -30366
rect 35992 -30372 36052 -30366
rect 38030 -30370 38090 -30366
rect 40060 -30370 40120 -30364
rect 42102 -30368 42162 -30364
rect 43112 -30368 43172 -30362
rect 44134 -30368 44194 -30362
rect 46170 -30368 46230 -30362
rect 31774 -31238 31834 -31232
rect 32938 -31238 32998 -31232
rect 39048 -31238 39108 -31232
rect 31834 -31298 32938 -31238
rect 32998 -31298 39048 -31238
rect 31774 -31304 31834 -31298
rect 32938 -31304 32998 -31298
rect 39048 -31304 39108 -31298
rect 41082 -31238 41142 -31232
rect 47190 -31238 47250 -31232
rect 48440 -31238 48500 -31232
rect 41142 -31298 47190 -31238
rect 47250 -31298 48440 -31238
rect 41082 -31304 41142 -31298
rect 47190 -31304 47250 -31298
rect 48440 -31304 48500 -31298
rect 34974 -31342 35034 -31336
rect 37010 -31342 37070 -31336
rect 43116 -31342 43176 -31336
rect 45150 -31342 45210 -31336
rect 35034 -31402 37010 -31342
rect 37070 -31350 37488 -31342
rect 37704 -31350 43116 -31342
rect 37070 -31396 43116 -31350
rect 37070 -31400 39504 -31396
rect 37070 -31402 38478 -31400
rect 38716 -31402 39504 -31400
rect 39720 -31402 43116 -31396
rect 43176 -31402 45150 -31342
rect 34974 -31408 35034 -31402
rect 37010 -31408 37070 -31402
rect 43116 -31408 43176 -31402
rect 45150 -31408 45210 -31402
rect 31644 -31442 31704 -31436
rect 32938 -31442 32998 -31436
rect 39044 -31442 39104 -31436
rect 41080 -31442 41140 -31436
rect 31704 -31502 32938 -31442
rect 32998 -31502 39044 -31442
rect 39104 -31502 41080 -31442
rect 31644 -31508 31704 -31502
rect 32938 -31508 32998 -31502
rect 39044 -31508 39104 -31502
rect 41080 -31508 41140 -31502
rect 41582 -31442 41642 -31436
rect 42602 -31442 42662 -31436
rect 43628 -31442 43688 -31436
rect 41642 -31502 42602 -31442
rect 42662 -31502 43628 -31442
rect 41582 -31508 41642 -31502
rect 42602 -31508 42662 -31502
rect 43628 -31508 43688 -31502
rect 44134 -31446 44194 -31440
rect 44648 -31446 44708 -31440
rect 45152 -31446 45212 -31440
rect 45658 -31446 45718 -31440
rect 44194 -31506 44648 -31446
rect 44708 -31506 45152 -31446
rect 45212 -31506 45658 -31446
rect 45718 -31506 46178 -31446
rect 46238 -31506 46244 -31446
rect 44134 -31512 44194 -31506
rect 44648 -31512 44708 -31506
rect 45152 -31512 45212 -31506
rect 45658 -31512 45718 -31506
rect 35990 -32376 36050 -32370
rect 38024 -32376 38084 -32370
rect 40062 -32376 40122 -32372
rect 35474 -32436 35480 -32376
rect 35540 -32436 35990 -32376
rect 36050 -32436 38024 -32376
rect 38084 -32378 40266 -32376
rect 42098 -32378 42158 -32372
rect 42598 -32378 42658 -32372
rect 43112 -32378 43172 -32372
rect 43636 -32378 43696 -32372
rect 44134 -32378 44194 -32372
rect 44636 -32378 44696 -32372
rect 38084 -32436 40062 -32378
rect 35990 -32442 36050 -32436
rect 38024 -32442 38084 -32436
rect 40122 -32438 42098 -32378
rect 42158 -32438 42598 -32378
rect 42658 -32438 43112 -32378
rect 43172 -32438 43636 -32378
rect 43696 -32438 44134 -32378
rect 44194 -32438 44636 -32378
rect 44696 -32380 45004 -32378
rect 45150 -32380 45210 -32374
rect 45658 -32380 45718 -32374
rect 46168 -32380 46228 -32374
rect 44696 -32438 45150 -32380
rect 40062 -32444 40122 -32438
rect 42098 -32444 42158 -32438
rect 42598 -32444 42658 -32438
rect 43112 -32444 43172 -32438
rect 43636 -32444 43696 -32438
rect 44033 -32440 44548 -32438
rect 44134 -32444 44194 -32440
rect 44636 -32444 44696 -32438
rect 44798 -32440 45150 -32438
rect 45210 -32440 45658 -32380
rect 45718 -32440 46168 -32380
rect 45150 -32446 45210 -32440
rect 45658 -32446 45718 -32440
rect 46168 -32446 46228 -32440
rect 34972 -32474 35036 -32468
rect 36848 -32474 36912 -32468
rect 35036 -32538 36848 -32474
rect 34972 -32544 35036 -32538
rect 36848 -32544 36912 -32538
rect 41082 -32476 41142 -32470
rect 47190 -32476 47250 -32470
rect 41142 -32536 47190 -32476
rect 41082 -32542 41142 -32536
rect 47190 -32542 47250 -32536
rect 36484 -32584 36544 -32578
rect 37508 -32584 37568 -32578
rect 38536 -32584 38596 -32578
rect 34462 -32592 34522 -32586
rect 35474 -32592 35534 -32586
rect 33418 -32652 33424 -32592
rect 33484 -32652 34462 -32592
rect 34522 -32652 35474 -32592
rect 36544 -32644 37508 -32584
rect 37568 -32644 38536 -32584
rect 36484 -32650 36544 -32644
rect 37508 -32650 37568 -32644
rect 38536 -32650 38596 -32644
rect 44640 -32592 44700 -32586
rect 45652 -32592 45712 -32586
rect 46654 -32592 46714 -32586
rect 34462 -32658 34522 -32652
rect 35474 -32658 35534 -32652
rect 44700 -32652 45652 -32592
rect 45712 -32652 46654 -32592
rect 44640 -32658 44700 -32652
rect 45652 -32658 45712 -32652
rect 46654 -32658 46714 -32652
rect 33954 -33514 34014 -33508
rect 35990 -33514 36050 -33508
rect 36512 -33514 36572 -33508
rect 37010 -33514 37070 -33508
rect 38024 -33514 38084 -33508
rect 38484 -33514 38544 -33508
rect 39522 -33514 39528 -33512
rect 34014 -33574 35990 -33514
rect 36050 -33574 36512 -33514
rect 36572 -33574 37010 -33514
rect 37070 -33516 38024 -33514
rect 37070 -33518 37992 -33516
rect 37070 -33574 37484 -33518
rect 33954 -33580 34014 -33574
rect 35990 -33580 36050 -33574
rect 36512 -33580 36572 -33574
rect 37010 -33580 37070 -33574
rect 37478 -33578 37484 -33574
rect 37544 -33574 37992 -33518
rect 38084 -33574 38484 -33514
rect 38544 -33572 39528 -33514
rect 39588 -33514 39594 -33512
rect 40060 -33514 40120 -33508
rect 41566 -33514 41572 -33512
rect 39588 -33572 40060 -33514
rect 38544 -33574 40060 -33572
rect 40120 -33572 41572 -33514
rect 41632 -33514 41638 -33512
rect 41632 -33516 41944 -33514
rect 42098 -33516 42158 -33510
rect 44134 -33516 44194 -33512
rect 41632 -33518 42098 -33516
rect 42158 -33518 44322 -33516
rect 46168 -33518 46228 -33512
rect 41632 -33572 42066 -33518
rect 40120 -33574 42066 -33572
rect 37544 -33578 37550 -33574
rect 37986 -33576 37992 -33574
rect 38052 -33576 38084 -33574
rect 38024 -33580 38084 -33576
rect 38484 -33580 38544 -33574
rect 40060 -33580 40120 -33574
rect 40204 -33576 41530 -33574
rect 41736 -33576 42066 -33574
rect 42158 -33522 43082 -33518
rect 43142 -33520 44134 -33518
rect 42158 -33576 42594 -33522
rect 42060 -33578 42066 -33576
rect 42126 -33578 42158 -33576
rect 42098 -33582 42158 -33578
rect 42588 -33582 42594 -33576
rect 42654 -33576 43082 -33522
rect 42654 -33582 42660 -33576
rect 43076 -33578 43082 -33576
rect 43176 -33522 44134 -33520
rect 43176 -33576 43594 -33522
rect 43110 -33580 43116 -33578
rect 43176 -33580 43182 -33576
rect 43588 -33582 43594 -33576
rect 43654 -33576 44134 -33522
rect 43654 -33582 43660 -33576
rect 44194 -33578 46168 -33518
rect 44134 -33584 44194 -33578
rect 46168 -33584 46228 -33578
rect 29636 -33624 29696 -33620
rect 34970 -33624 35034 -33618
rect 45150 -33624 45214 -33618
rect 29634 -33626 34970 -33624
rect 29634 -33686 29636 -33626
rect 29696 -33686 34970 -33626
rect 29634 -33688 34970 -33686
rect 35034 -33688 45150 -33624
rect 29636 -33692 29696 -33688
rect 34970 -33694 35034 -33688
rect 45150 -33694 45214 -33688
rect 32932 -33762 32996 -33756
rect 32996 -33766 48436 -33762
rect 32996 -33826 39042 -33766
rect 32932 -33832 32996 -33826
rect 39036 -33830 39042 -33826
rect 39106 -33826 48436 -33766
rect 48500 -33826 48506 -33762
rect 39106 -33830 39112 -33826
rect 31774 -33912 31834 -33906
rect 41078 -33908 41142 -33902
rect 31834 -33972 32756 -33912
rect 32816 -33972 41078 -33912
rect 47184 -33912 47244 -33906
rect 41142 -33972 47184 -33912
rect 31774 -33978 31834 -33972
rect 41078 -33978 41142 -33972
rect 47184 -33978 47244 -33972
rect 32872 -34018 32932 -34012
rect 33434 -34018 33494 -34012
rect 34476 -34018 34536 -34012
rect 35476 -34018 35536 -34012
rect 38638 -34018 38698 -34012
rect 39648 -34018 39708 -34012
rect 40590 -34018 40650 -34012
rect 32932 -34078 33434 -34018
rect 33494 -34078 34476 -34018
rect 34536 -34078 35476 -34018
rect 35536 -34078 38638 -34018
rect 38698 -34078 39648 -34018
rect 39708 -34078 40590 -34018
rect 32872 -34084 32932 -34078
rect 33434 -34084 33494 -34078
rect 34476 -34084 34536 -34078
rect 35476 -34084 35536 -34078
rect 38638 -34084 38698 -34078
rect 39648 -34084 39708 -34078
rect 40590 -34084 40650 -34078
rect 32986 -34220 33046 -34214
rect 36164 -34220 36224 -34214
rect 40232 -34220 40292 -34214
rect 44308 -34220 44368 -34214
rect 47504 -34220 47564 -34214
rect 33046 -34280 36164 -34220
rect 36224 -34280 40232 -34220
rect 40292 -34280 44308 -34220
rect 44368 -34280 47504 -34220
rect 32986 -34286 33046 -34280
rect 36164 -34286 36224 -34280
rect 40232 -34286 40292 -34280
rect 44308 -34286 44368 -34280
rect 47504 -34286 47564 -34280
rect 34130 -35156 34190 -35150
rect 36164 -35156 36224 -35150
rect 38206 -35156 38266 -35150
rect 40232 -35156 40292 -35150
rect 42274 -35156 42334 -35150
rect 44310 -35156 44370 -35150
rect 46346 -35156 46406 -35150
rect 34190 -35216 36164 -35156
rect 36224 -35216 38206 -35156
rect 38266 -35216 40232 -35156
rect 40292 -35216 42274 -35156
rect 42334 -35216 44310 -35156
rect 44370 -35216 46346 -35156
rect 34130 -35222 34190 -35216
rect 36164 -35222 36224 -35216
rect 38206 -35222 38266 -35216
rect 40232 -35222 40292 -35216
rect 42274 -35222 42334 -35216
rect 44310 -35222 44370 -35216
rect 46346 -35222 46406 -35216
rect 34634 -35264 34694 -35258
rect 34694 -35324 35656 -35264
rect 35716 -35324 36674 -35264
rect 36734 -35324 37698 -35264
rect 37758 -35324 38712 -35264
rect 38772 -35324 39730 -35264
rect 39790 -35324 40740 -35264
rect 40800 -35324 41762 -35264
rect 41822 -35324 42776 -35264
rect 42836 -35324 43808 -35264
rect 43868 -35324 44818 -35264
rect 44878 -35324 45840 -35264
rect 45900 -35324 45906 -35264
rect 34634 -35330 34694 -35324
rect 34126 -36188 34186 -36182
rect 38206 -36188 38266 -36182
rect 42274 -36188 42334 -36182
rect 46342 -36188 46402 -36182
rect 48734 -36188 48794 -36182
rect 26594 -36248 34126 -36188
rect 34186 -36248 38206 -36188
rect 38266 -36248 42274 -36188
rect 42334 -36248 46342 -36188
rect 46402 -36248 48734 -36188
rect -14318 -40774 -14218 -40765
rect -7399 -40852 -7309 -40848
rect -15855 -41124 -15765 -41120
rect -14318 -41124 -14218 -40874
rect -7404 -40857 -5210 -40852
rect -7404 -40947 -7399 -40857
rect -7309 -40947 -5210 -40857
rect -7404 -40952 -5210 -40947
rect -7399 -40956 -7309 -40952
rect -7973 -41094 -7883 -41090
rect -15860 -41129 -14218 -41124
rect -15860 -41219 -15855 -41129
rect -15765 -41219 -14218 -41129
rect -13177 -41194 -13168 -41094
rect -13068 -41099 -7878 -41094
rect -13068 -41189 -7973 -41099
rect -7883 -41189 -7878 -41099
rect -13068 -41194 -7878 -41189
rect -5310 -41146 -5210 -40952
rect -7973 -41198 -7883 -41194
rect -15860 -41224 -14218 -41219
rect -15855 -41228 -15765 -41224
rect -5310 -41255 -5210 -41246
rect 11452 -42356 22722 -42100
rect -14632 -42469 -14532 -42464
rect -14636 -42559 -14627 -42469
rect -14537 -42559 -14528 -42469
rect -6432 -42537 -6332 -42532
rect -14632 -47424 -14532 -42559
rect -6436 -42627 -6427 -42537
rect -6337 -42627 -6328 -42537
rect -11643 -42836 -11553 -42832
rect -9531 -42836 -9441 -42832
rect -13746 -42841 -11548 -42836
rect -13746 -42931 -11643 -42841
rect -11553 -42931 -11548 -42841
rect -13746 -42936 -11548 -42931
rect -9536 -42841 -7342 -42836
rect -9536 -42931 -9531 -42841
rect -9441 -42931 -7342 -42841
rect -9536 -42936 -7342 -42931
rect -13746 -43120 -13646 -42936
rect -11643 -42940 -11553 -42936
rect -9531 -42940 -9441 -42936
rect -13746 -43229 -13646 -43220
rect -7442 -43112 -7342 -42936
rect -7442 -43221 -7342 -43212
rect -10917 -44832 -10827 -44828
rect -10922 -44837 -10064 -44832
rect -10922 -44927 -10917 -44837
rect -10827 -44927 -10064 -44837
rect -10922 -44932 -10064 -44927
rect -10917 -44936 -10827 -44932
rect -10164 -45124 -10064 -44932
rect -10164 -45233 -10064 -45224
rect -7444 -46758 -7344 -46749
rect -13741 -46836 -13651 -46832
rect -13746 -46841 -11544 -46836
rect -13746 -46931 -13741 -46841
rect -13651 -46931 -11544 -46841
rect -13746 -46936 -11544 -46931
rect -13741 -46940 -13651 -46936
rect -11644 -47134 -11544 -46936
rect -9537 -47104 -9447 -47100
rect -7444 -47104 -7344 -46858
rect -9542 -47109 -7344 -47104
rect -9542 -47199 -9537 -47109
rect -9447 -47199 -7344 -47109
rect -9542 -47204 -7344 -47199
rect -9537 -47208 -9447 -47204
rect -11644 -47243 -11544 -47234
rect -14632 -47533 -14532 -47524
rect -6432 -47530 -6332 -42627
rect 11452 -42648 11814 -42356
rect 22578 -42648 22722 -42356
rect 11452 -42956 22722 -42648
rect 11452 -43278 23804 -42956
rect 26594 -43600 26654 -36248
rect 34126 -36254 34186 -36248
rect 38206 -36254 38266 -36248
rect 42274 -36254 42334 -36248
rect 46342 -36254 46402 -36248
rect 48734 -36254 48794 -36248
rect 32130 -36320 32190 -36314
rect 36672 -36320 36678 -36318
rect 32190 -36322 36678 -36320
rect 32190 -36380 34632 -36322
rect 32130 -36386 32190 -36380
rect 34626 -36382 34632 -36380
rect 34692 -36326 36678 -36322
rect 34692 -36380 35646 -36326
rect 34692 -36382 34698 -36380
rect 35640 -36386 35646 -36380
rect 35706 -36378 36678 -36326
rect 36738 -36320 36744 -36318
rect 37670 -36320 37676 -36318
rect 36738 -36378 37676 -36320
rect 37736 -36320 37742 -36318
rect 38714 -36320 38720 -36318
rect 37736 -36378 38720 -36320
rect 38780 -36320 38786 -36318
rect 42770 -36320 42776 -36318
rect 38780 -36322 42776 -36320
rect 38780 -36378 39724 -36322
rect 35706 -36380 39724 -36378
rect 35706 -36386 35712 -36380
rect 39718 -36382 39724 -36380
rect 39784 -36380 40740 -36322
rect 39784 -36382 39790 -36380
rect 40734 -36382 40740 -36380
rect 40800 -36380 41744 -36322
rect 40800 -36382 40806 -36380
rect 41738 -36382 41744 -36380
rect 41804 -36378 42776 -36322
rect 42836 -36320 42842 -36318
rect 48298 -36320 48358 -36314
rect 42836 -36322 48298 -36320
rect 42836 -36378 43792 -36322
rect 41804 -36380 43792 -36378
rect 41804 -36382 41810 -36380
rect 43786 -36382 43792 -36380
rect 43852 -36380 44820 -36322
rect 43852 -36382 43858 -36380
rect 44814 -36382 44820 -36380
rect 44880 -36380 45840 -36322
rect 44880 -36382 44886 -36380
rect 45834 -36382 45840 -36380
rect 45900 -36380 48298 -36322
rect 45900 -36382 45906 -36380
rect 48298 -36386 48358 -36380
rect 39524 -36530 39584 -36524
rect 39584 -36590 41260 -36530
rect 41320 -36590 41326 -36530
rect 47158 -36544 47218 -36540
rect 47156 -36546 48500 -36544
rect 39524 -36596 39584 -36590
rect 47156 -36606 47158 -36546
rect 47218 -36548 48500 -36546
rect 47218 -36606 48440 -36548
rect 47156 -36608 48440 -36606
rect 48500 -36608 48506 -36548
rect 47158 -36612 47218 -36608
rect 40540 -36726 40604 -36720
rect 44604 -36726 44668 -36720
rect 45628 -36726 45692 -36720
rect 46640 -36726 46704 -36720
rect 40604 -36790 44604 -36726
rect 44668 -36790 45628 -36726
rect 45692 -36790 46640 -36726
rect 40540 -36796 40604 -36790
rect 44604 -36796 44668 -36790
rect 45628 -36796 45692 -36790
rect 46640 -36796 46704 -36790
rect 32756 -36848 32816 -36842
rect 33922 -36848 33982 -36842
rect 35958 -36848 36018 -36842
rect 32816 -36908 33922 -36848
rect 33982 -36908 35958 -36848
rect 32756 -36914 32816 -36908
rect 33922 -36914 33982 -36908
rect 35958 -36914 36018 -36908
rect 36466 -36848 36530 -36842
rect 40542 -36848 40606 -36842
rect 36530 -36912 40542 -36848
rect 36466 -36918 36530 -36912
rect 40542 -36918 40606 -36912
rect 44104 -36848 44164 -36842
rect 46138 -36848 46198 -36842
rect 48582 -36848 48642 -36842
rect 44164 -36908 46138 -36848
rect 46198 -36908 48582 -36848
rect 44104 -36914 44164 -36908
rect 46138 -36914 46198 -36908
rect 48582 -36914 48642 -36908
rect 32004 -36930 32064 -36924
rect 32246 -36930 32306 -36924
rect 32064 -36990 32246 -36930
rect 32004 -36996 32064 -36990
rect 32246 -36996 32306 -36990
rect 34940 -37796 35000 -37790
rect 36976 -37796 37036 -37790
rect 35000 -37856 36976 -37796
rect 34940 -37862 35000 -37856
rect 36976 -37862 37036 -37856
rect 37318 -37794 37378 -37788
rect 40032 -37794 40092 -37788
rect 37378 -37854 40032 -37794
rect 37318 -37860 37378 -37854
rect 40032 -37860 40092 -37854
rect 45120 -37796 45180 -37790
rect 47156 -37796 47216 -37790
rect 45180 -37856 47156 -37796
rect 45120 -37862 45180 -37856
rect 29120 -37884 29180 -37878
rect 30142 -37884 30202 -37878
rect 29180 -37944 30142 -37884
rect 29120 -37950 29180 -37944
rect 30142 -37950 30202 -37944
rect 32488 -37894 32548 -37888
rect 45228 -37894 45288 -37856
rect 47156 -37862 47216 -37856
rect 32548 -37954 45288 -37894
rect 32488 -37960 32548 -37954
rect 29228 -37996 29288 -37990
rect 30012 -37996 30072 -37990
rect 29288 -38056 30012 -37996
rect 29228 -38062 29288 -38056
rect 30012 -38062 30072 -38056
rect 32624 -37992 32684 -37986
rect 34940 -37992 35000 -37986
rect 32684 -38052 34940 -37992
rect 32624 -38058 32684 -38052
rect 34940 -38058 35000 -38052
rect 35960 -37990 36020 -37984
rect 41050 -37990 41110 -37984
rect 48422 -37990 48482 -37984
rect 36020 -38050 41050 -37990
rect 41110 -38050 48422 -37990
rect 35960 -38056 36020 -38050
rect 41050 -38056 41110 -38050
rect 48422 -38056 48482 -38050
rect 33926 -38102 33986 -38096
rect 35960 -38102 36020 -38096
rect 33986 -38162 35960 -38102
rect 33926 -38168 33986 -38162
rect 35960 -38168 36020 -38162
rect 39016 -38104 39076 -38098
rect 41050 -38104 41110 -38098
rect 39076 -38164 41050 -38104
rect 39016 -38170 39076 -38164
rect 41050 -38170 41110 -38164
rect 44106 -38104 44166 -38098
rect 46140 -38102 46200 -38098
rect 46072 -38104 46200 -38102
rect 48734 -38104 48794 -38098
rect 44166 -38164 46140 -38104
rect 46200 -38164 48734 -38104
rect 44106 -38170 44166 -38164
rect 46072 -38166 46200 -38164
rect 46140 -38170 46200 -38166
rect 48734 -38170 48794 -38164
rect 27458 -38918 27518 -38912
rect 30652 -38918 30712 -38912
rect 27518 -38978 30652 -38918
rect 27458 -38984 27518 -38978
rect 30652 -38984 30712 -38978
rect 28618 -39028 28678 -39022
rect 31804 -39028 31864 -39022
rect 28678 -39088 31804 -39028
rect 44970 -39038 45030 -39032
rect 28618 -39094 28678 -39088
rect 31804 -39094 31864 -39088
rect 32246 -39052 32306 -39046
rect 39012 -39052 39072 -39046
rect 40032 -39052 40092 -39046
rect 42068 -39052 42128 -39046
rect 32306 -39112 39012 -39052
rect 39072 -39112 40032 -39052
rect 40092 -39112 42068 -39052
rect 45030 -39098 49392 -39038
rect 44970 -39104 45030 -39098
rect 32246 -39118 32306 -39112
rect 39012 -39118 39072 -39112
rect 40032 -39118 40092 -39112
rect 42068 -39118 42128 -39112
rect 45118 -39148 45178 -39142
rect 47158 -39148 47218 -39142
rect 48298 -39148 48358 -39142
rect 31996 -39156 32056 -39150
rect 36978 -39156 37038 -39150
rect 44102 -39156 44162 -39150
rect 32056 -39216 34942 -39156
rect 35002 -39216 36978 -39156
rect 37038 -39216 44102 -39156
rect 45178 -39208 47158 -39148
rect 47218 -39208 48298 -39148
rect 45118 -39214 45178 -39208
rect 47158 -39214 47218 -39208
rect 48298 -39214 48358 -39208
rect 31996 -39222 32056 -39216
rect 36978 -39222 37038 -39216
rect 44102 -39222 44162 -39216
rect 36976 -39258 37036 -39252
rect 46138 -39258 46198 -39252
rect 32242 -39266 32302 -39260
rect 32908 -39266 32968 -39260
rect 32302 -39326 32908 -39266
rect 37036 -39318 46138 -39258
rect 36976 -39324 37036 -39318
rect 46138 -39324 46198 -39318
rect 32242 -39332 32302 -39326
rect 32908 -39332 32968 -39326
rect 34942 -39360 35002 -39354
rect 36976 -39360 37036 -39354
rect 35002 -39420 36976 -39360
rect 34942 -39426 35002 -39420
rect 36976 -39426 37036 -39420
rect 40032 -39358 40092 -39352
rect 41050 -39358 41110 -39352
rect 42066 -39358 42126 -39352
rect 44970 -39358 45030 -39352
rect 40092 -39418 41050 -39358
rect 41110 -39418 42066 -39358
rect 42126 -39418 44970 -39358
rect 40032 -39424 40092 -39418
rect 41050 -39424 41110 -39418
rect 42066 -39424 42126 -39418
rect 44970 -39424 45030 -39418
rect 45122 -39356 45182 -39350
rect 47156 -39356 47216 -39350
rect 48422 -39356 48482 -39350
rect 45182 -39416 47156 -39356
rect 47216 -39416 48422 -39356
rect 48482 -39416 49264 -39356
rect 45122 -39422 45182 -39416
rect 47156 -39422 47216 -39416
rect 48422 -39422 48482 -39416
rect 29134 -39952 29194 -39946
rect 30144 -39952 30204 -39946
rect 27326 -40066 27332 -40006
rect 27392 -40066 27398 -40006
rect 29194 -40012 30144 -39952
rect 29134 -40018 29194 -40012
rect 30144 -40018 30204 -40012
rect 29240 -40052 29300 -40046
rect 30026 -40052 30086 -40046
rect 26840 -41122 26846 -41062
rect 26906 -41122 26912 -41062
rect 26720 -41622 26726 -41562
rect 26786 -41622 26792 -41562
rect 26726 -43472 26786 -41622
rect 26726 -43538 26786 -43532
rect 26846 -43470 26906 -41122
rect 26980 -41298 26986 -41238
rect 27046 -41298 27052 -41238
rect 26986 -42942 27046 -41298
rect 27208 -42120 27214 -42060
rect 27274 -42120 27280 -42060
rect 26986 -43452 27046 -43002
rect 27214 -43436 27274 -42120
rect 27332 -43336 27392 -40066
rect 29300 -40112 30026 -40052
rect 29240 -40118 29300 -40112
rect 30026 -40118 30086 -40112
rect 36978 -40300 37038 -40294
rect 38780 -40300 38840 -40294
rect 32130 -40308 32190 -40302
rect 33924 -40308 33984 -40302
rect 35960 -40308 36020 -40302
rect 32190 -40368 33924 -40308
rect 33984 -40368 35960 -40308
rect 37038 -40360 38780 -40300
rect 36978 -40366 37038 -40360
rect 38780 -40366 38840 -40360
rect 39014 -40306 39074 -40300
rect 41050 -40306 41110 -40300
rect 39074 -40366 41050 -40306
rect 32130 -40374 32190 -40368
rect 30126 -41300 30132 -41240
rect 30192 -41300 30198 -41240
rect 27880 -41472 27886 -41412
rect 27946 -41472 27952 -41412
rect 27774 -41884 27780 -41824
rect 27840 -41884 27846 -41824
rect 27654 -42002 27660 -41942
rect 27720 -42002 27726 -41942
rect 27660 -43326 27720 -42002
rect 27780 -42918 27840 -41884
rect 27763 -42927 27853 -42918
rect 27763 -43026 27853 -43017
rect 27326 -43396 27332 -43336
rect 27392 -43396 27398 -43336
rect 27780 -43334 27840 -43026
rect 27660 -43392 27720 -43386
rect 27774 -43394 27780 -43334
rect 27840 -43394 27846 -43334
rect 27886 -43470 27946 -41472
rect 30132 -41822 30192 -41300
rect 30126 -41882 30132 -41822
rect 30192 -41882 30198 -41822
rect 27214 -43502 27274 -43496
rect 26986 -43518 27046 -43512
rect 27880 -43530 27886 -43470
rect 27946 -43530 27952 -43470
rect 26846 -43536 26906 -43530
rect 27104 -43590 27164 -43584
rect 32358 -43590 32418 -40368
rect 33924 -40374 33984 -40368
rect 35960 -40374 36020 -40368
rect 39014 -40372 39074 -40366
rect 41050 -40372 41110 -40366
rect 44104 -40304 44164 -40298
rect 46140 -40304 46200 -40298
rect 44164 -40364 46140 -40304
rect 44104 -40370 44164 -40364
rect 46140 -40370 46200 -40364
rect 35960 -40416 36020 -40410
rect 41048 -40416 41108 -40410
rect 48298 -40416 48358 -40410
rect 36020 -40476 41048 -40416
rect 41108 -40476 48298 -40416
rect 35960 -40482 36020 -40476
rect 41048 -40482 41108 -40476
rect 48298 -40482 48358 -40476
rect 32756 -40516 32816 -40510
rect 32816 -40576 45340 -40516
rect 32756 -40582 32816 -40576
rect 34938 -40618 34998 -40612
rect 36972 -40618 37032 -40612
rect 34998 -40678 36972 -40618
rect 45126 -40618 45186 -40612
rect 45280 -40618 45340 -40576
rect 47160 -40618 47220 -40612
rect 34938 -40684 34998 -40678
rect 36972 -40684 37032 -40678
rect 37176 -40630 37236 -40624
rect 37236 -40690 40538 -40630
rect 40598 -40690 41554 -40630
rect 41614 -40690 44614 -40630
rect 44674 -40690 44680 -40630
rect 45186 -40678 47160 -40618
rect 45126 -40684 45186 -40678
rect 47160 -40684 47220 -40678
rect 37176 -40696 37236 -40690
rect 49204 -41091 49264 -39416
rect 49182 -41181 49191 -41091
rect 49281 -41181 49290 -41091
rect 32488 -41566 32548 -41560
rect 33920 -41566 33980 -41560
rect 35956 -41566 36016 -41560
rect 32548 -41626 33920 -41566
rect 33980 -41626 35956 -41566
rect 32488 -41632 32548 -41626
rect 33920 -41632 33980 -41626
rect 35956 -41632 36016 -41626
rect 44108 -41566 44168 -41560
rect 46144 -41566 46204 -41560
rect 44168 -41626 46144 -41566
rect 44108 -41632 44168 -41626
rect 32624 -41696 32684 -41690
rect 44238 -41696 44298 -41626
rect 46144 -41632 46204 -41626
rect 32684 -41756 44298 -41696
rect 32624 -41762 32684 -41756
rect 36978 -41836 37038 -41830
rect 48582 -41836 48642 -41830
rect 37038 -41896 48582 -41836
rect 36978 -41902 37038 -41896
rect 27164 -43650 32418 -43590
rect 27104 -43656 27164 -43650
rect 26594 -43666 26654 -43660
rect 38698 -43820 38758 -41896
rect 38698 -43886 38758 -43880
rect 43802 -43820 43862 -41896
rect 47862 -43826 47922 -41896
rect 48582 -41902 48642 -41896
rect 43802 -43886 43862 -43880
rect 47856 -43886 47862 -43826
rect 47922 -43886 47928 -43826
rect 23882 -44198 23942 -44192
rect 27660 -44198 27720 -44192
rect 23942 -44258 27660 -44198
rect 23882 -44264 23942 -44258
rect 27660 -44264 27720 -44258
rect 25408 -44332 25468 -44326
rect 27214 -44332 27274 -44326
rect 25468 -44392 27214 -44332
rect 25408 -44398 25468 -44392
rect 27214 -44398 27274 -44392
rect 26986 -45104 27046 -45098
rect 27780 -45104 27840 -45098
rect 27046 -45164 27780 -45104
rect 26986 -45170 27046 -45164
rect 27780 -45170 27840 -45164
rect 27456 -45556 27516 -45550
rect 27516 -45616 29030 -45556
rect 29090 -45616 29096 -45556
rect 27456 -45622 27516 -45616
rect 30044 -45772 30104 -45766
rect 32084 -45772 32144 -45766
rect 34124 -45772 34184 -45766
rect 36154 -45772 36214 -45766
rect 38194 -45772 38254 -45766
rect 40226 -45772 40286 -45766
rect 42266 -45772 42326 -45766
rect 44302 -45772 44362 -45766
rect 46336 -45772 46396 -45766
rect 30104 -45832 32084 -45772
rect 32144 -45832 34124 -45772
rect 34184 -45832 36154 -45772
rect 36214 -45832 38194 -45772
rect 38254 -45832 40226 -45772
rect 40286 -45832 42266 -45772
rect 42326 -45832 44302 -45772
rect 44362 -45832 46336 -45772
rect 30044 -45838 30104 -45832
rect 32084 -45838 32144 -45832
rect 34124 -45838 34184 -45832
rect 36154 -45838 36214 -45832
rect 38194 -45838 38254 -45832
rect 40226 -45838 40286 -45832
rect 42266 -45838 42326 -45832
rect 44302 -45838 44362 -45832
rect 46336 -45838 46396 -45832
rect 27668 -45892 27728 -45886
rect 28012 -45892 28072 -45886
rect 27728 -45952 28012 -45892
rect 27668 -45958 27728 -45952
rect 28012 -45958 28072 -45952
rect 29536 -45898 29596 -45892
rect 37680 -45898 37740 -45892
rect 29596 -45958 30550 -45898
rect 30610 -45958 31572 -45898
rect 31632 -45958 32586 -45898
rect 32646 -45958 33612 -45898
rect 33672 -45958 34624 -45898
rect 34684 -45958 35660 -45898
rect 35720 -45958 36666 -45898
rect 36726 -45958 37680 -45898
rect 37740 -45958 38696 -45898
rect 38756 -45958 39704 -45898
rect 39764 -45958 40720 -45898
rect 40780 -45958 41744 -45898
rect 41804 -45958 42766 -45898
rect 42826 -45958 43788 -45898
rect 43848 -45958 44806 -45898
rect 44866 -45958 45820 -45898
rect 45880 -45958 46844 -45898
rect 46904 -45958 46910 -45898
rect 29536 -45964 29596 -45958
rect 37680 -45964 37740 -45958
rect 27886 -46014 27946 -46008
rect 33100 -46014 33160 -46008
rect 43288 -46014 43348 -46008
rect 47360 -46014 47420 -46008
rect 48492 -46014 48552 -46008
rect 27946 -46074 33100 -46014
rect 33160 -46074 43288 -46014
rect 43348 -46074 47360 -46014
rect 47420 -46074 48492 -46014
rect 27886 -46080 27946 -46074
rect 33100 -46080 33160 -46074
rect 43288 -46080 43348 -46074
rect 47360 -46080 47420 -46074
rect 48492 -46080 48552 -46074
rect 26986 -46860 27046 -46854
rect 27780 -46860 27840 -46854
rect 27046 -46920 27780 -46860
rect 26986 -46926 27046 -46920
rect 27780 -46926 27840 -46920
rect 30048 -46936 30108 -46930
rect 32088 -46936 32148 -46930
rect 34120 -46936 34180 -46930
rect 36152 -46936 36212 -46930
rect 38188 -46936 38248 -46930
rect 40224 -46936 40284 -46930
rect 42262 -46936 42322 -46930
rect 44300 -46936 44360 -46930
rect 46336 -46936 46396 -46930
rect 30108 -46996 32088 -46936
rect 32148 -46996 34120 -46936
rect 34180 -46996 36152 -46936
rect 36212 -46996 38188 -46936
rect 38248 -46996 40224 -46936
rect 40284 -46996 42262 -46936
rect 42322 -46996 44300 -46936
rect 44360 -46996 46336 -46936
rect 30048 -47002 30108 -46996
rect 32088 -47002 32148 -46996
rect 34120 -47002 34180 -46996
rect 36152 -47002 36212 -46996
rect 38188 -47002 38248 -46996
rect 40224 -47002 40284 -46996
rect 42262 -47002 42322 -46996
rect 44300 -47002 44360 -46996
rect 46336 -47002 46396 -46996
rect 29540 -47046 29600 -47040
rect 30562 -47046 30622 -47040
rect 31576 -47046 31636 -47040
rect 32590 -47046 32650 -47040
rect 33608 -47046 33668 -47040
rect 34634 -47046 34694 -47040
rect 35654 -47046 35714 -47040
rect 36674 -47046 36734 -47040
rect 37676 -47046 37736 -47040
rect 38702 -47046 38762 -47040
rect 39720 -47046 39780 -47040
rect 40728 -47046 40788 -47040
rect 41740 -47046 41800 -47040
rect 42772 -47046 42832 -47040
rect 43786 -47046 43846 -47040
rect 44804 -47046 44864 -47040
rect 45828 -47046 45888 -47040
rect 46848 -47046 46908 -47040
rect 29600 -47106 30562 -47046
rect 30622 -47106 31576 -47046
rect 31636 -47106 32590 -47046
rect 32650 -47106 33608 -47046
rect 33668 -47106 34634 -47046
rect 34694 -47106 35654 -47046
rect 35714 -47106 36674 -47046
rect 36734 -47106 37676 -47046
rect 37736 -47106 38702 -47046
rect 38762 -47106 39720 -47046
rect 39780 -47106 40728 -47046
rect 40788 -47106 41740 -47046
rect 41800 -47106 42772 -47046
rect 42832 -47106 43786 -47046
rect 43846 -47106 44804 -47046
rect 44864 -47106 45828 -47046
rect 45888 -47106 46848 -47046
rect 29540 -47112 29600 -47106
rect 30562 -47112 30622 -47106
rect 31576 -47112 31636 -47106
rect 32590 -47112 32650 -47106
rect 33608 -47112 33668 -47106
rect 34634 -47112 34694 -47106
rect 35654 -47112 35714 -47106
rect 36674 -47112 36734 -47106
rect 37676 -47112 37736 -47106
rect 38702 -47112 38762 -47106
rect 39720 -47112 39780 -47106
rect 40728 -47112 40788 -47106
rect 41740 -47112 41800 -47106
rect 42772 -47112 42832 -47106
rect 43786 -47112 43846 -47106
rect 44804 -47112 44864 -47106
rect 45828 -47112 45888 -47106
rect 46848 -47112 46908 -47106
rect 27564 -47152 27624 -47146
rect 29030 -47152 29090 -47146
rect 31070 -47152 31130 -47146
rect 33100 -47152 33160 -47146
rect 35140 -47152 35200 -47146
rect 37174 -47152 37234 -47146
rect 39210 -47152 39270 -47146
rect 41246 -47152 41306 -47146
rect 43286 -47152 43346 -47146
rect 45316 -47152 45376 -47146
rect 47356 -47152 47416 -47146
rect 27624 -47212 29030 -47152
rect 29090 -47212 31070 -47152
rect 31130 -47212 33100 -47152
rect 33160 -47212 35140 -47152
rect 35200 -47212 37174 -47152
rect 37234 -47212 39210 -47152
rect 39270 -47212 41246 -47152
rect 41306 -47212 43286 -47152
rect 43346 -47212 45316 -47152
rect 45376 -47212 47356 -47152
rect 27564 -47218 27624 -47212
rect 29030 -47218 29090 -47212
rect 31070 -47218 31130 -47212
rect 33100 -47218 33160 -47212
rect 35140 -47218 35200 -47212
rect 37174 -47218 37234 -47212
rect 39210 -47218 39270 -47212
rect 41246 -47218 41306 -47212
rect 43286 -47218 43346 -47212
rect 45316 -47218 45376 -47212
rect 47356 -47218 47416 -47212
rect 28016 -47258 28076 -47252
rect 28514 -47258 28574 -47252
rect 29026 -47258 29086 -47252
rect 35306 -47258 35366 -47252
rect 37174 -47258 37234 -47252
rect 39212 -47258 39272 -47252
rect 41092 -47258 41152 -47252
rect 27324 -47318 27330 -47258
rect 27390 -47318 28016 -47258
rect 28076 -47318 28514 -47258
rect 28574 -47318 29026 -47258
rect 29086 -47318 35306 -47258
rect 35366 -47318 37174 -47258
rect 37234 -47318 39212 -47258
rect 39272 -47318 41092 -47258
rect 28016 -47324 28076 -47318
rect 28514 -47324 28574 -47318
rect 29026 -47324 29086 -47318
rect 35306 -47324 35366 -47318
rect 37174 -47324 37234 -47318
rect 39212 -47324 39272 -47318
rect 41092 -47324 41152 -47318
rect 45316 -47256 45376 -47250
rect 48492 -47256 48552 -47250
rect 45376 -47316 48492 -47256
rect 45316 -47322 45376 -47316
rect 48492 -47322 48552 -47316
rect -6432 -47639 -6332 -47630
rect 27886 -48148 27946 -48142
rect 31064 -48148 31124 -48142
rect 34120 -48148 34180 -48142
rect 40226 -48148 40286 -48142
rect 45320 -48148 45380 -48142
rect 27946 -48208 31064 -48148
rect 31124 -48208 34120 -48148
rect 34180 -48208 40226 -48148
rect 40286 -48208 45320 -48148
rect 27886 -48214 27946 -48208
rect 31064 -48214 31124 -48208
rect 34120 -48214 34180 -48208
rect 40226 -48214 40286 -48208
rect 45320 -48214 45380 -48208
rect 27456 -48252 27516 -48246
rect 28010 -48252 28070 -48246
rect 29530 -48252 29590 -48246
rect 27516 -48312 28010 -48252
rect 28070 -48312 29530 -48252
rect 27456 -48318 27516 -48312
rect 28010 -48318 28070 -48312
rect 29530 -48318 29590 -48312
rect 30042 -48252 30102 -48246
rect 31066 -48252 31126 -48246
rect 32078 -48252 32138 -48246
rect 33098 -48252 33158 -48246
rect 36156 -48252 36216 -48246
rect 38194 -48252 38254 -48246
rect 41244 -48252 41304 -48246
rect 42262 -48252 42322 -48246
rect 43282 -48252 43342 -48246
rect 44298 -48252 44358 -48246
rect 46334 -48252 46394 -48246
rect 30102 -48312 31066 -48252
rect 31126 -48312 32078 -48252
rect 32138 -48312 33098 -48252
rect 33158 -48312 36156 -48252
rect 36216 -48312 38194 -48252
rect 38254 -48312 41244 -48252
rect 41304 -48312 42262 -48252
rect 42322 -48312 43282 -48252
rect 43342 -48312 44298 -48252
rect 44358 -48312 46334 -48252
rect 30042 -48318 30102 -48312
rect 31066 -48318 31126 -48312
rect 32078 -48318 32138 -48312
rect 33098 -48318 33158 -48312
rect 36156 -48318 36216 -48312
rect 38194 -48318 38254 -48312
rect 41244 -48318 41304 -48312
rect 42262 -48318 42322 -48312
rect 43282 -48318 43342 -48312
rect 44298 -48318 44358 -48312
rect 46334 -48318 46394 -48312
rect 26986 -48374 27046 -48368
rect 27780 -48374 27840 -48368
rect 35140 -48374 35200 -48368
rect 37174 -48374 37234 -48368
rect 39204 -48374 39264 -48368
rect 49204 -48374 49264 -41181
rect 27046 -48434 27780 -48374
rect 27840 -48434 35140 -48374
rect 35200 -48434 37174 -48374
rect 37234 -48434 39204 -48374
rect 39264 -48434 49264 -48374
rect 26986 -48440 27046 -48434
rect 27780 -48440 27840 -48434
rect 35140 -48440 35200 -48434
rect 37174 -48440 37234 -48434
rect 39204 -48440 39264 -48434
rect 27668 -48488 27728 -48482
rect 28516 -48488 28576 -48482
rect 27728 -48548 28516 -48488
rect 27668 -48554 27728 -48548
rect 28516 -48554 28576 -48548
rect 30048 -48486 30108 -48480
rect 32084 -48486 32144 -48480
rect 48478 -48486 48538 -48480
rect 30108 -48546 32084 -48486
rect 32144 -48546 48478 -48486
rect 30048 -48552 30108 -48546
rect 32084 -48552 32144 -48546
rect 48478 -48552 48538 -48546
rect 48606 -48504 48666 -48498
rect 49206 -48504 49266 -48498
rect 48666 -48564 49206 -48504
rect 48606 -48570 48666 -48564
rect 49206 -48570 49266 -48564
rect -5312 -48778 -5212 -48769
rect -15855 -48852 -15765 -48848
rect -12999 -48850 -12909 -48846
rect -8060 -48850 -7960 -48841
rect -15860 -48857 -13656 -48852
rect -15860 -48947 -15855 -48857
rect -15765 -48947 -13656 -48857
rect -15860 -48952 -13656 -48947
rect -13004 -48855 -8060 -48850
rect -13004 -48945 -12999 -48855
rect -12909 -48945 -8060 -48855
rect -13004 -48950 -8060 -48945
rect -15855 -48956 -15765 -48952
rect -13756 -49148 -13656 -48952
rect -12999 -48954 -12909 -48950
rect -8060 -48959 -7960 -48950
rect -7431 -49046 -7341 -49042
rect -5312 -49046 -5212 -48878
rect -7436 -49051 -5212 -49046
rect -7436 -49141 -7431 -49051
rect -7341 -49141 -5212 -49051
rect -7436 -49146 -5212 -49141
rect -7431 -49150 -7341 -49146
rect -13756 -49257 -13656 -49248
rect 48372 -49374 48432 -49368
rect 49332 -49374 49392 -39098
rect 52262 -39086 55130 -39076
rect 56534 -39086 58154 -39076
rect 55130 -39386 55366 -39320
rect 52262 -39396 55366 -39386
rect 56534 -39396 58154 -39386
rect 53114 -40017 53174 -40011
rect 52006 -40077 53114 -40017
rect 53114 -40083 53174 -40077
rect 53264 -40256 53324 -40250
rect 54294 -40256 54354 -40250
rect 55186 -40256 55246 -40250
rect 53324 -40316 54294 -40256
rect 54354 -40316 55186 -40256
rect 53264 -40322 53324 -40316
rect 54294 -40322 54354 -40316
rect 55186 -40322 55246 -40316
rect 52380 -40374 52440 -40368
rect 53134 -40374 53194 -40368
rect 53392 -40374 53452 -40368
rect 54166 -40374 54226 -40368
rect 54426 -40374 54486 -40368
rect 52440 -40434 53134 -40374
rect 53194 -40434 53392 -40374
rect 53452 -40434 54166 -40374
rect 54226 -40434 54426 -40374
rect 52380 -40440 52440 -40434
rect 53134 -40440 53194 -40434
rect 53392 -40440 53452 -40434
rect 54166 -40440 54226 -40434
rect 54426 -40440 54486 -40434
rect 55004 -40374 55064 -40368
rect 55306 -40374 55366 -39396
rect 56318 -39666 56378 -39660
rect 56704 -39666 56764 -39660
rect 56962 -39666 57022 -39660
rect 57346 -39666 57406 -39660
rect 57986 -39666 58046 -39660
rect 56378 -39726 56704 -39666
rect 56764 -39726 56962 -39666
rect 57022 -39726 57346 -39666
rect 57406 -39726 57986 -39666
rect 56318 -39732 56378 -39726
rect 56704 -39732 56764 -39726
rect 56962 -39732 57022 -39726
rect 57346 -39732 57406 -39726
rect 57986 -39732 58046 -39726
rect 55064 -40434 55366 -40374
rect 55004 -40440 55064 -40434
rect 57474 -40476 57534 -40470
rect 57465 -40536 57474 -40476
rect 57534 -40536 57543 -40476
rect 55732 -40544 55792 -40538
rect 56318 -40544 56378 -40538
rect 56442 -40544 56502 -40538
rect 56704 -40544 56764 -40538
rect 56832 -40544 56892 -40538
rect 56958 -40544 57018 -40538
rect 57216 -40544 57276 -40538
rect 57346 -40544 57406 -40538
rect 57474 -40542 57534 -40536
rect 55792 -40604 56318 -40544
rect 56378 -40604 56442 -40544
rect 56502 -40604 56704 -40544
rect 56764 -40604 56832 -40544
rect 56892 -40604 56958 -40544
rect 57018 -40604 57216 -40544
rect 57276 -40604 57346 -40544
rect 55732 -40610 55792 -40604
rect 56318 -40610 56378 -40604
rect 56442 -40610 56502 -40604
rect 56704 -40610 56764 -40604
rect 56832 -40610 56892 -40604
rect 56958 -40610 57018 -40604
rect 57216 -40610 57276 -40604
rect 57346 -40610 57406 -40604
rect 52878 -41106 52938 -41100
rect 53132 -41106 53192 -41100
rect 53392 -41106 53452 -41100
rect 53650 -41106 53710 -41100
rect 53908 -41106 53968 -41100
rect 54166 -41106 54226 -41100
rect 54424 -41106 54484 -41100
rect 54682 -41106 54742 -41100
rect 51909 -41166 51918 -41106
rect 51978 -41166 52878 -41106
rect 52938 -41166 53132 -41106
rect 53192 -41166 53392 -41106
rect 53452 -41166 53650 -41106
rect 53710 -41166 53908 -41106
rect 53968 -41166 54166 -41106
rect 54226 -41166 54424 -41106
rect 54484 -41166 54682 -41106
rect 52878 -41172 52938 -41166
rect 53132 -41172 53192 -41166
rect 53392 -41172 53452 -41166
rect 53650 -41172 53710 -41166
rect 53908 -41172 53968 -41166
rect 54166 -41172 54226 -41166
rect 54424 -41172 54484 -41166
rect 54682 -41172 54742 -41166
rect 52748 -41226 52808 -41220
rect 53262 -41226 53322 -41220
rect 53778 -41226 53838 -41220
rect 54294 -41226 54354 -41220
rect 54806 -41226 54866 -41220
rect 55586 -41226 55646 -41220
rect 52808 -41286 53262 -41226
rect 53322 -41286 53778 -41226
rect 53838 -41286 54294 -41226
rect 54354 -41286 54806 -41226
rect 54866 -41286 55586 -41226
rect 52748 -41292 52808 -41286
rect 53262 -41292 53322 -41286
rect 53778 -41292 53838 -41286
rect 54294 -41292 54354 -41286
rect 54806 -41292 54866 -41286
rect 55586 -41292 55646 -41286
rect 56438 -41298 56498 -41292
rect 56828 -41298 56888 -41292
rect 57216 -41298 57276 -41292
rect 57986 -41298 58046 -41292
rect 56498 -41358 56828 -41298
rect 56888 -41358 57216 -41298
rect 57276 -41358 57986 -41298
rect 58046 -41358 58316 -41298
rect 56438 -41364 56498 -41358
rect 56828 -41364 56888 -41358
rect 57216 -41364 57276 -41358
rect 57986 -41364 58046 -41358
rect 56962 -41540 58094 -41480
rect 56962 -41874 57022 -41540
rect 57136 -41874 57196 -41868
rect 56962 -41934 57136 -41874
rect 52380 -41962 52440 -41953
rect 52874 -41962 52934 -41956
rect 53650 -41962 53710 -41956
rect 53906 -41962 53966 -41956
rect 54678 -41962 54738 -41956
rect 52440 -42022 52874 -41962
rect 52934 -42022 53650 -41962
rect 53710 -42022 53906 -41962
rect 53966 -42022 54678 -41962
rect 52380 -42031 52440 -42022
rect 52874 -42028 52934 -42022
rect 53650 -42028 53710 -42022
rect 53906 -42028 53966 -42022
rect 54678 -42028 54738 -42022
rect 56856 -41984 56916 -41978
rect 56962 -41984 57022 -41934
rect 57136 -41940 57196 -41934
rect 58034 -41932 58094 -41540
rect 58256 -41590 58316 -41358
rect 58256 -41656 58316 -41650
rect 56916 -42044 57022 -41984
rect 57128 -42044 57134 -41984
rect 57194 -42044 57200 -41984
rect 58034 -41992 58452 -41932
rect 56856 -42050 56916 -42044
rect 52746 -42078 52806 -42072
rect 52806 -42080 56064 -42078
rect 52806 -42138 53778 -42080
rect 52746 -42144 52806 -42138
rect 53772 -42140 53778 -42138
rect 53838 -42138 54808 -42080
rect 53838 -42140 53844 -42138
rect 53914 -42368 53974 -42138
rect 54802 -42140 54808 -42138
rect 54868 -42138 55186 -42080
rect 54868 -42140 54874 -42138
rect 55180 -42140 55186 -42138
rect 55246 -42138 56064 -42080
rect 55246 -42140 55252 -42138
rect 56004 -42178 56064 -42138
rect 57134 -42132 57194 -42044
rect 56004 -42238 56496 -42178
rect 57134 -42192 58450 -42132
rect 53914 -42434 53974 -42428
rect 54200 -42476 54260 -42470
rect 55295 -42471 55365 -42465
rect 51994 -42542 53314 -42482
rect 53374 -42542 53383 -42482
rect 54191 -42548 54200 -42476
rect 54260 -42548 54269 -42476
rect 54200 -42554 54260 -42548
rect 55286 -42553 55295 -42471
rect 55365 -42553 55374 -42471
rect 56436 -42502 56496 -42238
rect 55295 -42559 55365 -42553
rect 56436 -42562 56608 -42502
rect 56668 -42562 56674 -42502
rect 56042 -42572 56142 -42566
rect 56038 -42667 56042 -42577
rect 56142 -42667 56146 -42577
rect 56042 -42678 56142 -42672
rect 54846 -42716 54906 -42710
rect 54588 -42726 54648 -42720
rect 54332 -42736 54392 -42730
rect 54332 -43048 54392 -42796
rect 54332 -43114 54392 -43108
rect 54588 -43046 54648 -42786
rect 54588 -43112 54648 -43106
rect 54846 -43046 54906 -42776
rect 55098 -42718 55158 -42712
rect 55098 -43046 55158 -42778
rect 55232 -42716 55292 -42710
rect 55092 -43106 55098 -43046
rect 55158 -43106 55164 -43046
rect 55232 -43068 55292 -42776
rect 55732 -42958 55792 -42952
rect 56004 -42958 56064 -42952
rect 56120 -42958 56180 -42952
rect 56436 -42958 56496 -42562
rect 57946 -42574 58046 -42568
rect 57942 -42669 57946 -42579
rect 58046 -42669 58050 -42579
rect 57946 -42680 58046 -42674
rect 56912 -42928 56918 -42868
rect 56978 -42928 57138 -42868
rect 57198 -42928 57204 -42868
rect 55792 -43018 56004 -42958
rect 56114 -43018 56120 -42958
rect 56180 -43018 56496 -42958
rect 55732 -43024 55792 -43018
rect 56004 -43024 56064 -43018
rect 56120 -43024 56180 -43018
rect 55580 -43068 55586 -43066
rect 54846 -43112 54906 -43106
rect 55232 -43126 55586 -43068
rect 55646 -43068 55652 -43066
rect 56666 -43068 56726 -43062
rect 57020 -43068 57080 -42928
rect 58024 -42968 58084 -42962
rect 58256 -42968 58316 -42962
rect 58084 -43028 58256 -42968
rect 58024 -43034 58084 -43028
rect 58256 -43034 58316 -43028
rect 57374 -43068 57434 -43062
rect 57904 -43068 57964 -43062
rect 55646 -43126 56666 -43068
rect 55232 -43128 56666 -43126
rect 56726 -43128 57374 -43068
rect 57434 -43128 57904 -43068
rect 56666 -43134 56726 -43128
rect 57904 -43134 57964 -43128
rect 55824 -43278 58268 -43268
rect 55824 -43594 58268 -43584
rect 31064 -49392 31124 -49386
rect 33100 -49392 33160 -49386
rect 41244 -49392 41304 -49386
rect 43280 -49392 43340 -49386
rect 47354 -49392 47414 -49386
rect 27892 -49416 27952 -49410
rect 29030 -49416 29090 -49410
rect 27952 -49476 29030 -49416
rect 29090 -49476 29912 -49416
rect 31124 -49452 33100 -49392
rect 33160 -49452 41244 -49392
rect 41304 -49452 43280 -49392
rect 43340 -49452 47354 -49392
rect 48432 -49434 49392 -49374
rect 48372 -49440 48432 -49434
rect 31064 -49458 31124 -49452
rect 33100 -49458 33160 -49452
rect 41244 -49458 41304 -49452
rect 43280 -49458 43340 -49452
rect 47354 -49458 47414 -49452
rect 27892 -49482 27952 -49476
rect 29030 -49482 29090 -49476
rect 26982 -49616 27042 -49610
rect 27780 -49616 27840 -49610
rect 29028 -49616 29088 -49610
rect 27042 -49676 27780 -49616
rect 27840 -49676 29028 -49616
rect 29852 -49612 29912 -49476
rect 30046 -49496 30106 -49490
rect 32086 -49496 32146 -49490
rect 34118 -49496 34178 -49490
rect 36152 -49496 36212 -49490
rect 38192 -49496 38252 -49490
rect 40226 -49496 40286 -49490
rect 30106 -49556 32086 -49496
rect 32146 -49556 34118 -49496
rect 34178 -49556 36152 -49496
rect 36212 -49556 38192 -49496
rect 38252 -49556 40226 -49496
rect 30046 -49562 30106 -49556
rect 32086 -49562 32146 -49556
rect 34118 -49562 34178 -49556
rect 36152 -49562 36212 -49556
rect 38192 -49562 38252 -49556
rect 40226 -49562 40286 -49556
rect 40422 -49500 40482 -49494
rect 45314 -49500 45374 -49494
rect 40482 -49560 45314 -49500
rect 48972 -49504 49032 -49498
rect 40422 -49566 40482 -49560
rect 45314 -49566 45374 -49560
rect 45812 -49564 45818 -49504
rect 45878 -49564 48972 -49504
rect 48972 -49570 49032 -49564
rect 30560 -49610 30620 -49604
rect 34118 -49608 34178 -49602
rect 36154 -49608 36214 -49602
rect 38190 -49608 38250 -49602
rect 40226 -49608 40286 -49602
rect 42260 -49608 42320 -49602
rect 44298 -49608 44358 -49602
rect 46338 -49608 46398 -49602
rect 48722 -49608 48782 -49602
rect 29852 -49670 30560 -49612
rect 30620 -49670 31564 -49610
rect 31624 -49670 32576 -49610
rect 32636 -49670 33596 -49610
rect 33656 -49670 33662 -49610
rect 34178 -49668 36154 -49608
rect 36214 -49668 38190 -49608
rect 38250 -49668 40226 -49608
rect 40286 -49668 42260 -49608
rect 42320 -49668 44298 -49608
rect 44358 -49668 46338 -49608
rect 46398 -49668 48722 -49608
rect 29852 -49672 30902 -49670
rect 30560 -49676 30620 -49672
rect 34118 -49674 34178 -49668
rect 36154 -49674 36214 -49668
rect 38190 -49674 38250 -49668
rect 40226 -49674 40286 -49668
rect 42260 -49674 42320 -49668
rect 44298 -49674 44358 -49668
rect 46338 -49674 46398 -49668
rect 48722 -49674 48782 -49668
rect 26982 -49682 27042 -49676
rect 27780 -49682 27840 -49676
rect 29028 -49682 29088 -49676
rect 27104 -49718 27164 -49712
rect 27674 -49718 27734 -49712
rect 35136 -49718 35196 -49712
rect 37170 -49718 37230 -49712
rect 39210 -49718 39270 -49712
rect 40422 -49718 40482 -49712
rect 27164 -49778 27674 -49718
rect 27734 -49778 35136 -49718
rect 35196 -49778 37170 -49718
rect 37230 -49778 39210 -49718
rect 39270 -49778 40422 -49718
rect 27104 -49784 27164 -49778
rect 27674 -49784 27734 -49778
rect 35136 -49784 35196 -49778
rect 37170 -49784 37230 -49778
rect 39210 -49784 39270 -49778
rect 40422 -49784 40482 -49778
rect 40716 -49716 40776 -49710
rect 40776 -49776 41744 -49716
rect 41804 -49776 41810 -49716
rect 42262 -49722 42322 -49716
rect 44298 -49722 44358 -49716
rect 46336 -49722 46396 -49716
rect 48478 -49722 48538 -49716
rect 40716 -49782 40776 -49776
rect 42322 -49782 44298 -49722
rect 44358 -49782 46336 -49722
rect 46396 -49782 48478 -49722
rect 42262 -49788 42322 -49782
rect 44298 -49788 44358 -49782
rect 46336 -49788 46396 -49782
rect 48478 -49788 48538 -49782
rect 44810 -50636 44870 -50630
rect 29028 -50648 29088 -50642
rect 31066 -50648 31126 -50642
rect 33102 -50648 33162 -50642
rect 35134 -50648 35194 -50642
rect 29088 -50708 31066 -50648
rect 31126 -50708 33102 -50648
rect 33162 -50708 35134 -50648
rect 39710 -50696 39716 -50636
rect 39776 -50696 44810 -50636
rect 44810 -50702 44870 -50696
rect 44948 -50632 45008 -50626
rect 45830 -50632 45890 -50626
rect 46836 -50632 46896 -50626
rect 45008 -50692 45830 -50632
rect 45890 -50692 46836 -50632
rect 44948 -50698 45008 -50692
rect 45830 -50698 45890 -50692
rect 46836 -50698 46896 -50692
rect 47354 -50636 47414 -50630
rect 48606 -50636 48666 -50630
rect 47414 -50696 48606 -50636
rect 47354 -50702 47414 -50696
rect 48606 -50702 48666 -50696
rect 29028 -50714 29088 -50708
rect 31066 -50714 31126 -50708
rect 33102 -50714 33162 -50708
rect 35134 -50714 35194 -50708
rect 29534 -50750 29594 -50744
rect 34626 -50750 34686 -50744
rect 26594 -50800 26654 -50794
rect 29594 -50810 34626 -50750
rect 29534 -50816 29594 -50810
rect 34626 -50816 34686 -50810
rect 39210 -50764 39270 -50758
rect 47354 -50764 47414 -50758
rect 39270 -50824 47354 -50764
rect 39210 -50830 39270 -50824
rect 47354 -50830 47414 -50824
rect 22046 -51726 22106 -51720
rect 26594 -51726 26654 -50860
rect 26986 -50852 27046 -50846
rect 27780 -50852 27840 -50846
rect 31064 -50852 31124 -50846
rect 27046 -50912 27780 -50852
rect 27840 -50912 31064 -50852
rect 26986 -50918 27046 -50912
rect 27780 -50918 27840 -50912
rect 31064 -50918 31124 -50912
rect 31572 -50858 31632 -50852
rect 32594 -50858 32654 -50852
rect 33608 -50858 33668 -50852
rect 34626 -50858 34686 -50852
rect 35646 -50858 35706 -50852
rect 42758 -50858 42818 -50852
rect 43788 -50858 43848 -50852
rect 44948 -50858 45008 -50852
rect 31632 -50918 32594 -50858
rect 32654 -50918 33608 -50858
rect 33668 -50918 34626 -50858
rect 34686 -50918 35646 -50858
rect 35706 -50918 42758 -50858
rect 42818 -50918 43788 -50858
rect 43848 -50918 44948 -50858
rect 31572 -50924 31632 -50918
rect 32594 -50924 32654 -50918
rect 33608 -50924 33668 -50918
rect 34626 -50924 34686 -50918
rect 35646 -50924 35706 -50918
rect 42758 -50924 42818 -50918
rect 43788 -50924 43848 -50918
rect 44948 -50924 45008 -50918
rect 45316 -50858 45376 -50852
rect 48844 -50858 48904 -50852
rect 45376 -50918 48844 -50858
rect 45316 -50924 45376 -50918
rect 48844 -50924 48904 -50918
rect 30048 -50952 30108 -50946
rect 32082 -50952 32142 -50946
rect 34118 -50952 34178 -50946
rect 30108 -51012 32082 -50952
rect 32142 -51012 34118 -50952
rect 30048 -51018 30108 -51012
rect 32082 -51018 32142 -51012
rect 34118 -51018 34178 -51012
rect 41246 -50962 41306 -50956
rect 45316 -50962 45376 -50956
rect 41306 -51022 45316 -50962
rect 41246 -51028 41306 -51022
rect 45316 -51028 45376 -51022
rect 46332 -50960 46392 -50954
rect 48722 -50960 48782 -50954
rect 46392 -51020 48722 -50960
rect 46332 -51026 46392 -51020
rect 48722 -51026 48782 -51020
rect 22106 -51786 26654 -51726
rect 22046 -51792 22106 -51786
rect 20016 -51872 20076 -51866
rect 24076 -51872 24136 -51866
rect 26260 -51872 26320 -51866
rect 26726 -51872 26786 -51866
rect 36154 -51870 36214 -51864
rect 38190 -51870 38250 -51864
rect 40226 -51870 40286 -51864
rect 42264 -51870 42324 -51864
rect 15930 -51932 15936 -51872
rect 15996 -51932 20016 -51872
rect 20076 -51932 24076 -51872
rect 24136 -51932 26260 -51872
rect 26320 -51932 26726 -51872
rect 20016 -51938 20076 -51932
rect 24076 -51938 24136 -51932
rect 26260 -51938 26320 -51932
rect 26726 -51938 26786 -51932
rect 29530 -51876 29590 -51870
rect 30440 -51876 30500 -51870
rect 31442 -51876 31502 -51870
rect 32594 -51876 32654 -51870
rect 33604 -51876 33664 -51870
rect 34610 -51876 34670 -51870
rect 35654 -51876 35714 -51870
rect 29590 -51936 30440 -51876
rect 30500 -51936 31442 -51876
rect 31502 -51936 32594 -51876
rect 32654 -51936 33604 -51876
rect 33664 -51936 34610 -51876
rect 34670 -51936 35654 -51876
rect 36214 -51930 38190 -51870
rect 38250 -51930 40226 -51870
rect 40286 -51930 42264 -51870
rect 36154 -51936 36214 -51930
rect 38190 -51936 38250 -51930
rect 40226 -51936 40286 -51930
rect 42264 -51936 42324 -51930
rect 44300 -51870 44360 -51864
rect 46338 -51870 46398 -51864
rect 44360 -51930 46338 -51870
rect 44300 -51936 44360 -51930
rect 46338 -51936 46398 -51930
rect 29530 -51942 29590 -51936
rect 30440 -51942 30500 -51936
rect 31442 -51942 31502 -51936
rect 32594 -51942 32654 -51936
rect 33604 -51942 33664 -51936
rect 34610 -51942 34670 -51936
rect 35654 -51942 35714 -51936
rect 32082 -51978 32142 -51972
rect 42256 -51978 42316 -51972
rect 44296 -51978 44356 -51972
rect 46334 -51978 46394 -51972
rect 14775 -51987 14865 -51978
rect 17460 -52000 17520 -51994
rect 18492 -52000 18552 -51994
rect 21552 -52000 21612 -51994
rect 22548 -52000 22608 -51994
rect 26846 -52000 26906 -51994
rect 14865 -52060 17460 -52000
rect 17520 -52060 18492 -52000
rect 18552 -52060 21552 -52000
rect 21612 -52060 22548 -52000
rect 22608 -52060 26846 -52000
rect 32142 -52038 42256 -51978
rect 42316 -52038 44296 -51978
rect 44356 -52038 46334 -51978
rect 32082 -52044 32142 -52038
rect 42256 -52044 42316 -52038
rect 44296 -52044 44356 -52038
rect 46334 -52044 46394 -52038
rect 17460 -52066 17520 -52060
rect 18492 -52066 18552 -52060
rect 21552 -52066 21612 -52060
rect 22548 -52066 22608 -52060
rect 26846 -52066 26906 -52060
rect 14775 -52086 14865 -52077
rect 29530 -52092 29590 -52086
rect 31582 -52092 31642 -52086
rect 34608 -52092 34668 -52086
rect 35648 -52092 35708 -52086
rect 36662 -52092 36722 -52086
rect 37670 -52092 37730 -52086
rect 38714 -52092 38774 -52086
rect 39704 -52092 39764 -52086
rect 40722 -52092 40782 -52086
rect 41756 -52092 41816 -52086
rect 44788 -52092 44848 -52086
rect 45826 -52092 45886 -52086
rect 46852 -52092 46912 -52086
rect 29590 -52152 30568 -52092
rect 30628 -52152 31582 -52092
rect 31642 -52152 34608 -52092
rect 34668 -52152 35648 -52092
rect 35708 -52152 36662 -52092
rect 36722 -52152 37670 -52092
rect 37730 -52152 38714 -52092
rect 38774 -52152 39704 -52092
rect 39764 -52152 40722 -52092
rect 40782 -52152 41756 -52092
rect 41816 -52152 44788 -52092
rect 44848 -52152 45826 -52092
rect 45886 -52152 46852 -52092
rect 46912 -52152 48970 -52092
rect 49030 -52152 49036 -52092
rect 29530 -52158 29590 -52152
rect 31582 -52158 31642 -52152
rect 34608 -52158 34668 -52152
rect 35648 -52158 35708 -52152
rect 36662 -52158 36722 -52152
rect 37670 -52158 37730 -52152
rect 38714 -52158 38774 -52152
rect 39704 -52158 39764 -52152
rect 40722 -52158 40782 -52152
rect 41756 -52158 41816 -52152
rect 44788 -52158 44848 -52152
rect 45826 -52158 45886 -52152
rect 46852 -52158 46912 -52152
rect 35132 -52196 35192 -52190
rect 37174 -52196 37234 -52190
rect 39212 -52196 39272 -52190
rect 41246 -52196 41306 -52190
rect 43280 -52194 43340 -52188
rect 45314 -52194 45374 -52188
rect 47356 -52194 47416 -52188
rect 48606 -52194 48666 -52188
rect 27888 -52256 27894 -52196
rect 27954 -52256 35132 -52196
rect 35192 -52256 37174 -52196
rect 37234 -52256 39212 -52196
rect 39272 -52256 41246 -52196
rect 35132 -52262 35192 -52256
rect 37174 -52262 37234 -52256
rect 39212 -52262 39272 -52256
rect 41246 -52262 41306 -52256
rect 41758 -52200 41818 -52194
rect 42780 -52200 42840 -52194
rect 41818 -52260 42780 -52200
rect 43340 -52254 45314 -52194
rect 45374 -52254 47356 -52194
rect 47416 -52254 48606 -52194
rect 43280 -52260 43340 -52254
rect 45314 -52260 45374 -52254
rect 47356 -52260 47416 -52254
rect 48606 -52260 48666 -52254
rect 41758 -52266 41818 -52260
rect 42780 -52266 42840 -52260
rect 14767 -52948 14857 -52944
rect 14756 -53048 14762 -52948
rect 14862 -53048 14868 -52948
rect 16440 -52962 16500 -52956
rect 17464 -52962 17524 -52956
rect 18496 -52962 18556 -52956
rect 19496 -52962 19556 -52956
rect 20516 -52962 20576 -52956
rect 21536 -52962 21596 -52956
rect 23560 -52962 23620 -52956
rect 26380 -52962 26440 -52956
rect 26986 -52962 27046 -52956
rect 27782 -52962 27842 -52956
rect 16500 -53022 17464 -52962
rect 17524 -53022 18496 -52962
rect 18556 -53022 19496 -52962
rect 19556 -53022 20516 -52962
rect 20576 -53022 21536 -52962
rect 21596 -53022 22546 -52962
rect 22606 -53022 23560 -52962
rect 23620 -53022 24578 -52962
rect 24638 -53022 26380 -52962
rect 26440 -53022 26986 -52962
rect 27046 -53022 27782 -52962
rect 16440 -53028 16500 -53022
rect 17464 -53028 17524 -53022
rect 18496 -53028 18556 -53022
rect 19496 -53028 19556 -53022
rect 20516 -53028 20576 -53022
rect 21536 -53028 21596 -53022
rect 23560 -53028 23620 -53022
rect 26380 -53028 26440 -53022
rect 26986 -53028 27046 -53022
rect 27782 -53028 27842 -53022
rect 14767 -53052 14857 -53048
rect 15940 -53066 16000 -53060
rect 17976 -53066 18036 -53060
rect 20012 -53066 20072 -53060
rect 22046 -53066 22106 -53060
rect 24082 -53066 24142 -53060
rect 16000 -53126 17976 -53066
rect 18036 -53126 20012 -53066
rect 20072 -53126 22046 -53066
rect 22106 -53126 24082 -53066
rect 34122 -53098 34182 -53092
rect 38190 -53098 38250 -53092
rect 40224 -53098 40284 -53092
rect 15940 -53132 16000 -53126
rect 17976 -53132 18036 -53126
rect 20012 -53132 20072 -53126
rect 22046 -53132 22106 -53126
rect 24082 -53132 24142 -53126
rect 29528 -53104 29588 -53098
rect 30536 -53104 30596 -53098
rect 31550 -53104 31610 -53098
rect 32588 -53104 32648 -53098
rect 33606 -53104 33666 -53098
rect 29588 -53164 30536 -53104
rect 30596 -53164 31550 -53104
rect 31610 -53164 32588 -53104
rect 32648 -53164 33606 -53104
rect 34182 -53158 36158 -53098
rect 36218 -53158 38190 -53098
rect 38250 -53158 40224 -53098
rect 34122 -53164 34182 -53158
rect 38190 -53164 38250 -53158
rect 40224 -53164 40284 -53158
rect 41246 -53096 41306 -53090
rect 41600 -53096 41660 -53090
rect 41306 -53156 41600 -53096
rect 41246 -53162 41306 -53156
rect 41600 -53162 41660 -53156
rect 45318 -53096 45378 -53090
rect 48602 -53096 48662 -53090
rect 45378 -53156 48602 -53096
rect 45318 -53162 45378 -53156
rect 48602 -53162 48662 -53156
rect 21026 -53170 21086 -53164
rect 27564 -53170 27624 -53164
rect 29528 -53170 29588 -53164
rect 30536 -53170 30596 -53164
rect 31550 -53170 31610 -53164
rect 32588 -53170 32648 -53164
rect 33606 -53170 33666 -53164
rect 16952 -53230 16958 -53170
rect 17018 -53230 18994 -53170
rect 19054 -53230 21026 -53170
rect 21086 -53230 23060 -53170
rect 23120 -53230 25104 -53170
rect 25164 -53230 27564 -53170
rect 21026 -53236 21086 -53230
rect 27564 -53236 27624 -53230
rect 27674 -53208 27734 -53202
rect 29030 -53208 29090 -53202
rect 37174 -53208 37234 -53202
rect 39210 -53208 39270 -53202
rect 41242 -53208 41302 -53202
rect 27734 -53268 29030 -53208
rect 29090 -53268 37174 -53208
rect 37234 -53268 39210 -53208
rect 39270 -53268 41242 -53208
rect 27674 -53274 27734 -53268
rect 29030 -53274 29090 -53268
rect 37174 -53274 37234 -53268
rect 39210 -53274 39270 -53268
rect 41242 -53274 41302 -53268
rect 40752 -53306 40812 -53300
rect 41790 -53306 41850 -53300
rect 42766 -53306 42826 -53300
rect 43782 -53306 43842 -53300
rect 45808 -53306 45868 -53300
rect 46838 -53306 46898 -53300
rect 27332 -53320 27392 -53314
rect 30046 -53320 30106 -53314
rect 32084 -53320 32144 -53314
rect 36156 -53320 36216 -53314
rect 27392 -53380 30046 -53320
rect 30106 -53380 32084 -53320
rect 32144 -53380 36156 -53320
rect 40812 -53366 41790 -53306
rect 41850 -53366 42766 -53306
rect 42826 -53366 43782 -53306
rect 43842 -53366 45808 -53306
rect 45868 -53366 46838 -53306
rect 40752 -53372 40812 -53366
rect 41790 -53372 41850 -53366
rect 42766 -53372 42826 -53366
rect 43782 -53372 43842 -53366
rect 45808 -53372 45868 -53366
rect 46838 -53372 46898 -53366
rect 27332 -53386 27392 -53380
rect 30046 -53386 30106 -53380
rect 32084 -53386 32144 -53380
rect 36156 -53386 36216 -53380
rect 29026 -53418 29086 -53412
rect 31064 -53418 31124 -53412
rect 33104 -53418 33164 -53412
rect 35140 -53418 35200 -53412
rect 41244 -53418 41304 -53412
rect 41594 -53418 41600 -53414
rect 29086 -53478 31064 -53418
rect 31124 -53478 33104 -53418
rect 33164 -53478 35140 -53418
rect 35200 -53474 41600 -53418
rect 41660 -53418 41666 -53414
rect 43280 -53418 43340 -53412
rect 45316 -53418 45376 -53412
rect 47352 -53418 47412 -53412
rect 41660 -53474 43280 -53418
rect 35200 -53478 43280 -53474
rect 43340 -53478 45316 -53418
rect 45376 -53478 47352 -53418
rect 29026 -53484 29086 -53478
rect 31064 -53484 31124 -53478
rect 33104 -53484 33164 -53478
rect 35140 -53484 35200 -53478
rect 41244 -53484 41304 -53478
rect 43280 -53484 43340 -53478
rect 45316 -53484 45376 -53478
rect 47352 -53484 47412 -53478
rect 26380 -53564 26440 -53558
rect 27780 -53564 27840 -53558
rect 26440 -53624 27780 -53564
rect 26380 -53630 26440 -53624
rect 27780 -53630 27840 -53624
rect 14769 -53942 14859 -53938
rect 14758 -54042 14764 -53942
rect 14864 -54042 14870 -53942
rect 14769 -54046 14859 -54042
rect 17970 -54112 18030 -54106
rect 22046 -54112 22106 -54106
rect 26260 -54112 26320 -54106
rect 18030 -54172 22046 -54112
rect 22106 -54172 26260 -54112
rect 17970 -54178 18030 -54172
rect 22046 -54178 22106 -54172
rect 26260 -54178 26320 -54172
rect 14782 -54232 14842 -54226
rect 16432 -54232 16492 -54226
rect 19502 -54232 19562 -54226
rect 20510 -54232 20570 -54226
rect 23572 -54232 23632 -54226
rect 24598 -54232 24658 -54226
rect 14842 -54292 16432 -54232
rect 16492 -54292 19502 -54232
rect 19562 -54292 20510 -54232
rect 20570 -54292 23572 -54232
rect 23632 -54292 24598 -54232
rect 14782 -54298 14842 -54292
rect 16432 -54298 16492 -54292
rect 19502 -54298 19562 -54292
rect 20510 -54298 20570 -54292
rect 23572 -54298 23632 -54292
rect 24598 -54298 24658 -54292
rect 36152 -54322 36212 -54316
rect 38194 -54322 38254 -54316
rect 40226 -54322 40286 -54316
rect 42266 -54322 42326 -54316
rect 48722 -54322 48782 -54316
rect 30046 -54342 30106 -54336
rect 32082 -54342 32142 -54336
rect 34120 -54342 34180 -54336
rect 30106 -54402 32082 -54342
rect 32142 -54402 34120 -54342
rect 35976 -54382 35982 -54322
rect 36042 -54382 36152 -54322
rect 36212 -54382 38194 -54322
rect 38254 -54382 40226 -54322
rect 40286 -54382 42266 -54322
rect 42326 -54382 48722 -54322
rect 36152 -54388 36212 -54382
rect 38194 -54388 38254 -54382
rect 40226 -54388 40286 -54382
rect 42266 -54388 42326 -54382
rect 48722 -54388 48782 -54382
rect 30046 -54408 30106 -54402
rect 32082 -54408 32142 -54402
rect 34120 -54408 34180 -54402
rect 41244 -54420 41304 -54414
rect 47350 -54420 47410 -54414
rect 48602 -54420 48662 -54414
rect 27892 -54440 27952 -54434
rect 31064 -54440 31124 -54434
rect 27952 -54500 31064 -54440
rect 27892 -54506 27952 -54500
rect 31064 -54506 31124 -54500
rect 32588 -54440 32648 -54434
rect 35636 -54440 35696 -54434
rect 32648 -54500 33610 -54440
rect 33670 -54500 34632 -54440
rect 34692 -54500 35636 -54440
rect 41304 -54480 47350 -54420
rect 47410 -54480 48602 -54420
rect 41244 -54486 41304 -54480
rect 47350 -54486 47410 -54480
rect 48602 -54486 48662 -54480
rect 32588 -54506 32648 -54500
rect 35636 -54506 35696 -54500
rect 36158 -54530 36218 -54524
rect 38186 -54530 38246 -54524
rect 40230 -54530 40290 -54524
rect 42258 -54530 42318 -54524
rect 44296 -54530 44356 -54524
rect 46336 -54530 46396 -54524
rect 30050 -54536 30110 -54530
rect 32086 -54536 32146 -54530
rect 34114 -54536 34174 -54530
rect 35982 -54536 36042 -54530
rect 30110 -54596 32086 -54536
rect 32146 -54596 34114 -54536
rect 34174 -54596 35982 -54536
rect 36218 -54590 38186 -54530
rect 38246 -54590 40230 -54530
rect 40290 -54590 42258 -54530
rect 42318 -54590 44296 -54530
rect 44356 -54590 46336 -54530
rect 36158 -54596 36218 -54590
rect 38186 -54596 38246 -54590
rect 40230 -54596 40290 -54590
rect 42258 -54596 42318 -54590
rect 44296 -54596 44356 -54590
rect 46336 -54596 46396 -54590
rect 46854 -54526 46914 -54520
rect 48366 -54526 48426 -54520
rect 48972 -54526 49032 -54520
rect 46914 -54586 48366 -54526
rect 48426 -54586 48972 -54526
rect 46854 -54592 46914 -54586
rect 48366 -54592 48426 -54586
rect 48972 -54592 49032 -54586
rect 30050 -54602 30110 -54596
rect 32086 -54602 32146 -54596
rect 34114 -54602 34174 -54596
rect 35982 -54602 36042 -54596
rect 29032 -54656 29092 -54650
rect 33100 -54656 33160 -54650
rect 35134 -54656 35194 -54650
rect 43284 -54656 43344 -54650
rect 45314 -54656 45374 -54650
rect 47354 -54654 47414 -54648
rect 48844 -54654 48904 -54648
rect 29092 -54716 33100 -54656
rect 33160 -54716 35134 -54656
rect 35194 -54716 43284 -54656
rect 43344 -54716 45314 -54656
rect 45834 -54714 45840 -54654
rect 45900 -54714 47354 -54654
rect 47414 -54714 48844 -54654
rect 29032 -54722 29092 -54716
rect 33100 -54722 33160 -54716
rect 35134 -54722 35194 -54716
rect 43284 -54722 43344 -54716
rect 45314 -54722 45374 -54716
rect 47354 -54720 47414 -54714
rect 48844 -54720 48904 -54714
rect 14769 -54948 14859 -54944
rect 14758 -55048 14764 -54948
rect 14864 -55048 14870 -54948
rect 14769 -55052 14859 -55048
rect 25104 -55176 25164 -55170
rect 16952 -55236 16958 -55176
rect 17018 -55236 18994 -55176
rect 19054 -55236 21026 -55176
rect 21086 -55236 23060 -55176
rect 23120 -55236 25104 -55176
rect 25104 -55242 25164 -55236
rect 15944 -55284 16004 -55278
rect 17980 -55284 18040 -55278
rect 20016 -55284 20076 -55278
rect 22050 -55284 22110 -55278
rect 24086 -55284 24146 -55278
rect 16004 -55344 17980 -55284
rect 18040 -55344 20016 -55284
rect 20076 -55344 22050 -55284
rect 22110 -55344 24086 -55284
rect 15944 -55350 16004 -55344
rect 17980 -55350 18040 -55344
rect 20016 -55350 20076 -55344
rect 22050 -55350 22110 -55344
rect 24086 -55350 24146 -55344
rect 16438 -55396 16498 -55390
rect 17462 -55396 17522 -55390
rect 18494 -55396 18554 -55390
rect 19494 -55396 19554 -55390
rect 20514 -55396 20574 -55390
rect 21534 -55396 21594 -55390
rect 23558 -55396 23618 -55390
rect 26380 -55396 26440 -55390
rect 27780 -55396 27840 -55390
rect 16498 -55456 17462 -55396
rect 17522 -55456 18494 -55396
rect 18554 -55456 19494 -55396
rect 19554 -55456 20514 -55396
rect 20574 -55456 21534 -55396
rect 21594 -55456 22544 -55396
rect 22604 -55456 23558 -55396
rect 23618 -55456 24576 -55396
rect 24636 -55456 26380 -55396
rect 26440 -55456 27780 -55396
rect 16438 -55462 16498 -55456
rect 17462 -55462 17522 -55456
rect 18494 -55462 18554 -55456
rect 19494 -55462 19554 -55456
rect 20514 -55462 20574 -55456
rect 21534 -55462 21594 -55456
rect 23558 -55462 23618 -55456
rect 26380 -55462 26440 -55456
rect 27780 -55462 27840 -55456
rect 27780 -55572 27840 -55566
rect 37168 -55572 37228 -55566
rect 39210 -55572 39270 -55566
rect 41246 -55572 41306 -55566
rect 27840 -55632 37168 -55572
rect 37228 -55632 39210 -55572
rect 39270 -55632 41246 -55572
rect 27780 -55638 27840 -55632
rect 37168 -55638 37228 -55632
rect 39210 -55638 39270 -55632
rect 41246 -55638 41306 -55632
rect 44300 -55572 44360 -55566
rect 46332 -55572 46392 -55566
rect 48478 -55572 48538 -55566
rect 44360 -55632 46332 -55572
rect 46392 -55632 48478 -55572
rect 44300 -55638 44360 -55632
rect 46332 -55638 46392 -55632
rect 48478 -55638 48538 -55632
rect 31584 -55686 31644 -55680
rect 36664 -55686 36724 -55680
rect 27674 -55698 27734 -55692
rect 31064 -55698 31124 -55692
rect 27734 -55758 31064 -55698
rect 31644 -55746 36664 -55686
rect 31584 -55752 31644 -55746
rect 36664 -55752 36724 -55746
rect 41752 -55682 41812 -55676
rect 46852 -55682 46912 -55676
rect 41812 -55742 46852 -55682
rect 41752 -55748 41812 -55742
rect 46852 -55748 46912 -55742
rect 47860 -55682 47920 -55676
rect 49094 -55682 49154 -55676
rect 47920 -55742 49094 -55682
rect 47860 -55748 47920 -55742
rect 49094 -55748 49154 -55742
rect 27674 -55764 27734 -55758
rect 31064 -55764 31124 -55758
rect 30046 -55800 30106 -55794
rect 32082 -55800 32142 -55794
rect 33102 -55800 33162 -55794
rect 34118 -55800 34178 -55794
rect 35138 -55800 35198 -55794
rect 36156 -55800 36216 -55794
rect 38186 -55800 38246 -55794
rect 40224 -55800 40284 -55794
rect 42260 -55800 42320 -55794
rect 43282 -55800 43342 -55794
rect 44302 -55800 44362 -55794
rect 45316 -55800 45376 -55794
rect 46338 -55800 46398 -55794
rect 30106 -55860 32082 -55800
rect 32142 -55860 33102 -55800
rect 33162 -55860 34118 -55800
rect 34178 -55860 35138 -55800
rect 35198 -55860 36156 -55800
rect 36216 -55860 38186 -55800
rect 38246 -55860 40224 -55800
rect 40284 -55860 42260 -55800
rect 42320 -55860 43282 -55800
rect 43342 -55860 44302 -55800
rect 44362 -55860 45316 -55800
rect 45376 -55860 46338 -55800
rect 30046 -55866 30106 -55860
rect 32082 -55866 32142 -55860
rect 33102 -55866 33162 -55860
rect 34118 -55866 34178 -55860
rect 35138 -55866 35198 -55860
rect 36156 -55866 36216 -55860
rect 38186 -55866 38246 -55860
rect 40224 -55866 40284 -55860
rect 42260 -55866 42320 -55860
rect 43282 -55866 43342 -55860
rect 44302 -55866 44362 -55860
rect 45316 -55866 45376 -55860
rect 46338 -55866 46398 -55860
rect 31064 -55904 31124 -55898
rect 36000 -55904 36060 -55898
rect 42406 -55904 42466 -55898
rect 45316 -55904 45376 -55898
rect 48498 -55904 48558 -55898
rect 31124 -55964 36000 -55904
rect 36060 -55964 42406 -55904
rect 42466 -55964 45316 -55904
rect 45376 -55964 48498 -55904
rect 31064 -55970 31124 -55964
rect 36000 -55970 36060 -55964
rect 42406 -55970 42466 -55964
rect 45316 -55970 45376 -55964
rect 48498 -55970 48558 -55964
rect 14779 -56339 14869 -56330
rect 17452 -56358 17512 -56352
rect 18484 -56358 18544 -56352
rect 21544 -56358 21604 -56352
rect 22540 -56358 22600 -56352
rect 14869 -56418 17452 -56358
rect 17512 -56418 18484 -56358
rect 18544 -56418 21544 -56358
rect 21604 -56418 22540 -56358
rect 17452 -56424 17512 -56418
rect 18484 -56424 18544 -56418
rect 21544 -56424 21604 -56418
rect 22540 -56424 22600 -56418
rect 14779 -56438 14869 -56429
rect 20018 -56488 20078 -56482
rect 24078 -56488 24138 -56482
rect 26260 -56488 26320 -56482
rect 15932 -56548 15938 -56488
rect 15998 -56548 20018 -56488
rect 20078 -56548 24078 -56488
rect 24138 -56548 26260 -56488
rect 20018 -56554 20078 -56548
rect 24078 -56554 24138 -56548
rect 26260 -56554 26320 -56548
rect 9350 -56724 9452 -56700
rect 9350 -57518 9372 -56724
rect 9436 -57518 9452 -56724
rect 11554 -56780 11560 -56720
rect 11620 -56780 12236 -56720
rect 9350 -57536 9452 -57518
rect 10912 -57486 10972 -57480
rect 11430 -57486 11490 -57480
rect 10972 -57546 11430 -57486
rect 12176 -57532 12236 -56780
rect 27892 -56802 27952 -56796
rect 31062 -56802 31122 -56796
rect 27952 -56862 31062 -56802
rect 27892 -56868 27952 -56862
rect 31062 -56868 31122 -56862
rect 35292 -56800 35352 -56794
rect 37170 -56800 37230 -56794
rect 39208 -56800 39268 -56794
rect 41078 -56800 41138 -56794
rect 47354 -56800 47414 -56794
rect 35352 -56860 37170 -56800
rect 37230 -56860 39208 -56800
rect 39268 -56860 41078 -56800
rect 41138 -56860 47354 -56800
rect 35292 -56866 35352 -56860
rect 37170 -56866 37230 -56860
rect 39208 -56866 39268 -56860
rect 41078 -56866 41138 -56860
rect 47354 -56866 47414 -56860
rect 27564 -56906 27624 -56900
rect 29028 -56906 29088 -56900
rect 31068 -56906 31128 -56900
rect 33098 -56906 33158 -56900
rect 35138 -56906 35198 -56900
rect 37174 -56906 37234 -56900
rect 39210 -56906 39270 -56900
rect 41244 -56906 41304 -56900
rect 43284 -56906 43344 -56900
rect 45314 -56906 45374 -56900
rect 47354 -56906 47414 -56900
rect 49206 -56906 49266 -56900
rect 27624 -56966 29028 -56906
rect 29088 -56966 31068 -56906
rect 31128 -56966 33098 -56906
rect 33158 -56966 35138 -56906
rect 35198 -56966 37174 -56906
rect 37234 -56966 39210 -56906
rect 39270 -56966 41244 -56906
rect 41304 -56966 43284 -56906
rect 43344 -56966 45314 -56906
rect 45374 -56966 47354 -56906
rect 47414 -56966 49206 -56906
rect 27564 -56972 27624 -56966
rect 29028 -56972 29088 -56966
rect 31068 -56972 31128 -56966
rect 33098 -56972 33158 -56966
rect 35138 -56972 35198 -56966
rect 37174 -56972 37234 -56966
rect 39210 -56972 39270 -56966
rect 41244 -56972 41304 -56966
rect 43284 -56972 43344 -56966
rect 45314 -56972 45374 -56966
rect 47354 -56972 47414 -56966
rect 49206 -56972 49266 -56966
rect 29536 -57012 29596 -57006
rect 30556 -57012 30616 -57006
rect 31580 -57012 31640 -57006
rect 32598 -57012 32658 -57006
rect 33612 -57012 33672 -57006
rect 34644 -57012 34704 -57006
rect 35656 -57012 35716 -57006
rect 36664 -57012 36724 -57006
rect 37682 -57012 37742 -57006
rect 38708 -57012 38768 -57006
rect 39710 -57012 39770 -57006
rect 40730 -57012 40790 -57006
rect 41750 -57012 41810 -57006
rect 42776 -57012 42836 -57006
rect 43794 -57012 43854 -57006
rect 44808 -57012 44868 -57006
rect 45822 -57012 45882 -57006
rect 46844 -57012 46904 -57006
rect 29596 -57072 30556 -57012
rect 30616 -57072 31580 -57012
rect 31640 -57072 32598 -57012
rect 32658 -57072 33612 -57012
rect 33672 -57072 34644 -57012
rect 34704 -57072 35656 -57012
rect 35716 -57072 36664 -57012
rect 36724 -57072 37682 -57012
rect 37742 -57072 38708 -57012
rect 38768 -57072 39710 -57012
rect 39770 -57072 40730 -57012
rect 40790 -57072 41750 -57012
rect 41810 -57072 42776 -57012
rect 42836 -57072 43794 -57012
rect 43854 -57072 44808 -57012
rect 44868 -57072 45822 -57012
rect 45882 -57072 46844 -57012
rect 29536 -57078 29596 -57072
rect 30556 -57078 30616 -57072
rect 31580 -57078 31640 -57072
rect 32598 -57078 32658 -57072
rect 33612 -57078 33672 -57072
rect 34644 -57078 34704 -57072
rect 35656 -57078 35716 -57072
rect 36664 -57078 36724 -57072
rect 37682 -57078 37742 -57072
rect 38708 -57078 38768 -57072
rect 39710 -57078 39770 -57072
rect 40730 -57078 40790 -57072
rect 41750 -57078 41810 -57072
rect 42776 -57078 42836 -57072
rect 43794 -57078 43854 -57072
rect 44808 -57078 44868 -57072
rect 45822 -57078 45882 -57072
rect 46844 -57078 46904 -57072
rect 30048 -57122 30108 -57116
rect 32084 -57122 32144 -57116
rect 34122 -57122 34182 -57116
rect 36160 -57122 36220 -57116
rect 38196 -57122 38256 -57116
rect 40232 -57122 40292 -57116
rect 42264 -57122 42324 -57116
rect 44296 -57122 44356 -57116
rect 46336 -57122 46396 -57116
rect 30108 -57182 32084 -57122
rect 32144 -57182 34122 -57122
rect 34182 -57182 36160 -57122
rect 36220 -57182 38196 -57122
rect 38256 -57182 40232 -57122
rect 40292 -57182 42264 -57122
rect 42324 -57182 44296 -57122
rect 44356 -57182 46336 -57122
rect 30048 -57188 30108 -57182
rect 32084 -57188 32144 -57182
rect 34122 -57188 34182 -57182
rect 36160 -57188 36220 -57182
rect 38196 -57188 38256 -57182
rect 40232 -57188 40292 -57182
rect 42264 -57188 42324 -57182
rect 44296 -57188 44356 -57182
rect 46336 -57188 46396 -57182
rect 12524 -57532 12584 -57523
rect 10912 -57552 10972 -57546
rect 11430 -57552 11490 -57546
rect 12170 -57592 12176 -57532
rect 12236 -57592 12242 -57532
rect 12518 -57592 12524 -57532
rect 12584 -57592 12590 -57532
rect 12524 -57601 12584 -57592
rect 10654 -57635 10714 -57629
rect 11170 -57635 11230 -57629
rect 10643 -57695 10652 -57635
rect 10714 -57695 11170 -57635
rect 11230 -57695 11688 -57635
rect 11748 -57695 11754 -57635
rect 10654 -57701 10714 -57695
rect 11170 -57701 11230 -57695
rect 17416 -57854 17476 -57848
rect 19454 -57854 19514 -57848
rect 21490 -57854 21550 -57848
rect 23526 -57854 23586 -57848
rect 17476 -57914 19454 -57854
rect 19514 -57914 21490 -57854
rect 21550 -57914 23526 -57854
rect 17416 -57920 17476 -57914
rect 19454 -57920 19514 -57914
rect 21490 -57920 21550 -57914
rect 23526 -57920 23586 -57914
rect 18434 -57966 18494 -57960
rect 22508 -57966 22568 -57960
rect 26514 -57966 26574 -57960
rect 18494 -58026 22508 -57966
rect 22568 -58026 26514 -57966
rect 18434 -58032 18494 -58026
rect 22508 -58032 22568 -58026
rect 26514 -58032 26574 -58026
rect 27892 -58044 27952 -58038
rect 29028 -58044 29088 -58038
rect 33098 -58044 33158 -58038
rect 43278 -58044 43338 -58038
rect 48498 -58044 48558 -58038
rect 10914 -58074 10974 -58068
rect 10914 -58286 10974 -58134
rect 11430 -58074 11490 -58068
rect 27952 -58104 29028 -58044
rect 29088 -58104 33098 -58044
rect 33158 -58104 43278 -58044
rect 43338 -58104 48498 -58044
rect 27892 -58110 27952 -58104
rect 29028 -58110 29088 -58104
rect 33098 -58110 33158 -58104
rect 43278 -58110 43338 -58104
rect 48498 -58110 48558 -58104
rect 11430 -58286 11490 -58134
rect 29540 -58152 29600 -58146
rect 37684 -58152 37744 -58146
rect 11558 -58183 11618 -58177
rect 11618 -58243 12526 -58183
rect 12586 -58243 12595 -58183
rect 29600 -58212 30554 -58152
rect 30614 -58212 31576 -58152
rect 31636 -58212 32590 -58152
rect 32650 -58212 33616 -58152
rect 33676 -58212 34628 -58152
rect 34688 -58212 35664 -58152
rect 35724 -58212 36670 -58152
rect 36730 -58212 37684 -58152
rect 37744 -58212 38700 -58152
rect 38760 -58212 39708 -58152
rect 39768 -58212 40724 -58152
rect 40784 -58212 41748 -58152
rect 41808 -58212 42770 -58152
rect 42830 -58212 43792 -58152
rect 43852 -58212 44810 -58152
rect 44870 -58212 45824 -58152
rect 45884 -58212 46848 -58152
rect 46908 -58212 46914 -58152
rect 29540 -58218 29600 -58212
rect 37684 -58218 37744 -58212
rect 11558 -58249 11618 -58243
rect 10914 -58346 13076 -58286
rect 10276 -58408 12130 -58390
rect 10276 -58514 10294 -58408
rect 12110 -58514 12130 -58408
rect 10276 -58528 12130 -58514
rect 13016 -59714 13076 -58346
rect 17326 -58454 49412 -58408
rect 17326 -58608 17372 -58454
rect 49372 -58608 49412 -58454
rect 17326 -58654 49412 -58608
rect 13228 -58794 13828 -58784
rect 13228 -59104 13828 -59094
rect 49660 -58794 50260 -58784
rect 49660 -59104 50260 -59094
rect 13007 -59774 13016 -59714
rect 13076 -59774 13085 -59714
rect -9207 -64086 -9198 -64026
rect -9138 -64086 -9129 -64026
rect -27578 -64532 -26978 -64522
rect -27578 -64842 -26978 -64832
rect -26066 -64532 -25466 -64522
rect -26066 -64842 -25466 -64832
rect -23578 -64532 -22978 -64522
rect -23578 -64842 -22978 -64832
rect -22066 -64532 -21466 -64522
rect -22066 -64842 -21466 -64832
rect -19578 -64532 -18978 -64522
rect -19578 -64842 -18978 -64832
rect -18066 -64532 -17466 -64522
rect -18066 -64842 -17466 -64832
rect -15578 -64532 -14978 -64522
rect -15578 -64842 -14978 -64832
rect -14066 -64532 -13466 -64522
rect -14066 -64842 -13466 -64832
rect -11578 -64532 -10978 -64522
rect -11578 -64842 -10978 -64832
rect -10066 -64532 -9466 -64522
rect -10066 -64842 -9466 -64832
rect -27422 -65036 -25520 -65006
rect -27422 -65100 -27388 -65036
rect -25564 -65100 -25520 -65036
rect -27422 -65130 -25520 -65100
rect -23422 -65036 -21520 -65006
rect -23422 -65100 -23388 -65036
rect -21564 -65100 -21520 -65036
rect -23422 -65130 -21520 -65100
rect -19422 -65036 -17520 -65006
rect -19422 -65100 -19388 -65036
rect -17564 -65100 -17520 -65036
rect -19422 -65130 -17520 -65100
rect -15422 -65036 -13520 -65006
rect -15422 -65100 -15388 -65036
rect -13564 -65100 -13520 -65036
rect -15422 -65130 -13520 -65100
rect -11422 -65036 -9520 -65006
rect -11422 -65100 -11388 -65036
rect -9564 -65100 -9520 -65036
rect -11422 -65130 -9520 -65100
rect -25195 -65195 -25105 -65186
rect -26834 -65214 -26774 -65208
rect -26316 -65214 -26256 -65208
rect -26774 -65274 -26316 -65214
rect -26256 -65274 -25195 -65214
rect -26834 -65280 -26774 -65274
rect -26316 -65280 -26256 -65274
rect -21031 -65197 -20941 -65188
rect -22834 -65214 -22774 -65208
rect -22316 -65214 -22256 -65208
rect -22774 -65274 -22316 -65214
rect -22256 -65274 -21031 -65214
rect -22834 -65280 -22774 -65274
rect -22316 -65280 -22256 -65274
rect -25195 -65294 -25105 -65285
rect -17109 -65197 -17019 -65188
rect -18834 -65214 -18774 -65208
rect -18316 -65214 -18256 -65208
rect -18774 -65274 -18316 -65214
rect -18256 -65274 -17109 -65214
rect -18834 -65280 -18774 -65274
rect -18316 -65280 -18256 -65274
rect -21031 -65296 -20941 -65287
rect -17109 -65296 -17019 -65287
rect -16087 -65197 -15997 -65188
rect -14834 -65214 -14774 -65208
rect -14316 -65214 -14256 -65208
rect -15997 -65274 -14834 -65214
rect -14774 -65274 -14316 -65214
rect -14834 -65280 -14774 -65274
rect -14316 -65280 -14256 -65274
rect -10834 -65214 -10774 -65208
rect -10316 -65214 -10256 -65208
rect -9198 -65214 -9138 -64086
rect -7578 -64532 -6978 -64522
rect -7578 -64842 -6978 -64832
rect -6066 -64532 -5466 -64522
rect -6066 -64842 -5466 -64832
rect -3578 -64532 -2978 -64522
rect -3578 -64842 -2978 -64832
rect -2066 -64532 -1466 -64522
rect -2066 -64842 -1466 -64832
rect 422 -64532 1022 -64522
rect 422 -64842 1022 -64832
rect 1934 -64532 2534 -64522
rect 1934 -64842 2534 -64832
rect 4422 -64532 5022 -64522
rect 4422 -64842 5022 -64832
rect 5934 -64532 6534 -64522
rect 5934 -64842 6534 -64832
rect -7422 -65036 -5520 -65006
rect -7422 -65100 -7388 -65036
rect -5564 -65100 -5520 -65036
rect -7422 -65130 -5520 -65100
rect -3422 -65036 -1520 -65006
rect -3422 -65100 -3388 -65036
rect -1564 -65100 -1520 -65036
rect -3422 -65130 -1520 -65100
rect 578 -65036 2480 -65006
rect 578 -65100 612 -65036
rect 2436 -65100 2480 -65036
rect 578 -65130 2480 -65100
rect 4578 -65036 6480 -65006
rect 4578 -65100 4612 -65036
rect 6436 -65100 6480 -65036
rect 4578 -65130 6480 -65100
rect -4097 -65197 -4007 -65188
rect -6834 -65214 -6774 -65208
rect -6316 -65214 -6256 -65208
rect -10774 -65274 -10316 -65214
rect -10256 -65274 -9138 -65214
rect -7965 -65274 -7956 -65214
rect -7896 -65274 -6834 -65214
rect -6774 -65274 -6316 -65214
rect -10834 -65280 -10774 -65274
rect -10316 -65280 -10256 -65274
rect -6834 -65280 -6774 -65274
rect -6316 -65280 -6256 -65274
rect -16087 -65296 -15997 -65287
rect -39 -65201 51 -65192
rect -2834 -65214 -2774 -65208
rect -2316 -65214 -2256 -65208
rect -4007 -65274 -2834 -65214
rect -2774 -65274 -2316 -65214
rect -2834 -65280 -2774 -65274
rect -2316 -65280 -2256 -65274
rect -4097 -65296 -4007 -65287
rect 4015 -65199 4105 -65190
rect 1166 -65214 1226 -65208
rect 1684 -65214 1744 -65208
rect 51 -65274 1166 -65214
rect 1226 -65274 1684 -65214
rect 1166 -65280 1226 -65274
rect 1684 -65280 1744 -65274
rect -39 -65300 51 -65291
rect 5166 -65214 5226 -65208
rect 5684 -65214 5744 -65208
rect 4105 -65274 5166 -65214
rect 5226 -65274 5684 -65214
rect 5166 -65280 5226 -65274
rect 5684 -65280 5744 -65274
rect 4015 -65298 4105 -65289
rect -26578 -65326 -26518 -65320
rect -25648 -65326 -25588 -65320
rect -26518 -65386 -25648 -65326
rect -26578 -65392 -26518 -65386
rect -25648 -65392 -25588 -65386
rect -22578 -65326 -22518 -65320
rect -21648 -65326 -21588 -65320
rect -22518 -65386 -21648 -65326
rect -22578 -65392 -22518 -65386
rect -21648 -65392 -21588 -65386
rect -18578 -65326 -18518 -65320
rect -17648 -65326 -17588 -65320
rect -18518 -65386 -17648 -65326
rect -18578 -65392 -18518 -65386
rect -17648 -65392 -17588 -65386
rect -14578 -65326 -14518 -65320
rect -13648 -65326 -13588 -65320
rect -14518 -65386 -13648 -65326
rect -14578 -65392 -14518 -65386
rect -13648 -65392 -13588 -65386
rect -10578 -65326 -10518 -65320
rect -9648 -65326 -9588 -65320
rect -10518 -65386 -9648 -65326
rect -10578 -65392 -10518 -65386
rect -9648 -65392 -9588 -65386
rect -6578 -65326 -6518 -65320
rect -5648 -65326 -5588 -65320
rect -6518 -65386 -5648 -65326
rect -6578 -65392 -6518 -65386
rect -5648 -65392 -5588 -65386
rect -2578 -65326 -2518 -65320
rect -1648 -65326 -1588 -65320
rect -2518 -65386 -1648 -65326
rect -2578 -65392 -2518 -65386
rect -1648 -65392 -1588 -65386
rect 1422 -65326 1482 -65320
rect 2352 -65326 2412 -65320
rect 1482 -65386 2352 -65326
rect 1422 -65392 1482 -65386
rect 2352 -65392 2412 -65386
rect 5422 -65326 5482 -65320
rect 6352 -65326 6412 -65320
rect 5482 -65386 6352 -65326
rect 5422 -65392 5482 -65386
rect 6352 -65392 6412 -65386
rect -27496 -65446 -27436 -65440
rect -26706 -65446 -26646 -65440
rect -26450 -65446 -26390 -65440
rect -23496 -65446 -23436 -65440
rect -22706 -65446 -22646 -65440
rect -22450 -65446 -22390 -65440
rect -19496 -65446 -19436 -65440
rect -18706 -65446 -18646 -65440
rect -18450 -65446 -18390 -65440
rect -15496 -65446 -15436 -65440
rect -14706 -65446 -14646 -65440
rect -14450 -65446 -14390 -65440
rect -11496 -65446 -11436 -65440
rect -10706 -65446 -10646 -65440
rect -10450 -65446 -10390 -65440
rect -7496 -65446 -7436 -65440
rect -6706 -65446 -6646 -65440
rect -6450 -65446 -6390 -65440
rect -3496 -65446 -3436 -65440
rect -2706 -65446 -2646 -65440
rect -2450 -65446 -2390 -65440
rect 504 -65446 564 -65440
rect 1294 -65446 1354 -65440
rect 1550 -65446 1610 -65440
rect 4504 -65446 4564 -65440
rect 5294 -65446 5354 -65440
rect 5550 -65446 5610 -65440
rect -27436 -65506 -26706 -65446
rect -26646 -65506 -26450 -65446
rect -26388 -65506 -26379 -65446
rect -23436 -65506 -22706 -65446
rect -22646 -65506 -22450 -65446
rect -22388 -65506 -22379 -65446
rect -19436 -65506 -18706 -65446
rect -18646 -65506 -18450 -65446
rect -18390 -65506 -18381 -65446
rect -15436 -65506 -14706 -65446
rect -14646 -65506 -14450 -65446
rect -14390 -65506 -14381 -65446
rect -11436 -65506 -10706 -65446
rect -10646 -65506 -10450 -65446
rect -10390 -65506 -10381 -65446
rect -7436 -65506 -6706 -65446
rect -6646 -65506 -6450 -65446
rect -6388 -65506 -6379 -65446
rect -3436 -65506 -2706 -65446
rect -2646 -65506 -2452 -65446
rect -2390 -65506 -2383 -65446
rect 564 -65506 1294 -65446
rect 1354 -65506 1550 -65446
rect 1612 -65506 1621 -65446
rect 4564 -65506 5294 -65446
rect 5354 -65506 5550 -65446
rect 5614 -65506 5623 -65446
rect -27496 -65512 -27436 -65506
rect -26706 -65512 -26646 -65506
rect -26450 -65512 -26390 -65506
rect -23496 -65512 -23436 -65506
rect -22706 -65512 -22646 -65506
rect -22450 -65512 -22390 -65506
rect -19496 -65512 -19436 -65506
rect -18706 -65512 -18646 -65506
rect -18450 -65512 -18390 -65506
rect -15496 -65512 -15436 -65506
rect -14706 -65512 -14646 -65506
rect -14450 -65512 -14390 -65506
rect -11496 -65512 -11436 -65506
rect -10706 -65512 -10646 -65506
rect -10450 -65512 -10390 -65506
rect -7496 -65512 -7436 -65506
rect -6706 -65512 -6646 -65506
rect -6450 -65512 -6390 -65506
rect -3496 -65512 -3436 -65506
rect -2706 -65512 -2646 -65506
rect -2450 -65512 -2390 -65506
rect 504 -65512 564 -65506
rect 1294 -65512 1354 -65506
rect 1550 -65512 1610 -65506
rect 4504 -65512 4564 -65506
rect 5294 -65512 5354 -65506
rect 5550 -65512 5610 -65506
rect -28230 -66100 -27496 -66040
rect -27436 -66100 -27430 -66040
rect -24230 -66100 -23496 -66040
rect -23436 -66100 -23430 -66040
rect -20230 -66100 -19496 -66040
rect -19436 -66100 -19430 -66040
rect -16230 -66100 -15496 -66040
rect -15436 -66100 -15430 -66040
rect -12230 -66100 -11496 -66040
rect -11436 -66100 -11430 -66040
rect -8230 -66100 -7496 -66040
rect -7436 -66100 -7430 -66040
rect -4230 -66100 -3496 -66040
rect -3436 -66100 -3430 -66040
rect -230 -66100 504 -66040
rect 564 -66100 570 -66040
rect 3770 -66100 4504 -66040
rect 4564 -66100 4570 -66040
rect -28230 -67556 -28170 -66100
rect -26962 -66170 -26902 -66164
rect -26704 -66170 -26644 -66164
rect -26446 -66170 -26386 -66164
rect -26188 -66170 -26128 -66164
rect -27494 -66230 -26962 -66170
rect -26902 -66230 -26704 -66170
rect -26644 -66230 -26446 -66170
rect -26386 -66230 -26188 -66170
rect -28236 -67616 -28230 -67556
rect -28170 -67616 -28164 -67556
rect -27494 -67614 -27434 -66230
rect -26962 -66236 -26902 -66230
rect -26704 -66236 -26644 -66230
rect -26446 -66236 -26386 -66230
rect -26188 -66236 -26128 -66230
rect -27092 -66284 -27032 -66278
rect -26574 -66284 -26514 -66278
rect -26058 -66284 -25998 -66278
rect -27032 -66344 -26574 -66284
rect -26514 -66344 -26058 -66284
rect -27092 -66350 -27032 -66344
rect -26574 -66350 -26514 -66344
rect -26058 -66350 -25998 -66344
rect -27914 -67674 -27908 -67614
rect -27848 -67674 -27434 -67614
rect -27494 -68838 -27434 -67674
rect -27246 -67020 -27186 -67014
rect -26962 -67020 -26902 -67014
rect -26186 -67020 -26126 -67014
rect -27186 -67080 -26962 -67020
rect -26902 -67080 -26186 -67020
rect -27246 -68142 -27186 -67080
rect -26962 -67086 -26902 -67080
rect -26186 -67086 -26126 -67080
rect -27094 -67132 -27034 -67126
rect -26058 -67132 -25998 -67126
rect -25648 -67132 -25588 -67126
rect -27034 -67192 -26058 -67132
rect -25998 -67192 -25648 -67132
rect -27094 -67986 -27034 -67192
rect -26058 -67198 -25998 -67192
rect -25648 -67198 -25588 -67192
rect -26320 -67240 -26260 -67234
rect -26578 -67280 -26518 -67274
rect -26578 -67920 -26518 -67340
rect -26587 -67980 -26578 -67920
rect -26518 -67980 -26509 -67920
rect -27094 -68052 -27034 -68046
rect -26840 -68030 -26780 -68024
rect -26320 -68030 -26260 -67300
rect -24230 -67556 -24170 -66100
rect -22962 -66170 -22902 -66164
rect -22704 -66170 -22644 -66164
rect -22446 -66170 -22386 -66164
rect -22188 -66170 -22128 -66164
rect -23494 -66230 -22962 -66170
rect -22902 -66230 -22704 -66170
rect -22644 -66230 -22446 -66170
rect -22386 -66230 -22188 -66170
rect -24236 -67616 -24230 -67556
rect -24170 -67616 -24164 -67556
rect -23494 -67614 -23434 -66230
rect -22962 -66236 -22902 -66230
rect -22704 -66236 -22644 -66230
rect -22446 -66236 -22386 -66230
rect -22188 -66236 -22128 -66230
rect -23092 -66284 -23032 -66278
rect -22574 -66284 -22514 -66278
rect -22058 -66284 -21998 -66278
rect -23032 -66344 -22574 -66284
rect -22514 -66344 -22058 -66284
rect -23092 -66350 -23032 -66344
rect -22574 -66350 -22514 -66344
rect -22058 -66350 -21998 -66344
rect -23914 -67674 -23908 -67614
rect -23848 -67674 -23434 -67614
rect -26780 -68090 -26320 -68030
rect -26840 -68096 -26780 -68090
rect -26320 -68096 -26260 -68090
rect -26708 -68142 -26648 -68136
rect -26452 -68142 -26392 -68136
rect -27246 -68202 -26708 -68142
rect -26648 -68202 -26452 -68142
rect -26708 -68208 -26648 -68202
rect -26452 -68208 -26392 -68202
rect -26966 -68838 -26906 -68832
rect -26192 -68838 -26132 -68832
rect -27494 -68898 -26966 -68838
rect -26906 -68898 -26192 -68838
rect -23494 -68838 -23434 -67674
rect -23246 -67020 -23186 -67014
rect -22962 -67020 -22902 -67014
rect -22186 -67020 -22126 -67014
rect -23186 -67080 -22962 -67020
rect -22902 -67080 -22186 -67020
rect -23246 -68142 -23186 -67080
rect -22962 -67086 -22902 -67080
rect -22186 -67086 -22126 -67080
rect -23094 -67132 -23034 -67126
rect -22058 -67132 -21998 -67126
rect -21648 -67132 -21588 -67126
rect -23034 -67192 -22058 -67132
rect -21998 -67192 -21648 -67132
rect -23094 -67986 -23034 -67192
rect -22058 -67198 -21998 -67192
rect -21648 -67198 -21588 -67192
rect -22320 -67240 -22260 -67234
rect -22578 -67280 -22518 -67274
rect -22578 -67920 -22518 -67340
rect -22587 -67980 -22578 -67920
rect -22518 -67980 -22509 -67920
rect -23094 -68052 -23034 -68046
rect -22840 -68030 -22780 -68024
rect -22320 -68030 -22260 -67300
rect -20230 -67556 -20170 -66100
rect -18962 -66170 -18902 -66164
rect -18704 -66170 -18644 -66164
rect -18446 -66170 -18386 -66164
rect -18188 -66170 -18128 -66164
rect -19494 -66230 -18962 -66170
rect -18902 -66230 -18704 -66170
rect -18644 -66230 -18446 -66170
rect -18386 -66230 -18188 -66170
rect -20236 -67616 -20230 -67556
rect -20170 -67616 -20164 -67556
rect -19494 -67614 -19434 -66230
rect -18962 -66236 -18902 -66230
rect -18704 -66236 -18644 -66230
rect -18446 -66236 -18386 -66230
rect -18188 -66236 -18128 -66230
rect -19092 -66284 -19032 -66278
rect -18574 -66284 -18514 -66278
rect -18058 -66284 -17998 -66278
rect -19032 -66344 -18574 -66284
rect -18514 -66344 -18058 -66284
rect -19092 -66350 -19032 -66344
rect -18574 -66350 -18514 -66344
rect -18058 -66350 -17998 -66344
rect -19914 -67674 -19908 -67614
rect -19848 -67674 -19434 -67614
rect -22780 -68090 -22320 -68030
rect -22840 -68096 -22780 -68090
rect -22320 -68096 -22260 -68090
rect -22708 -68142 -22648 -68136
rect -22452 -68142 -22392 -68136
rect -23246 -68202 -22708 -68142
rect -22648 -68202 -22452 -68142
rect -22708 -68208 -22648 -68202
rect -22452 -68208 -22392 -68202
rect -22966 -68838 -22906 -68832
rect -22192 -68838 -22132 -68832
rect -23494 -68898 -22966 -68838
rect -22906 -68898 -22192 -68838
rect -19494 -68838 -19434 -67674
rect -19246 -67020 -19186 -67014
rect -18962 -67020 -18902 -67014
rect -18186 -67020 -18126 -67014
rect -19186 -67080 -18962 -67020
rect -18902 -67080 -18186 -67020
rect -19246 -68142 -19186 -67080
rect -18962 -67086 -18902 -67080
rect -18186 -67086 -18126 -67080
rect -19094 -67132 -19034 -67126
rect -18058 -67132 -17998 -67126
rect -17648 -67132 -17588 -67126
rect -19034 -67192 -18058 -67132
rect -17998 -67192 -17648 -67132
rect -19094 -67986 -19034 -67192
rect -18058 -67198 -17998 -67192
rect -17648 -67198 -17588 -67192
rect -18320 -67240 -18260 -67234
rect -18578 -67280 -18518 -67274
rect -18578 -67920 -18518 -67340
rect -18587 -67980 -18578 -67920
rect -18518 -67980 -18509 -67920
rect -19094 -68052 -19034 -68046
rect -18840 -68030 -18780 -68024
rect -18320 -68030 -18260 -67300
rect -16230 -67556 -16170 -66100
rect -14962 -66170 -14902 -66164
rect -14704 -66170 -14644 -66164
rect -14446 -66170 -14386 -66164
rect -14188 -66170 -14128 -66164
rect -15494 -66230 -14962 -66170
rect -14902 -66230 -14704 -66170
rect -14644 -66230 -14446 -66170
rect -14386 -66230 -14188 -66170
rect -16236 -67616 -16230 -67556
rect -16170 -67616 -16164 -67556
rect -15494 -67614 -15434 -66230
rect -14962 -66236 -14902 -66230
rect -14704 -66236 -14644 -66230
rect -14446 -66236 -14386 -66230
rect -14188 -66236 -14128 -66230
rect -15092 -66284 -15032 -66278
rect -14574 -66284 -14514 -66278
rect -14058 -66284 -13998 -66278
rect -15032 -66344 -14574 -66284
rect -14514 -66344 -14058 -66284
rect -15092 -66350 -15032 -66344
rect -14574 -66350 -14514 -66344
rect -14058 -66350 -13998 -66344
rect -15914 -67674 -15908 -67614
rect -15848 -67674 -15434 -67614
rect -18780 -68090 -18320 -68030
rect -18840 -68096 -18780 -68090
rect -18320 -68096 -18260 -68090
rect -18708 -68142 -18648 -68136
rect -18452 -68142 -18392 -68136
rect -19246 -68202 -18708 -68142
rect -18648 -68202 -18452 -68142
rect -18708 -68208 -18648 -68202
rect -18452 -68208 -18392 -68202
rect -18966 -68838 -18906 -68832
rect -18192 -68838 -18132 -68832
rect -19494 -68898 -18966 -68838
rect -18906 -68898 -18192 -68838
rect -15494 -68838 -15434 -67674
rect -15246 -67020 -15186 -67014
rect -14962 -67020 -14902 -67014
rect -14186 -67020 -14126 -67014
rect -15186 -67080 -14962 -67020
rect -14902 -67080 -14186 -67020
rect -15246 -68142 -15186 -67080
rect -14962 -67086 -14902 -67080
rect -14186 -67086 -14126 -67080
rect -15094 -67132 -15034 -67126
rect -14058 -67132 -13998 -67126
rect -13648 -67132 -13588 -67126
rect -15034 -67192 -14058 -67132
rect -13998 -67192 -13648 -67132
rect -15094 -67986 -15034 -67192
rect -14058 -67198 -13998 -67192
rect -13648 -67198 -13588 -67192
rect -14320 -67240 -14260 -67234
rect -14578 -67280 -14518 -67274
rect -14578 -67920 -14518 -67340
rect -14587 -67980 -14578 -67920
rect -14518 -67980 -14509 -67920
rect -15094 -68052 -15034 -68046
rect -14840 -68030 -14780 -68024
rect -14320 -68030 -14260 -67300
rect -12230 -67556 -12170 -66100
rect -10962 -66170 -10902 -66164
rect -10704 -66170 -10644 -66164
rect -10446 -66170 -10386 -66164
rect -10188 -66170 -10128 -66164
rect -11494 -66230 -10962 -66170
rect -10902 -66230 -10704 -66170
rect -10644 -66230 -10446 -66170
rect -10386 -66230 -10188 -66170
rect -12236 -67616 -12230 -67556
rect -12170 -67616 -12164 -67556
rect -11494 -67614 -11434 -66230
rect -10962 -66236 -10902 -66230
rect -10704 -66236 -10644 -66230
rect -10446 -66236 -10386 -66230
rect -10188 -66236 -10128 -66230
rect -11092 -66284 -11032 -66278
rect -10574 -66284 -10514 -66278
rect -10058 -66284 -9998 -66278
rect -11032 -66344 -10574 -66284
rect -10514 -66344 -10058 -66284
rect -11092 -66350 -11032 -66344
rect -10574 -66350 -10514 -66344
rect -10058 -66350 -9998 -66344
rect -11914 -67674 -11908 -67614
rect -11848 -67674 -11434 -67614
rect -14780 -68090 -14320 -68030
rect -14840 -68096 -14780 -68090
rect -14320 -68096 -14260 -68090
rect -14708 -68142 -14648 -68136
rect -14452 -68142 -14392 -68136
rect -15246 -68202 -14708 -68142
rect -14648 -68202 -14452 -68142
rect -14708 -68208 -14648 -68202
rect -14452 -68208 -14392 -68202
rect -14966 -68838 -14906 -68832
rect -14192 -68838 -14132 -68832
rect -15494 -68898 -14966 -68838
rect -14906 -68898 -14192 -68838
rect -11494 -68838 -11434 -67674
rect -11246 -67020 -11186 -67014
rect -10962 -67020 -10902 -67014
rect -10186 -67020 -10126 -67014
rect -11186 -67080 -10962 -67020
rect -10902 -67080 -10186 -67020
rect -11246 -68142 -11186 -67080
rect -10962 -67086 -10902 -67080
rect -10186 -67086 -10126 -67080
rect -11094 -67132 -11034 -67126
rect -10058 -67132 -9998 -67126
rect -9648 -67132 -9588 -67126
rect -11034 -67192 -10058 -67132
rect -9998 -67192 -9648 -67132
rect -11094 -67986 -11034 -67192
rect -10058 -67198 -9998 -67192
rect -9648 -67198 -9588 -67192
rect -10320 -67240 -10260 -67234
rect -10578 -67280 -10518 -67274
rect -10578 -67920 -10518 -67340
rect -10587 -67980 -10578 -67920
rect -10518 -67980 -10509 -67920
rect -11094 -68052 -11034 -68046
rect -10840 -68030 -10780 -68024
rect -10320 -68030 -10260 -67300
rect -8230 -67556 -8170 -66100
rect -6962 -66170 -6902 -66164
rect -6704 -66170 -6644 -66164
rect -6446 -66170 -6386 -66164
rect -6188 -66170 -6128 -66164
rect -7494 -66230 -6962 -66170
rect -6902 -66230 -6704 -66170
rect -6644 -66230 -6446 -66170
rect -6386 -66230 -6188 -66170
rect -8236 -67616 -8230 -67556
rect -8170 -67616 -8164 -67556
rect -7494 -67614 -7434 -66230
rect -6962 -66236 -6902 -66230
rect -6704 -66236 -6644 -66230
rect -6446 -66236 -6386 -66230
rect -6188 -66236 -6128 -66230
rect -7092 -66284 -7032 -66278
rect -6574 -66284 -6514 -66278
rect -6058 -66284 -5998 -66278
rect -7032 -66344 -6574 -66284
rect -6514 -66344 -6058 -66284
rect -7092 -66350 -7032 -66344
rect -6574 -66350 -6514 -66344
rect -6058 -66350 -5998 -66344
rect -7914 -67674 -7908 -67614
rect -7848 -67674 -7434 -67614
rect -10780 -68090 -10320 -68030
rect -10840 -68096 -10780 -68090
rect -10320 -68096 -10260 -68090
rect -10708 -68142 -10648 -68136
rect -10452 -68142 -10392 -68136
rect -11246 -68202 -10708 -68142
rect -10648 -68202 -10452 -68142
rect -10708 -68208 -10648 -68202
rect -10452 -68208 -10392 -68202
rect -10966 -68838 -10906 -68832
rect -10192 -68838 -10132 -68832
rect -11494 -68898 -10966 -68838
rect -10906 -68898 -10192 -68838
rect -7494 -68838 -7434 -67674
rect -7246 -67020 -7186 -67014
rect -6962 -67020 -6902 -67014
rect -6186 -67020 -6126 -67014
rect -7186 -67080 -6962 -67020
rect -6902 -67080 -6186 -67020
rect -7246 -68142 -7186 -67080
rect -6962 -67086 -6902 -67080
rect -6186 -67086 -6126 -67080
rect -7094 -67132 -7034 -67126
rect -6058 -67132 -5998 -67126
rect -5648 -67132 -5588 -67126
rect -7034 -67192 -6058 -67132
rect -5998 -67192 -5648 -67132
rect -7094 -67986 -7034 -67192
rect -6058 -67198 -5998 -67192
rect -5648 -67198 -5588 -67192
rect -6320 -67240 -6260 -67234
rect -6578 -67280 -6518 -67274
rect -6578 -67920 -6518 -67340
rect -6587 -67980 -6578 -67920
rect -6518 -67980 -6509 -67920
rect -7094 -68052 -7034 -68046
rect -6840 -68030 -6780 -68024
rect -6320 -68030 -6260 -67300
rect -4230 -67556 -4170 -66100
rect -2962 -66170 -2902 -66164
rect -2704 -66170 -2644 -66164
rect -2446 -66170 -2386 -66164
rect -2188 -66170 -2128 -66164
rect -3494 -66230 -2962 -66170
rect -2902 -66230 -2704 -66170
rect -2644 -66230 -2446 -66170
rect -2386 -66230 -2188 -66170
rect -4236 -67616 -4230 -67556
rect -4170 -67616 -4164 -67556
rect -3494 -67614 -3434 -66230
rect -2962 -66236 -2902 -66230
rect -2704 -66236 -2644 -66230
rect -2446 -66236 -2386 -66230
rect -2188 -66236 -2128 -66230
rect -3092 -66284 -3032 -66278
rect -2574 -66284 -2514 -66278
rect -2058 -66284 -1998 -66278
rect -3032 -66344 -2574 -66284
rect -2514 -66344 -2058 -66284
rect -3092 -66350 -3032 -66344
rect -2574 -66350 -2514 -66344
rect -2058 -66350 -1998 -66344
rect -3914 -67674 -3908 -67614
rect -3848 -67674 -3434 -67614
rect -6780 -68090 -6320 -68030
rect -6840 -68096 -6780 -68090
rect -6320 -68096 -6260 -68090
rect -6708 -68142 -6648 -68136
rect -6452 -68142 -6392 -68136
rect -7246 -68202 -6708 -68142
rect -6648 -68202 -6452 -68142
rect -6708 -68208 -6648 -68202
rect -6452 -68208 -6392 -68202
rect -6966 -68838 -6906 -68832
rect -6192 -68838 -6132 -68832
rect -7494 -68898 -6966 -68838
rect -6906 -68898 -6192 -68838
rect -3494 -68838 -3434 -67674
rect -3246 -67020 -3186 -67014
rect -2962 -67020 -2902 -67014
rect -2186 -67020 -2126 -67014
rect -3186 -67080 -2962 -67020
rect -2902 -67080 -2186 -67020
rect -3246 -68142 -3186 -67080
rect -2962 -67086 -2902 -67080
rect -2186 -67086 -2126 -67080
rect -3094 -67132 -3034 -67126
rect -2058 -67132 -1998 -67126
rect -1648 -67132 -1588 -67126
rect -3034 -67192 -2058 -67132
rect -1998 -67192 -1648 -67132
rect -3094 -67986 -3034 -67192
rect -2058 -67198 -1998 -67192
rect -1648 -67198 -1588 -67192
rect -2320 -67240 -2260 -67234
rect -2578 -67280 -2518 -67274
rect -2578 -67920 -2518 -67340
rect -2587 -67980 -2578 -67920
rect -2518 -67980 -2509 -67920
rect -3094 -68052 -3034 -68046
rect -2840 -68030 -2780 -68024
rect -2320 -68030 -2260 -67300
rect -230 -67556 -170 -66100
rect 1038 -66170 1098 -66164
rect 1296 -66170 1356 -66164
rect 1554 -66170 1614 -66164
rect 1812 -66170 1872 -66164
rect 506 -66230 1038 -66170
rect 1098 -66230 1296 -66170
rect 1356 -66230 1554 -66170
rect 1614 -66230 1812 -66170
rect -236 -67616 -230 -67556
rect -170 -67616 -164 -67556
rect 506 -67614 566 -66230
rect 1038 -66236 1098 -66230
rect 1296 -66236 1356 -66230
rect 1554 -66236 1614 -66230
rect 1812 -66236 1872 -66230
rect 908 -66284 968 -66278
rect 1426 -66284 1486 -66278
rect 1942 -66284 2002 -66278
rect 968 -66344 1426 -66284
rect 1486 -66344 1942 -66284
rect 908 -66350 968 -66344
rect 1426 -66350 1486 -66344
rect 1942 -66350 2002 -66344
rect 86 -67674 92 -67614
rect 152 -67674 566 -67614
rect -2780 -68090 -2320 -68030
rect -2840 -68096 -2780 -68090
rect -2320 -68096 -2260 -68090
rect -2708 -68142 -2648 -68136
rect -2452 -68142 -2392 -68136
rect -3246 -68202 -2708 -68142
rect -2648 -68202 -2452 -68142
rect -2708 -68208 -2648 -68202
rect -2452 -68208 -2392 -68202
rect -2966 -68838 -2906 -68832
rect -2192 -68838 -2132 -68832
rect -3494 -68898 -2966 -68838
rect -2906 -68898 -2192 -68838
rect 506 -68838 566 -67674
rect 754 -67020 814 -67014
rect 1038 -67020 1098 -67014
rect 1814 -67020 1874 -67014
rect 814 -67080 1038 -67020
rect 1098 -67080 1814 -67020
rect 754 -68142 814 -67080
rect 1038 -67086 1098 -67080
rect 1814 -67086 1874 -67080
rect 906 -67132 966 -67126
rect 1942 -67132 2002 -67126
rect 2352 -67132 2412 -67126
rect 966 -67192 1942 -67132
rect 2002 -67192 2352 -67132
rect 906 -67986 966 -67192
rect 1942 -67198 2002 -67192
rect 2352 -67198 2412 -67192
rect 1680 -67240 1740 -67234
rect 1422 -67280 1482 -67274
rect 1422 -67920 1482 -67340
rect 1413 -67980 1422 -67920
rect 1482 -67980 1491 -67920
rect 906 -68052 966 -68046
rect 1160 -68030 1220 -68024
rect 1680 -68030 1740 -67300
rect 3770 -67556 3830 -66100
rect 5038 -66170 5098 -66164
rect 5296 -66170 5356 -66164
rect 5554 -66170 5614 -66164
rect 5812 -66170 5872 -66164
rect 4506 -66230 5038 -66170
rect 5098 -66230 5296 -66170
rect 5356 -66230 5554 -66170
rect 5614 -66230 5812 -66170
rect 3764 -67616 3770 -67556
rect 3830 -67616 3836 -67556
rect 4506 -67614 4566 -66230
rect 5038 -66236 5098 -66230
rect 5296 -66236 5356 -66230
rect 5554 -66236 5614 -66230
rect 5812 -66236 5872 -66230
rect 4908 -66284 4968 -66278
rect 5426 -66284 5486 -66278
rect 5942 -66284 6002 -66278
rect 4968 -66344 5426 -66284
rect 5486 -66344 5942 -66284
rect 4908 -66350 4968 -66344
rect 5426 -66350 5486 -66344
rect 5942 -66350 6002 -66344
rect 4086 -67674 4092 -67614
rect 4152 -67674 4566 -67614
rect 1220 -68090 1680 -68030
rect 1160 -68096 1220 -68090
rect 1680 -68096 1740 -68090
rect 1292 -68142 1352 -68136
rect 1548 -68142 1608 -68136
rect 754 -68202 1292 -68142
rect 1352 -68202 1548 -68142
rect 1292 -68208 1352 -68202
rect 1548 -68208 1608 -68202
rect 1034 -68838 1094 -68832
rect 1808 -68838 1868 -68832
rect 506 -68898 1034 -68838
rect 1094 -68898 1808 -68838
rect 4506 -68838 4566 -67674
rect 4754 -67020 4814 -67014
rect 5038 -67020 5098 -67014
rect 5814 -67020 5874 -67014
rect 4814 -67080 5038 -67020
rect 5098 -67080 5814 -67020
rect 4754 -68142 4814 -67080
rect 5038 -67086 5098 -67080
rect 5814 -67086 5874 -67080
rect 4906 -67132 4966 -67126
rect 5942 -67132 6002 -67126
rect 6352 -67132 6412 -67126
rect 4966 -67192 5942 -67132
rect 6002 -67192 6352 -67132
rect 4906 -67986 4966 -67192
rect 5942 -67198 6002 -67192
rect 6352 -67198 6412 -67192
rect 5680 -67240 5740 -67234
rect 5422 -67280 5482 -67274
rect 5422 -67920 5482 -67340
rect 5416 -67922 5422 -67920
rect 5482 -67922 5488 -67920
rect 5413 -67982 5422 -67922
rect 5482 -67982 5491 -67922
rect 4906 -68052 4966 -68046
rect 5160 -68030 5220 -68024
rect 5680 -68030 5740 -67300
rect 5220 -68090 5680 -68030
rect 5160 -68096 5220 -68090
rect 5680 -68096 5740 -68090
rect 5292 -68142 5352 -68136
rect 5548 -68142 5608 -68136
rect 4754 -68202 5292 -68142
rect 5352 -68202 5548 -68142
rect 5292 -68208 5352 -68202
rect 5548 -68208 5608 -68202
rect 5034 -68838 5094 -68832
rect 5808 -68838 5868 -68832
rect 4506 -68898 5034 -68838
rect 5094 -68898 5808 -68838
rect -26966 -68904 -26906 -68898
rect -26192 -68904 -26132 -68898
rect -22966 -68904 -22906 -68898
rect -22192 -68904 -22132 -68898
rect -18966 -68904 -18906 -68898
rect -18192 -68904 -18132 -68898
rect -14966 -68904 -14906 -68898
rect -14192 -68904 -14132 -68898
rect -10966 -68904 -10906 -68898
rect -10192 -68904 -10132 -68898
rect -6966 -68904 -6906 -68898
rect -6192 -68904 -6132 -68898
rect -2966 -68904 -2906 -68898
rect -2192 -68904 -2132 -68898
rect 1034 -68904 1094 -68898
rect 1808 -68904 1868 -68898
rect 5034 -68904 5094 -68898
rect 5808 -68904 5868 -68898
rect -27100 -68952 -27040 -68946
rect -26064 -68952 -26004 -68946
rect -23100 -68952 -23040 -68946
rect -22064 -68952 -22004 -68946
rect -19100 -68952 -19040 -68946
rect -18064 -68952 -18004 -68946
rect -15100 -68952 -15040 -68946
rect -14064 -68952 -14004 -68946
rect -11100 -68952 -11040 -68946
rect -10064 -68952 -10004 -68946
rect -7100 -68952 -7040 -68946
rect -6064 -68952 -6004 -68946
rect -3100 -68952 -3040 -68946
rect -2064 -68952 -2004 -68946
rect 900 -68952 960 -68946
rect 1936 -68952 1996 -68946
rect 4900 -68952 4960 -68946
rect 5936 -68952 5996 -68946
rect -27040 -69012 -26064 -68952
rect -26004 -69012 -25232 -68952
rect -25172 -69012 -25163 -68952
rect -23040 -69012 -22064 -68952
rect -22004 -69012 -21232 -68952
rect -21172 -69012 -21163 -68952
rect -19040 -69012 -18064 -68952
rect -18004 -69012 -17232 -68952
rect -17172 -69012 -17163 -68952
rect -15040 -69012 -14064 -68952
rect -14004 -69012 -13232 -68952
rect -13172 -69012 -13163 -68952
rect -11040 -69012 -10064 -68952
rect -10004 -69012 -9232 -68952
rect -9172 -69012 -9163 -68952
rect -7040 -69012 -6064 -68952
rect -6004 -69012 -5232 -68952
rect -5172 -69012 -5163 -68952
rect -3040 -69012 -2064 -68952
rect -2004 -69012 -1232 -68952
rect -1172 -69012 -1163 -68952
rect 960 -69012 1936 -68952
rect 1996 -69012 2768 -68952
rect 2828 -69012 2837 -68952
rect 4960 -69012 5936 -68952
rect 5996 -69012 6768 -68952
rect 6828 -69012 6837 -68952
rect -27100 -69018 -27040 -69012
rect -26064 -69018 -26004 -69012
rect -23100 -69018 -23040 -69012
rect -22064 -69018 -22004 -69012
rect -19100 -69018 -19040 -69012
rect -18064 -69018 -18004 -69012
rect -15100 -69018 -15040 -69012
rect -14064 -69018 -14004 -69012
rect -11100 -69018 -11040 -69012
rect -10064 -69018 -10004 -69012
rect -7100 -69018 -7040 -69012
rect -6064 -69018 -6004 -69012
rect -3100 -69018 -3040 -69012
rect -2064 -69018 -2004 -69012
rect 900 -69018 960 -69012
rect 1936 -69018 1996 -69012
rect 4900 -69018 4960 -69012
rect 5936 -69018 5996 -69012
rect -27466 -69154 -25688 -69122
rect -27466 -69222 -27430 -69154
rect -25722 -69222 -25688 -69154
rect -27466 -69252 -25688 -69222
rect -23466 -69154 -21688 -69122
rect -23466 -69222 -23430 -69154
rect -21722 -69222 -21688 -69154
rect -23466 -69252 -21688 -69222
rect -19466 -69154 -17688 -69122
rect -19466 -69222 -19430 -69154
rect -17722 -69222 -17688 -69154
rect -19466 -69252 -17688 -69222
rect -15466 -69154 -13688 -69122
rect -15466 -69222 -15430 -69154
rect -13722 -69222 -13688 -69154
rect -15466 -69252 -13688 -69222
rect -11466 -69154 -9688 -69122
rect -11466 -69222 -11430 -69154
rect -9722 -69222 -9688 -69154
rect -11466 -69252 -9688 -69222
rect -7466 -69154 -5688 -69122
rect -7466 -69222 -7430 -69154
rect -5722 -69222 -5688 -69154
rect -7466 -69252 -5688 -69222
rect -3466 -69154 -1688 -69122
rect -3466 -69222 -3430 -69154
rect -1722 -69222 -1688 -69154
rect -3466 -69252 -1688 -69222
rect 534 -69154 2312 -69122
rect 534 -69222 570 -69154
rect 2278 -69222 2312 -69154
rect 534 -69252 2312 -69222
rect 4534 -69154 6312 -69122
rect 4534 -69222 4570 -69154
rect 6278 -69222 6312 -69154
rect 4534 -69252 6312 -69222
rect -27578 -69404 -26978 -69394
rect -27578 -69714 -26978 -69704
rect -26066 -69404 -25466 -69394
rect -26066 -69714 -25466 -69704
rect -23578 -69404 -22978 -69394
rect -23578 -69714 -22978 -69704
rect -22066 -69404 -21466 -69394
rect -22066 -69714 -21466 -69704
rect -19578 -69404 -18978 -69394
rect -19578 -69714 -18978 -69704
rect -18066 -69404 -17466 -69394
rect -18066 -69714 -17466 -69704
rect -15578 -69404 -14978 -69394
rect -15578 -69714 -14978 -69704
rect -14066 -69404 -13466 -69394
rect -14066 -69714 -13466 -69704
rect -11578 -69404 -10978 -69394
rect -11578 -69714 -10978 -69704
rect -10066 -69404 -9466 -69394
rect -10066 -69714 -9466 -69704
rect -7578 -69404 -6978 -69394
rect -7578 -69714 -6978 -69704
rect -6066 -69404 -5466 -69394
rect -6066 -69714 -5466 -69704
rect -3578 -69404 -2978 -69394
rect -3578 -69714 -2978 -69704
rect -2066 -69404 -1466 -69394
rect -2066 -69714 -1466 -69704
rect 422 -69404 1022 -69394
rect 422 -69714 1022 -69704
rect 1934 -69404 2534 -69394
rect 1934 -69714 2534 -69704
rect 4422 -69404 5022 -69394
rect 4422 -69714 5022 -69704
rect 5934 -69404 6534 -69394
rect 5934 -69714 6534 -69704
rect -27578 -70492 -26978 -70482
rect -27578 -70802 -26978 -70792
rect -26066 -70492 -25466 -70482
rect -26066 -70802 -25466 -70792
rect -23578 -70492 -22978 -70482
rect -23578 -70802 -22978 -70792
rect -22066 -70492 -21466 -70482
rect -22066 -70802 -21466 -70792
rect -19578 -70492 -18978 -70482
rect -19578 -70802 -18978 -70792
rect -18066 -70492 -17466 -70482
rect -18066 -70802 -17466 -70792
rect -15578 -70492 -14978 -70482
rect -15578 -70802 -14978 -70792
rect -14066 -70492 -13466 -70482
rect -14066 -70802 -13466 -70792
rect -11578 -70492 -10978 -70482
rect -11578 -70802 -10978 -70792
rect -10066 -70492 -9466 -70482
rect -10066 -70802 -9466 -70792
rect -7578 -70492 -6978 -70482
rect -7578 -70802 -6978 -70792
rect -6066 -70492 -5466 -70482
rect -6066 -70802 -5466 -70792
rect -3578 -70492 -2978 -70482
rect -3578 -70802 -2978 -70792
rect -2066 -70492 -1466 -70482
rect -2066 -70802 -1466 -70792
rect 422 -70492 1022 -70482
rect 422 -70802 1022 -70792
rect 1934 -70492 2534 -70482
rect 1934 -70802 2534 -70792
rect 4422 -70492 5022 -70482
rect 4422 -70802 5022 -70792
rect 5934 -70492 6534 -70482
rect 5934 -70802 6534 -70792
rect -27466 -70974 -25688 -70944
rect -27466 -71042 -27430 -70974
rect -25722 -71042 -25688 -70974
rect -27466 -71074 -25688 -71042
rect -23466 -70974 -21688 -70944
rect -23466 -71042 -23430 -70974
rect -21722 -71042 -21688 -70974
rect -23466 -71074 -21688 -71042
rect -19466 -70974 -17688 -70944
rect -19466 -71042 -19430 -70974
rect -17722 -71042 -17688 -70974
rect -19466 -71074 -17688 -71042
rect -15466 -70974 -13688 -70944
rect -15466 -71042 -15430 -70974
rect -13722 -71042 -13688 -70974
rect -15466 -71074 -13688 -71042
rect -11466 -70974 -9688 -70944
rect -11466 -71042 -11430 -70974
rect -9722 -71042 -9688 -70974
rect -11466 -71074 -9688 -71042
rect -7466 -70974 -5688 -70944
rect -7466 -71042 -7430 -70974
rect -5722 -71042 -5688 -70974
rect -7466 -71074 -5688 -71042
rect -3466 -70974 -1688 -70944
rect -3466 -71042 -3430 -70974
rect -1722 -71042 -1688 -70974
rect -3466 -71074 -1688 -71042
rect 534 -70974 2312 -70944
rect 534 -71042 570 -70974
rect 2278 -71042 2312 -70974
rect 534 -71074 2312 -71042
rect 4534 -70974 6312 -70944
rect 4534 -71042 4570 -70974
rect 6278 -71042 6312 -70974
rect 4534 -71074 6312 -71042
rect -27100 -71184 -27040 -71178
rect -26064 -71184 -26004 -71178
rect -27040 -71244 -26064 -71184
rect -27100 -71250 -27040 -71244
rect -26064 -71250 -26004 -71244
rect -23100 -71184 -23040 -71178
rect -22064 -71184 -22004 -71178
rect -23040 -71244 -22064 -71184
rect -23100 -71250 -23040 -71244
rect -22064 -71250 -22004 -71244
rect -19100 -71184 -19040 -71178
rect -18064 -71184 -18004 -71178
rect -19040 -71244 -18064 -71184
rect -19100 -71250 -19040 -71244
rect -18064 -71250 -18004 -71244
rect -15100 -71184 -15040 -71178
rect -14064 -71184 -14004 -71178
rect -15040 -71244 -14064 -71184
rect -15100 -71250 -15040 -71244
rect -14064 -71250 -14004 -71244
rect -11100 -71184 -11040 -71178
rect -10064 -71184 -10004 -71178
rect -11040 -71244 -10064 -71184
rect -11100 -71250 -11040 -71244
rect -10064 -71250 -10004 -71244
rect -7100 -71184 -7040 -71178
rect -6064 -71184 -6004 -71178
rect -7040 -71244 -6064 -71184
rect -7100 -71250 -7040 -71244
rect -6064 -71250 -6004 -71244
rect -3100 -71184 -3040 -71178
rect -2064 -71184 -2004 -71178
rect -3040 -71244 -2064 -71184
rect -3100 -71250 -3040 -71244
rect -2064 -71250 -2004 -71244
rect 900 -71184 960 -71178
rect 1936 -71184 1996 -71178
rect 960 -71244 1936 -71184
rect 900 -71250 960 -71244
rect 1936 -71250 1996 -71244
rect 4900 -71184 4960 -71178
rect 5936 -71184 5996 -71178
rect 4960 -71244 5936 -71184
rect 4900 -71250 4960 -71244
rect 5936 -71250 5996 -71244
rect -26966 -71298 -26906 -71292
rect -26192 -71298 -26132 -71292
rect -22966 -71298 -22906 -71292
rect -22192 -71298 -22132 -71292
rect -18966 -71298 -18906 -71292
rect -18192 -71298 -18132 -71292
rect -14966 -71298 -14906 -71292
rect -14192 -71298 -14132 -71292
rect -10966 -71298 -10906 -71292
rect -10192 -71298 -10132 -71292
rect -6966 -71298 -6906 -71292
rect -6192 -71298 -6132 -71292
rect -2966 -71298 -2906 -71292
rect -2192 -71298 -2132 -71292
rect 1034 -71298 1094 -71292
rect 1808 -71298 1868 -71292
rect 5034 -71298 5094 -71292
rect 5808 -71298 5868 -71292
rect -27494 -71358 -26966 -71298
rect -26906 -71358 -26192 -71298
rect -27494 -72522 -27434 -71358
rect -26966 -71364 -26906 -71358
rect -26192 -71364 -26132 -71358
rect -23494 -71358 -22966 -71298
rect -22906 -71358 -22192 -71298
rect -26708 -71994 -26648 -71988
rect -26452 -71994 -26392 -71988
rect -28236 -72640 -28230 -72580
rect -28170 -72640 -28164 -72580
rect -27914 -72582 -27908 -72522
rect -27848 -72582 -27434 -72522
rect -28230 -74096 -28170 -72640
rect -27494 -73966 -27434 -72582
rect -27246 -72054 -26708 -71994
rect -26648 -72054 -26452 -71994
rect -27246 -73116 -27186 -72054
rect -26708 -72060 -26648 -72054
rect -26452 -72060 -26392 -72054
rect -26840 -72106 -26780 -72100
rect -26320 -72106 -26260 -72100
rect -25238 -72106 -25178 -72097
rect -27094 -72150 -27034 -72144
rect -26780 -72166 -26320 -72106
rect -26260 -72166 -25238 -72106
rect -26840 -72172 -26780 -72166
rect -27094 -72882 -27034 -72210
rect -26584 -72276 -26578 -72216
rect -26518 -72276 -26512 -72216
rect -26578 -72856 -26518 -72276
rect -27103 -72942 -27094 -72882
rect -27034 -72942 -27025 -72882
rect -26578 -72922 -26518 -72916
rect -26320 -72896 -26260 -72166
rect -25238 -72175 -25178 -72166
rect -23494 -72522 -23434 -71358
rect -22966 -71364 -22906 -71358
rect -22192 -71364 -22132 -71358
rect -19494 -71358 -18966 -71298
rect -18906 -71358 -18192 -71298
rect -22708 -71994 -22648 -71988
rect -22452 -71994 -22392 -71988
rect -24236 -72640 -24230 -72580
rect -24170 -72640 -24164 -72580
rect -23914 -72582 -23908 -72522
rect -23848 -72582 -23434 -72522
rect -27094 -73004 -27034 -72942
rect -26320 -72962 -26260 -72956
rect -26058 -73004 -25998 -72998
rect -25648 -73004 -25588 -72998
rect -27034 -73064 -26058 -73004
rect -25998 -73064 -25648 -73004
rect -27094 -73070 -27034 -73064
rect -26058 -73070 -25998 -73064
rect -25648 -73070 -25588 -73064
rect -26962 -73116 -26902 -73110
rect -26186 -73116 -26126 -73110
rect -27186 -73176 -26962 -73116
rect -26902 -73176 -26186 -73116
rect -27246 -73182 -27186 -73176
rect -26962 -73182 -26902 -73176
rect -26186 -73182 -26126 -73176
rect -27092 -73852 -27032 -73846
rect -26574 -73852 -26514 -73846
rect -26058 -73852 -25998 -73846
rect -27032 -73912 -26574 -73852
rect -26514 -73912 -26058 -73852
rect -27092 -73918 -27032 -73912
rect -26574 -73918 -26514 -73912
rect -26058 -73918 -25998 -73912
rect -26962 -73966 -26902 -73960
rect -26704 -73966 -26644 -73960
rect -26446 -73966 -26386 -73960
rect -26188 -73966 -26128 -73960
rect -27494 -74026 -26962 -73966
rect -26902 -74026 -26704 -73966
rect -26644 -74026 -26446 -73966
rect -26386 -74026 -26188 -73966
rect -26962 -74032 -26902 -74026
rect -26704 -74032 -26644 -74026
rect -26446 -74032 -26386 -74026
rect -26188 -74032 -26128 -74026
rect -24230 -74096 -24170 -72640
rect -23494 -73966 -23434 -72582
rect -23246 -72054 -22708 -71994
rect -22648 -72054 -22452 -71994
rect -23246 -73116 -23186 -72054
rect -22708 -72060 -22648 -72054
rect -22452 -72060 -22392 -72054
rect -22840 -72106 -22780 -72100
rect -22320 -72106 -22260 -72100
rect -21238 -72106 -21178 -72097
rect -23094 -72150 -23034 -72144
rect -22780 -72166 -22320 -72106
rect -22260 -72166 -21238 -72106
rect -22840 -72172 -22780 -72166
rect -23094 -72882 -23034 -72210
rect -22584 -72276 -22578 -72216
rect -22518 -72276 -22512 -72216
rect -22578 -72856 -22518 -72276
rect -23103 -72942 -23094 -72882
rect -23034 -72942 -23025 -72882
rect -22578 -72922 -22518 -72916
rect -22320 -72896 -22260 -72166
rect -21238 -72175 -21178 -72166
rect -19494 -72522 -19434 -71358
rect -18966 -71364 -18906 -71358
rect -18192 -71364 -18132 -71358
rect -15494 -71358 -14966 -71298
rect -14906 -71358 -14192 -71298
rect -18708 -71994 -18648 -71988
rect -18452 -71994 -18392 -71988
rect -20236 -72640 -20230 -72580
rect -20170 -72640 -20164 -72580
rect -19914 -72582 -19908 -72522
rect -19848 -72582 -19434 -72522
rect -23094 -73004 -23034 -72942
rect -22320 -72962 -22260 -72956
rect -22058 -73004 -21998 -72998
rect -21648 -73004 -21588 -72998
rect -23034 -73064 -22058 -73004
rect -21998 -73064 -21648 -73004
rect -23094 -73070 -23034 -73064
rect -22058 -73070 -21998 -73064
rect -21648 -73070 -21588 -73064
rect -22962 -73116 -22902 -73110
rect -22186 -73116 -22126 -73110
rect -23186 -73176 -22962 -73116
rect -22902 -73176 -22186 -73116
rect -23246 -73182 -23186 -73176
rect -22962 -73182 -22902 -73176
rect -22186 -73182 -22126 -73176
rect -23092 -73852 -23032 -73846
rect -22574 -73852 -22514 -73846
rect -22058 -73852 -21998 -73846
rect -23032 -73912 -22574 -73852
rect -22514 -73912 -22058 -73852
rect -23092 -73918 -23032 -73912
rect -22574 -73918 -22514 -73912
rect -22058 -73918 -21998 -73912
rect -22962 -73966 -22902 -73960
rect -22704 -73966 -22644 -73960
rect -22446 -73966 -22386 -73960
rect -22188 -73966 -22128 -73960
rect -23494 -74026 -22962 -73966
rect -22902 -74026 -22704 -73966
rect -22644 -74026 -22446 -73966
rect -22386 -74026 -22188 -73966
rect -22962 -74032 -22902 -74026
rect -22704 -74032 -22644 -74026
rect -22446 -74032 -22386 -74026
rect -22188 -74032 -22128 -74026
rect -20230 -74096 -20170 -72640
rect -19494 -73966 -19434 -72582
rect -19246 -72054 -18708 -71994
rect -18648 -72054 -18452 -71994
rect -19246 -73116 -19186 -72054
rect -18708 -72060 -18648 -72054
rect -18452 -72060 -18392 -72054
rect -18840 -72106 -18780 -72100
rect -18320 -72106 -18260 -72100
rect -17238 -72106 -17178 -72097
rect -19094 -72150 -19034 -72144
rect -18780 -72166 -18320 -72106
rect -18260 -72166 -17238 -72106
rect -18840 -72172 -18780 -72166
rect -19094 -72882 -19034 -72210
rect -18584 -72276 -18578 -72216
rect -18518 -72276 -18512 -72216
rect -18578 -72856 -18518 -72276
rect -19103 -72942 -19094 -72882
rect -19034 -72942 -19025 -72882
rect -18578 -72922 -18518 -72916
rect -18320 -72896 -18260 -72166
rect -17238 -72175 -17178 -72166
rect -15494 -72522 -15434 -71358
rect -14966 -71364 -14906 -71358
rect -14192 -71364 -14132 -71358
rect -11494 -71358 -10966 -71298
rect -10906 -71358 -10192 -71298
rect -14708 -71994 -14648 -71988
rect -14452 -71994 -14392 -71988
rect -16236 -72640 -16230 -72580
rect -16170 -72640 -16164 -72580
rect -15914 -72582 -15908 -72522
rect -15848 -72582 -15434 -72522
rect -19094 -73004 -19034 -72942
rect -18320 -72962 -18260 -72956
rect -18058 -73004 -17998 -72998
rect -17648 -73004 -17588 -72998
rect -19034 -73064 -18058 -73004
rect -17998 -73064 -17648 -73004
rect -19094 -73070 -19034 -73064
rect -18058 -73070 -17998 -73064
rect -17648 -73070 -17588 -73064
rect -18962 -73116 -18902 -73110
rect -18186 -73116 -18126 -73110
rect -19186 -73176 -18962 -73116
rect -18902 -73176 -18186 -73116
rect -19246 -73182 -19186 -73176
rect -18962 -73182 -18902 -73176
rect -18186 -73182 -18126 -73176
rect -19092 -73852 -19032 -73846
rect -18574 -73852 -18514 -73846
rect -18058 -73852 -17998 -73846
rect -19032 -73912 -18574 -73852
rect -18514 -73912 -18058 -73852
rect -19092 -73918 -19032 -73912
rect -18574 -73918 -18514 -73912
rect -18058 -73918 -17998 -73912
rect -18962 -73966 -18902 -73960
rect -18704 -73966 -18644 -73960
rect -18446 -73966 -18386 -73960
rect -18188 -73966 -18128 -73960
rect -19494 -74026 -18962 -73966
rect -18902 -74026 -18704 -73966
rect -18644 -74026 -18446 -73966
rect -18386 -74026 -18188 -73966
rect -18962 -74032 -18902 -74026
rect -18704 -74032 -18644 -74026
rect -18446 -74032 -18386 -74026
rect -18188 -74032 -18128 -74026
rect -16230 -74096 -16170 -72640
rect -15494 -73966 -15434 -72582
rect -15246 -72054 -14708 -71994
rect -14648 -72054 -14452 -71994
rect -15246 -73116 -15186 -72054
rect -14708 -72060 -14648 -72054
rect -14452 -72060 -14392 -72054
rect -14840 -72106 -14780 -72100
rect -14320 -72106 -14260 -72100
rect -13238 -72106 -13178 -72097
rect -15094 -72150 -15034 -72144
rect -14780 -72166 -14320 -72106
rect -14260 -72166 -13238 -72106
rect -14840 -72172 -14780 -72166
rect -15094 -72882 -15034 -72210
rect -14584 -72276 -14578 -72216
rect -14518 -72276 -14512 -72216
rect -14578 -72856 -14518 -72276
rect -15103 -72942 -15094 -72882
rect -15034 -72942 -15025 -72882
rect -14578 -72922 -14518 -72916
rect -14320 -72896 -14260 -72166
rect -13238 -72175 -13178 -72166
rect -11494 -72522 -11434 -71358
rect -10966 -71364 -10906 -71358
rect -10192 -71364 -10132 -71358
rect -7494 -71358 -6966 -71298
rect -6906 -71358 -6192 -71298
rect -10708 -71994 -10648 -71988
rect -10452 -71994 -10392 -71988
rect -12236 -72640 -12230 -72580
rect -12170 -72640 -12164 -72580
rect -11914 -72582 -11908 -72522
rect -11848 -72582 -11434 -72522
rect -15094 -73004 -15034 -72942
rect -14320 -72962 -14260 -72956
rect -14058 -73004 -13998 -72998
rect -13648 -73004 -13588 -72998
rect -15034 -73064 -14058 -73004
rect -13998 -73064 -13648 -73004
rect -15094 -73070 -15034 -73064
rect -14058 -73070 -13998 -73064
rect -13648 -73070 -13588 -73064
rect -14962 -73116 -14902 -73110
rect -14186 -73116 -14126 -73110
rect -15186 -73176 -14962 -73116
rect -14902 -73176 -14186 -73116
rect -15246 -73182 -15186 -73176
rect -14962 -73182 -14902 -73176
rect -14186 -73182 -14126 -73176
rect -15092 -73852 -15032 -73846
rect -14574 -73852 -14514 -73846
rect -14058 -73852 -13998 -73846
rect -15032 -73912 -14574 -73852
rect -14514 -73912 -14058 -73852
rect -15092 -73918 -15032 -73912
rect -14574 -73918 -14514 -73912
rect -14058 -73918 -13998 -73912
rect -14962 -73966 -14902 -73960
rect -14704 -73966 -14644 -73960
rect -14446 -73966 -14386 -73960
rect -14188 -73966 -14128 -73960
rect -15494 -74026 -14962 -73966
rect -14902 -74026 -14704 -73966
rect -14644 -74026 -14446 -73966
rect -14386 -74026 -14188 -73966
rect -14962 -74032 -14902 -74026
rect -14704 -74032 -14644 -74026
rect -14446 -74032 -14386 -74026
rect -14188 -74032 -14128 -74026
rect -12230 -74096 -12170 -72640
rect -11494 -73966 -11434 -72582
rect -11246 -72054 -10708 -71994
rect -10648 -72054 -10452 -71994
rect -11246 -73116 -11186 -72054
rect -10708 -72060 -10648 -72054
rect -10452 -72060 -10392 -72054
rect -10840 -72106 -10780 -72100
rect -10320 -72106 -10260 -72100
rect -9238 -72106 -9178 -72097
rect -11094 -72150 -11034 -72144
rect -10780 -72166 -10320 -72106
rect -10260 -72166 -9238 -72106
rect -10840 -72172 -10780 -72166
rect -11094 -72880 -11034 -72210
rect -10584 -72276 -10578 -72216
rect -10518 -72276 -10512 -72216
rect -10578 -72856 -10518 -72276
rect -11103 -72940 -11094 -72880
rect -11034 -72940 -11025 -72880
rect -10578 -72922 -10518 -72916
rect -10320 -72896 -10260 -72166
rect -9238 -72175 -9178 -72166
rect -7494 -72522 -7434 -71358
rect -6966 -71364 -6906 -71358
rect -6192 -71364 -6132 -71358
rect -3494 -71358 -2966 -71298
rect -2906 -71358 -2192 -71298
rect -6708 -71994 -6648 -71988
rect -6452 -71994 -6392 -71988
rect -8236 -72640 -8230 -72580
rect -8170 -72640 -8164 -72580
rect -7914 -72582 -7908 -72522
rect -7848 -72582 -7434 -72522
rect -11094 -73004 -11034 -72940
rect -10320 -72962 -10260 -72956
rect -10058 -73004 -9998 -72998
rect -9648 -73004 -9588 -72998
rect -11034 -73064 -10058 -73004
rect -9998 -73064 -9648 -73004
rect -11094 -73070 -11034 -73064
rect -10058 -73070 -9998 -73064
rect -9648 -73070 -9588 -73064
rect -10962 -73116 -10902 -73110
rect -10186 -73116 -10126 -73110
rect -11186 -73176 -10962 -73116
rect -10902 -73176 -10186 -73116
rect -11246 -73182 -11186 -73176
rect -10962 -73182 -10902 -73176
rect -10186 -73182 -10126 -73176
rect -11092 -73852 -11032 -73846
rect -10574 -73852 -10514 -73846
rect -10058 -73852 -9998 -73846
rect -11032 -73912 -10574 -73852
rect -10514 -73912 -10058 -73852
rect -11092 -73918 -11032 -73912
rect -10574 -73918 -10514 -73912
rect -10058 -73918 -9998 -73912
rect -10962 -73966 -10902 -73960
rect -10704 -73966 -10644 -73960
rect -10446 -73966 -10386 -73960
rect -10188 -73966 -10128 -73960
rect -11494 -74026 -10962 -73966
rect -10902 -74026 -10704 -73966
rect -10644 -74026 -10446 -73966
rect -10386 -74026 -10188 -73966
rect -10962 -74032 -10902 -74026
rect -10704 -74032 -10644 -74026
rect -10446 -74032 -10386 -74026
rect -10188 -74032 -10128 -74026
rect -8230 -74096 -8170 -72640
rect -7494 -73966 -7434 -72582
rect -7246 -72054 -6708 -71994
rect -6648 -72054 -6452 -71994
rect -7246 -73116 -7186 -72054
rect -6708 -72060 -6648 -72054
rect -6452 -72060 -6392 -72054
rect -6840 -72106 -6780 -72100
rect -6320 -72106 -6260 -72100
rect -5238 -72106 -5178 -72097
rect -7094 -72150 -7034 -72144
rect -6780 -72166 -6320 -72106
rect -6260 -72166 -5238 -72106
rect -6840 -72172 -6780 -72166
rect -7094 -72882 -7034 -72210
rect -6584 -72276 -6578 -72216
rect -6518 -72276 -6512 -72216
rect -6578 -72856 -6518 -72276
rect -7103 -72942 -7094 -72882
rect -7034 -72942 -7025 -72882
rect -6578 -72922 -6518 -72916
rect -6320 -72896 -6260 -72166
rect -5238 -72175 -5178 -72166
rect -3494 -72522 -3434 -71358
rect -2966 -71364 -2906 -71358
rect -2192 -71364 -2132 -71358
rect 506 -71358 1034 -71298
rect 1094 -71358 1808 -71298
rect -2708 -71994 -2648 -71988
rect -2452 -71994 -2392 -71988
rect -4236 -72640 -4230 -72580
rect -4170 -72640 -4164 -72580
rect -3914 -72582 -3908 -72522
rect -3848 -72582 -3434 -72522
rect -7094 -73004 -7034 -72942
rect -6320 -72962 -6260 -72956
rect -6058 -73004 -5998 -72998
rect -5648 -73004 -5588 -72998
rect -7034 -73064 -6058 -73004
rect -5998 -73064 -5648 -73004
rect -7094 -73070 -7034 -73064
rect -6058 -73070 -5998 -73064
rect -5648 -73070 -5588 -73064
rect -6962 -73116 -6902 -73110
rect -6186 -73116 -6126 -73110
rect -7186 -73176 -6962 -73116
rect -6902 -73176 -6186 -73116
rect -7246 -73182 -7186 -73176
rect -6962 -73182 -6902 -73176
rect -6186 -73182 -6126 -73176
rect -7092 -73852 -7032 -73846
rect -6574 -73852 -6514 -73846
rect -6058 -73852 -5998 -73846
rect -7032 -73912 -6574 -73852
rect -6514 -73912 -6058 -73852
rect -7092 -73918 -7032 -73912
rect -6574 -73918 -6514 -73912
rect -6058 -73918 -5998 -73912
rect -6962 -73966 -6902 -73960
rect -6704 -73966 -6644 -73960
rect -6446 -73966 -6386 -73960
rect -6188 -73966 -6128 -73960
rect -7494 -74026 -6962 -73966
rect -6902 -74026 -6704 -73966
rect -6644 -74026 -6446 -73966
rect -6386 -74026 -6188 -73966
rect -6962 -74032 -6902 -74026
rect -6704 -74032 -6644 -74026
rect -6446 -74032 -6386 -74026
rect -6188 -74032 -6128 -74026
rect -4230 -74096 -4170 -72640
rect -3494 -73966 -3434 -72582
rect -3246 -72054 -2708 -71994
rect -2648 -72054 -2452 -71994
rect -3246 -72332 -3186 -72054
rect -2708 -72060 -2648 -72054
rect -2452 -72060 -2392 -72054
rect -2840 -72106 -2780 -72100
rect -2320 -72106 -2260 -72100
rect -1238 -72106 -1178 -72097
rect -3246 -73116 -3186 -72392
rect -3094 -72150 -3034 -72144
rect -2780 -72166 -2320 -72106
rect -2260 -72166 -1238 -72106
rect -2840 -72172 -2780 -72166
rect -3094 -72882 -3034 -72210
rect -2584 -72276 -2578 -72216
rect -2518 -72276 -2512 -72216
rect -2578 -72856 -2518 -72276
rect -3103 -72942 -3094 -72882
rect -3034 -72942 -3025 -72882
rect -2578 -72922 -2518 -72916
rect -2320 -72896 -2260 -72166
rect -1238 -72175 -1178 -72166
rect 506 -72522 566 -71358
rect 1034 -71364 1094 -71358
rect 1808 -71364 1868 -71358
rect 4506 -71358 5034 -71298
rect 5094 -71358 5808 -71298
rect 1292 -71994 1352 -71988
rect 1548 -71994 1608 -71988
rect -236 -72640 -230 -72580
rect -170 -72640 -164 -72580
rect 86 -72582 92 -72522
rect 152 -72582 566 -72522
rect -3094 -73004 -3034 -72942
rect -2320 -72962 -2260 -72956
rect -2058 -73004 -1998 -72998
rect -1648 -73004 -1588 -72998
rect -3034 -73064 -2058 -73004
rect -1998 -73064 -1648 -73004
rect -3094 -73070 -3034 -73064
rect -2058 -73070 -1998 -73064
rect -1648 -73070 -1588 -73064
rect -2962 -73116 -2902 -73110
rect -2186 -73116 -2126 -73110
rect -3186 -73176 -2962 -73116
rect -2902 -73176 -2186 -73116
rect -3246 -73182 -3186 -73176
rect -2962 -73182 -2902 -73176
rect -2186 -73182 -2126 -73176
rect -3092 -73852 -3032 -73846
rect -2574 -73852 -2514 -73846
rect -2058 -73852 -1998 -73846
rect -3032 -73912 -2574 -73852
rect -2514 -73912 -2058 -73852
rect -3092 -73918 -3032 -73912
rect -2574 -73918 -2514 -73912
rect -2058 -73918 -1998 -73912
rect -2962 -73966 -2902 -73960
rect -2704 -73966 -2644 -73960
rect -2446 -73966 -2386 -73960
rect -2188 -73966 -2128 -73960
rect -3494 -74026 -2962 -73966
rect -2902 -74026 -2704 -73966
rect -2644 -74026 -2446 -73966
rect -2386 -74026 -2188 -73966
rect -2962 -74032 -2902 -74026
rect -2704 -74032 -2644 -74026
rect -2446 -74032 -2386 -74026
rect -2188 -74032 -2128 -74026
rect -230 -74096 -170 -72640
rect 506 -73966 566 -72582
rect 754 -72054 1292 -71994
rect 1352 -72054 1548 -71994
rect 754 -73116 814 -72054
rect 1292 -72060 1352 -72054
rect 1548 -72060 1608 -72054
rect 1160 -72106 1220 -72100
rect 1680 -72106 1740 -72100
rect 2762 -72106 2822 -72097
rect 906 -72150 966 -72144
rect 1220 -72166 1680 -72106
rect 1740 -72166 2762 -72106
rect 1160 -72172 1220 -72166
rect 906 -72882 966 -72210
rect 1416 -72276 1422 -72216
rect 1482 -72276 1488 -72216
rect 1422 -72856 1482 -72276
rect 897 -72942 906 -72882
rect 966 -72942 975 -72882
rect 1422 -72922 1482 -72916
rect 1680 -72896 1740 -72166
rect 2762 -72175 2822 -72166
rect 4506 -72522 4566 -71358
rect 5034 -71364 5094 -71358
rect 5808 -71364 5868 -71358
rect 5292 -71994 5352 -71988
rect 5548 -71994 5608 -71988
rect 3764 -72640 3770 -72580
rect 3830 -72640 3836 -72580
rect 4086 -72582 4092 -72522
rect 4152 -72582 4566 -72522
rect 906 -73004 966 -72942
rect 1680 -72962 1740 -72956
rect 1942 -73004 2002 -72998
rect 2352 -73004 2412 -72998
rect 966 -73064 1942 -73004
rect 2002 -73064 2352 -73004
rect 906 -73070 966 -73064
rect 1942 -73070 2002 -73064
rect 2352 -73070 2412 -73064
rect 1038 -73116 1098 -73110
rect 1814 -73116 1874 -73110
rect 814 -73176 1038 -73116
rect 1098 -73176 1814 -73116
rect 754 -73182 814 -73176
rect 1038 -73182 1098 -73176
rect 1814 -73182 1874 -73176
rect 908 -73852 968 -73846
rect 1426 -73852 1486 -73846
rect 1942 -73852 2002 -73846
rect 968 -73912 1426 -73852
rect 1486 -73912 1942 -73852
rect 908 -73918 968 -73912
rect 1426 -73918 1486 -73912
rect 1942 -73918 2002 -73912
rect 1038 -73966 1098 -73960
rect 1296 -73966 1356 -73960
rect 1554 -73966 1614 -73960
rect 1812 -73966 1872 -73960
rect 506 -74026 1038 -73966
rect 1098 -74026 1296 -73966
rect 1356 -74026 1554 -73966
rect 1614 -74026 1812 -73966
rect 1038 -74032 1098 -74026
rect 1296 -74032 1356 -74026
rect 1554 -74032 1614 -74026
rect 1812 -74032 1872 -74026
rect 3770 -74096 3830 -72640
rect 4506 -73966 4566 -72582
rect 4754 -72054 5292 -71994
rect 5352 -72054 5548 -71994
rect 4754 -73116 4814 -72054
rect 5292 -72060 5352 -72054
rect 5548 -72060 5608 -72054
rect 5160 -72106 5220 -72100
rect 5680 -72106 5740 -72100
rect 6762 -72106 6822 -72097
rect 4906 -72150 4966 -72144
rect 5220 -72166 5680 -72106
rect 5740 -72166 6762 -72106
rect 5160 -72172 5220 -72166
rect 4906 -72882 4966 -72210
rect 5416 -72276 5422 -72216
rect 5482 -72276 5488 -72216
rect 5422 -72856 5482 -72276
rect 4897 -72942 4906 -72882
rect 4966 -72942 4975 -72882
rect 5422 -72922 5482 -72916
rect 5680 -72896 5740 -72166
rect 6762 -72175 6822 -72166
rect 4906 -73004 4966 -72942
rect 5680 -72962 5740 -72956
rect 5942 -73004 6002 -72998
rect 6352 -73004 6412 -72998
rect 4966 -73064 5942 -73004
rect 6002 -73064 6352 -73004
rect 4906 -73070 4966 -73064
rect 5942 -73070 6002 -73064
rect 6352 -73070 6412 -73064
rect 5038 -73116 5098 -73110
rect 5814 -73116 5874 -73110
rect 4814 -73176 5038 -73116
rect 5098 -73176 5814 -73116
rect 4754 -73182 4814 -73176
rect 5038 -73182 5098 -73176
rect 5814 -73182 5874 -73176
rect 4908 -73852 4968 -73846
rect 5426 -73852 5486 -73846
rect 5942 -73852 6002 -73846
rect 4968 -73912 5426 -73852
rect 5486 -73912 5942 -73852
rect 4908 -73918 4968 -73912
rect 5426 -73918 5486 -73912
rect 5942 -73918 6002 -73912
rect 5038 -73966 5098 -73960
rect 5296 -73966 5356 -73960
rect 5554 -73966 5614 -73960
rect 5812 -73966 5872 -73960
rect 4506 -74026 5038 -73966
rect 5098 -74026 5296 -73966
rect 5356 -74026 5554 -73966
rect 5614 -74026 5812 -73966
rect 5038 -74032 5098 -74026
rect 5296 -74032 5356 -74026
rect 5554 -74032 5614 -74026
rect 5812 -74032 5872 -74026
rect -28230 -74156 -27496 -74096
rect -27436 -74156 -27430 -74096
rect -24230 -74156 -23496 -74096
rect -23436 -74156 -23430 -74096
rect -20230 -74156 -19496 -74096
rect -19436 -74156 -19430 -74096
rect -16230 -74156 -15496 -74096
rect -15436 -74156 -15430 -74096
rect -12230 -74156 -11496 -74096
rect -11436 -74156 -11430 -74096
rect -8230 -74156 -7496 -74096
rect -7436 -74156 -7430 -74096
rect -4230 -74156 -3496 -74096
rect -3436 -74156 -3430 -74096
rect -230 -74156 504 -74096
rect 564 -74156 570 -74096
rect 3770 -74156 4504 -74096
rect 4564 -74156 4570 -74096
rect -27496 -74690 -27436 -74684
rect -26706 -74690 -26646 -74684
rect -26450 -74690 -26390 -74684
rect -27436 -74750 -26706 -74690
rect -26646 -74750 -26450 -74690
rect -27496 -74756 -27436 -74750
rect -26706 -74756 -26646 -74750
rect -26450 -74756 -26390 -74750
rect -23496 -74690 -23436 -74684
rect -22706 -74690 -22646 -74684
rect -22450 -74690 -22390 -74684
rect -23436 -74750 -22706 -74690
rect -22646 -74750 -22450 -74690
rect -23496 -74756 -23436 -74750
rect -22706 -74756 -22646 -74750
rect -22450 -74756 -22390 -74750
rect -19496 -74690 -19436 -74684
rect -18706 -74690 -18646 -74684
rect -18450 -74690 -18390 -74684
rect -19436 -74750 -18706 -74690
rect -18646 -74750 -18450 -74690
rect -19496 -74756 -19436 -74750
rect -18706 -74756 -18646 -74750
rect -18450 -74756 -18390 -74750
rect -15496 -74690 -15436 -74684
rect -14706 -74690 -14646 -74684
rect -14450 -74690 -14390 -74684
rect -15436 -74750 -14706 -74690
rect -14646 -74750 -14450 -74690
rect -15496 -74756 -15436 -74750
rect -14706 -74756 -14646 -74750
rect -14450 -74756 -14390 -74750
rect -11496 -74690 -11436 -74684
rect -10706 -74690 -10646 -74684
rect -10450 -74690 -10390 -74684
rect -11436 -74750 -10706 -74690
rect -10646 -74750 -10450 -74690
rect -11496 -74756 -11436 -74750
rect -10706 -74756 -10646 -74750
rect -10450 -74756 -10390 -74750
rect -7496 -74690 -7436 -74684
rect -6706 -74690 -6646 -74684
rect -6450 -74690 -6390 -74684
rect -7436 -74750 -6706 -74690
rect -6646 -74750 -6450 -74690
rect -7496 -74756 -7436 -74750
rect -6706 -74756 -6646 -74750
rect -6450 -74756 -6390 -74750
rect -3496 -74690 -3436 -74684
rect -2706 -74690 -2646 -74684
rect -2450 -74690 -2390 -74684
rect -3436 -74750 -2706 -74690
rect -2646 -74750 -2450 -74690
rect -3496 -74756 -3436 -74750
rect -2706 -74756 -2646 -74750
rect -2450 -74756 -2390 -74750
rect 504 -74690 564 -74684
rect 1294 -74690 1354 -74684
rect 1550 -74690 1610 -74684
rect 564 -74750 1294 -74690
rect 1354 -74750 1550 -74690
rect 504 -74756 564 -74750
rect 1294 -74756 1354 -74750
rect 1550 -74756 1610 -74750
rect 4504 -74690 4564 -74684
rect 5294 -74690 5354 -74684
rect 5550 -74690 5610 -74684
rect 4564 -74750 5294 -74690
rect 5354 -74750 5550 -74690
rect 4504 -74756 4564 -74750
rect 5294 -74756 5354 -74750
rect 5550 -74756 5610 -74750
rect -26578 -74810 -26518 -74804
rect -25648 -74810 -25588 -74804
rect -27092 -74870 -27032 -74864
rect -26518 -74870 -25648 -74810
rect -22578 -74810 -22518 -74804
rect -21648 -74810 -21588 -74804
rect -23092 -74868 -23032 -74862
rect -27101 -74930 -27092 -74870
rect -27032 -74930 -27023 -74870
rect -26578 -74876 -26518 -74870
rect -25648 -74876 -25588 -74870
rect -26834 -74922 -26774 -74916
rect -26316 -74922 -26256 -74916
rect -27092 -74936 -27032 -74930
rect -26774 -74982 -26316 -74922
rect -23101 -74928 -23092 -74868
rect -23032 -74928 -23023 -74868
rect -22518 -74870 -21648 -74810
rect -18578 -74810 -18518 -74804
rect -17648 -74810 -17588 -74804
rect -19092 -74868 -19032 -74862
rect -22578 -74876 -22518 -74870
rect -21648 -74876 -21588 -74870
rect -22834 -74922 -22774 -74916
rect -22316 -74922 -22256 -74916
rect -23092 -74934 -23032 -74928
rect -26834 -74988 -26774 -74982
rect -26316 -74988 -26256 -74982
rect -22774 -74982 -22316 -74922
rect -19101 -74928 -19092 -74868
rect -19032 -74928 -19023 -74868
rect -18518 -74870 -17648 -74810
rect -14578 -74810 -14518 -74804
rect -13648 -74810 -13588 -74804
rect -15092 -74868 -15032 -74862
rect -18578 -74876 -18518 -74870
rect -17648 -74876 -17588 -74870
rect -18834 -74922 -18774 -74916
rect -18316 -74922 -18256 -74916
rect -19092 -74934 -19032 -74928
rect -22834 -74988 -22774 -74982
rect -22316 -74988 -22256 -74982
rect -18774 -74982 -18316 -74922
rect -15101 -74928 -15092 -74868
rect -15032 -74928 -15023 -74868
rect -14518 -74870 -13648 -74810
rect -10578 -74810 -10518 -74804
rect -9648 -74810 -9588 -74804
rect -11092 -74870 -11032 -74864
rect -10518 -74870 -9648 -74810
rect -6578 -74810 -6518 -74804
rect -5648 -74810 -5588 -74804
rect -7092 -74870 -7032 -74864
rect -6518 -74870 -5648 -74810
rect -2578 -74810 -2518 -74804
rect -1648 -74810 -1588 -74804
rect -3092 -74868 -3032 -74862
rect -14578 -74876 -14518 -74870
rect -13648 -74876 -13588 -74870
rect -14834 -74922 -14774 -74916
rect -14316 -74922 -14256 -74916
rect -15092 -74934 -15032 -74928
rect -18834 -74988 -18774 -74982
rect -18316 -74988 -18256 -74982
rect -14774 -74982 -14316 -74922
rect -11101 -74930 -11092 -74870
rect -11032 -74930 -11023 -74870
rect -10578 -74876 -10518 -74870
rect -9648 -74876 -9588 -74870
rect -10834 -74922 -10774 -74916
rect -10316 -74922 -10256 -74916
rect -11092 -74936 -11032 -74930
rect -14834 -74988 -14774 -74982
rect -14316 -74988 -14256 -74982
rect -10774 -74982 -10316 -74922
rect -7101 -74930 -7092 -74870
rect -7032 -74930 -7023 -74870
rect -6578 -74876 -6518 -74870
rect -5648 -74876 -5588 -74870
rect -6834 -74922 -6774 -74916
rect -6316 -74922 -6256 -74916
rect -7092 -74936 -7032 -74930
rect -10834 -74988 -10774 -74982
rect -10316 -74988 -10256 -74982
rect -6774 -74982 -6316 -74922
rect -3101 -74928 -3092 -74868
rect -3032 -74928 -3023 -74868
rect -2518 -74870 -1648 -74810
rect 1422 -74810 1482 -74804
rect 2352 -74810 2412 -74804
rect 908 -74868 968 -74862
rect -2578 -74876 -2518 -74870
rect -1648 -74876 -1588 -74870
rect -2834 -74922 -2774 -74916
rect -2316 -74922 -2256 -74916
rect -3092 -74934 -3032 -74928
rect -6834 -74988 -6774 -74982
rect -6316 -74988 -6256 -74982
rect -2774 -74982 -2316 -74922
rect 899 -74928 908 -74868
rect 968 -74928 977 -74868
rect 1482 -74870 2352 -74810
rect 5422 -74810 5482 -74804
rect 6352 -74810 6412 -74804
rect 4908 -74866 4968 -74860
rect 1422 -74876 1482 -74870
rect 2352 -74876 2412 -74870
rect 1166 -74922 1226 -74916
rect 1684 -74922 1744 -74916
rect 908 -74934 968 -74928
rect -2834 -74988 -2774 -74982
rect -2316 -74988 -2256 -74982
rect 1226 -74982 1684 -74922
rect 4899 -74926 4908 -74866
rect 4968 -74926 4977 -74866
rect 5482 -74870 6352 -74810
rect 5422 -74876 5482 -74870
rect 6352 -74876 6412 -74870
rect 5166 -74922 5226 -74916
rect 5684 -74922 5744 -74916
rect 4908 -74932 4968 -74926
rect 1166 -74988 1226 -74982
rect 1684 -74988 1744 -74982
rect 5226 -74982 5684 -74922
rect 5166 -74988 5226 -74982
rect 5684 -74988 5744 -74982
rect -27422 -75096 -25520 -75066
rect -27422 -75160 -27388 -75096
rect -25564 -75160 -25520 -75096
rect -27422 -75190 -25520 -75160
rect -23422 -75096 -21520 -75066
rect -23422 -75160 -23388 -75096
rect -21564 -75160 -21520 -75096
rect -23422 -75190 -21520 -75160
rect -19422 -75096 -17520 -75066
rect -19422 -75160 -19388 -75096
rect -17564 -75160 -17520 -75096
rect -19422 -75190 -17520 -75160
rect -15422 -75096 -13520 -75066
rect -15422 -75160 -15388 -75096
rect -13564 -75160 -13520 -75096
rect -15422 -75190 -13520 -75160
rect -11422 -75096 -9520 -75066
rect -11422 -75160 -11388 -75096
rect -9564 -75160 -9520 -75096
rect -11422 -75190 -9520 -75160
rect -7422 -75096 -5520 -75066
rect -7422 -75160 -7388 -75096
rect -5564 -75160 -5520 -75096
rect -7422 -75190 -5520 -75160
rect -3422 -75096 -1520 -75066
rect -3422 -75160 -3388 -75096
rect -1564 -75160 -1520 -75096
rect -3422 -75190 -1520 -75160
rect 578 -75096 2480 -75066
rect 578 -75160 612 -75096
rect 2436 -75160 2480 -75096
rect 578 -75190 2480 -75160
rect 4578 -75096 6480 -75066
rect 4578 -75160 4612 -75096
rect 6436 -75160 6480 -75096
rect 4578 -75190 6480 -75160
rect -27578 -75364 -26978 -75354
rect -27578 -75674 -26978 -75664
rect -26066 -75364 -25466 -75354
rect -26066 -75674 -25466 -75664
rect -23578 -75364 -22978 -75354
rect -23578 -75674 -22978 -75664
rect -22066 -75364 -21466 -75354
rect -22066 -75674 -21466 -75664
rect -19578 -75364 -18978 -75354
rect -19578 -75674 -18978 -75664
rect -18066 -75364 -17466 -75354
rect -18066 -75674 -17466 -75664
rect -15578 -75364 -14978 -75354
rect -15578 -75674 -14978 -75664
rect -14066 -75364 -13466 -75354
rect -14066 -75674 -13466 -75664
rect -11578 -75364 -10978 -75354
rect -11578 -75674 -10978 -75664
rect -10066 -75364 -9466 -75354
rect -10066 -75674 -9466 -75664
rect -7578 -75364 -6978 -75354
rect -7578 -75674 -6978 -75664
rect -6066 -75364 -5466 -75354
rect -6066 -75674 -5466 -75664
rect -3578 -75364 -2978 -75354
rect -3578 -75674 -2978 -75664
rect -2066 -75364 -1466 -75354
rect -2066 -75674 -1466 -75664
rect 422 -75364 1022 -75354
rect 422 -75674 1022 -75664
rect 1934 -75364 2534 -75354
rect 1934 -75674 2534 -75664
rect 4422 -75364 5022 -75354
rect 4422 -75674 5022 -75664
rect 5934 -75364 6534 -75354
rect 5934 -75674 6534 -75664
<< via2 >>
rect 25928 -28062 26528 -27762
rect 49560 -28062 50160 -27762
rect 29505 -28358 46290 -28144
rect -14318 -40874 -14218 -40774
rect -7399 -40947 -7309 -40857
rect -15855 -41219 -15765 -41129
rect -13168 -41194 -13068 -41094
rect -7973 -41189 -7883 -41099
rect -5310 -41246 -5210 -41146
rect -14627 -42559 -14537 -42469
rect -6427 -42627 -6337 -42537
rect -11643 -42931 -11553 -42841
rect -9531 -42931 -9441 -42841
rect -13746 -43220 -13646 -43120
rect -7442 -43212 -7342 -43112
rect -10917 -44927 -10827 -44837
rect -10164 -45224 -10064 -45124
rect -13741 -46931 -13651 -46841
rect -7444 -46858 -7344 -46758
rect -11644 -47234 -11544 -47134
rect -9537 -47199 -9447 -47109
rect -14632 -47524 -14532 -47424
rect 11814 -42648 22576 -42356
rect 26986 -43002 27046 -42942
rect 27763 -43017 27853 -42927
rect 49191 -41181 49281 -41091
rect -6432 -47630 -6332 -47530
rect -15855 -48947 -15765 -48857
rect -12999 -48945 -12909 -48855
rect -8060 -48950 -7960 -48850
rect -5312 -48878 -5212 -48778
rect -7431 -49141 -7341 -49051
rect -13756 -49248 -13656 -49148
rect 52262 -39386 55130 -39086
rect 56534 -39386 58154 -39086
rect 57474 -40536 57534 -40476
rect 51918 -41166 51978 -41106
rect 52380 -42022 52440 -41962
rect 53314 -42542 53374 -42482
rect 54200 -42548 54260 -42476
rect 55295 -42553 55365 -42471
rect 56047 -42667 56137 -42577
rect 57951 -42669 58041 -42579
rect 55824 -43584 58268 -43278
rect 14775 -52000 14865 -51987
rect 14775 -52060 14782 -52000
rect 14782 -52060 14842 -52000
rect 14842 -52060 14865 -52000
rect 14775 -52077 14865 -52060
rect 14767 -53043 14857 -52953
rect 14769 -54037 14859 -53947
rect 14769 -55043 14859 -54953
rect 14779 -56358 14869 -56339
rect 14779 -56418 14782 -56358
rect 14782 -56418 14842 -56358
rect 14842 -56418 14869 -56358
rect 14779 -56429 14869 -56418
rect 9372 -57518 9436 -56724
rect 12524 -57592 12584 -57532
rect 10652 -57695 10654 -57635
rect 10654 -57695 10712 -57635
rect 12526 -58243 12586 -58183
rect 10294 -58514 12110 -58408
rect 17372 -58608 49372 -58454
rect 13228 -59094 13828 -58794
rect 49660 -59094 50260 -58794
rect 13016 -59774 13076 -59714
rect -9198 -64086 -9138 -64026
rect -27578 -64832 -26978 -64532
rect -26066 -64832 -25466 -64532
rect -23578 -64832 -22978 -64532
rect -22066 -64832 -21466 -64532
rect -19578 -64832 -18978 -64532
rect -18066 -64832 -17466 -64532
rect -15578 -64832 -14978 -64532
rect -14066 -64832 -13466 -64532
rect -11578 -64832 -10978 -64532
rect -10066 -64832 -9466 -64532
rect -27388 -65100 -25564 -65036
rect -23388 -65100 -21564 -65036
rect -19388 -65100 -17564 -65036
rect -15388 -65100 -13564 -65036
rect -11388 -65100 -9564 -65036
rect -25195 -65285 -25105 -65195
rect -21031 -65287 -20941 -65197
rect -17109 -65287 -17019 -65197
rect -16087 -65287 -15997 -65197
rect -7578 -64832 -6978 -64532
rect -6066 -64832 -5466 -64532
rect -3578 -64832 -2978 -64532
rect -2066 -64832 -1466 -64532
rect 422 -64832 1022 -64532
rect 1934 -64832 2534 -64532
rect 4422 -64832 5022 -64532
rect 5934 -64832 6534 -64532
rect -7388 -65100 -5564 -65036
rect -3388 -65100 -1564 -65036
rect 612 -65100 2436 -65036
rect 4612 -65100 6436 -65036
rect -7956 -65274 -7896 -65214
rect -4097 -65287 -4007 -65197
rect -39 -65291 51 -65201
rect 4015 -65289 4105 -65199
rect -26448 -65506 -26390 -65446
rect -26390 -65506 -26388 -65446
rect -22448 -65506 -22390 -65446
rect -22390 -65506 -22388 -65446
rect -18450 -65506 -18390 -65446
rect -14450 -65506 -14390 -65446
rect -10450 -65506 -10390 -65446
rect -6448 -65506 -6390 -65446
rect -6390 -65506 -6388 -65446
rect -2452 -65506 -2450 -65446
rect -2450 -65506 -2392 -65446
rect 1552 -65506 1610 -65446
rect 1610 -65506 1612 -65446
rect 5554 -65506 5610 -65446
rect 5610 -65506 5614 -65446
rect -26578 -67980 -26518 -67920
rect -22578 -67980 -22518 -67920
rect -18578 -67980 -18518 -67920
rect -14578 -67980 -14518 -67920
rect -10578 -67980 -10518 -67920
rect -6578 -67980 -6518 -67920
rect -2578 -67980 -2518 -67920
rect 1422 -67980 1482 -67920
rect 5422 -67980 5482 -67922
rect 5422 -67982 5482 -67980
rect -25232 -69012 -25172 -68952
rect -21232 -69012 -21172 -68952
rect -17232 -69012 -17172 -68952
rect -13232 -69012 -13172 -68952
rect -9232 -69012 -9172 -68952
rect -5232 -69012 -5172 -68952
rect -1232 -69012 -1172 -68952
rect 2768 -69012 2828 -68952
rect 6768 -69012 6828 -68952
rect -27430 -69222 -25722 -69154
rect -23430 -69222 -21722 -69154
rect -19430 -69222 -17722 -69154
rect -15430 -69222 -13722 -69154
rect -11430 -69222 -9722 -69154
rect -7430 -69222 -5722 -69154
rect -3430 -69222 -1722 -69154
rect 570 -69222 2278 -69154
rect 4570 -69222 6278 -69154
rect -27578 -69704 -26978 -69404
rect -26066 -69704 -25466 -69404
rect -23578 -69704 -22978 -69404
rect -22066 -69704 -21466 -69404
rect -19578 -69704 -18978 -69404
rect -18066 -69704 -17466 -69404
rect -15578 -69704 -14978 -69404
rect -14066 -69704 -13466 -69404
rect -11578 -69704 -10978 -69404
rect -10066 -69704 -9466 -69404
rect -7578 -69704 -6978 -69404
rect -6066 -69704 -5466 -69404
rect -3578 -69704 -2978 -69404
rect -2066 -69704 -1466 -69404
rect 422 -69704 1022 -69404
rect 1934 -69704 2534 -69404
rect 4422 -69704 5022 -69404
rect 5934 -69704 6534 -69404
rect -27578 -70792 -26978 -70492
rect -26066 -70792 -25466 -70492
rect -23578 -70792 -22978 -70492
rect -22066 -70792 -21466 -70492
rect -19578 -70792 -18978 -70492
rect -18066 -70792 -17466 -70492
rect -15578 -70792 -14978 -70492
rect -14066 -70792 -13466 -70492
rect -11578 -70792 -10978 -70492
rect -10066 -70792 -9466 -70492
rect -7578 -70792 -6978 -70492
rect -6066 -70792 -5466 -70492
rect -3578 -70792 -2978 -70492
rect -2066 -70792 -1466 -70492
rect 422 -70792 1022 -70492
rect 1934 -70792 2534 -70492
rect 4422 -70792 5022 -70492
rect 5934 -70792 6534 -70492
rect -27430 -71042 -25722 -70974
rect -23430 -71042 -21722 -70974
rect -19430 -71042 -17722 -70974
rect -15430 -71042 -13722 -70974
rect -11430 -71042 -9722 -70974
rect -7430 -71042 -5722 -70974
rect -3430 -71042 -1722 -70974
rect 570 -71042 2278 -70974
rect 4570 -71042 6278 -70974
rect -25238 -72166 -25178 -72106
rect -27094 -72942 -27034 -72882
rect -21238 -72166 -21178 -72106
rect -23094 -72942 -23034 -72882
rect -17238 -72166 -17178 -72106
rect -19094 -72942 -19034 -72882
rect -13238 -72166 -13178 -72106
rect -15094 -72942 -15034 -72882
rect -9238 -72166 -9178 -72106
rect -11094 -72940 -11034 -72880
rect -5238 -72166 -5178 -72106
rect -7094 -72942 -7034 -72882
rect -1238 -72166 -1178 -72106
rect -3094 -72942 -3034 -72882
rect 2762 -72166 2822 -72106
rect 906 -72942 966 -72882
rect 6762 -72166 6822 -72106
rect 4906 -72942 4966 -72882
rect -27092 -74930 -27032 -74870
rect -23092 -74928 -23032 -74868
rect -19092 -74928 -19032 -74868
rect -15092 -74928 -15032 -74868
rect -11092 -74930 -11032 -74870
rect -7092 -74930 -7032 -74870
rect -3092 -74928 -3032 -74868
rect 908 -74928 968 -74868
rect 4908 -74926 4968 -74866
rect -27388 -75160 -25564 -75096
rect -23388 -75160 -21564 -75096
rect -19388 -75160 -17564 -75096
rect -15388 -75160 -13564 -75096
rect -11388 -75160 -9564 -75096
rect -7388 -75160 -5564 -75096
rect -3388 -75160 -1564 -75096
rect 612 -75160 2436 -75096
rect 4612 -75160 6436 -75096
rect -27578 -75664 -26978 -75364
rect -26066 -75664 -25466 -75364
rect -23578 -75664 -22978 -75364
rect -22066 -75664 -21466 -75364
rect -19578 -75664 -18978 -75364
rect -18066 -75664 -17466 -75364
rect -15578 -75664 -14978 -75364
rect -14066 -75664 -13466 -75364
rect -11578 -75664 -10978 -75364
rect -10066 -75664 -9466 -75364
rect -7578 -75664 -6978 -75364
rect -6066 -75664 -5466 -75364
rect -3578 -75664 -2978 -75364
rect -2066 -75664 -1466 -75364
rect 422 -75664 1022 -75364
rect 1934 -75664 2534 -75364
rect 4422 -75664 5022 -75364
rect 5934 -75664 6534 -75364
<< metal3 >>
rect -29235 -27370 -27536 -27206
rect -29235 -28652 -27620 -27370
rect -27556 -28652 -27536 -27370
rect -29235 -28806 -27536 -28652
rect -27129 -27370 -25430 -27206
rect -27129 -28652 -25514 -27370
rect -25450 -28652 -25430 -27370
rect -27129 -28806 -25430 -28652
rect -25023 -27370 -23324 -27206
rect -25023 -28652 -23408 -27370
rect -23344 -28652 -23324 -27370
rect -25023 -28806 -23324 -28652
rect -22917 -27370 -21218 -27206
rect -22917 -28652 -21302 -27370
rect -21238 -28652 -21218 -27370
rect -22917 -28806 -21218 -28652
rect -20811 -27370 -19112 -27206
rect -20811 -28652 -19196 -27370
rect -19132 -28652 -19112 -27370
rect -20811 -28806 -19112 -28652
rect -18705 -27370 -17006 -27206
rect -18705 -28652 -17090 -27370
rect -17026 -28652 -17006 -27370
rect -18705 -28806 -17006 -28652
rect -16599 -27370 -14900 -27206
rect -16599 -28652 -14984 -27370
rect -14920 -28652 -14900 -27370
rect -16599 -28806 -14900 -28652
rect -14493 -27370 -12794 -27206
rect -14493 -28652 -12878 -27370
rect -12814 -28652 -12794 -27370
rect -14493 -28806 -12794 -28652
rect -12387 -27370 -10688 -27206
rect -12387 -28652 -10772 -27370
rect -10708 -28652 -10688 -27370
rect -12387 -28806 -10688 -28652
rect -10281 -27370 -8582 -27206
rect -10281 -28652 -8666 -27370
rect -8602 -28652 -8582 -27370
rect -10281 -28806 -8582 -28652
rect -8175 -27370 -6476 -27206
rect -8175 -28652 -6560 -27370
rect -6496 -28652 -6476 -27370
rect -8175 -28806 -6476 -28652
rect -6069 -27370 -4370 -27206
rect -6069 -28652 -4454 -27370
rect -4390 -28652 -4370 -27370
rect -6069 -28806 -4370 -28652
rect -3963 -27370 -2264 -27206
rect -3963 -28652 -2348 -27370
rect -2284 -28652 -2264 -27370
rect -3963 -28806 -2264 -28652
rect -1857 -27370 -158 -27206
rect -1857 -28652 -242 -27370
rect -178 -28652 -158 -27370
rect -1857 -28806 -158 -28652
rect 249 -27370 1948 -27206
rect 249 -28652 1864 -27370
rect 1928 -28652 1948 -27370
rect 249 -28806 1948 -28652
rect 2355 -27370 4054 -27206
rect 2355 -28652 3970 -27370
rect 4034 -28652 4054 -27370
rect 2355 -28806 4054 -28652
rect 4461 -27370 6160 -27206
rect 4461 -28652 6076 -27370
rect 6140 -28652 6160 -27370
rect 4461 -28806 6160 -28652
rect 6567 -27370 8266 -27206
rect 6567 -28652 8182 -27370
rect 8246 -28652 8266 -27370
rect 25918 -27762 26538 -27757
rect 25918 -28062 25928 -27762
rect 26528 -28062 26538 -27762
rect 25918 -28067 26538 -28062
rect 49550 -27762 50170 -27757
rect 49550 -28062 49560 -27762
rect 50160 -28062 50170 -27762
rect 49550 -28067 50170 -28062
rect 29442 -28144 46322 -28112
rect 29442 -28358 29505 -28144
rect 46290 -28358 46322 -28144
rect 29442 -28378 46322 -28358
rect 29442 -28380 33796 -28378
rect 6567 -28806 8266 -28652
rect 10276 -29038 25316 -28892
rect 10276 -29048 24470 -29038
rect -29235 -29370 -27536 -29206
rect -29235 -30652 -27620 -29370
rect -27556 -30652 -27536 -29370
rect -29235 -30806 -27536 -30652
rect -27129 -29370 -25430 -29206
rect -27129 -30652 -25514 -29370
rect -25450 -29944 -25430 -29370
rect -25023 -29370 -23324 -29206
rect -25023 -29944 -23408 -29370
rect -25450 -30044 -23408 -29944
rect -25450 -30652 -25430 -30044
rect -27129 -30806 -25430 -30652
rect -25023 -30652 -23408 -30044
rect -23344 -29944 -23324 -29370
rect -22917 -29370 -21218 -29206
rect -22917 -29944 -21302 -29370
rect -23344 -30044 -21302 -29944
rect -23344 -30652 -23324 -30044
rect -25023 -30806 -23324 -30652
rect -22917 -30652 -21302 -30044
rect -21238 -29944 -21218 -29370
rect -20811 -29370 -19112 -29206
rect -20811 -29944 -19196 -29370
rect -21238 -30044 -19196 -29944
rect -21238 -30652 -21218 -30044
rect -22917 -30806 -21218 -30652
rect -20811 -30652 -19196 -30044
rect -19132 -29944 -19112 -29370
rect -18705 -29370 -17006 -29206
rect -18705 -29944 -17090 -29370
rect -19132 -30044 -17090 -29944
rect -19132 -30652 -19112 -30044
rect -20811 -30806 -19112 -30652
rect -18705 -30652 -17090 -30044
rect -17026 -29944 -17006 -29370
rect -16599 -29370 -14900 -29206
rect -16599 -29944 -14984 -29370
rect -17026 -30044 -14984 -29944
rect -17026 -30652 -17006 -30044
rect -18705 -30806 -17006 -30652
rect -16599 -30652 -14984 -30044
rect -14920 -29944 -14900 -29370
rect -14493 -29370 -12794 -29206
rect -14493 -29944 -12878 -29370
rect -14920 -30044 -12878 -29944
rect -14920 -30652 -14900 -30044
rect -16599 -30806 -14900 -30652
rect -14493 -30652 -12878 -30044
rect -12814 -29944 -12794 -29370
rect -12387 -29370 -10688 -29206
rect -12387 -29944 -10772 -29370
rect -12814 -30044 -10772 -29944
rect -12814 -30652 -12794 -30044
rect -14493 -30806 -12794 -30652
rect -12387 -30652 -10772 -30044
rect -10708 -29944 -10688 -29370
rect -10281 -29370 -8582 -29206
rect -10281 -29944 -8666 -29370
rect -10708 -30044 -8666 -29944
rect -10708 -30652 -10688 -30044
rect -12387 -30806 -10688 -30652
rect -10281 -30652 -8666 -30044
rect -8602 -29944 -8582 -29370
rect -8175 -29370 -6476 -29206
rect -8175 -29944 -6560 -29370
rect -8602 -30044 -6560 -29944
rect -8602 -30652 -8582 -30044
rect -10281 -30806 -8582 -30652
rect -8175 -30652 -6560 -30044
rect -6496 -29944 -6476 -29370
rect -6069 -29370 -4370 -29206
rect -6069 -29944 -4454 -29370
rect -6496 -30044 -4454 -29944
rect -6496 -30652 -6476 -30044
rect -8175 -30806 -6476 -30652
rect -6069 -30652 -4454 -30044
rect -4390 -29944 -4370 -29370
rect -3963 -29370 -2264 -29206
rect -3963 -29944 -2348 -29370
rect -4390 -30044 -2348 -29944
rect -4390 -30652 -4370 -30044
rect -6069 -30806 -4370 -30652
rect -3963 -30652 -2348 -30044
rect -2284 -29944 -2264 -29370
rect -1857 -29370 -158 -29206
rect -1857 -29944 -242 -29370
rect -2284 -30044 -242 -29944
rect -2284 -30652 -2264 -30044
rect -3963 -30806 -2264 -30652
rect -1857 -30652 -242 -30044
rect -178 -29944 -158 -29370
rect 249 -29370 1948 -29206
rect 249 -29944 1864 -29370
rect -178 -30044 1864 -29944
rect -178 -30652 -158 -30044
rect -1857 -30806 -158 -30652
rect 249 -30652 1864 -30044
rect 1928 -29944 1948 -29370
rect 2355 -29370 4054 -29206
rect 2355 -29944 3970 -29370
rect 1928 -30044 3970 -29944
rect 1928 -30652 1948 -30044
rect 249 -30806 1948 -30652
rect 2355 -30652 3970 -30044
rect 4034 -29944 4054 -29370
rect 4461 -29370 6160 -29206
rect 4461 -29944 6076 -29370
rect 4034 -30044 6076 -29944
rect 4034 -30652 4054 -30044
rect 2355 -30806 4054 -30652
rect 4461 -30652 6076 -30044
rect 6140 -30652 6160 -29370
rect 4461 -30806 6160 -30652
rect 6567 -29370 8266 -29206
rect 6567 -30652 8182 -29370
rect 8246 -30652 8266 -29370
rect 6567 -30806 8266 -30652
rect 10276 -29738 10428 -29048
rect 11124 -29736 24470 -29048
rect 25160 -29736 25316 -29038
rect 11124 -29738 25316 -29736
rect -26392 -31206 -26292 -30806
rect -24286 -31206 -24178 -30806
rect -22172 -31206 -22072 -30806
rect -20066 -31206 -19966 -30806
rect -17960 -31206 -17860 -30806
rect -15854 -31206 -15754 -30806
rect -13748 -31206 -13648 -30806
rect -11642 -31206 -11542 -30806
rect -9536 -31206 -9436 -30806
rect -7430 -31206 -7330 -30806
rect -5324 -31206 -5224 -30806
rect -3218 -31206 -3118 -30806
rect -1112 -31206 -1012 -30806
rect 994 -31206 1094 -30806
rect 3060 -31206 3160 -30806
rect 5228 -31206 5328 -30806
rect -29235 -31370 -27536 -31206
rect -29235 -32652 -27620 -31370
rect -27556 -32652 -27536 -31370
rect -29235 -32806 -27536 -32652
rect -27129 -31370 -25430 -31206
rect -27129 -32652 -25514 -31370
rect -25450 -31934 -25430 -31370
rect -25023 -31370 -23324 -31206
rect -25023 -31934 -23408 -31370
rect -25450 -32034 -23408 -31934
rect -25450 -32652 -25430 -32034
rect -27129 -32806 -25430 -32652
rect -25023 -32652 -23408 -32034
rect -23344 -31934 -23324 -31370
rect -22917 -31370 -21218 -31206
rect -22917 -31934 -21302 -31370
rect -23344 -32034 -21302 -31934
rect -23344 -32652 -23324 -32034
rect -25023 -32806 -23324 -32652
rect -22917 -32652 -21302 -32034
rect -21238 -31934 -21218 -31370
rect -20811 -31370 -19112 -31206
rect -20811 -31934 -19196 -31370
rect -21238 -32034 -19196 -31934
rect -21238 -32652 -21218 -32034
rect -22917 -32806 -21218 -32652
rect -20811 -32652 -19196 -32034
rect -19132 -31934 -19112 -31370
rect -18705 -31370 -17006 -31206
rect -18705 -31934 -17090 -31370
rect -19132 -32034 -17090 -31934
rect -19132 -32652 -19112 -32034
rect -20811 -32806 -19112 -32652
rect -18705 -32652 -17090 -32034
rect -17026 -31934 -17006 -31370
rect -16599 -31370 -14900 -31206
rect -16599 -31934 -14984 -31370
rect -17026 -32034 -14984 -31934
rect -17026 -32652 -17006 -32034
rect -18705 -32806 -17006 -32652
rect -16599 -32652 -14984 -32034
rect -14920 -31934 -14900 -31370
rect -14493 -31370 -12794 -31206
rect -14493 -31934 -12878 -31370
rect -14920 -32034 -12878 -31934
rect -14920 -32652 -14900 -32034
rect -16599 -32806 -14900 -32652
rect -14493 -32652 -12878 -32034
rect -12814 -31934 -12794 -31370
rect -12387 -31370 -10688 -31206
rect -12387 -31934 -10772 -31370
rect -12814 -32034 -10772 -31934
rect -12814 -32652 -12794 -32034
rect -14493 -32806 -12794 -32652
rect -12387 -32652 -10772 -32034
rect -10708 -31934 -10688 -31370
rect -10281 -31370 -8582 -31206
rect -10281 -31934 -8666 -31370
rect -10708 -32034 -8666 -31934
rect -10708 -32652 -10688 -32034
rect -12387 -32806 -10688 -32652
rect -10281 -32652 -8666 -32034
rect -8602 -31934 -8582 -31370
rect -8175 -31370 -6476 -31206
rect -8175 -31934 -6560 -31370
rect -8602 -32034 -6560 -31934
rect -8602 -32652 -8582 -32034
rect -10281 -32806 -8582 -32652
rect -8175 -32652 -6560 -32034
rect -6496 -31934 -6476 -31370
rect -6069 -31370 -4370 -31206
rect -6069 -31934 -4454 -31370
rect -6496 -32034 -4454 -31934
rect -6496 -32652 -6476 -32034
rect -8175 -32806 -6476 -32652
rect -6069 -32652 -4454 -32034
rect -4390 -31934 -4370 -31370
rect -3963 -31370 -2264 -31206
rect -3963 -31934 -2348 -31370
rect -4390 -32034 -2348 -31934
rect -4390 -32652 -4370 -32034
rect -6069 -32806 -4370 -32652
rect -3963 -32652 -2348 -32034
rect -2284 -31934 -2264 -31370
rect -1857 -31370 -158 -31206
rect -1857 -31934 -242 -31370
rect -2284 -32034 -242 -31934
rect -2284 -32652 -2264 -32034
rect -3963 -32806 -2264 -32652
rect -1857 -32652 -242 -32034
rect -178 -31934 -158 -31370
rect 249 -31370 1948 -31206
rect 249 -31934 1864 -31370
rect -178 -32034 1864 -31934
rect -178 -32652 -158 -32034
rect -1857 -32806 -158 -32652
rect 249 -32652 1864 -32034
rect 1928 -31934 1948 -31370
rect 2355 -31370 4054 -31206
rect 2355 -31934 3970 -31370
rect 1928 -32034 3970 -31934
rect 1928 -32652 1948 -32034
rect 249 -32806 1948 -32652
rect 2355 -32652 3970 -32034
rect 4034 -31950 4054 -31370
rect 4461 -31370 6160 -31206
rect 4461 -31950 6076 -31370
rect 4034 -32050 6076 -31950
rect 4034 -32652 4054 -32050
rect 2355 -32806 4054 -32652
rect 4461 -32652 6076 -32050
rect 6140 -32652 6160 -31370
rect 4461 -32806 6160 -32652
rect 6567 -31370 8266 -31206
rect 6567 -32652 8182 -31370
rect 8246 -32652 8266 -31370
rect 6567 -32806 8266 -32652
rect -26392 -33206 -26292 -32806
rect -24286 -33206 -24186 -32806
rect -22134 -33206 -22034 -32806
rect -20036 -33206 -19936 -32806
rect -17892 -33206 -17792 -32806
rect -1134 -33206 -1034 -32806
rect 964 -33206 1064 -32806
rect 3060 -33206 3160 -32806
rect 5228 -33206 5328 -32806
rect -29235 -33370 -27536 -33206
rect -29235 -34652 -27620 -33370
rect -27556 -34652 -27536 -33370
rect -29235 -34806 -27536 -34652
rect -27129 -33370 -25430 -33206
rect -27129 -34652 -25514 -33370
rect -25450 -33956 -25430 -33370
rect -25023 -33370 -23324 -33206
rect -25023 -33956 -23408 -33370
rect -25450 -34056 -23408 -33956
rect -25450 -34652 -25430 -34056
rect -27129 -34806 -25430 -34652
rect -25023 -34652 -23408 -34056
rect -23344 -33956 -23324 -33370
rect -22917 -33370 -21218 -33206
rect -22917 -33956 -21302 -33370
rect -23344 -34056 -21302 -33956
rect -23344 -34652 -23324 -34056
rect -25023 -34806 -23324 -34652
rect -22917 -34652 -21302 -34056
rect -21238 -33956 -21218 -33370
rect -20811 -33370 -19112 -33206
rect -20811 -33956 -19196 -33370
rect -21238 -34056 -19196 -33956
rect -21238 -34652 -21218 -34056
rect -22917 -34806 -21218 -34652
rect -20811 -34652 -19196 -34056
rect -19132 -33956 -19112 -33370
rect -18705 -33370 -17006 -33206
rect -18705 -33956 -17090 -33370
rect -19132 -34056 -17090 -33956
rect -19132 -34652 -19112 -34056
rect -20811 -34806 -19112 -34652
rect -18705 -34652 -17090 -34056
rect -17026 -34652 -17006 -33370
rect -18705 -34806 -17006 -34652
rect -16599 -33370 -14900 -33206
rect -16599 -34652 -14984 -33370
rect -14920 -33920 -14900 -33370
rect -14493 -33370 -12794 -33206
rect -14493 -33920 -12878 -33370
rect -14920 -34020 -12878 -33920
rect -14920 -34652 -14900 -34020
rect -16599 -34806 -14900 -34652
rect -14493 -34652 -12878 -34020
rect -12814 -33920 -12794 -33370
rect -12387 -33370 -10688 -33206
rect -12387 -33920 -10772 -33370
rect -12814 -34020 -10772 -33920
rect -12814 -34652 -12794 -34020
rect -14493 -34806 -12794 -34652
rect -12387 -34652 -10772 -34020
rect -10708 -33920 -10688 -33370
rect -10281 -33370 -8582 -33206
rect -10281 -33920 -8666 -33370
rect -10708 -34020 -8666 -33920
rect -10708 -34652 -10688 -34020
rect -12387 -34806 -10688 -34652
rect -10281 -34652 -8666 -34020
rect -8602 -33920 -8582 -33370
rect -8175 -33370 -6476 -33206
rect -8175 -33920 -6560 -33370
rect -8602 -34020 -6560 -33920
rect -8602 -34652 -8582 -34020
rect -10281 -34806 -8582 -34652
rect -8175 -34652 -6560 -34020
rect -6496 -33920 -6476 -33370
rect -6069 -33370 -4370 -33206
rect -6069 -33920 -4454 -33370
rect -6496 -34020 -4454 -33920
rect -6496 -34652 -6476 -34020
rect -8175 -34806 -6476 -34652
rect -6069 -34652 -4454 -34020
rect -4390 -33920 -4370 -33370
rect -3963 -33370 -2264 -33206
rect -3963 -33920 -2348 -33370
rect -4390 -34020 -2348 -33920
rect -4390 -34652 -4370 -34020
rect -6069 -34806 -4370 -34652
rect -3963 -34652 -2348 -34020
rect -2284 -34652 -2264 -33370
rect -3963 -34806 -2264 -34652
rect -1857 -33370 -158 -33206
rect -1857 -34652 -242 -33370
rect -178 -33950 -158 -33370
rect 249 -33370 1948 -33206
rect 249 -33950 1864 -33370
rect -178 -34050 1864 -33950
rect -178 -34652 -158 -34050
rect -1857 -34806 -158 -34652
rect 249 -34652 1864 -34050
rect 1928 -33950 1948 -33370
rect 2355 -33370 4054 -33206
rect 2355 -33950 3970 -33370
rect 1928 -34050 3970 -33950
rect 1928 -34652 1948 -34050
rect 249 -34806 1948 -34652
rect 2355 -34652 3970 -34050
rect 4034 -33950 4054 -33370
rect 4461 -33370 6160 -33206
rect 4461 -33950 6076 -33370
rect 4034 -34050 6076 -33950
rect 4034 -34652 4054 -34050
rect 2355 -34806 4054 -34652
rect 4461 -34652 6076 -34050
rect 6140 -34652 6160 -33370
rect 4461 -34806 6160 -34652
rect 6567 -33370 8266 -33206
rect 6567 -34652 8182 -33370
rect 8246 -34652 8266 -33370
rect 6567 -34806 8266 -34652
rect -26392 -35206 -26292 -34806
rect -24286 -35206 -24186 -34806
rect -22180 -35206 -22080 -34806
rect -15854 -35206 -15754 -34806
rect -13748 -35206 -13648 -34806
rect -11642 -35206 -11542 -34806
rect -9536 -35206 -9436 -34806
rect -7430 -35206 -7330 -34806
rect -5324 -35206 -5224 -34806
rect -3264 -35206 -3164 -34806
rect 964 -35206 1064 -34806
rect 3060 -35206 3160 -34806
rect 5228 -35206 5328 -34806
rect -29235 -35370 -27536 -35206
rect -29235 -36652 -27620 -35370
rect -27556 -36652 -27536 -35370
rect -29235 -36806 -27536 -36652
rect -27129 -35370 -25430 -35206
rect -27129 -36652 -25514 -35370
rect -25450 -35916 -25430 -35370
rect -25023 -35370 -23324 -35206
rect -25023 -35916 -23408 -35370
rect -25450 -36016 -23408 -35916
rect -25450 -36652 -25430 -36016
rect -27129 -36806 -25430 -36652
rect -25023 -36652 -23408 -36016
rect -23344 -35916 -23324 -35370
rect -22917 -35370 -21218 -35206
rect -22917 -35916 -21302 -35370
rect -23344 -36016 -21302 -35916
rect -23344 -36652 -23324 -36016
rect -25023 -36806 -23324 -36652
rect -22917 -36652 -21302 -36016
rect -21238 -36652 -21218 -35370
rect -22917 -36806 -21218 -36652
rect -20811 -35370 -19112 -35206
rect -20811 -36652 -19196 -35370
rect -19132 -35958 -19112 -35370
rect -18705 -35370 -17006 -35206
rect -18705 -35958 -17090 -35370
rect -19132 -36058 -17090 -35958
rect -19132 -36652 -19112 -36058
rect -20811 -36806 -19112 -36652
rect -18705 -36652 -17090 -36058
rect -17026 -35958 -17006 -35370
rect -16599 -35370 -14900 -35206
rect -16599 -35958 -14984 -35370
rect -17026 -36058 -14984 -35958
rect -17026 -36652 -17006 -36058
rect -18705 -36806 -17006 -36652
rect -16599 -36652 -14984 -36058
rect -14920 -35958 -14900 -35370
rect -14493 -35370 -12794 -35206
rect -14493 -35958 -12878 -35370
rect -14920 -36058 -12878 -35958
rect -14920 -36652 -14900 -36058
rect -16599 -36806 -14900 -36652
rect -14493 -36652 -12878 -36058
rect -12814 -35958 -12794 -35370
rect -12387 -35370 -10688 -35206
rect -12387 -35958 -10772 -35370
rect -12814 -36058 -10772 -35958
rect -12814 -36652 -12794 -36058
rect -14493 -36806 -12794 -36652
rect -12387 -36652 -10772 -36058
rect -10708 -35958 -10688 -35370
rect -10281 -35370 -8582 -35206
rect -10281 -35958 -8666 -35370
rect -10708 -36058 -8666 -35958
rect -10708 -36652 -10688 -36058
rect -12387 -36806 -10688 -36652
rect -10281 -36652 -8666 -36058
rect -8602 -35958 -8582 -35370
rect -8175 -35370 -6476 -35206
rect -8175 -35958 -6560 -35370
rect -8602 -36058 -6560 -35958
rect -8602 -36652 -8582 -36058
rect -10281 -36806 -8582 -36652
rect -8175 -36652 -6560 -36058
rect -6496 -35958 -6476 -35370
rect -6069 -35370 -4370 -35206
rect -6069 -35958 -4454 -35370
rect -6496 -36058 -4454 -35958
rect -6496 -36652 -6476 -36058
rect -8175 -36806 -6476 -36652
rect -6069 -36652 -4454 -36058
rect -4390 -35958 -4370 -35370
rect -3963 -35370 -2264 -35206
rect -3963 -35958 -2348 -35370
rect -4390 -36058 -2348 -35958
rect -4390 -36652 -4370 -36058
rect -6069 -36806 -4370 -36652
rect -3963 -36652 -2348 -36058
rect -2284 -35958 -2264 -35370
rect -1857 -35370 -158 -35206
rect -1857 -35958 -242 -35370
rect -2284 -36058 -242 -35958
rect -2284 -36652 -2264 -36058
rect -3963 -36806 -2264 -36652
rect -1857 -36652 -242 -36058
rect -178 -36652 -158 -35370
rect -1857 -36806 -158 -36652
rect 249 -35370 1948 -35206
rect 249 -36652 1864 -35370
rect 1928 -35934 1948 -35370
rect 2355 -35370 4054 -35206
rect 2355 -35934 3970 -35370
rect 1928 -36034 3970 -35934
rect 1928 -36652 1948 -36034
rect 249 -36806 1948 -36652
rect 2355 -36652 3970 -36034
rect 4034 -35950 4054 -35370
rect 4461 -35370 6160 -35206
rect 4461 -35950 6076 -35370
rect 4034 -36050 6076 -35950
rect 4034 -36652 4054 -36050
rect 2355 -36806 4054 -36652
rect 4461 -36652 6076 -36050
rect 6140 -36652 6160 -35370
rect 4461 -36806 6160 -36652
rect 6567 -35370 8266 -35206
rect 6567 -36652 8182 -35370
rect 8246 -36652 8266 -35370
rect 6567 -36806 8266 -36652
rect -26392 -37206 -26292 -36806
rect -24286 -37206 -24186 -36806
rect -20078 -37206 -19978 -36806
rect -1110 -37206 -1010 -36806
rect 964 -37206 1064 -36806
rect 3060 -37206 3160 -36806
rect 5228 -37206 5328 -36806
rect -29235 -37370 -27536 -37206
rect -29235 -38652 -27620 -37370
rect -27556 -38652 -27536 -37370
rect -29235 -38806 -27536 -38652
rect -27129 -37370 -25430 -37206
rect -27129 -38652 -25514 -37370
rect -25450 -37942 -25430 -37370
rect -25023 -37370 -23324 -37206
rect -25023 -37942 -23408 -37370
rect -25450 -38042 -23408 -37942
rect -25450 -38652 -25430 -38042
rect -27129 -38806 -25430 -38652
rect -25023 -38652 -23408 -38042
rect -23344 -38652 -23324 -37370
rect -25023 -38806 -23324 -38652
rect -22917 -37370 -21218 -37206
rect -22917 -38652 -21302 -37370
rect -21238 -37980 -21218 -37370
rect -20811 -37370 -19112 -37206
rect -20811 -37980 -19196 -37370
rect -21238 -38080 -19196 -37980
rect -21238 -38652 -21218 -38080
rect -22917 -38806 -21218 -38652
rect -20811 -38652 -19196 -38080
rect -19132 -38652 -19112 -37370
rect -20811 -38806 -19112 -38652
rect -18705 -37370 -17006 -37206
rect -18705 -38652 -17090 -37370
rect -17026 -37936 -17006 -37370
rect -16599 -37370 -14900 -37206
rect -16599 -37936 -14984 -37370
rect -17026 -38036 -14984 -37936
rect -17026 -38652 -17006 -38036
rect -18705 -38806 -17006 -38652
rect -16599 -38652 -14984 -38036
rect -14920 -37936 -14900 -37370
rect -14493 -37370 -12794 -37206
rect -14493 -37936 -12878 -37370
rect -14920 -38036 -12878 -37936
rect -14920 -38652 -14900 -38036
rect -16599 -38806 -14900 -38652
rect -14493 -38652 -12878 -38036
rect -12814 -37936 -12794 -37370
rect -12387 -37370 -10688 -37206
rect -12387 -37936 -10772 -37370
rect -12814 -38036 -10772 -37936
rect -12814 -38652 -12794 -38036
rect -14493 -38806 -12794 -38652
rect -12387 -38652 -10772 -38036
rect -10708 -37936 -10688 -37370
rect -10281 -37370 -8582 -37206
rect -10281 -37936 -8666 -37370
rect -10708 -38036 -8666 -37936
rect -10708 -38652 -10688 -38036
rect -12387 -38806 -10688 -38652
rect -10281 -38652 -8666 -38036
rect -8602 -37936 -8582 -37370
rect -8175 -37370 -6476 -37206
rect -8175 -37936 -6560 -37370
rect -8602 -38036 -6560 -37936
rect -8602 -38652 -8582 -38036
rect -10281 -38806 -8582 -38652
rect -8175 -38652 -6560 -38036
rect -6496 -37936 -6476 -37370
rect -6069 -37370 -4370 -37206
rect -6069 -37936 -4454 -37370
rect -6496 -38036 -4454 -37936
rect -6496 -38652 -6476 -38036
rect -8175 -38806 -6476 -38652
rect -6069 -38652 -4454 -38036
rect -4390 -37936 -4370 -37370
rect -3963 -37370 -2264 -37206
rect -3963 -37936 -2348 -37370
rect -4390 -38036 -2348 -37936
rect -4390 -38652 -4370 -38036
rect -6069 -38806 -4370 -38652
rect -3963 -38652 -2348 -38036
rect -2284 -38652 -2264 -37370
rect -3963 -38806 -2264 -38652
rect -1857 -37370 -158 -37206
rect -1857 -38652 -242 -37370
rect -178 -38652 -158 -37370
rect -1857 -38806 -158 -38652
rect 249 -37370 1948 -37206
rect 249 -38652 1864 -37370
rect 1928 -37918 1948 -37370
rect 2355 -37370 4054 -37206
rect 2355 -37918 3970 -37370
rect 1928 -38018 3970 -37918
rect 1928 -38652 1948 -38018
rect 249 -38806 1948 -38652
rect 2355 -38652 3970 -38018
rect 4034 -37950 4054 -37370
rect 4461 -37370 6160 -37206
rect 4461 -37950 6076 -37370
rect 4034 -38050 6076 -37950
rect 4034 -38652 4054 -38050
rect 2355 -38806 4054 -38652
rect 4461 -38652 6076 -38050
rect 6140 -38652 6160 -37370
rect 4461 -38806 6160 -38652
rect 6567 -37370 8266 -37206
rect 6567 -38652 8182 -37370
rect 8246 -38652 8266 -37370
rect 6567 -38806 8266 -38652
rect -26392 -39206 -26292 -38806
rect -24286 -39206 -24186 -38806
rect -22154 -39206 -22054 -38806
rect -20078 -39206 -19978 -38806
rect -17986 -39206 -17886 -38806
rect -15882 -39206 -15782 -38806
rect -5340 -39206 -5240 -38806
rect -3180 -39206 -3080 -38806
rect -1110 -39206 -1010 -38806
rect 3060 -39206 3160 -38806
rect 5228 -39206 5328 -38806
rect -29235 -39370 -27536 -39206
rect -29235 -40652 -27620 -39370
rect -27556 -40652 -27536 -39370
rect -29235 -40806 -27536 -40652
rect -27129 -39370 -25430 -39206
rect -27129 -40652 -25514 -39370
rect -25450 -39962 -25430 -39370
rect -25023 -39370 -23324 -39206
rect -25023 -39962 -23408 -39370
rect -25450 -40062 -23408 -39962
rect -25450 -40652 -25430 -40062
rect -27129 -40806 -25430 -40652
rect -25023 -40652 -23408 -40062
rect -23344 -40652 -23324 -39370
rect -25023 -40806 -23324 -40652
rect -22917 -39370 -21218 -39206
rect -22917 -40652 -21302 -39370
rect -21238 -39980 -21218 -39370
rect -20811 -39370 -19112 -39206
rect -20811 -39980 -19196 -39370
rect -21238 -40080 -19196 -39980
rect -21238 -40652 -21218 -40080
rect -22917 -40806 -21218 -40652
rect -20811 -40652 -19196 -40080
rect -19132 -40652 -19112 -39370
rect -20811 -40806 -19112 -40652
rect -18705 -39370 -17006 -39206
rect -18705 -40652 -17090 -39370
rect -17026 -39928 -17006 -39370
rect -16599 -39370 -14900 -39206
rect -16599 -39928 -14984 -39370
rect -17026 -40028 -14984 -39928
rect -17026 -40652 -17006 -40028
rect -18705 -40806 -17006 -40652
rect -16599 -40652 -14984 -40028
rect -14920 -40652 -14900 -39370
rect -16599 -40806 -14900 -40652
rect -14493 -39370 -12794 -39206
rect -14493 -40652 -12878 -39370
rect -12814 -39906 -12794 -39370
rect -12387 -39370 -10688 -39206
rect -12387 -39906 -10772 -39370
rect -12814 -40006 -10772 -39906
rect -12814 -40652 -12794 -40006
rect -14493 -40774 -12794 -40652
rect -14493 -40806 -14318 -40774
rect -26392 -41206 -26292 -40806
rect -24286 -41206 -24186 -40806
rect -22154 -41206 -22054 -40806
rect -20078 -41206 -19978 -40806
rect -17986 -41206 -17886 -40806
rect -14323 -40874 -14318 -40806
rect -14218 -40806 -12794 -40774
rect -12387 -40652 -10772 -40006
rect -10708 -39906 -10688 -39370
rect -10281 -39370 -8582 -39206
rect -10281 -39906 -8666 -39370
rect -10708 -40006 -8666 -39906
rect -10708 -40652 -10688 -40006
rect -12387 -40806 -10688 -40652
rect -10281 -40652 -8666 -40006
rect -8602 -39906 -8582 -39370
rect -8175 -39370 -6476 -39206
rect -8175 -39906 -6560 -39370
rect -8602 -40006 -6560 -39906
rect -8602 -40652 -8582 -40006
rect -10281 -40806 -8582 -40652
rect -8175 -40652 -6560 -40006
rect -6496 -40652 -6476 -39370
rect -8175 -40806 -6476 -40652
rect -6069 -39370 -4370 -39206
rect -6069 -40652 -4454 -39370
rect -4390 -39968 -4370 -39370
rect -3963 -39370 -2264 -39206
rect -3963 -39968 -2348 -39370
rect -4390 -40068 -2348 -39968
rect -4390 -40652 -4370 -40068
rect -6069 -40806 -4370 -40652
rect -3963 -40652 -2348 -40068
rect -2284 -40652 -2264 -39370
rect -3963 -40806 -2264 -40652
rect -1857 -39370 -158 -39206
rect -1857 -40652 -242 -39370
rect -178 -39950 -158 -39370
rect 249 -39370 1948 -39206
rect 249 -39950 1864 -39370
rect -178 -40050 1864 -39950
rect -178 -40652 -158 -40050
rect -1857 -40806 -158 -40652
rect 249 -40652 1864 -40050
rect 1928 -40652 1948 -39370
rect 249 -40806 1948 -40652
rect 2355 -39370 4054 -39206
rect 2355 -40652 3970 -39370
rect 4034 -39950 4054 -39370
rect 4461 -39370 6160 -39206
rect 4461 -39950 6076 -39370
rect 4034 -40050 6076 -39950
rect 4034 -40652 4054 -40050
rect 2355 -40806 4054 -40652
rect 4461 -40652 6076 -40050
rect 6140 -40652 6160 -39370
rect 4461 -40806 6160 -40652
rect 6567 -39370 8266 -39206
rect 6567 -40652 8182 -39370
rect 8246 -40652 8266 -39370
rect 6567 -40806 8266 -40652
rect -14218 -40874 -14213 -40806
rect -14323 -40879 -14213 -40874
rect -7404 -40857 -7304 -40806
rect -7404 -40947 -7399 -40857
rect -7309 -40947 -7304 -40857
rect -7404 -40952 -7304 -40947
rect -13180 -41094 -13048 -41088
rect -15860 -41129 -15760 -41124
rect -15860 -41206 -15855 -41129
rect -29235 -41370 -27536 -41206
rect -29235 -42652 -27620 -41370
rect -27556 -42652 -27536 -41370
rect -29235 -42806 -27536 -42652
rect -27129 -41370 -25430 -41206
rect -27129 -42652 -25514 -41370
rect -25450 -41954 -25430 -41370
rect -25023 -41370 -23324 -41206
rect -25023 -41954 -23408 -41370
rect -25450 -42054 -23408 -41954
rect -25450 -42652 -25430 -42054
rect -27129 -42806 -25430 -42652
rect -25023 -42652 -23408 -42054
rect -23344 -42652 -23324 -41370
rect -25023 -42806 -23324 -42652
rect -22917 -41370 -21218 -41206
rect -22917 -42652 -21302 -41370
rect -21238 -41980 -21218 -41370
rect -20811 -41370 -19112 -41206
rect -20811 -41980 -19196 -41370
rect -21238 -42080 -19196 -41980
rect -21238 -42652 -21218 -42080
rect -22917 -42806 -21218 -42652
rect -20811 -42652 -19196 -42080
rect -19132 -42652 -19112 -41370
rect -20811 -42806 -19112 -42652
rect -18705 -41370 -17006 -41206
rect -18705 -42652 -17090 -41370
rect -17026 -42652 -17006 -41370
rect -18705 -42806 -17006 -42652
rect -16599 -41219 -15855 -41206
rect -15765 -41206 -15760 -41129
rect -13180 -41194 -13168 -41094
rect -13068 -41194 -13048 -41094
rect -13180 -41206 -13048 -41194
rect -7978 -41099 -7878 -41094
rect -7978 -41189 -7973 -41099
rect -7883 -41189 -7878 -41099
rect -7978 -41206 -7878 -41189
rect -5315 -41146 -5205 -41141
rect -5315 -41206 -5310 -41146
rect -15765 -41219 -14900 -41206
rect -16599 -41370 -14900 -41219
rect -16599 -42652 -14984 -41370
rect -14920 -42652 -14900 -41370
rect -14493 -41370 -12794 -41206
rect -14493 -42464 -12878 -41370
rect -14632 -42469 -12878 -42464
rect -14632 -42559 -14627 -42469
rect -14537 -42559 -12878 -42469
rect -14632 -42564 -12878 -42559
rect -16599 -42806 -14900 -42652
rect -14493 -42652 -12878 -42564
rect -12814 -42652 -12794 -41370
rect -14493 -42806 -12794 -42652
rect -12387 -41370 -10688 -41206
rect -12387 -42652 -10772 -41370
rect -10708 -41924 -10688 -41370
rect -10281 -41370 -8582 -41206
rect -10281 -41924 -8666 -41370
rect -10708 -42024 -8666 -41924
rect -10708 -42652 -10688 -42024
rect -12387 -42806 -10688 -42652
rect -10281 -42652 -8666 -42024
rect -8602 -42652 -8582 -41370
rect -10281 -42806 -8582 -42652
rect -8175 -41370 -6476 -41206
rect -8175 -42652 -6560 -41370
rect -6496 -42532 -6476 -41370
rect -6069 -41246 -5310 -41206
rect -5210 -41206 -5205 -41146
rect -3180 -41206 -3080 -40806
rect -1110 -41206 -1010 -40806
rect 1010 -41206 1110 -40806
rect 3060 -41206 3160 -40806
rect 5228 -41206 5328 -40806
rect -5210 -41246 -4370 -41206
rect -6069 -41370 -4370 -41246
rect -6496 -42537 -6332 -42532
rect -6496 -42627 -6427 -42537
rect -6337 -42627 -6332 -42537
rect -6496 -42632 -6332 -42627
rect -6496 -42652 -6476 -42632
rect -8175 -42806 -6476 -42652
rect -6069 -42652 -4454 -41370
rect -4390 -42652 -4370 -41370
rect -6069 -42806 -4370 -42652
rect -3963 -41370 -2264 -41206
rect -3963 -42652 -2348 -41370
rect -2284 -42652 -2264 -41370
rect -3963 -42806 -2264 -42652
rect -1857 -41370 -158 -41206
rect -1857 -42652 -242 -41370
rect -178 -41946 -158 -41370
rect 249 -41370 1948 -41206
rect 249 -41946 1864 -41370
rect -178 -42046 1864 -41946
rect -178 -42652 -158 -42046
rect -1857 -42806 -158 -42652
rect 249 -42652 1864 -42046
rect 1928 -42652 1948 -41370
rect 249 -42806 1948 -42652
rect 2355 -41370 4054 -41206
rect 2355 -42652 3970 -41370
rect 4034 -41950 4054 -41370
rect 4461 -41370 6160 -41206
rect 4461 -41950 6076 -41370
rect 4034 -42050 6076 -41950
rect 4034 -42652 4054 -42050
rect 2355 -42806 4054 -42652
rect 4461 -42652 6076 -42050
rect 6140 -42652 6160 -41370
rect 4461 -42806 6160 -42652
rect 6567 -41370 8266 -41206
rect 6567 -42652 8182 -41370
rect 8246 -42652 8266 -41370
rect 6567 -42806 8266 -42652
rect 10276 -42356 25316 -29738
rect 52252 -39086 55140 -39081
rect 52252 -39386 52262 -39086
rect 55130 -39386 55140 -39086
rect 52252 -39391 55140 -39386
rect 56524 -39086 58164 -39081
rect 56524 -39386 56534 -39086
rect 58154 -39386 58164 -39086
rect 56524 -39391 58164 -39386
rect 57456 -40471 57556 -40454
rect 57456 -40476 57475 -40471
rect 57456 -40536 57474 -40476
rect 57456 -40541 57475 -40536
rect 57539 -40541 57556 -40471
rect 57456 -40554 57556 -40541
rect 49186 -41091 52004 -41086
rect 49186 -41181 49191 -41091
rect 49281 -41106 52004 -41091
rect 49281 -41166 51918 -41106
rect 51978 -41166 52004 -41106
rect 49281 -41181 52004 -41166
rect 49186 -41186 52004 -41181
rect 10276 -42648 11814 -42356
rect 22576 -42648 25316 -42356
rect -26392 -43206 -26292 -42806
rect -24286 -43206 -24186 -42806
rect -22154 -43206 -22054 -42806
rect -20078 -43206 -19978 -42806
rect -17986 -43206 -17886 -42806
rect -15860 -43206 -15760 -42806
rect -11648 -42841 -11548 -42806
rect -11648 -42931 -11643 -42841
rect -11553 -42931 -11548 -42841
rect -11648 -42936 -11548 -42931
rect -9536 -42841 -9436 -42806
rect -9536 -42931 -9531 -42841
rect -9441 -42931 -9436 -42841
rect -9536 -42936 -9436 -42931
rect -7447 -43112 -7337 -43107
rect -13751 -43120 -13641 -43115
rect -13751 -43206 -13746 -43120
rect -29235 -43370 -27536 -43206
rect -29235 -44652 -27620 -43370
rect -27556 -44652 -27536 -43370
rect -29235 -44806 -27536 -44652
rect -27129 -43370 -25430 -43206
rect -27129 -44652 -25514 -43370
rect -25450 -43954 -25430 -43370
rect -25023 -43370 -23324 -43206
rect -25023 -43954 -23408 -43370
rect -25450 -44054 -23408 -43954
rect -25450 -44652 -25430 -44054
rect -27129 -44806 -25430 -44652
rect -25023 -44652 -23408 -44054
rect -23344 -44652 -23324 -43370
rect -25023 -44806 -23324 -44652
rect -22917 -43370 -21218 -43206
rect -22917 -44652 -21302 -43370
rect -21238 -43980 -21218 -43370
rect -20811 -43370 -19112 -43206
rect -20811 -43980 -19196 -43370
rect -21238 -44080 -19196 -43980
rect -21238 -44652 -21218 -44080
rect -22917 -44806 -21218 -44652
rect -20811 -44652 -19196 -44080
rect -19132 -44652 -19112 -43370
rect -20811 -44806 -19112 -44652
rect -18705 -43370 -17006 -43206
rect -18705 -44652 -17090 -43370
rect -17026 -44652 -17006 -43370
rect -18705 -44806 -17006 -44652
rect -16599 -43370 -14900 -43206
rect -16599 -44652 -14984 -43370
rect -14920 -44652 -14900 -43370
rect -16599 -44806 -14900 -44652
rect -14493 -43220 -13746 -43206
rect -13646 -43206 -13641 -43120
rect -7447 -43206 -7442 -43112
rect -13646 -43220 -12794 -43206
rect -14493 -43370 -12794 -43220
rect -14493 -44652 -12878 -43370
rect -12814 -44652 -12794 -43370
rect -14493 -44806 -12794 -44652
rect -12387 -43370 -10688 -43206
rect -12387 -44652 -10772 -43370
rect -10708 -44652 -10688 -43370
rect -12387 -44806 -10688 -44652
rect -10281 -43370 -8582 -43206
rect -10281 -44652 -8666 -43370
rect -8602 -44652 -8582 -43370
rect -10281 -44806 -8582 -44652
rect -8175 -43212 -7442 -43206
rect -7342 -43206 -7337 -43112
rect -5306 -43206 -5206 -42806
rect -3180 -43206 -3080 -42806
rect -1110 -43206 -1010 -42806
rect 1010 -43206 1110 -42806
rect 3060 -43206 3160 -42806
rect 5228 -43206 5328 -42806
rect 10276 -42956 25316 -42648
rect 52310 -41962 52510 -41908
rect 52310 -42022 52380 -41962
rect 52440 -42022 52510 -41962
rect 27759 -42922 27857 -42917
rect 27758 -42923 27858 -42922
rect 26958 -42937 27090 -42924
rect -7342 -43212 -6476 -43206
rect -8175 -43370 -6476 -43212
rect -8175 -44652 -6560 -43370
rect -6496 -44652 -6476 -43370
rect -8175 -44806 -6476 -44652
rect -6069 -43370 -4370 -43206
rect -6069 -44652 -4454 -43370
rect -4390 -44652 -4370 -43370
rect -6069 -44806 -4370 -44652
rect -3963 -43370 -2264 -43206
rect -3963 -44652 -2348 -43370
rect -2284 -44652 -2264 -43370
rect -3963 -44806 -2264 -44652
rect -1857 -43370 -158 -43206
rect -1857 -44652 -242 -43370
rect -178 -43916 -158 -43370
rect 249 -43370 1948 -43206
rect 249 -43916 1864 -43370
rect -178 -44016 1864 -43916
rect -178 -44652 -158 -44016
rect -1857 -44806 -158 -44652
rect 249 -44652 1864 -44016
rect 1928 -44652 1948 -43370
rect 249 -44806 1948 -44652
rect 2355 -43370 4054 -43206
rect 2355 -44652 3970 -43370
rect 4034 -43950 4054 -43370
rect 4461 -43370 6160 -43206
rect 4461 -43950 6076 -43370
rect 4034 -44050 6076 -43950
rect 4034 -44652 4054 -44050
rect 2355 -44806 4054 -44652
rect 4461 -44652 6076 -44050
rect 6140 -44652 6160 -43370
rect 4461 -44806 6160 -44652
rect 6567 -43370 8266 -43206
rect 6567 -44652 8182 -43370
rect 8246 -44652 8266 -43370
rect 10276 -43450 24066 -42956
rect 26958 -43001 26981 -42937
rect 27051 -43001 27090 -42937
rect 26958 -43002 26986 -43001
rect 27046 -43002 27090 -43001
rect 26958 -43018 27090 -43002
rect 27758 -43021 27759 -42923
rect 27857 -43021 27858 -42923
rect 27758 -43022 27858 -43021
rect 27759 -43027 27857 -43022
rect 10276 -43894 24068 -43450
rect 23730 -43896 24068 -43894
rect 6567 -44806 8266 -44652
rect -26392 -45206 -26292 -44806
rect -24286 -45206 -24186 -44806
rect -22154 -45206 -22054 -44806
rect -20078 -45206 -19978 -44806
rect -17986 -45206 -17886 -44806
rect -15860 -45206 -15760 -44806
rect -13746 -45206 -13646 -44806
rect -10922 -44837 -10822 -44806
rect -10922 -44927 -10917 -44837
rect -10827 -44927 -10822 -44837
rect -10922 -44932 -10822 -44927
rect -10169 -45124 -10059 -45119
rect -10169 -45206 -10164 -45124
rect -29235 -45370 -27536 -45206
rect -29235 -46652 -27620 -45370
rect -27556 -46652 -27536 -45370
rect -29235 -46806 -27536 -46652
rect -27129 -45370 -25430 -45206
rect -27129 -46652 -25514 -45370
rect -25450 -45954 -25430 -45370
rect -25023 -45370 -23324 -45206
rect -25023 -45954 -23408 -45370
rect -25450 -46054 -23408 -45954
rect -25450 -46652 -25430 -46054
rect -27129 -46806 -25430 -46652
rect -25023 -46652 -23408 -46054
rect -23344 -46652 -23324 -45370
rect -25023 -46806 -23324 -46652
rect -22917 -45370 -21218 -45206
rect -22917 -46652 -21302 -45370
rect -21238 -45980 -21218 -45370
rect -20811 -45370 -19112 -45206
rect -20811 -45980 -19196 -45370
rect -21238 -46080 -19196 -45980
rect -21238 -46652 -21218 -46080
rect -22917 -46806 -21218 -46652
rect -20811 -46652 -19196 -46080
rect -19132 -46652 -19112 -45370
rect -20811 -46806 -19112 -46652
rect -18705 -45370 -17006 -45206
rect -18705 -46652 -17090 -45370
rect -17026 -46652 -17006 -45370
rect -18705 -46806 -17006 -46652
rect -16599 -45370 -14900 -45206
rect -16599 -46652 -14984 -45370
rect -14920 -46652 -14900 -45370
rect -16599 -46806 -14900 -46652
rect -14493 -45370 -12794 -45206
rect -14493 -46652 -12878 -45370
rect -12814 -46652 -12794 -45370
rect -14493 -46806 -12794 -46652
rect -12387 -45370 -10688 -45206
rect -12387 -46652 -10772 -45370
rect -10708 -46652 -10688 -45370
rect -12387 -46806 -10688 -46652
rect -10281 -45224 -10164 -45206
rect -10064 -45206 -10059 -45124
rect -7444 -45206 -7344 -44806
rect -5306 -45206 -5206 -44806
rect -3180 -45206 -3080 -44806
rect -1110 -45206 -1010 -44806
rect 1010 -45206 1110 -44806
rect 3060 -45206 3160 -44806
rect 5228 -45206 5328 -44806
rect -10064 -45224 -8582 -45206
rect -10281 -45370 -8582 -45224
rect -10281 -46652 -8666 -45370
rect -8602 -46652 -8582 -45370
rect -10281 -46806 -8582 -46652
rect -8175 -45370 -6476 -45206
rect -8175 -46652 -6560 -45370
rect -6496 -46652 -6476 -45370
rect -8175 -46758 -6476 -46652
rect -8175 -46806 -7444 -46758
rect -26392 -47206 -26292 -46806
rect -24286 -47206 -24186 -46806
rect -22154 -47206 -22054 -46806
rect -20078 -47206 -19978 -46806
rect -17986 -47206 -17886 -46806
rect -15860 -47206 -15760 -46806
rect -13746 -46841 -13646 -46806
rect -13746 -46931 -13741 -46841
rect -13651 -46931 -13646 -46841
rect -7449 -46858 -7444 -46806
rect -7344 -46806 -6476 -46758
rect -6069 -45370 -4370 -45206
rect -6069 -46652 -4454 -45370
rect -4390 -46652 -4370 -45370
rect -6069 -46806 -4370 -46652
rect -3963 -45370 -2264 -45206
rect -3963 -46652 -2348 -45370
rect -2284 -46652 -2264 -45370
rect -3963 -46806 -2264 -46652
rect -1857 -45370 -158 -45206
rect -1857 -46652 -242 -45370
rect -178 -45948 -158 -45370
rect 249 -45370 1948 -45206
rect 249 -45948 1864 -45370
rect -178 -46048 1864 -45948
rect -178 -46652 -158 -46048
rect -1857 -46806 -158 -46652
rect 249 -46652 1864 -46048
rect 1928 -46652 1948 -45370
rect 249 -46806 1948 -46652
rect 2355 -45370 4054 -45206
rect 2355 -46652 3970 -45370
rect 4034 -45950 4054 -45370
rect 4461 -45370 6160 -45206
rect 4461 -45950 6076 -45370
rect 4034 -46050 6076 -45950
rect 4034 -46652 4054 -46050
rect 2355 -46806 4054 -46652
rect 4461 -46652 6076 -46050
rect 6140 -46652 6160 -45370
rect 4461 -46806 6160 -46652
rect 6567 -45370 8266 -45206
rect 6567 -46652 8182 -45370
rect 8246 -46652 8266 -45370
rect 6567 -46806 8266 -46652
rect -7344 -46858 -7339 -46806
rect -7449 -46863 -7339 -46858
rect -13746 -46936 -13646 -46931
rect -9542 -47109 -9442 -47104
rect -11649 -47134 -11539 -47129
rect -11649 -47206 -11644 -47134
rect -29235 -47370 -27536 -47206
rect -29235 -48652 -27620 -47370
rect -27556 -48652 -27536 -47370
rect -29235 -48806 -27536 -48652
rect -27129 -47370 -25430 -47206
rect -27129 -48652 -25514 -47370
rect -25450 -47954 -25430 -47370
rect -25023 -47370 -23324 -47206
rect -25023 -47954 -23408 -47370
rect -25450 -48054 -23408 -47954
rect -25450 -48652 -25430 -48054
rect -27129 -48806 -25430 -48652
rect -25023 -48652 -23408 -48054
rect -23344 -48652 -23324 -47370
rect -25023 -48806 -23324 -48652
rect -22917 -47370 -21218 -47206
rect -22917 -48652 -21302 -47370
rect -21238 -47980 -21218 -47370
rect -20811 -47370 -19112 -47206
rect -20811 -47980 -19196 -47370
rect -21238 -48080 -19196 -47980
rect -21238 -48652 -21218 -48080
rect -22917 -48806 -21218 -48652
rect -20811 -48652 -19196 -48080
rect -19132 -48652 -19112 -47370
rect -20811 -48806 -19112 -48652
rect -18705 -47370 -17006 -47206
rect -18705 -48652 -17090 -47370
rect -17026 -48652 -17006 -47370
rect -18705 -48806 -17006 -48652
rect -16599 -47370 -14900 -47206
rect -16599 -48652 -14984 -47370
rect -14920 -48652 -14900 -47370
rect -14493 -47370 -12794 -47206
rect -14493 -47406 -12878 -47370
rect -14654 -47424 -12878 -47406
rect -14654 -47524 -14632 -47424
rect -14532 -47524 -12878 -47424
rect -14654 -47554 -12878 -47524
rect -16599 -48806 -14900 -48652
rect -14493 -48652 -12878 -47554
rect -12814 -48652 -12794 -47370
rect -14493 -48806 -12794 -48652
rect -12387 -47234 -11644 -47206
rect -11544 -47206 -11539 -47134
rect -9542 -47199 -9537 -47109
rect -9447 -47199 -9442 -47109
rect -9542 -47206 -9442 -47199
rect -5306 -47206 -5206 -46806
rect -3180 -47206 -3080 -46806
rect -1110 -47206 -1010 -46806
rect 1010 -47206 1110 -46806
rect 3060 -47206 3160 -46806
rect 5228 -47206 5328 -46806
rect -11544 -47234 -10688 -47206
rect -12387 -47370 -10688 -47234
rect -12387 -48652 -10772 -47370
rect -10708 -47914 -10688 -47370
rect -10281 -47370 -8582 -47206
rect -10281 -47914 -8666 -47370
rect -10708 -48014 -8666 -47914
rect -10708 -48652 -10688 -48014
rect -12387 -48806 -10688 -48652
rect -10281 -48652 -8666 -48014
rect -8602 -48652 -8582 -47370
rect -10281 -48806 -8582 -48652
rect -8175 -47370 -6476 -47206
rect -8175 -48652 -6560 -47370
rect -6496 -47516 -6476 -47370
rect -6069 -47370 -4370 -47206
rect -6496 -47530 -6320 -47516
rect -6496 -47630 -6432 -47530
rect -6332 -47630 -6320 -47530
rect -6496 -47648 -6320 -47630
rect -6496 -48652 -6476 -47648
rect -8175 -48806 -6476 -48652
rect -6069 -48652 -4454 -47370
rect -4390 -48652 -4370 -47370
rect -6069 -48778 -4370 -48652
rect -6069 -48806 -5312 -48778
rect -26392 -49206 -26292 -48806
rect -24286 -49206 -24186 -48806
rect -22154 -49206 -22054 -48806
rect -20078 -49206 -19978 -48806
rect -17986 -49206 -17886 -48806
rect -15860 -48857 -15760 -48806
rect -15860 -48947 -15855 -48857
rect -15765 -48947 -15760 -48857
rect -15860 -48952 -15760 -48947
rect -13004 -48855 -12904 -48806
rect -13004 -48945 -12999 -48855
rect -12909 -48945 -12904 -48855
rect -13004 -48950 -12904 -48945
rect -8074 -48850 -7938 -48806
rect -8074 -48950 -8060 -48850
rect -7960 -48950 -7938 -48850
rect -5317 -48878 -5312 -48806
rect -5212 -48806 -4370 -48778
rect -3963 -47370 -2264 -47206
rect -3963 -48652 -2348 -47370
rect -2284 -48652 -2264 -47370
rect -3963 -48806 -2264 -48652
rect -1857 -47370 -158 -47206
rect -1857 -48652 -242 -47370
rect -178 -47944 -158 -47370
rect 249 -47370 1948 -47206
rect 249 -47944 1864 -47370
rect -178 -48044 1864 -47944
rect -178 -48652 -158 -48044
rect -1857 -48806 -158 -48652
rect 249 -48652 1864 -48044
rect 1928 -48652 1948 -47370
rect 249 -48806 1948 -48652
rect 2355 -47370 4054 -47206
rect 2355 -48652 3970 -47370
rect 4034 -47950 4054 -47370
rect 4461 -47370 6160 -47206
rect 4461 -47950 6076 -47370
rect 4034 -48050 6076 -47950
rect 4034 -48652 4054 -48050
rect 2355 -48806 4054 -48652
rect 4461 -48652 6076 -48050
rect 6140 -48652 6160 -47370
rect 4461 -48806 6160 -48652
rect 6567 -47370 8266 -47206
rect 6567 -48652 8182 -47370
rect 8246 -48652 8266 -47370
rect 6567 -48806 8266 -48652
rect -5212 -48878 -5207 -48806
rect -5317 -48883 -5207 -48878
rect -8074 -48966 -7938 -48950
rect -7436 -49051 -7336 -49046
rect -7436 -49141 -7431 -49051
rect -7341 -49141 -7336 -49051
rect -13761 -49148 -13651 -49143
rect -13761 -49206 -13756 -49148
rect -29235 -49370 -27536 -49206
rect -29235 -50652 -27620 -49370
rect -27556 -50652 -27536 -49370
rect -29235 -50806 -27536 -50652
rect -27129 -49370 -25430 -49206
rect -27129 -50652 -25514 -49370
rect -25450 -49954 -25430 -49370
rect -25023 -49370 -23324 -49206
rect -25023 -49954 -23408 -49370
rect -25450 -50054 -23408 -49954
rect -25450 -50652 -25430 -50054
rect -27129 -50806 -25430 -50652
rect -25023 -50652 -23408 -50054
rect -23344 -50652 -23324 -49370
rect -25023 -50806 -23324 -50652
rect -22917 -49370 -21218 -49206
rect -22917 -50652 -21302 -49370
rect -21238 -49980 -21218 -49370
rect -20811 -49370 -19112 -49206
rect -20811 -49980 -19196 -49370
rect -21238 -50080 -19196 -49980
rect -21238 -50652 -21218 -50080
rect -22917 -50806 -21218 -50652
rect -20811 -50652 -19196 -50080
rect -19132 -50652 -19112 -49370
rect -20811 -50806 -19112 -50652
rect -18705 -49370 -17006 -49206
rect -18705 -50652 -17090 -49370
rect -17026 -49922 -17006 -49370
rect -16599 -49370 -14900 -49206
rect -16599 -49922 -14984 -49370
rect -17026 -50022 -14984 -49922
rect -17026 -50652 -17006 -50022
rect -18705 -50806 -17006 -50652
rect -16599 -50652 -14984 -50022
rect -14920 -50652 -14900 -49370
rect -16599 -50806 -14900 -50652
rect -14493 -49248 -13756 -49206
rect -13656 -49206 -13651 -49148
rect -7436 -49206 -7336 -49141
rect -3180 -49206 -3080 -48806
rect -1110 -49206 -1010 -48806
rect 1010 -49206 1110 -48806
rect 3060 -49206 3160 -48806
rect 5228 -49206 5328 -48806
rect -13656 -49248 -12794 -49206
rect -14493 -49370 -12794 -49248
rect -14493 -50652 -12878 -49370
rect -12814 -49906 -12794 -49370
rect -12387 -49370 -10688 -49206
rect -12387 -49906 -10772 -49370
rect -12814 -50006 -10772 -49906
rect -12814 -50652 -12794 -50006
rect -14493 -50806 -12794 -50652
rect -12387 -50652 -10772 -50006
rect -10708 -49906 -10688 -49370
rect -10281 -49370 -8582 -49206
rect -10281 -49906 -8666 -49370
rect -10708 -50006 -8666 -49906
rect -10708 -50652 -10688 -50006
rect -12387 -50806 -10688 -50652
rect -10281 -50652 -8666 -50006
rect -8602 -49906 -8582 -49370
rect -8175 -49370 -6476 -49206
rect -8175 -49906 -6560 -49370
rect -8602 -50006 -6560 -49906
rect -8602 -50652 -8582 -50006
rect -10281 -50806 -8582 -50652
rect -8175 -50652 -6560 -50006
rect -6496 -50652 -6476 -49370
rect -8175 -50806 -6476 -50652
rect -6069 -49370 -4370 -49206
rect -6069 -50652 -4454 -49370
rect -4390 -49940 -4370 -49370
rect -3963 -49370 -2264 -49206
rect -3963 -49940 -2348 -49370
rect -4390 -50040 -2348 -49940
rect -4390 -50652 -4370 -50040
rect -6069 -50806 -4370 -50652
rect -3963 -50652 -2348 -50040
rect -2284 -50652 -2264 -49370
rect -3963 -50806 -2264 -50652
rect -1857 -49370 -158 -49206
rect -1857 -50652 -242 -49370
rect -178 -49926 -158 -49370
rect 249 -49370 1948 -49206
rect 249 -49926 1864 -49370
rect -178 -50026 1864 -49926
rect -178 -50652 -158 -50026
rect -1857 -50806 -158 -50652
rect 249 -50652 1864 -50026
rect 1928 -50652 1948 -49370
rect 249 -50806 1948 -50652
rect 2355 -49370 4054 -49206
rect 2355 -50652 3970 -49370
rect 4034 -49950 4054 -49370
rect 4461 -49370 6160 -49206
rect 4461 -49950 6076 -49370
rect 4034 -50050 6076 -49950
rect 4034 -50652 4054 -50050
rect 2355 -50806 4054 -50652
rect 4461 -50652 6076 -50050
rect 6140 -50652 6160 -49370
rect 4461 -50806 6160 -50652
rect 6567 -49370 8266 -49206
rect 6567 -50652 8182 -49370
rect 8246 -50652 8266 -49370
rect 6567 -50806 8266 -50652
rect -26392 -51206 -26292 -50806
rect -24286 -51206 -24186 -50806
rect -20078 -51206 -19978 -50806
rect -17986 -51206 -17886 -50806
rect -15868 -51206 -15768 -50806
rect -5324 -51206 -5224 -50806
rect -3180 -51206 -3080 -50806
rect -1110 -51206 -1010 -50806
rect 1010 -51206 1110 -50806
rect 3060 -51206 3160 -50806
rect 5228 -51206 5328 -50806
rect -29235 -51370 -27536 -51206
rect -29235 -52652 -27620 -51370
rect -27556 -52652 -27536 -51370
rect -29235 -52806 -27536 -52652
rect -27129 -51370 -25430 -51206
rect -27129 -52652 -25514 -51370
rect -25450 -51954 -25430 -51370
rect -25023 -51370 -23324 -51206
rect -25023 -51954 -23408 -51370
rect -25450 -52054 -23408 -51954
rect -25450 -52652 -25430 -52054
rect -27129 -52806 -25430 -52652
rect -25023 -52652 -23408 -52054
rect -23344 -51956 -23324 -51370
rect -22917 -51370 -21218 -51206
rect -22917 -51956 -21302 -51370
rect -23344 -52056 -21302 -51956
rect -23344 -52652 -23324 -52056
rect -25023 -52806 -23324 -52652
rect -22917 -52652 -21302 -52056
rect -21238 -52652 -21218 -51370
rect -22917 -52806 -21218 -52652
rect -20811 -51370 -19112 -51206
rect -20811 -52652 -19196 -51370
rect -19132 -52652 -19112 -51370
rect -20811 -52806 -19112 -52652
rect -18705 -51370 -17006 -51206
rect -18705 -52652 -17090 -51370
rect -17026 -51980 -17006 -51370
rect -16599 -51370 -14900 -51206
rect -16599 -51980 -14984 -51370
rect -17026 -52080 -14984 -51980
rect -17026 -52652 -17006 -52080
rect -18705 -52806 -17006 -52652
rect -16599 -52652 -14984 -52080
rect -14920 -51980 -14900 -51370
rect -14493 -51370 -12794 -51206
rect -14493 -51980 -12878 -51370
rect -14920 -52080 -12878 -51980
rect -14920 -52652 -14900 -52080
rect -16599 -52806 -14900 -52652
rect -14493 -52652 -12878 -52080
rect -12814 -51980 -12794 -51370
rect -12387 -51370 -10688 -51206
rect -12387 -51980 -10772 -51370
rect -12814 -52080 -10772 -51980
rect -12814 -52652 -12794 -52080
rect -14493 -52806 -12794 -52652
rect -12387 -52652 -10772 -52080
rect -10708 -51980 -10688 -51370
rect -10281 -51370 -8582 -51206
rect -10281 -51980 -8666 -51370
rect -10708 -52080 -8666 -51980
rect -10708 -52652 -10688 -52080
rect -12387 -52806 -10688 -52652
rect -10281 -52652 -8666 -52080
rect -8602 -51980 -8582 -51370
rect -8175 -51370 -6476 -51206
rect -8175 -51980 -6560 -51370
rect -8602 -52080 -6560 -51980
rect -8602 -52652 -8582 -52080
rect -10281 -52806 -8582 -52652
rect -8175 -52652 -6560 -52080
rect -6496 -51980 -6476 -51370
rect -6069 -51370 -4370 -51206
rect -6069 -51980 -4454 -51370
rect -6496 -52080 -4454 -51980
rect -6496 -52652 -6476 -52080
rect -8175 -52806 -6476 -52652
rect -6069 -52652 -4454 -52080
rect -4390 -51980 -4370 -51370
rect -3963 -51370 -2264 -51206
rect -3963 -51980 -2348 -51370
rect -4390 -52080 -2348 -51980
rect -4390 -52652 -4370 -52080
rect -6069 -52806 -4370 -52652
rect -3963 -52652 -2348 -52080
rect -2284 -52652 -2264 -51370
rect -3963 -52806 -2264 -52652
rect -1857 -51370 -158 -51206
rect -1857 -52652 -242 -51370
rect -178 -51970 -158 -51370
rect 249 -51370 1948 -51206
rect 249 -51970 1864 -51370
rect -178 -52070 1864 -51970
rect -178 -52652 -158 -52070
rect -1857 -52806 -158 -52652
rect 249 -52652 1864 -52070
rect 1928 -52652 1948 -51370
rect 249 -52806 1948 -52652
rect 2355 -51370 4054 -51206
rect 2355 -52652 3970 -51370
rect 4034 -51950 4054 -51370
rect 4461 -51370 6160 -51206
rect 4461 -51950 6076 -51370
rect 4034 -52050 6076 -51950
rect 4034 -52652 4054 -52050
rect 2355 -52806 4054 -52652
rect 4461 -52652 6076 -52050
rect 6140 -52652 6160 -51370
rect 4461 -52806 6160 -52652
rect 6567 -51370 8266 -51206
rect 6567 -52652 8182 -51370
rect 8246 -51982 8266 -51370
rect 8246 -51987 14870 -51982
rect 8246 -52077 14775 -51987
rect 14865 -52077 14870 -51987
rect 8246 -52082 14870 -52077
rect 8246 -52652 8266 -52082
rect 6567 -52806 8266 -52652
rect -26392 -53206 -26292 -52806
rect -24286 -53206 -24186 -52806
rect -22226 -53206 -22126 -52806
rect -20078 -53206 -19978 -52806
rect -1110 -53206 -1010 -52806
rect 3060 -53206 3160 -52806
rect 5228 -53206 5328 -52806
rect 8165 -52948 8263 -52943
rect 8164 -52949 14862 -52948
rect 8164 -53047 8165 -52949
rect 8263 -52953 14862 -52949
rect 8263 -53043 14767 -52953
rect 14857 -53043 14862 -52953
rect 8263 -53047 14862 -53043
rect 8164 -53048 14862 -53047
rect 8165 -53053 8263 -53048
rect -29235 -53370 -27536 -53206
rect -29235 -54652 -27620 -53370
rect -27556 -54652 -27536 -53370
rect -29235 -54806 -27536 -54652
rect -27129 -53370 -25430 -53206
rect -27129 -54652 -25514 -53370
rect -25450 -53954 -25430 -53370
rect -25023 -53370 -23324 -53206
rect -25023 -53954 -23408 -53370
rect -25450 -54054 -23408 -53954
rect -25450 -54652 -25430 -54054
rect -27129 -54806 -25430 -54652
rect -25023 -54652 -23408 -54054
rect -23344 -53954 -23324 -53370
rect -22917 -53370 -21218 -53206
rect -22917 -53954 -21302 -53370
rect -23344 -54054 -21302 -53954
rect -23344 -54652 -23324 -54054
rect -25023 -54806 -23324 -54652
rect -22917 -54652 -21302 -54054
rect -21238 -54652 -21218 -53370
rect -22917 -54806 -21218 -54652
rect -20811 -53370 -19112 -53206
rect -20811 -54652 -19196 -53370
rect -19132 -53970 -19112 -53370
rect -18705 -53370 -17006 -53206
rect -18705 -53970 -17090 -53370
rect -19132 -54070 -17090 -53970
rect -19132 -54652 -19112 -54070
rect -20811 -54806 -19112 -54652
rect -18705 -54652 -17090 -54070
rect -17026 -53970 -17006 -53370
rect -16599 -53370 -14900 -53206
rect -16599 -53970 -14984 -53370
rect -17026 -54070 -14984 -53970
rect -17026 -54652 -17006 -54070
rect -18705 -54806 -17006 -54652
rect -16599 -54652 -14984 -54070
rect -14920 -53970 -14900 -53370
rect -14493 -53370 -12794 -53206
rect -14493 -53970 -12878 -53370
rect -14920 -54070 -12878 -53970
rect -14920 -54652 -14900 -54070
rect -16599 -54806 -14900 -54652
rect -14493 -54652 -12878 -54070
rect -12814 -53970 -12794 -53370
rect -12387 -53370 -10688 -53206
rect -12387 -53970 -10772 -53370
rect -12814 -54070 -10772 -53970
rect -12814 -54652 -12794 -54070
rect -14493 -54806 -12794 -54652
rect -12387 -54652 -10772 -54070
rect -10708 -53970 -10688 -53370
rect -10281 -53370 -8582 -53206
rect -10281 -53970 -8666 -53370
rect -10708 -54070 -8666 -53970
rect -10708 -54652 -10688 -54070
rect -12387 -54806 -10688 -54652
rect -10281 -54652 -8666 -54070
rect -8602 -53970 -8582 -53370
rect -8175 -53370 -6476 -53206
rect -8175 -53970 -6560 -53370
rect -8602 -54070 -6560 -53970
rect -8602 -54652 -8582 -54070
rect -10281 -54806 -8582 -54652
rect -8175 -54652 -6560 -54070
rect -6496 -53970 -6476 -53370
rect -6069 -53370 -4370 -53206
rect -6069 -53970 -4454 -53370
rect -6496 -54070 -4454 -53970
rect -6496 -54652 -6476 -54070
rect -8175 -54806 -6476 -54652
rect -6069 -54652 -4454 -54070
rect -4390 -53970 -4370 -53370
rect -3963 -53370 -2264 -53206
rect -3963 -53970 -2348 -53370
rect -4390 -54070 -2348 -53970
rect -4390 -54652 -4370 -54070
rect -6069 -54806 -4370 -54652
rect -3963 -54652 -2348 -54070
rect -2284 -53970 -2264 -53370
rect -1857 -53370 -158 -53206
rect -1857 -53970 -242 -53370
rect -2284 -54070 -242 -53970
rect -2284 -54652 -2264 -54070
rect -3963 -54806 -2264 -54652
rect -1857 -54652 -242 -54070
rect -178 -54652 -158 -53370
rect -1857 -54806 -158 -54652
rect 249 -53370 1948 -53206
rect 249 -54652 1864 -53370
rect 1928 -53950 1948 -53370
rect 2355 -53370 4054 -53206
rect 2355 -53950 3970 -53370
rect 1928 -54050 3970 -53950
rect 1928 -54652 1948 -54050
rect 249 -54806 1948 -54652
rect 2355 -54652 3970 -54050
rect 4034 -53950 4054 -53370
rect 4461 -53370 6160 -53206
rect 4461 -53950 6076 -53370
rect 4034 -54050 6076 -53950
rect 4034 -54652 4054 -54050
rect 2355 -54806 4054 -54652
rect 4461 -54652 6076 -54050
rect 6140 -54652 6160 -53370
rect 4461 -54806 6160 -54652
rect 6567 -53370 8266 -53206
rect 6567 -54652 8182 -53370
rect 8246 -53942 8266 -53370
rect 8246 -53947 14864 -53942
rect 8246 -54037 14769 -53947
rect 14859 -54037 14864 -53947
rect 8246 -54042 14864 -54037
rect 8246 -54652 8266 -54042
rect 6567 -54806 8266 -54652
rect -26392 -55206 -26292 -54806
rect -24286 -55206 -24186 -54806
rect -22180 -55206 -22080 -54806
rect -17970 -55206 -17870 -54806
rect -15864 -55206 -15764 -54806
rect -13758 -55206 -13658 -54806
rect -11652 -55206 -11552 -54806
rect -9546 -55206 -9446 -54806
rect -7440 -55206 -7340 -54806
rect -5340 -55206 -5240 -54806
rect 1010 -55206 1110 -54806
rect 3060 -55206 3160 -54806
rect 5228 -55206 5328 -54806
rect 8163 -54948 8261 -54943
rect 8162 -54949 14864 -54948
rect 8162 -55047 8163 -54949
rect 8261 -54953 14864 -54949
rect 8261 -55043 14769 -54953
rect 14859 -55043 14864 -54953
rect 8261 -55047 14864 -55043
rect 8162 -55048 14864 -55047
rect 8163 -55053 8261 -55048
rect -29235 -55370 -27536 -55206
rect -29235 -56652 -27620 -55370
rect -27556 -56652 -27536 -55370
rect -29235 -56806 -27536 -56652
rect -27129 -55370 -25430 -55206
rect -27129 -56652 -25514 -55370
rect -25450 -55954 -25430 -55370
rect -25023 -55370 -23324 -55206
rect -25023 -55954 -23408 -55370
rect -25450 -56054 -23408 -55954
rect -25450 -56652 -25430 -56054
rect -27129 -56806 -25430 -56652
rect -25023 -56652 -23408 -56054
rect -23344 -55954 -23324 -55370
rect -22917 -55370 -21218 -55206
rect -22917 -55954 -21302 -55370
rect -23344 -56054 -21302 -55954
rect -23344 -56652 -23324 -56054
rect -25023 -56806 -23324 -56652
rect -22917 -56652 -21302 -56054
rect -21238 -55954 -21218 -55370
rect -20811 -55370 -19112 -55206
rect -20811 -55954 -19196 -55370
rect -21238 -56054 -19196 -55954
rect -21238 -56652 -21218 -56054
rect -22917 -56806 -21218 -56652
rect -20811 -56652 -19196 -56054
rect -19132 -56652 -19112 -55370
rect -20811 -56806 -19112 -56652
rect -18705 -55370 -17006 -55206
rect -18705 -56652 -17090 -55370
rect -17026 -55976 -17006 -55370
rect -16599 -55370 -14900 -55206
rect -16599 -55976 -14984 -55370
rect -17026 -56076 -14984 -55976
rect -17026 -56652 -17006 -56076
rect -18705 -56806 -17006 -56652
rect -16599 -56652 -14984 -56076
rect -14920 -55976 -14900 -55370
rect -14493 -55370 -12794 -55206
rect -14493 -55976 -12878 -55370
rect -14920 -56076 -12878 -55976
rect -14920 -56652 -14900 -56076
rect -16599 -56806 -14900 -56652
rect -14493 -56652 -12878 -56076
rect -12814 -55976 -12794 -55370
rect -12387 -55370 -10688 -55206
rect -12387 -55976 -10772 -55370
rect -12814 -56076 -10772 -55976
rect -12814 -56652 -12794 -56076
rect -14493 -56806 -12794 -56652
rect -12387 -56652 -10772 -56076
rect -10708 -55976 -10688 -55370
rect -10281 -55370 -8582 -55206
rect -10281 -55976 -8666 -55370
rect -10708 -56076 -8666 -55976
rect -10708 -56652 -10688 -56076
rect -12387 -56806 -10688 -56652
rect -10281 -56652 -8666 -56076
rect -8602 -55976 -8582 -55370
rect -8175 -55370 -6476 -55206
rect -8175 -55976 -6560 -55370
rect -8602 -56076 -6560 -55976
rect -8602 -56652 -8582 -56076
rect -10281 -56806 -8582 -56652
rect -8175 -56652 -6560 -56076
rect -6496 -55976 -6476 -55370
rect -6069 -55370 -4370 -55206
rect -6069 -55976 -4454 -55370
rect -6496 -56076 -4454 -55976
rect -6496 -56652 -6476 -56076
rect -8175 -56806 -6476 -56652
rect -6069 -56652 -4454 -56076
rect -4390 -56652 -4370 -55370
rect -6069 -56806 -4370 -56652
rect -3963 -55370 -2264 -55206
rect -3963 -56652 -2348 -55370
rect -2284 -55950 -2264 -55370
rect -1857 -55370 -158 -55206
rect -1857 -55950 -242 -55370
rect -2284 -56050 -242 -55950
rect -2284 -56652 -2264 -56050
rect -3963 -56806 -2264 -56652
rect -1857 -56652 -242 -56050
rect -178 -55950 -158 -55370
rect 249 -55370 1948 -55206
rect 249 -55950 1864 -55370
rect -178 -56050 1864 -55950
rect -178 -56652 -158 -56050
rect -1857 -56806 -158 -56652
rect 249 -56652 1864 -56050
rect 1928 -55950 1948 -55370
rect 2355 -55370 4054 -55206
rect 2355 -55950 3970 -55370
rect 1928 -56050 3970 -55950
rect 1928 -56652 1948 -56050
rect 249 -56806 1948 -56652
rect 2355 -56652 3970 -56050
rect 4034 -55950 4054 -55370
rect 4461 -55370 6160 -55206
rect 4461 -55950 6076 -55370
rect 4034 -56050 6076 -55950
rect 4034 -56652 4054 -56050
rect 2355 -56806 4054 -56652
rect 4461 -56652 6076 -56050
rect 6140 -56652 6160 -55370
rect 4461 -56806 6160 -56652
rect 6567 -55370 8266 -55206
rect 6567 -56652 8182 -55370
rect 8246 -56334 8266 -55370
rect 8246 -56339 14874 -56334
rect 8246 -56429 14779 -56339
rect 14869 -56429 14874 -56339
rect 8246 -56434 14874 -56429
rect 8246 -56652 8266 -56434
rect 6567 -56806 8266 -56652
rect 9350 -56724 9452 -56700
rect -26392 -57206 -26292 -56806
rect -24286 -57206 -24186 -56806
rect -22156 -57206 -22056 -56806
rect -20012 -57206 -19912 -56806
rect -3278 -57206 -3178 -56806
rect -1156 -57206 -1056 -56806
rect 1010 -57206 1110 -56806
rect 3060 -57206 3160 -56806
rect 5228 -57206 5328 -56806
rect -29235 -57370 -27536 -57206
rect -29235 -58652 -27620 -57370
rect -27556 -58652 -27536 -57370
rect -29235 -58806 -27536 -58652
rect -27129 -57370 -25430 -57206
rect -27129 -58652 -25514 -57370
rect -25450 -57954 -25430 -57370
rect -25023 -57370 -23324 -57206
rect -25023 -57954 -23408 -57370
rect -25450 -58054 -23408 -57954
rect -25450 -58652 -25430 -58054
rect -27129 -58806 -25430 -58652
rect -25023 -58652 -23408 -58054
rect -23344 -57930 -23324 -57370
rect -22917 -57370 -21218 -57206
rect -22917 -57930 -21302 -57370
rect -23344 -58030 -21302 -57930
rect -23344 -58652 -23324 -58030
rect -25023 -58806 -23324 -58652
rect -22917 -58652 -21302 -58030
rect -21238 -57930 -21218 -57370
rect -20811 -57370 -19112 -57206
rect -20811 -57930 -19196 -57370
rect -21238 -58030 -19196 -57930
rect -21238 -58652 -21218 -58030
rect -22917 -58806 -21218 -58652
rect -20811 -58652 -19196 -58030
rect -19132 -57930 -19112 -57370
rect -18705 -57370 -17006 -57206
rect -18705 -57930 -17090 -57370
rect -19132 -58030 -17090 -57930
rect -19132 -58652 -19112 -58030
rect -20811 -58806 -19112 -58652
rect -18705 -58652 -17090 -58030
rect -17026 -57930 -17006 -57370
rect -16599 -57370 -14900 -57206
rect -16599 -57930 -14984 -57370
rect -17026 -58030 -14984 -57930
rect -17026 -58652 -17006 -58030
rect -18705 -58806 -17006 -58652
rect -16599 -58652 -14984 -58030
rect -14920 -57930 -14900 -57370
rect -14493 -57370 -12794 -57206
rect -14493 -57930 -12878 -57370
rect -14920 -58030 -12878 -57930
rect -14920 -58652 -14900 -58030
rect -16599 -58806 -14900 -58652
rect -14493 -58652 -12878 -58030
rect -12814 -57930 -12794 -57370
rect -12387 -57370 -10688 -57206
rect -12387 -57930 -10772 -57370
rect -12814 -58030 -10772 -57930
rect -12814 -58652 -12794 -58030
rect -14493 -58806 -12794 -58652
rect -12387 -58652 -10772 -58030
rect -10708 -57930 -10688 -57370
rect -10281 -57370 -8582 -57206
rect -10281 -57930 -8666 -57370
rect -10708 -58030 -8666 -57930
rect -10708 -58652 -10688 -58030
rect -12387 -58806 -10688 -58652
rect -10281 -58652 -8666 -58030
rect -8602 -57930 -8582 -57370
rect -8175 -57370 -6476 -57206
rect -8175 -57930 -6560 -57370
rect -8602 -58030 -6560 -57930
rect -8602 -58652 -8582 -58030
rect -10281 -58806 -8582 -58652
rect -8175 -58652 -6560 -58030
rect -6496 -57930 -6476 -57370
rect -6069 -57370 -4370 -57206
rect -6069 -57930 -4454 -57370
rect -6496 -58030 -4454 -57930
rect -6496 -58652 -6476 -58030
rect -8175 -58806 -6476 -58652
rect -6069 -58652 -4454 -58030
rect -4390 -57930 -4370 -57370
rect -3963 -57370 -2264 -57206
rect -3963 -57930 -2348 -57370
rect -4390 -58030 -2348 -57930
rect -4390 -58652 -4370 -58030
rect -6069 -58806 -4370 -58652
rect -3963 -58652 -2348 -58030
rect -2284 -57930 -2264 -57370
rect -1857 -57370 -158 -57206
rect -1857 -57930 -242 -57370
rect -2284 -58030 -242 -57930
rect -2284 -58652 -2264 -58030
rect -3963 -58806 -2264 -58652
rect -1857 -58652 -242 -58030
rect -178 -57930 -158 -57370
rect 249 -57370 1948 -57206
rect 249 -57930 1864 -57370
rect -178 -58030 1864 -57930
rect -178 -58652 -158 -58030
rect -1857 -58806 -158 -58652
rect 249 -58652 1864 -58030
rect 1928 -57930 1948 -57370
rect 2355 -57370 4054 -57206
rect 2355 -57930 3970 -57370
rect 1928 -58030 3970 -57930
rect 1928 -58652 1948 -58030
rect 249 -58806 1948 -58652
rect 2355 -58652 3970 -58030
rect 4034 -57930 4054 -57370
rect 4461 -57370 6160 -57206
rect 4461 -57930 6076 -57370
rect 4034 -58030 6076 -57930
rect 4034 -58652 4054 -58030
rect 2355 -58806 4054 -58652
rect 4461 -58652 6076 -58030
rect 6140 -58652 6160 -57370
rect 4461 -58806 6160 -58652
rect 6567 -57370 8266 -57206
rect 6567 -58652 8182 -57370
rect 8246 -57614 8266 -57370
rect 9350 -57518 9372 -56724
rect 9436 -57518 9452 -56724
rect 9350 -57536 9452 -57518
rect 12504 -57532 12604 -57512
rect 12504 -57592 12524 -57532
rect 12584 -57592 12604 -57532
rect 8246 -57635 10734 -57614
rect 8246 -57695 10652 -57635
rect 10712 -57695 10734 -57635
rect 8246 -57712 10734 -57695
rect 8246 -57714 10652 -57712
rect 8246 -58652 8266 -57714
rect 12504 -58183 12604 -57592
rect 12504 -58243 12526 -58183
rect 12586 -58243 12604 -58183
rect 10276 -58408 12130 -58390
rect 10276 -58514 10294 -58408
rect 12110 -58514 12130 -58408
rect 10276 -58528 12130 -58514
rect 6567 -58806 8266 -58652
rect -26392 -59206 -26292 -58806
rect -24286 -59206 -24186 -58806
rect -22166 -59206 -22066 -58806
rect -20060 -59206 -19960 -58806
rect -17954 -59206 -17854 -58806
rect -15848 -59206 -15748 -58806
rect -13742 -59206 -13642 -58806
rect -11636 -59206 -11536 -58806
rect -9530 -59206 -9430 -58806
rect -7424 -59206 -7324 -58806
rect -5318 -59206 -5218 -58806
rect -3212 -59206 -3112 -58806
rect -1106 -59206 -1006 -58806
rect 1000 -59206 1100 -58806
rect 3106 -59206 3206 -58806
rect 5228 -59206 5328 -58806
rect -29235 -59370 -27536 -59206
rect -29235 -60652 -27620 -59370
rect -27556 -60652 -27536 -59370
rect -29235 -60806 -27536 -60652
rect -27129 -59370 -25430 -59206
rect -27129 -60652 -25514 -59370
rect -25450 -59946 -25430 -59370
rect -25023 -59370 -23324 -59206
rect -25023 -59946 -23408 -59370
rect -25450 -60046 -23408 -59946
rect -25450 -60652 -25430 -60046
rect -27129 -60806 -25430 -60652
rect -25023 -60652 -23408 -60046
rect -23344 -59946 -23324 -59370
rect -22917 -59370 -21218 -59206
rect -22917 -59946 -21302 -59370
rect -23344 -60046 -21302 -59946
rect -23344 -60652 -23324 -60046
rect -25023 -60806 -23324 -60652
rect -22917 -60652 -21302 -60046
rect -21238 -59946 -21218 -59370
rect -20811 -59370 -19112 -59206
rect -20811 -59946 -19196 -59370
rect -21238 -60046 -19196 -59946
rect -21238 -60652 -21218 -60046
rect -22917 -60806 -21218 -60652
rect -20811 -60652 -19196 -60046
rect -19132 -59946 -19112 -59370
rect -18705 -59370 -17006 -59206
rect -18705 -59946 -17090 -59370
rect -19132 -60046 -17090 -59946
rect -19132 -60652 -19112 -60046
rect -20811 -60806 -19112 -60652
rect -18705 -60652 -17090 -60046
rect -17026 -59946 -17006 -59370
rect -16599 -59370 -14900 -59206
rect -16599 -59946 -14984 -59370
rect -17026 -60046 -14984 -59946
rect -17026 -60652 -17006 -60046
rect -18705 -60806 -17006 -60652
rect -16599 -60652 -14984 -60046
rect -14920 -59946 -14900 -59370
rect -14493 -59370 -12794 -59206
rect -14493 -59946 -12878 -59370
rect -14920 -60046 -12878 -59946
rect -14920 -60652 -14900 -60046
rect -16599 -60806 -14900 -60652
rect -14493 -60652 -12878 -60046
rect -12814 -59946 -12794 -59370
rect -12387 -59370 -10688 -59206
rect -12387 -59946 -10772 -59370
rect -12814 -60046 -10772 -59946
rect -12814 -60652 -12794 -60046
rect -14493 -60806 -12794 -60652
rect -12387 -60652 -10772 -60046
rect -10708 -59946 -10688 -59370
rect -10281 -59370 -8582 -59206
rect -10281 -59946 -8666 -59370
rect -10708 -60046 -8666 -59946
rect -10708 -60652 -10688 -60046
rect -12387 -60806 -10688 -60652
rect -10281 -60652 -8666 -60046
rect -8602 -59946 -8582 -59370
rect -8175 -59370 -6476 -59206
rect -8175 -59946 -6560 -59370
rect -8602 -60046 -6560 -59946
rect -8602 -60652 -8582 -60046
rect -10281 -60806 -8582 -60652
rect -8175 -60652 -6560 -60046
rect -6496 -59946 -6476 -59370
rect -6069 -59370 -4370 -59206
rect -6069 -59946 -4454 -59370
rect -6496 -60046 -4454 -59946
rect -6496 -60652 -6476 -60046
rect -8175 -60806 -6476 -60652
rect -6069 -60652 -4454 -60046
rect -4390 -59946 -4370 -59370
rect -3963 -59370 -2264 -59206
rect -3963 -59946 -2348 -59370
rect -4390 -60046 -2348 -59946
rect -4390 -60652 -4370 -60046
rect -6069 -60806 -4370 -60652
rect -3963 -60652 -2348 -60046
rect -2284 -59946 -2264 -59370
rect -1857 -59370 -158 -59206
rect -1857 -59946 -242 -59370
rect -2284 -60046 -242 -59946
rect -2284 -60652 -2264 -60046
rect -3963 -60806 -2264 -60652
rect -1857 -60652 -242 -60046
rect -178 -59946 -158 -59370
rect 249 -59370 1948 -59206
rect 249 -59946 1864 -59370
rect -178 -60046 1864 -59946
rect -178 -60652 -158 -60046
rect -1857 -60806 -158 -60652
rect 249 -60652 1864 -60046
rect 1928 -59946 1948 -59370
rect 2355 -59370 4054 -59206
rect 2355 -59946 3970 -59370
rect 1928 -60046 3970 -59946
rect 1928 -60652 1948 -60046
rect 249 -60806 1948 -60652
rect 2355 -60652 3970 -60046
rect 4034 -59946 4054 -59370
rect 4461 -59370 6160 -59206
rect 4461 -59946 6076 -59370
rect 4034 -60046 6076 -59946
rect 4034 -60652 4054 -60046
rect 2355 -60806 4054 -60652
rect 4461 -60652 6076 -60046
rect 6140 -60652 6160 -59370
rect 4461 -60806 6160 -60652
rect 6567 -59370 8266 -59206
rect 6567 -60652 8182 -59370
rect 8246 -60652 8266 -59370
rect 6567 -60806 8266 -60652
rect -29235 -61370 -27536 -61206
rect -29235 -62652 -27620 -61370
rect -27556 -62652 -27536 -61370
rect -29235 -62806 -27536 -62652
rect -27129 -61370 -25430 -61206
rect -27129 -62652 -25514 -61370
rect -25450 -61936 -25430 -61370
rect -25023 -61370 -23324 -61206
rect -25023 -61936 -23408 -61370
rect -25450 -62040 -23408 -61936
rect -25450 -62652 -25430 -62040
rect -27129 -62806 -25430 -62652
rect -25023 -62652 -23408 -62040
rect -23344 -62652 -23324 -61370
rect -25023 -62806 -23324 -62652
rect -22917 -61370 -21218 -61206
rect -22917 -62652 -21302 -61370
rect -21238 -62652 -21218 -61370
rect -22917 -62806 -21218 -62652
rect -20811 -61370 -19112 -61206
rect -20811 -62652 -19196 -61370
rect -19132 -62652 -19112 -61370
rect -20811 -62806 -19112 -62652
rect -18705 -61370 -17006 -61206
rect -18705 -62652 -17090 -61370
rect -17026 -62652 -17006 -61370
rect -18705 -62806 -17006 -62652
rect -16599 -61370 -14900 -61206
rect -16599 -62652 -14984 -61370
rect -14920 -62652 -14900 -61370
rect -16599 -62806 -14900 -62652
rect -14493 -61370 -12794 -61206
rect -14493 -62652 -12878 -61370
rect -12814 -62652 -12794 -61370
rect -14493 -62806 -12794 -62652
rect -12387 -61370 -10688 -61206
rect -12387 -62652 -10772 -61370
rect -10708 -62652 -10688 -61370
rect -12387 -62806 -10688 -62652
rect -10281 -61370 -8582 -61206
rect -10281 -62652 -8666 -61370
rect -8602 -62652 -8582 -61370
rect -10281 -62806 -8582 -62652
rect -8175 -61370 -6476 -61206
rect -8175 -62652 -6560 -61370
rect -6496 -62652 -6476 -61370
rect -8175 -62806 -6476 -62652
rect -6069 -61370 -4370 -61206
rect -6069 -62652 -4454 -61370
rect -4390 -62652 -4370 -61370
rect -6069 -62806 -4370 -62652
rect -3963 -61370 -2264 -61206
rect -3963 -62652 -2348 -61370
rect -2284 -62652 -2264 -61370
rect -3963 -62806 -2264 -62652
rect -1857 -61370 -158 -61206
rect -1857 -62652 -242 -61370
rect -178 -62652 -158 -61370
rect -1857 -62806 -158 -62652
rect 249 -61370 1948 -61206
rect 249 -62652 1864 -61370
rect 1928 -62652 1948 -61370
rect 249 -62806 1948 -62652
rect 2355 -61370 4054 -61206
rect 2355 -62652 3970 -61370
rect 4034 -62652 4054 -61370
rect 2355 -62806 4054 -62652
rect 4461 -61370 6160 -61206
rect 4461 -62652 6076 -61370
rect 6140 -62652 6160 -61370
rect 4461 -62806 6160 -62652
rect 6567 -61370 8266 -61206
rect 6567 -62652 8182 -61370
rect 8246 -62652 8266 -61370
rect 6567 -62806 8266 -62652
rect -9938 -63001 -9838 -63000
rect -14752 -63009 -14652 -63008
rect -16848 -63011 -16748 -63010
rect -18964 -63015 -18864 -63014
rect -18969 -63113 -18963 -63015
rect -18865 -63113 -18859 -63015
rect -16853 -63109 -16847 -63011
rect -16749 -63109 -16743 -63011
rect -14757 -63107 -14751 -63009
rect -14653 -63107 -14647 -63009
rect -10592 -63011 -10492 -63010
rect -12628 -63019 -12528 -63018
rect -25200 -63278 -25100 -63272
rect -18964 -63326 -18864 -63113
rect -16848 -63310 -16748 -63109
rect -27588 -64532 -26968 -64527
rect -27588 -64832 -27578 -64532
rect -26978 -64832 -26968 -64532
rect -27588 -64837 -26968 -64832
rect -26076 -64532 -25456 -64527
rect -26076 -64832 -26066 -64532
rect -25466 -64832 -25456 -64532
rect -26076 -64837 -25456 -64832
rect -27422 -65036 -25520 -65006
rect -27422 -65100 -27388 -65036
rect -25564 -65100 -25520 -65036
rect -27422 -65130 -25520 -65100
rect -25200 -65195 -25100 -63378
rect -21036 -63426 -18864 -63326
rect -17114 -63410 -16748 -63310
rect -23588 -64532 -22968 -64527
rect -23588 -64832 -23578 -64532
rect -22978 -64832 -22968 -64532
rect -23588 -64837 -22968 -64832
rect -22076 -64532 -21456 -64527
rect -22076 -64832 -22066 -64532
rect -21466 -64832 -21456 -64532
rect -22076 -64837 -21456 -64832
rect -23422 -65036 -21520 -65006
rect -23422 -65100 -23388 -65036
rect -21564 -65100 -21520 -65036
rect -23422 -65130 -21520 -65100
rect -25200 -65285 -25195 -65195
rect -25105 -65285 -25100 -65195
rect -25200 -65290 -25100 -65285
rect -21036 -65197 -20936 -63426
rect -19588 -64532 -18968 -64527
rect -19588 -64832 -19578 -64532
rect -18978 -64832 -18968 -64532
rect -19588 -64837 -18968 -64832
rect -18076 -64532 -17456 -64527
rect -18076 -64832 -18066 -64532
rect -17466 -64832 -17456 -64532
rect -18076 -64837 -17456 -64832
rect -19422 -65036 -17520 -65006
rect -19422 -65100 -19388 -65036
rect -17564 -65100 -17520 -65036
rect -19422 -65130 -17520 -65100
rect -21036 -65287 -21031 -65197
rect -20941 -65287 -20936 -65197
rect -21036 -65292 -20936 -65287
rect -17114 -65197 -17014 -63410
rect -14752 -63634 -14652 -63107
rect -12633 -63117 -12627 -63019
rect -12529 -63117 -12523 -63019
rect -10597 -63109 -10591 -63011
rect -10493 -63109 -10487 -63011
rect -9943 -63099 -9937 -63001
rect -9839 -63099 -9833 -63001
rect -8496 -63019 -8396 -63018
rect -17114 -65287 -17109 -65197
rect -17019 -65287 -17014 -65197
rect -17114 -65292 -17014 -65287
rect -16092 -63734 -14652 -63634
rect -16092 -65197 -15992 -63734
rect -12628 -64188 -12528 -63117
rect -10592 -64004 -10492 -63109
rect -9938 -63640 -9838 -63099
rect -8501 -63117 -8495 -63019
rect -8397 -63117 -8391 -63019
rect -7927 -63022 -7829 -63017
rect -7928 -63023 4110 -63022
rect -8496 -63322 -8396 -63117
rect -7928 -63121 -7927 -63023
rect -7829 -63121 4110 -63023
rect -7928 -63122 4110 -63121
rect -7927 -63127 -7829 -63122
rect -8496 -63422 56 -63322
rect -9938 -63740 -4002 -63640
rect -10592 -64026 -9114 -64004
rect -10592 -64086 -9198 -64026
rect -9138 -64086 -9114 -64026
rect -10592 -64104 -9114 -64086
rect -12628 -64288 -7874 -64188
rect -15588 -64532 -14968 -64527
rect -15588 -64832 -15578 -64532
rect -14978 -64832 -14968 -64532
rect -15588 -64837 -14968 -64832
rect -14076 -64532 -13456 -64527
rect -14076 -64832 -14066 -64532
rect -13466 -64832 -13456 -64532
rect -14076 -64837 -13456 -64832
rect -11588 -64532 -10968 -64527
rect -11588 -64832 -11578 -64532
rect -10978 -64832 -10968 -64532
rect -11588 -64837 -10968 -64832
rect -10076 -64532 -9456 -64527
rect -10076 -64832 -10066 -64532
rect -9466 -64832 -9456 -64532
rect -10076 -64837 -9456 -64832
rect -15422 -65036 -13520 -65006
rect -15422 -65100 -15388 -65036
rect -13564 -65100 -13520 -65036
rect -15422 -65130 -13520 -65100
rect -11422 -65036 -9520 -65006
rect -11422 -65100 -11388 -65036
rect -9564 -65100 -9520 -65036
rect -11422 -65130 -9520 -65100
rect -16092 -65287 -16087 -65197
rect -15997 -65287 -15992 -65197
rect -16092 -65292 -15992 -65287
rect -7974 -65214 -7874 -64288
rect -7588 -64532 -6968 -64527
rect -7588 -64832 -7578 -64532
rect -6978 -64832 -6968 -64532
rect -7588 -64837 -6968 -64832
rect -6076 -64532 -5456 -64527
rect -6076 -64832 -6066 -64532
rect -5466 -64832 -5456 -64532
rect -6076 -64837 -5456 -64832
rect -7422 -65036 -5520 -65006
rect -7422 -65100 -7388 -65036
rect -5564 -65100 -5520 -65036
rect -7422 -65130 -5520 -65100
rect -7974 -65274 -7956 -65214
rect -7896 -65274 -7874 -65214
rect -7974 -65298 -7874 -65274
rect -4102 -65197 -4002 -63740
rect -3588 -64532 -2968 -64527
rect -3588 -64832 -3578 -64532
rect -2978 -64832 -2968 -64532
rect -3588 -64837 -2968 -64832
rect -2076 -64532 -1456 -64527
rect -2076 -64832 -2066 -64532
rect -1466 -64832 -1456 -64532
rect -2076 -64837 -1456 -64832
rect -3422 -65036 -1520 -65006
rect -3422 -65100 -3388 -65036
rect -1564 -65100 -1520 -65036
rect -3422 -65130 -1520 -65100
rect -4102 -65287 -4097 -65197
rect -4007 -65287 -4002 -65197
rect -4102 -65292 -4002 -65287
rect -44 -65201 56 -63422
rect 412 -64532 1032 -64527
rect 412 -64832 422 -64532
rect 1022 -64832 1032 -64532
rect 412 -64837 1032 -64832
rect 1924 -64532 2544 -64527
rect 1924 -64832 1934 -64532
rect 2534 -64832 2544 -64532
rect 1924 -64837 2544 -64832
rect 578 -65036 2480 -65006
rect 578 -65100 612 -65036
rect 2436 -65100 2480 -65036
rect 578 -65130 2480 -65100
rect -44 -65291 -39 -65201
rect 51 -65291 56 -65201
rect -44 -65296 56 -65291
rect 4010 -65199 4110 -63122
rect 4412 -64532 5032 -64527
rect 4412 -64832 4422 -64532
rect 5022 -64832 5032 -64532
rect 4412 -64837 5032 -64832
rect 5924 -64532 6544 -64527
rect 5924 -64832 5934 -64532
rect 6534 -64832 6544 -64532
rect 5924 -64837 6544 -64832
rect 4578 -65036 6480 -65006
rect 4578 -65100 4612 -65036
rect 6436 -65100 6480 -65036
rect 4578 -65130 6480 -65100
rect 4010 -65289 4015 -65199
rect 4105 -65289 4110 -65199
rect 4010 -65294 4110 -65289
rect 12504 -65426 12604 -58243
rect 17326 -58454 49412 -58408
rect 17326 -58608 17372 -58454
rect 49372 -58608 49412 -58454
rect 17326 -58654 49412 -58608
rect 13218 -58794 13838 -58789
rect 13218 -59094 13228 -58794
rect 13828 -59094 13838 -58794
rect 13218 -59099 13838 -59094
rect 49650 -58794 50270 -58789
rect 49650 -59094 49660 -58794
rect 50260 -59094 50270 -58794
rect 49650 -59099 50270 -59094
rect 52310 -59666 52510 -42022
rect 58424 -42208 58524 -42202
rect 53290 -42560 53296 -42460
rect 53396 -42560 53402 -42460
rect 54180 -42471 54282 -42462
rect 54180 -42553 54195 -42471
rect 54259 -42476 54282 -42471
rect 54260 -42548 54282 -42476
rect 54259 -42553 54282 -42548
rect 53296 -43828 53396 -42560
rect 54180 -42562 54282 -42553
rect 55276 -42466 55382 -42458
rect 55276 -42471 55300 -42466
rect 55276 -42553 55295 -42471
rect 55276 -42558 55300 -42553
rect 55370 -42558 55382 -42466
rect 55276 -42566 55382 -42558
rect 56042 -42573 56142 -42572
rect 56037 -42671 56043 -42573
rect 56141 -42671 56147 -42573
rect 57946 -42575 58046 -42574
rect 56042 -42672 56142 -42671
rect 57941 -42673 57947 -42575
rect 58045 -42673 58051 -42575
rect 57946 -42674 58046 -42673
rect 55814 -43278 58278 -43273
rect 55814 -43584 55824 -43278
rect 58268 -43584 58278 -43278
rect 55814 -43589 58278 -43584
rect 58424 -43828 58524 -42308
rect 53296 -43928 58524 -43828
rect -26472 -65446 12604 -65426
rect -26472 -65506 -26448 -65446
rect -26388 -65506 -22448 -65446
rect -22388 -65506 -18450 -65446
rect -18390 -65506 -14450 -65446
rect -14390 -65506 -10450 -65446
rect -10390 -65506 -6448 -65446
rect -6388 -65506 -2452 -65446
rect -2392 -65506 1552 -65446
rect 1612 -65506 5554 -65446
rect 5614 -65506 12604 -65446
rect -26472 -65526 12604 -65506
rect 12962 -59714 52510 -59666
rect 12962 -59774 13016 -59714
rect 13076 -59774 52510 -59714
rect 12962 -59866 52510 -59774
rect -28296 -67920 5506 -67902
rect -28296 -67980 -26578 -67920
rect -26518 -67980 -22578 -67920
rect -22518 -67980 -18578 -67920
rect -18518 -67980 -14578 -67920
rect -14518 -67980 -10578 -67920
rect -10518 -67980 -6578 -67920
rect -6518 -67980 -2578 -67920
rect -2518 -67980 1422 -67920
rect 1482 -67922 5506 -67920
rect 1482 -67980 5422 -67922
rect -28296 -67982 5422 -67980
rect 5482 -67982 5506 -67922
rect -28296 -68002 5506 -67982
rect -25254 -68952 -25154 -68924
rect -25254 -69012 -25232 -68952
rect -25172 -69012 -25154 -68952
rect -27466 -69154 -25688 -69122
rect -27466 -69222 -27430 -69154
rect -25722 -69222 -25688 -69154
rect -27466 -69252 -25688 -69222
rect -27588 -69404 -26968 -69399
rect -27588 -69704 -27578 -69404
rect -26978 -69704 -26968 -69404
rect -27588 -69709 -26968 -69704
rect -26076 -69404 -25456 -69399
rect -26076 -69704 -26066 -69404
rect -25466 -69704 -25456 -69404
rect -26076 -69709 -25456 -69704
rect -27588 -70492 -26968 -70487
rect -27588 -70792 -27578 -70492
rect -26978 -70792 -26968 -70492
rect -27588 -70797 -26968 -70792
rect -26076 -70492 -25456 -70487
rect -26076 -70792 -26066 -70492
rect -25466 -70792 -25456 -70492
rect -26076 -70797 -25456 -70792
rect -27466 -70974 -25688 -70944
rect -27466 -71042 -27430 -70974
rect -25722 -71042 -25688 -70974
rect -27466 -71074 -25688 -71042
rect -25254 -72106 -25154 -69012
rect -21254 -68952 -21154 -68924
rect -21254 -69012 -21232 -68952
rect -21172 -69012 -21154 -68952
rect -23466 -69154 -21688 -69122
rect -23466 -69222 -23430 -69154
rect -21722 -69222 -21688 -69154
rect -23466 -69252 -21688 -69222
rect -23588 -69404 -22968 -69399
rect -23588 -69704 -23578 -69404
rect -22978 -69704 -22968 -69404
rect -23588 -69709 -22968 -69704
rect -22076 -69404 -21456 -69399
rect -22076 -69704 -22066 -69404
rect -21466 -69704 -21456 -69404
rect -22076 -69709 -21456 -69704
rect -23588 -70492 -22968 -70487
rect -23588 -70792 -23578 -70492
rect -22978 -70792 -22968 -70492
rect -23588 -70797 -22968 -70792
rect -22076 -70492 -21456 -70487
rect -22076 -70792 -22066 -70492
rect -21466 -70792 -21456 -70492
rect -22076 -70797 -21456 -70792
rect -23466 -70974 -21688 -70944
rect -23466 -71042 -23430 -70974
rect -21722 -71042 -21688 -70974
rect -23466 -71074 -21688 -71042
rect -25254 -72166 -25238 -72106
rect -25178 -72166 -25154 -72106
rect -25254 -72192 -25154 -72166
rect -21254 -72106 -21154 -69012
rect -17254 -68952 -17154 -68924
rect -17254 -69012 -17232 -68952
rect -17172 -69012 -17154 -68952
rect -19466 -69154 -17688 -69122
rect -19466 -69222 -19430 -69154
rect -17722 -69222 -17688 -69154
rect -19466 -69252 -17688 -69222
rect -19588 -69404 -18968 -69399
rect -19588 -69704 -19578 -69404
rect -18978 -69704 -18968 -69404
rect -19588 -69709 -18968 -69704
rect -18076 -69404 -17456 -69399
rect -18076 -69704 -18066 -69404
rect -17466 -69704 -17456 -69404
rect -18076 -69709 -17456 -69704
rect -19588 -70492 -18968 -70487
rect -19588 -70792 -19578 -70492
rect -18978 -70792 -18968 -70492
rect -19588 -70797 -18968 -70792
rect -18076 -70492 -17456 -70487
rect -18076 -70792 -18066 -70492
rect -17466 -70792 -17456 -70492
rect -18076 -70797 -17456 -70792
rect -19466 -70974 -17688 -70944
rect -19466 -71042 -19430 -70974
rect -17722 -71042 -17688 -70974
rect -19466 -71074 -17688 -71042
rect -21254 -72166 -21238 -72106
rect -21178 -72166 -21154 -72106
rect -21254 -72192 -21154 -72166
rect -17254 -72106 -17154 -69012
rect -13254 -68952 -13154 -68924
rect -13254 -69012 -13232 -68952
rect -13172 -69012 -13154 -68952
rect -15466 -69154 -13688 -69122
rect -15466 -69222 -15430 -69154
rect -13722 -69222 -13688 -69154
rect -15466 -69252 -13688 -69222
rect -15588 -69404 -14968 -69399
rect -15588 -69704 -15578 -69404
rect -14978 -69704 -14968 -69404
rect -15588 -69709 -14968 -69704
rect -14076 -69404 -13456 -69399
rect -14076 -69704 -14066 -69404
rect -13466 -69704 -13456 -69404
rect -14076 -69709 -13456 -69704
rect -15588 -70492 -14968 -70487
rect -15588 -70792 -15578 -70492
rect -14978 -70792 -14968 -70492
rect -15588 -70797 -14968 -70792
rect -14076 -70492 -13456 -70487
rect -14076 -70792 -14066 -70492
rect -13466 -70792 -13456 -70492
rect -14076 -70797 -13456 -70792
rect -15466 -70974 -13688 -70944
rect -15466 -71042 -15430 -70974
rect -13722 -71042 -13688 -70974
rect -15466 -71074 -13688 -71042
rect -17254 -72166 -17238 -72106
rect -17178 -72166 -17154 -72106
rect -17254 -72192 -17154 -72166
rect -13254 -72106 -13154 -69012
rect -9254 -68952 -9154 -68924
rect -9254 -69012 -9232 -68952
rect -9172 -69012 -9154 -68952
rect -11466 -69154 -9688 -69122
rect -11466 -69222 -11430 -69154
rect -9722 -69222 -9688 -69154
rect -11466 -69252 -9688 -69222
rect -11588 -69404 -10968 -69399
rect -11588 -69704 -11578 -69404
rect -10978 -69704 -10968 -69404
rect -11588 -69709 -10968 -69704
rect -10076 -69404 -9456 -69399
rect -10076 -69704 -10066 -69404
rect -9466 -69704 -9456 -69404
rect -10076 -69709 -9456 -69704
rect -11588 -70492 -10968 -70487
rect -11588 -70792 -11578 -70492
rect -10978 -70792 -10968 -70492
rect -11588 -70797 -10968 -70792
rect -10076 -70492 -9456 -70487
rect -10076 -70792 -10066 -70492
rect -9466 -70792 -9456 -70492
rect -10076 -70797 -9456 -70792
rect -11466 -70974 -9688 -70944
rect -11466 -71042 -11430 -70974
rect -9722 -71042 -9688 -70974
rect -11466 -71074 -9688 -71042
rect -13254 -72166 -13238 -72106
rect -13178 -72166 -13154 -72106
rect -13254 -72192 -13154 -72166
rect -9254 -72106 -9154 -69012
rect -5254 -68952 -5154 -68924
rect -5254 -69012 -5232 -68952
rect -5172 -69012 -5154 -68952
rect -7466 -69154 -5688 -69122
rect -7466 -69222 -7430 -69154
rect -5722 -69222 -5688 -69154
rect -7466 -69252 -5688 -69222
rect -7588 -69404 -6968 -69399
rect -7588 -69704 -7578 -69404
rect -6978 -69704 -6968 -69404
rect -7588 -69709 -6968 -69704
rect -6076 -69404 -5456 -69399
rect -6076 -69704 -6066 -69404
rect -5466 -69704 -5456 -69404
rect -6076 -69709 -5456 -69704
rect -7588 -70492 -6968 -70487
rect -7588 -70792 -7578 -70492
rect -6978 -70792 -6968 -70492
rect -7588 -70797 -6968 -70792
rect -6076 -70492 -5456 -70487
rect -6076 -70792 -6066 -70492
rect -5466 -70792 -5456 -70492
rect -6076 -70797 -5456 -70792
rect -7466 -70974 -5688 -70944
rect -7466 -71042 -7430 -70974
rect -5722 -71042 -5688 -70974
rect -7466 -71074 -5688 -71042
rect -9254 -72166 -9238 -72106
rect -9178 -72166 -9154 -72106
rect -9254 -72192 -9154 -72166
rect -5254 -72106 -5154 -69012
rect -1254 -68952 -1154 -68924
rect -1254 -69012 -1232 -68952
rect -1172 -69012 -1154 -68952
rect -3466 -69154 -1688 -69122
rect -3466 -69222 -3430 -69154
rect -1722 -69222 -1688 -69154
rect -3466 -69252 -1688 -69222
rect -3588 -69404 -2968 -69399
rect -3588 -69704 -3578 -69404
rect -2978 -69704 -2968 -69404
rect -3588 -69709 -2968 -69704
rect -2076 -69404 -1456 -69399
rect -2076 -69704 -2066 -69404
rect -1466 -69704 -1456 -69404
rect -2076 -69709 -1456 -69704
rect -3588 -70492 -2968 -70487
rect -3588 -70792 -3578 -70492
rect -2978 -70792 -2968 -70492
rect -3588 -70797 -2968 -70792
rect -2076 -70492 -1456 -70487
rect -2076 -70792 -2066 -70492
rect -1466 -70792 -1456 -70492
rect -2076 -70797 -1456 -70792
rect -3466 -70974 -1688 -70944
rect -3466 -71042 -3430 -70974
rect -1722 -71042 -1688 -70974
rect -3466 -71074 -1688 -71042
rect -5254 -72166 -5238 -72106
rect -5178 -72166 -5154 -72106
rect -5254 -72192 -5154 -72166
rect -1254 -72106 -1154 -69012
rect 2746 -68952 2846 -68924
rect 2746 -69012 2768 -68952
rect 2828 -69012 2846 -68952
rect 534 -69154 2312 -69122
rect 534 -69222 570 -69154
rect 2278 -69222 2312 -69154
rect 534 -69252 2312 -69222
rect 412 -69404 1032 -69399
rect 412 -69704 422 -69404
rect 1022 -69704 1032 -69404
rect 412 -69709 1032 -69704
rect 1924 -69404 2544 -69399
rect 1924 -69704 1934 -69404
rect 2534 -69704 2544 -69404
rect 1924 -69709 2544 -69704
rect 412 -70492 1032 -70487
rect 412 -70792 422 -70492
rect 1022 -70792 1032 -70492
rect 412 -70797 1032 -70792
rect 1924 -70492 2544 -70487
rect 1924 -70792 1934 -70492
rect 2534 -70792 2544 -70492
rect 1924 -70797 2544 -70792
rect 534 -70974 2312 -70944
rect 534 -71042 570 -70974
rect 2278 -71042 2312 -70974
rect 534 -71074 2312 -71042
rect -1254 -72166 -1238 -72106
rect -1178 -72166 -1154 -72106
rect -1254 -72192 -1154 -72166
rect 2746 -72106 2846 -69012
rect 6746 -68952 6846 -68924
rect 6746 -69012 6768 -68952
rect 6828 -69012 6846 -68952
rect 4534 -69154 6312 -69122
rect 4534 -69222 4570 -69154
rect 6278 -69222 6312 -69154
rect 4534 -69252 6312 -69222
rect 4412 -69404 5032 -69399
rect 4412 -69704 4422 -69404
rect 5022 -69704 5032 -69404
rect 4412 -69709 5032 -69704
rect 5924 -69404 6544 -69399
rect 5924 -69704 5934 -69404
rect 6534 -69704 6544 -69404
rect 5924 -69709 6544 -69704
rect 4412 -70492 5032 -70487
rect 4412 -70792 4422 -70492
rect 5022 -70792 5032 -70492
rect 4412 -70797 5032 -70792
rect 5924 -70492 6544 -70487
rect 5924 -70792 5934 -70492
rect 6534 -70792 6544 -70492
rect 5924 -70797 6544 -70792
rect 4534 -70974 6312 -70944
rect 4534 -71042 4570 -70974
rect 6278 -71042 6312 -70974
rect 4534 -71074 6312 -71042
rect 2746 -72166 2762 -72106
rect 2822 -72166 2846 -72106
rect 2746 -72192 2846 -72166
rect 6746 -72106 6846 -69012
rect 6746 -72166 6762 -72106
rect 6822 -72166 6846 -72106
rect 6746 -72192 6846 -72166
rect 12962 -72808 13162 -59866
rect 4844 -72864 13162 -72808
rect -28500 -72880 13162 -72864
rect -28500 -72882 -11094 -72880
rect -28500 -72942 -27094 -72882
rect -27034 -72942 -23094 -72882
rect -23034 -72942 -19094 -72882
rect -19034 -72942 -15094 -72882
rect -15034 -72940 -11094 -72882
rect -11034 -72882 13162 -72880
rect -11034 -72940 -7094 -72882
rect -15034 -72942 -7094 -72940
rect -7034 -72942 -3094 -72882
rect -3034 -72942 906 -72882
rect 966 -72942 4906 -72882
rect 4966 -72942 13162 -72882
rect -28500 -72964 13162 -72942
rect 4844 -73008 13162 -72964
rect -28238 -74866 4986 -74848
rect -28238 -74868 4908 -74866
rect -28238 -74870 -23092 -74868
rect -28238 -74930 -27092 -74870
rect -27032 -74928 -23092 -74870
rect -23032 -74928 -19092 -74868
rect -19032 -74928 -15092 -74868
rect -15032 -74870 -3092 -74868
rect -15032 -74928 -11092 -74870
rect -27032 -74930 -11092 -74928
rect -11032 -74930 -7092 -74870
rect -7032 -74928 -3092 -74870
rect -3032 -74928 908 -74868
rect 968 -74926 4908 -74868
rect 4968 -74926 4986 -74866
rect 968 -74928 4986 -74926
rect -7032 -74930 4986 -74928
rect -28238 -74948 4986 -74930
rect -27422 -75096 -25520 -75066
rect -27422 -75160 -27388 -75096
rect -25564 -75160 -25520 -75096
rect -27422 -75190 -25520 -75160
rect -23422 -75096 -21520 -75066
rect -23422 -75160 -23388 -75096
rect -21564 -75160 -21520 -75096
rect -23422 -75190 -21520 -75160
rect -19422 -75096 -17520 -75066
rect -19422 -75160 -19388 -75096
rect -17564 -75160 -17520 -75096
rect -19422 -75190 -17520 -75160
rect -15422 -75096 -13520 -75066
rect -15422 -75160 -15388 -75096
rect -13564 -75160 -13520 -75096
rect -15422 -75190 -13520 -75160
rect -11422 -75096 -9520 -75066
rect -11422 -75160 -11388 -75096
rect -9564 -75160 -9520 -75096
rect -11422 -75190 -9520 -75160
rect -7422 -75096 -5520 -75066
rect -7422 -75160 -7388 -75096
rect -5564 -75160 -5520 -75096
rect -7422 -75190 -5520 -75160
rect -3422 -75096 -1520 -75066
rect -3422 -75160 -3388 -75096
rect -1564 -75160 -1520 -75096
rect -3422 -75190 -1520 -75160
rect 578 -75096 2480 -75066
rect 578 -75160 612 -75096
rect 2436 -75160 2480 -75096
rect 578 -75190 2480 -75160
rect 4578 -75096 6480 -75066
rect 4578 -75160 4612 -75096
rect 6436 -75160 6480 -75096
rect 4578 -75190 6480 -75160
rect -27588 -75364 -26968 -75359
rect -27588 -75664 -27578 -75364
rect -26978 -75664 -26968 -75364
rect -27588 -75669 -26968 -75664
rect -26076 -75364 -25456 -75359
rect -26076 -75664 -26066 -75364
rect -25466 -75664 -25456 -75364
rect -26076 -75669 -25456 -75664
rect -23588 -75364 -22968 -75359
rect -23588 -75664 -23578 -75364
rect -22978 -75664 -22968 -75364
rect -23588 -75669 -22968 -75664
rect -22076 -75364 -21456 -75359
rect -22076 -75664 -22066 -75364
rect -21466 -75664 -21456 -75364
rect -22076 -75669 -21456 -75664
rect -19588 -75364 -18968 -75359
rect -19588 -75664 -19578 -75364
rect -18978 -75664 -18968 -75364
rect -19588 -75669 -18968 -75664
rect -18076 -75364 -17456 -75359
rect -18076 -75664 -18066 -75364
rect -17466 -75664 -17456 -75364
rect -18076 -75669 -17456 -75664
rect -15588 -75364 -14968 -75359
rect -15588 -75664 -15578 -75364
rect -14978 -75664 -14968 -75364
rect -15588 -75669 -14968 -75664
rect -14076 -75364 -13456 -75359
rect -14076 -75664 -14066 -75364
rect -13466 -75664 -13456 -75364
rect -14076 -75669 -13456 -75664
rect -11588 -75364 -10968 -75359
rect -11588 -75664 -11578 -75364
rect -10978 -75664 -10968 -75364
rect -11588 -75669 -10968 -75664
rect -10076 -75364 -9456 -75359
rect -10076 -75664 -10066 -75364
rect -9466 -75664 -9456 -75364
rect -10076 -75669 -9456 -75664
rect -7588 -75364 -6968 -75359
rect -7588 -75664 -7578 -75364
rect -6978 -75664 -6968 -75364
rect -7588 -75669 -6968 -75664
rect -6076 -75364 -5456 -75359
rect -6076 -75664 -6066 -75364
rect -5466 -75664 -5456 -75364
rect -6076 -75669 -5456 -75664
rect -3588 -75364 -2968 -75359
rect -3588 -75664 -3578 -75364
rect -2978 -75664 -2968 -75364
rect -3588 -75669 -2968 -75664
rect -2076 -75364 -1456 -75359
rect -2076 -75664 -2066 -75364
rect -1466 -75664 -1456 -75364
rect -2076 -75669 -1456 -75664
rect 412 -75364 1032 -75359
rect 412 -75664 422 -75364
rect 1022 -75664 1032 -75364
rect 412 -75669 1032 -75664
rect 1924 -75364 2544 -75359
rect 1924 -75664 1934 -75364
rect 2534 -75664 2544 -75364
rect 1924 -75669 2544 -75664
rect 4412 -75364 5032 -75359
rect 4412 -75664 4422 -75364
rect 5022 -75664 5032 -75364
rect 4412 -75669 5032 -75664
rect 5924 -75364 6544 -75359
rect 5924 -75664 5934 -75364
rect 6534 -75664 6544 -75364
rect 5924 -75669 6544 -75664
<< via3 >>
rect -27620 -28652 -27556 -27370
rect -25514 -28652 -25450 -27370
rect -23408 -28652 -23344 -27370
rect -21302 -28652 -21238 -27370
rect -19196 -28652 -19132 -27370
rect -17090 -28652 -17026 -27370
rect -14984 -28652 -14920 -27370
rect -12878 -28652 -12814 -27370
rect -10772 -28652 -10708 -27370
rect -8666 -28652 -8602 -27370
rect -6560 -28652 -6496 -27370
rect -4454 -28652 -4390 -27370
rect -2348 -28652 -2284 -27370
rect -242 -28652 -178 -27370
rect 1864 -28652 1928 -27370
rect 3970 -28652 4034 -27370
rect 6076 -28652 6140 -27370
rect 8182 -28652 8246 -27370
rect 25928 -28062 26528 -27762
rect 49560 -28062 50160 -27762
rect 29505 -28358 46290 -28144
rect -27620 -30652 -27556 -29370
rect -25514 -30652 -25450 -29370
rect -23408 -30652 -23344 -29370
rect -21302 -30652 -21238 -29370
rect -19196 -30652 -19132 -29370
rect -17090 -30652 -17026 -29370
rect -14984 -30652 -14920 -29370
rect -12878 -30652 -12814 -29370
rect -10772 -30652 -10708 -29370
rect -8666 -30652 -8602 -29370
rect -6560 -30652 -6496 -29370
rect -4454 -30652 -4390 -29370
rect -2348 -30652 -2284 -29370
rect -242 -30652 -178 -29370
rect 1864 -30652 1928 -29370
rect 3970 -30652 4034 -29370
rect 6076 -30652 6140 -29370
rect 8182 -30652 8246 -29370
rect 10428 -29738 11124 -29048
rect 24470 -29736 25160 -29038
rect -27620 -32652 -27556 -31370
rect -25514 -32652 -25450 -31370
rect -23408 -32652 -23344 -31370
rect -21302 -32652 -21238 -31370
rect -19196 -32652 -19132 -31370
rect -17090 -32652 -17026 -31370
rect -14984 -32652 -14920 -31370
rect -12878 -32652 -12814 -31370
rect -10772 -32652 -10708 -31370
rect -8666 -32652 -8602 -31370
rect -6560 -32652 -6496 -31370
rect -4454 -32652 -4390 -31370
rect -2348 -32652 -2284 -31370
rect -242 -32652 -178 -31370
rect 1864 -32652 1928 -31370
rect 3970 -32652 4034 -31370
rect 6076 -32652 6140 -31370
rect 8182 -32652 8246 -31370
rect -27620 -34652 -27556 -33370
rect -25514 -34652 -25450 -33370
rect -23408 -34652 -23344 -33370
rect -21302 -34652 -21238 -33370
rect -19196 -34652 -19132 -33370
rect -17090 -34652 -17026 -33370
rect -14984 -34652 -14920 -33370
rect -12878 -34652 -12814 -33370
rect -10772 -34652 -10708 -33370
rect -8666 -34652 -8602 -33370
rect -6560 -34652 -6496 -33370
rect -4454 -34652 -4390 -33370
rect -2348 -34652 -2284 -33370
rect -242 -34652 -178 -33370
rect 1864 -34652 1928 -33370
rect 3970 -34652 4034 -33370
rect 6076 -34652 6140 -33370
rect 8182 -34652 8246 -33370
rect -27620 -36652 -27556 -35370
rect -25514 -36652 -25450 -35370
rect -23408 -36652 -23344 -35370
rect -21302 -36652 -21238 -35370
rect -19196 -36652 -19132 -35370
rect -17090 -36652 -17026 -35370
rect -14984 -36652 -14920 -35370
rect -12878 -36652 -12814 -35370
rect -10772 -36652 -10708 -35370
rect -8666 -36652 -8602 -35370
rect -6560 -36652 -6496 -35370
rect -4454 -36652 -4390 -35370
rect -2348 -36652 -2284 -35370
rect -242 -36652 -178 -35370
rect 1864 -36652 1928 -35370
rect 3970 -36652 4034 -35370
rect 6076 -36652 6140 -35370
rect 8182 -36652 8246 -35370
rect -27620 -38652 -27556 -37370
rect -25514 -38652 -25450 -37370
rect -23408 -38652 -23344 -37370
rect -21302 -38652 -21238 -37370
rect -19196 -38652 -19132 -37370
rect -17090 -38652 -17026 -37370
rect -14984 -38652 -14920 -37370
rect -12878 -38652 -12814 -37370
rect -10772 -38652 -10708 -37370
rect -8666 -38652 -8602 -37370
rect -6560 -38652 -6496 -37370
rect -4454 -38652 -4390 -37370
rect -2348 -38652 -2284 -37370
rect -242 -38652 -178 -37370
rect 1864 -38652 1928 -37370
rect 3970 -38652 4034 -37370
rect 6076 -38652 6140 -37370
rect 8182 -38652 8246 -37370
rect -27620 -40652 -27556 -39370
rect -25514 -40652 -25450 -39370
rect -23408 -40652 -23344 -39370
rect -21302 -40652 -21238 -39370
rect -19196 -40652 -19132 -39370
rect -17090 -40652 -17026 -39370
rect -14984 -40652 -14920 -39370
rect -12878 -40652 -12814 -39370
rect -10772 -40652 -10708 -39370
rect -8666 -40652 -8602 -39370
rect -6560 -40652 -6496 -39370
rect -4454 -40652 -4390 -39370
rect -2348 -40652 -2284 -39370
rect -242 -40652 -178 -39370
rect 1864 -40652 1928 -39370
rect 3970 -40652 4034 -39370
rect 6076 -40652 6140 -39370
rect 8182 -40652 8246 -39370
rect -27620 -42652 -27556 -41370
rect -25514 -42652 -25450 -41370
rect -23408 -42652 -23344 -41370
rect -21302 -42652 -21238 -41370
rect -19196 -42652 -19132 -41370
rect -17090 -42652 -17026 -41370
rect -14984 -42652 -14920 -41370
rect -12878 -42652 -12814 -41370
rect -10772 -42652 -10708 -41370
rect -8666 -42652 -8602 -41370
rect -6560 -42652 -6496 -41370
rect -4454 -42652 -4390 -41370
rect -2348 -42652 -2284 -41370
rect -242 -42652 -178 -41370
rect 1864 -42652 1928 -41370
rect 3970 -42652 4034 -41370
rect 6076 -42652 6140 -41370
rect 8182 -42652 8246 -41370
rect 52262 -39386 55130 -39086
rect 56534 -39386 58154 -39086
rect 57475 -40476 57539 -40471
rect 57475 -40536 57534 -40476
rect 57534 -40536 57539 -40476
rect 57475 -40541 57539 -40536
rect -27620 -44652 -27556 -43370
rect -25514 -44652 -25450 -43370
rect -23408 -44652 -23344 -43370
rect -21302 -44652 -21238 -43370
rect -19196 -44652 -19132 -43370
rect -17090 -44652 -17026 -43370
rect -14984 -44652 -14920 -43370
rect -12878 -44652 -12814 -43370
rect -10772 -44652 -10708 -43370
rect -8666 -44652 -8602 -43370
rect -6560 -44652 -6496 -43370
rect -4454 -44652 -4390 -43370
rect -2348 -44652 -2284 -43370
rect -242 -44652 -178 -43370
rect 1864 -44652 1928 -43370
rect 3970 -44652 4034 -43370
rect 6076 -44652 6140 -43370
rect 8182 -44652 8246 -43370
rect 26981 -42942 27051 -42937
rect 26981 -43001 26986 -42942
rect 26986 -43001 27046 -42942
rect 27046 -43001 27051 -42942
rect 27759 -42927 27857 -42923
rect 27759 -43017 27763 -42927
rect 27763 -43017 27853 -42927
rect 27853 -43017 27857 -42927
rect 27759 -43021 27857 -43017
rect -27620 -46652 -27556 -45370
rect -25514 -46652 -25450 -45370
rect -23408 -46652 -23344 -45370
rect -21302 -46652 -21238 -45370
rect -19196 -46652 -19132 -45370
rect -17090 -46652 -17026 -45370
rect -14984 -46652 -14920 -45370
rect -12878 -46652 -12814 -45370
rect -10772 -46652 -10708 -45370
rect -8666 -46652 -8602 -45370
rect -6560 -46652 -6496 -45370
rect -4454 -46652 -4390 -45370
rect -2348 -46652 -2284 -45370
rect -242 -46652 -178 -45370
rect 1864 -46652 1928 -45370
rect 3970 -46652 4034 -45370
rect 6076 -46652 6140 -45370
rect 8182 -46652 8246 -45370
rect -27620 -48652 -27556 -47370
rect -25514 -48652 -25450 -47370
rect -23408 -48652 -23344 -47370
rect -21302 -48652 -21238 -47370
rect -19196 -48652 -19132 -47370
rect -17090 -48652 -17026 -47370
rect -14984 -48652 -14920 -47370
rect -12878 -48652 -12814 -47370
rect -10772 -48652 -10708 -47370
rect -8666 -48652 -8602 -47370
rect -6560 -48652 -6496 -47370
rect -4454 -48652 -4390 -47370
rect -2348 -48652 -2284 -47370
rect -242 -48652 -178 -47370
rect 1864 -48652 1928 -47370
rect 3970 -48652 4034 -47370
rect 6076 -48652 6140 -47370
rect 8182 -48652 8246 -47370
rect -27620 -50652 -27556 -49370
rect -25514 -50652 -25450 -49370
rect -23408 -50652 -23344 -49370
rect -21302 -50652 -21238 -49370
rect -19196 -50652 -19132 -49370
rect -17090 -50652 -17026 -49370
rect -14984 -50652 -14920 -49370
rect -12878 -50652 -12814 -49370
rect -10772 -50652 -10708 -49370
rect -8666 -50652 -8602 -49370
rect -6560 -50652 -6496 -49370
rect -4454 -50652 -4390 -49370
rect -2348 -50652 -2284 -49370
rect -242 -50652 -178 -49370
rect 1864 -50652 1928 -49370
rect 3970 -50652 4034 -49370
rect 6076 -50652 6140 -49370
rect 8182 -50652 8246 -49370
rect -27620 -52652 -27556 -51370
rect -25514 -52652 -25450 -51370
rect -23408 -52652 -23344 -51370
rect -21302 -52652 -21238 -51370
rect -19196 -52652 -19132 -51370
rect -17090 -52652 -17026 -51370
rect -14984 -52652 -14920 -51370
rect -12878 -52652 -12814 -51370
rect -10772 -52652 -10708 -51370
rect -8666 -52652 -8602 -51370
rect -6560 -52652 -6496 -51370
rect -4454 -52652 -4390 -51370
rect -2348 -52652 -2284 -51370
rect -242 -52652 -178 -51370
rect 1864 -52652 1928 -51370
rect 3970 -52652 4034 -51370
rect 6076 -52652 6140 -51370
rect 8182 -52652 8246 -51370
rect 8165 -53047 8263 -52949
rect -27620 -54652 -27556 -53370
rect -25514 -54652 -25450 -53370
rect -23408 -54652 -23344 -53370
rect -21302 -54652 -21238 -53370
rect -19196 -54652 -19132 -53370
rect -17090 -54652 -17026 -53370
rect -14984 -54652 -14920 -53370
rect -12878 -54652 -12814 -53370
rect -10772 -54652 -10708 -53370
rect -8666 -54652 -8602 -53370
rect -6560 -54652 -6496 -53370
rect -4454 -54652 -4390 -53370
rect -2348 -54652 -2284 -53370
rect -242 -54652 -178 -53370
rect 1864 -54652 1928 -53370
rect 3970 -54652 4034 -53370
rect 6076 -54652 6140 -53370
rect 8182 -54652 8246 -53370
rect 8163 -55047 8261 -54949
rect -27620 -56652 -27556 -55370
rect -25514 -56652 -25450 -55370
rect -23408 -56652 -23344 -55370
rect -21302 -56652 -21238 -55370
rect -19196 -56652 -19132 -55370
rect -17090 -56652 -17026 -55370
rect -14984 -56652 -14920 -55370
rect -12878 -56652 -12814 -55370
rect -10772 -56652 -10708 -55370
rect -8666 -56652 -8602 -55370
rect -6560 -56652 -6496 -55370
rect -4454 -56652 -4390 -55370
rect -2348 -56652 -2284 -55370
rect -242 -56652 -178 -55370
rect 1864 -56652 1928 -55370
rect 3970 -56652 4034 -55370
rect 6076 -56652 6140 -55370
rect 8182 -56652 8246 -55370
rect -27620 -58652 -27556 -57370
rect -25514 -58652 -25450 -57370
rect -23408 -58652 -23344 -57370
rect -21302 -58652 -21238 -57370
rect -19196 -58652 -19132 -57370
rect -17090 -58652 -17026 -57370
rect -14984 -58652 -14920 -57370
rect -12878 -58652 -12814 -57370
rect -10772 -58652 -10708 -57370
rect -8666 -58652 -8602 -57370
rect -6560 -58652 -6496 -57370
rect -4454 -58652 -4390 -57370
rect -2348 -58652 -2284 -57370
rect -242 -58652 -178 -57370
rect 1864 -58652 1928 -57370
rect 3970 -58652 4034 -57370
rect 6076 -58652 6140 -57370
rect 8182 -58652 8246 -57370
rect 9372 -57518 9436 -56724
rect 10294 -58514 12110 -58408
rect -27620 -60652 -27556 -59370
rect -25514 -60652 -25450 -59370
rect -23408 -60652 -23344 -59370
rect -21302 -60652 -21238 -59370
rect -19196 -60652 -19132 -59370
rect -17090 -60652 -17026 -59370
rect -14984 -60652 -14920 -59370
rect -12878 -60652 -12814 -59370
rect -10772 -60652 -10708 -59370
rect -8666 -60652 -8602 -59370
rect -6560 -60652 -6496 -59370
rect -4454 -60652 -4390 -59370
rect -2348 -60652 -2284 -59370
rect -242 -60652 -178 -59370
rect 1864 -60652 1928 -59370
rect 3970 -60652 4034 -59370
rect 6076 -60652 6140 -59370
rect 8182 -60652 8246 -59370
rect -27620 -62652 -27556 -61370
rect -25514 -62652 -25450 -61370
rect -23408 -62652 -23344 -61370
rect -21302 -62652 -21238 -61370
rect -19196 -62652 -19132 -61370
rect -17090 -62652 -17026 -61370
rect -14984 -62652 -14920 -61370
rect -12878 -62652 -12814 -61370
rect -10772 -62652 -10708 -61370
rect -8666 -62652 -8602 -61370
rect -6560 -62652 -6496 -61370
rect -4454 -62652 -4390 -61370
rect -2348 -62652 -2284 -61370
rect -242 -62652 -178 -61370
rect 1864 -62652 1928 -61370
rect 3970 -62652 4034 -61370
rect 6076 -62652 6140 -61370
rect 8182 -62652 8246 -61370
rect -18963 -63113 -18865 -63015
rect -16847 -63109 -16749 -63011
rect -14751 -63107 -14653 -63009
rect -25200 -63378 -25100 -63278
rect -27578 -64832 -26978 -64532
rect -26066 -64832 -25466 -64532
rect -27388 -65100 -25564 -65036
rect -23578 -64832 -22978 -64532
rect -22066 -64832 -21466 -64532
rect -23388 -65100 -21564 -65036
rect -19578 -64832 -18978 -64532
rect -18066 -64832 -17466 -64532
rect -19388 -65100 -17564 -65036
rect -12627 -63117 -12529 -63019
rect -10591 -63109 -10493 -63011
rect -9937 -63099 -9839 -63001
rect -8495 -63117 -8397 -63019
rect -7927 -63121 -7829 -63023
rect -15578 -64832 -14978 -64532
rect -14066 -64832 -13466 -64532
rect -11578 -64832 -10978 -64532
rect -10066 -64832 -9466 -64532
rect -15388 -65100 -13564 -65036
rect -11388 -65100 -9564 -65036
rect -7578 -64832 -6978 -64532
rect -6066 -64832 -5466 -64532
rect -7388 -65100 -5564 -65036
rect -3578 -64832 -2978 -64532
rect -2066 -64832 -1466 -64532
rect -3388 -65100 -1564 -65036
rect 422 -64832 1022 -64532
rect 1934 -64832 2534 -64532
rect 612 -65100 2436 -65036
rect 4422 -64832 5022 -64532
rect 5934 -64832 6534 -64532
rect 4612 -65100 6436 -65036
rect 17372 -58608 49372 -58454
rect 13228 -59094 13828 -58794
rect 49660 -59094 50260 -58794
rect 58424 -42308 58524 -42208
rect 53296 -42482 53396 -42460
rect 53296 -42542 53314 -42482
rect 53314 -42542 53374 -42482
rect 53374 -42542 53396 -42482
rect 53296 -42560 53396 -42542
rect 54195 -42476 54259 -42471
rect 54195 -42548 54200 -42476
rect 54200 -42548 54259 -42476
rect 54195 -42553 54259 -42548
rect 55300 -42471 55370 -42466
rect 55300 -42553 55365 -42471
rect 55365 -42553 55370 -42471
rect 55300 -42558 55370 -42553
rect 56043 -42577 56141 -42573
rect 56043 -42667 56047 -42577
rect 56047 -42667 56137 -42577
rect 56137 -42667 56141 -42577
rect 56043 -42671 56141 -42667
rect 57947 -42579 58045 -42575
rect 57947 -42669 57951 -42579
rect 57951 -42669 58041 -42579
rect 58041 -42669 58045 -42579
rect 57947 -42673 58045 -42669
rect 55824 -43584 58268 -43278
rect -27430 -69222 -25722 -69154
rect -27578 -69704 -26978 -69404
rect -26066 -69704 -25466 -69404
rect -27578 -70792 -26978 -70492
rect -26066 -70792 -25466 -70492
rect -27430 -71042 -25722 -70974
rect -23430 -69222 -21722 -69154
rect -23578 -69704 -22978 -69404
rect -22066 -69704 -21466 -69404
rect -23578 -70792 -22978 -70492
rect -22066 -70792 -21466 -70492
rect -23430 -71042 -21722 -70974
rect -19430 -69222 -17722 -69154
rect -19578 -69704 -18978 -69404
rect -18066 -69704 -17466 -69404
rect -19578 -70792 -18978 -70492
rect -18066 -70792 -17466 -70492
rect -19430 -71042 -17722 -70974
rect -15430 -69222 -13722 -69154
rect -15578 -69704 -14978 -69404
rect -14066 -69704 -13466 -69404
rect -15578 -70792 -14978 -70492
rect -14066 -70792 -13466 -70492
rect -15430 -71042 -13722 -70974
rect -11430 -69222 -9722 -69154
rect -11578 -69704 -10978 -69404
rect -10066 -69704 -9466 -69404
rect -11578 -70792 -10978 -70492
rect -10066 -70792 -9466 -70492
rect -11430 -71042 -9722 -70974
rect -7430 -69222 -5722 -69154
rect -7578 -69704 -6978 -69404
rect -6066 -69704 -5466 -69404
rect -7578 -70792 -6978 -70492
rect -6066 -70792 -5466 -70492
rect -7430 -71042 -5722 -70974
rect -3430 -69222 -1722 -69154
rect -3578 -69704 -2978 -69404
rect -2066 -69704 -1466 -69404
rect -3578 -70792 -2978 -70492
rect -2066 -70792 -1466 -70492
rect -3430 -71042 -1722 -70974
rect 570 -69222 2278 -69154
rect 422 -69704 1022 -69404
rect 1934 -69704 2534 -69404
rect 422 -70792 1022 -70492
rect 1934 -70792 2534 -70492
rect 570 -71042 2278 -70974
rect 4570 -69222 6278 -69154
rect 4422 -69704 5022 -69404
rect 5934 -69704 6534 -69404
rect 4422 -70792 5022 -70492
rect 5934 -70792 6534 -70492
rect 4570 -71042 6278 -70974
rect -27388 -75160 -25564 -75096
rect -23388 -75160 -21564 -75096
rect -19388 -75160 -17564 -75096
rect -15388 -75160 -13564 -75096
rect -11388 -75160 -9564 -75096
rect -7388 -75160 -5564 -75096
rect -3388 -75160 -1564 -75096
rect 612 -75160 2436 -75096
rect 4612 -75160 6436 -75096
rect -27578 -75664 -26978 -75364
rect -26066 -75664 -25466 -75364
rect -23578 -75664 -22978 -75364
rect -22066 -75664 -21466 -75364
rect -19578 -75664 -18978 -75364
rect -18066 -75664 -17466 -75364
rect -15578 -75664 -14978 -75364
rect -14066 -75664 -13466 -75364
rect -11578 -75664 -10978 -75364
rect -10066 -75664 -9466 -75364
rect -7578 -75664 -6978 -75364
rect -6066 -75664 -5466 -75364
rect -3578 -75664 -2978 -75364
rect -2066 -75664 -1466 -75364
rect 422 -75664 1022 -75364
rect 1934 -75664 2534 -75364
rect 4422 -75664 5022 -75364
rect 5934 -75664 6534 -75364
<< mimcap >>
rect -29135 -27346 -27735 -27306
rect -29135 -28666 -29095 -27346
rect -27775 -28666 -27735 -27346
rect -29135 -28706 -27735 -28666
rect -27029 -27346 -25629 -27306
rect -27029 -28666 -26989 -27346
rect -25669 -28666 -25629 -27346
rect -27029 -28706 -25629 -28666
rect -24923 -27346 -23523 -27306
rect -24923 -28666 -24883 -27346
rect -23563 -28666 -23523 -27346
rect -24923 -28706 -23523 -28666
rect -22817 -27346 -21417 -27306
rect -22817 -28666 -22777 -27346
rect -21457 -28666 -21417 -27346
rect -22817 -28706 -21417 -28666
rect -20711 -27346 -19311 -27306
rect -20711 -28666 -20671 -27346
rect -19351 -28666 -19311 -27346
rect -20711 -28706 -19311 -28666
rect -18605 -27346 -17205 -27306
rect -18605 -28666 -18565 -27346
rect -17245 -28666 -17205 -27346
rect -18605 -28706 -17205 -28666
rect -16499 -27346 -15099 -27306
rect -16499 -28666 -16459 -27346
rect -15139 -28666 -15099 -27346
rect -16499 -28706 -15099 -28666
rect -14393 -27346 -12993 -27306
rect -14393 -28666 -14353 -27346
rect -13033 -28666 -12993 -27346
rect -14393 -28706 -12993 -28666
rect -12287 -27346 -10887 -27306
rect -12287 -28666 -12247 -27346
rect -10927 -28666 -10887 -27346
rect -12287 -28706 -10887 -28666
rect -10181 -27346 -8781 -27306
rect -10181 -28666 -10141 -27346
rect -8821 -28666 -8781 -27346
rect -10181 -28706 -8781 -28666
rect -8075 -27346 -6675 -27306
rect -8075 -28666 -8035 -27346
rect -6715 -28666 -6675 -27346
rect -8075 -28706 -6675 -28666
rect -5969 -27346 -4569 -27306
rect -5969 -28666 -5929 -27346
rect -4609 -28666 -4569 -27346
rect -5969 -28706 -4569 -28666
rect -3863 -27346 -2463 -27306
rect -3863 -28666 -3823 -27346
rect -2503 -28666 -2463 -27346
rect -3863 -28706 -2463 -28666
rect -1757 -27346 -357 -27306
rect -1757 -28666 -1717 -27346
rect -397 -28666 -357 -27346
rect -1757 -28706 -357 -28666
rect 349 -27346 1749 -27306
rect 349 -28666 389 -27346
rect 1709 -28666 1749 -27346
rect 349 -28706 1749 -28666
rect 2455 -27346 3855 -27306
rect 2455 -28666 2495 -27346
rect 3815 -28666 3855 -27346
rect 2455 -28706 3855 -28666
rect 4561 -27346 5961 -27306
rect 4561 -28666 4601 -27346
rect 5921 -28666 5961 -27346
rect 4561 -28706 5961 -28666
rect 6667 -27346 8067 -27306
rect 6667 -28666 6707 -27346
rect 8027 -28666 8067 -27346
rect 6667 -28706 8067 -28666
rect 11462 -29042 17662 -28992
rect -29135 -29346 -27735 -29306
rect -29135 -30666 -29095 -29346
rect -27775 -30666 -27735 -29346
rect -29135 -30706 -27735 -30666
rect -27029 -29346 -25629 -29306
rect -27029 -30666 -26989 -29346
rect -25669 -30666 -25629 -29346
rect -27029 -30706 -25629 -30666
rect -24923 -29346 -23523 -29306
rect -24923 -30666 -24883 -29346
rect -23563 -30666 -23523 -29346
rect -24923 -30706 -23523 -30666
rect -22817 -29346 -21417 -29306
rect -22817 -30666 -22777 -29346
rect -21457 -30666 -21417 -29346
rect -22817 -30706 -21417 -30666
rect -20711 -29346 -19311 -29306
rect -20711 -30666 -20671 -29346
rect -19351 -30666 -19311 -29346
rect -20711 -30706 -19311 -30666
rect -18605 -29346 -17205 -29306
rect -18605 -30666 -18565 -29346
rect -17245 -30666 -17205 -29346
rect -18605 -30706 -17205 -30666
rect -16499 -29346 -15099 -29306
rect -16499 -30666 -16459 -29346
rect -15139 -30666 -15099 -29346
rect -16499 -30706 -15099 -30666
rect -14393 -29346 -12993 -29306
rect -14393 -30666 -14353 -29346
rect -13033 -30666 -12993 -29346
rect -14393 -30706 -12993 -30666
rect -12287 -29346 -10887 -29306
rect -12287 -30666 -12247 -29346
rect -10927 -30666 -10887 -29346
rect -12287 -30706 -10887 -30666
rect -10181 -29346 -8781 -29306
rect -10181 -30666 -10141 -29346
rect -8821 -30666 -8781 -29346
rect -10181 -30706 -8781 -30666
rect -8075 -29346 -6675 -29306
rect -8075 -30666 -8035 -29346
rect -6715 -30666 -6675 -29346
rect -8075 -30706 -6675 -30666
rect -5969 -29346 -4569 -29306
rect -5969 -30666 -5929 -29346
rect -4609 -30666 -4569 -29346
rect -5969 -30706 -4569 -30666
rect -3863 -29346 -2463 -29306
rect -3863 -30666 -3823 -29346
rect -2503 -30666 -2463 -29346
rect -3863 -30706 -2463 -30666
rect -1757 -29346 -357 -29306
rect -1757 -30666 -1717 -29346
rect -397 -30666 -357 -29346
rect -1757 -30706 -357 -30666
rect 349 -29346 1749 -29306
rect 349 -30666 389 -29346
rect 1709 -30666 1749 -29346
rect 349 -30706 1749 -30666
rect 2455 -29346 3855 -29306
rect 2455 -30666 2495 -29346
rect 3815 -30666 3855 -29346
rect 2455 -30706 3855 -30666
rect 4561 -29346 5961 -29306
rect 4561 -30666 4601 -29346
rect 5921 -30666 5961 -29346
rect 4561 -30706 5961 -30666
rect 6667 -29346 8067 -29306
rect 6667 -30666 6707 -29346
rect 8027 -30666 8067 -29346
rect 11462 -29342 17312 -29042
rect 17612 -29342 17662 -29042
rect 11462 -29392 17662 -29342
rect 17862 -29042 24062 -28992
rect 17862 -29342 23712 -29042
rect 24012 -29342 24062 -29042
rect 17862 -29392 24062 -29342
rect 6667 -30706 8067 -30666
rect 10376 -30124 11176 -30074
rect -29135 -31346 -27735 -31306
rect -29135 -32666 -29095 -31346
rect -27775 -32666 -27735 -31346
rect -29135 -32706 -27735 -32666
rect -27029 -31346 -25629 -31306
rect -27029 -32666 -26989 -31346
rect -25669 -32666 -25629 -31346
rect -27029 -32706 -25629 -32666
rect -24923 -31346 -23523 -31306
rect -24923 -32666 -24883 -31346
rect -23563 -32666 -23523 -31346
rect -24923 -32706 -23523 -32666
rect -22817 -31346 -21417 -31306
rect -22817 -32666 -22777 -31346
rect -21457 -32666 -21417 -31346
rect -22817 -32706 -21417 -32666
rect -20711 -31346 -19311 -31306
rect -20711 -32666 -20671 -31346
rect -19351 -32666 -19311 -31346
rect -20711 -32706 -19311 -32666
rect -18605 -31346 -17205 -31306
rect -18605 -32666 -18565 -31346
rect -17245 -32666 -17205 -31346
rect -18605 -32706 -17205 -32666
rect -16499 -31346 -15099 -31306
rect -16499 -32666 -16459 -31346
rect -15139 -32666 -15099 -31346
rect -16499 -32706 -15099 -32666
rect -14393 -31346 -12993 -31306
rect -14393 -32666 -14353 -31346
rect -13033 -32666 -12993 -31346
rect -14393 -32706 -12993 -32666
rect -12287 -31346 -10887 -31306
rect -12287 -32666 -12247 -31346
rect -10927 -32666 -10887 -31346
rect -12287 -32706 -10887 -32666
rect -10181 -31346 -8781 -31306
rect -10181 -32666 -10141 -31346
rect -8821 -32666 -8781 -31346
rect -10181 -32706 -8781 -32666
rect -8075 -31346 -6675 -31306
rect -8075 -32666 -8035 -31346
rect -6715 -32666 -6675 -31346
rect -8075 -32706 -6675 -32666
rect -5969 -31346 -4569 -31306
rect -5969 -32666 -5929 -31346
rect -4609 -32666 -4569 -31346
rect -5969 -32706 -4569 -32666
rect -3863 -31346 -2463 -31306
rect -3863 -32666 -3823 -31346
rect -2503 -32666 -2463 -31346
rect -3863 -32706 -2463 -32666
rect -1757 -31346 -357 -31306
rect -1757 -32666 -1717 -31346
rect -397 -32666 -357 -31346
rect -1757 -32706 -357 -32666
rect 349 -31346 1749 -31306
rect 349 -32666 389 -31346
rect 1709 -32666 1749 -31346
rect 349 -32706 1749 -32666
rect 2455 -31346 3855 -31306
rect 2455 -32666 2495 -31346
rect 3815 -32666 3855 -31346
rect 2455 -32706 3855 -32666
rect 4561 -31346 5961 -31306
rect 4561 -32666 4601 -31346
rect 5921 -32666 5961 -31346
rect 4561 -32706 5961 -32666
rect 6667 -31346 8067 -31306
rect 6667 -32666 6707 -31346
rect 8027 -32666 8067 -31346
rect 6667 -32706 8067 -32666
rect -29135 -33346 -27735 -33306
rect -29135 -34666 -29095 -33346
rect -27775 -34666 -27735 -33346
rect -29135 -34706 -27735 -34666
rect -27029 -33346 -25629 -33306
rect -27029 -34666 -26989 -33346
rect -25669 -34666 -25629 -33346
rect -27029 -34706 -25629 -34666
rect -24923 -33346 -23523 -33306
rect -24923 -34666 -24883 -33346
rect -23563 -34666 -23523 -33346
rect -24923 -34706 -23523 -34666
rect -22817 -33346 -21417 -33306
rect -22817 -34666 -22777 -33346
rect -21457 -34666 -21417 -33346
rect -22817 -34706 -21417 -34666
rect -20711 -33346 -19311 -33306
rect -20711 -34666 -20671 -33346
rect -19351 -34666 -19311 -33346
rect -20711 -34706 -19311 -34666
rect -18605 -33346 -17205 -33306
rect -18605 -34666 -18565 -33346
rect -17245 -34666 -17205 -33346
rect -18605 -34706 -17205 -34666
rect -16499 -33346 -15099 -33306
rect -16499 -34666 -16459 -33346
rect -15139 -34666 -15099 -33346
rect -16499 -34706 -15099 -34666
rect -14393 -33346 -12993 -33306
rect -14393 -34666 -14353 -33346
rect -13033 -34666 -12993 -33346
rect -14393 -34706 -12993 -34666
rect -12287 -33346 -10887 -33306
rect -12287 -34666 -12247 -33346
rect -10927 -34666 -10887 -33346
rect -12287 -34706 -10887 -34666
rect -10181 -33346 -8781 -33306
rect -10181 -34666 -10141 -33346
rect -8821 -34666 -8781 -33346
rect -10181 -34706 -8781 -34666
rect -8075 -33346 -6675 -33306
rect -8075 -34666 -8035 -33346
rect -6715 -34666 -6675 -33346
rect -8075 -34706 -6675 -34666
rect -5969 -33346 -4569 -33306
rect -5969 -34666 -5929 -33346
rect -4609 -34666 -4569 -33346
rect -5969 -34706 -4569 -34666
rect -3863 -33346 -2463 -33306
rect -3863 -34666 -3823 -33346
rect -2503 -34666 -2463 -33346
rect -3863 -34706 -2463 -34666
rect -1757 -33346 -357 -33306
rect -1757 -34666 -1717 -33346
rect -397 -34666 -357 -33346
rect -1757 -34706 -357 -34666
rect 349 -33346 1749 -33306
rect 349 -34666 389 -33346
rect 1709 -34666 1749 -33346
rect 349 -34706 1749 -34666
rect 2455 -33346 3855 -33306
rect 2455 -34666 2495 -33346
rect 3815 -34666 3855 -33346
rect 2455 -34706 3855 -34666
rect 4561 -33346 5961 -33306
rect 4561 -34666 4601 -33346
rect 5921 -34666 5961 -33346
rect 4561 -34706 5961 -34666
rect 6667 -33346 8067 -33306
rect 6667 -34666 6707 -33346
rect 8027 -34666 8067 -33346
rect 6667 -34706 8067 -34666
rect -29135 -35346 -27735 -35306
rect -29135 -36666 -29095 -35346
rect -27775 -36666 -27735 -35346
rect -29135 -36706 -27735 -36666
rect -27029 -35346 -25629 -35306
rect -27029 -36666 -26989 -35346
rect -25669 -36666 -25629 -35346
rect -27029 -36706 -25629 -36666
rect -24923 -35346 -23523 -35306
rect -24923 -36666 -24883 -35346
rect -23563 -36666 -23523 -35346
rect -24923 -36706 -23523 -36666
rect -22817 -35346 -21417 -35306
rect -22817 -36666 -22777 -35346
rect -21457 -36666 -21417 -35346
rect -22817 -36706 -21417 -36666
rect -20711 -35346 -19311 -35306
rect -20711 -36666 -20671 -35346
rect -19351 -36666 -19311 -35346
rect -20711 -36706 -19311 -36666
rect -18605 -35346 -17205 -35306
rect -18605 -36666 -18565 -35346
rect -17245 -36666 -17205 -35346
rect -18605 -36706 -17205 -36666
rect -16499 -35346 -15099 -35306
rect -16499 -36666 -16459 -35346
rect -15139 -36666 -15099 -35346
rect -16499 -36706 -15099 -36666
rect -14393 -35346 -12993 -35306
rect -14393 -36666 -14353 -35346
rect -13033 -36666 -12993 -35346
rect -14393 -36706 -12993 -36666
rect -12287 -35346 -10887 -35306
rect -12287 -36666 -12247 -35346
rect -10927 -36666 -10887 -35346
rect -12287 -36706 -10887 -36666
rect -10181 -35346 -8781 -35306
rect -10181 -36666 -10141 -35346
rect -8821 -36666 -8781 -35346
rect -10181 -36706 -8781 -36666
rect -8075 -35346 -6675 -35306
rect -8075 -36666 -8035 -35346
rect -6715 -36666 -6675 -35346
rect -8075 -36706 -6675 -36666
rect -5969 -35346 -4569 -35306
rect -5969 -36666 -5929 -35346
rect -4609 -36666 -4569 -35346
rect -5969 -36706 -4569 -36666
rect -3863 -35346 -2463 -35306
rect -3863 -36666 -3823 -35346
rect -2503 -36666 -2463 -35346
rect -3863 -36706 -2463 -36666
rect -1757 -35346 -357 -35306
rect -1757 -36666 -1717 -35346
rect -397 -36666 -357 -35346
rect -1757 -36706 -357 -36666
rect 349 -35346 1749 -35306
rect 349 -36666 389 -35346
rect 1709 -36666 1749 -35346
rect 349 -36706 1749 -36666
rect 2455 -35346 3855 -35306
rect 2455 -36666 2495 -35346
rect 3815 -36666 3855 -35346
rect 2455 -36706 3855 -36666
rect 4561 -35346 5961 -35306
rect 4561 -36666 4601 -35346
rect 5921 -36666 5961 -35346
rect 4561 -36706 5961 -36666
rect 6667 -35346 8067 -35306
rect 6667 -36666 6707 -35346
rect 8027 -36666 8067 -35346
rect 10376 -35824 10826 -30124
rect 11126 -35824 11176 -30124
rect 24420 -30124 25220 -30074
rect 12316 -31042 17516 -30992
rect 12316 -35742 17166 -31042
rect 17466 -35742 17516 -31042
rect 12316 -35792 17516 -35742
rect 17916 -31042 23116 -30992
rect 17916 -35742 22766 -31042
rect 23066 -35742 23116 -31042
rect 17916 -35792 23116 -35742
rect 10376 -35874 11176 -35824
rect 24420 -35824 24870 -30124
rect 25170 -35824 25220 -30124
rect 24420 -35874 25220 -35824
rect 6667 -36706 8067 -36666
rect 10376 -36616 11176 -36566
rect -29135 -37346 -27735 -37306
rect -29135 -38666 -29095 -37346
rect -27775 -38666 -27735 -37346
rect -29135 -38706 -27735 -38666
rect -27029 -37346 -25629 -37306
rect -27029 -38666 -26989 -37346
rect -25669 -38666 -25629 -37346
rect -27029 -38706 -25629 -38666
rect -24923 -37346 -23523 -37306
rect -24923 -38666 -24883 -37346
rect -23563 -38666 -23523 -37346
rect -24923 -38706 -23523 -38666
rect -22817 -37346 -21417 -37306
rect -22817 -38666 -22777 -37346
rect -21457 -38666 -21417 -37346
rect -22817 -38706 -21417 -38666
rect -20711 -37346 -19311 -37306
rect -20711 -38666 -20671 -37346
rect -19351 -38666 -19311 -37346
rect -20711 -38706 -19311 -38666
rect -18605 -37346 -17205 -37306
rect -18605 -38666 -18565 -37346
rect -17245 -38666 -17205 -37346
rect -18605 -38706 -17205 -38666
rect -16499 -37346 -15099 -37306
rect -16499 -38666 -16459 -37346
rect -15139 -38666 -15099 -37346
rect -16499 -38706 -15099 -38666
rect -14393 -37346 -12993 -37306
rect -14393 -38666 -14353 -37346
rect -13033 -38666 -12993 -37346
rect -14393 -38706 -12993 -38666
rect -12287 -37346 -10887 -37306
rect -12287 -38666 -12247 -37346
rect -10927 -38666 -10887 -37346
rect -12287 -38706 -10887 -38666
rect -10181 -37346 -8781 -37306
rect -10181 -38666 -10141 -37346
rect -8821 -38666 -8781 -37346
rect -10181 -38706 -8781 -38666
rect -8075 -37346 -6675 -37306
rect -8075 -38666 -8035 -37346
rect -6715 -38666 -6675 -37346
rect -8075 -38706 -6675 -38666
rect -5969 -37346 -4569 -37306
rect -5969 -38666 -5929 -37346
rect -4609 -38666 -4569 -37346
rect -5969 -38706 -4569 -38666
rect -3863 -37346 -2463 -37306
rect -3863 -38666 -3823 -37346
rect -2503 -38666 -2463 -37346
rect -3863 -38706 -2463 -38666
rect -1757 -37346 -357 -37306
rect -1757 -38666 -1717 -37346
rect -397 -38666 -357 -37346
rect -1757 -38706 -357 -38666
rect 349 -37346 1749 -37306
rect 349 -38666 389 -37346
rect 1709 -38666 1749 -37346
rect 349 -38706 1749 -38666
rect 2455 -37346 3855 -37306
rect 2455 -38666 2495 -37346
rect 3815 -38666 3855 -37346
rect 2455 -38706 3855 -38666
rect 4561 -37346 5961 -37306
rect 4561 -38666 4601 -37346
rect 5921 -38666 5961 -37346
rect 4561 -38706 5961 -38666
rect 6667 -37346 8067 -37306
rect 6667 -38666 6707 -37346
rect 8027 -38666 8067 -37346
rect 6667 -38706 8067 -38666
rect -29135 -39346 -27735 -39306
rect -29135 -40666 -29095 -39346
rect -27775 -40666 -27735 -39346
rect -29135 -40706 -27735 -40666
rect -27029 -39346 -25629 -39306
rect -27029 -40666 -26989 -39346
rect -25669 -40666 -25629 -39346
rect -27029 -40706 -25629 -40666
rect -24923 -39346 -23523 -39306
rect -24923 -40666 -24883 -39346
rect -23563 -40666 -23523 -39346
rect -24923 -40706 -23523 -40666
rect -22817 -39346 -21417 -39306
rect -22817 -40666 -22777 -39346
rect -21457 -40666 -21417 -39346
rect -22817 -40706 -21417 -40666
rect -20711 -39346 -19311 -39306
rect -20711 -40666 -20671 -39346
rect -19351 -40666 -19311 -39346
rect -20711 -40706 -19311 -40666
rect -18605 -39346 -17205 -39306
rect -18605 -40666 -18565 -39346
rect -17245 -40666 -17205 -39346
rect -18605 -40706 -17205 -40666
rect -16499 -39346 -15099 -39306
rect -16499 -40666 -16459 -39346
rect -15139 -40666 -15099 -39346
rect -16499 -40706 -15099 -40666
rect -14393 -39346 -12993 -39306
rect -14393 -40666 -14353 -39346
rect -13033 -40666 -12993 -39346
rect -14393 -40706 -12993 -40666
rect -12287 -39346 -10887 -39306
rect -12287 -40666 -12247 -39346
rect -10927 -40666 -10887 -39346
rect -12287 -40706 -10887 -40666
rect -10181 -39346 -8781 -39306
rect -10181 -40666 -10141 -39346
rect -8821 -40666 -8781 -39346
rect -10181 -40706 -8781 -40666
rect -8075 -39346 -6675 -39306
rect -8075 -40666 -8035 -39346
rect -6715 -40666 -6675 -39346
rect -8075 -40706 -6675 -40666
rect -5969 -39346 -4569 -39306
rect -5969 -40666 -5929 -39346
rect -4609 -40666 -4569 -39346
rect -5969 -40706 -4569 -40666
rect -3863 -39346 -2463 -39306
rect -3863 -40666 -3823 -39346
rect -2503 -40666 -2463 -39346
rect -3863 -40706 -2463 -40666
rect -1757 -39346 -357 -39306
rect -1757 -40666 -1717 -39346
rect -397 -40666 -357 -39346
rect -1757 -40706 -357 -40666
rect 349 -39346 1749 -39306
rect 349 -40666 389 -39346
rect 1709 -40666 1749 -39346
rect 349 -40706 1749 -40666
rect 2455 -39346 3855 -39306
rect 2455 -40666 2495 -39346
rect 3815 -40666 3855 -39346
rect 2455 -40706 3855 -40666
rect 4561 -39346 5961 -39306
rect 4561 -40666 4601 -39346
rect 5921 -40666 5961 -39346
rect 4561 -40706 5961 -40666
rect 6667 -39346 8067 -39306
rect 6667 -40666 6707 -39346
rect 8027 -40666 8067 -39346
rect 6667 -40706 8067 -40666
rect -29135 -41346 -27735 -41306
rect -29135 -42666 -29095 -41346
rect -27775 -42666 -27735 -41346
rect -29135 -42706 -27735 -42666
rect -27029 -41346 -25629 -41306
rect -27029 -42666 -26989 -41346
rect -25669 -42666 -25629 -41346
rect -27029 -42706 -25629 -42666
rect -24923 -41346 -23523 -41306
rect -24923 -42666 -24883 -41346
rect -23563 -42666 -23523 -41346
rect -24923 -42706 -23523 -42666
rect -22817 -41346 -21417 -41306
rect -22817 -42666 -22777 -41346
rect -21457 -42666 -21417 -41346
rect -22817 -42706 -21417 -42666
rect -20711 -41346 -19311 -41306
rect -20711 -42666 -20671 -41346
rect -19351 -42666 -19311 -41346
rect -20711 -42706 -19311 -42666
rect -18605 -41346 -17205 -41306
rect -18605 -42666 -18565 -41346
rect -17245 -42666 -17205 -41346
rect -18605 -42706 -17205 -42666
rect -16499 -41346 -15099 -41306
rect -16499 -42666 -16459 -41346
rect -15139 -42666 -15099 -41346
rect -16499 -42706 -15099 -42666
rect -14393 -41346 -12993 -41306
rect -14393 -42666 -14353 -41346
rect -13033 -42666 -12993 -41346
rect -14393 -42706 -12993 -42666
rect -12287 -41346 -10887 -41306
rect -12287 -42666 -12247 -41346
rect -10927 -42666 -10887 -41346
rect -12287 -42706 -10887 -42666
rect -10181 -41346 -8781 -41306
rect -10181 -42666 -10141 -41346
rect -8821 -42666 -8781 -41346
rect -10181 -42706 -8781 -42666
rect -8075 -41346 -6675 -41306
rect -8075 -42666 -8035 -41346
rect -6715 -42666 -6675 -41346
rect -8075 -42706 -6675 -42666
rect -5969 -41346 -4569 -41306
rect -5969 -42666 -5929 -41346
rect -4609 -42666 -4569 -41346
rect -5969 -42706 -4569 -42666
rect -3863 -41346 -2463 -41306
rect -3863 -42666 -3823 -41346
rect -2503 -42666 -2463 -41346
rect -3863 -42706 -2463 -42666
rect -1757 -41346 -357 -41306
rect -1757 -42666 -1717 -41346
rect -397 -42666 -357 -41346
rect -1757 -42706 -357 -42666
rect 349 -41346 1749 -41306
rect 349 -42666 389 -41346
rect 1709 -42666 1749 -41346
rect 349 -42706 1749 -42666
rect 2455 -41346 3855 -41306
rect 2455 -42666 2495 -41346
rect 3815 -42666 3855 -41346
rect 2455 -42706 3855 -42666
rect 4561 -41346 5961 -41306
rect 4561 -42666 4601 -41346
rect 5921 -42666 5961 -41346
rect 4561 -42706 5961 -42666
rect 6667 -41346 8067 -41306
rect 6667 -42666 6707 -41346
rect 8027 -42666 8067 -41346
rect 10376 -42316 10826 -36616
rect 11126 -42316 11176 -36616
rect 12316 -36642 17516 -36592
rect 12316 -41342 17166 -36642
rect 17466 -41342 17516 -36642
rect 12316 -41392 17516 -41342
rect 17916 -36642 23116 -36592
rect 17916 -41342 22766 -36642
rect 23066 -41342 23116 -36642
rect 17916 -41392 23116 -41342
rect 24420 -36616 25220 -36566
rect 10376 -42366 11176 -42316
rect 24420 -42316 24870 -36616
rect 25170 -42316 25220 -36616
rect 24420 -42366 25220 -42316
rect 6667 -42706 8067 -42666
rect 10962 -43042 17162 -42992
rect -29135 -43346 -27735 -43306
rect -29135 -44666 -29095 -43346
rect -27775 -44666 -27735 -43346
rect -29135 -44706 -27735 -44666
rect -27029 -43346 -25629 -43306
rect -27029 -44666 -26989 -43346
rect -25669 -44666 -25629 -43346
rect -27029 -44706 -25629 -44666
rect -24923 -43346 -23523 -43306
rect -24923 -44666 -24883 -43346
rect -23563 -44666 -23523 -43346
rect -24923 -44706 -23523 -44666
rect -22817 -43346 -21417 -43306
rect -22817 -44666 -22777 -43346
rect -21457 -44666 -21417 -43346
rect -22817 -44706 -21417 -44666
rect -20711 -43346 -19311 -43306
rect -20711 -44666 -20671 -43346
rect -19351 -44666 -19311 -43346
rect -20711 -44706 -19311 -44666
rect -18605 -43346 -17205 -43306
rect -18605 -44666 -18565 -43346
rect -17245 -44666 -17205 -43346
rect -18605 -44706 -17205 -44666
rect -16499 -43346 -15099 -43306
rect -16499 -44666 -16459 -43346
rect -15139 -44666 -15099 -43346
rect -16499 -44706 -15099 -44666
rect -14393 -43346 -12993 -43306
rect -14393 -44666 -14353 -43346
rect -13033 -44666 -12993 -43346
rect -14393 -44706 -12993 -44666
rect -12287 -43346 -10887 -43306
rect -12287 -44666 -12247 -43346
rect -10927 -44666 -10887 -43346
rect -12287 -44706 -10887 -44666
rect -10181 -43346 -8781 -43306
rect -10181 -44666 -10141 -43346
rect -8821 -44666 -8781 -43346
rect -10181 -44706 -8781 -44666
rect -8075 -43346 -6675 -43306
rect -8075 -44666 -8035 -43346
rect -6715 -44666 -6675 -43346
rect -8075 -44706 -6675 -44666
rect -5969 -43346 -4569 -43306
rect -5969 -44666 -5929 -43346
rect -4609 -44666 -4569 -43346
rect -5969 -44706 -4569 -44666
rect -3863 -43346 -2463 -43306
rect -3863 -44666 -3823 -43346
rect -2503 -44666 -2463 -43346
rect -3863 -44706 -2463 -44666
rect -1757 -43346 -357 -43306
rect -1757 -44666 -1717 -43346
rect -397 -44666 -357 -43346
rect -1757 -44706 -357 -44666
rect 349 -43346 1749 -43306
rect 349 -44666 389 -43346
rect 1709 -44666 1749 -43346
rect 349 -44706 1749 -44666
rect 2455 -43346 3855 -43306
rect 2455 -44666 2495 -43346
rect 3815 -44666 3855 -43346
rect 2455 -44706 3855 -44666
rect 4561 -43346 5961 -43306
rect 4561 -44666 4601 -43346
rect 5921 -44666 5961 -43346
rect 4561 -44706 5961 -44666
rect 6667 -43346 8067 -43306
rect 6667 -44666 6707 -43346
rect 8027 -44666 8067 -43346
rect 10962 -43342 16812 -43042
rect 17112 -43342 17162 -43042
rect 10962 -43392 17162 -43342
rect 17362 -43042 23562 -42992
rect 17362 -43342 23212 -43042
rect 23512 -43342 23562 -43042
rect 17362 -43392 23562 -43342
rect 6667 -44706 8067 -44666
rect -29135 -45346 -27735 -45306
rect -29135 -46666 -29095 -45346
rect -27775 -46666 -27735 -45346
rect -29135 -46706 -27735 -46666
rect -27029 -45346 -25629 -45306
rect -27029 -46666 -26989 -45346
rect -25669 -46666 -25629 -45346
rect -27029 -46706 -25629 -46666
rect -24923 -45346 -23523 -45306
rect -24923 -46666 -24883 -45346
rect -23563 -46666 -23523 -45346
rect -24923 -46706 -23523 -46666
rect -22817 -45346 -21417 -45306
rect -22817 -46666 -22777 -45346
rect -21457 -46666 -21417 -45346
rect -22817 -46706 -21417 -46666
rect -20711 -45346 -19311 -45306
rect -20711 -46666 -20671 -45346
rect -19351 -46666 -19311 -45346
rect -20711 -46706 -19311 -46666
rect -18605 -45346 -17205 -45306
rect -18605 -46666 -18565 -45346
rect -17245 -46666 -17205 -45346
rect -18605 -46706 -17205 -46666
rect -16499 -45346 -15099 -45306
rect -16499 -46666 -16459 -45346
rect -15139 -46666 -15099 -45346
rect -16499 -46706 -15099 -46666
rect -14393 -45346 -12993 -45306
rect -14393 -46666 -14353 -45346
rect -13033 -46666 -12993 -45346
rect -14393 -46706 -12993 -46666
rect -12287 -45346 -10887 -45306
rect -12287 -46666 -12247 -45346
rect -10927 -46666 -10887 -45346
rect -12287 -46706 -10887 -46666
rect -10181 -45346 -8781 -45306
rect -10181 -46666 -10141 -45346
rect -8821 -46666 -8781 -45346
rect -10181 -46706 -8781 -46666
rect -8075 -45346 -6675 -45306
rect -8075 -46666 -8035 -45346
rect -6715 -46666 -6675 -45346
rect -8075 -46706 -6675 -46666
rect -5969 -45346 -4569 -45306
rect -5969 -46666 -5929 -45346
rect -4609 -46666 -4569 -45346
rect -5969 -46706 -4569 -46666
rect -3863 -45346 -2463 -45306
rect -3863 -46666 -3823 -45346
rect -2503 -46666 -2463 -45346
rect -3863 -46706 -2463 -46666
rect -1757 -45346 -357 -45306
rect -1757 -46666 -1717 -45346
rect -397 -46666 -357 -45346
rect -1757 -46706 -357 -46666
rect 349 -45346 1749 -45306
rect 349 -46666 389 -45346
rect 1709 -46666 1749 -45346
rect 349 -46706 1749 -46666
rect 2455 -45346 3855 -45306
rect 2455 -46666 2495 -45346
rect 3815 -46666 3855 -45346
rect 2455 -46706 3855 -46666
rect 4561 -45346 5961 -45306
rect 4561 -46666 4601 -45346
rect 5921 -46666 5961 -45346
rect 4561 -46706 5961 -46666
rect 6667 -45346 8067 -45306
rect 6667 -46666 6707 -45346
rect 8027 -46666 8067 -45346
rect 6667 -46706 8067 -46666
rect -29135 -47346 -27735 -47306
rect -29135 -48666 -29095 -47346
rect -27775 -48666 -27735 -47346
rect -29135 -48706 -27735 -48666
rect -27029 -47346 -25629 -47306
rect -27029 -48666 -26989 -47346
rect -25669 -48666 -25629 -47346
rect -27029 -48706 -25629 -48666
rect -24923 -47346 -23523 -47306
rect -24923 -48666 -24883 -47346
rect -23563 -48666 -23523 -47346
rect -24923 -48706 -23523 -48666
rect -22817 -47346 -21417 -47306
rect -22817 -48666 -22777 -47346
rect -21457 -48666 -21417 -47346
rect -22817 -48706 -21417 -48666
rect -20711 -47346 -19311 -47306
rect -20711 -48666 -20671 -47346
rect -19351 -48666 -19311 -47346
rect -20711 -48706 -19311 -48666
rect -18605 -47346 -17205 -47306
rect -18605 -48666 -18565 -47346
rect -17245 -48666 -17205 -47346
rect -18605 -48706 -17205 -48666
rect -16499 -47346 -15099 -47306
rect -16499 -48666 -16459 -47346
rect -15139 -48666 -15099 -47346
rect -16499 -48706 -15099 -48666
rect -14393 -47346 -12993 -47306
rect -14393 -48666 -14353 -47346
rect -13033 -48666 -12993 -47346
rect -14393 -48706 -12993 -48666
rect -12287 -47346 -10887 -47306
rect -12287 -48666 -12247 -47346
rect -10927 -48666 -10887 -47346
rect -12287 -48706 -10887 -48666
rect -10181 -47346 -8781 -47306
rect -10181 -48666 -10141 -47346
rect -8821 -48666 -8781 -47346
rect -10181 -48706 -8781 -48666
rect -8075 -47346 -6675 -47306
rect -8075 -48666 -8035 -47346
rect -6715 -48666 -6675 -47346
rect -8075 -48706 -6675 -48666
rect -5969 -47346 -4569 -47306
rect -5969 -48666 -5929 -47346
rect -4609 -48666 -4569 -47346
rect -5969 -48706 -4569 -48666
rect -3863 -47346 -2463 -47306
rect -3863 -48666 -3823 -47346
rect -2503 -48666 -2463 -47346
rect -3863 -48706 -2463 -48666
rect -1757 -47346 -357 -47306
rect -1757 -48666 -1717 -47346
rect -397 -48666 -357 -47346
rect -1757 -48706 -357 -48666
rect 349 -47346 1749 -47306
rect 349 -48666 389 -47346
rect 1709 -48666 1749 -47346
rect 349 -48706 1749 -48666
rect 2455 -47346 3855 -47306
rect 2455 -48666 2495 -47346
rect 3815 -48666 3855 -47346
rect 2455 -48706 3855 -48666
rect 4561 -47346 5961 -47306
rect 4561 -48666 4601 -47346
rect 5921 -48666 5961 -47346
rect 4561 -48706 5961 -48666
rect 6667 -47346 8067 -47306
rect 6667 -48666 6707 -47346
rect 8027 -48666 8067 -47346
rect 6667 -48706 8067 -48666
rect -29135 -49346 -27735 -49306
rect -29135 -50666 -29095 -49346
rect -27775 -50666 -27735 -49346
rect -29135 -50706 -27735 -50666
rect -27029 -49346 -25629 -49306
rect -27029 -50666 -26989 -49346
rect -25669 -50666 -25629 -49346
rect -27029 -50706 -25629 -50666
rect -24923 -49346 -23523 -49306
rect -24923 -50666 -24883 -49346
rect -23563 -50666 -23523 -49346
rect -24923 -50706 -23523 -50666
rect -22817 -49346 -21417 -49306
rect -22817 -50666 -22777 -49346
rect -21457 -50666 -21417 -49346
rect -22817 -50706 -21417 -50666
rect -20711 -49346 -19311 -49306
rect -20711 -50666 -20671 -49346
rect -19351 -50666 -19311 -49346
rect -20711 -50706 -19311 -50666
rect -18605 -49346 -17205 -49306
rect -18605 -50666 -18565 -49346
rect -17245 -50666 -17205 -49346
rect -18605 -50706 -17205 -50666
rect -16499 -49346 -15099 -49306
rect -16499 -50666 -16459 -49346
rect -15139 -50666 -15099 -49346
rect -16499 -50706 -15099 -50666
rect -14393 -49346 -12993 -49306
rect -14393 -50666 -14353 -49346
rect -13033 -50666 -12993 -49346
rect -14393 -50706 -12993 -50666
rect -12287 -49346 -10887 -49306
rect -12287 -50666 -12247 -49346
rect -10927 -50666 -10887 -49346
rect -12287 -50706 -10887 -50666
rect -10181 -49346 -8781 -49306
rect -10181 -50666 -10141 -49346
rect -8821 -50666 -8781 -49346
rect -10181 -50706 -8781 -50666
rect -8075 -49346 -6675 -49306
rect -8075 -50666 -8035 -49346
rect -6715 -50666 -6675 -49346
rect -8075 -50706 -6675 -50666
rect -5969 -49346 -4569 -49306
rect -5969 -50666 -5929 -49346
rect -4609 -50666 -4569 -49346
rect -5969 -50706 -4569 -50666
rect -3863 -49346 -2463 -49306
rect -3863 -50666 -3823 -49346
rect -2503 -50666 -2463 -49346
rect -3863 -50706 -2463 -50666
rect -1757 -49346 -357 -49306
rect -1757 -50666 -1717 -49346
rect -397 -50666 -357 -49346
rect -1757 -50706 -357 -50666
rect 349 -49346 1749 -49306
rect 349 -50666 389 -49346
rect 1709 -50666 1749 -49346
rect 349 -50706 1749 -50666
rect 2455 -49346 3855 -49306
rect 2455 -50666 2495 -49346
rect 3815 -50666 3855 -49346
rect 2455 -50706 3855 -50666
rect 4561 -49346 5961 -49306
rect 4561 -50666 4601 -49346
rect 5921 -50666 5961 -49346
rect 4561 -50706 5961 -50666
rect 6667 -49346 8067 -49306
rect 6667 -50666 6707 -49346
rect 8027 -50666 8067 -49346
rect 6667 -50706 8067 -50666
rect -29135 -51346 -27735 -51306
rect -29135 -52666 -29095 -51346
rect -27775 -52666 -27735 -51346
rect -29135 -52706 -27735 -52666
rect -27029 -51346 -25629 -51306
rect -27029 -52666 -26989 -51346
rect -25669 -52666 -25629 -51346
rect -27029 -52706 -25629 -52666
rect -24923 -51346 -23523 -51306
rect -24923 -52666 -24883 -51346
rect -23563 -52666 -23523 -51346
rect -24923 -52706 -23523 -52666
rect -22817 -51346 -21417 -51306
rect -22817 -52666 -22777 -51346
rect -21457 -52666 -21417 -51346
rect -22817 -52706 -21417 -52666
rect -20711 -51346 -19311 -51306
rect -20711 -52666 -20671 -51346
rect -19351 -52666 -19311 -51346
rect -20711 -52706 -19311 -52666
rect -18605 -51346 -17205 -51306
rect -18605 -52666 -18565 -51346
rect -17245 -52666 -17205 -51346
rect -18605 -52706 -17205 -52666
rect -16499 -51346 -15099 -51306
rect -16499 -52666 -16459 -51346
rect -15139 -52666 -15099 -51346
rect -16499 -52706 -15099 -52666
rect -14393 -51346 -12993 -51306
rect -14393 -52666 -14353 -51346
rect -13033 -52666 -12993 -51346
rect -14393 -52706 -12993 -52666
rect -12287 -51346 -10887 -51306
rect -12287 -52666 -12247 -51346
rect -10927 -52666 -10887 -51346
rect -12287 -52706 -10887 -52666
rect -10181 -51346 -8781 -51306
rect -10181 -52666 -10141 -51346
rect -8821 -52666 -8781 -51346
rect -10181 -52706 -8781 -52666
rect -8075 -51346 -6675 -51306
rect -8075 -52666 -8035 -51346
rect -6715 -52666 -6675 -51346
rect -8075 -52706 -6675 -52666
rect -5969 -51346 -4569 -51306
rect -5969 -52666 -5929 -51346
rect -4609 -52666 -4569 -51346
rect -5969 -52706 -4569 -52666
rect -3863 -51346 -2463 -51306
rect -3863 -52666 -3823 -51346
rect -2503 -52666 -2463 -51346
rect -3863 -52706 -2463 -52666
rect -1757 -51346 -357 -51306
rect -1757 -52666 -1717 -51346
rect -397 -52666 -357 -51346
rect -1757 -52706 -357 -52666
rect 349 -51346 1749 -51306
rect 349 -52666 389 -51346
rect 1709 -52666 1749 -51346
rect 349 -52706 1749 -52666
rect 2455 -51346 3855 -51306
rect 2455 -52666 2495 -51346
rect 3815 -52666 3855 -51346
rect 2455 -52706 3855 -52666
rect 4561 -51346 5961 -51306
rect 4561 -52666 4601 -51346
rect 5921 -52666 5961 -51346
rect 4561 -52706 5961 -52666
rect 6667 -51346 8067 -51306
rect 6667 -52666 6707 -51346
rect 8027 -52666 8067 -51346
rect 6667 -52706 8067 -52666
rect -29135 -53346 -27735 -53306
rect -29135 -54666 -29095 -53346
rect -27775 -54666 -27735 -53346
rect -29135 -54706 -27735 -54666
rect -27029 -53346 -25629 -53306
rect -27029 -54666 -26989 -53346
rect -25669 -54666 -25629 -53346
rect -27029 -54706 -25629 -54666
rect -24923 -53346 -23523 -53306
rect -24923 -54666 -24883 -53346
rect -23563 -54666 -23523 -53346
rect -24923 -54706 -23523 -54666
rect -22817 -53346 -21417 -53306
rect -22817 -54666 -22777 -53346
rect -21457 -54666 -21417 -53346
rect -22817 -54706 -21417 -54666
rect -20711 -53346 -19311 -53306
rect -20711 -54666 -20671 -53346
rect -19351 -54666 -19311 -53346
rect -20711 -54706 -19311 -54666
rect -18605 -53346 -17205 -53306
rect -18605 -54666 -18565 -53346
rect -17245 -54666 -17205 -53346
rect -18605 -54706 -17205 -54666
rect -16499 -53346 -15099 -53306
rect -16499 -54666 -16459 -53346
rect -15139 -54666 -15099 -53346
rect -16499 -54706 -15099 -54666
rect -14393 -53346 -12993 -53306
rect -14393 -54666 -14353 -53346
rect -13033 -54666 -12993 -53346
rect -14393 -54706 -12993 -54666
rect -12287 -53346 -10887 -53306
rect -12287 -54666 -12247 -53346
rect -10927 -54666 -10887 -53346
rect -12287 -54706 -10887 -54666
rect -10181 -53346 -8781 -53306
rect -10181 -54666 -10141 -53346
rect -8821 -54666 -8781 -53346
rect -10181 -54706 -8781 -54666
rect -8075 -53346 -6675 -53306
rect -8075 -54666 -8035 -53346
rect -6715 -54666 -6675 -53346
rect -8075 -54706 -6675 -54666
rect -5969 -53346 -4569 -53306
rect -5969 -54666 -5929 -53346
rect -4609 -54666 -4569 -53346
rect -5969 -54706 -4569 -54666
rect -3863 -53346 -2463 -53306
rect -3863 -54666 -3823 -53346
rect -2503 -54666 -2463 -53346
rect -3863 -54706 -2463 -54666
rect -1757 -53346 -357 -53306
rect -1757 -54666 -1717 -53346
rect -397 -54666 -357 -53346
rect -1757 -54706 -357 -54666
rect 349 -53346 1749 -53306
rect 349 -54666 389 -53346
rect 1709 -54666 1749 -53346
rect 349 -54706 1749 -54666
rect 2455 -53346 3855 -53306
rect 2455 -54666 2495 -53346
rect 3815 -54666 3855 -53346
rect 2455 -54706 3855 -54666
rect 4561 -53346 5961 -53306
rect 4561 -54666 4601 -53346
rect 5921 -54666 5961 -53346
rect 4561 -54706 5961 -54666
rect 6667 -53346 8067 -53306
rect 6667 -54666 6707 -53346
rect 8027 -54666 8067 -53346
rect 6667 -54706 8067 -54666
rect -29135 -55346 -27735 -55306
rect -29135 -56666 -29095 -55346
rect -27775 -56666 -27735 -55346
rect -29135 -56706 -27735 -56666
rect -27029 -55346 -25629 -55306
rect -27029 -56666 -26989 -55346
rect -25669 -56666 -25629 -55346
rect -27029 -56706 -25629 -56666
rect -24923 -55346 -23523 -55306
rect -24923 -56666 -24883 -55346
rect -23563 -56666 -23523 -55346
rect -24923 -56706 -23523 -56666
rect -22817 -55346 -21417 -55306
rect -22817 -56666 -22777 -55346
rect -21457 -56666 -21417 -55346
rect -22817 -56706 -21417 -56666
rect -20711 -55346 -19311 -55306
rect -20711 -56666 -20671 -55346
rect -19351 -56666 -19311 -55346
rect -20711 -56706 -19311 -56666
rect -18605 -55346 -17205 -55306
rect -18605 -56666 -18565 -55346
rect -17245 -56666 -17205 -55346
rect -18605 -56706 -17205 -56666
rect -16499 -55346 -15099 -55306
rect -16499 -56666 -16459 -55346
rect -15139 -56666 -15099 -55346
rect -16499 -56706 -15099 -56666
rect -14393 -55346 -12993 -55306
rect -14393 -56666 -14353 -55346
rect -13033 -56666 -12993 -55346
rect -14393 -56706 -12993 -56666
rect -12287 -55346 -10887 -55306
rect -12287 -56666 -12247 -55346
rect -10927 -56666 -10887 -55346
rect -12287 -56706 -10887 -56666
rect -10181 -55346 -8781 -55306
rect -10181 -56666 -10141 -55346
rect -8821 -56666 -8781 -55346
rect -10181 -56706 -8781 -56666
rect -8075 -55346 -6675 -55306
rect -8075 -56666 -8035 -55346
rect -6715 -56666 -6675 -55346
rect -8075 -56706 -6675 -56666
rect -5969 -55346 -4569 -55306
rect -5969 -56666 -5929 -55346
rect -4609 -56666 -4569 -55346
rect -5969 -56706 -4569 -56666
rect -3863 -55346 -2463 -55306
rect -3863 -56666 -3823 -55346
rect -2503 -56666 -2463 -55346
rect -3863 -56706 -2463 -56666
rect -1757 -55346 -357 -55306
rect -1757 -56666 -1717 -55346
rect -397 -56666 -357 -55346
rect -1757 -56706 -357 -56666
rect 349 -55346 1749 -55306
rect 349 -56666 389 -55346
rect 1709 -56666 1749 -55346
rect 349 -56706 1749 -56666
rect 2455 -55346 3855 -55306
rect 2455 -56666 2495 -55346
rect 3815 -56666 3855 -55346
rect 2455 -56706 3855 -56666
rect 4561 -55346 5961 -55306
rect 4561 -56666 4601 -55346
rect 5921 -56666 5961 -55346
rect 4561 -56706 5961 -56666
rect 6667 -55346 8067 -55306
rect 6667 -56666 6707 -55346
rect 8027 -56666 8067 -55346
rect 6667 -56706 8067 -56666
rect -29135 -57346 -27735 -57306
rect -29135 -58666 -29095 -57346
rect -27775 -58666 -27735 -57346
rect -29135 -58706 -27735 -58666
rect -27029 -57346 -25629 -57306
rect -27029 -58666 -26989 -57346
rect -25669 -58666 -25629 -57346
rect -27029 -58706 -25629 -58666
rect -24923 -57346 -23523 -57306
rect -24923 -58666 -24883 -57346
rect -23563 -58666 -23523 -57346
rect -24923 -58706 -23523 -58666
rect -22817 -57346 -21417 -57306
rect -22817 -58666 -22777 -57346
rect -21457 -58666 -21417 -57346
rect -22817 -58706 -21417 -58666
rect -20711 -57346 -19311 -57306
rect -20711 -58666 -20671 -57346
rect -19351 -58666 -19311 -57346
rect -20711 -58706 -19311 -58666
rect -18605 -57346 -17205 -57306
rect -18605 -58666 -18565 -57346
rect -17245 -58666 -17205 -57346
rect -18605 -58706 -17205 -58666
rect -16499 -57346 -15099 -57306
rect -16499 -58666 -16459 -57346
rect -15139 -58666 -15099 -57346
rect -16499 -58706 -15099 -58666
rect -14393 -57346 -12993 -57306
rect -14393 -58666 -14353 -57346
rect -13033 -58666 -12993 -57346
rect -14393 -58706 -12993 -58666
rect -12287 -57346 -10887 -57306
rect -12287 -58666 -12247 -57346
rect -10927 -58666 -10887 -57346
rect -12287 -58706 -10887 -58666
rect -10181 -57346 -8781 -57306
rect -10181 -58666 -10141 -57346
rect -8821 -58666 -8781 -57346
rect -10181 -58706 -8781 -58666
rect -8075 -57346 -6675 -57306
rect -8075 -58666 -8035 -57346
rect -6715 -58666 -6675 -57346
rect -8075 -58706 -6675 -58666
rect -5969 -57346 -4569 -57306
rect -5969 -58666 -5929 -57346
rect -4609 -58666 -4569 -57346
rect -5969 -58706 -4569 -58666
rect -3863 -57346 -2463 -57306
rect -3863 -58666 -3823 -57346
rect -2503 -58666 -2463 -57346
rect -3863 -58706 -2463 -58666
rect -1757 -57346 -357 -57306
rect -1757 -58666 -1717 -57346
rect -397 -58666 -357 -57346
rect -1757 -58706 -357 -58666
rect 349 -57346 1749 -57306
rect 349 -58666 389 -57346
rect 1709 -58666 1749 -57346
rect 349 -58706 1749 -58666
rect 2455 -57346 3855 -57306
rect 2455 -58666 2495 -57346
rect 3815 -58666 3855 -57346
rect 2455 -58706 3855 -58666
rect 4561 -57346 5961 -57306
rect 4561 -58666 4601 -57346
rect 5921 -58666 5961 -57346
rect 4561 -58706 5961 -58666
rect 6667 -57346 8067 -57306
rect 6667 -58666 6707 -57346
rect 8027 -58666 8067 -57346
rect 6667 -58706 8067 -58666
rect -29135 -59346 -27735 -59306
rect -29135 -60666 -29095 -59346
rect -27775 -60666 -27735 -59346
rect -29135 -60706 -27735 -60666
rect -27029 -59346 -25629 -59306
rect -27029 -60666 -26989 -59346
rect -25669 -60666 -25629 -59346
rect -27029 -60706 -25629 -60666
rect -24923 -59346 -23523 -59306
rect -24923 -60666 -24883 -59346
rect -23563 -60666 -23523 -59346
rect -24923 -60706 -23523 -60666
rect -22817 -59346 -21417 -59306
rect -22817 -60666 -22777 -59346
rect -21457 -60666 -21417 -59346
rect -22817 -60706 -21417 -60666
rect -20711 -59346 -19311 -59306
rect -20711 -60666 -20671 -59346
rect -19351 -60666 -19311 -59346
rect -20711 -60706 -19311 -60666
rect -18605 -59346 -17205 -59306
rect -18605 -60666 -18565 -59346
rect -17245 -60666 -17205 -59346
rect -18605 -60706 -17205 -60666
rect -16499 -59346 -15099 -59306
rect -16499 -60666 -16459 -59346
rect -15139 -60666 -15099 -59346
rect -16499 -60706 -15099 -60666
rect -14393 -59346 -12993 -59306
rect -14393 -60666 -14353 -59346
rect -13033 -60666 -12993 -59346
rect -14393 -60706 -12993 -60666
rect -12287 -59346 -10887 -59306
rect -12287 -60666 -12247 -59346
rect -10927 -60666 -10887 -59346
rect -12287 -60706 -10887 -60666
rect -10181 -59346 -8781 -59306
rect -10181 -60666 -10141 -59346
rect -8821 -60666 -8781 -59346
rect -10181 -60706 -8781 -60666
rect -8075 -59346 -6675 -59306
rect -8075 -60666 -8035 -59346
rect -6715 -60666 -6675 -59346
rect -8075 -60706 -6675 -60666
rect -5969 -59346 -4569 -59306
rect -5969 -60666 -5929 -59346
rect -4609 -60666 -4569 -59346
rect -5969 -60706 -4569 -60666
rect -3863 -59346 -2463 -59306
rect -3863 -60666 -3823 -59346
rect -2503 -60666 -2463 -59346
rect -3863 -60706 -2463 -60666
rect -1757 -59346 -357 -59306
rect -1757 -60666 -1717 -59346
rect -397 -60666 -357 -59346
rect -1757 -60706 -357 -60666
rect 349 -59346 1749 -59306
rect 349 -60666 389 -59346
rect 1709 -60666 1749 -59346
rect 349 -60706 1749 -60666
rect 2455 -59346 3855 -59306
rect 2455 -60666 2495 -59346
rect 3815 -60666 3855 -59346
rect 2455 -60706 3855 -60666
rect 4561 -59346 5961 -59306
rect 4561 -60666 4601 -59346
rect 5921 -60666 5961 -59346
rect 4561 -60706 5961 -60666
rect 6667 -59346 8067 -59306
rect 6667 -60666 6707 -59346
rect 8027 -60666 8067 -59346
rect 6667 -60706 8067 -60666
rect -29135 -61346 -27735 -61306
rect -29135 -62666 -29095 -61346
rect -27775 -62666 -27735 -61346
rect -29135 -62706 -27735 -62666
rect -27029 -61346 -25629 -61306
rect -27029 -62666 -26989 -61346
rect -25669 -62666 -25629 -61346
rect -27029 -62706 -25629 -62666
rect -24923 -61346 -23523 -61306
rect -24923 -62666 -24883 -61346
rect -23563 -62666 -23523 -61346
rect -24923 -62706 -23523 -62666
rect -22817 -61346 -21417 -61306
rect -22817 -62666 -22777 -61346
rect -21457 -62666 -21417 -61346
rect -22817 -62706 -21417 -62666
rect -20711 -61346 -19311 -61306
rect -20711 -62666 -20671 -61346
rect -19351 -62666 -19311 -61346
rect -20711 -62706 -19311 -62666
rect -18605 -61346 -17205 -61306
rect -18605 -62666 -18565 -61346
rect -17245 -62666 -17205 -61346
rect -18605 -62706 -17205 -62666
rect -16499 -61346 -15099 -61306
rect -16499 -62666 -16459 -61346
rect -15139 -62666 -15099 -61346
rect -16499 -62706 -15099 -62666
rect -14393 -61346 -12993 -61306
rect -14393 -62666 -14353 -61346
rect -13033 -62666 -12993 -61346
rect -14393 -62706 -12993 -62666
rect -12287 -61346 -10887 -61306
rect -12287 -62666 -12247 -61346
rect -10927 -62666 -10887 -61346
rect -12287 -62706 -10887 -62666
rect -10181 -61346 -8781 -61306
rect -10181 -62666 -10141 -61346
rect -8821 -62666 -8781 -61346
rect -10181 -62706 -8781 -62666
rect -8075 -61346 -6675 -61306
rect -8075 -62666 -8035 -61346
rect -6715 -62666 -6675 -61346
rect -8075 -62706 -6675 -62666
rect -5969 -61346 -4569 -61306
rect -5969 -62666 -5929 -61346
rect -4609 -62666 -4569 -61346
rect -5969 -62706 -4569 -62666
rect -3863 -61346 -2463 -61306
rect -3863 -62666 -3823 -61346
rect -2503 -62666 -2463 -61346
rect -3863 -62706 -2463 -62666
rect -1757 -61346 -357 -61306
rect -1757 -62666 -1717 -61346
rect -397 -62666 -357 -61346
rect -1757 -62706 -357 -62666
rect 349 -61346 1749 -61306
rect 349 -62666 389 -61346
rect 1709 -62666 1749 -61346
rect 349 -62706 1749 -62666
rect 2455 -61346 3855 -61306
rect 2455 -62666 2495 -61346
rect 3815 -62666 3855 -61346
rect 2455 -62706 3855 -62666
rect 4561 -61346 5961 -61306
rect 4561 -62666 4601 -61346
rect 5921 -62666 5961 -61346
rect 4561 -62706 5961 -62666
rect 6667 -61346 8067 -61306
rect 6667 -62666 6707 -61346
rect 8027 -62666 8067 -61346
rect 6667 -62706 8067 -62666
<< mimcapcontact >>
rect -29095 -28666 -27775 -27346
rect -26989 -28666 -25669 -27346
rect -24883 -28666 -23563 -27346
rect -22777 -28666 -21457 -27346
rect -20671 -28666 -19351 -27346
rect -18565 -28666 -17245 -27346
rect -16459 -28666 -15139 -27346
rect -14353 -28666 -13033 -27346
rect -12247 -28666 -10927 -27346
rect -10141 -28666 -8821 -27346
rect -8035 -28666 -6715 -27346
rect -5929 -28666 -4609 -27346
rect -3823 -28666 -2503 -27346
rect -1717 -28666 -397 -27346
rect 389 -28666 1709 -27346
rect 2495 -28666 3815 -27346
rect 4601 -28666 5921 -27346
rect 6707 -28666 8027 -27346
rect -29095 -30666 -27775 -29346
rect -26989 -30666 -25669 -29346
rect -24883 -30666 -23563 -29346
rect -22777 -30666 -21457 -29346
rect -20671 -30666 -19351 -29346
rect -18565 -30666 -17245 -29346
rect -16459 -30666 -15139 -29346
rect -14353 -30666 -13033 -29346
rect -12247 -30666 -10927 -29346
rect -10141 -30666 -8821 -29346
rect -8035 -30666 -6715 -29346
rect -5929 -30666 -4609 -29346
rect -3823 -30666 -2503 -29346
rect -1717 -30666 -397 -29346
rect 389 -30666 1709 -29346
rect 2495 -30666 3815 -29346
rect 4601 -30666 5921 -29346
rect 6707 -30666 8027 -29346
rect 17312 -29342 17612 -29042
rect 23712 -29342 24012 -29042
rect -29095 -32666 -27775 -31346
rect -26989 -32666 -25669 -31346
rect -24883 -32666 -23563 -31346
rect -22777 -32666 -21457 -31346
rect -20671 -32666 -19351 -31346
rect -18565 -32666 -17245 -31346
rect -16459 -32666 -15139 -31346
rect -14353 -32666 -13033 -31346
rect -12247 -32666 -10927 -31346
rect -10141 -32666 -8821 -31346
rect -8035 -32666 -6715 -31346
rect -5929 -32666 -4609 -31346
rect -3823 -32666 -2503 -31346
rect -1717 -32666 -397 -31346
rect 389 -32666 1709 -31346
rect 2495 -32666 3815 -31346
rect 4601 -32666 5921 -31346
rect 6707 -32666 8027 -31346
rect -29095 -34666 -27775 -33346
rect -26989 -34666 -25669 -33346
rect -24883 -34666 -23563 -33346
rect -22777 -34666 -21457 -33346
rect -20671 -34666 -19351 -33346
rect -18565 -34666 -17245 -33346
rect -16459 -34666 -15139 -33346
rect -14353 -34666 -13033 -33346
rect -12247 -34666 -10927 -33346
rect -10141 -34666 -8821 -33346
rect -8035 -34666 -6715 -33346
rect -5929 -34666 -4609 -33346
rect -3823 -34666 -2503 -33346
rect -1717 -34666 -397 -33346
rect 389 -34666 1709 -33346
rect 2495 -34666 3815 -33346
rect 4601 -34666 5921 -33346
rect 6707 -34666 8027 -33346
rect -29095 -36666 -27775 -35346
rect -26989 -36666 -25669 -35346
rect -24883 -36666 -23563 -35346
rect -22777 -36666 -21457 -35346
rect -20671 -36666 -19351 -35346
rect -18565 -36666 -17245 -35346
rect -16459 -36666 -15139 -35346
rect -14353 -36666 -13033 -35346
rect -12247 -36666 -10927 -35346
rect -10141 -36666 -8821 -35346
rect -8035 -36666 -6715 -35346
rect -5929 -36666 -4609 -35346
rect -3823 -36666 -2503 -35346
rect -1717 -36666 -397 -35346
rect 389 -36666 1709 -35346
rect 2495 -36666 3815 -35346
rect 4601 -36666 5921 -35346
rect 6707 -36666 8027 -35346
rect 10826 -35824 11126 -30124
rect 17166 -35742 17466 -31042
rect 22766 -35742 23066 -31042
rect 24870 -35824 25170 -30124
rect -29095 -38666 -27775 -37346
rect -26989 -38666 -25669 -37346
rect -24883 -38666 -23563 -37346
rect -22777 -38666 -21457 -37346
rect -20671 -38666 -19351 -37346
rect -18565 -38666 -17245 -37346
rect -16459 -38666 -15139 -37346
rect -14353 -38666 -13033 -37346
rect -12247 -38666 -10927 -37346
rect -10141 -38666 -8821 -37346
rect -8035 -38666 -6715 -37346
rect -5929 -38666 -4609 -37346
rect -3823 -38666 -2503 -37346
rect -1717 -38666 -397 -37346
rect 389 -38666 1709 -37346
rect 2495 -38666 3815 -37346
rect 4601 -38666 5921 -37346
rect 6707 -38666 8027 -37346
rect -29095 -40666 -27775 -39346
rect -26989 -40666 -25669 -39346
rect -24883 -40666 -23563 -39346
rect -22777 -40666 -21457 -39346
rect -20671 -40666 -19351 -39346
rect -18565 -40666 -17245 -39346
rect -16459 -40666 -15139 -39346
rect -14353 -40666 -13033 -39346
rect -12247 -40666 -10927 -39346
rect -10141 -40666 -8821 -39346
rect -8035 -40666 -6715 -39346
rect -5929 -40666 -4609 -39346
rect -3823 -40666 -2503 -39346
rect -1717 -40666 -397 -39346
rect 389 -40666 1709 -39346
rect 2495 -40666 3815 -39346
rect 4601 -40666 5921 -39346
rect 6707 -40666 8027 -39346
rect -29095 -42666 -27775 -41346
rect -26989 -42666 -25669 -41346
rect -24883 -42666 -23563 -41346
rect -22777 -42666 -21457 -41346
rect -20671 -42666 -19351 -41346
rect -18565 -42666 -17245 -41346
rect -16459 -42666 -15139 -41346
rect -14353 -42666 -13033 -41346
rect -12247 -42666 -10927 -41346
rect -10141 -42666 -8821 -41346
rect -8035 -42666 -6715 -41346
rect -5929 -42666 -4609 -41346
rect -3823 -42666 -2503 -41346
rect -1717 -42666 -397 -41346
rect 389 -42666 1709 -41346
rect 2495 -42666 3815 -41346
rect 4601 -42666 5921 -41346
rect 6707 -42666 8027 -41346
rect 10826 -42316 11126 -36616
rect 17166 -41342 17466 -36642
rect 22766 -41342 23066 -36642
rect 24870 -42316 25170 -36616
rect -29095 -44666 -27775 -43346
rect -26989 -44666 -25669 -43346
rect -24883 -44666 -23563 -43346
rect -22777 -44666 -21457 -43346
rect -20671 -44666 -19351 -43346
rect -18565 -44666 -17245 -43346
rect -16459 -44666 -15139 -43346
rect -14353 -44666 -13033 -43346
rect -12247 -44666 -10927 -43346
rect -10141 -44666 -8821 -43346
rect -8035 -44666 -6715 -43346
rect -5929 -44666 -4609 -43346
rect -3823 -44666 -2503 -43346
rect -1717 -44666 -397 -43346
rect 389 -44666 1709 -43346
rect 2495 -44666 3815 -43346
rect 4601 -44666 5921 -43346
rect 6707 -44666 8027 -43346
rect 16812 -43342 17112 -43042
rect 23212 -43342 23512 -43042
rect -29095 -46666 -27775 -45346
rect -26989 -46666 -25669 -45346
rect -24883 -46666 -23563 -45346
rect -22777 -46666 -21457 -45346
rect -20671 -46666 -19351 -45346
rect -18565 -46666 -17245 -45346
rect -16459 -46666 -15139 -45346
rect -14353 -46666 -13033 -45346
rect -12247 -46666 -10927 -45346
rect -10141 -46666 -8821 -45346
rect -8035 -46666 -6715 -45346
rect -5929 -46666 -4609 -45346
rect -3823 -46666 -2503 -45346
rect -1717 -46666 -397 -45346
rect 389 -46666 1709 -45346
rect 2495 -46666 3815 -45346
rect 4601 -46666 5921 -45346
rect 6707 -46666 8027 -45346
rect -29095 -48666 -27775 -47346
rect -26989 -48666 -25669 -47346
rect -24883 -48666 -23563 -47346
rect -22777 -48666 -21457 -47346
rect -20671 -48666 -19351 -47346
rect -18565 -48666 -17245 -47346
rect -16459 -48666 -15139 -47346
rect -14353 -48666 -13033 -47346
rect -12247 -48666 -10927 -47346
rect -10141 -48666 -8821 -47346
rect -8035 -48666 -6715 -47346
rect -5929 -48666 -4609 -47346
rect -3823 -48666 -2503 -47346
rect -1717 -48666 -397 -47346
rect 389 -48666 1709 -47346
rect 2495 -48666 3815 -47346
rect 4601 -48666 5921 -47346
rect 6707 -48666 8027 -47346
rect -29095 -50666 -27775 -49346
rect -26989 -50666 -25669 -49346
rect -24883 -50666 -23563 -49346
rect -22777 -50666 -21457 -49346
rect -20671 -50666 -19351 -49346
rect -18565 -50666 -17245 -49346
rect -16459 -50666 -15139 -49346
rect -14353 -50666 -13033 -49346
rect -12247 -50666 -10927 -49346
rect -10141 -50666 -8821 -49346
rect -8035 -50666 -6715 -49346
rect -5929 -50666 -4609 -49346
rect -3823 -50666 -2503 -49346
rect -1717 -50666 -397 -49346
rect 389 -50666 1709 -49346
rect 2495 -50666 3815 -49346
rect 4601 -50666 5921 -49346
rect 6707 -50666 8027 -49346
rect -29095 -52666 -27775 -51346
rect -26989 -52666 -25669 -51346
rect -24883 -52666 -23563 -51346
rect -22777 -52666 -21457 -51346
rect -20671 -52666 -19351 -51346
rect -18565 -52666 -17245 -51346
rect -16459 -52666 -15139 -51346
rect -14353 -52666 -13033 -51346
rect -12247 -52666 -10927 -51346
rect -10141 -52666 -8821 -51346
rect -8035 -52666 -6715 -51346
rect -5929 -52666 -4609 -51346
rect -3823 -52666 -2503 -51346
rect -1717 -52666 -397 -51346
rect 389 -52666 1709 -51346
rect 2495 -52666 3815 -51346
rect 4601 -52666 5921 -51346
rect 6707 -52666 8027 -51346
rect -29095 -54666 -27775 -53346
rect -26989 -54666 -25669 -53346
rect -24883 -54666 -23563 -53346
rect -22777 -54666 -21457 -53346
rect -20671 -54666 -19351 -53346
rect -18565 -54666 -17245 -53346
rect -16459 -54666 -15139 -53346
rect -14353 -54666 -13033 -53346
rect -12247 -54666 -10927 -53346
rect -10141 -54666 -8821 -53346
rect -8035 -54666 -6715 -53346
rect -5929 -54666 -4609 -53346
rect -3823 -54666 -2503 -53346
rect -1717 -54666 -397 -53346
rect 389 -54666 1709 -53346
rect 2495 -54666 3815 -53346
rect 4601 -54666 5921 -53346
rect 6707 -54666 8027 -53346
rect -29095 -56666 -27775 -55346
rect -26989 -56666 -25669 -55346
rect -24883 -56666 -23563 -55346
rect -22777 -56666 -21457 -55346
rect -20671 -56666 -19351 -55346
rect -18565 -56666 -17245 -55346
rect -16459 -56666 -15139 -55346
rect -14353 -56666 -13033 -55346
rect -12247 -56666 -10927 -55346
rect -10141 -56666 -8821 -55346
rect -8035 -56666 -6715 -55346
rect -5929 -56666 -4609 -55346
rect -3823 -56666 -2503 -55346
rect -1717 -56666 -397 -55346
rect 389 -56666 1709 -55346
rect 2495 -56666 3815 -55346
rect 4601 -56666 5921 -55346
rect 6707 -56666 8027 -55346
rect -29095 -58666 -27775 -57346
rect -26989 -58666 -25669 -57346
rect -24883 -58666 -23563 -57346
rect -22777 -58666 -21457 -57346
rect -20671 -58666 -19351 -57346
rect -18565 -58666 -17245 -57346
rect -16459 -58666 -15139 -57346
rect -14353 -58666 -13033 -57346
rect -12247 -58666 -10927 -57346
rect -10141 -58666 -8821 -57346
rect -8035 -58666 -6715 -57346
rect -5929 -58666 -4609 -57346
rect -3823 -58666 -2503 -57346
rect -1717 -58666 -397 -57346
rect 389 -58666 1709 -57346
rect 2495 -58666 3815 -57346
rect 4601 -58666 5921 -57346
rect 6707 -58666 8027 -57346
rect -29095 -60666 -27775 -59346
rect -26989 -60666 -25669 -59346
rect -24883 -60666 -23563 -59346
rect -22777 -60666 -21457 -59346
rect -20671 -60666 -19351 -59346
rect -18565 -60666 -17245 -59346
rect -16459 -60666 -15139 -59346
rect -14353 -60666 -13033 -59346
rect -12247 -60666 -10927 -59346
rect -10141 -60666 -8821 -59346
rect -8035 -60666 -6715 -59346
rect -5929 -60666 -4609 -59346
rect -3823 -60666 -2503 -59346
rect -1717 -60666 -397 -59346
rect 389 -60666 1709 -59346
rect 2495 -60666 3815 -59346
rect 4601 -60666 5921 -59346
rect 6707 -60666 8027 -59346
rect -29095 -62666 -27775 -61346
rect -26989 -62666 -25669 -61346
rect -24883 -62666 -23563 -61346
rect -22777 -62666 -21457 -61346
rect -20671 -62666 -19351 -61346
rect -18565 -62666 -17245 -61346
rect -16459 -62666 -15139 -61346
rect -14353 -62666 -13033 -61346
rect -12247 -62666 -10927 -61346
rect -10141 -62666 -8821 -61346
rect -8035 -62666 -6715 -61346
rect -5929 -62666 -4609 -61346
rect -3823 -62666 -2503 -61346
rect -1717 -62666 -397 -61346
rect 389 -62666 1709 -61346
rect 2495 -62666 3815 -61346
rect 4601 -62666 5921 -61346
rect 6707 -62666 8027 -61346
<< metal4 >>
rect -29096 -27346 -27774 -27345
rect -29096 -28666 -29095 -27346
rect -27775 -27958 -27774 -27346
rect -27636 -27370 -27540 -27344
rect -27636 -27958 -27620 -27370
rect -27775 -28058 -27620 -27958
rect -27775 -28666 -27774 -28058
rect -29096 -28667 -27774 -28666
rect -27640 -28652 -27620 -28058
rect -27556 -27958 -27540 -27370
rect -26990 -27346 -25668 -27345
rect -26990 -27958 -26989 -27346
rect -27556 -28058 -26989 -27958
rect -27556 -28652 -27540 -28058
rect -28470 -28948 -28370 -28667
rect -27640 -28948 -27540 -28652
rect -26990 -28666 -26989 -28058
rect -25669 -27958 -25668 -27346
rect -25530 -27370 -25434 -27344
rect -25530 -27958 -25514 -27370
rect -25669 -28058 -25514 -27958
rect -25669 -28666 -25668 -28058
rect -26990 -28667 -25668 -28666
rect -25530 -28652 -25514 -28058
rect -25450 -27958 -25434 -27370
rect -24884 -27346 -23562 -27345
rect -24884 -27958 -24883 -27346
rect -25450 -28058 -24883 -27958
rect -25450 -28652 -25434 -28058
rect -26348 -28948 -26248 -28667
rect -25530 -28668 -25434 -28652
rect -24884 -28666 -24883 -28058
rect -23563 -27958 -23562 -27346
rect -23424 -27370 -23328 -27344
rect -23424 -27958 -23408 -27370
rect -23563 -28058 -23408 -27958
rect -23563 -28666 -23562 -28058
rect -24884 -28667 -23562 -28666
rect -23424 -28652 -23408 -28058
rect -23344 -27958 -23328 -27370
rect -22778 -27346 -21456 -27345
rect -22778 -27958 -22777 -27346
rect -23344 -28058 -22777 -27958
rect -23344 -28652 -23328 -28058
rect -24242 -28948 -24142 -28667
rect -23424 -28668 -23328 -28652
rect -22778 -28666 -22777 -28058
rect -21457 -27958 -21456 -27346
rect -21318 -27370 -21222 -27344
rect -21318 -27958 -21302 -27370
rect -21457 -28058 -21302 -27958
rect -21457 -28666 -21456 -28058
rect -22778 -28667 -21456 -28666
rect -21318 -28652 -21302 -28058
rect -21238 -27958 -21222 -27370
rect -20672 -27346 -19350 -27345
rect -20672 -27958 -20671 -27346
rect -21238 -28058 -20671 -27958
rect -21238 -28652 -21222 -28058
rect -22136 -28948 -22036 -28667
rect -21318 -28668 -21222 -28652
rect -20672 -28666 -20671 -28058
rect -19351 -27958 -19350 -27346
rect -19212 -27370 -19116 -27344
rect -19212 -27958 -19196 -27370
rect -19351 -28058 -19196 -27958
rect -19351 -28666 -19350 -28058
rect -20672 -28667 -19350 -28666
rect -19212 -28652 -19196 -28058
rect -19132 -27958 -19116 -27370
rect -18566 -27346 -17244 -27345
rect -18566 -27958 -18565 -27346
rect -19132 -28058 -18565 -27958
rect -19132 -28652 -19116 -28058
rect -20030 -28948 -19930 -28667
rect -19212 -28668 -19116 -28652
rect -18566 -28666 -18565 -28058
rect -17245 -27958 -17244 -27346
rect -17106 -27370 -17010 -27344
rect -17106 -27958 -17090 -27370
rect -17245 -28058 -17090 -27958
rect -17245 -28666 -17244 -28058
rect -18566 -28667 -17244 -28666
rect -17106 -28652 -17090 -28058
rect -17026 -27958 -17010 -27370
rect -16460 -27346 -15138 -27345
rect -16460 -27958 -16459 -27346
rect -17026 -28058 -16459 -27958
rect -17026 -28652 -17010 -28058
rect -17924 -28948 -17824 -28667
rect -17106 -28668 -17010 -28652
rect -16460 -28666 -16459 -28058
rect -15139 -27958 -15138 -27346
rect -15000 -27370 -14904 -27344
rect -15000 -27958 -14984 -27370
rect -15139 -28058 -14984 -27958
rect -15139 -28666 -15138 -28058
rect -16460 -28667 -15138 -28666
rect -15000 -28652 -14984 -28058
rect -14920 -27958 -14904 -27370
rect -14354 -27346 -13032 -27345
rect -14354 -27958 -14353 -27346
rect -14920 -28058 -14353 -27958
rect -14920 -28652 -14904 -28058
rect -15818 -28948 -15718 -28667
rect -15000 -28668 -14904 -28652
rect -14354 -28666 -14353 -28058
rect -13033 -27958 -13032 -27346
rect -12894 -27370 -12798 -27344
rect -12894 -27958 -12878 -27370
rect -13033 -28058 -12878 -27958
rect -13033 -28666 -13032 -28058
rect -14354 -28667 -13032 -28666
rect -12894 -28652 -12878 -28058
rect -12814 -27958 -12798 -27370
rect -12248 -27346 -10926 -27345
rect -12248 -27958 -12247 -27346
rect -12814 -28058 -12247 -27958
rect -12814 -28652 -12798 -28058
rect -13712 -28948 -13612 -28667
rect -12894 -28668 -12798 -28652
rect -12248 -28666 -12247 -28058
rect -10927 -27958 -10926 -27346
rect -10788 -27370 -10692 -27344
rect -10788 -27958 -10772 -27370
rect -10927 -28058 -10772 -27958
rect -10927 -28666 -10926 -28058
rect -12248 -28667 -10926 -28666
rect -10788 -28652 -10772 -28058
rect -10708 -27958 -10692 -27370
rect -10142 -27346 -8820 -27345
rect -10142 -27958 -10141 -27346
rect -10708 -28058 -10141 -27958
rect -10708 -28652 -10692 -28058
rect -11606 -28948 -11506 -28667
rect -10788 -28668 -10692 -28652
rect -10142 -28666 -10141 -28058
rect -8821 -27958 -8820 -27346
rect -8682 -27370 -8586 -27344
rect -8682 -27958 -8666 -27370
rect -8821 -28058 -8666 -27958
rect -8821 -28666 -8820 -28058
rect -10142 -28667 -8820 -28666
rect -8682 -28652 -8666 -28058
rect -8602 -27958 -8586 -27370
rect -8036 -27346 -6714 -27345
rect -8036 -27958 -8035 -27346
rect -8602 -28058 -8035 -27958
rect -8602 -28652 -8586 -28058
rect -9500 -28948 -9400 -28667
rect -8682 -28668 -8586 -28652
rect -8036 -28666 -8035 -28058
rect -6715 -27958 -6714 -27346
rect -6576 -27370 -6480 -27344
rect -6576 -27958 -6560 -27370
rect -6715 -28058 -6560 -27958
rect -6715 -28666 -6714 -28058
rect -8036 -28667 -6714 -28666
rect -6576 -28652 -6560 -28058
rect -6496 -27958 -6480 -27370
rect -5930 -27346 -4608 -27345
rect -5930 -27958 -5929 -27346
rect -6496 -28058 -5929 -27958
rect -6496 -28652 -6480 -28058
rect -7394 -28948 -7294 -28667
rect -6576 -28668 -6480 -28652
rect -5930 -28666 -5929 -28058
rect -4609 -27958 -4608 -27346
rect -4470 -27370 -4374 -27344
rect -4470 -27958 -4454 -27370
rect -4609 -28058 -4454 -27958
rect -4609 -28666 -4608 -28058
rect -5930 -28667 -4608 -28666
rect -4470 -28652 -4454 -28058
rect -4390 -27958 -4374 -27370
rect -3824 -27346 -2502 -27345
rect -3824 -27958 -3823 -27346
rect -4390 -28058 -3823 -27958
rect -4390 -28652 -4374 -28058
rect -5288 -28948 -5188 -28667
rect -4470 -28668 -4374 -28652
rect -3824 -28666 -3823 -28058
rect -2503 -27958 -2502 -27346
rect -2364 -27370 -2268 -27344
rect -2364 -27958 -2348 -27370
rect -2503 -28058 -2348 -27958
rect -2503 -28666 -2502 -28058
rect -3824 -28667 -2502 -28666
rect -2364 -28652 -2348 -28058
rect -2284 -27958 -2268 -27370
rect -1718 -27346 -396 -27345
rect -1718 -27958 -1717 -27346
rect -2284 -28058 -1717 -27958
rect -2284 -28652 -2268 -28058
rect -3182 -28948 -3082 -28667
rect -2364 -28668 -2268 -28652
rect -1718 -28666 -1717 -28058
rect -397 -27958 -396 -27346
rect -258 -27370 -162 -27344
rect -258 -27958 -242 -27370
rect -397 -28058 -242 -27958
rect -397 -28666 -396 -28058
rect -1718 -28667 -396 -28666
rect -258 -28652 -242 -28058
rect -178 -27958 -162 -27370
rect 388 -27346 1710 -27345
rect 388 -27958 389 -27346
rect -178 -28058 389 -27958
rect -178 -28652 -162 -28058
rect -1076 -28948 -976 -28667
rect -258 -28668 -162 -28652
rect 388 -28666 389 -28058
rect 1709 -27958 1710 -27346
rect 1848 -27370 1944 -27344
rect 1848 -27958 1864 -27370
rect 1709 -28058 1864 -27958
rect 1709 -28666 1710 -28058
rect 388 -28667 1710 -28666
rect 1848 -28652 1864 -28058
rect 1928 -27958 1944 -27370
rect 2494 -27346 3816 -27345
rect 2494 -27958 2495 -27346
rect 1928 -28058 2495 -27958
rect 1928 -28652 1944 -28058
rect 1030 -28948 1130 -28667
rect 1848 -28668 1944 -28652
rect 2494 -28666 2495 -28058
rect 3815 -27958 3816 -27346
rect 3954 -27370 4050 -27344
rect 3954 -27958 3970 -27370
rect 3815 -28058 3970 -27958
rect 3815 -28666 3816 -28058
rect 2494 -28667 3816 -28666
rect 3954 -28652 3970 -28058
rect 4034 -27958 4050 -27370
rect 4600 -27346 5922 -27345
rect 4600 -27958 4601 -27346
rect 4034 -28058 4601 -27958
rect 4034 -28652 4050 -28058
rect 3136 -28948 3236 -28667
rect 3954 -28668 4050 -28652
rect 4600 -28666 4601 -28058
rect 5921 -27958 5922 -27346
rect 6060 -27370 6156 -27344
rect 6060 -27958 6076 -27370
rect 5921 -28058 6076 -27958
rect 5921 -28666 5922 -28058
rect 4600 -28667 5922 -28666
rect 6060 -28652 6076 -28058
rect 6140 -27958 6156 -27370
rect 6706 -27346 8028 -27345
rect 6706 -27958 6707 -27346
rect 6140 -28058 6707 -27958
rect 6140 -28652 6156 -28058
rect 5242 -28948 5342 -28667
rect 6060 -28668 6156 -28652
rect 6706 -28666 6707 -28058
rect 8027 -27942 8028 -27346
rect 8166 -27370 8262 -27344
rect 8166 -27942 8182 -27370
rect 8027 -28058 8182 -27942
rect 8027 -28666 8028 -28058
rect 6706 -28667 8028 -28666
rect 8160 -28652 8182 -28058
rect 8246 -27958 8262 -27370
rect 8246 -28058 8276 -27958
rect 8246 -28652 8262 -28058
rect 9588 -27762 50552 -27578
rect 9588 -28062 25928 -27762
rect 26528 -28062 49560 -27762
rect 50160 -28062 50552 -27762
rect 9588 -28144 50552 -28062
rect 9588 -28358 29505 -28144
rect 46290 -28358 50552 -28144
rect 9588 -28378 50552 -28358
rect 7368 -28948 7468 -28667
rect 8160 -28668 8262 -28652
rect 8160 -28948 8260 -28668
rect -28470 -29048 8260 -28948
rect -28470 -29345 -28370 -29048
rect -29096 -29346 -27774 -29345
rect -29096 -30666 -29095 -29346
rect -27775 -29938 -27774 -29346
rect -27640 -29370 -27540 -29048
rect -26348 -29345 -26248 -29048
rect -27640 -29938 -27620 -29370
rect -27775 -30038 -27620 -29938
rect -27775 -30666 -27774 -30038
rect -29096 -30667 -27774 -30666
rect -27640 -30652 -27620 -30038
rect -27556 -30652 -27540 -29370
rect -28470 -30948 -28370 -30667
rect -27640 -30948 -27540 -30652
rect -26990 -29346 -25668 -29345
rect -26990 -30666 -26989 -29346
rect -25669 -30666 -25668 -29346
rect -26990 -30667 -25668 -30666
rect -25530 -29370 -25434 -29344
rect -24242 -29345 -24142 -29048
rect -25530 -30652 -25514 -29370
rect -25450 -30652 -25434 -29370
rect -26348 -30948 -26248 -30667
rect -25530 -30668 -25434 -30652
rect -24884 -29346 -23562 -29345
rect -24884 -30666 -24883 -29346
rect -23563 -30666 -23562 -29346
rect -24884 -30667 -23562 -30666
rect -23424 -29370 -23328 -29344
rect -22136 -29345 -22036 -29048
rect -23424 -30652 -23408 -29370
rect -23344 -30652 -23328 -29370
rect -24242 -30948 -24142 -30667
rect -23424 -30668 -23328 -30652
rect -22778 -29346 -21456 -29345
rect -22778 -30666 -22777 -29346
rect -21457 -30666 -21456 -29346
rect -22778 -30667 -21456 -30666
rect -21318 -29370 -21222 -29344
rect -20030 -29345 -19930 -29048
rect -21318 -30652 -21302 -29370
rect -21238 -30652 -21222 -29370
rect -22136 -30948 -22036 -30667
rect -21318 -30668 -21222 -30652
rect -20672 -29346 -19350 -29345
rect -20672 -30666 -20671 -29346
rect -19351 -30666 -19350 -29346
rect -20672 -30667 -19350 -30666
rect -19212 -29370 -19116 -29344
rect -17924 -29345 -17824 -29048
rect -19212 -30652 -19196 -29370
rect -19132 -30652 -19116 -29370
rect -20030 -30948 -19930 -30667
rect -19212 -30668 -19116 -30652
rect -18566 -29346 -17244 -29345
rect -18566 -30666 -18565 -29346
rect -17245 -30666 -17244 -29346
rect -18566 -30667 -17244 -30666
rect -17106 -29370 -17010 -29344
rect -15818 -29345 -15718 -29048
rect -17106 -30652 -17090 -29370
rect -17026 -30652 -17010 -29370
rect -17924 -30948 -17824 -30667
rect -17106 -30668 -17010 -30652
rect -16460 -29346 -15138 -29345
rect -16460 -30666 -16459 -29346
rect -15139 -30666 -15138 -29346
rect -16460 -30667 -15138 -30666
rect -15000 -29370 -14904 -29344
rect -13712 -29345 -13612 -29048
rect -15000 -30652 -14984 -29370
rect -14920 -30652 -14904 -29370
rect -15818 -30948 -15718 -30667
rect -15000 -30668 -14904 -30652
rect -14354 -29346 -13032 -29345
rect -14354 -30666 -14353 -29346
rect -13033 -30666 -13032 -29346
rect -14354 -30667 -13032 -30666
rect -12894 -29370 -12798 -29344
rect -11606 -29345 -11506 -29048
rect -12894 -30652 -12878 -29370
rect -12814 -30652 -12798 -29370
rect -13712 -30948 -13612 -30667
rect -12894 -30668 -12798 -30652
rect -12248 -29346 -10926 -29345
rect -12248 -30666 -12247 -29346
rect -10927 -30666 -10926 -29346
rect -12248 -30667 -10926 -30666
rect -10788 -29370 -10692 -29344
rect -9500 -29345 -9400 -29048
rect -10788 -30652 -10772 -29370
rect -10708 -30652 -10692 -29370
rect -11606 -30948 -11506 -30667
rect -10788 -30668 -10692 -30652
rect -10142 -29346 -8820 -29345
rect -10142 -30666 -10141 -29346
rect -8821 -30666 -8820 -29346
rect -10142 -30667 -8820 -30666
rect -8682 -29370 -8586 -29344
rect -7394 -29345 -7294 -29048
rect -8682 -30652 -8666 -29370
rect -8602 -30652 -8586 -29370
rect -9500 -30948 -9400 -30667
rect -8682 -30668 -8586 -30652
rect -8036 -29346 -6714 -29345
rect -8036 -30666 -8035 -29346
rect -6715 -30666 -6714 -29346
rect -8036 -30667 -6714 -30666
rect -6576 -29370 -6480 -29344
rect -5288 -29345 -5188 -29048
rect -6576 -30652 -6560 -29370
rect -6496 -30652 -6480 -29370
rect -7394 -30948 -7294 -30667
rect -6576 -30668 -6480 -30652
rect -5930 -29346 -4608 -29345
rect -5930 -30666 -5929 -29346
rect -4609 -30666 -4608 -29346
rect -5930 -30667 -4608 -30666
rect -4470 -29370 -4374 -29344
rect -3182 -29345 -3082 -29048
rect -4470 -30652 -4454 -29370
rect -4390 -30652 -4374 -29370
rect -5288 -30948 -5188 -30667
rect -4470 -30668 -4374 -30652
rect -3824 -29346 -2502 -29345
rect -3824 -30666 -3823 -29346
rect -2503 -30666 -2502 -29346
rect -3824 -30667 -2502 -30666
rect -2364 -29370 -2268 -29344
rect -1076 -29345 -976 -29048
rect -2364 -30652 -2348 -29370
rect -2284 -30652 -2268 -29370
rect -3182 -30948 -3082 -30667
rect -2364 -30668 -2268 -30652
rect -1718 -29346 -396 -29345
rect -1718 -30666 -1717 -29346
rect -397 -30666 -396 -29346
rect -1718 -30667 -396 -30666
rect -258 -29370 -162 -29344
rect 1030 -29345 1130 -29048
rect -258 -30652 -242 -29370
rect -178 -30652 -162 -29370
rect -1076 -30948 -976 -30667
rect -258 -30668 -162 -30652
rect 388 -29346 1710 -29345
rect 388 -30666 389 -29346
rect 1709 -30666 1710 -29346
rect 388 -30667 1710 -30666
rect 1848 -29370 1944 -29344
rect 3136 -29345 3236 -29048
rect 1848 -30652 1864 -29370
rect 1928 -30652 1944 -29370
rect 1030 -30948 1130 -30667
rect 1848 -30668 1944 -30652
rect 2494 -29346 3816 -29345
rect 2494 -30666 2495 -29346
rect 3815 -30666 3816 -29346
rect 2494 -30667 3816 -30666
rect 3954 -29370 4050 -29344
rect 5242 -29345 5342 -29048
rect 3954 -30652 3970 -29370
rect 4034 -30652 4050 -29370
rect 3136 -30948 3236 -30667
rect 3954 -30668 4050 -30652
rect 4600 -29346 5922 -29345
rect 4600 -30666 4601 -29346
rect 5921 -30666 5922 -29346
rect 4600 -30667 5922 -30666
rect 6060 -29370 6156 -29344
rect 7368 -29345 7468 -29048
rect 8160 -29344 8260 -29048
rect 10276 -29038 25316 -28892
rect 10276 -29042 24470 -29038
rect 10276 -29048 17312 -29042
rect 6060 -30652 6076 -29370
rect 6140 -30652 6156 -29370
rect 5242 -30948 5342 -30667
rect 6060 -30668 6156 -30652
rect 6706 -29346 8028 -29345
rect 6706 -30666 6707 -29346
rect 8027 -29942 8028 -29346
rect 8160 -29370 8262 -29344
rect 8160 -29942 8182 -29370
rect 8027 -30042 8182 -29942
rect 8027 -30666 8028 -30042
rect 6706 -30667 8028 -30666
rect 8160 -30652 8182 -30042
rect 8246 -30652 8262 -29370
rect 7368 -30948 7468 -30667
rect 8160 -30668 8262 -30652
rect 10276 -29738 10428 -29048
rect 11124 -29342 17312 -29048
rect 17612 -29342 23712 -29042
rect 24012 -29342 24470 -29042
rect 11124 -29736 24470 -29342
rect 25160 -29736 25316 -29038
rect 11124 -29738 25316 -29736
rect 10276 -30068 25316 -29738
rect 10276 -30124 11458 -30068
rect 8160 -30948 8260 -30668
rect -28470 -31048 8260 -30948
rect -28470 -31345 -28370 -31048
rect -29096 -31346 -27774 -31345
rect -29096 -32666 -29095 -31346
rect -27775 -31938 -27774 -31346
rect -27640 -31370 -27540 -31048
rect -26348 -31345 -26248 -31048
rect -27640 -31938 -27620 -31370
rect -27775 -32038 -27620 -31938
rect -27775 -32666 -27774 -32038
rect -29096 -32667 -27774 -32666
rect -27640 -32652 -27620 -32038
rect -27556 -32652 -27540 -31370
rect -28470 -32948 -28370 -32667
rect -27640 -32948 -27540 -32652
rect -26990 -31346 -25668 -31345
rect -26990 -32666 -26989 -31346
rect -25669 -32666 -25668 -31346
rect -26990 -32667 -25668 -32666
rect -25530 -31370 -25434 -31344
rect -24242 -31345 -24142 -31048
rect -25530 -32652 -25514 -31370
rect -25450 -32652 -25434 -31370
rect -26348 -32948 -26248 -32667
rect -25530 -32668 -25434 -32652
rect -24884 -31346 -23562 -31345
rect -24884 -32666 -24883 -31346
rect -23563 -32666 -23562 -31346
rect -24884 -32667 -23562 -32666
rect -23424 -31370 -23328 -31344
rect -22136 -31345 -22036 -31048
rect -23424 -32652 -23408 -31370
rect -23344 -32652 -23328 -31370
rect -24242 -32948 -24142 -32667
rect -23424 -32668 -23328 -32652
rect -22778 -31346 -21456 -31345
rect -22778 -32666 -22777 -31346
rect -21457 -32666 -21456 -31346
rect -22778 -32667 -21456 -32666
rect -21318 -31370 -21222 -31344
rect -20030 -31345 -19930 -31048
rect -21318 -32652 -21302 -31370
rect -21238 -32652 -21222 -31370
rect -22136 -32948 -22036 -32667
rect -21318 -32668 -21222 -32652
rect -20672 -31346 -19350 -31345
rect -20672 -32666 -20671 -31346
rect -19351 -32666 -19350 -31346
rect -20672 -32667 -19350 -32666
rect -19212 -31370 -19116 -31344
rect -17924 -31345 -17824 -31048
rect -19212 -32652 -19196 -31370
rect -19132 -32652 -19116 -31370
rect -20030 -32948 -19930 -32667
rect -19212 -32668 -19116 -32652
rect -18566 -31346 -17244 -31345
rect -18566 -32666 -18565 -31346
rect -17245 -32666 -17244 -31346
rect -18566 -32667 -17244 -32666
rect -17106 -31370 -17010 -31344
rect -15818 -31345 -15718 -31048
rect -17106 -32652 -17090 -31370
rect -17026 -32652 -17010 -31370
rect -17924 -32948 -17824 -32667
rect -17106 -32668 -17010 -32652
rect -16460 -31346 -15138 -31345
rect -16460 -32666 -16459 -31346
rect -15139 -32666 -15138 -31346
rect -16460 -32667 -15138 -32666
rect -15000 -31370 -14904 -31344
rect -13712 -31345 -13612 -31048
rect -15000 -32652 -14984 -31370
rect -14920 -32652 -14904 -31370
rect -15818 -32948 -15718 -32667
rect -15000 -32668 -14904 -32652
rect -14354 -31346 -13032 -31345
rect -14354 -32666 -14353 -31346
rect -13033 -32666 -13032 -31346
rect -14354 -32667 -13032 -32666
rect -12894 -31370 -12798 -31344
rect -11606 -31345 -11506 -31048
rect -12894 -32652 -12878 -31370
rect -12814 -32652 -12798 -31370
rect -13712 -32948 -13612 -32667
rect -12894 -32668 -12798 -32652
rect -12248 -31346 -10926 -31345
rect -12248 -32666 -12247 -31346
rect -10927 -32666 -10926 -31346
rect -12248 -32667 -10926 -32666
rect -10788 -31370 -10692 -31344
rect -9500 -31345 -9400 -31048
rect -10788 -32652 -10772 -31370
rect -10708 -32652 -10692 -31370
rect -11606 -32948 -11506 -32667
rect -10788 -32668 -10692 -32652
rect -10142 -31346 -8820 -31345
rect -10142 -32666 -10141 -31346
rect -8821 -32666 -8820 -31346
rect -10142 -32667 -8820 -32666
rect -8682 -31370 -8586 -31344
rect -7394 -31345 -7294 -31048
rect -8682 -32652 -8666 -31370
rect -8602 -32652 -8586 -31370
rect -9500 -32948 -9400 -32667
rect -8682 -32668 -8586 -32652
rect -8036 -31346 -6714 -31345
rect -8036 -32666 -8035 -31346
rect -6715 -32666 -6714 -31346
rect -8036 -32667 -6714 -32666
rect -6576 -31370 -6480 -31344
rect -5288 -31345 -5188 -31048
rect -6576 -32652 -6560 -31370
rect -6496 -32652 -6480 -31370
rect -7394 -32948 -7294 -32667
rect -6576 -32668 -6480 -32652
rect -5930 -31346 -4608 -31345
rect -5930 -32666 -5929 -31346
rect -4609 -32666 -4608 -31346
rect -5930 -32667 -4608 -32666
rect -4470 -31370 -4374 -31344
rect -3182 -31345 -3082 -31048
rect -4470 -32652 -4454 -31370
rect -4390 -32652 -4374 -31370
rect -5288 -32948 -5188 -32667
rect -4470 -32668 -4374 -32652
rect -3824 -31346 -2502 -31345
rect -3824 -32666 -3823 -31346
rect -2503 -32666 -2502 -31346
rect -3824 -32667 -2502 -32666
rect -2364 -31370 -2268 -31344
rect -1076 -31345 -976 -31048
rect -2364 -32652 -2348 -31370
rect -2284 -32652 -2268 -31370
rect -3182 -32948 -3082 -32667
rect -2364 -32668 -2268 -32652
rect -1718 -31346 -396 -31345
rect -1718 -32666 -1717 -31346
rect -397 -32666 -396 -31346
rect -1718 -32667 -396 -32666
rect -258 -31370 -162 -31344
rect 1030 -31345 1130 -31048
rect -258 -32652 -242 -31370
rect -178 -32652 -162 -31370
rect -1076 -32948 -976 -32667
rect -258 -32668 -162 -32652
rect 388 -31346 1710 -31345
rect 388 -32666 389 -31346
rect 1709 -32666 1710 -31346
rect 388 -32667 1710 -32666
rect 1848 -31370 1944 -31344
rect 3136 -31345 3236 -31048
rect 1848 -32652 1864 -31370
rect 1928 -32652 1944 -31370
rect 1030 -32948 1130 -32667
rect 1848 -32668 1944 -32652
rect 2494 -31346 3816 -31345
rect 2494 -32666 2495 -31346
rect 3815 -32666 3816 -31346
rect 2494 -32667 3816 -32666
rect 3954 -31370 4050 -31344
rect 5242 -31345 5342 -31048
rect 3954 -32652 3970 -31370
rect 4034 -32652 4050 -31370
rect 3136 -32948 3236 -32667
rect 3954 -32668 4050 -32652
rect 4600 -31346 5922 -31345
rect 4600 -32666 4601 -31346
rect 5921 -32666 5922 -31346
rect 4600 -32667 5922 -32666
rect 6060 -31370 6156 -31344
rect 7368 -31345 7468 -31048
rect 8160 -31344 8260 -31048
rect 6060 -32652 6076 -31370
rect 6140 -32652 6156 -31370
rect 5242 -32948 5342 -32667
rect 6060 -32668 6156 -32652
rect 6706 -31346 8028 -31345
rect 6706 -32666 6707 -31346
rect 8027 -31942 8028 -31346
rect 8160 -31370 8262 -31344
rect 8160 -31942 8182 -31370
rect 8027 -32042 8182 -31942
rect 8027 -32666 8028 -32042
rect 6706 -32667 8028 -32666
rect 8160 -32652 8182 -32042
rect 8246 -32652 8262 -31370
rect 7368 -32948 7468 -32667
rect 8160 -32668 8262 -32652
rect 8160 -32948 8260 -32668
rect -28470 -33048 8260 -32948
rect -28470 -33345 -28370 -33048
rect -29096 -33346 -27774 -33345
rect -29096 -34666 -29095 -33346
rect -27775 -33938 -27774 -33346
rect -27640 -33370 -27540 -33048
rect -26348 -33345 -26248 -33048
rect -27640 -33938 -27620 -33370
rect -27775 -34038 -27620 -33938
rect -27775 -34666 -27774 -34038
rect -29096 -34667 -27774 -34666
rect -27640 -34652 -27620 -34038
rect -27556 -34652 -27540 -33370
rect -28470 -34948 -28370 -34667
rect -27640 -34948 -27540 -34652
rect -26990 -33346 -25668 -33345
rect -26990 -34666 -26989 -33346
rect -25669 -34666 -25668 -33346
rect -26990 -34667 -25668 -34666
rect -25530 -33370 -25434 -33344
rect -24242 -33345 -24142 -33048
rect -25530 -34652 -25514 -33370
rect -25450 -34652 -25434 -33370
rect -26348 -34948 -26248 -34667
rect -25530 -34668 -25434 -34652
rect -24884 -33346 -23562 -33345
rect -24884 -34666 -24883 -33346
rect -23563 -34666 -23562 -33346
rect -24884 -34667 -23562 -34666
rect -23424 -33370 -23328 -33344
rect -22136 -33345 -22036 -33048
rect -23424 -34652 -23408 -33370
rect -23344 -34652 -23328 -33370
rect -24242 -34948 -24142 -34667
rect -23424 -34668 -23328 -34652
rect -22778 -33346 -21456 -33345
rect -22778 -34666 -22777 -33346
rect -21457 -34666 -21456 -33346
rect -22778 -34667 -21456 -34666
rect -21318 -33370 -21222 -33344
rect -20030 -33345 -19930 -33048
rect -21318 -34652 -21302 -33370
rect -21238 -34652 -21222 -33370
rect -22136 -34948 -22036 -34667
rect -21318 -34668 -21222 -34652
rect -20672 -33346 -19350 -33345
rect -20672 -34666 -20671 -33346
rect -19351 -34666 -19350 -33346
rect -20672 -34667 -19350 -34666
rect -19212 -33370 -19116 -33344
rect -17924 -33345 -17824 -33048
rect -19212 -34652 -19196 -33370
rect -19132 -34652 -19116 -33370
rect -20030 -34948 -19930 -34667
rect -19212 -34668 -19116 -34652
rect -18566 -33346 -17244 -33345
rect -18566 -34666 -18565 -33346
rect -17245 -34666 -17244 -33346
rect -18566 -34667 -17244 -34666
rect -17106 -33370 -17010 -33344
rect -15818 -33345 -15718 -33048
rect -17106 -34652 -17090 -33370
rect -17026 -34652 -17010 -33370
rect -17924 -34948 -17824 -34667
rect -17106 -34668 -17010 -34652
rect -16460 -33346 -15138 -33345
rect -16460 -34666 -16459 -33346
rect -15139 -34666 -15138 -33346
rect -16460 -34667 -15138 -34666
rect -15000 -33370 -14904 -33344
rect -13712 -33345 -13612 -33048
rect -15000 -34652 -14984 -33370
rect -14920 -34652 -14904 -33370
rect -15818 -34948 -15718 -34667
rect -15000 -34668 -14904 -34652
rect -14354 -33346 -13032 -33345
rect -14354 -34666 -14353 -33346
rect -13033 -34666 -13032 -33346
rect -14354 -34667 -13032 -34666
rect -12894 -33370 -12798 -33344
rect -11606 -33345 -11506 -33048
rect -12894 -34652 -12878 -33370
rect -12814 -34652 -12798 -33370
rect -13712 -34948 -13612 -34667
rect -12894 -34668 -12798 -34652
rect -12248 -33346 -10926 -33345
rect -12248 -34666 -12247 -33346
rect -10927 -34666 -10926 -33346
rect -12248 -34667 -10926 -34666
rect -10788 -33370 -10692 -33344
rect -9500 -33345 -9400 -33048
rect -10788 -34652 -10772 -33370
rect -10708 -34652 -10692 -33370
rect -11606 -34948 -11506 -34667
rect -10788 -34668 -10692 -34652
rect -10142 -33346 -8820 -33345
rect -10142 -34666 -10141 -33346
rect -8821 -34666 -8820 -33346
rect -10142 -34667 -8820 -34666
rect -8682 -33370 -8586 -33344
rect -7394 -33345 -7294 -33048
rect -8682 -34652 -8666 -33370
rect -8602 -34652 -8586 -33370
rect -9500 -34948 -9400 -34667
rect -8682 -34668 -8586 -34652
rect -8036 -33346 -6714 -33345
rect -8036 -34666 -8035 -33346
rect -6715 -34666 -6714 -33346
rect -8036 -34667 -6714 -34666
rect -6576 -33370 -6480 -33344
rect -5288 -33345 -5188 -33048
rect -6576 -34652 -6560 -33370
rect -6496 -34652 -6480 -33370
rect -7394 -34948 -7294 -34667
rect -6576 -34668 -6480 -34652
rect -5930 -33346 -4608 -33345
rect -5930 -34666 -5929 -33346
rect -4609 -34666 -4608 -33346
rect -5930 -34667 -4608 -34666
rect -4470 -33370 -4374 -33344
rect -3182 -33345 -3082 -33048
rect -4470 -34652 -4454 -33370
rect -4390 -34652 -4374 -33370
rect -5288 -34948 -5188 -34667
rect -4470 -34668 -4374 -34652
rect -3824 -33346 -2502 -33345
rect -3824 -34666 -3823 -33346
rect -2503 -34666 -2502 -33346
rect -3824 -34667 -2502 -34666
rect -2364 -33370 -2268 -33344
rect -1076 -33345 -976 -33048
rect -2364 -34652 -2348 -33370
rect -2284 -34652 -2268 -33370
rect -3182 -34948 -3082 -34667
rect -2364 -34668 -2268 -34652
rect -1718 -33346 -396 -33345
rect -1718 -34666 -1717 -33346
rect -397 -34666 -396 -33346
rect -1718 -34667 -396 -34666
rect -258 -33370 -162 -33344
rect 1030 -33345 1130 -33048
rect -258 -34652 -242 -33370
rect -178 -34652 -162 -33370
rect -1076 -34948 -976 -34667
rect -258 -34668 -162 -34652
rect 388 -33346 1710 -33345
rect 388 -34666 389 -33346
rect 1709 -34666 1710 -33346
rect 388 -34667 1710 -34666
rect 1848 -33370 1944 -33344
rect 3136 -33345 3236 -33048
rect 1848 -34652 1864 -33370
rect 1928 -34652 1944 -33370
rect 1030 -34948 1130 -34667
rect 1848 -34668 1944 -34652
rect 2494 -33346 3816 -33345
rect 2494 -34666 2495 -33346
rect 3815 -34666 3816 -33346
rect 2494 -34667 3816 -34666
rect 3954 -33370 4050 -33344
rect 5242 -33345 5342 -33048
rect 3954 -34652 3970 -33370
rect 4034 -34652 4050 -33370
rect 3136 -34948 3236 -34667
rect 3954 -34668 4050 -34652
rect 4600 -33346 5922 -33345
rect 4600 -34666 4601 -33346
rect 5921 -34666 5922 -33346
rect 4600 -34667 5922 -34666
rect 6060 -33370 6156 -33344
rect 7368 -33345 7468 -33048
rect 8160 -33344 8260 -33048
rect 6060 -34652 6076 -33370
rect 6140 -34652 6156 -33370
rect 5242 -34948 5342 -34667
rect 6060 -34668 6156 -34652
rect 6706 -33346 8028 -33345
rect 6706 -34666 6707 -33346
rect 8027 -33942 8028 -33346
rect 8160 -33370 8262 -33344
rect 8160 -33942 8182 -33370
rect 8027 -34042 8182 -33942
rect 8027 -34666 8028 -34042
rect 6706 -34667 8028 -34666
rect 8160 -34652 8182 -34042
rect 8246 -34652 8262 -33370
rect 7368 -34948 7468 -34667
rect 8160 -34668 8262 -34652
rect 8160 -34948 8260 -34668
rect -28470 -35048 8260 -34948
rect -28470 -35345 -28370 -35048
rect -29096 -35346 -27774 -35345
rect -29096 -36666 -29095 -35346
rect -27775 -35938 -27774 -35346
rect -27640 -35370 -27540 -35048
rect -26348 -35345 -26248 -35048
rect -27640 -35938 -27620 -35370
rect -27775 -36038 -27620 -35938
rect -27775 -36666 -27774 -36038
rect -29096 -36667 -27774 -36666
rect -27640 -36652 -27620 -36038
rect -27556 -36652 -27540 -35370
rect -28470 -36948 -28370 -36667
rect -27640 -36948 -27540 -36652
rect -26990 -35346 -25668 -35345
rect -26990 -36666 -26989 -35346
rect -25669 -36666 -25668 -35346
rect -26990 -36667 -25668 -36666
rect -25530 -35370 -25434 -35344
rect -24242 -35345 -24142 -35048
rect -25530 -36652 -25514 -35370
rect -25450 -36652 -25434 -35370
rect -26348 -36948 -26248 -36667
rect -25530 -36668 -25434 -36652
rect -24884 -35346 -23562 -35345
rect -24884 -36666 -24883 -35346
rect -23563 -36666 -23562 -35346
rect -24884 -36667 -23562 -36666
rect -23424 -35370 -23328 -35344
rect -22136 -35345 -22036 -35048
rect -23424 -36652 -23408 -35370
rect -23344 -36652 -23328 -35370
rect -24242 -36948 -24142 -36667
rect -23424 -36668 -23328 -36652
rect -22778 -35346 -21456 -35345
rect -22778 -36666 -22777 -35346
rect -21457 -36666 -21456 -35346
rect -22778 -36667 -21456 -36666
rect -21318 -35370 -21222 -35344
rect -20030 -35345 -19930 -35048
rect -21318 -36652 -21302 -35370
rect -21238 -36652 -21222 -35370
rect -22136 -36948 -22036 -36667
rect -21318 -36668 -21222 -36652
rect -20672 -35346 -19350 -35345
rect -20672 -36666 -20671 -35346
rect -19351 -36666 -19350 -35346
rect -20672 -36667 -19350 -36666
rect -19212 -35370 -19116 -35344
rect -17924 -35345 -17824 -35048
rect -19212 -36652 -19196 -35370
rect -19132 -36652 -19116 -35370
rect -20030 -36948 -19930 -36667
rect -19212 -36668 -19116 -36652
rect -18566 -35346 -17244 -35345
rect -18566 -36666 -18565 -35346
rect -17245 -36666 -17244 -35346
rect -18566 -36667 -17244 -36666
rect -17106 -35370 -17010 -35344
rect -15818 -35345 -15718 -35048
rect -17106 -36652 -17090 -35370
rect -17026 -36652 -17010 -35370
rect -17924 -36948 -17824 -36667
rect -17106 -36668 -17010 -36652
rect -16460 -35346 -15138 -35345
rect -16460 -36666 -16459 -35346
rect -15139 -36666 -15138 -35346
rect -16460 -36667 -15138 -36666
rect -15000 -35370 -14904 -35344
rect -13712 -35345 -13612 -35048
rect -15000 -36652 -14984 -35370
rect -14920 -36652 -14904 -35370
rect -15818 -36948 -15718 -36667
rect -15000 -36668 -14904 -36652
rect -14354 -35346 -13032 -35345
rect -14354 -36666 -14353 -35346
rect -13033 -36666 -13032 -35346
rect -14354 -36667 -13032 -36666
rect -12894 -35370 -12798 -35344
rect -11606 -35345 -11506 -35048
rect -12894 -36652 -12878 -35370
rect -12814 -36652 -12798 -35370
rect -13712 -36948 -13612 -36667
rect -12894 -36668 -12798 -36652
rect -12248 -35346 -10926 -35345
rect -12248 -36666 -12247 -35346
rect -10927 -36666 -10926 -35346
rect -12248 -36667 -10926 -36666
rect -10788 -35370 -10692 -35344
rect -9500 -35345 -9400 -35048
rect -10788 -36652 -10772 -35370
rect -10708 -36652 -10692 -35370
rect -11606 -36948 -11506 -36667
rect -10788 -36668 -10692 -36652
rect -10142 -35346 -8820 -35345
rect -10142 -36666 -10141 -35346
rect -8821 -36666 -8820 -35346
rect -10142 -36667 -8820 -36666
rect -8682 -35370 -8586 -35344
rect -7394 -35345 -7294 -35048
rect -8682 -36652 -8666 -35370
rect -8602 -36652 -8586 -35370
rect -9500 -36948 -9400 -36667
rect -8682 -36668 -8586 -36652
rect -8036 -35346 -6714 -35345
rect -8036 -36666 -8035 -35346
rect -6715 -36666 -6714 -35346
rect -8036 -36667 -6714 -36666
rect -6576 -35370 -6480 -35344
rect -5288 -35345 -5188 -35048
rect -6576 -36652 -6560 -35370
rect -6496 -36652 -6480 -35370
rect -7394 -36948 -7294 -36667
rect -6576 -36668 -6480 -36652
rect -5930 -35346 -4608 -35345
rect -5930 -36666 -5929 -35346
rect -4609 -36666 -4608 -35346
rect -5930 -36667 -4608 -36666
rect -4470 -35370 -4374 -35344
rect -3182 -35345 -3082 -35048
rect -4470 -36652 -4454 -35370
rect -4390 -36652 -4374 -35370
rect -5288 -36948 -5188 -36667
rect -4470 -36668 -4374 -36652
rect -3824 -35346 -2502 -35345
rect -3824 -36666 -3823 -35346
rect -2503 -36666 -2502 -35346
rect -3824 -36667 -2502 -36666
rect -2364 -35370 -2268 -35344
rect -1076 -35345 -976 -35048
rect -2364 -36652 -2348 -35370
rect -2284 -36652 -2268 -35370
rect -3182 -36948 -3082 -36667
rect -2364 -36668 -2268 -36652
rect -1718 -35346 -396 -35345
rect -1718 -36666 -1717 -35346
rect -397 -36666 -396 -35346
rect -1718 -36667 -396 -36666
rect -258 -35370 -162 -35344
rect 1030 -35345 1130 -35048
rect -258 -36652 -242 -35370
rect -178 -36652 -162 -35370
rect -1076 -36948 -976 -36667
rect -258 -36668 -162 -36652
rect 388 -35346 1710 -35345
rect 388 -36666 389 -35346
rect 1709 -36666 1710 -35346
rect 388 -36667 1710 -36666
rect 1848 -35370 1944 -35344
rect 3136 -35345 3236 -35048
rect 1848 -36652 1864 -35370
rect 1928 -36652 1944 -35370
rect 1030 -36948 1130 -36667
rect 1848 -36668 1944 -36652
rect 2494 -35346 3816 -35345
rect 2494 -36666 2495 -35346
rect 3815 -36666 3816 -35346
rect 2494 -36667 3816 -36666
rect 3954 -35370 4050 -35344
rect 5242 -35345 5342 -35048
rect 3954 -36652 3970 -35370
rect 4034 -36652 4050 -35370
rect 3136 -36948 3236 -36667
rect 3954 -36668 4050 -36652
rect 4600 -35346 5922 -35345
rect 4600 -36666 4601 -35346
rect 5921 -36666 5922 -35346
rect 4600 -36667 5922 -36666
rect 6060 -35370 6156 -35344
rect 7368 -35345 7468 -35048
rect 8160 -35344 8260 -35048
rect 6060 -36652 6076 -35370
rect 6140 -36652 6156 -35370
rect 5242 -36948 5342 -36667
rect 6060 -36668 6156 -36652
rect 6706 -35346 8028 -35345
rect 6706 -36666 6707 -35346
rect 8027 -35942 8028 -35346
rect 8160 -35370 8262 -35344
rect 8160 -35942 8182 -35370
rect 8027 -36042 8182 -35942
rect 8027 -36666 8028 -36042
rect 6706 -36667 8028 -36666
rect 8160 -36652 8182 -36042
rect 8246 -36652 8262 -35370
rect 7368 -36948 7468 -36667
rect 8160 -36668 8262 -36652
rect 10276 -35824 10826 -30124
rect 11126 -35824 11458 -30124
rect 24016 -30124 25316 -30068
rect 10276 -36616 11458 -35824
rect 8160 -36948 8260 -36668
rect -28470 -37048 8260 -36948
rect -28470 -37345 -28370 -37048
rect -29096 -37346 -27774 -37345
rect -29096 -38666 -29095 -37346
rect -27775 -37938 -27774 -37346
rect -27640 -37370 -27540 -37048
rect -26348 -37345 -26248 -37048
rect -27640 -37938 -27620 -37370
rect -27775 -38038 -27620 -37938
rect -27775 -38666 -27774 -38038
rect -29096 -38667 -27774 -38666
rect -27640 -38652 -27620 -38038
rect -27556 -38652 -27540 -37370
rect -28470 -38948 -28370 -38667
rect -27640 -38948 -27540 -38652
rect -26990 -37346 -25668 -37345
rect -26990 -38666 -26989 -37346
rect -25669 -38666 -25668 -37346
rect -26990 -38667 -25668 -38666
rect -25530 -37370 -25434 -37344
rect -24242 -37345 -24142 -37048
rect -25530 -38652 -25514 -37370
rect -25450 -38652 -25434 -37370
rect -26348 -38948 -26248 -38667
rect -25530 -38668 -25434 -38652
rect -24884 -37346 -23562 -37345
rect -24884 -38666 -24883 -37346
rect -23563 -38666 -23562 -37346
rect -24884 -38667 -23562 -38666
rect -23424 -37370 -23328 -37344
rect -22136 -37345 -22036 -37048
rect -23424 -38652 -23408 -37370
rect -23344 -38652 -23328 -37370
rect -24242 -38948 -24142 -38667
rect -23424 -38668 -23328 -38652
rect -22778 -37346 -21456 -37345
rect -22778 -38666 -22777 -37346
rect -21457 -38666 -21456 -37346
rect -22778 -38667 -21456 -38666
rect -21318 -37370 -21222 -37344
rect -20030 -37345 -19930 -37048
rect -21318 -38652 -21302 -37370
rect -21238 -38652 -21222 -37370
rect -22136 -38948 -22036 -38667
rect -21318 -38668 -21222 -38652
rect -20672 -37346 -19350 -37345
rect -20672 -38666 -20671 -37346
rect -19351 -38666 -19350 -37346
rect -20672 -38667 -19350 -38666
rect -19212 -37370 -19116 -37344
rect -17924 -37345 -17824 -37048
rect -19212 -38652 -19196 -37370
rect -19132 -38652 -19116 -37370
rect -20030 -38948 -19930 -38667
rect -19212 -38668 -19116 -38652
rect -18566 -37346 -17244 -37345
rect -18566 -38666 -18565 -37346
rect -17245 -38666 -17244 -37346
rect -18566 -38667 -17244 -38666
rect -17106 -37370 -17010 -37344
rect -15818 -37345 -15718 -37048
rect -17106 -38652 -17090 -37370
rect -17026 -38652 -17010 -37370
rect -17924 -38948 -17824 -38667
rect -17106 -38668 -17010 -38652
rect -16460 -37346 -15138 -37345
rect -16460 -38666 -16459 -37346
rect -15139 -38666 -15138 -37346
rect -16460 -38667 -15138 -38666
rect -15000 -37370 -14904 -37344
rect -13712 -37345 -13612 -37048
rect -15000 -38652 -14984 -37370
rect -14920 -38652 -14904 -37370
rect -15818 -38948 -15718 -38667
rect -15000 -38668 -14904 -38652
rect -14354 -37346 -13032 -37345
rect -14354 -38666 -14353 -37346
rect -13033 -38666 -13032 -37346
rect -14354 -38667 -13032 -38666
rect -12894 -37370 -12798 -37344
rect -11606 -37345 -11506 -37048
rect -12894 -38652 -12878 -37370
rect -12814 -38652 -12798 -37370
rect -13712 -38948 -13612 -38667
rect -12894 -38668 -12798 -38652
rect -12248 -37346 -10926 -37345
rect -12248 -38666 -12247 -37346
rect -10927 -38666 -10926 -37346
rect -12248 -38667 -10926 -38666
rect -10788 -37370 -10692 -37344
rect -9500 -37345 -9400 -37048
rect -10788 -38652 -10772 -37370
rect -10708 -38652 -10692 -37370
rect -11606 -38948 -11506 -38667
rect -10788 -38668 -10692 -38652
rect -10142 -37346 -8820 -37345
rect -10142 -38666 -10141 -37346
rect -8821 -38666 -8820 -37346
rect -10142 -38667 -8820 -38666
rect -8682 -37370 -8586 -37344
rect -7394 -37345 -7294 -37048
rect -8682 -38652 -8666 -37370
rect -8602 -38652 -8586 -37370
rect -9500 -38948 -9400 -38667
rect -8682 -38668 -8586 -38652
rect -8036 -37346 -6714 -37345
rect -8036 -38666 -8035 -37346
rect -6715 -38666 -6714 -37346
rect -8036 -38667 -6714 -38666
rect -6576 -37370 -6480 -37344
rect -5288 -37345 -5188 -37048
rect -6576 -38652 -6560 -37370
rect -6496 -38652 -6480 -37370
rect -7394 -38948 -7294 -38667
rect -6576 -38668 -6480 -38652
rect -5930 -37346 -4608 -37345
rect -5930 -38666 -5929 -37346
rect -4609 -38666 -4608 -37346
rect -5930 -38667 -4608 -38666
rect -4470 -37370 -4374 -37344
rect -3182 -37345 -3082 -37048
rect -4470 -38652 -4454 -37370
rect -4390 -38652 -4374 -37370
rect -5288 -38948 -5188 -38667
rect -4470 -38668 -4374 -38652
rect -3824 -37346 -2502 -37345
rect -3824 -38666 -3823 -37346
rect -2503 -38666 -2502 -37346
rect -3824 -38667 -2502 -38666
rect -2364 -37370 -2268 -37344
rect -1076 -37345 -976 -37048
rect -2364 -38652 -2348 -37370
rect -2284 -38652 -2268 -37370
rect -3182 -38948 -3082 -38667
rect -2364 -38668 -2268 -38652
rect -1718 -37346 -396 -37345
rect -1718 -38666 -1717 -37346
rect -397 -38666 -396 -37346
rect -1718 -38667 -396 -38666
rect -258 -37370 -162 -37344
rect 1030 -37345 1130 -37048
rect -258 -38652 -242 -37370
rect -178 -38652 -162 -37370
rect -1076 -38948 -976 -38667
rect -258 -38668 -162 -38652
rect 388 -37346 1710 -37345
rect 388 -38666 389 -37346
rect 1709 -38666 1710 -37346
rect 388 -38667 1710 -38666
rect 1848 -37370 1944 -37344
rect 3136 -37345 3236 -37048
rect 1848 -38652 1864 -37370
rect 1928 -38652 1944 -37370
rect 1030 -38948 1130 -38667
rect 1848 -38668 1944 -38652
rect 2494 -37346 3816 -37345
rect 2494 -38666 2495 -37346
rect 3815 -38666 3816 -37346
rect 2494 -38667 3816 -38666
rect 3954 -37370 4050 -37344
rect 5242 -37345 5342 -37048
rect 3954 -38652 3970 -37370
rect 4034 -38652 4050 -37370
rect 3136 -38948 3236 -38667
rect 3954 -38668 4050 -38652
rect 4600 -37346 5922 -37345
rect 4600 -38666 4601 -37346
rect 5921 -38666 5922 -37346
rect 4600 -38667 5922 -38666
rect 6060 -37370 6156 -37344
rect 7368 -37345 7468 -37048
rect 8160 -37344 8260 -37048
rect 6060 -38652 6076 -37370
rect 6140 -38652 6156 -37370
rect 5242 -38948 5342 -38667
rect 6060 -38668 6156 -38652
rect 6706 -37346 8028 -37345
rect 6706 -38666 6707 -37346
rect 8027 -37942 8028 -37346
rect 8160 -37370 8262 -37344
rect 8160 -37942 8182 -37370
rect 8027 -38042 8182 -37942
rect 8027 -38666 8028 -38042
rect 6706 -38667 8028 -38666
rect 8160 -38652 8182 -38042
rect 8246 -38652 8262 -37370
rect 7368 -38948 7468 -38667
rect 8160 -38668 8262 -38652
rect 8160 -38948 8260 -38668
rect -28470 -39048 8260 -38948
rect -28470 -39345 -28370 -39048
rect -29096 -39346 -27774 -39345
rect -29096 -40666 -29095 -39346
rect -27775 -39938 -27774 -39346
rect -27640 -39370 -27540 -39048
rect -26348 -39345 -26248 -39048
rect -27640 -39938 -27620 -39370
rect -27775 -40038 -27620 -39938
rect -27775 -40666 -27774 -40038
rect -29096 -40667 -27774 -40666
rect -27640 -40652 -27620 -40038
rect -27556 -40652 -27540 -39370
rect -28470 -40948 -28370 -40667
rect -27640 -40948 -27540 -40652
rect -26990 -39346 -25668 -39345
rect -26990 -40666 -26989 -39346
rect -25669 -40666 -25668 -39346
rect -26990 -40667 -25668 -40666
rect -25530 -39370 -25434 -39344
rect -24242 -39345 -24142 -39048
rect -25530 -40652 -25514 -39370
rect -25450 -40652 -25434 -39370
rect -26348 -40948 -26248 -40667
rect -25530 -40668 -25434 -40652
rect -24884 -39346 -23562 -39345
rect -24884 -40666 -24883 -39346
rect -23563 -40666 -23562 -39346
rect -24884 -40667 -23562 -40666
rect -23424 -39370 -23328 -39344
rect -22136 -39345 -22036 -39048
rect -23424 -40652 -23408 -39370
rect -23344 -40652 -23328 -39370
rect -24242 -40948 -24142 -40667
rect -23424 -40668 -23328 -40652
rect -22778 -39346 -21456 -39345
rect -22778 -40666 -22777 -39346
rect -21457 -40666 -21456 -39346
rect -22778 -40667 -21456 -40666
rect -21318 -39370 -21222 -39344
rect -20030 -39345 -19930 -39048
rect -21318 -40652 -21302 -39370
rect -21238 -40652 -21222 -39370
rect -22136 -40948 -22036 -40667
rect -21318 -40668 -21222 -40652
rect -20672 -39346 -19350 -39345
rect -20672 -40666 -20671 -39346
rect -19351 -40666 -19350 -39346
rect -20672 -40667 -19350 -40666
rect -19212 -39370 -19116 -39344
rect -17924 -39345 -17824 -39048
rect -19212 -40652 -19196 -39370
rect -19132 -40652 -19116 -39370
rect -20030 -40948 -19930 -40667
rect -19212 -40668 -19116 -40652
rect -18566 -39346 -17244 -39345
rect -18566 -40666 -18565 -39346
rect -17245 -40666 -17244 -39346
rect -18566 -40667 -17244 -40666
rect -17106 -39370 -17010 -39344
rect -15818 -39345 -15718 -39048
rect -17106 -40652 -17090 -39370
rect -17026 -40652 -17010 -39370
rect -17924 -40948 -17824 -40667
rect -17106 -40668 -17010 -40652
rect -16460 -39346 -15138 -39345
rect -16460 -40666 -16459 -39346
rect -15139 -40666 -15138 -39346
rect -16460 -40667 -15138 -40666
rect -15000 -39370 -14904 -39344
rect -13712 -39345 -13612 -39048
rect -15000 -40652 -14984 -39370
rect -14920 -40652 -14904 -39370
rect -15818 -40948 -15718 -40667
rect -15000 -40668 -14904 -40652
rect -14354 -39346 -13032 -39345
rect -14354 -40666 -14353 -39346
rect -13033 -40666 -13032 -39346
rect -14354 -40667 -13032 -40666
rect -12894 -39370 -12798 -39344
rect -11606 -39345 -11506 -39048
rect -12894 -40652 -12878 -39370
rect -12814 -40652 -12798 -39370
rect -13712 -40948 -13612 -40667
rect -12894 -40668 -12798 -40652
rect -12248 -39346 -10926 -39345
rect -12248 -40666 -12247 -39346
rect -10927 -40666 -10926 -39346
rect -12248 -40667 -10926 -40666
rect -10788 -39370 -10692 -39344
rect -9500 -39345 -9400 -39048
rect -10788 -40652 -10772 -39370
rect -10708 -40652 -10692 -39370
rect -11606 -40948 -11506 -40667
rect -10788 -40668 -10692 -40652
rect -10142 -39346 -8820 -39345
rect -10142 -40666 -10141 -39346
rect -8821 -40666 -8820 -39346
rect -10142 -40667 -8820 -40666
rect -8682 -39370 -8586 -39344
rect -7394 -39345 -7294 -39048
rect -8682 -40652 -8666 -39370
rect -8602 -40652 -8586 -39370
rect -9500 -40948 -9400 -40667
rect -8682 -40668 -8586 -40652
rect -8036 -39346 -6714 -39345
rect -8036 -40666 -8035 -39346
rect -6715 -40666 -6714 -39346
rect -8036 -40667 -6714 -40666
rect -6576 -39370 -6480 -39344
rect -5288 -39345 -5188 -39048
rect -6576 -40652 -6560 -39370
rect -6496 -40652 -6480 -39370
rect -7394 -40948 -7294 -40667
rect -6576 -40668 -6480 -40652
rect -5930 -39346 -4608 -39345
rect -5930 -40666 -5929 -39346
rect -4609 -40666 -4608 -39346
rect -5930 -40667 -4608 -40666
rect -4470 -39370 -4374 -39344
rect -3182 -39345 -3082 -39048
rect -4470 -40652 -4454 -39370
rect -4390 -40652 -4374 -39370
rect -5288 -40948 -5188 -40667
rect -4470 -40668 -4374 -40652
rect -3824 -39346 -2502 -39345
rect -3824 -40666 -3823 -39346
rect -2503 -40666 -2502 -39346
rect -3824 -40667 -2502 -40666
rect -2364 -39370 -2268 -39344
rect -1076 -39345 -976 -39048
rect -2364 -40652 -2348 -39370
rect -2284 -40652 -2268 -39370
rect -3182 -40948 -3082 -40667
rect -2364 -40668 -2268 -40652
rect -1718 -39346 -396 -39345
rect -1718 -40666 -1717 -39346
rect -397 -40666 -396 -39346
rect -1718 -40667 -396 -40666
rect -258 -39370 -162 -39344
rect 1030 -39345 1130 -39048
rect -258 -40652 -242 -39370
rect -178 -40652 -162 -39370
rect -1076 -40948 -976 -40667
rect -258 -40668 -162 -40652
rect 388 -39346 1710 -39345
rect 388 -40666 389 -39346
rect 1709 -40666 1710 -39346
rect 388 -40667 1710 -40666
rect 1848 -39370 1944 -39344
rect 3136 -39345 3236 -39048
rect 1848 -40652 1864 -39370
rect 1928 -40652 1944 -39370
rect 1030 -40948 1130 -40667
rect 1848 -40668 1944 -40652
rect 2494 -39346 3816 -39345
rect 2494 -40666 2495 -39346
rect 3815 -40666 3816 -39346
rect 2494 -40667 3816 -40666
rect 3954 -39370 4050 -39344
rect 5242 -39345 5342 -39048
rect 3954 -40652 3970 -39370
rect 4034 -40652 4050 -39370
rect 3136 -40948 3236 -40667
rect 3954 -40668 4050 -40652
rect 4600 -39346 5922 -39345
rect 4600 -40666 4601 -39346
rect 5921 -40666 5922 -39346
rect 4600 -40667 5922 -40666
rect 6060 -39370 6156 -39344
rect 7368 -39345 7468 -39048
rect 8160 -39344 8260 -39048
rect 6060 -40652 6076 -39370
rect 6140 -40652 6156 -39370
rect 5242 -40948 5342 -40667
rect 6060 -40668 6156 -40652
rect 6706 -39346 8028 -39345
rect 6706 -40666 6707 -39346
rect 8027 -39942 8028 -39346
rect 8160 -39370 8262 -39344
rect 8160 -39942 8182 -39370
rect 8027 -40042 8182 -39942
rect 8027 -40666 8028 -40042
rect 6706 -40667 8028 -40666
rect 8160 -40652 8182 -40042
rect 8246 -40652 8262 -39370
rect 7368 -40948 7468 -40667
rect 8160 -40668 8262 -40652
rect 8160 -40948 8260 -40668
rect -28470 -41048 8260 -40948
rect -28470 -41345 -28370 -41048
rect -29096 -41346 -27774 -41345
rect -29096 -42666 -29095 -41346
rect -27775 -41938 -27774 -41346
rect -27640 -41370 -27540 -41048
rect -26348 -41345 -26248 -41048
rect -27640 -41938 -27620 -41370
rect -27775 -42038 -27620 -41938
rect -27775 -42666 -27774 -42038
rect -29096 -42667 -27774 -42666
rect -27640 -42652 -27620 -42038
rect -27556 -42652 -27540 -41370
rect -28470 -42948 -28370 -42667
rect -27640 -42948 -27540 -42652
rect -26990 -41346 -25668 -41345
rect -26990 -42666 -26989 -41346
rect -25669 -42666 -25668 -41346
rect -26990 -42667 -25668 -42666
rect -25530 -41370 -25434 -41344
rect -24242 -41345 -24142 -41048
rect -25530 -42652 -25514 -41370
rect -25450 -42652 -25434 -41370
rect -26348 -42948 -26248 -42667
rect -25530 -42668 -25434 -42652
rect -24884 -41346 -23562 -41345
rect -24884 -42666 -24883 -41346
rect -23563 -42666 -23562 -41346
rect -24884 -42667 -23562 -42666
rect -23424 -41370 -23328 -41344
rect -22136 -41345 -22036 -41048
rect -23424 -42652 -23408 -41370
rect -23344 -42652 -23328 -41370
rect -24242 -42948 -24142 -42667
rect -23424 -42668 -23328 -42652
rect -22778 -41346 -21456 -41345
rect -22778 -42666 -22777 -41346
rect -21457 -42666 -21456 -41346
rect -22778 -42667 -21456 -42666
rect -21318 -41370 -21222 -41344
rect -20030 -41345 -19930 -41048
rect -21318 -42652 -21302 -41370
rect -21238 -42652 -21222 -41370
rect -22136 -42948 -22036 -42667
rect -21318 -42668 -21222 -42652
rect -20672 -41346 -19350 -41345
rect -20672 -42666 -20671 -41346
rect -19351 -42666 -19350 -41346
rect -20672 -42667 -19350 -42666
rect -19212 -41370 -19116 -41344
rect -17924 -41345 -17824 -41048
rect -19212 -42652 -19196 -41370
rect -19132 -42652 -19116 -41370
rect -20030 -42948 -19930 -42667
rect -19212 -42668 -19116 -42652
rect -18566 -41346 -17244 -41345
rect -18566 -42666 -18565 -41346
rect -17245 -42666 -17244 -41346
rect -18566 -42667 -17244 -42666
rect -17106 -41370 -17010 -41344
rect -15818 -41345 -15718 -41048
rect -17106 -42652 -17090 -41370
rect -17026 -42652 -17010 -41370
rect -17924 -42948 -17824 -42667
rect -17106 -42668 -17010 -42652
rect -16460 -41346 -15138 -41345
rect -16460 -42666 -16459 -41346
rect -15139 -42666 -15138 -41346
rect -16460 -42667 -15138 -42666
rect -15000 -41370 -14904 -41344
rect -13712 -41345 -13612 -41048
rect -15000 -42652 -14984 -41370
rect -14920 -42652 -14904 -41370
rect -15818 -42948 -15718 -42667
rect -15000 -42668 -14904 -42652
rect -14354 -41346 -13032 -41345
rect -14354 -42666 -14353 -41346
rect -13033 -42666 -13032 -41346
rect -14354 -42667 -13032 -42666
rect -12894 -41370 -12798 -41344
rect -11606 -41345 -11506 -41048
rect -12894 -42652 -12878 -41370
rect -12814 -42652 -12798 -41370
rect -13712 -42948 -13612 -42667
rect -12894 -42668 -12798 -42652
rect -12248 -41346 -10926 -41345
rect -12248 -42666 -12247 -41346
rect -10927 -42666 -10926 -41346
rect -12248 -42667 -10926 -42666
rect -10788 -41370 -10692 -41344
rect -9500 -41345 -9400 -41048
rect -10788 -42652 -10772 -41370
rect -10708 -42652 -10692 -41370
rect -11606 -42948 -11506 -42667
rect -10788 -42668 -10692 -42652
rect -10142 -41346 -8820 -41345
rect -10142 -42666 -10141 -41346
rect -8821 -42666 -8820 -41346
rect -10142 -42667 -8820 -42666
rect -8682 -41370 -8586 -41344
rect -7394 -41345 -7294 -41048
rect -8682 -42652 -8666 -41370
rect -8602 -42652 -8586 -41370
rect -9500 -42948 -9400 -42667
rect -8682 -42668 -8586 -42652
rect -8036 -41346 -6714 -41345
rect -8036 -42666 -8035 -41346
rect -6715 -42666 -6714 -41346
rect -8036 -42667 -6714 -42666
rect -6576 -41370 -6480 -41344
rect -5288 -41345 -5188 -41048
rect -6576 -42652 -6560 -41370
rect -6496 -42652 -6480 -41370
rect -7394 -42948 -7294 -42667
rect -6576 -42668 -6480 -42652
rect -5930 -41346 -4608 -41345
rect -5930 -42666 -5929 -41346
rect -4609 -42666 -4608 -41346
rect -5930 -42667 -4608 -42666
rect -4470 -41370 -4374 -41344
rect -3182 -41345 -3082 -41048
rect -4470 -42652 -4454 -41370
rect -4390 -42652 -4374 -41370
rect -5288 -42948 -5188 -42667
rect -4470 -42668 -4374 -42652
rect -3824 -41346 -2502 -41345
rect -3824 -42666 -3823 -41346
rect -2503 -42666 -2502 -41346
rect -3824 -42667 -2502 -42666
rect -2364 -41370 -2268 -41344
rect -1076 -41345 -976 -41048
rect -2364 -42652 -2348 -41370
rect -2284 -42652 -2268 -41370
rect -3182 -42948 -3082 -42667
rect -2364 -42668 -2268 -42652
rect -1718 -41346 -396 -41345
rect -1718 -42666 -1717 -41346
rect -397 -42666 -396 -41346
rect -1718 -42667 -396 -42666
rect -258 -41370 -162 -41344
rect 1030 -41345 1130 -41048
rect -258 -42652 -242 -41370
rect -178 -42652 -162 -41370
rect -1076 -42948 -976 -42667
rect -258 -42668 -162 -42652
rect 388 -41346 1710 -41345
rect 388 -42666 389 -41346
rect 1709 -42666 1710 -41346
rect 388 -42667 1710 -42666
rect 1848 -41370 1944 -41344
rect 3136 -41345 3236 -41048
rect 1848 -42652 1864 -41370
rect 1928 -42652 1944 -41370
rect 1030 -42948 1130 -42667
rect 1848 -42668 1944 -42652
rect 2494 -41346 3816 -41345
rect 2494 -42666 2495 -41346
rect 3815 -42666 3816 -41346
rect 2494 -42667 3816 -42666
rect 3954 -41370 4050 -41344
rect 5242 -41345 5342 -41048
rect 3954 -42652 3970 -41370
rect 4034 -42652 4050 -41370
rect 3136 -42948 3236 -42667
rect 3954 -42668 4050 -42652
rect 4600 -41346 5922 -41345
rect 4600 -42666 4601 -41346
rect 5921 -42666 5922 -41346
rect 4600 -42667 5922 -42666
rect 6060 -41370 6156 -41344
rect 7368 -41345 7468 -41048
rect 8160 -41344 8260 -41048
rect 6060 -42652 6076 -41370
rect 6140 -42652 6156 -41370
rect 5242 -42948 5342 -42667
rect 6060 -42668 6156 -42652
rect 6706 -41346 8028 -41345
rect 6706 -42666 6707 -41346
rect 8027 -41942 8028 -41346
rect 8160 -41370 8262 -41344
rect 8160 -41942 8182 -41370
rect 8027 -42042 8182 -41942
rect 8027 -42666 8028 -42042
rect 6706 -42667 8028 -42666
rect 8160 -42652 8182 -42042
rect 8246 -42652 8262 -41370
rect 7368 -42948 7468 -42667
rect 8160 -42668 8262 -42652
rect 10276 -42316 10826 -36616
rect 11126 -42316 11458 -36616
rect 12216 -31042 23216 -30892
rect 12216 -35742 17166 -31042
rect 17466 -35742 22766 -31042
rect 23066 -35742 23216 -31042
rect 12216 -36642 23216 -35742
rect 12216 -41342 17166 -36642
rect 17466 -41342 22766 -36642
rect 23066 -41342 23216 -36642
rect 12216 -41794 23216 -41342
rect 24016 -35824 24870 -30124
rect 25170 -35824 25316 -30124
rect 24016 -36616 25316 -35824
rect 24016 -41414 24870 -36616
rect 12216 -41891 24117 -41794
rect 12216 -41892 23216 -41891
rect 8160 -42948 8260 -42668
rect 10276 -42730 11458 -42316
rect 10276 -42816 22722 -42730
rect -28470 -43048 8260 -42948
rect -28470 -43345 -28370 -43048
rect -29096 -43346 -27774 -43345
rect -29096 -44666 -29095 -43346
rect -27775 -43938 -27774 -43346
rect -27640 -43370 -27540 -43048
rect -26348 -43345 -26248 -43048
rect -27640 -43938 -27620 -43370
rect -27775 -44038 -27620 -43938
rect -27775 -44666 -27774 -44038
rect -29096 -44667 -27774 -44666
rect -27640 -44652 -27620 -44038
rect -27556 -44652 -27540 -43370
rect -28470 -44942 -28370 -44667
rect -27640 -44942 -27540 -44652
rect -26990 -43346 -25668 -43345
rect -26990 -44666 -26989 -43346
rect -25669 -44666 -25668 -43346
rect -26990 -44667 -25668 -44666
rect -25530 -43370 -25434 -43344
rect -24242 -43345 -24142 -43048
rect -25530 -44652 -25514 -43370
rect -25450 -44652 -25434 -43370
rect -26348 -44942 -26248 -44667
rect -25530 -44668 -25434 -44652
rect -24884 -43346 -23562 -43345
rect -24884 -44666 -24883 -43346
rect -23563 -44666 -23562 -43346
rect -24884 -44667 -23562 -44666
rect -23424 -43370 -23328 -43344
rect -22136 -43345 -22036 -43048
rect -23424 -44652 -23408 -43370
rect -23344 -44652 -23328 -43370
rect -24242 -44942 -24142 -44667
rect -23424 -44668 -23328 -44652
rect -22778 -43346 -21456 -43345
rect -22778 -44666 -22777 -43346
rect -21457 -44666 -21456 -43346
rect -22778 -44667 -21456 -44666
rect -21318 -43370 -21222 -43344
rect -20030 -43345 -19930 -43048
rect -21318 -44652 -21302 -43370
rect -21238 -44652 -21222 -43370
rect -22136 -44942 -22036 -44667
rect -21318 -44668 -21222 -44652
rect -20672 -43346 -19350 -43345
rect -20672 -44666 -20671 -43346
rect -19351 -44666 -19350 -43346
rect -20672 -44667 -19350 -44666
rect -19212 -43370 -19116 -43344
rect -17924 -43345 -17824 -43048
rect -19212 -44652 -19196 -43370
rect -19132 -44652 -19116 -43370
rect -20030 -44942 -19930 -44667
rect -19212 -44668 -19116 -44652
rect -18566 -43346 -17244 -43345
rect -18566 -44666 -18565 -43346
rect -17245 -44666 -17244 -43346
rect -18566 -44667 -17244 -44666
rect -17106 -43370 -17010 -43344
rect -15818 -43345 -15718 -43048
rect -17106 -44652 -17090 -43370
rect -17026 -44652 -17010 -43370
rect -17924 -44942 -17824 -44667
rect -17106 -44668 -17010 -44652
rect -16460 -43346 -15138 -43345
rect -16460 -44666 -16459 -43346
rect -15139 -44666 -15138 -43346
rect -16460 -44667 -15138 -44666
rect -15000 -43370 -14904 -43344
rect -15000 -44652 -14984 -43370
rect -14920 -44652 -14904 -43370
rect -15818 -44942 -15718 -44667
rect -15000 -44668 -14904 -44652
rect -14354 -43346 -13032 -43345
rect -14354 -44666 -14353 -43346
rect -13033 -44666 -13032 -43346
rect -14354 -44667 -13032 -44666
rect -12894 -43370 -12798 -43344
rect -11606 -43345 -11506 -43048
rect -12894 -44652 -12878 -43370
rect -12814 -44652 -12798 -43370
rect -13712 -44942 -13612 -44667
rect -12894 -44668 -12798 -44652
rect -12248 -43346 -10926 -43345
rect -12248 -44666 -12247 -43346
rect -10927 -44666 -10926 -43346
rect -12248 -44667 -10926 -44666
rect -10788 -43370 -10692 -43344
rect -9500 -43345 -9400 -43048
rect -10788 -44652 -10772 -43370
rect -10708 -44652 -10692 -43370
rect -11606 -44942 -11506 -44667
rect -10788 -44668 -10692 -44652
rect -10142 -43346 -8820 -43345
rect -10142 -44666 -10141 -43346
rect -8821 -44666 -8820 -43346
rect -8682 -43370 -8586 -43344
rect -8682 -44560 -8666 -43370
rect -10142 -44667 -8820 -44666
rect -8684 -44652 -8666 -44560
rect -8602 -44560 -8586 -43370
rect -8036 -43346 -6714 -43345
rect -8602 -44652 -8584 -44560
rect -9500 -44942 -9400 -44667
rect -28470 -45042 -9400 -44942
rect -8684 -44864 -8584 -44652
rect -8036 -44666 -8035 -43346
rect -6715 -44666 -6714 -43346
rect -8036 -44667 -6714 -44666
rect -6576 -43370 -6480 -43344
rect -5288 -43345 -5188 -43048
rect -6576 -44652 -6560 -43370
rect -6496 -44652 -6480 -43370
rect -8684 -44964 -8182 -44864
rect -7394 -44948 -7294 -44667
rect -6576 -44668 -6480 -44652
rect -5930 -43346 -4608 -43345
rect -5930 -44666 -5929 -43346
rect -4609 -44666 -4608 -43346
rect -5930 -44667 -4608 -44666
rect -4470 -43370 -4374 -43344
rect -3182 -43345 -3082 -43048
rect -4470 -44652 -4454 -43370
rect -4390 -44652 -4374 -43370
rect -5288 -44948 -5188 -44667
rect -4470 -44668 -4374 -44652
rect -3824 -43346 -2502 -43345
rect -3824 -44666 -3823 -43346
rect -2503 -44666 -2502 -43346
rect -3824 -44667 -2502 -44666
rect -2364 -43370 -2268 -43344
rect -1076 -43345 -976 -43048
rect -2364 -44652 -2348 -43370
rect -2284 -44652 -2268 -43370
rect -3182 -44948 -3082 -44667
rect -2364 -44668 -2268 -44652
rect -1718 -43346 -396 -43345
rect -1718 -44666 -1717 -43346
rect -397 -44666 -396 -43346
rect -1718 -44667 -396 -44666
rect -258 -43370 -162 -43344
rect 1030 -43345 1130 -43048
rect -258 -44652 -242 -43370
rect -178 -44652 -162 -43370
rect -1076 -44948 -976 -44667
rect -258 -44668 -162 -44652
rect 388 -43346 1710 -43345
rect 388 -44666 389 -43346
rect 1709 -44666 1710 -43346
rect 388 -44667 1710 -44666
rect 1848 -43370 1944 -43344
rect 3136 -43345 3236 -43048
rect 1848 -44652 1864 -43370
rect 1928 -44652 1944 -43370
rect 1030 -44948 1130 -44667
rect 1848 -44668 1944 -44652
rect 2494 -43346 3816 -43345
rect 2494 -44666 2495 -43346
rect 3815 -44666 3816 -43346
rect 2494 -44667 3816 -44666
rect 3954 -43370 4050 -43344
rect 5242 -43345 5342 -43048
rect 3954 -44652 3970 -43370
rect 4034 -44652 4050 -43370
rect 3136 -44948 3236 -44667
rect 3954 -44668 4050 -44652
rect 4600 -43346 5922 -43345
rect 4600 -44666 4601 -43346
rect 5921 -44666 5922 -43346
rect 4600 -44667 5922 -44666
rect 6060 -43370 6156 -43344
rect 7368 -43345 7468 -43048
rect 8160 -43344 8260 -43048
rect 10278 -42956 22722 -42816
rect 10278 -43042 23722 -42956
rect 10278 -43342 16812 -43042
rect 17112 -43342 23212 -43042
rect 23512 -43342 23722 -43042
rect 6060 -44652 6076 -43370
rect 6140 -44652 6156 -43370
rect 5242 -44948 5342 -44667
rect 6060 -44668 6156 -44652
rect 6706 -43346 8028 -43345
rect 6706 -44666 6707 -43346
rect 8027 -43942 8028 -43346
rect 8160 -43370 8262 -43344
rect 8160 -43942 8182 -43370
rect 8027 -44042 8182 -43942
rect 8027 -44666 8028 -44042
rect 6706 -44667 8028 -44666
rect 8160 -44652 8182 -44042
rect 8246 -44652 8262 -43370
rect 10278 -43894 23722 -43342
rect 24020 -43378 24117 -41891
rect 24386 -42316 24870 -41414
rect 25170 -42316 25316 -36616
rect 50552 -38692 52664 -38680
rect 50552 -38704 58368 -38692
rect 50552 -39456 50576 -38704
rect 51328 -39086 58368 -38704
rect 51328 -39386 52262 -39086
rect 55130 -39386 56534 -39086
rect 58154 -39386 58368 -39086
rect 51328 -39456 58368 -39386
rect 50552 -39480 58368 -39456
rect 52078 -39492 58368 -39480
rect 57454 -40471 58522 -40454
rect 57454 -40541 57475 -40471
rect 57539 -40541 58522 -40471
rect 57454 -40554 58522 -40541
rect 58422 -42207 58522 -40554
rect 58422 -42208 58525 -42207
rect 58422 -42214 58424 -42208
rect 24386 -42826 25316 -42316
rect 57946 -42308 58424 -42214
rect 58524 -42308 58525 -42208
rect 57946 -42309 58525 -42308
rect 57946 -42314 58522 -42309
rect 53295 -42460 53397 -42459
rect 53295 -42462 53296 -42460
rect 53288 -42560 53296 -42462
rect 53396 -42462 53397 -42460
rect 53396 -42466 56146 -42462
rect 53396 -42471 55300 -42466
rect 53396 -42553 54195 -42471
rect 54259 -42553 55300 -42471
rect 53396 -42558 55300 -42553
rect 55370 -42558 56146 -42466
rect 53396 -42560 56146 -42558
rect 53288 -42562 56146 -42560
rect 56042 -42573 56146 -42562
rect 56042 -42671 56043 -42573
rect 56141 -42671 56146 -42573
rect 56042 -42672 56146 -42671
rect 56046 -42676 56146 -42672
rect 57946 -42575 58046 -42314
rect 57946 -42673 57947 -42575
rect 58045 -42673 58046 -42575
rect 57946 -42674 58046 -42673
rect 25670 -42923 27858 -42922
rect 25670 -42937 27759 -42923
rect 25670 -43001 26981 -42937
rect 27051 -43001 27759 -42937
rect 25670 -43021 27759 -43001
rect 27857 -43021 27858 -42923
rect 25670 -43022 27858 -43021
rect 25670 -43378 25770 -43022
rect 24020 -43478 25770 -43378
rect 51344 -43278 58368 -43184
rect 51344 -43584 55824 -43278
rect 58268 -43584 58368 -43278
rect 51344 -43984 58368 -43584
rect 7368 -44948 7468 -44667
rect 8160 -44668 8262 -44652
rect 8160 -44948 8260 -44668
rect -28470 -45345 -28370 -45042
rect -29096 -45346 -27774 -45345
rect -29096 -46666 -29095 -45346
rect -27775 -45938 -27774 -45346
rect -27640 -45370 -27540 -45042
rect -26348 -45345 -26248 -45042
rect -27640 -45938 -27620 -45370
rect -27775 -46038 -27620 -45938
rect -27775 -46666 -27774 -46038
rect -29096 -46667 -27774 -46666
rect -27640 -46652 -27620 -46038
rect -27556 -46652 -27540 -45370
rect -28470 -46950 -28370 -46667
rect -27640 -46950 -27540 -46652
rect -26990 -45346 -25668 -45345
rect -26990 -46666 -26989 -45346
rect -25669 -46666 -25668 -45346
rect -26990 -46667 -25668 -46666
rect -25530 -45370 -25434 -45344
rect -24242 -45345 -24142 -45042
rect -25530 -46652 -25514 -45370
rect -25450 -46652 -25434 -45370
rect -26348 -46950 -26248 -46667
rect -25530 -46668 -25434 -46652
rect -24884 -45346 -23562 -45345
rect -24884 -46666 -24883 -45346
rect -23563 -46666 -23562 -45346
rect -24884 -46667 -23562 -46666
rect -23424 -45370 -23328 -45344
rect -22136 -45345 -22036 -45042
rect -23424 -46652 -23408 -45370
rect -23344 -46652 -23328 -45370
rect -24242 -46950 -24142 -46667
rect -23424 -46668 -23328 -46652
rect -22778 -45346 -21456 -45345
rect -22778 -46666 -22777 -45346
rect -21457 -46666 -21456 -45346
rect -22778 -46667 -21456 -46666
rect -21318 -45370 -21222 -45344
rect -20030 -45345 -19930 -45042
rect -21318 -46652 -21302 -45370
rect -21238 -46652 -21222 -45370
rect -22136 -46950 -22036 -46667
rect -21318 -46668 -21222 -46652
rect -20672 -45346 -19350 -45345
rect -20672 -46666 -20671 -45346
rect -19351 -46666 -19350 -45346
rect -20672 -46667 -19350 -46666
rect -19212 -45370 -19116 -45344
rect -17924 -45345 -17824 -45042
rect -19212 -46652 -19196 -45370
rect -19132 -46652 -19116 -45370
rect -20030 -46950 -19930 -46667
rect -19212 -46668 -19116 -46652
rect -18566 -45346 -17244 -45345
rect -18566 -46666 -18565 -45346
rect -17245 -46666 -17244 -45346
rect -18566 -46667 -17244 -46666
rect -17106 -45370 -17010 -45344
rect -15818 -45345 -15718 -45042
rect -17106 -46652 -17090 -45370
rect -17026 -46652 -17010 -45370
rect -17924 -46950 -17824 -46667
rect -17106 -46668 -17010 -46652
rect -16460 -45346 -15138 -45345
rect -16460 -46666 -16459 -45346
rect -15139 -46666 -15138 -45346
rect -16460 -46667 -15138 -46666
rect -15000 -45370 -14904 -45344
rect -13712 -45345 -13612 -45042
rect -15000 -46652 -14984 -45370
rect -14920 -46652 -14904 -45370
rect -15818 -46950 -15718 -46667
rect -15000 -46668 -14904 -46652
rect -14354 -45346 -13032 -45345
rect -14354 -46666 -14353 -45346
rect -13033 -46666 -13032 -45346
rect -14354 -46667 -13032 -46666
rect -12894 -45370 -12798 -45344
rect -11606 -45345 -11506 -45042
rect -12894 -46652 -12878 -45370
rect -12814 -46652 -12798 -45370
rect -13712 -46950 -13612 -46667
rect -12894 -46668 -12798 -46652
rect -12248 -45346 -10926 -45345
rect -12248 -46666 -12247 -45346
rect -10927 -46666 -10926 -45346
rect -10788 -45370 -10692 -45344
rect -9500 -45345 -9400 -45042
rect -10788 -46420 -10772 -45370
rect -12248 -46667 -10926 -46666
rect -10794 -46652 -10772 -46420
rect -10708 -46652 -10692 -45370
rect -11606 -46950 -11506 -46667
rect -28470 -47050 -11506 -46950
rect -10794 -46668 -10692 -46652
rect -10142 -45346 -8820 -45345
rect -10142 -46666 -10141 -45346
rect -8821 -46666 -8820 -45346
rect -8682 -45370 -8586 -45344
rect -8682 -46382 -8666 -45370
rect -10142 -46667 -8820 -46666
rect -8688 -46652 -8666 -46382
rect -8602 -46652 -8586 -45370
rect -10794 -46922 -10694 -46668
rect -10794 -47022 -10292 -46922
rect -28470 -47345 -28370 -47050
rect -29096 -47346 -27774 -47345
rect -29096 -48666 -29095 -47346
rect -27775 -47938 -27774 -47346
rect -27640 -47370 -27540 -47050
rect -26348 -47345 -26248 -47050
rect -27640 -47938 -27620 -47370
rect -27775 -48038 -27620 -47938
rect -27775 -48666 -27774 -48038
rect -29096 -48667 -27774 -48666
rect -27640 -48652 -27620 -48038
rect -27556 -48652 -27540 -47370
rect -28470 -48952 -28370 -48667
rect -27640 -48952 -27540 -48652
rect -26990 -47346 -25668 -47345
rect -26990 -48666 -26989 -47346
rect -25669 -48666 -25668 -47346
rect -26990 -48667 -25668 -48666
rect -25530 -47370 -25434 -47344
rect -24242 -47345 -24142 -47050
rect -25530 -48652 -25514 -47370
rect -25450 -48652 -25434 -47370
rect -26348 -48952 -26248 -48667
rect -25530 -48668 -25434 -48652
rect -24884 -47346 -23562 -47345
rect -24884 -48666 -24883 -47346
rect -23563 -48666 -23562 -47346
rect -24884 -48667 -23562 -48666
rect -23424 -47370 -23328 -47344
rect -22136 -47345 -22036 -47050
rect -23424 -48652 -23408 -47370
rect -23344 -48652 -23328 -47370
rect -24242 -48952 -24142 -48667
rect -23424 -48668 -23328 -48652
rect -22778 -47346 -21456 -47345
rect -22778 -48666 -22777 -47346
rect -21457 -48666 -21456 -47346
rect -22778 -48667 -21456 -48666
rect -21318 -47370 -21222 -47344
rect -20030 -47345 -19930 -47050
rect -21318 -48652 -21302 -47370
rect -21238 -48652 -21222 -47370
rect -22136 -48952 -22036 -48667
rect -21318 -48668 -21222 -48652
rect -20672 -47346 -19350 -47345
rect -20672 -48666 -20671 -47346
rect -19351 -48666 -19350 -47346
rect -20672 -48667 -19350 -48666
rect -19212 -47370 -19116 -47344
rect -17924 -47345 -17824 -47050
rect -19212 -48652 -19196 -47370
rect -19132 -48652 -19116 -47370
rect -20030 -48952 -19930 -48667
rect -19212 -48668 -19116 -48652
rect -18566 -47346 -17244 -47345
rect -18566 -48666 -18565 -47346
rect -17245 -48666 -17244 -47346
rect -18566 -48667 -17244 -48666
rect -17106 -47370 -17010 -47344
rect -15818 -47345 -15718 -47050
rect -17106 -48652 -17090 -47370
rect -17026 -48652 -17010 -47370
rect -17924 -48952 -17824 -48667
rect -17106 -48668 -17010 -48652
rect -16460 -47346 -15138 -47345
rect -16460 -48666 -16459 -47346
rect -15139 -48666 -15138 -47346
rect -16460 -48667 -15138 -48666
rect -15000 -47370 -14904 -47344
rect -13712 -47345 -13612 -47050
rect -15000 -48652 -14984 -47370
rect -14920 -48486 -14904 -47370
rect -14354 -47346 -13032 -47345
rect -14920 -48652 -14900 -48486
rect -15818 -48952 -15718 -48667
rect -28470 -49052 -15718 -48952
rect -15000 -48900 -14900 -48652
rect -14354 -48666 -14353 -47346
rect -13033 -48666 -13032 -47346
rect -12894 -47370 -12798 -47344
rect -11606 -47345 -11506 -47050
rect -12894 -48394 -12878 -47370
rect -14354 -48667 -13032 -48666
rect -12906 -48652 -12878 -48394
rect -12814 -48652 -12798 -47370
rect -15000 -49000 -14652 -48900
rect -28470 -49345 -28370 -49052
rect -29096 -49346 -27774 -49345
rect -29096 -50666 -29095 -49346
rect -27775 -49938 -27774 -49346
rect -27640 -49370 -27540 -49052
rect -26348 -49345 -26248 -49052
rect -27640 -49938 -27620 -49370
rect -27775 -50038 -27620 -49938
rect -27775 -50666 -27774 -50038
rect -29096 -50667 -27774 -50666
rect -27640 -50652 -27620 -50038
rect -27556 -50652 -27540 -49370
rect -28470 -50966 -28370 -50667
rect -27640 -50966 -27540 -50652
rect -26990 -49346 -25668 -49345
rect -26990 -50666 -26989 -49346
rect -25669 -50666 -25668 -49346
rect -26990 -50667 -25668 -50666
rect -25530 -49370 -25434 -49344
rect -24242 -49345 -24142 -49052
rect -25530 -50652 -25514 -49370
rect -25450 -50652 -25434 -49370
rect -26348 -50966 -26248 -50667
rect -25530 -50668 -25434 -50652
rect -24884 -49346 -23562 -49345
rect -24884 -50666 -24883 -49346
rect -23563 -50666 -23562 -49346
rect -24884 -50667 -23562 -50666
rect -23424 -49370 -23328 -49344
rect -22136 -49345 -22036 -49052
rect -23424 -50652 -23408 -49370
rect -23344 -50652 -23328 -49370
rect -24242 -50966 -24142 -50667
rect -23424 -50668 -23328 -50652
rect -22778 -49346 -21456 -49345
rect -22778 -50666 -22777 -49346
rect -21457 -50666 -21456 -49346
rect -22778 -50667 -21456 -50666
rect -21318 -49370 -21222 -49344
rect -20030 -49345 -19930 -49052
rect -21318 -50652 -21302 -49370
rect -21238 -50652 -21222 -49370
rect -22136 -50966 -22036 -50667
rect -21318 -50668 -21222 -50652
rect -20672 -49346 -19350 -49345
rect -20672 -50666 -20671 -49346
rect -19351 -50666 -19350 -49346
rect -20672 -50667 -19350 -50666
rect -19212 -49370 -19116 -49344
rect -17924 -49345 -17824 -49052
rect -19212 -50652 -19196 -49370
rect -19132 -50652 -19116 -49370
rect -20030 -50966 -19930 -50667
rect -19212 -50668 -19116 -50652
rect -18566 -49346 -17244 -49345
rect -18566 -50666 -18565 -49346
rect -17245 -50666 -17244 -49346
rect -18566 -50667 -17244 -50666
rect -17106 -49370 -17010 -49344
rect -15818 -49345 -15718 -49052
rect -17106 -50652 -17090 -49370
rect -17026 -50652 -17010 -49370
rect -17924 -50966 -17824 -50667
rect -17106 -50668 -17010 -50652
rect -16460 -49346 -15138 -49345
rect -16460 -50666 -16459 -49346
rect -15139 -50666 -15138 -49346
rect -16460 -50667 -15138 -50666
rect -15000 -49370 -14904 -49344
rect -15000 -50652 -14984 -49370
rect -14920 -50652 -14904 -49370
rect -15818 -50966 -15718 -50667
rect -15000 -50668 -14904 -50652
rect -28470 -51066 -15718 -50966
rect -28470 -51345 -28370 -51066
rect -29096 -51346 -27774 -51345
rect -29096 -52666 -29095 -51346
rect -27775 -51938 -27774 -51346
rect -27640 -51370 -27540 -51066
rect -26348 -51345 -26248 -51066
rect -27640 -51938 -27620 -51370
rect -27775 -52038 -27620 -51938
rect -27775 -52666 -27774 -52038
rect -29096 -52667 -27774 -52666
rect -27640 -52652 -27620 -52038
rect -27556 -52652 -27540 -51370
rect -28470 -52962 -28370 -52667
rect -27640 -52962 -27540 -52652
rect -26990 -51346 -25668 -51345
rect -26990 -52666 -26989 -51346
rect -25669 -52666 -25668 -51346
rect -26990 -52667 -25668 -52666
rect -25530 -51370 -25434 -51344
rect -24242 -51345 -24142 -51066
rect -25530 -52652 -25514 -51370
rect -25450 -52652 -25434 -51370
rect -26348 -52962 -26248 -52667
rect -25530 -52668 -25434 -52652
rect -24884 -51346 -23562 -51345
rect -24884 -52666 -24883 -51346
rect -23563 -52666 -23562 -51346
rect -24884 -52667 -23562 -52666
rect -23424 -51370 -23328 -51344
rect -22136 -51345 -22036 -51066
rect -23424 -52652 -23408 -51370
rect -23344 -52652 -23328 -51370
rect -24242 -52962 -24142 -52667
rect -23424 -52668 -23328 -52652
rect -22778 -51346 -21456 -51345
rect -22778 -52666 -22777 -51346
rect -21457 -52666 -21456 -51346
rect -22778 -52667 -21456 -52666
rect -21318 -51370 -21222 -51344
rect -20030 -51345 -19930 -51066
rect -21318 -52652 -21302 -51370
rect -21238 -52652 -21222 -51370
rect -22136 -52962 -22036 -52667
rect -21318 -52668 -21222 -52652
rect -20672 -51346 -19350 -51345
rect -20672 -52666 -20671 -51346
rect -19351 -52666 -19350 -51346
rect -20672 -52667 -19350 -52666
rect -19212 -51370 -19116 -51344
rect -17924 -51345 -17824 -51066
rect -19212 -52652 -19196 -51370
rect -19132 -52652 -19116 -51370
rect -20030 -52962 -19930 -52667
rect -19212 -52668 -19116 -52652
rect -18566 -51346 -17244 -51345
rect -18566 -52666 -18565 -51346
rect -17245 -52666 -17244 -51346
rect -17106 -51370 -17010 -51344
rect -15818 -51345 -15718 -51066
rect -17106 -52416 -17090 -51370
rect -18566 -52667 -17244 -52666
rect -17114 -52652 -17090 -52416
rect -17026 -52652 -17010 -51370
rect -17924 -52962 -17824 -52667
rect -28470 -53062 -17824 -52962
rect -28470 -53345 -28370 -53062
rect -29096 -53346 -27774 -53345
rect -29096 -54666 -29095 -53346
rect -27775 -53938 -27774 -53346
rect -27640 -53370 -27540 -53062
rect -26348 -53345 -26248 -53062
rect -27640 -53938 -27620 -53370
rect -27775 -54038 -27620 -53938
rect -27775 -54666 -27774 -54038
rect -29096 -54667 -27774 -54666
rect -27640 -54652 -27620 -54038
rect -27556 -54652 -27540 -53370
rect -28470 -54956 -28370 -54667
rect -27640 -54956 -27540 -54652
rect -26990 -53346 -25668 -53345
rect -26990 -54666 -26989 -53346
rect -25669 -54666 -25668 -53346
rect -26990 -54667 -25668 -54666
rect -25530 -53370 -25434 -53344
rect -24242 -53345 -24142 -53062
rect -25530 -54652 -25514 -53370
rect -25450 -54652 -25434 -53370
rect -26348 -54956 -26248 -54667
rect -25530 -54668 -25434 -54652
rect -24884 -53346 -23562 -53345
rect -24884 -54666 -24883 -53346
rect -23563 -54666 -23562 -53346
rect -24884 -54667 -23562 -54666
rect -23424 -53370 -23328 -53344
rect -22136 -53345 -22036 -53062
rect -23424 -54652 -23408 -53370
rect -23344 -54652 -23328 -53370
rect -24242 -54956 -24142 -54667
rect -23424 -54668 -23328 -54652
rect -22778 -53346 -21456 -53345
rect -22778 -54666 -22777 -53346
rect -21457 -54666 -21456 -53346
rect -22778 -54667 -21456 -54666
rect -21318 -53370 -21222 -53344
rect -20030 -53345 -19930 -53062
rect -21318 -54652 -21302 -53370
rect -21238 -54652 -21222 -53370
rect -22136 -54956 -22036 -54667
rect -21318 -54668 -21222 -54652
rect -20672 -53346 -19350 -53345
rect -20672 -54666 -20671 -53346
rect -19351 -54666 -19350 -53346
rect -20672 -54667 -19350 -54666
rect -19212 -53370 -19116 -53344
rect -17924 -53345 -17824 -53062
rect -17114 -52668 -17010 -52652
rect -16460 -51346 -15138 -51345
rect -16460 -52666 -16459 -51346
rect -15139 -52666 -15138 -51346
rect -16460 -52667 -15138 -52666
rect -15000 -51370 -14904 -51344
rect -15000 -52652 -14984 -51370
rect -14920 -52652 -14904 -51370
rect -17114 -52968 -17014 -52668
rect -17114 -53068 -16748 -52968
rect -19212 -54652 -19196 -53370
rect -19132 -54450 -19116 -53370
rect -18566 -53346 -17244 -53345
rect -19132 -54652 -19112 -54450
rect -20030 -54956 -19930 -54667
rect -28470 -55056 -19930 -54956
rect -19212 -54926 -19112 -54652
rect -18566 -54666 -18565 -53346
rect -17245 -54666 -17244 -53346
rect -18566 -54667 -17244 -54666
rect -17106 -53370 -17010 -53344
rect -17106 -54652 -17090 -53370
rect -17026 -54652 -17010 -53370
rect -19212 -55026 -18864 -54926
rect -28470 -55345 -28370 -55056
rect -29096 -55346 -27774 -55345
rect -29096 -56666 -29095 -55346
rect -27775 -55938 -27774 -55346
rect -27640 -55370 -27540 -55056
rect -26348 -55345 -26248 -55056
rect -27640 -55938 -27620 -55370
rect -27775 -56038 -27620 -55938
rect -27775 -56666 -27774 -56038
rect -29096 -56667 -27774 -56666
rect -27640 -56652 -27620 -56038
rect -27556 -56652 -27540 -55370
rect -28470 -56966 -28370 -56667
rect -27640 -56966 -27540 -56652
rect -26990 -55346 -25668 -55345
rect -26990 -56666 -26989 -55346
rect -25669 -56666 -25668 -55346
rect -26990 -56667 -25668 -56666
rect -25530 -55370 -25434 -55344
rect -24242 -55345 -24142 -55056
rect -25530 -56652 -25514 -55370
rect -25450 -56652 -25434 -55370
rect -26348 -56966 -26248 -56667
rect -25530 -56668 -25434 -56652
rect -24884 -55346 -23562 -55345
rect -24884 -56666 -24883 -55346
rect -23563 -56666 -23562 -55346
rect -24884 -56667 -23562 -56666
rect -23424 -55370 -23328 -55344
rect -22136 -55345 -22036 -55056
rect -23424 -56652 -23408 -55370
rect -23344 -56652 -23328 -55370
rect -24242 -56966 -24142 -56667
rect -23424 -56668 -23328 -56652
rect -22778 -55346 -21456 -55345
rect -22778 -56666 -22777 -55346
rect -21457 -56666 -21456 -55346
rect -22778 -56667 -21456 -56666
rect -21318 -55370 -21222 -55344
rect -20030 -55345 -19930 -55056
rect -21318 -56652 -21302 -55370
rect -21238 -56652 -21222 -55370
rect -22136 -56966 -22036 -56667
rect -21318 -56668 -21222 -56652
rect -20672 -55346 -19350 -55345
rect -20672 -56666 -20671 -55346
rect -19351 -56666 -19350 -55346
rect -20672 -56667 -19350 -56666
rect -19212 -55370 -19116 -55344
rect -19212 -56652 -19196 -55370
rect -19132 -56652 -19116 -55370
rect -20030 -56966 -19930 -56667
rect -19212 -56668 -19116 -56652
rect -28470 -57066 -19930 -56966
rect -28470 -57345 -28370 -57066
rect -29096 -57346 -27774 -57345
rect -29096 -58666 -29095 -57346
rect -27775 -57938 -27774 -57346
rect -27640 -57370 -27540 -57066
rect -26348 -57345 -26248 -57066
rect -27640 -57938 -27620 -57370
rect -27775 -58038 -27620 -57938
rect -27775 -58666 -27774 -58038
rect -29096 -58667 -27774 -58666
rect -27640 -58652 -27620 -58038
rect -27556 -58652 -27540 -57370
rect -28470 -58934 -28370 -58667
rect -27640 -58934 -27540 -58652
rect -26990 -57346 -25668 -57345
rect -26990 -58666 -26989 -57346
rect -25669 -58666 -25668 -57346
rect -26990 -58667 -25668 -58666
rect -25530 -57370 -25434 -57344
rect -24242 -57345 -24142 -57066
rect -25530 -58652 -25514 -57370
rect -25450 -58652 -25434 -57370
rect -26348 -58934 -26248 -58667
rect -25530 -58668 -25434 -58652
rect -24884 -57346 -23562 -57345
rect -24884 -58666 -24883 -57346
rect -23563 -58666 -23562 -57346
rect -24884 -58667 -23562 -58666
rect -23424 -57370 -23328 -57344
rect -22136 -57345 -22036 -57066
rect -23424 -58652 -23408 -57370
rect -23344 -58652 -23328 -57370
rect -24242 -58934 -24142 -58667
rect -23424 -58668 -23328 -58652
rect -22778 -57346 -21456 -57345
rect -22778 -58666 -22777 -57346
rect -21457 -58666 -21456 -57346
rect -22778 -58667 -21456 -58666
rect -21318 -57370 -21222 -57344
rect -20030 -57345 -19930 -57066
rect -21318 -58652 -21302 -57370
rect -21238 -58652 -21222 -57370
rect -22136 -58934 -22036 -58667
rect -21318 -58668 -21222 -58652
rect -20672 -57346 -19350 -57345
rect -20672 -58666 -20671 -57346
rect -19351 -58666 -19350 -57346
rect -20672 -58667 -19350 -58666
rect -19212 -57370 -19116 -57344
rect -19212 -58652 -19196 -57370
rect -19132 -58652 -19116 -57370
rect -20030 -58934 -19930 -58667
rect -19212 -58668 -19116 -58652
rect -28470 -59034 -19930 -58934
rect -28470 -59345 -28370 -59034
rect -29096 -59346 -27774 -59345
rect -29096 -60666 -29095 -59346
rect -27775 -59938 -27774 -59346
rect -27640 -59370 -27540 -59034
rect -26348 -59345 -26248 -59034
rect -27640 -59938 -27620 -59370
rect -27775 -60038 -27620 -59938
rect -27775 -60666 -27774 -60038
rect -29096 -60667 -27774 -60666
rect -27640 -60652 -27620 -60038
rect -27556 -60652 -27540 -59370
rect -28470 -60942 -28370 -60667
rect -27640 -60942 -27540 -60652
rect -26990 -59346 -25668 -59345
rect -26990 -60666 -26989 -59346
rect -25669 -60666 -25668 -59346
rect -26990 -60667 -25668 -60666
rect -25530 -59370 -25434 -59344
rect -24242 -59345 -24142 -59034
rect -25530 -60652 -25514 -59370
rect -25450 -60652 -25434 -59370
rect -26348 -60942 -26248 -60667
rect -28470 -61042 -26248 -60942
rect -25530 -60938 -25434 -60652
rect -24884 -59346 -23562 -59345
rect -24884 -60666 -24883 -59346
rect -23563 -60666 -23562 -59346
rect -24884 -60667 -23562 -60666
rect -23424 -59370 -23328 -59344
rect -22136 -59345 -22036 -59034
rect -23424 -60652 -23408 -59370
rect -23344 -60652 -23328 -59370
rect -25530 -61034 -25104 -60938
rect -28470 -61345 -28370 -61042
rect -29096 -61346 -27774 -61345
rect -29096 -62666 -29095 -61346
rect -27775 -61936 -27774 -61346
rect -27640 -61370 -27540 -61042
rect -26348 -61345 -26248 -61042
rect -27640 -61936 -27620 -61370
rect -27775 -62036 -27620 -61936
rect -27775 -62666 -27774 -62036
rect -29096 -62667 -27774 -62666
rect -27636 -62652 -27620 -62036
rect -27556 -61936 -27540 -61370
rect -26990 -61346 -25668 -61345
rect -26990 -61936 -26989 -61346
rect -27556 -62036 -26989 -61936
rect -27556 -62652 -27540 -62036
rect -27636 -62668 -27540 -62652
rect -26990 -62666 -26989 -62036
rect -25669 -61936 -25668 -61346
rect -25530 -61370 -25434 -61344
rect -25530 -61936 -25514 -61370
rect -25669 -62036 -25514 -61936
rect -25669 -62666 -25668 -62036
rect -26990 -62667 -25668 -62666
rect -25530 -62652 -25514 -62036
rect -25450 -62652 -25434 -61370
rect -25530 -62668 -25434 -62652
rect -25200 -63050 -25104 -61034
rect -24242 -60942 -24142 -60667
rect -23424 -60668 -23328 -60652
rect -22778 -59346 -21456 -59345
rect -22778 -60666 -22777 -59346
rect -21457 -60666 -21456 -59346
rect -22778 -60667 -21456 -60666
rect -21318 -59370 -21222 -59344
rect -20030 -59345 -19930 -59034
rect -21318 -60652 -21302 -59370
rect -21238 -60652 -21222 -59370
rect -22136 -60942 -22036 -60667
rect -21318 -60668 -21222 -60652
rect -20672 -59346 -19350 -59345
rect -20672 -60666 -20671 -59346
rect -19351 -60666 -19350 -59346
rect -20672 -60667 -19350 -60666
rect -19212 -59370 -19116 -59344
rect -19212 -60652 -19196 -59370
rect -19132 -60652 -19116 -59370
rect -20030 -60942 -19930 -60667
rect -19212 -60668 -19116 -60652
rect -24242 -61042 -19930 -60942
rect -24242 -61345 -24142 -61042
rect -24884 -61346 -23562 -61345
rect -24884 -62666 -24883 -61346
rect -23563 -61930 -23562 -61346
rect -23424 -61370 -23328 -61344
rect -22136 -61345 -22036 -61042
rect -23424 -61930 -23408 -61370
rect -23563 -62036 -23408 -61930
rect -23563 -62666 -23562 -62036
rect -24884 -62667 -23562 -62666
rect -23424 -62652 -23408 -62036
rect -23344 -61936 -23328 -61370
rect -22778 -61346 -21456 -61345
rect -22778 -61936 -22777 -61346
rect -23344 -62036 -22777 -61936
rect -23344 -62652 -23328 -62036
rect -23424 -62668 -23328 -62652
rect -22778 -62666 -22777 -62036
rect -21457 -61930 -21456 -61346
rect -21318 -61370 -21222 -61344
rect -20030 -61345 -19930 -61042
rect -21318 -61930 -21302 -61370
rect -21457 -62036 -21302 -61930
rect -21457 -62666 -21456 -62036
rect -22778 -62667 -21456 -62666
rect -21318 -62652 -21302 -62036
rect -21238 -61936 -21222 -61370
rect -20672 -61346 -19350 -61345
rect -20672 -61936 -20671 -61346
rect -21238 -62036 -20671 -61936
rect -21238 -62652 -21222 -62036
rect -21318 -62668 -21222 -62652
rect -20672 -62666 -20671 -62036
rect -19351 -61930 -19350 -61346
rect -19212 -61370 -19116 -61344
rect -19212 -61930 -19196 -61370
rect -19351 -62030 -19196 -61930
rect -19351 -62666 -19350 -62030
rect -20672 -62667 -19350 -62666
rect -19212 -62652 -19196 -62030
rect -19132 -62652 -19116 -61370
rect -19212 -62668 -19116 -62652
rect -18964 -63015 -18864 -55026
rect -17924 -55345 -17824 -54667
rect -17106 -54668 -17010 -54652
rect -18566 -55346 -17244 -55345
rect -18566 -56666 -18565 -55346
rect -17245 -56666 -17244 -55346
rect -18566 -56667 -17244 -56666
rect -17106 -55370 -17010 -55344
rect -17106 -56652 -17090 -55370
rect -17026 -56652 -17010 -55370
rect -17924 -57345 -17824 -56667
rect -17106 -56668 -17010 -56652
rect -18566 -57346 -17244 -57345
rect -18566 -58666 -18565 -57346
rect -17245 -58666 -17244 -57346
rect -18566 -58667 -17244 -58666
rect -17106 -57370 -17010 -57344
rect -17106 -58652 -17090 -57370
rect -17026 -58652 -17010 -57370
rect -17924 -59345 -17824 -58667
rect -17106 -58668 -17010 -58652
rect -18566 -59346 -17244 -59345
rect -18566 -60666 -18565 -59346
rect -17245 -60666 -17244 -59346
rect -18566 -60667 -17244 -60666
rect -17106 -59370 -17010 -59344
rect -17106 -60652 -17090 -59370
rect -17026 -60652 -17010 -59370
rect -17924 -61345 -17824 -60667
rect -17106 -60668 -17010 -60652
rect -18566 -61346 -17244 -61345
rect -18566 -62666 -18565 -61346
rect -17245 -61930 -17244 -61346
rect -17106 -61370 -17010 -61344
rect -17106 -61930 -17090 -61370
rect -17245 -62030 -17090 -61930
rect -17245 -62666 -17244 -62030
rect -18566 -62667 -17244 -62666
rect -17106 -62652 -17090 -62030
rect -17026 -62652 -17010 -61370
rect -17106 -62668 -17010 -62652
rect -25200 -63277 -25100 -63050
rect -18964 -63113 -18963 -63015
rect -18865 -63113 -18864 -63015
rect -16848 -63011 -16748 -53068
rect -15818 -53345 -15718 -52667
rect -15000 -52668 -14904 -52652
rect -16460 -53346 -15138 -53345
rect -16460 -54666 -16459 -53346
rect -15139 -54666 -15138 -53346
rect -16460 -54667 -15138 -54666
rect -15000 -53370 -14904 -53344
rect -15000 -54652 -14984 -53370
rect -14920 -54652 -14904 -53370
rect -15818 -55345 -15718 -54667
rect -15000 -54668 -14904 -54652
rect -16460 -55346 -15138 -55345
rect -16460 -56666 -16459 -55346
rect -15139 -56666 -15138 -55346
rect -16460 -56667 -15138 -56666
rect -15000 -55370 -14904 -55344
rect -15000 -56652 -14984 -55370
rect -14920 -56652 -14904 -55370
rect -15818 -57345 -15718 -56667
rect -15000 -56668 -14904 -56652
rect -16460 -57346 -15138 -57345
rect -16460 -58666 -16459 -57346
rect -15139 -58666 -15138 -57346
rect -16460 -58667 -15138 -58666
rect -15000 -57370 -14904 -57344
rect -15000 -58652 -14984 -57370
rect -14920 -58652 -14904 -57370
rect -15818 -59345 -15718 -58667
rect -15000 -58668 -14904 -58652
rect -16460 -59346 -15138 -59345
rect -16460 -60666 -16459 -59346
rect -15139 -60666 -15138 -59346
rect -16460 -60667 -15138 -60666
rect -15000 -59370 -14904 -59344
rect -15000 -60652 -14984 -59370
rect -14920 -60652 -14904 -59370
rect -15818 -61345 -15718 -60667
rect -15000 -60668 -14904 -60652
rect -16460 -61346 -15138 -61345
rect -16460 -62666 -16459 -61346
rect -15139 -61930 -15138 -61346
rect -15000 -61370 -14904 -61344
rect -15000 -61930 -14984 -61370
rect -15139 -62030 -14984 -61930
rect -15139 -62666 -15138 -62030
rect -16460 -62667 -15138 -62666
rect -15000 -62652 -14984 -62030
rect -14920 -62652 -14904 -61370
rect -15000 -62668 -14904 -62652
rect -16848 -63109 -16847 -63011
rect -16749 -63109 -16748 -63011
rect -14752 -63009 -14652 -49000
rect -13712 -49345 -13612 -48667
rect -12906 -48668 -12798 -48652
rect -12248 -47346 -10926 -47345
rect -12248 -48666 -12247 -47346
rect -10927 -48666 -10926 -47346
rect -10788 -47370 -10692 -47344
rect -10788 -48326 -10772 -47370
rect -12248 -48667 -10926 -48666
rect -10794 -48652 -10772 -48326
rect -10708 -48652 -10692 -47370
rect -12906 -48898 -12806 -48668
rect -12906 -48998 -12528 -48898
rect -14354 -49346 -13032 -49345
rect -14354 -50666 -14353 -49346
rect -13033 -50666 -13032 -49346
rect -14354 -50667 -13032 -50666
rect -12894 -49370 -12798 -49344
rect -12894 -50652 -12878 -49370
rect -12814 -50652 -12798 -49370
rect -13712 -51345 -13612 -50667
rect -12894 -50668 -12798 -50652
rect -14354 -51346 -13032 -51345
rect -14354 -52666 -14353 -51346
rect -13033 -52666 -13032 -51346
rect -14354 -52667 -13032 -52666
rect -12894 -51370 -12798 -51344
rect -12894 -52652 -12878 -51370
rect -12814 -52652 -12798 -51370
rect -13712 -53345 -13612 -52667
rect -12894 -52668 -12798 -52652
rect -14354 -53346 -13032 -53345
rect -14354 -54666 -14353 -53346
rect -13033 -54666 -13032 -53346
rect -14354 -54667 -13032 -54666
rect -12894 -53370 -12798 -53344
rect -12894 -54652 -12878 -53370
rect -12814 -54652 -12798 -53370
rect -13712 -55345 -13612 -54667
rect -12894 -54668 -12798 -54652
rect -14354 -55346 -13032 -55345
rect -14354 -56666 -14353 -55346
rect -13033 -56666 -13032 -55346
rect -14354 -56667 -13032 -56666
rect -12894 -55370 -12798 -55344
rect -12894 -56652 -12878 -55370
rect -12814 -56652 -12798 -55370
rect -13712 -57345 -13612 -56667
rect -12894 -56668 -12798 -56652
rect -14354 -57346 -13032 -57345
rect -14354 -58666 -14353 -57346
rect -13033 -58666 -13032 -57346
rect -14354 -58667 -13032 -58666
rect -12894 -57370 -12798 -57344
rect -12894 -58652 -12878 -57370
rect -12814 -58652 -12798 -57370
rect -13712 -59345 -13612 -58667
rect -12894 -58668 -12798 -58652
rect -14354 -59346 -13032 -59345
rect -14354 -60666 -14353 -59346
rect -13033 -60666 -13032 -59346
rect -14354 -60667 -13032 -60666
rect -12894 -59370 -12798 -59344
rect -12894 -60652 -12878 -59370
rect -12814 -60652 -12798 -59370
rect -13712 -61345 -13612 -60667
rect -12894 -60668 -12798 -60652
rect -14354 -61346 -13032 -61345
rect -14354 -62666 -14353 -61346
rect -13033 -61930 -13032 -61346
rect -12894 -61370 -12798 -61344
rect -12894 -61930 -12878 -61370
rect -13033 -62030 -12878 -61930
rect -13033 -62666 -13032 -62030
rect -14354 -62667 -13032 -62666
rect -12894 -62652 -12878 -62030
rect -12814 -62652 -12798 -61370
rect -12894 -62668 -12798 -62652
rect -14752 -63107 -14751 -63009
rect -14653 -63107 -14652 -63009
rect -14752 -63108 -14652 -63107
rect -12628 -63019 -12528 -48998
rect -11606 -49345 -11506 -48667
rect -10794 -48668 -10692 -48652
rect -10794 -48956 -10694 -48668
rect -10794 -49056 -10492 -48956
rect -12248 -49346 -10926 -49345
rect -12248 -50666 -12247 -49346
rect -10927 -50666 -10926 -49346
rect -12248 -50667 -10926 -50666
rect -10788 -49370 -10692 -49344
rect -10788 -50652 -10772 -49370
rect -10708 -50652 -10692 -49370
rect -11606 -51345 -11506 -50667
rect -10788 -50668 -10692 -50652
rect -12248 -51346 -10926 -51345
rect -12248 -52666 -12247 -51346
rect -10927 -52666 -10926 -51346
rect -12248 -52667 -10926 -52666
rect -10788 -51370 -10692 -51344
rect -10788 -52652 -10772 -51370
rect -10708 -52652 -10692 -51370
rect -11606 -53345 -11506 -52667
rect -10788 -52668 -10692 -52652
rect -12248 -53346 -10926 -53345
rect -12248 -54666 -12247 -53346
rect -10927 -54666 -10926 -53346
rect -12248 -54667 -10926 -54666
rect -10788 -53370 -10692 -53344
rect -10788 -54652 -10772 -53370
rect -10708 -54652 -10692 -53370
rect -11606 -55345 -11506 -54667
rect -10788 -54668 -10692 -54652
rect -12248 -55346 -10926 -55345
rect -12248 -56666 -12247 -55346
rect -10927 -56666 -10926 -55346
rect -12248 -56667 -10926 -56666
rect -10788 -55370 -10692 -55344
rect -10788 -56652 -10772 -55370
rect -10708 -56652 -10692 -55370
rect -11606 -57345 -11506 -56667
rect -10788 -56668 -10692 -56652
rect -12248 -57346 -10926 -57345
rect -12248 -58666 -12247 -57346
rect -10927 -58666 -10926 -57346
rect -12248 -58667 -10926 -58666
rect -10788 -57370 -10692 -57344
rect -10788 -58652 -10772 -57370
rect -10708 -58652 -10692 -57370
rect -11606 -59345 -11506 -58667
rect -10788 -58668 -10692 -58652
rect -12248 -59346 -10926 -59345
rect -12248 -60666 -12247 -59346
rect -10927 -60666 -10926 -59346
rect -12248 -60667 -10926 -60666
rect -10788 -59370 -10692 -59344
rect -10788 -60652 -10772 -59370
rect -10708 -60652 -10692 -59370
rect -11606 -61345 -11506 -60667
rect -10788 -60668 -10692 -60652
rect -12248 -61346 -10926 -61345
rect -12248 -62666 -12247 -61346
rect -10927 -61930 -10926 -61346
rect -10788 -61370 -10692 -61344
rect -10788 -61930 -10772 -61370
rect -10927 -62030 -10772 -61930
rect -10927 -62666 -10926 -62030
rect -12248 -62667 -10926 -62666
rect -10788 -62652 -10772 -62030
rect -10708 -62652 -10692 -61370
rect -10788 -62668 -10692 -62652
rect -16848 -63110 -16748 -63109
rect -18964 -63114 -18864 -63113
rect -12628 -63117 -12627 -63019
rect -12529 -63117 -12528 -63019
rect -10592 -63011 -10492 -49056
rect -10592 -63109 -10591 -63011
rect -10493 -63109 -10492 -63011
rect -10392 -63000 -10292 -47022
rect -9500 -47345 -9400 -46667
rect -8688 -46668 -8586 -46652
rect -8688 -47012 -8588 -46668
rect -8688 -47112 -8396 -47012
rect -10142 -47346 -8820 -47345
rect -10142 -48666 -10141 -47346
rect -8821 -48666 -8820 -47346
rect -10142 -48667 -8820 -48666
rect -8682 -47370 -8586 -47344
rect -8682 -48652 -8666 -47370
rect -8602 -48652 -8586 -47370
rect -9500 -49345 -9400 -48667
rect -8682 -48668 -8586 -48652
rect -10142 -49346 -8820 -49345
rect -10142 -50666 -10141 -49346
rect -8821 -50666 -8820 -49346
rect -10142 -50667 -8820 -50666
rect -8682 -49370 -8586 -49344
rect -8682 -50652 -8666 -49370
rect -8602 -50652 -8586 -49370
rect -9500 -51345 -9400 -50667
rect -8682 -50668 -8586 -50652
rect -10142 -51346 -8820 -51345
rect -10142 -52666 -10141 -51346
rect -8821 -52666 -8820 -51346
rect -10142 -52667 -8820 -52666
rect -8682 -51370 -8586 -51344
rect -8682 -52652 -8666 -51370
rect -8602 -52652 -8586 -51370
rect -9500 -53345 -9400 -52667
rect -8682 -52668 -8586 -52652
rect -10142 -53346 -8820 -53345
rect -10142 -54666 -10141 -53346
rect -8821 -54666 -8820 -53346
rect -10142 -54667 -8820 -54666
rect -8682 -53370 -8586 -53344
rect -8682 -54652 -8666 -53370
rect -8602 -54652 -8586 -53370
rect -9500 -55345 -9400 -54667
rect -8682 -54668 -8586 -54652
rect -10142 -55346 -8820 -55345
rect -10142 -56666 -10141 -55346
rect -8821 -56666 -8820 -55346
rect -10142 -56667 -8820 -56666
rect -8682 -55370 -8586 -55344
rect -8682 -56652 -8666 -55370
rect -8602 -56652 -8586 -55370
rect -9500 -57345 -9400 -56667
rect -8682 -56668 -8586 -56652
rect -10142 -57346 -8820 -57345
rect -10142 -58666 -10141 -57346
rect -8821 -58666 -8820 -57346
rect -10142 -58667 -8820 -58666
rect -8682 -57370 -8586 -57344
rect -8682 -58652 -8666 -57370
rect -8602 -58652 -8586 -57370
rect -9500 -59345 -9400 -58667
rect -8682 -58668 -8586 -58652
rect -10142 -59346 -8820 -59345
rect -10142 -60666 -10141 -59346
rect -8821 -60666 -8820 -59346
rect -10142 -60667 -8820 -60666
rect -8682 -59370 -8586 -59344
rect -8682 -60652 -8666 -59370
rect -8602 -60652 -8586 -59370
rect -9500 -61345 -9400 -60667
rect -8682 -60668 -8586 -60652
rect -10142 -61346 -8820 -61345
rect -10142 -62666 -10141 -61346
rect -8821 -61930 -8820 -61346
rect -8682 -61370 -8586 -61344
rect -8682 -61930 -8666 -61370
rect -8821 -62030 -8666 -61930
rect -8821 -62666 -8820 -62030
rect -10142 -62667 -8820 -62666
rect -8682 -62652 -8666 -62030
rect -8602 -62652 -8586 -61370
rect -8682 -62668 -8586 -62652
rect -10392 -63001 -9838 -63000
rect -10392 -63099 -9937 -63001
rect -9839 -63099 -9838 -63001
rect -10392 -63100 -9838 -63099
rect -8496 -63019 -8396 -47112
rect -10592 -63110 -10492 -63109
rect -12628 -63118 -12528 -63117
rect -8496 -63117 -8495 -63019
rect -8397 -63117 -8396 -63019
rect -8496 -63118 -8396 -63117
rect -8282 -63022 -8182 -44964
rect -7408 -45048 8260 -44948
rect -7394 -45345 -7294 -45048
rect -8036 -45346 -6714 -45345
rect -8036 -46666 -8035 -45346
rect -6715 -46666 -6714 -45346
rect -8036 -46667 -6714 -46666
rect -6576 -45370 -6480 -45344
rect -5288 -45345 -5188 -45048
rect -6576 -46652 -6560 -45370
rect -6496 -46652 -6480 -45370
rect -7394 -46948 -7294 -46667
rect -6576 -46668 -6480 -46652
rect -5930 -45346 -4608 -45345
rect -5930 -46666 -5929 -45346
rect -4609 -46666 -4608 -45346
rect -5930 -46667 -4608 -46666
rect -4470 -45370 -4374 -45344
rect -3182 -45345 -3082 -45048
rect -4470 -46652 -4454 -45370
rect -4390 -46652 -4374 -45370
rect -5288 -46948 -5188 -46667
rect -4470 -46668 -4374 -46652
rect -3824 -45346 -2502 -45345
rect -3824 -46666 -3823 -45346
rect -2503 -46666 -2502 -45346
rect -3824 -46667 -2502 -46666
rect -2364 -45370 -2268 -45344
rect -1076 -45345 -976 -45048
rect -2364 -46652 -2348 -45370
rect -2284 -46652 -2268 -45370
rect -3182 -46948 -3082 -46667
rect -2364 -46668 -2268 -46652
rect -1718 -45346 -396 -45345
rect -1718 -46666 -1717 -45346
rect -397 -46666 -396 -45346
rect -1718 -46667 -396 -46666
rect -258 -45370 -162 -45344
rect 1030 -45345 1130 -45048
rect -258 -46652 -242 -45370
rect -178 -46652 -162 -45370
rect -1076 -46948 -976 -46667
rect -258 -46668 -162 -46652
rect 388 -45346 1710 -45345
rect 388 -46666 389 -45346
rect 1709 -46666 1710 -45346
rect 388 -46667 1710 -46666
rect 1848 -45370 1944 -45344
rect 3136 -45345 3236 -45048
rect 1848 -46652 1864 -45370
rect 1928 -46652 1944 -45370
rect 1030 -46948 1130 -46667
rect 1848 -46668 1944 -46652
rect 2494 -45346 3816 -45345
rect 2494 -46666 2495 -45346
rect 3815 -46666 3816 -45346
rect 2494 -46667 3816 -46666
rect 3954 -45370 4050 -45344
rect 5242 -45345 5342 -45048
rect 3954 -46652 3970 -45370
rect 4034 -46652 4050 -45370
rect 3136 -46948 3236 -46667
rect 3954 -46668 4050 -46652
rect 4600 -45346 5922 -45345
rect 4600 -46666 4601 -45346
rect 5921 -46666 5922 -45346
rect 4600 -46667 5922 -46666
rect 6060 -45370 6156 -45344
rect 7368 -45345 7468 -45048
rect 8160 -45344 8260 -45048
rect 6060 -46652 6076 -45370
rect 6140 -46652 6156 -45370
rect 5242 -46948 5342 -46667
rect 6060 -46668 6156 -46652
rect 6706 -45346 8028 -45345
rect 6706 -46666 6707 -45346
rect 8027 -45942 8028 -45346
rect 8160 -45370 8262 -45344
rect 8160 -45942 8182 -45370
rect 8027 -46042 8182 -45942
rect 8027 -46666 8028 -46042
rect 6706 -46667 8028 -46666
rect 8160 -46652 8182 -46042
rect 8246 -46652 8262 -45370
rect 7368 -46948 7468 -46667
rect 8160 -46668 8262 -46652
rect 8160 -46948 8260 -46668
rect -7394 -47048 8260 -46948
rect -7394 -47345 -7294 -47048
rect -8036 -47346 -6714 -47345
rect -8036 -48666 -8035 -47346
rect -6715 -48666 -6714 -47346
rect -8036 -48667 -6714 -48666
rect -6576 -47370 -6480 -47344
rect -5288 -47345 -5188 -47048
rect -6576 -48652 -6560 -47370
rect -6496 -48652 -6480 -47370
rect -7394 -48948 -7294 -48667
rect -6576 -48668 -6480 -48652
rect -5930 -47346 -4608 -47345
rect -5930 -48666 -5929 -47346
rect -4609 -48666 -4608 -47346
rect -5930 -48667 -4608 -48666
rect -4470 -47370 -4374 -47344
rect -3182 -47345 -3082 -47048
rect -4470 -48652 -4454 -47370
rect -4390 -48652 -4374 -47370
rect -5288 -48948 -5188 -48667
rect -4470 -48668 -4374 -48652
rect -3824 -47346 -2502 -47345
rect -3824 -48666 -3823 -47346
rect -2503 -48666 -2502 -47346
rect -3824 -48667 -2502 -48666
rect -2364 -47370 -2268 -47344
rect -1076 -47345 -976 -47048
rect -2364 -48652 -2348 -47370
rect -2284 -48652 -2268 -47370
rect -3182 -48948 -3082 -48667
rect -2364 -48668 -2268 -48652
rect -1718 -47346 -396 -47345
rect -1718 -48666 -1717 -47346
rect -397 -48666 -396 -47346
rect -1718 -48667 -396 -48666
rect -258 -47370 -162 -47344
rect 1030 -47345 1130 -47048
rect -258 -48652 -242 -47370
rect -178 -48652 -162 -47370
rect -1076 -48948 -976 -48667
rect -258 -48668 -162 -48652
rect 388 -47346 1710 -47345
rect 388 -48666 389 -47346
rect 1709 -48666 1710 -47346
rect 388 -48667 1710 -48666
rect 1848 -47370 1944 -47344
rect 3136 -47345 3236 -47048
rect 1848 -48652 1864 -47370
rect 1928 -48652 1944 -47370
rect 1030 -48948 1130 -48667
rect 1848 -48668 1944 -48652
rect 2494 -47346 3816 -47345
rect 2494 -48666 2495 -47346
rect 3815 -48666 3816 -47346
rect 2494 -48667 3816 -48666
rect 3954 -47370 4050 -47344
rect 5242 -47345 5342 -47048
rect 3954 -48652 3970 -47370
rect 4034 -48652 4050 -47370
rect 3136 -48948 3236 -48667
rect 3954 -48668 4050 -48652
rect 4600 -47346 5922 -47345
rect 4600 -48666 4601 -47346
rect 5921 -48666 5922 -47346
rect 4600 -48667 5922 -48666
rect 6060 -47370 6156 -47344
rect 7368 -47345 7468 -47048
rect 8160 -47344 8260 -47048
rect 6060 -48652 6076 -47370
rect 6140 -48652 6156 -47370
rect 5242 -48948 5342 -48667
rect 6060 -48668 6156 -48652
rect 6706 -47346 8028 -47345
rect 6706 -48666 6707 -47346
rect 8027 -47942 8028 -47346
rect 8160 -47370 8262 -47344
rect 8160 -47942 8182 -47370
rect 8027 -48042 8182 -47942
rect 8027 -48666 8028 -48042
rect 6706 -48667 8028 -48666
rect 8160 -48652 8182 -48042
rect 8246 -48652 8262 -47370
rect 7368 -48948 7468 -48667
rect 8160 -48668 8262 -48652
rect 8160 -48948 8260 -48668
rect -7394 -49048 8260 -48948
rect -7394 -49345 -7294 -49048
rect -8036 -49346 -6714 -49345
rect -8036 -50666 -8035 -49346
rect -6715 -50666 -6714 -49346
rect -8036 -50667 -6714 -50666
rect -6576 -49370 -6480 -49344
rect -5288 -49345 -5188 -49048
rect -6576 -50652 -6560 -49370
rect -6496 -50652 -6480 -49370
rect -7394 -51345 -7294 -50667
rect -6576 -50668 -6480 -50652
rect -5930 -49346 -4608 -49345
rect -5930 -50666 -5929 -49346
rect -4609 -50666 -4608 -49346
rect -5930 -50667 -4608 -50666
rect -4470 -49370 -4374 -49344
rect -3182 -49345 -3082 -49048
rect -4470 -50652 -4454 -49370
rect -4390 -50652 -4374 -49370
rect -5288 -50948 -5188 -50667
rect -4470 -50668 -4374 -50652
rect -3824 -49346 -2502 -49345
rect -3824 -50666 -3823 -49346
rect -2503 -50666 -2502 -49346
rect -3824 -50667 -2502 -50666
rect -2364 -49370 -2268 -49344
rect -1076 -49345 -976 -49048
rect -2364 -50652 -2348 -49370
rect -2284 -50652 -2268 -49370
rect -3182 -50948 -3082 -50667
rect -2364 -50668 -2268 -50652
rect -1718 -49346 -396 -49345
rect -1718 -50666 -1717 -49346
rect -397 -50666 -396 -49346
rect -1718 -50667 -396 -50666
rect -258 -49370 -162 -49344
rect 1030 -49345 1130 -49048
rect -258 -50652 -242 -49370
rect -178 -50652 -162 -49370
rect -1076 -50948 -976 -50667
rect -258 -50668 -162 -50652
rect 388 -49346 1710 -49345
rect 388 -50666 389 -49346
rect 1709 -50666 1710 -49346
rect 388 -50667 1710 -50666
rect 1848 -49370 1944 -49344
rect 3136 -49345 3236 -49048
rect 1848 -50652 1864 -49370
rect 1928 -50652 1944 -49370
rect 1030 -50948 1130 -50667
rect 1848 -50668 1944 -50652
rect 2494 -49346 3816 -49345
rect 2494 -50666 2495 -49346
rect 3815 -50666 3816 -49346
rect 2494 -50667 3816 -50666
rect 3954 -49370 4050 -49344
rect 5242 -49345 5342 -49048
rect 3954 -50652 3970 -49370
rect 4034 -50652 4050 -49370
rect 3136 -50948 3236 -50667
rect 3954 -50668 4050 -50652
rect 4600 -49346 5922 -49345
rect 4600 -50666 4601 -49346
rect 5921 -50666 5922 -49346
rect 4600 -50667 5922 -50666
rect 6060 -49370 6156 -49344
rect 7368 -49345 7468 -49048
rect 8160 -49344 8260 -49048
rect 6060 -50652 6076 -49370
rect 6140 -50652 6156 -49370
rect 5242 -50948 5342 -50667
rect 6060 -50668 6156 -50652
rect 6706 -49346 8028 -49345
rect 6706 -50666 6707 -49346
rect 8027 -49942 8028 -49346
rect 8160 -49370 8262 -49344
rect 8160 -49942 8182 -49370
rect 8027 -50042 8182 -49942
rect 8027 -50666 8028 -50042
rect 6706 -50667 8028 -50666
rect 8160 -50652 8182 -50042
rect 8246 -50652 8262 -49370
rect 7368 -50948 7468 -50667
rect 8160 -50668 8262 -50652
rect 8160 -50948 8260 -50668
rect -5288 -51048 8260 -50948
rect -8036 -51346 -6714 -51345
rect -8036 -52666 -8035 -51346
rect -6715 -52666 -6714 -51346
rect -8036 -52667 -6714 -52666
rect -6576 -51370 -6480 -51344
rect -5288 -51345 -5188 -51048
rect -6576 -52652 -6560 -51370
rect -6496 -52652 -6480 -51370
rect -7394 -53345 -7294 -52667
rect -6576 -52668 -6480 -52652
rect -5930 -51346 -4608 -51345
rect -5930 -52666 -5929 -51346
rect -4609 -52666 -4608 -51346
rect -5930 -52667 -4608 -52666
rect -4470 -51370 -4374 -51344
rect -3182 -51345 -3082 -51048
rect -4470 -52652 -4454 -51370
rect -4390 -52652 -4374 -51370
rect -5288 -52948 -5188 -52667
rect -4470 -52668 -4374 -52652
rect -3824 -51346 -2502 -51345
rect -3824 -52666 -3823 -51346
rect -2503 -52666 -2502 -51346
rect -3824 -52667 -2502 -52666
rect -2364 -51370 -2268 -51344
rect -1076 -51345 -976 -51048
rect -2364 -52652 -2348 -51370
rect -2284 -52652 -2268 -51370
rect -3182 -52948 -3082 -52667
rect -2364 -52668 -2268 -52652
rect -1718 -51346 -396 -51345
rect -1718 -52666 -1717 -51346
rect -397 -52666 -396 -51346
rect -1718 -52667 -396 -52666
rect -258 -51370 -162 -51344
rect 1030 -51345 1130 -51048
rect -258 -52652 -242 -51370
rect -178 -52652 -162 -51370
rect -1076 -52948 -976 -52667
rect -258 -52668 -162 -52652
rect 388 -51346 1710 -51345
rect 388 -52666 389 -51346
rect 1709 -52666 1710 -51346
rect 388 -52667 1710 -52666
rect 1848 -51370 1944 -51344
rect 3136 -51345 3236 -51048
rect 1848 -52652 1864 -51370
rect 1928 -52652 1944 -51370
rect 1030 -52948 1130 -52667
rect 1848 -52668 1944 -52652
rect 2494 -51346 3816 -51345
rect 2494 -52666 2495 -51346
rect 3815 -52666 3816 -51346
rect 2494 -52667 3816 -52666
rect 3954 -51370 4050 -51344
rect 5242 -51345 5342 -51048
rect 3954 -52652 3970 -51370
rect 4034 -52652 4050 -51370
rect 3136 -52948 3236 -52667
rect 3954 -52668 4050 -52652
rect 4600 -51346 5922 -51345
rect 4600 -52666 4601 -51346
rect 5921 -52666 5922 -51346
rect 4600 -52667 5922 -52666
rect 6060 -51370 6156 -51344
rect 7368 -51345 7468 -51048
rect 8160 -51344 8260 -51048
rect 6060 -52652 6076 -51370
rect 6140 -52652 6156 -51370
rect 5242 -52948 5342 -52667
rect 6060 -52668 6156 -52652
rect 6706 -51346 8028 -51345
rect 6706 -52666 6707 -51346
rect 8027 -51942 8028 -51346
rect 8160 -51370 8262 -51344
rect 8160 -51942 8182 -51370
rect 8027 -52042 8182 -51942
rect 8027 -52666 8028 -52042
rect 6706 -52667 8028 -52666
rect 8160 -52652 8182 -52042
rect 8246 -52652 8262 -51370
rect 7368 -52948 7468 -52667
rect 8160 -52668 8262 -52652
rect 8160 -52948 8260 -52668
rect -5288 -52949 8264 -52948
rect -5288 -53047 8165 -52949
rect 8263 -53047 8264 -52949
rect -5288 -53048 8264 -53047
rect -8036 -53346 -6714 -53345
rect -8036 -54666 -8035 -53346
rect -6715 -54666 -6714 -53346
rect -8036 -54667 -6714 -54666
rect -6576 -53370 -6480 -53344
rect -5288 -53345 -5188 -53048
rect -6576 -54652 -6560 -53370
rect -6496 -54652 -6480 -53370
rect -7394 -55345 -7294 -54667
rect -6576 -54668 -6480 -54652
rect -5930 -53346 -4608 -53345
rect -5930 -54666 -5929 -53346
rect -4609 -54666 -4608 -53346
rect -5930 -54667 -4608 -54666
rect -4470 -53370 -4374 -53344
rect -3182 -53345 -3082 -53048
rect -4470 -54652 -4454 -53370
rect -4390 -54652 -4374 -53370
rect -5288 -54948 -5188 -54667
rect -4470 -54668 -4374 -54652
rect -3824 -53346 -2502 -53345
rect -3824 -54666 -3823 -53346
rect -2503 -54666 -2502 -53346
rect -3824 -54667 -2502 -54666
rect -2364 -53370 -2268 -53344
rect -1076 -53345 -976 -53048
rect -2364 -54652 -2348 -53370
rect -2284 -54652 -2268 -53370
rect -3182 -54948 -3082 -54667
rect -2364 -54668 -2268 -54652
rect -1718 -53346 -396 -53345
rect -1718 -54666 -1717 -53346
rect -397 -54666 -396 -53346
rect -1718 -54667 -396 -54666
rect -258 -53370 -162 -53344
rect 1030 -53345 1130 -53048
rect -258 -54652 -242 -53370
rect -178 -54652 -162 -53370
rect -1076 -54948 -976 -54667
rect -258 -54668 -162 -54652
rect 388 -53346 1710 -53345
rect 388 -54666 389 -53346
rect 1709 -54666 1710 -53346
rect 388 -54667 1710 -54666
rect 1848 -53370 1944 -53344
rect 3136 -53345 3236 -53048
rect 1848 -54652 1864 -53370
rect 1928 -54652 1944 -53370
rect 1030 -54948 1130 -54667
rect 1848 -54668 1944 -54652
rect 2494 -53346 3816 -53345
rect 2494 -54666 2495 -53346
rect 3815 -54666 3816 -53346
rect 2494 -54667 3816 -54666
rect 3954 -53370 4050 -53344
rect 5242 -53345 5342 -53048
rect 3954 -54652 3970 -53370
rect 4034 -54652 4050 -53370
rect 3136 -54948 3236 -54667
rect 3954 -54668 4050 -54652
rect 4600 -53346 5922 -53345
rect 4600 -54666 4601 -53346
rect 5921 -54666 5922 -53346
rect 4600 -54667 5922 -54666
rect 6060 -53370 6156 -53344
rect 7368 -53345 7468 -53048
rect 8160 -53344 8260 -53048
rect 6060 -54652 6076 -53370
rect 6140 -54652 6156 -53370
rect 5242 -54948 5342 -54667
rect 6060 -54668 6156 -54652
rect 6706 -53346 8028 -53345
rect 6706 -54666 6707 -53346
rect 8027 -53942 8028 -53346
rect 8160 -53370 8262 -53344
rect 8160 -53942 8182 -53370
rect 8027 -54042 8182 -53942
rect 8027 -54666 8028 -54042
rect 6706 -54667 8028 -54666
rect 8160 -54652 8182 -54042
rect 8246 -54652 8262 -53370
rect 7368 -54948 7468 -54667
rect 8160 -54668 8262 -54652
rect 8160 -54948 8260 -54668
rect -5288 -54949 8262 -54948
rect -5288 -55047 8163 -54949
rect 8261 -55047 8262 -54949
rect -5288 -55048 8262 -55047
rect -8036 -55346 -6714 -55345
rect -8036 -56666 -8035 -55346
rect -6715 -56666 -6714 -55346
rect -8036 -56667 -6714 -56666
rect -6576 -55370 -6480 -55344
rect -5288 -55345 -5188 -55048
rect -6576 -56652 -6560 -55370
rect -6496 -56652 -6480 -55370
rect -7394 -57345 -7294 -56667
rect -6576 -56668 -6480 -56652
rect -5930 -55346 -4608 -55345
rect -5930 -56666 -5929 -55346
rect -4609 -56666 -4608 -55346
rect -5930 -56667 -4608 -56666
rect -4470 -55370 -4374 -55344
rect -3182 -55345 -3082 -55048
rect -4470 -56652 -4454 -55370
rect -4390 -56652 -4374 -55370
rect -5288 -56948 -5188 -56667
rect -4470 -56668 -4374 -56652
rect -3824 -55346 -2502 -55345
rect -3824 -56666 -3823 -55346
rect -2503 -56666 -2502 -55346
rect -3824 -56667 -2502 -56666
rect -2364 -55370 -2268 -55344
rect -1076 -55345 -976 -55048
rect -2364 -56652 -2348 -55370
rect -2284 -56652 -2268 -55370
rect -3182 -56948 -3082 -56667
rect -2364 -56668 -2268 -56652
rect -1718 -55346 -396 -55345
rect -1718 -56666 -1717 -55346
rect -397 -56666 -396 -55346
rect -1718 -56667 -396 -56666
rect -258 -55370 -162 -55344
rect 1030 -55345 1130 -55048
rect -258 -56652 -242 -55370
rect -178 -56652 -162 -55370
rect -1076 -56948 -976 -56667
rect -258 -56668 -162 -56652
rect 388 -55346 1710 -55345
rect 388 -56666 389 -55346
rect 1709 -56666 1710 -55346
rect 388 -56667 1710 -56666
rect 1848 -55370 1944 -55344
rect 3136 -55345 3236 -55048
rect 1848 -56652 1864 -55370
rect 1928 -56652 1944 -55370
rect 1030 -56948 1130 -56667
rect 1848 -56668 1944 -56652
rect 2494 -55346 3816 -55345
rect 2494 -56666 2495 -55346
rect 3815 -56666 3816 -55346
rect 2494 -56667 3816 -56666
rect 3954 -55370 4050 -55344
rect 5242 -55345 5342 -55048
rect 3954 -56652 3970 -55370
rect 4034 -56652 4050 -55370
rect 3136 -56948 3236 -56667
rect 3954 -56668 4050 -56652
rect 4600 -55346 5922 -55345
rect 4600 -56666 4601 -55346
rect 5921 -56666 5922 -55346
rect 4600 -56667 5922 -56666
rect 6060 -55370 6156 -55344
rect 7368 -55345 7468 -55048
rect 8160 -55344 8260 -55048
rect 6060 -56652 6076 -55370
rect 6140 -56652 6156 -55370
rect 5242 -56948 5342 -56667
rect 6060 -56668 6156 -56652
rect 6706 -55346 8028 -55345
rect 6706 -56666 6707 -55346
rect 8027 -55942 8028 -55346
rect 8160 -55370 8262 -55344
rect 8160 -55942 8182 -55370
rect 8027 -56042 8182 -55942
rect 8027 -56666 8028 -56042
rect 6706 -56667 8028 -56666
rect 8160 -56652 8182 -56042
rect 8246 -56652 8262 -55370
rect 7368 -56948 7468 -56667
rect 8160 -56668 8262 -56652
rect 8160 -56948 8260 -56668
rect -5288 -57048 8260 -56948
rect -8036 -57346 -6714 -57345
rect -8036 -58666 -8035 -57346
rect -6715 -58666 -6714 -57346
rect -8036 -58667 -6714 -58666
rect -6576 -57370 -6480 -57344
rect -5288 -57345 -5188 -57048
rect -6576 -58652 -6560 -57370
rect -6496 -58652 -6480 -57370
rect -7394 -59345 -7294 -58667
rect -6576 -58668 -6480 -58652
rect -5930 -57346 -4608 -57345
rect -5930 -58666 -5929 -57346
rect -4609 -58666 -4608 -57346
rect -5930 -58667 -4608 -58666
rect -4470 -57370 -4374 -57344
rect -3182 -57345 -3082 -57048
rect -4470 -58652 -4454 -57370
rect -4390 -58652 -4374 -57370
rect -5288 -58948 -5188 -58667
rect -4470 -58668 -4374 -58652
rect -3824 -57346 -2502 -57345
rect -3824 -58666 -3823 -57346
rect -2503 -58666 -2502 -57346
rect -3824 -58667 -2502 -58666
rect -2364 -57370 -2268 -57344
rect -1076 -57345 -976 -57048
rect -2364 -58652 -2348 -57370
rect -2284 -58652 -2268 -57370
rect -3182 -58948 -3082 -58667
rect -2364 -58668 -2268 -58652
rect -1718 -57346 -396 -57345
rect -1718 -58666 -1717 -57346
rect -397 -58666 -396 -57346
rect -1718 -58667 -396 -58666
rect -258 -57370 -162 -57344
rect 1030 -57345 1130 -57048
rect -258 -58652 -242 -57370
rect -178 -58652 -162 -57370
rect -1076 -58948 -976 -58667
rect -258 -58668 -162 -58652
rect 388 -57346 1710 -57345
rect 388 -58666 389 -57346
rect 1709 -58666 1710 -57346
rect 388 -58667 1710 -58666
rect 1848 -57370 1944 -57344
rect 3136 -57345 3236 -57048
rect 1848 -58652 1864 -57370
rect 1928 -58652 1944 -57370
rect 1030 -58948 1130 -58667
rect 1848 -58668 1944 -58652
rect 2494 -57346 3816 -57345
rect 2494 -58666 2495 -57346
rect 3815 -58666 3816 -57346
rect 2494 -58667 3816 -58666
rect 3954 -57370 4050 -57344
rect 5242 -57345 5342 -57048
rect 3954 -58652 3970 -57370
rect 4034 -58652 4050 -57370
rect 3136 -58948 3236 -58667
rect 3954 -58668 4050 -58652
rect 4600 -57346 5922 -57345
rect 4600 -58666 4601 -57346
rect 5921 -58666 5922 -57346
rect 4600 -58667 5922 -58666
rect 6060 -57370 6156 -57344
rect 7368 -57345 7468 -57048
rect 8160 -57344 8260 -57048
rect 6060 -58652 6076 -57370
rect 6140 -58652 6156 -57370
rect 5242 -58948 5342 -58667
rect 6060 -58668 6156 -58652
rect 6706 -57346 8028 -57345
rect 6706 -58666 6707 -57346
rect 8027 -57942 8028 -57346
rect 8160 -57370 8262 -57344
rect 8160 -57942 8182 -57370
rect 8027 -58042 8182 -57942
rect 8027 -58666 8028 -58042
rect 6706 -58667 8028 -58666
rect 8160 -58652 8182 -58042
rect 8246 -58652 8262 -57370
rect 7368 -58948 7468 -58667
rect 8160 -58668 8262 -58652
rect 11076 -58380 50444 -58378
rect 11076 -58404 51344 -58380
rect 11076 -58408 50568 -58404
rect 12110 -58454 50568 -58408
rect 12110 -58514 17372 -58454
rect 8160 -58948 8260 -58668
rect -5288 -59048 8260 -58948
rect -8036 -59346 -6714 -59345
rect -8036 -60666 -8035 -59346
rect -6715 -60666 -6714 -59346
rect -8036 -60667 -6714 -60666
rect -6576 -59370 -6480 -59344
rect -5288 -59345 -5188 -59048
rect -6576 -60652 -6560 -59370
rect -6496 -60652 -6480 -59370
rect -7394 -61345 -7294 -60667
rect -6576 -60668 -6480 -60652
rect -5930 -59346 -4608 -59345
rect -5930 -60666 -5929 -59346
rect -4609 -60666 -4608 -59346
rect -5930 -60667 -4608 -60666
rect -4470 -59370 -4374 -59344
rect -3182 -59345 -3082 -59048
rect -4470 -60652 -4454 -59370
rect -4390 -60652 -4374 -59370
rect -5288 -60968 -5188 -60667
rect -4470 -60668 -4374 -60652
rect -3824 -59346 -2502 -59345
rect -3824 -60666 -3823 -59346
rect -2503 -60666 -2502 -59346
rect -3824 -60667 -2502 -60666
rect -2364 -59370 -2268 -59344
rect -1076 -59345 -976 -59048
rect -2364 -60652 -2348 -59370
rect -2284 -60652 -2268 -59370
rect -3182 -60968 -3082 -60667
rect -2364 -60668 -2268 -60652
rect -1718 -59346 -396 -59345
rect -1718 -60666 -1717 -59346
rect -397 -60666 -396 -59346
rect -1718 -60667 -396 -60666
rect -258 -59370 -162 -59344
rect 1030 -59345 1130 -59048
rect -258 -60652 -242 -59370
rect -178 -60652 -162 -59370
rect -1076 -60968 -976 -60667
rect -258 -60668 -162 -60652
rect 388 -59346 1710 -59345
rect 388 -60666 389 -59346
rect 1709 -60666 1710 -59346
rect 388 -60667 1710 -60666
rect 1848 -59370 1944 -59344
rect 3136 -59345 3236 -59048
rect 1848 -60652 1864 -59370
rect 1928 -60652 1944 -59370
rect 1030 -60968 1130 -60667
rect 1848 -60668 1944 -60652
rect 2494 -59346 3816 -59345
rect 2494 -60666 2495 -59346
rect 3815 -60666 3816 -59346
rect 2494 -60667 3816 -60666
rect 3954 -59370 4050 -59344
rect 5242 -59345 5342 -59048
rect 3954 -60652 3970 -59370
rect 4034 -60652 4050 -59370
rect 3136 -60968 3236 -60667
rect 3954 -60668 4050 -60652
rect 4600 -59346 5922 -59345
rect 4600 -60666 4601 -59346
rect 5921 -60666 5922 -59346
rect 4600 -60667 5922 -60666
rect 6060 -59370 6156 -59344
rect 7368 -59345 7468 -59048
rect 8160 -59344 8260 -59048
rect 11076 -58608 17372 -58514
rect 49372 -58608 50568 -58454
rect 11076 -58794 50568 -58608
rect 11076 -59094 13228 -58794
rect 13828 -59094 49660 -58794
rect 50260 -59094 50568 -58794
rect 11076 -59156 50568 -59094
rect 51320 -59156 51344 -58404
rect 11076 -59178 51344 -59156
rect 49716 -59180 51344 -59178
rect 6060 -60652 6076 -59370
rect 6140 -60652 6156 -59370
rect 5242 -60968 5342 -60667
rect 6060 -60668 6156 -60652
rect 6706 -59346 8028 -59345
rect 6706 -60666 6707 -59346
rect 8027 -59942 8028 -59346
rect 8160 -59370 8262 -59344
rect 8160 -59942 8182 -59370
rect 8027 -60042 8182 -59942
rect 8027 -60666 8028 -60042
rect 6706 -60667 8028 -60666
rect 8160 -60652 8182 -60042
rect 8246 -60652 8262 -59370
rect 7368 -60968 7468 -60667
rect 8160 -60668 8262 -60652
rect 8160 -60968 8260 -60668
rect -5288 -61068 8260 -60968
rect -8036 -61346 -6714 -61345
rect -8036 -62666 -8035 -61346
rect -6715 -61930 -6714 -61346
rect -6576 -61370 -6480 -61344
rect -5288 -61345 -5188 -61068
rect -6576 -61930 -6560 -61370
rect -6715 -62030 -6560 -61930
rect -6715 -62666 -6714 -62030
rect -8036 -62667 -6714 -62666
rect -6576 -62652 -6560 -62030
rect -6496 -62652 -6480 -61370
rect -6576 -62668 -6480 -62652
rect -5930 -61346 -4608 -61345
rect -5930 -62666 -5929 -61346
rect -4609 -61930 -4608 -61346
rect -4470 -61370 -4374 -61344
rect -3182 -61345 -3082 -61068
rect -4470 -61930 -4454 -61370
rect -4609 -62030 -4454 -61930
rect -4609 -62666 -4608 -62030
rect -5930 -62667 -4608 -62666
rect -4470 -62652 -4454 -62030
rect -4390 -61930 -4374 -61370
rect -3824 -61346 -2502 -61345
rect -3824 -61930 -3823 -61346
rect -4390 -62030 -3823 -61930
rect -4390 -62652 -4374 -62030
rect -4470 -62668 -4374 -62652
rect -3824 -62666 -3823 -62030
rect -2503 -61930 -2502 -61346
rect -2364 -61370 -2268 -61344
rect -1076 -61345 -976 -61068
rect -2364 -61930 -2348 -61370
rect -2503 -62030 -2348 -61930
rect -2503 -62666 -2502 -62030
rect -3824 -62667 -2502 -62666
rect -2364 -62652 -2348 -62030
rect -2284 -61930 -2268 -61370
rect -1718 -61346 -396 -61345
rect -1718 -61930 -1717 -61346
rect -2284 -62030 -1717 -61930
rect -2284 -62652 -2268 -62030
rect -2364 -62668 -2268 -62652
rect -1718 -62666 -1717 -62030
rect -397 -61930 -396 -61346
rect -258 -61370 -162 -61344
rect 1030 -61345 1130 -61068
rect -258 -61930 -242 -61370
rect -397 -62030 -242 -61930
rect -397 -62666 -396 -62030
rect -1718 -62667 -396 -62666
rect -258 -62652 -242 -62030
rect -178 -61930 -162 -61370
rect 388 -61346 1710 -61345
rect 388 -61930 389 -61346
rect -178 -62030 389 -61930
rect -178 -62652 -162 -62030
rect -258 -62668 -162 -62652
rect 388 -62666 389 -62030
rect 1709 -61930 1710 -61346
rect 1848 -61370 1944 -61344
rect 3136 -61345 3236 -61068
rect 1848 -61930 1864 -61370
rect 1709 -62030 1864 -61930
rect 1709 -62666 1710 -62030
rect 388 -62667 1710 -62666
rect 1848 -62652 1864 -62030
rect 1928 -61930 1944 -61370
rect 2494 -61346 3816 -61345
rect 2494 -61930 2495 -61346
rect 1928 -62030 2495 -61930
rect 1928 -62652 1944 -62030
rect 1848 -62668 1944 -62652
rect 2494 -62666 2495 -62030
rect 3815 -61930 3816 -61346
rect 3954 -61370 4050 -61344
rect 5242 -61345 5342 -61068
rect 3954 -61930 3970 -61370
rect 3815 -62030 3970 -61930
rect 3815 -62666 3816 -62030
rect 2494 -62667 3816 -62666
rect 3954 -62652 3970 -62030
rect 4034 -61930 4050 -61370
rect 4600 -61346 5922 -61345
rect 4600 -61930 4601 -61346
rect 4034 -62030 4601 -61930
rect 4034 -62652 4050 -62030
rect 3954 -62668 4050 -62652
rect 4600 -62666 4601 -62030
rect 5921 -61930 5922 -61346
rect 6060 -61370 6156 -61344
rect 7368 -61345 7468 -61068
rect 8160 -61344 8260 -61068
rect 6060 -61930 6076 -61370
rect 5921 -62036 6076 -61930
rect 5921 -62666 5922 -62036
rect 4600 -62667 5922 -62666
rect 6060 -62652 6076 -62036
rect 6140 -61930 6156 -61370
rect 6706 -61346 8028 -61345
rect 6706 -61930 6707 -61346
rect 6140 -62036 6707 -61930
rect 6140 -62652 6156 -62036
rect 6060 -62668 6156 -62652
rect 6706 -62666 6707 -62036
rect 8027 -61936 8028 -61346
rect 8160 -61370 8262 -61344
rect 8160 -61936 8182 -61370
rect 8027 -62036 8182 -61936
rect 8027 -62666 8028 -62036
rect 8160 -62122 8182 -62036
rect 6706 -62667 8028 -62666
rect 8166 -62652 8182 -62122
rect 8246 -62652 8262 -61370
rect 8166 -62668 8262 -62652
rect -8282 -63023 -7828 -63022
rect -8282 -63121 -7927 -63023
rect -7829 -63121 -7828 -63023
rect -8282 -63122 -7828 -63121
rect -25201 -63278 -25099 -63277
rect -25201 -63378 -25200 -63278
rect -25100 -63378 -25099 -63278
rect -25201 -63379 -25099 -63378
rect -27764 -64532 7040 -64348
rect -27764 -64832 -27578 -64532
rect -26978 -64832 -26066 -64532
rect -25466 -64832 -23578 -64532
rect -22978 -64832 -22066 -64532
rect -21466 -64832 -19578 -64532
rect -18978 -64832 -18066 -64532
rect -17466 -64832 -15578 -64532
rect -14978 -64832 -14066 -64532
rect -13466 -64832 -11578 -64532
rect -10978 -64832 -10066 -64532
rect -9466 -64832 -7578 -64532
rect -6978 -64832 -6066 -64532
rect -5466 -64832 -3578 -64532
rect -2978 -64832 -2066 -64532
rect -1466 -64832 422 -64532
rect 1022 -64832 1934 -64532
rect 2534 -64832 4422 -64532
rect 5022 -64832 5934 -64532
rect 6534 -64832 7040 -64532
rect -27764 -65036 7040 -64832
rect 7728 -65036 8854 -64348
rect -27762 -65100 -27388 -65036
rect -25564 -65100 -25282 -65036
rect -27762 -65148 -25282 -65100
rect -23762 -65100 -23388 -65036
rect -21564 -65100 -21282 -65036
rect -23762 -65148 -21282 -65100
rect -19762 -65100 -19388 -65036
rect -17564 -65100 -17282 -65036
rect -19762 -65148 -17282 -65100
rect -15762 -65100 -15388 -65036
rect -13564 -65100 -13282 -65036
rect -15762 -65148 -13282 -65100
rect -11762 -65100 -11388 -65036
rect -9564 -65100 -9282 -65036
rect -11762 -65148 -9282 -65100
rect -7762 -65100 -7388 -65036
rect -5564 -65100 -5282 -65036
rect -7762 -65148 -5282 -65100
rect -3762 -65100 -3388 -65036
rect -1564 -65100 -1282 -65036
rect -3762 -65148 -1282 -65100
rect 238 -65100 612 -65036
rect 2436 -65100 2718 -65036
rect 238 -65148 2718 -65100
rect 4238 -65100 4612 -65036
rect 6436 -65100 6718 -65036
rect 4238 -65148 6718 -65100
rect -27762 -69154 -25282 -69088
rect -27762 -69222 -27430 -69154
rect -25722 -69222 -25282 -69154
rect -27762 -69404 -25282 -69222
rect -27762 -69704 -27578 -69404
rect -26978 -69704 -26066 -69404
rect -25466 -69704 -25282 -69404
rect -27762 -69716 -25282 -69704
rect -23762 -69154 -21282 -69088
rect -23762 -69222 -23430 -69154
rect -21722 -69222 -21282 -69154
rect -23762 -69404 -21282 -69222
rect -23762 -69704 -23578 -69404
rect -22978 -69704 -22066 -69404
rect -21466 -69704 -21282 -69404
rect -23762 -69716 -21282 -69704
rect -19762 -69154 -17282 -69088
rect -19762 -69222 -19430 -69154
rect -17722 -69222 -17282 -69154
rect -19762 -69404 -17282 -69222
rect -19762 -69704 -19578 -69404
rect -18978 -69704 -18066 -69404
rect -17466 -69704 -17282 -69404
rect -19762 -69716 -17282 -69704
rect -15762 -69154 -13282 -69088
rect -15762 -69222 -15430 -69154
rect -13722 -69222 -13282 -69154
rect -15762 -69404 -13282 -69222
rect -15762 -69704 -15578 -69404
rect -14978 -69704 -14066 -69404
rect -13466 -69704 -13282 -69404
rect -15762 -69716 -13282 -69704
rect -11762 -69154 -9282 -69088
rect -11762 -69222 -11430 -69154
rect -9722 -69222 -9282 -69154
rect -11762 -69404 -9282 -69222
rect -11762 -69704 -11578 -69404
rect -10978 -69704 -10066 -69404
rect -9466 -69704 -9282 -69404
rect -11762 -69716 -9282 -69704
rect -7762 -69154 -5282 -69088
rect -7762 -69222 -7430 -69154
rect -5722 -69222 -5282 -69154
rect -7762 -69404 -5282 -69222
rect -7762 -69704 -7578 -69404
rect -6978 -69704 -6066 -69404
rect -5466 -69704 -5282 -69404
rect -7762 -69716 -5282 -69704
rect -3762 -69154 -1282 -69088
rect -3762 -69222 -3430 -69154
rect -1722 -69222 -1282 -69154
rect -3762 -69404 -1282 -69222
rect -3762 -69704 -3578 -69404
rect -2978 -69704 -2066 -69404
rect -1466 -69704 -1282 -69404
rect -3762 -69716 -1282 -69704
rect 238 -69154 2718 -69088
rect 238 -69222 570 -69154
rect 2278 -69222 2718 -69154
rect 238 -69404 2718 -69222
rect 238 -69704 422 -69404
rect 1022 -69704 1934 -69404
rect 2534 -69704 2718 -69404
rect 238 -69716 2718 -69704
rect 4238 -69154 6718 -69088
rect 4238 -69222 4570 -69154
rect 6278 -69222 6718 -69154
rect 4238 -69404 6718 -69222
rect 4238 -69704 4422 -69404
rect 5022 -69704 5934 -69404
rect 6534 -69704 6718 -69404
rect 4238 -69716 6718 -69704
rect 9356 -69716 11076 -69714
rect -27762 -69738 11076 -69716
rect -27762 -70490 10300 -69738
rect 11052 -70490 11076 -69738
rect -27762 -70492 11076 -70490
rect -27762 -70792 -27578 -70492
rect -26978 -70792 -26066 -70492
rect -25466 -70516 -23578 -70492
rect -25466 -70792 -25282 -70516
rect -27762 -70974 -25282 -70792
rect -27762 -71042 -27430 -70974
rect -25722 -71042 -25282 -70974
rect -27762 -71108 -25282 -71042
rect -23762 -70792 -23578 -70516
rect -22978 -70792 -22066 -70492
rect -21466 -70516 -19578 -70492
rect -21466 -70792 -21282 -70516
rect -23762 -70974 -21282 -70792
rect -23762 -71042 -23430 -70974
rect -21722 -71042 -21282 -70974
rect -23762 -71108 -21282 -71042
rect -19762 -70792 -19578 -70516
rect -18978 -70792 -18066 -70492
rect -17466 -70516 -15578 -70492
rect -17466 -70792 -17282 -70516
rect -19762 -70974 -17282 -70792
rect -19762 -71042 -19430 -70974
rect -17722 -71042 -17282 -70974
rect -19762 -71108 -17282 -71042
rect -15762 -70792 -15578 -70516
rect -14978 -70792 -14066 -70492
rect -13466 -70516 -11578 -70492
rect -13466 -70792 -13282 -70516
rect -15762 -70974 -13282 -70792
rect -15762 -71042 -15430 -70974
rect -13722 -71042 -13282 -70974
rect -15762 -71108 -13282 -71042
rect -11762 -70792 -11578 -70516
rect -10978 -70792 -10066 -70492
rect -9466 -70516 -7578 -70492
rect -9466 -70792 -9282 -70516
rect -11762 -70974 -9282 -70792
rect -11762 -71042 -11430 -70974
rect -9722 -71042 -9282 -70974
rect -11762 -71108 -9282 -71042
rect -7762 -70792 -7578 -70516
rect -6978 -70792 -6066 -70492
rect -5466 -70516 -3578 -70492
rect -5466 -70792 -5282 -70516
rect -7762 -70974 -5282 -70792
rect -7762 -71042 -7430 -70974
rect -5722 -71042 -5282 -70974
rect -7762 -71108 -5282 -71042
rect -3762 -70792 -3578 -70516
rect -2978 -70792 -2066 -70492
rect -1466 -70516 422 -70492
rect -1466 -70792 -1282 -70516
rect -3762 -70974 -1282 -70792
rect -3762 -71042 -3430 -70974
rect -1722 -71042 -1282 -70974
rect -3762 -71108 -1282 -71042
rect 238 -70792 422 -70516
rect 1022 -70792 1934 -70492
rect 2534 -70516 4422 -70492
rect 2534 -70792 2718 -70516
rect 238 -70974 2718 -70792
rect 238 -71042 570 -70974
rect 2278 -71042 2718 -70974
rect 238 -71108 2718 -71042
rect 4238 -70792 4422 -70516
rect 5022 -70792 5934 -70492
rect 6534 -70514 11076 -70492
rect 6534 -70516 10276 -70514
rect 6534 -70792 6718 -70516
rect 4238 -70974 6718 -70792
rect 4238 -71042 4570 -70974
rect 6278 -71042 6718 -70974
rect 4238 -71108 6718 -71042
rect -27762 -75096 -25282 -75048
rect -27762 -75160 -27388 -75096
rect -25564 -75160 -25282 -75096
rect -23762 -75096 -21282 -75048
rect -23762 -75160 -23388 -75096
rect -21564 -75160 -21282 -75096
rect -19762 -75096 -17282 -75048
rect -19762 -75160 -19388 -75096
rect -17564 -75160 -17282 -75096
rect -15762 -75096 -13282 -75048
rect -15762 -75160 -15388 -75096
rect -13564 -75160 -13282 -75096
rect -11762 -75096 -9282 -75048
rect -11762 -75160 -11388 -75096
rect -9564 -75160 -9282 -75096
rect -7762 -75096 -5282 -75048
rect -7762 -75160 -7388 -75096
rect -5564 -75160 -5282 -75096
rect -3762 -75096 -1282 -75048
rect -3762 -75160 -3388 -75096
rect -1564 -75160 -1282 -75096
rect 238 -75096 2718 -75048
rect 238 -75160 612 -75096
rect 2436 -75160 2718 -75096
rect 4238 -75096 6718 -75048
rect 4238 -75160 4612 -75096
rect 6436 -75160 6718 -75096
rect -27762 -75178 7728 -75160
rect -27762 -75364 7064 -75178
rect -27762 -75664 -27578 -75364
rect -26978 -75664 -26066 -75364
rect -25466 -75664 -23578 -75364
rect -22978 -75664 -22066 -75364
rect -21466 -75664 -19578 -75364
rect -18978 -75664 -18066 -75364
rect -17466 -75664 -15578 -75364
rect -14978 -75664 -14066 -75364
rect -13466 -75664 -11578 -75364
rect -10978 -75664 -10066 -75364
rect -9466 -75664 -7578 -75364
rect -6978 -75664 -6066 -75364
rect -5466 -75664 -3578 -75364
rect -2978 -75664 -2066 -75364
rect -1466 -75664 422 -75364
rect 1022 -75664 1934 -75364
rect 2534 -75664 4422 -75364
rect 5022 -75664 5934 -75364
rect 6534 -75664 7064 -75364
rect -27762 -75818 7064 -75664
rect 7704 -75818 7728 -75178
rect -27762 -75848 7728 -75818
<< via4 >>
rect 8788 -28378 9588 -27578
rect 50552 -28378 51352 -27578
rect 10428 -29738 11124 -29048
rect 24470 -29736 25160 -29038
rect 50576 -39456 51328 -38704
rect 50544 -43984 51344 -43184
rect 9250 -56724 9554 -56598
rect 9250 -57518 9372 -56724
rect 9372 -57518 9436 -56724
rect 9436 -57518 9554 -56724
rect 9250 -57594 9554 -57518
rect 10276 -58408 11076 -58378
rect 10276 -58514 10294 -58408
rect 10294 -58514 11076 -58408
rect 10276 -59178 11076 -58514
rect 50568 -59156 51320 -58404
rect 7040 -65036 7728 -64348
rect 8854 -65036 9542 -64348
rect 10300 -70490 11052 -69738
rect 7064 -75818 7704 -75178
<< mimcap2 >>
rect 11462 -29442 17262 -28992
rect 11462 -29742 11512 -29442
rect 17212 -29742 17262 -29442
rect 11462 -29792 17262 -29742
rect 17862 -29442 23662 -28992
rect 17862 -29742 17912 -29442
rect 23612 -29742 23662 -29442
rect 17862 -29792 23662 -29742
rect 10376 -35924 10776 -30074
rect 10376 -36224 10426 -35924
rect 10726 -36224 10776 -35924
rect 12316 -35842 17116 -30992
rect 12316 -36142 12366 -35842
rect 17066 -36142 17116 -35842
rect 12316 -36192 17116 -36142
rect 17916 -35842 22716 -30992
rect 17916 -36142 17966 -35842
rect 22666 -36142 22716 -35842
rect 17916 -36192 22716 -36142
rect 24420 -35924 24820 -30074
rect 10376 -36274 10776 -36224
rect 24420 -36224 24470 -35924
rect 24770 -36224 24820 -35924
rect 24420 -36274 24820 -36224
rect 10376 -42416 10776 -36566
rect 12316 -41442 17116 -36592
rect 12316 -41742 12366 -41442
rect 17066 -41742 17116 -41442
rect 12316 -41792 17116 -41742
rect 17916 -41442 22716 -36592
rect 17916 -41742 17966 -41442
rect 22666 -41742 22716 -41442
rect 17916 -41792 22716 -41742
rect 10376 -42716 10426 -42416
rect 10726 -42716 10776 -42416
rect 10376 -42766 10776 -42716
rect 24420 -42416 24820 -36566
rect 24420 -42702 24470 -42416
rect 24770 -42702 24820 -42416
rect 24420 -42766 24820 -42702
rect 10962 -43442 16762 -42992
rect 10962 -43742 11012 -43442
rect 16712 -43742 16762 -43442
rect 10962 -43792 16762 -43742
rect 17362 -43442 23162 -42992
rect 17362 -43742 17412 -43442
rect 23112 -43742 23162 -43442
rect 17362 -43792 23162 -43742
<< mimcap2contact >>
rect 11512 -29742 17212 -29442
rect 17912 -29742 23612 -29442
rect 10426 -36224 10726 -35924
rect 12366 -36142 17066 -35842
rect 17966 -36142 22666 -35842
rect 24470 -36224 24770 -35924
rect 12366 -41742 17066 -41442
rect 17966 -41742 22666 -41442
rect 10426 -42716 10726 -42416
rect 24470 -42702 24770 -42416
rect 11012 -43742 16712 -43442
rect 17412 -43742 23112 -43442
<< metal5 >>
rect 8764 -27578 9612 -27554
rect 8764 -28378 8788 -27578
rect 9588 -28378 9612 -27578
rect 8764 -28402 9612 -28378
rect 50528 -27578 51376 -27554
rect 50528 -28378 50552 -27578
rect 51352 -28378 51376 -27578
rect 50528 -28402 51376 -28378
rect 8788 -56598 9588 -28402
rect 10276 -29038 25316 -28892
rect 10276 -29048 24470 -29038
rect 10276 -29738 10428 -29048
rect 11124 -29442 24470 -29048
rect 11124 -29738 11512 -29442
rect 10276 -29742 11512 -29738
rect 17212 -29742 17912 -29442
rect 23612 -29736 24470 -29442
rect 25160 -29736 25316 -29038
rect 23612 -29742 25316 -29736
rect 10276 -35842 25316 -29742
rect 10276 -35924 12366 -35842
rect 10276 -36224 10426 -35924
rect 10726 -36142 12366 -35924
rect 17066 -36142 17966 -35842
rect 22666 -35924 25316 -35842
rect 22666 -36142 24470 -35924
rect 10726 -36224 24470 -36142
rect 24770 -36224 25316 -35924
rect 10276 -41442 25316 -36224
rect 50552 -38704 51352 -28402
rect 50552 -39456 50576 -38704
rect 51328 -39456 51352 -38704
rect 50552 -39480 51352 -39456
rect 10276 -41742 12366 -41442
rect 17066 -41742 17966 -41442
rect 22666 -41742 25316 -41442
rect 10276 -42416 25316 -41742
rect 10276 -42716 10426 -42416
rect 10726 -42702 24470 -42416
rect 24770 -42702 25316 -42416
rect 10726 -42716 25316 -42702
rect 10276 -42742 25316 -42716
rect 10276 -43442 25314 -42742
rect 10276 -43742 11012 -43442
rect 16712 -43742 17412 -43442
rect 23112 -43742 25314 -43442
rect 10276 -43894 25314 -43742
rect 50520 -43184 51368 -43160
rect 50520 -43984 50544 -43184
rect 51344 -43984 51368 -43184
rect 50520 -44008 51368 -43984
rect 8788 -57594 9250 -56598
rect 9554 -57594 9588 -56598
rect 7016 -64348 7752 -64324
rect 7016 -65036 7040 -64348
rect 7728 -65036 7752 -64348
rect 7016 -65060 7752 -65036
rect 8788 -64348 9588 -57594
rect 10252 -58378 11100 -58354
rect 10252 -59178 10276 -58378
rect 11076 -59178 11100 -58378
rect 10252 -59202 11100 -59178
rect 50544 -58404 51344 -44008
rect 50544 -59156 50568 -58404
rect 51320 -59156 51344 -58404
rect 50544 -59180 51344 -59156
rect 8788 -65036 8854 -64348
rect 9542 -65036 9588 -64348
rect 7040 -75178 7728 -65060
rect 8788 -65088 9588 -65036
rect 10276 -69738 11076 -59202
rect 10276 -70490 10300 -69738
rect 11052 -70490 11076 -69738
rect 10276 -70514 11076 -70490
rect 7040 -75818 7064 -75178
rect 7704 -75818 7728 -75178
rect 7040 -75842 7728 -75818
<< labels >>
flabel metal3 -18928 -63224 -18910 -63206 1 FreeSans 480 0 0 0 c6m
flabel metal3 -16804 -63244 -16796 -63228 1 FreeSans 480 0 0 0 c5m
flabel metal3 -14718 -63246 -14704 -63230 1 FreeSans 480 0 0 0 c4m
flabel metal3 -8458 -63254 -8442 -63236 1 FreeSans 480 0 0 0 c1m
flabel metal3 -9900 -63276 -9878 -63242 1 FreeSans 480 0 0 0 cdumm
flabel metal3 -7508 -63088 -7478 -63062 1 FreeSans 480 0 0 0 c0m
flabel metal4 -27544 -70138 -27514 -70094 1 FreeSans 480 0 0 0 VSS
port 3 n ground bidirectional
flabel metal4 -27740 -64374 -27728 -64364 1 FreeSans 480 0 0 0 VDD
port 2 n power bidirectional
flabel metal3 -28160 -74900 -28146 -74892 1 FreeSans 480 0 0 0 vref
port 5 n
flabel metal3 -28452 -72922 -28438 -72906 1 FreeSans 480 0 0 0 vlow
port 4 n
flabel metal3 -28232 -67966 -28214 -67946 1 FreeSans 480 0 0 0 vin
port 6 n
flabel metal3 12544 -58056 12562 -58044 1 FreeSans 480 0 0 0 sample
port 1 n
flabel metal2 12200 -57048 12212 -57040 1 FreeSans 480 0 0 0 adc_run
flabel metal1 -28342 -72610 -28336 -72600 1 FreeSans 480 0 0 0 q7
port 7 n
flabel metal1 -24328 -72616 -24316 -72604 1 FreeSans 480 0 0 0 q6
port 8 n
flabel metal1 -20346 -72616 -20340 -72608 1 FreeSans 480 0 0 0 q5
port 9 n
flabel metal1 -16352 -72620 -16346 -72608 1 FreeSans 480 0 0 0 q4
port 10 n
flabel metal1 -12382 -72614 -12370 -72604 1 FreeSans 480 0 0 0 q3
port 11 n
flabel metal1 -8362 -72620 -8352 -72608 1 FreeSans 480 0 0 0 q2
port 12 n
flabel metal1 -356 -72608 -350 -72602 1 FreeSans 480 0 0 0 q1
port 13 n
flabel metal1 3634 -72616 3644 -72606 1 FreeSans 480 0 0 0 q0
port 14 n
flabel metal1 15262 -56936 15270 -56922 1 FreeSans 480 0 0 0 ibiasn
port 15 n
flabel metal3 10682 -52044 10722 -52028 1 FreeSans 480 0 0 0 vcom
port 20 n
flabel metal2 27012 -43058 27020 -43048 1 FreeSans 480 0 0 0 vcom_buf
flabel metal2 52036 -40050 52042 -40042 1 FreeSans 480 0 0 0 ibiasp
port 16 n
flabel metal2 52026 -42516 52034 -42508 1 FreeSans 480 0 0 0 adc_clk
port 17 n
flabel metal2 58410 -41968 58422 -41960 1 FreeSans 480 0 0 0 comp_out
port 18 n
flabel metal2 58400 -42168 58406 -42162 1 FreeSans 480 0 0 0 comp_outm
port 19 n
flabel metal3 -25158 -63656 -25132 -63634 1 FreeSans 480 0 0 0 c7m
flabel metal3 -12584 -63246 -12564 -63222 1 FreeSans 480 0 0 0 c2m
flabel metal3 -10558 -63254 -10540 -63232 1 FreeSans 480 0 0 0 c3m
flabel metal1 -28148 -72606 -28142 -72602 5 FreeSans 480 0 0 0 amux_2to1_17/SEL
flabel metal2 -26552 -72536 -26544 -72528 5 FreeSans 480 0 0 0 amux_2to1_17/A
flabel metal2 -26298 -72554 -26290 -72548 5 FreeSans 480 0 0 0 amux_2to1_17/Y
flabel metal2 -27074 -72556 -27064 -72550 5 FreeSans 480 0 0 0 amux_2to1_17/B
flabel metal2 -27688 -72560 -27678 -72550 5 FreeSans 480 0 0 0 amux_2to1_17/SELB
flabel metal4 -26812 -75832 -26800 -75822 5 FreeSans 480 0 0 0 amux_2to1_17/VDD
flabel metal4 -26740 -70332 -26726 -70324 5 FreeSans 480 0 0 0 amux_2to1_17/VSS
flabel locali -27908 -72693 -27874 -72659 0 FreeSans 340 0 0 0 amux_2to1_17/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -27908 -72625 -27874 -72591 0 FreeSans 340 0 0 0 amux_2to1_17/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -28000 -72625 -27966 -72591 0 FreeSans 340 0 0 0 amux_2to1_17/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -28043 -72931 -28009 -72897 0 FreeSans 200 0 0 0 amux_2to1_17/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -28043 -72387 -28009 -72353 0 FreeSans 200 0 0 0 amux_2to1_17/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -28043 -72387 -28009 -72353 0 FreeSans 200 0 0 0 amux_2to1_17/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -28043 -72931 -28009 -72897 0 FreeSans 200 0 0 0 amux_2to1_17/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -28072 -72370 -28072 -72370 2 amux_2to1_17/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -24148 -72606 -24142 -72602 5 FreeSans 480 0 0 0 amux_2to1_16/SEL
flabel metal2 -22552 -72536 -22544 -72528 5 FreeSans 480 0 0 0 amux_2to1_16/A
flabel metal2 -22298 -72554 -22290 -72548 5 FreeSans 480 0 0 0 amux_2to1_16/Y
flabel metal2 -23074 -72556 -23064 -72550 5 FreeSans 480 0 0 0 amux_2to1_16/B
flabel metal2 -23688 -72560 -23678 -72550 5 FreeSans 480 0 0 0 amux_2to1_16/SELB
flabel metal4 -22812 -75832 -22800 -75822 5 FreeSans 480 0 0 0 amux_2to1_16/VDD
flabel metal4 -22740 -70332 -22726 -70324 5 FreeSans 480 0 0 0 amux_2to1_16/VSS
flabel locali -23908 -72693 -23874 -72659 0 FreeSans 340 0 0 0 amux_2to1_16/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -23908 -72625 -23874 -72591 0 FreeSans 340 0 0 0 amux_2to1_16/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -24000 -72625 -23966 -72591 0 FreeSans 340 0 0 0 amux_2to1_16/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -24043 -72931 -24009 -72897 0 FreeSans 200 0 0 0 amux_2to1_16/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -24043 -72387 -24009 -72353 0 FreeSans 200 0 0 0 amux_2to1_16/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -24043 -72387 -24009 -72353 0 FreeSans 200 0 0 0 amux_2to1_16/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -24043 -72931 -24009 -72897 0 FreeSans 200 0 0 0 amux_2to1_16/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -24072 -72370 -24072 -72370 2 amux_2to1_16/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -20148 -72606 -20142 -72602 5 FreeSans 480 0 0 0 amux_2to1_15/SEL
flabel metal2 -18552 -72536 -18544 -72528 5 FreeSans 480 0 0 0 amux_2to1_15/A
flabel metal2 -18298 -72554 -18290 -72548 5 FreeSans 480 0 0 0 amux_2to1_15/Y
flabel metal2 -19074 -72556 -19064 -72550 5 FreeSans 480 0 0 0 amux_2to1_15/B
flabel metal2 -19688 -72560 -19678 -72550 5 FreeSans 480 0 0 0 amux_2to1_15/SELB
flabel metal4 -18812 -75832 -18800 -75822 5 FreeSans 480 0 0 0 amux_2to1_15/VDD
flabel metal4 -18740 -70332 -18726 -70324 5 FreeSans 480 0 0 0 amux_2to1_15/VSS
flabel locali -19908 -72693 -19874 -72659 0 FreeSans 340 0 0 0 amux_2to1_15/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -19908 -72625 -19874 -72591 0 FreeSans 340 0 0 0 amux_2to1_15/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -20000 -72625 -19966 -72591 0 FreeSans 340 0 0 0 amux_2to1_15/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -20043 -72931 -20009 -72897 0 FreeSans 200 0 0 0 amux_2to1_15/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -20043 -72387 -20009 -72353 0 FreeSans 200 0 0 0 amux_2to1_15/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -20043 -72387 -20009 -72353 0 FreeSans 200 0 0 0 amux_2to1_15/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -20043 -72931 -20009 -72897 0 FreeSans 200 0 0 0 amux_2to1_15/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -20072 -72370 -20072 -72370 2 amux_2to1_15/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -16148 -72606 -16142 -72602 5 FreeSans 480 0 0 0 amux_2to1_14/SEL
flabel metal2 -14552 -72536 -14544 -72528 5 FreeSans 480 0 0 0 amux_2to1_14/A
flabel metal2 -14298 -72554 -14290 -72548 5 FreeSans 480 0 0 0 amux_2to1_14/Y
flabel metal2 -15074 -72556 -15064 -72550 5 FreeSans 480 0 0 0 amux_2to1_14/B
flabel metal2 -15688 -72560 -15678 -72550 5 FreeSans 480 0 0 0 amux_2to1_14/SELB
flabel metal4 -14812 -75832 -14800 -75822 5 FreeSans 480 0 0 0 amux_2to1_14/VDD
flabel metal4 -14740 -70332 -14726 -70324 5 FreeSans 480 0 0 0 amux_2to1_14/VSS
flabel locali -15908 -72693 -15874 -72659 0 FreeSans 340 0 0 0 amux_2to1_14/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -15908 -72625 -15874 -72591 0 FreeSans 340 0 0 0 amux_2to1_14/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -16000 -72625 -15966 -72591 0 FreeSans 340 0 0 0 amux_2to1_14/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -16043 -72931 -16009 -72897 0 FreeSans 200 0 0 0 amux_2to1_14/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -16043 -72387 -16009 -72353 0 FreeSans 200 0 0 0 amux_2to1_14/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -16043 -72387 -16009 -72353 0 FreeSans 200 0 0 0 amux_2to1_14/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -16043 -72931 -16009 -72897 0 FreeSans 200 0 0 0 amux_2to1_14/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -16072 -72370 -16072 -72370 2 amux_2to1_14/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -12148 -72606 -12142 -72602 5 FreeSans 480 0 0 0 amux_2to1_13/SEL
flabel metal2 -10552 -72536 -10544 -72528 5 FreeSans 480 0 0 0 amux_2to1_13/A
flabel metal2 -10298 -72554 -10290 -72548 5 FreeSans 480 0 0 0 amux_2to1_13/Y
flabel metal2 -11074 -72556 -11064 -72550 5 FreeSans 480 0 0 0 amux_2to1_13/B
flabel metal2 -11688 -72560 -11678 -72550 5 FreeSans 480 0 0 0 amux_2to1_13/SELB
flabel metal4 -10812 -75832 -10800 -75822 5 FreeSans 480 0 0 0 amux_2to1_13/VDD
flabel metal4 -10740 -70332 -10726 -70324 5 FreeSans 480 0 0 0 amux_2to1_13/VSS
flabel locali -11908 -72693 -11874 -72659 0 FreeSans 340 0 0 0 amux_2to1_13/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -11908 -72625 -11874 -72591 0 FreeSans 340 0 0 0 amux_2to1_13/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -12000 -72625 -11966 -72591 0 FreeSans 340 0 0 0 amux_2to1_13/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -12043 -72931 -12009 -72897 0 FreeSans 200 0 0 0 amux_2to1_13/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -12043 -72387 -12009 -72353 0 FreeSans 200 0 0 0 amux_2to1_13/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -12043 -72387 -12009 -72353 0 FreeSans 200 0 0 0 amux_2to1_13/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -12043 -72931 -12009 -72897 0 FreeSans 200 0 0 0 amux_2to1_13/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -12072 -72370 -12072 -72370 2 amux_2to1_13/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -8148 -72606 -8142 -72602 5 FreeSans 480 0 0 0 amux_2to1_12/SEL
flabel metal2 -6552 -72536 -6544 -72528 5 FreeSans 480 0 0 0 amux_2to1_12/A
flabel metal2 -6298 -72554 -6290 -72548 5 FreeSans 480 0 0 0 amux_2to1_12/Y
flabel metal2 -7074 -72556 -7064 -72550 5 FreeSans 480 0 0 0 amux_2to1_12/B
flabel metal2 -7688 -72560 -7678 -72550 5 FreeSans 480 0 0 0 amux_2to1_12/SELB
flabel metal4 -6812 -75832 -6800 -75822 5 FreeSans 480 0 0 0 amux_2to1_12/VDD
flabel metal4 -6740 -70332 -6726 -70324 5 FreeSans 480 0 0 0 amux_2to1_12/VSS
flabel locali -7908 -72693 -7874 -72659 0 FreeSans 340 0 0 0 amux_2to1_12/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -7908 -72625 -7874 -72591 0 FreeSans 340 0 0 0 amux_2to1_12/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -8000 -72625 -7966 -72591 0 FreeSans 340 0 0 0 amux_2to1_12/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -8043 -72931 -8009 -72897 0 FreeSans 200 0 0 0 amux_2to1_12/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -8043 -72387 -8009 -72353 0 FreeSans 200 0 0 0 amux_2to1_12/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -8043 -72387 -8009 -72353 0 FreeSans 200 0 0 0 amux_2to1_12/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -8043 -72931 -8009 -72897 0 FreeSans 200 0 0 0 amux_2to1_12/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -8072 -72370 -8072 -72370 2 amux_2to1_12/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -4148 -72606 -4142 -72602 5 FreeSans 480 0 0 0 amux_2to1_11/SEL
flabel metal2 -2552 -72536 -2544 -72528 5 FreeSans 480 0 0 0 amux_2to1_11/A
flabel metal2 -2298 -72554 -2290 -72548 5 FreeSans 480 0 0 0 amux_2to1_11/Y
flabel metal2 -3074 -72556 -3064 -72550 5 FreeSans 480 0 0 0 amux_2to1_11/B
flabel metal2 -3688 -72560 -3678 -72550 5 FreeSans 480 0 0 0 amux_2to1_11/SELB
flabel metal4 -2812 -75832 -2800 -75822 5 FreeSans 480 0 0 0 amux_2to1_11/VDD
flabel metal4 -2740 -70332 -2726 -70324 5 FreeSans 480 0 0 0 amux_2to1_11/VSS
flabel locali -3908 -72693 -3874 -72659 0 FreeSans 340 0 0 0 amux_2to1_11/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -3908 -72625 -3874 -72591 0 FreeSans 340 0 0 0 amux_2to1_11/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -4000 -72625 -3966 -72591 0 FreeSans 340 0 0 0 amux_2to1_11/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -4043 -72931 -4009 -72897 0 FreeSans 200 0 0 0 amux_2to1_11/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -4043 -72387 -4009 -72353 0 FreeSans 200 0 0 0 amux_2to1_11/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -4043 -72387 -4009 -72353 0 FreeSans 200 0 0 0 amux_2to1_11/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -4043 -72931 -4009 -72897 0 FreeSans 200 0 0 0 amux_2to1_11/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -4072 -72370 -4072 -72370 2 amux_2to1_11/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -148 -72606 -142 -72602 5 FreeSans 480 0 0 0 amux_2to1_10/SEL
flabel metal2 1448 -72536 1456 -72528 5 FreeSans 480 0 0 0 amux_2to1_10/A
flabel metal2 1702 -72554 1710 -72548 5 FreeSans 480 0 0 0 amux_2to1_10/Y
flabel metal2 926 -72556 936 -72550 5 FreeSans 480 0 0 0 amux_2to1_10/B
flabel metal2 312 -72560 322 -72550 5 FreeSans 480 0 0 0 amux_2to1_10/SELB
flabel metal4 1188 -75832 1200 -75822 5 FreeSans 480 0 0 0 amux_2to1_10/VDD
flabel metal4 1260 -70332 1274 -70324 5 FreeSans 480 0 0 0 amux_2to1_10/VSS
flabel locali 92 -72693 126 -72659 0 FreeSans 340 0 0 0 amux_2to1_10/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 92 -72625 126 -72591 0 FreeSans 340 0 0 0 amux_2to1_10/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 0 -72625 34 -72591 0 FreeSans 340 0 0 0 amux_2to1_10/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -43 -72931 -9 -72897 0 FreeSans 200 0 0 0 amux_2to1_10/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -43 -72387 -9 -72353 0 FreeSans 200 0 0 0 amux_2to1_10/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -43 -72387 -9 -72353 0 FreeSans 200 0 0 0 amux_2to1_10/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -43 -72931 -9 -72897 0 FreeSans 200 0 0 0 amux_2to1_10/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -72 -72370 -72 -72370 2 amux_2to1_10/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 3852 -72606 3858 -72602 5 FreeSans 480 0 0 0 amux_2to1_9/SEL
flabel metal2 5448 -72536 5456 -72528 5 FreeSans 480 0 0 0 amux_2to1_9/A
flabel metal2 5702 -72554 5710 -72548 5 FreeSans 480 0 0 0 amux_2to1_9/Y
flabel metal2 4926 -72556 4936 -72550 5 FreeSans 480 0 0 0 amux_2to1_9/B
flabel metal2 4312 -72560 4322 -72550 5 FreeSans 480 0 0 0 amux_2to1_9/SELB
flabel metal4 5188 -75832 5200 -75822 5 FreeSans 480 0 0 0 amux_2to1_9/VDD
flabel metal4 5260 -70332 5274 -70324 5 FreeSans 480 0 0 0 amux_2to1_9/VSS
flabel locali 4092 -72693 4126 -72659 0 FreeSans 340 0 0 0 amux_2to1_9/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 4092 -72625 4126 -72591 0 FreeSans 340 0 0 0 amux_2to1_9/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 4000 -72625 4034 -72591 0 FreeSans 340 0 0 0 amux_2to1_9/sky130_fd_sc_hd__inv_1_0/A
flabel nwell 3957 -72931 3991 -72897 0 FreeSans 200 0 0 0 amux_2to1_9/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 3957 -72387 3991 -72353 0 FreeSans 200 0 0 0 amux_2to1_9/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 3957 -72387 3991 -72353 0 FreeSans 200 0 0 0 amux_2to1_9/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 3957 -72931 3991 -72897 0 FreeSans 200 0 0 0 amux_2to1_9/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 3928 -72370 3928 -72370 2 amux_2to1_9/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -28148 -67594 -28142 -67590 1 FreeSans 480 0 0 0 amux_2to1_0/SEL
flabel metal2 -26552 -67668 -26544 -67660 1 FreeSans 480 0 0 0 amux_2to1_0/A
flabel metal2 -26298 -67648 -26290 -67642 1 FreeSans 480 0 0 0 amux_2to1_0/Y
flabel metal2 -27074 -67646 -27064 -67640 1 FreeSans 480 0 0 0 amux_2to1_0/B
flabel metal2 -27688 -67646 -27678 -67636 1 FreeSans 480 0 0 0 amux_2to1_0/SELB
flabel metal4 -26812 -64374 -26800 -64364 1 FreeSans 480 0 0 0 amux_2to1_0/VDD
flabel metal4 -26740 -69872 -26726 -69864 1 FreeSans 480 0 0 0 amux_2to1_0/VSS
flabel locali -27908 -67537 -27874 -67503 0 FreeSans 340 0 0 0 amux_2to1_0/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -27908 -67605 -27874 -67571 0 FreeSans 340 0 0 0 amux_2to1_0/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -28000 -67605 -27966 -67571 0 FreeSans 340 0 0 0 amux_2to1_0/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -28043 -67299 -28009 -67265 0 FreeSans 200 0 0 0 amux_2to1_0/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -28043 -67843 -28009 -67809 0 FreeSans 200 0 0 0 amux_2to1_0/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -28043 -67843 -28009 -67809 0 FreeSans 200 0 0 0 amux_2to1_0/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -28043 -67299 -28009 -67265 0 FreeSans 200 0 0 0 amux_2to1_0/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -28072 -67826 -28072 -67826 4 amux_2to1_0/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -24148 -67594 -24142 -67590 1 FreeSans 480 0 0 0 amux_2to1_1/SEL
flabel metal2 -22552 -67668 -22544 -67660 1 FreeSans 480 0 0 0 amux_2to1_1/A
flabel metal2 -22298 -67648 -22290 -67642 1 FreeSans 480 0 0 0 amux_2to1_1/Y
flabel metal2 -23074 -67646 -23064 -67640 1 FreeSans 480 0 0 0 amux_2to1_1/B
flabel metal2 -23688 -67646 -23678 -67636 1 FreeSans 480 0 0 0 amux_2to1_1/SELB
flabel metal4 -22812 -64374 -22800 -64364 1 FreeSans 480 0 0 0 amux_2to1_1/VDD
flabel metal4 -22740 -69872 -22726 -69864 1 FreeSans 480 0 0 0 amux_2to1_1/VSS
flabel locali -23908 -67537 -23874 -67503 0 FreeSans 340 0 0 0 amux_2to1_1/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -23908 -67605 -23874 -67571 0 FreeSans 340 0 0 0 amux_2to1_1/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -24000 -67605 -23966 -67571 0 FreeSans 340 0 0 0 amux_2to1_1/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -24043 -67299 -24009 -67265 0 FreeSans 200 0 0 0 amux_2to1_1/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -24043 -67843 -24009 -67809 0 FreeSans 200 0 0 0 amux_2to1_1/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -24043 -67843 -24009 -67809 0 FreeSans 200 0 0 0 amux_2to1_1/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -24043 -67299 -24009 -67265 0 FreeSans 200 0 0 0 amux_2to1_1/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -24072 -67826 -24072 -67826 4 amux_2to1_1/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -20148 -67594 -20142 -67590 1 FreeSans 480 0 0 0 amux_2to1_2/SEL
flabel metal2 -18552 -67668 -18544 -67660 1 FreeSans 480 0 0 0 amux_2to1_2/A
flabel metal2 -18298 -67648 -18290 -67642 1 FreeSans 480 0 0 0 amux_2to1_2/Y
flabel metal2 -19074 -67646 -19064 -67640 1 FreeSans 480 0 0 0 amux_2to1_2/B
flabel metal2 -19688 -67646 -19678 -67636 1 FreeSans 480 0 0 0 amux_2to1_2/SELB
flabel metal4 -18812 -64374 -18800 -64364 1 FreeSans 480 0 0 0 amux_2to1_2/VDD
flabel metal4 -18740 -69872 -18726 -69864 1 FreeSans 480 0 0 0 amux_2to1_2/VSS
flabel locali -19908 -67537 -19874 -67503 0 FreeSans 340 0 0 0 amux_2to1_2/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -19908 -67605 -19874 -67571 0 FreeSans 340 0 0 0 amux_2to1_2/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -20000 -67605 -19966 -67571 0 FreeSans 340 0 0 0 amux_2to1_2/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -20043 -67299 -20009 -67265 0 FreeSans 200 0 0 0 amux_2to1_2/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -20043 -67843 -20009 -67809 0 FreeSans 200 0 0 0 amux_2to1_2/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -20043 -67843 -20009 -67809 0 FreeSans 200 0 0 0 amux_2to1_2/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -20043 -67299 -20009 -67265 0 FreeSans 200 0 0 0 amux_2to1_2/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -20072 -67826 -20072 -67826 4 amux_2to1_2/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -16148 -67594 -16142 -67590 1 FreeSans 480 0 0 0 amux_2to1_3/SEL
flabel metal2 -14552 -67668 -14544 -67660 1 FreeSans 480 0 0 0 amux_2to1_3/A
flabel metal2 -14298 -67648 -14290 -67642 1 FreeSans 480 0 0 0 amux_2to1_3/Y
flabel metal2 -15074 -67646 -15064 -67640 1 FreeSans 480 0 0 0 amux_2to1_3/B
flabel metal2 -15688 -67646 -15678 -67636 1 FreeSans 480 0 0 0 amux_2to1_3/SELB
flabel metal4 -14812 -64374 -14800 -64364 1 FreeSans 480 0 0 0 amux_2to1_3/VDD
flabel metal4 -14740 -69872 -14726 -69864 1 FreeSans 480 0 0 0 amux_2to1_3/VSS
flabel locali -15908 -67537 -15874 -67503 0 FreeSans 340 0 0 0 amux_2to1_3/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -15908 -67605 -15874 -67571 0 FreeSans 340 0 0 0 amux_2to1_3/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -16000 -67605 -15966 -67571 0 FreeSans 340 0 0 0 amux_2to1_3/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -16043 -67299 -16009 -67265 0 FreeSans 200 0 0 0 amux_2to1_3/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -16043 -67843 -16009 -67809 0 FreeSans 200 0 0 0 amux_2to1_3/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -16043 -67843 -16009 -67809 0 FreeSans 200 0 0 0 amux_2to1_3/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -16043 -67299 -16009 -67265 0 FreeSans 200 0 0 0 amux_2to1_3/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -16072 -67826 -16072 -67826 4 amux_2to1_3/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -12148 -67594 -12142 -67590 1 FreeSans 480 0 0 0 amux_2to1_4/SEL
flabel metal2 -10552 -67668 -10544 -67660 1 FreeSans 480 0 0 0 amux_2to1_4/A
flabel metal2 -10298 -67648 -10290 -67642 1 FreeSans 480 0 0 0 amux_2to1_4/Y
flabel metal2 -11074 -67646 -11064 -67640 1 FreeSans 480 0 0 0 amux_2to1_4/B
flabel metal2 -11688 -67646 -11678 -67636 1 FreeSans 480 0 0 0 amux_2to1_4/SELB
flabel metal4 -10812 -64374 -10800 -64364 1 FreeSans 480 0 0 0 amux_2to1_4/VDD
flabel metal4 -10740 -69872 -10726 -69864 1 FreeSans 480 0 0 0 amux_2to1_4/VSS
flabel locali -11908 -67537 -11874 -67503 0 FreeSans 340 0 0 0 amux_2to1_4/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -11908 -67605 -11874 -67571 0 FreeSans 340 0 0 0 amux_2to1_4/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -12000 -67605 -11966 -67571 0 FreeSans 340 0 0 0 amux_2to1_4/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -12043 -67299 -12009 -67265 0 FreeSans 200 0 0 0 amux_2to1_4/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -12043 -67843 -12009 -67809 0 FreeSans 200 0 0 0 amux_2to1_4/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -12043 -67843 -12009 -67809 0 FreeSans 200 0 0 0 amux_2to1_4/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -12043 -67299 -12009 -67265 0 FreeSans 200 0 0 0 amux_2to1_4/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -12072 -67826 -12072 -67826 4 amux_2to1_4/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -8148 -67594 -8142 -67590 1 FreeSans 480 0 0 0 amux_2to1_5/SEL
flabel metal2 -6552 -67668 -6544 -67660 1 FreeSans 480 0 0 0 amux_2to1_5/A
flabel metal2 -6298 -67648 -6290 -67642 1 FreeSans 480 0 0 0 amux_2to1_5/Y
flabel metal2 -7074 -67646 -7064 -67640 1 FreeSans 480 0 0 0 amux_2to1_5/B
flabel metal2 -7688 -67646 -7678 -67636 1 FreeSans 480 0 0 0 amux_2to1_5/SELB
flabel metal4 -6812 -64374 -6800 -64364 1 FreeSans 480 0 0 0 amux_2to1_5/VDD
flabel metal4 -6740 -69872 -6726 -69864 1 FreeSans 480 0 0 0 amux_2to1_5/VSS
flabel locali -7908 -67537 -7874 -67503 0 FreeSans 340 0 0 0 amux_2to1_5/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -7908 -67605 -7874 -67571 0 FreeSans 340 0 0 0 amux_2to1_5/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -8000 -67605 -7966 -67571 0 FreeSans 340 0 0 0 amux_2to1_5/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -8043 -67299 -8009 -67265 0 FreeSans 200 0 0 0 amux_2to1_5/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -8043 -67843 -8009 -67809 0 FreeSans 200 0 0 0 amux_2to1_5/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -8043 -67843 -8009 -67809 0 FreeSans 200 0 0 0 amux_2to1_5/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -8043 -67299 -8009 -67265 0 FreeSans 200 0 0 0 amux_2to1_5/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -8072 -67826 -8072 -67826 4 amux_2to1_5/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -4148 -67594 -4142 -67590 1 FreeSans 480 0 0 0 amux_2to1_6/SEL
flabel metal2 -2552 -67668 -2544 -67660 1 FreeSans 480 0 0 0 amux_2to1_6/A
flabel metal2 -2298 -67648 -2290 -67642 1 FreeSans 480 0 0 0 amux_2to1_6/Y
flabel metal2 -3074 -67646 -3064 -67640 1 FreeSans 480 0 0 0 amux_2to1_6/B
flabel metal2 -3688 -67646 -3678 -67636 1 FreeSans 480 0 0 0 amux_2to1_6/SELB
flabel metal4 -2812 -64374 -2800 -64364 1 FreeSans 480 0 0 0 amux_2to1_6/VDD
flabel metal4 -2740 -69872 -2726 -69864 1 FreeSans 480 0 0 0 amux_2to1_6/VSS
flabel locali -3908 -67537 -3874 -67503 0 FreeSans 340 0 0 0 amux_2to1_6/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -3908 -67605 -3874 -67571 0 FreeSans 340 0 0 0 amux_2to1_6/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -4000 -67605 -3966 -67571 0 FreeSans 340 0 0 0 amux_2to1_6/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -4043 -67299 -4009 -67265 0 FreeSans 200 0 0 0 amux_2to1_6/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -4043 -67843 -4009 -67809 0 FreeSans 200 0 0 0 amux_2to1_6/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -4043 -67843 -4009 -67809 0 FreeSans 200 0 0 0 amux_2to1_6/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -4043 -67299 -4009 -67265 0 FreeSans 200 0 0 0 amux_2to1_6/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -4072 -67826 -4072 -67826 4 amux_2to1_6/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -148 -67594 -142 -67590 1 FreeSans 480 0 0 0 amux_2to1_7/SEL
flabel metal2 1448 -67668 1456 -67660 1 FreeSans 480 0 0 0 amux_2to1_7/A
flabel metal2 1702 -67648 1710 -67642 1 FreeSans 480 0 0 0 amux_2to1_7/Y
flabel metal2 926 -67646 936 -67640 1 FreeSans 480 0 0 0 amux_2to1_7/B
flabel metal2 312 -67646 322 -67636 1 FreeSans 480 0 0 0 amux_2to1_7/SELB
flabel metal4 1188 -64374 1200 -64364 1 FreeSans 480 0 0 0 amux_2to1_7/VDD
flabel metal4 1260 -69872 1274 -69864 1 FreeSans 480 0 0 0 amux_2to1_7/VSS
flabel locali 92 -67537 126 -67503 0 FreeSans 340 0 0 0 amux_2to1_7/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 92 -67605 126 -67571 0 FreeSans 340 0 0 0 amux_2to1_7/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 0 -67605 34 -67571 0 FreeSans 340 0 0 0 amux_2to1_7/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -43 -67299 -9 -67265 0 FreeSans 200 0 0 0 amux_2to1_7/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -43 -67843 -9 -67809 0 FreeSans 200 0 0 0 amux_2to1_7/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -43 -67843 -9 -67809 0 FreeSans 200 0 0 0 amux_2to1_7/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -43 -67299 -9 -67265 0 FreeSans 200 0 0 0 amux_2to1_7/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -72 -67826 -72 -67826 4 amux_2to1_7/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 3852 -67594 3858 -67590 1 FreeSans 480 0 0 0 amux_2to1_8/SEL
flabel metal2 5448 -67668 5456 -67660 1 FreeSans 480 0 0 0 amux_2to1_8/A
flabel metal2 5702 -67648 5710 -67642 1 FreeSans 480 0 0 0 amux_2to1_8/Y
flabel metal2 4926 -67646 4936 -67640 1 FreeSans 480 0 0 0 amux_2to1_8/B
flabel metal2 4312 -67646 4322 -67636 1 FreeSans 480 0 0 0 amux_2to1_8/SELB
flabel metal4 5188 -64374 5200 -64364 1 FreeSans 480 0 0 0 amux_2to1_8/VDD
flabel metal4 5260 -69872 5274 -69864 1 FreeSans 480 0 0 0 amux_2to1_8/VSS
flabel locali 4092 -67537 4126 -67503 0 FreeSans 340 0 0 0 amux_2to1_8/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 4092 -67605 4126 -67571 0 FreeSans 340 0 0 0 amux_2to1_8/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 4000 -67605 4034 -67571 0 FreeSans 340 0 0 0 amux_2to1_8/sky130_fd_sc_hd__inv_1_0/A
flabel nwell 3957 -67299 3991 -67265 0 FreeSans 200 0 0 0 amux_2to1_8/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 3957 -67843 3991 -67809 0 FreeSans 200 0 0 0 amux_2to1_8/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 3957 -67843 3991 -67809 0 FreeSans 200 0 0 0 amux_2to1_8/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 3957 -67299 3991 -67265 0 FreeSans 200 0 0 0 amux_2to1_8/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 3928 -67826 3928 -67826 4 amux_2to1_8/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 17366 -44330 17366 -44330 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias1
flabel metal1 19238 -51004 19238 -51004 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias2
flabel metal1 48624 -51296 48648 -51266 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/VSS
flabel metal1 49000 -50448 49000 -50448 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias3
flabel metal1 48744 -50242 48744 -50242 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascnm
flabel metal1 48880 -54474 48880 -54474 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias4
flabel metal1 27582 -50080 27610 -50050 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vtail_cascn
flabel metal1 27900 -46738 27932 -46698 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascnp
flabel metal1 28766 -43876 28856 -43846 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M8d
flabel metal1 27688 -50340 27726 -50304 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vmirror
flabel metal1 48382 -48608 48418 -48578 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M16d
flabel metal1 14798 -53518 14826 -53474 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vip
flabel metal1 26398 -53514 26430 -53476 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vim
flabel metal1 20242 -56944 20338 -56908 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/ibiasn
flabel metal1 25392 -54218 25440 -54194 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vtail_cascn
flabel metal4 14524 -58722 14550 -58700 1 FreeSans 3200 0 0 0 se_fold_casc_wide_swing_ota_0/VSS
flabel metal2 18880 -51912 18928 -51896 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpp
flabel metal1 15956 -54146 15988 -54118 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpm
flabel metal4 13740 -28068 13766 -27974 1 FreeSans 3200 0 0 0 se_fold_casc_wide_swing_ota_0/VDD
flabel metal4 26038 -42980 26058 -42960 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vo
flabel metal1 48052 -40350 48058 -40332 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vo
flabel metal1 32942 -33528 32974 -33496 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M9d
flabel metal1 28376 -36986 28448 -36956 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascnm
flabel metal1 31100 -36978 31142 -36956 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascnp
flabel metal1 29654 -37016 29680 -36978 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vtail_cascp
flabel metal1 29142 -41024 29172 -40998 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vip
flabel metal1 30150 -41028 30180 -40994 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vim
flabel metal2 45616 -36368 45678 -36340 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vmirror
flabel metal1 41654 -34164 41706 -34138 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/VDD
flabel metal2 35890 -35206 35958 -35176 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpp
flabel metal2 36114 -36238 36166 -36204 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpm
flabel metal2 33768 -30094 33768 -30094 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias1
flabel metal2 34746 -30356 34776 -30328 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/VDD
flabel metal1 31790 -31368 31824 -31346 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M7d
flabel metal2 33178 -31492 33236 -31456 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M13d
flabel metal2 35204 -33672 35282 -33638 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vtail_cascp
flabel metal1 42954 -37838 42990 -37810 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/VDD
flabel metal2 37310 -41886 37364 -41852 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M8d
flabel metal2 37734 -36898 37816 -36866 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias2
flabel metal2 42284 -39408 42346 -39378 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M16d
flabel metal2 41876 -39096 41940 -39064 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M13d
flabel metal1 32768 -37058 32808 -37024 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M7d
flabel metal2 47838 -39196 47900 -39164 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vmirror
flabel metal2 45952 -39306 46002 -39270 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpm
flabel metal2 46004 -40354 46096 -40322 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpp
flabel metal2 33062 -38026 33062 -38026 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias1
flabel metal2 32932 -41612 32988 -41578 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M9d
flabel locali 12258 -57513 12292 -57479 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 12258 -57581 12292 -57547 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 12350 -57581 12384 -57547 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/A
flabel nwell 12393 -57275 12427 -57241 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 12393 -57819 12427 -57785 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 12393 -57819 12427 -57785 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 12393 -57275 12427 -57241 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 12456 -57802 12456 -57802 6 sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal4 55802 -38836 55818 -38830 1 FreeSans 480 0 0 0 latched_comparator_folded_0/VDD
flabel metal1 52392 -41082 52406 -41070 1 FreeSans 480 0 0 0 latched_comparator_folded_0/vip
flabel metal1 53162 -41202 53172 -41192 1 FreeSans 480 0 0 0 latched_comparator_folded_0/vim
flabel metal1 55202 -40692 55216 -40672 1 FreeSans 480 0 0 0 latched_comparator_folded_0/vlatchm
flabel metal1 52768 -41158 52782 -41148 1 FreeSans 480 0 0 0 latched_comparator_folded_0/vlatchp
flabel metal1 53814 -40170 53832 -40156 1 FreeSans 480 0 0 0 latched_comparator_folded_0/vtailp
flabel metal1 53732 -40052 53752 -40040 1 FreeSans 480 0 0 0 latched_comparator_folded_0/ibiasp
flabel via1 56340 -40602 56356 -40586 1 FreeSans 480 0 0 0 latched_comparator_folded_0/vcompm
flabel metal1 58004 -40380 58024 -40356 1 FreeSans 480 0 0 0 latched_comparator_folded_0/vcompp
flabel metal4 55292 -43504 55318 -43484 1 FreeSans 480 0 0 0 latched_comparator_folded_0/VSS
flabel metal1 56838 -42538 56844 -42532 1 FreeSans 480 0 0 0 latched_comparator_folded_0/vlatchm
flabel metal2 56926 -43104 56934 -43096 1 FreeSans 480 0 0 0 latched_comparator_folded_0/vlatchp
flabel metal1 56634 -41904 56640 -41898 1 FreeSans 160 0 0 0 latched_comparator_folded_0/vcompm_buf
flabel metal1 56378 -41904 56384 -41900 1 FreeSans 160 0 0 0 latched_comparator_folded_0/vcompmb
flabel metal1 57402 -41900 57406 -41896 1 FreeSans 160 0 0 0 latched_comparator_folded_0/vcompp_buf
flabel metal1 57656 -41902 57662 -41898 1 FreeSans 160 0 0 0 latched_comparator_folded_0/vcomppb
flabel metal2 58152 -41960 58158 -41954 1 FreeSans 480 0 0 0 latched_comparator_folded_0/vop
flabel metal1 57084 -42022 57090 -42014 1 FreeSans 480 0 0 0 latched_comparator_folded_0/vom
flabel metal4 53930 -42522 53950 -42504 1 FreeSans 480 0 0 0 latched_comparator_folded_0/clk
flabel locali 57748 -41847 57782 -41813 0 FreeSans 340 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_3/Y
flabel locali 57748 -41915 57782 -41881 0 FreeSans 340 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_3/Y
flabel locali 57840 -41915 57874 -41881 0 FreeSans 340 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_3/A
flabel nwell 57883 -41609 57917 -41575 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_3/VPB
flabel pwell 57883 -42153 57917 -42119 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_3/VNB
flabel metal1 57883 -42153 57917 -42119 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_3/VGND
flabel metal1 57883 -41609 57917 -41575 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_3/VPWR
rlabel comment 57946 -42136 57946 -42136 6 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_3/inv_1
flabel locali 57472 -41847 57506 -41813 0 FreeSans 340 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_2/Y
flabel locali 57472 -41915 57506 -41881 0 FreeSans 340 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_2/Y
flabel locali 57564 -41915 57598 -41881 0 FreeSans 340 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_2/A
flabel nwell 57607 -41609 57641 -41575 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_2/VPB
flabel pwell 57607 -42153 57641 -42119 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_2/VNB
flabel metal1 57607 -42153 57641 -42119 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_2/VGND
flabel metal1 57607 -41609 57641 -41575 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_2/VPWR
rlabel comment 57670 -42136 57670 -42136 6 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_2/inv_1
flabel locali 56544 -41847 56578 -41813 0 FreeSans 340 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_1/Y
flabel locali 56544 -41915 56578 -41881 0 FreeSans 340 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_1/Y
flabel locali 56452 -41915 56486 -41881 0 FreeSans 340 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_1/A
flabel nwell 56409 -41609 56443 -41575 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_1/VPB
flabel pwell 56409 -42153 56443 -42119 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_1/VNB
flabel metal1 56409 -42153 56443 -42119 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_1/VGND
flabel metal1 56409 -41609 56443 -41575 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_1/VPWR
rlabel comment 56380 -42136 56380 -42136 4 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_1/inv_1
flabel locali 56268 -41847 56302 -41813 0 FreeSans 340 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 56268 -41915 56302 -41881 0 FreeSans 340 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 56176 -41915 56210 -41881 0 FreeSans 340 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_0/A
flabel nwell 56133 -41609 56167 -41575 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 56133 -42153 56167 -42119 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 56133 -42153 56167 -42119 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 56133 -41609 56167 -41575 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 56104 -42136 56104 -42136 4 latched_comparator_folded_0/sky130_fd_sc_hd__inv_1_0/inv_1
flabel locali 56776 -42051 56810 -42017 0 FreeSans 250 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_0/Y
flabel locali 56776 -41983 56810 -41949 0 FreeSans 250 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_0/Y
flabel locali 56776 -41915 56810 -41881 0 FreeSans 250 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_0/Y
flabel locali 56684 -41915 56718 -41881 0 FreeSans 250 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_0/B
flabel locali 56868 -41915 56902 -41881 0 FreeSans 250 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_0/A
flabel nwell 56684 -41609 56718 -41575 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_0/VPB
flabel pwell 56684 -42153 56718 -42119 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_0/VNB
flabel metal1 56684 -42153 56718 -42119 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_0/VGND
flabel metal1 56684 -41609 56718 -41575 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_0/VPWR
rlabel comment 56656 -42136 56656 -42136 4 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_0/nand2_1
flabel locali 57240 -42051 57274 -42017 0 FreeSans 250 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_1/Y
flabel locali 57240 -41983 57274 -41949 0 FreeSans 250 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_1/Y
flabel locali 57240 -41915 57274 -41881 0 FreeSans 250 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_1/Y
flabel locali 57332 -41915 57366 -41881 0 FreeSans 250 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_1/B
flabel locali 57148 -41915 57182 -41881 0 FreeSans 250 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_1/A
flabel nwell 57332 -41609 57366 -41575 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_1/VPB
flabel pwell 57332 -42153 57366 -42119 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_1/VNB
flabel metal1 57332 -42153 57366 -42119 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_1/VGND
flabel metal1 57332 -41609 57366 -41575 0 FreeSans 200 0 0 0 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_1/VPWR
rlabel comment 57394 -42136 57394 -42136 6 latched_comparator_folded_0/sky130_fd_sc_hd__nand2_1_1/nand2_1
<< end >>
