magic
tech sky130A
magscale 1 2
timestamp 1621819980
<< error_p >>
rect -410 400 -370 1000
rect -350 400 -310 1000
rect 309 400 349 1000
rect 369 400 409 1000
rect -410 -300 -370 300
rect -350 -300 -310 300
rect 309 -300 349 300
rect 369 -300 409 300
rect -410 -1000 -370 -400
rect -350 -1000 -310 -400
rect 309 -1000 349 -400
rect 369 -1000 409 -400
<< metal3 >>
rect -1069 972 -370 1000
rect -1069 428 -454 972
rect -390 428 -370 972
rect -1069 400 -370 428
rect -350 972 349 1000
rect -350 428 265 972
rect 329 428 349 972
rect -350 400 349 428
rect 369 972 1068 1000
rect 369 428 984 972
rect 1048 428 1068 972
rect 369 400 1068 428
rect -1069 272 -370 300
rect -1069 -272 -454 272
rect -390 -272 -370 272
rect -1069 -300 -370 -272
rect -350 272 349 300
rect -350 -272 265 272
rect 329 -272 349 272
rect -350 -300 349 -272
rect 369 272 1068 300
rect 369 -272 984 272
rect 1048 -272 1068 272
rect 369 -300 1068 -272
rect -1069 -428 -370 -400
rect -1069 -972 -454 -428
rect -390 -972 -370 -428
rect -1069 -1000 -370 -972
rect -350 -428 349 -400
rect -350 -972 265 -428
rect 329 -972 349 -428
rect -350 -1000 349 -972
rect 369 -428 1068 -400
rect 369 -972 984 -428
rect 1048 -972 1068 -428
rect 369 -1000 1068 -972
<< via3 >>
rect -454 428 -390 972
rect 265 428 329 972
rect 984 428 1048 972
rect -454 -272 -390 272
rect 265 -272 329 272
rect 984 -272 1048 272
rect -454 -972 -390 -428
rect 265 -972 329 -428
rect 984 -972 1048 -428
<< mimcap >>
rect -969 860 -569 900
rect -969 540 -929 860
rect -609 540 -569 860
rect -969 500 -569 540
rect -250 860 150 900
rect -250 540 -210 860
rect 110 540 150 860
rect -250 500 150 540
rect 469 860 869 900
rect 469 540 509 860
rect 829 540 869 860
rect 469 500 869 540
rect -969 160 -569 200
rect -969 -160 -929 160
rect -609 -160 -569 160
rect -969 -200 -569 -160
rect -250 160 150 200
rect -250 -160 -210 160
rect 110 -160 150 160
rect -250 -200 150 -160
rect 469 160 869 200
rect 469 -160 509 160
rect 829 -160 869 160
rect 469 -200 869 -160
rect -969 -540 -569 -500
rect -969 -860 -929 -540
rect -609 -860 -569 -540
rect -969 -900 -569 -860
rect -250 -540 150 -500
rect -250 -860 -210 -540
rect 110 -860 150 -540
rect -250 -900 150 -860
rect 469 -540 869 -500
rect 469 -860 509 -540
rect 829 -860 869 -540
rect 469 -900 869 -860
<< mimcapcontact >>
rect -929 540 -609 860
rect -210 540 110 860
rect 509 540 829 860
rect -929 -160 -609 160
rect -210 -160 110 160
rect 509 -160 829 160
rect -929 -860 -609 -540
rect -210 -860 110 -540
rect 509 -860 829 -540
<< metal4 >>
rect -470 972 -374 988
rect -930 860 -608 861
rect -930 540 -929 860
rect -609 540 -608 860
rect -930 539 -608 540
rect -470 428 -454 972
rect -390 428 -374 972
rect 249 972 345 988
rect -211 860 111 861
rect -211 540 -210 860
rect 110 540 111 860
rect -211 539 111 540
rect -470 412 -374 428
rect 249 428 265 972
rect 329 428 345 972
rect 968 972 1064 988
rect 508 860 830 861
rect 508 540 509 860
rect 829 540 830 860
rect 508 539 830 540
rect 249 412 345 428
rect 968 428 984 972
rect 1048 428 1064 972
rect 968 412 1064 428
rect -470 272 -374 288
rect -930 160 -608 161
rect -930 -160 -929 160
rect -609 -160 -608 160
rect -930 -161 -608 -160
rect -470 -272 -454 272
rect -390 -272 -374 272
rect 249 272 345 288
rect -211 160 111 161
rect -211 -160 -210 160
rect 110 -160 111 160
rect -211 -161 111 -160
rect -470 -288 -374 -272
rect 249 -272 265 272
rect 329 -272 345 272
rect 968 272 1064 288
rect 508 160 830 161
rect 508 -160 509 160
rect 829 -160 830 160
rect 508 -161 830 -160
rect 249 -288 345 -272
rect 968 -272 984 272
rect 1048 -272 1064 272
rect 968 -288 1064 -272
rect -470 -428 -374 -412
rect -930 -540 -608 -539
rect -930 -860 -929 -540
rect -609 -860 -608 -540
rect -930 -861 -608 -860
rect -470 -972 -454 -428
rect -390 -972 -374 -428
rect 249 -428 345 -412
rect -211 -540 111 -539
rect -211 -860 -210 -540
rect 110 -860 111 -540
rect -211 -861 111 -860
rect -470 -988 -374 -972
rect 249 -972 265 -428
rect 329 -972 345 -428
rect 968 -428 1064 -412
rect 508 -540 830 -539
rect 508 -860 509 -540
rect 829 -860 830 -540
rect 508 -861 830 -860
rect 249 -988 345 -972
rect 968 -972 984 -428
rect 1048 -972 1064 -428
rect 968 -988 1064 -972
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 369 400 969 1000
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 3 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
string library sky130
<< end >>
