magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1700 -12160 13960 4260
<< nwell >>
rect -398 -7578 12658 2958
<< pwell >>
rect -388 -7904 12648 -7752
rect -388 -10696 -236 -7904
rect 12496 -10696 12648 -7904
rect -388 -10848 12648 -10696
<< psubdiff >>
rect -362 -7811 12622 -7778
rect -362 -7845 -177 -7811
rect -143 -7845 -109 -7811
rect -75 -7845 -41 -7811
rect -7 -7845 27 -7811
rect 61 -7845 95 -7811
rect 129 -7845 163 -7811
rect 197 -7845 231 -7811
rect 265 -7845 299 -7811
rect 333 -7845 367 -7811
rect 401 -7845 435 -7811
rect 469 -7845 503 -7811
rect 537 -7845 571 -7811
rect 605 -7845 639 -7811
rect 673 -7845 707 -7811
rect 741 -7845 775 -7811
rect 809 -7845 843 -7811
rect 877 -7845 911 -7811
rect 945 -7845 979 -7811
rect 1013 -7845 1047 -7811
rect 1081 -7845 1115 -7811
rect 1149 -7845 1183 -7811
rect 1217 -7845 1251 -7811
rect 1285 -7845 1319 -7811
rect 1353 -7845 1387 -7811
rect 1421 -7845 1455 -7811
rect 1489 -7845 1523 -7811
rect 1557 -7845 1591 -7811
rect 1625 -7845 1659 -7811
rect 1693 -7845 1727 -7811
rect 1761 -7845 1795 -7811
rect 1829 -7845 1863 -7811
rect 1897 -7845 1931 -7811
rect 1965 -7845 1999 -7811
rect 2033 -7845 2067 -7811
rect 2101 -7845 2135 -7811
rect 2169 -7845 2203 -7811
rect 2237 -7845 2271 -7811
rect 2305 -7845 2339 -7811
rect 2373 -7845 2407 -7811
rect 2441 -7845 2475 -7811
rect 2509 -7845 2543 -7811
rect 2577 -7845 2611 -7811
rect 2645 -7845 2679 -7811
rect 2713 -7845 2747 -7811
rect 2781 -7845 2815 -7811
rect 2849 -7845 2883 -7811
rect 2917 -7845 2951 -7811
rect 2985 -7845 3019 -7811
rect 3053 -7845 3087 -7811
rect 3121 -7845 3155 -7811
rect 3189 -7845 3223 -7811
rect 3257 -7845 3291 -7811
rect 3325 -7845 3359 -7811
rect 3393 -7845 3427 -7811
rect 3461 -7845 3495 -7811
rect 3529 -7845 3563 -7811
rect 3597 -7845 3631 -7811
rect 3665 -7845 3699 -7811
rect 3733 -7845 3767 -7811
rect 3801 -7845 3835 -7811
rect 3869 -7845 3903 -7811
rect 3937 -7845 3971 -7811
rect 4005 -7845 4039 -7811
rect 4073 -7845 4107 -7811
rect 4141 -7845 4175 -7811
rect 4209 -7845 4243 -7811
rect 4277 -7845 4311 -7811
rect 4345 -7845 4379 -7811
rect 4413 -7845 4447 -7811
rect 4481 -7845 4515 -7811
rect 4549 -7845 4583 -7811
rect 4617 -7845 4651 -7811
rect 4685 -7845 4719 -7811
rect 4753 -7845 4787 -7811
rect 4821 -7845 4855 -7811
rect 4889 -7845 4923 -7811
rect 4957 -7845 4991 -7811
rect 5025 -7845 5059 -7811
rect 5093 -7845 5127 -7811
rect 5161 -7845 5195 -7811
rect 5229 -7845 5263 -7811
rect 5297 -7845 5331 -7811
rect 5365 -7845 5399 -7811
rect 5433 -7845 5467 -7811
rect 5501 -7845 5535 -7811
rect 5569 -7845 5603 -7811
rect 5637 -7845 5671 -7811
rect 5705 -7845 5739 -7811
rect 5773 -7845 5807 -7811
rect 5841 -7845 5875 -7811
rect 5909 -7845 5943 -7811
rect 5977 -7845 6011 -7811
rect 6045 -7845 6079 -7811
rect 6113 -7845 6147 -7811
rect 6181 -7845 6215 -7811
rect 6249 -7845 6283 -7811
rect 6317 -7845 6351 -7811
rect 6385 -7845 6419 -7811
rect 6453 -7845 6487 -7811
rect 6521 -7845 6555 -7811
rect 6589 -7845 6623 -7811
rect 6657 -7845 6691 -7811
rect 6725 -7845 6759 -7811
rect 6793 -7845 6827 -7811
rect 6861 -7845 6895 -7811
rect 6929 -7845 6963 -7811
rect 6997 -7845 7031 -7811
rect 7065 -7845 7099 -7811
rect 7133 -7845 7167 -7811
rect 7201 -7845 7235 -7811
rect 7269 -7845 7303 -7811
rect 7337 -7845 7371 -7811
rect 7405 -7845 7439 -7811
rect 7473 -7845 7507 -7811
rect 7541 -7845 7575 -7811
rect 7609 -7845 7643 -7811
rect 7677 -7845 7711 -7811
rect 7745 -7845 7779 -7811
rect 7813 -7845 7847 -7811
rect 7881 -7845 7915 -7811
rect 7949 -7845 7983 -7811
rect 8017 -7845 8051 -7811
rect 8085 -7845 8119 -7811
rect 8153 -7845 8187 -7811
rect 8221 -7845 8255 -7811
rect 8289 -7845 8323 -7811
rect 8357 -7845 8391 -7811
rect 8425 -7845 8459 -7811
rect 8493 -7845 8527 -7811
rect 8561 -7845 8595 -7811
rect 8629 -7845 8663 -7811
rect 8697 -7845 8731 -7811
rect 8765 -7845 8799 -7811
rect 8833 -7845 8867 -7811
rect 8901 -7845 8935 -7811
rect 8969 -7845 9003 -7811
rect 9037 -7845 9071 -7811
rect 9105 -7845 9139 -7811
rect 9173 -7845 9207 -7811
rect 9241 -7845 9275 -7811
rect 9309 -7845 9343 -7811
rect 9377 -7845 9411 -7811
rect 9445 -7845 9479 -7811
rect 9513 -7845 9547 -7811
rect 9581 -7845 9615 -7811
rect 9649 -7845 9683 -7811
rect 9717 -7845 9751 -7811
rect 9785 -7845 9819 -7811
rect 9853 -7845 9887 -7811
rect 9921 -7845 9955 -7811
rect 9989 -7845 10023 -7811
rect 10057 -7845 10091 -7811
rect 10125 -7845 10159 -7811
rect 10193 -7845 10227 -7811
rect 10261 -7845 10295 -7811
rect 10329 -7845 10363 -7811
rect 10397 -7845 10431 -7811
rect 10465 -7845 10499 -7811
rect 10533 -7845 10567 -7811
rect 10601 -7845 10635 -7811
rect 10669 -7845 10703 -7811
rect 10737 -7845 10771 -7811
rect 10805 -7845 10839 -7811
rect 10873 -7845 10907 -7811
rect 10941 -7845 10975 -7811
rect 11009 -7845 11043 -7811
rect 11077 -7845 11111 -7811
rect 11145 -7845 11179 -7811
rect 11213 -7845 11247 -7811
rect 11281 -7845 11315 -7811
rect 11349 -7845 11383 -7811
rect 11417 -7845 11451 -7811
rect 11485 -7845 11519 -7811
rect 11553 -7845 11587 -7811
rect 11621 -7845 11655 -7811
rect 11689 -7845 11723 -7811
rect 11757 -7845 11791 -7811
rect 11825 -7845 11859 -7811
rect 11893 -7845 11927 -7811
rect 11961 -7845 11995 -7811
rect 12029 -7845 12063 -7811
rect 12097 -7845 12131 -7811
rect 12165 -7845 12199 -7811
rect 12233 -7845 12267 -7811
rect 12301 -7845 12335 -7811
rect 12369 -7845 12403 -7811
rect 12437 -7845 12622 -7811
rect -362 -7878 12622 -7845
rect -362 -7957 -262 -7878
rect -362 -7991 -329 -7957
rect -295 -7991 -262 -7957
rect -362 -8025 -262 -7991
rect -362 -8059 -329 -8025
rect -295 -8059 -262 -8025
rect -362 -8093 -262 -8059
rect -362 -8127 -329 -8093
rect -295 -8127 -262 -8093
rect -362 -8161 -262 -8127
rect -362 -8195 -329 -8161
rect -295 -8195 -262 -8161
rect -362 -8229 -262 -8195
rect -362 -8263 -329 -8229
rect -295 -8263 -262 -8229
rect -362 -8297 -262 -8263
rect -362 -8331 -329 -8297
rect -295 -8331 -262 -8297
rect -362 -8365 -262 -8331
rect -362 -8399 -329 -8365
rect -295 -8399 -262 -8365
rect -362 -8433 -262 -8399
rect -362 -8467 -329 -8433
rect -295 -8467 -262 -8433
rect -362 -8501 -262 -8467
rect -362 -8535 -329 -8501
rect -295 -8535 -262 -8501
rect -362 -8569 -262 -8535
rect -362 -8603 -329 -8569
rect -295 -8603 -262 -8569
rect -362 -8637 -262 -8603
rect -362 -8671 -329 -8637
rect -295 -8671 -262 -8637
rect -362 -8705 -262 -8671
rect -362 -8739 -329 -8705
rect -295 -8739 -262 -8705
rect -362 -8773 -262 -8739
rect -362 -8807 -329 -8773
rect -295 -8807 -262 -8773
rect -362 -8841 -262 -8807
rect -362 -8875 -329 -8841
rect -295 -8875 -262 -8841
rect -362 -8909 -262 -8875
rect -362 -8943 -329 -8909
rect -295 -8943 -262 -8909
rect -362 -8977 -262 -8943
rect -362 -9011 -329 -8977
rect -295 -9011 -262 -8977
rect -362 -9045 -262 -9011
rect -362 -9079 -329 -9045
rect -295 -9079 -262 -9045
rect -362 -9113 -262 -9079
rect -362 -9147 -329 -9113
rect -295 -9147 -262 -9113
rect -362 -9181 -262 -9147
rect -362 -9215 -329 -9181
rect -295 -9215 -262 -9181
rect -362 -9249 -262 -9215
rect -362 -9283 -329 -9249
rect -295 -9283 -262 -9249
rect -362 -9317 -262 -9283
rect -362 -9351 -329 -9317
rect -295 -9351 -262 -9317
rect -362 -9385 -262 -9351
rect -362 -9419 -329 -9385
rect -295 -9419 -262 -9385
rect -362 -9453 -262 -9419
rect -362 -9487 -329 -9453
rect -295 -9487 -262 -9453
rect -362 -9521 -262 -9487
rect -362 -9555 -329 -9521
rect -295 -9555 -262 -9521
rect -362 -9589 -262 -9555
rect -362 -9623 -329 -9589
rect -295 -9623 -262 -9589
rect -362 -9657 -262 -9623
rect -362 -9691 -329 -9657
rect -295 -9691 -262 -9657
rect -362 -9725 -262 -9691
rect -362 -9759 -329 -9725
rect -295 -9759 -262 -9725
rect -362 -9793 -262 -9759
rect -362 -9827 -329 -9793
rect -295 -9827 -262 -9793
rect -362 -9861 -262 -9827
rect -362 -9895 -329 -9861
rect -295 -9895 -262 -9861
rect -362 -9929 -262 -9895
rect -362 -9963 -329 -9929
rect -295 -9963 -262 -9929
rect -362 -9997 -262 -9963
rect -362 -10031 -329 -9997
rect -295 -10031 -262 -9997
rect -362 -10065 -262 -10031
rect -362 -10099 -329 -10065
rect -295 -10099 -262 -10065
rect -362 -10133 -262 -10099
rect -362 -10167 -329 -10133
rect -295 -10167 -262 -10133
rect -362 -10201 -262 -10167
rect -362 -10235 -329 -10201
rect -295 -10235 -262 -10201
rect -362 -10269 -262 -10235
rect -362 -10303 -329 -10269
rect -295 -10303 -262 -10269
rect -362 -10337 -262 -10303
rect -362 -10371 -329 -10337
rect -295 -10371 -262 -10337
rect -362 -10405 -262 -10371
rect -362 -10439 -329 -10405
rect -295 -10439 -262 -10405
rect -362 -10473 -262 -10439
rect -362 -10507 -329 -10473
rect -295 -10507 -262 -10473
rect -362 -10541 -262 -10507
rect -362 -10575 -329 -10541
rect -295 -10575 -262 -10541
rect -362 -10609 -262 -10575
rect -362 -10643 -329 -10609
rect -295 -10643 -262 -10609
rect -362 -10722 -262 -10643
rect 12522 -7957 12622 -7878
rect 12522 -7991 12555 -7957
rect 12589 -7991 12622 -7957
rect 12522 -8025 12622 -7991
rect 12522 -8059 12555 -8025
rect 12589 -8059 12622 -8025
rect 12522 -8093 12622 -8059
rect 12522 -8127 12555 -8093
rect 12589 -8127 12622 -8093
rect 12522 -8161 12622 -8127
rect 12522 -8195 12555 -8161
rect 12589 -8195 12622 -8161
rect 12522 -8229 12622 -8195
rect 12522 -8263 12555 -8229
rect 12589 -8263 12622 -8229
rect 12522 -8297 12622 -8263
rect 12522 -8331 12555 -8297
rect 12589 -8331 12622 -8297
rect 12522 -8365 12622 -8331
rect 12522 -8399 12555 -8365
rect 12589 -8399 12622 -8365
rect 12522 -8433 12622 -8399
rect 12522 -8467 12555 -8433
rect 12589 -8467 12622 -8433
rect 12522 -8501 12622 -8467
rect 12522 -8535 12555 -8501
rect 12589 -8535 12622 -8501
rect 12522 -8569 12622 -8535
rect 12522 -8603 12555 -8569
rect 12589 -8603 12622 -8569
rect 12522 -8637 12622 -8603
rect 12522 -8671 12555 -8637
rect 12589 -8671 12622 -8637
rect 12522 -8705 12622 -8671
rect 12522 -8739 12555 -8705
rect 12589 -8739 12622 -8705
rect 12522 -8773 12622 -8739
rect 12522 -8807 12555 -8773
rect 12589 -8807 12622 -8773
rect 12522 -8841 12622 -8807
rect 12522 -8875 12555 -8841
rect 12589 -8875 12622 -8841
rect 12522 -8909 12622 -8875
rect 12522 -8943 12555 -8909
rect 12589 -8943 12622 -8909
rect 12522 -8977 12622 -8943
rect 12522 -9011 12555 -8977
rect 12589 -9011 12622 -8977
rect 12522 -9045 12622 -9011
rect 12522 -9079 12555 -9045
rect 12589 -9079 12622 -9045
rect 12522 -9113 12622 -9079
rect 12522 -9147 12555 -9113
rect 12589 -9147 12622 -9113
rect 12522 -9181 12622 -9147
rect 12522 -9215 12555 -9181
rect 12589 -9215 12622 -9181
rect 12522 -9249 12622 -9215
rect 12522 -9283 12555 -9249
rect 12589 -9283 12622 -9249
rect 12522 -9317 12622 -9283
rect 12522 -9351 12555 -9317
rect 12589 -9351 12622 -9317
rect 12522 -9385 12622 -9351
rect 12522 -9419 12555 -9385
rect 12589 -9419 12622 -9385
rect 12522 -9453 12622 -9419
rect 12522 -9487 12555 -9453
rect 12589 -9487 12622 -9453
rect 12522 -9521 12622 -9487
rect 12522 -9555 12555 -9521
rect 12589 -9555 12622 -9521
rect 12522 -9589 12622 -9555
rect 12522 -9623 12555 -9589
rect 12589 -9623 12622 -9589
rect 12522 -9657 12622 -9623
rect 12522 -9691 12555 -9657
rect 12589 -9691 12622 -9657
rect 12522 -9725 12622 -9691
rect 12522 -9759 12555 -9725
rect 12589 -9759 12622 -9725
rect 12522 -9793 12622 -9759
rect 12522 -9827 12555 -9793
rect 12589 -9827 12622 -9793
rect 12522 -9861 12622 -9827
rect 12522 -9895 12555 -9861
rect 12589 -9895 12622 -9861
rect 12522 -9929 12622 -9895
rect 12522 -9963 12555 -9929
rect 12589 -9963 12622 -9929
rect 12522 -9997 12622 -9963
rect 12522 -10031 12555 -9997
rect 12589 -10031 12622 -9997
rect 12522 -10065 12622 -10031
rect 12522 -10099 12555 -10065
rect 12589 -10099 12622 -10065
rect 12522 -10133 12622 -10099
rect 12522 -10167 12555 -10133
rect 12589 -10167 12622 -10133
rect 12522 -10201 12622 -10167
rect 12522 -10235 12555 -10201
rect 12589 -10235 12622 -10201
rect 12522 -10269 12622 -10235
rect 12522 -10303 12555 -10269
rect 12589 -10303 12622 -10269
rect 12522 -10337 12622 -10303
rect 12522 -10371 12555 -10337
rect 12589 -10371 12622 -10337
rect 12522 -10405 12622 -10371
rect 12522 -10439 12555 -10405
rect 12589 -10439 12622 -10405
rect 12522 -10473 12622 -10439
rect 12522 -10507 12555 -10473
rect 12589 -10507 12622 -10473
rect 12522 -10541 12622 -10507
rect 12522 -10575 12555 -10541
rect 12589 -10575 12622 -10541
rect 12522 -10609 12622 -10575
rect 12522 -10643 12555 -10609
rect 12589 -10643 12622 -10609
rect 12522 -10722 12622 -10643
rect -362 -10755 12622 -10722
rect -362 -10789 -177 -10755
rect -143 -10789 -109 -10755
rect -75 -10789 -41 -10755
rect -7 -10789 27 -10755
rect 61 -10789 95 -10755
rect 129 -10789 163 -10755
rect 197 -10789 231 -10755
rect 265 -10789 299 -10755
rect 333 -10789 367 -10755
rect 401 -10789 435 -10755
rect 469 -10789 503 -10755
rect 537 -10789 571 -10755
rect 605 -10789 639 -10755
rect 673 -10789 707 -10755
rect 741 -10789 775 -10755
rect 809 -10789 843 -10755
rect 877 -10789 911 -10755
rect 945 -10789 979 -10755
rect 1013 -10789 1047 -10755
rect 1081 -10789 1115 -10755
rect 1149 -10789 1183 -10755
rect 1217 -10789 1251 -10755
rect 1285 -10789 1319 -10755
rect 1353 -10789 1387 -10755
rect 1421 -10789 1455 -10755
rect 1489 -10789 1523 -10755
rect 1557 -10789 1591 -10755
rect 1625 -10789 1659 -10755
rect 1693 -10789 1727 -10755
rect 1761 -10789 1795 -10755
rect 1829 -10789 1863 -10755
rect 1897 -10789 1931 -10755
rect 1965 -10789 1999 -10755
rect 2033 -10789 2067 -10755
rect 2101 -10789 2135 -10755
rect 2169 -10789 2203 -10755
rect 2237 -10789 2271 -10755
rect 2305 -10789 2339 -10755
rect 2373 -10789 2407 -10755
rect 2441 -10789 2475 -10755
rect 2509 -10789 2543 -10755
rect 2577 -10789 2611 -10755
rect 2645 -10789 2679 -10755
rect 2713 -10789 2747 -10755
rect 2781 -10789 2815 -10755
rect 2849 -10789 2883 -10755
rect 2917 -10789 2951 -10755
rect 2985 -10789 3019 -10755
rect 3053 -10789 3087 -10755
rect 3121 -10789 3155 -10755
rect 3189 -10789 3223 -10755
rect 3257 -10789 3291 -10755
rect 3325 -10789 3359 -10755
rect 3393 -10789 3427 -10755
rect 3461 -10789 3495 -10755
rect 3529 -10789 3563 -10755
rect 3597 -10789 3631 -10755
rect 3665 -10789 3699 -10755
rect 3733 -10789 3767 -10755
rect 3801 -10789 3835 -10755
rect 3869 -10789 3903 -10755
rect 3937 -10789 3971 -10755
rect 4005 -10789 4039 -10755
rect 4073 -10789 4107 -10755
rect 4141 -10789 4175 -10755
rect 4209 -10789 4243 -10755
rect 4277 -10789 4311 -10755
rect 4345 -10789 4379 -10755
rect 4413 -10789 4447 -10755
rect 4481 -10789 4515 -10755
rect 4549 -10789 4583 -10755
rect 4617 -10789 4651 -10755
rect 4685 -10789 4719 -10755
rect 4753 -10789 4787 -10755
rect 4821 -10789 4855 -10755
rect 4889 -10789 4923 -10755
rect 4957 -10789 4991 -10755
rect 5025 -10789 5059 -10755
rect 5093 -10789 5127 -10755
rect 5161 -10789 5195 -10755
rect 5229 -10789 5263 -10755
rect 5297 -10789 5331 -10755
rect 5365 -10789 5399 -10755
rect 5433 -10789 5467 -10755
rect 5501 -10789 5535 -10755
rect 5569 -10789 5603 -10755
rect 5637 -10789 5671 -10755
rect 5705 -10789 5739 -10755
rect 5773 -10789 5807 -10755
rect 5841 -10789 5875 -10755
rect 5909 -10789 5943 -10755
rect 5977 -10789 6011 -10755
rect 6045 -10789 6079 -10755
rect 6113 -10789 6147 -10755
rect 6181 -10789 6215 -10755
rect 6249 -10789 6283 -10755
rect 6317 -10789 6351 -10755
rect 6385 -10789 6419 -10755
rect 6453 -10789 6487 -10755
rect 6521 -10789 6555 -10755
rect 6589 -10789 6623 -10755
rect 6657 -10789 6691 -10755
rect 6725 -10789 6759 -10755
rect 6793 -10789 6827 -10755
rect 6861 -10789 6895 -10755
rect 6929 -10789 6963 -10755
rect 6997 -10789 7031 -10755
rect 7065 -10789 7099 -10755
rect 7133 -10789 7167 -10755
rect 7201 -10789 7235 -10755
rect 7269 -10789 7303 -10755
rect 7337 -10789 7371 -10755
rect 7405 -10789 7439 -10755
rect 7473 -10789 7507 -10755
rect 7541 -10789 7575 -10755
rect 7609 -10789 7643 -10755
rect 7677 -10789 7711 -10755
rect 7745 -10789 7779 -10755
rect 7813 -10789 7847 -10755
rect 7881 -10789 7915 -10755
rect 7949 -10789 7983 -10755
rect 8017 -10789 8051 -10755
rect 8085 -10789 8119 -10755
rect 8153 -10789 8187 -10755
rect 8221 -10789 8255 -10755
rect 8289 -10789 8323 -10755
rect 8357 -10789 8391 -10755
rect 8425 -10789 8459 -10755
rect 8493 -10789 8527 -10755
rect 8561 -10789 8595 -10755
rect 8629 -10789 8663 -10755
rect 8697 -10789 8731 -10755
rect 8765 -10789 8799 -10755
rect 8833 -10789 8867 -10755
rect 8901 -10789 8935 -10755
rect 8969 -10789 9003 -10755
rect 9037 -10789 9071 -10755
rect 9105 -10789 9139 -10755
rect 9173 -10789 9207 -10755
rect 9241 -10789 9275 -10755
rect 9309 -10789 9343 -10755
rect 9377 -10789 9411 -10755
rect 9445 -10789 9479 -10755
rect 9513 -10789 9547 -10755
rect 9581 -10789 9615 -10755
rect 9649 -10789 9683 -10755
rect 9717 -10789 9751 -10755
rect 9785 -10789 9819 -10755
rect 9853 -10789 9887 -10755
rect 9921 -10789 9955 -10755
rect 9989 -10789 10023 -10755
rect 10057 -10789 10091 -10755
rect 10125 -10789 10159 -10755
rect 10193 -10789 10227 -10755
rect 10261 -10789 10295 -10755
rect 10329 -10789 10363 -10755
rect 10397 -10789 10431 -10755
rect 10465 -10789 10499 -10755
rect 10533 -10789 10567 -10755
rect 10601 -10789 10635 -10755
rect 10669 -10789 10703 -10755
rect 10737 -10789 10771 -10755
rect 10805 -10789 10839 -10755
rect 10873 -10789 10907 -10755
rect 10941 -10789 10975 -10755
rect 11009 -10789 11043 -10755
rect 11077 -10789 11111 -10755
rect 11145 -10789 11179 -10755
rect 11213 -10789 11247 -10755
rect 11281 -10789 11315 -10755
rect 11349 -10789 11383 -10755
rect 11417 -10789 11451 -10755
rect 11485 -10789 11519 -10755
rect 11553 -10789 11587 -10755
rect 11621 -10789 11655 -10755
rect 11689 -10789 11723 -10755
rect 11757 -10789 11791 -10755
rect 11825 -10789 11859 -10755
rect 11893 -10789 11927 -10755
rect 11961 -10789 11995 -10755
rect 12029 -10789 12063 -10755
rect 12097 -10789 12131 -10755
rect 12165 -10789 12199 -10755
rect 12233 -10789 12267 -10755
rect 12301 -10789 12335 -10755
rect 12369 -10789 12403 -10755
rect 12437 -10789 12622 -10755
rect -362 -10822 12622 -10789
<< nsubdiff >>
rect -362 2889 12622 2922
rect -362 2855 -177 2889
rect -143 2855 -109 2889
rect -75 2855 -41 2889
rect -7 2855 27 2889
rect 61 2855 95 2889
rect 129 2855 163 2889
rect 197 2855 231 2889
rect 265 2855 299 2889
rect 333 2855 367 2889
rect 401 2855 435 2889
rect 469 2855 503 2889
rect 537 2855 571 2889
rect 605 2855 639 2889
rect 673 2855 707 2889
rect 741 2855 775 2889
rect 809 2855 843 2889
rect 877 2855 911 2889
rect 945 2855 979 2889
rect 1013 2855 1047 2889
rect 1081 2855 1115 2889
rect 1149 2855 1183 2889
rect 1217 2855 1251 2889
rect 1285 2855 1319 2889
rect 1353 2855 1387 2889
rect 1421 2855 1455 2889
rect 1489 2855 1523 2889
rect 1557 2855 1591 2889
rect 1625 2855 1659 2889
rect 1693 2855 1727 2889
rect 1761 2855 1795 2889
rect 1829 2855 1863 2889
rect 1897 2855 1931 2889
rect 1965 2855 1999 2889
rect 2033 2855 2067 2889
rect 2101 2855 2135 2889
rect 2169 2855 2203 2889
rect 2237 2855 2271 2889
rect 2305 2855 2339 2889
rect 2373 2855 2407 2889
rect 2441 2855 2475 2889
rect 2509 2855 2543 2889
rect 2577 2855 2611 2889
rect 2645 2855 2679 2889
rect 2713 2855 2747 2889
rect 2781 2855 2815 2889
rect 2849 2855 2883 2889
rect 2917 2855 2951 2889
rect 2985 2855 3019 2889
rect 3053 2855 3087 2889
rect 3121 2855 3155 2889
rect 3189 2855 3223 2889
rect 3257 2855 3291 2889
rect 3325 2855 3359 2889
rect 3393 2855 3427 2889
rect 3461 2855 3495 2889
rect 3529 2855 3563 2889
rect 3597 2855 3631 2889
rect 3665 2855 3699 2889
rect 3733 2855 3767 2889
rect 3801 2855 3835 2889
rect 3869 2855 3903 2889
rect 3937 2855 3971 2889
rect 4005 2855 4039 2889
rect 4073 2855 4107 2889
rect 4141 2855 4175 2889
rect 4209 2855 4243 2889
rect 4277 2855 4311 2889
rect 4345 2855 4379 2889
rect 4413 2855 4447 2889
rect 4481 2855 4515 2889
rect 4549 2855 4583 2889
rect 4617 2855 4651 2889
rect 4685 2855 4719 2889
rect 4753 2855 4787 2889
rect 4821 2855 4855 2889
rect 4889 2855 4923 2889
rect 4957 2855 4991 2889
rect 5025 2855 5059 2889
rect 5093 2855 5127 2889
rect 5161 2855 5195 2889
rect 5229 2855 5263 2889
rect 5297 2855 5331 2889
rect 5365 2855 5399 2889
rect 5433 2855 5467 2889
rect 5501 2855 5535 2889
rect 5569 2855 5603 2889
rect 5637 2855 5671 2889
rect 5705 2855 5739 2889
rect 5773 2855 5807 2889
rect 5841 2855 5875 2889
rect 5909 2855 5943 2889
rect 5977 2855 6011 2889
rect 6045 2855 6079 2889
rect 6113 2855 6147 2889
rect 6181 2855 6215 2889
rect 6249 2855 6283 2889
rect 6317 2855 6351 2889
rect 6385 2855 6419 2889
rect 6453 2855 6487 2889
rect 6521 2855 6555 2889
rect 6589 2855 6623 2889
rect 6657 2855 6691 2889
rect 6725 2855 6759 2889
rect 6793 2855 6827 2889
rect 6861 2855 6895 2889
rect 6929 2855 6963 2889
rect 6997 2855 7031 2889
rect 7065 2855 7099 2889
rect 7133 2855 7167 2889
rect 7201 2855 7235 2889
rect 7269 2855 7303 2889
rect 7337 2855 7371 2889
rect 7405 2855 7439 2889
rect 7473 2855 7507 2889
rect 7541 2855 7575 2889
rect 7609 2855 7643 2889
rect 7677 2855 7711 2889
rect 7745 2855 7779 2889
rect 7813 2855 7847 2889
rect 7881 2855 7915 2889
rect 7949 2855 7983 2889
rect 8017 2855 8051 2889
rect 8085 2855 8119 2889
rect 8153 2855 8187 2889
rect 8221 2855 8255 2889
rect 8289 2855 8323 2889
rect 8357 2855 8391 2889
rect 8425 2855 8459 2889
rect 8493 2855 8527 2889
rect 8561 2855 8595 2889
rect 8629 2855 8663 2889
rect 8697 2855 8731 2889
rect 8765 2855 8799 2889
rect 8833 2855 8867 2889
rect 8901 2855 8935 2889
rect 8969 2855 9003 2889
rect 9037 2855 9071 2889
rect 9105 2855 9139 2889
rect 9173 2855 9207 2889
rect 9241 2855 9275 2889
rect 9309 2855 9343 2889
rect 9377 2855 9411 2889
rect 9445 2855 9479 2889
rect 9513 2855 9547 2889
rect 9581 2855 9615 2889
rect 9649 2855 9683 2889
rect 9717 2855 9751 2889
rect 9785 2855 9819 2889
rect 9853 2855 9887 2889
rect 9921 2855 9955 2889
rect 9989 2855 10023 2889
rect 10057 2855 10091 2889
rect 10125 2855 10159 2889
rect 10193 2855 10227 2889
rect 10261 2855 10295 2889
rect 10329 2855 10363 2889
rect 10397 2855 10431 2889
rect 10465 2855 10499 2889
rect 10533 2855 10567 2889
rect 10601 2855 10635 2889
rect 10669 2855 10703 2889
rect 10737 2855 10771 2889
rect 10805 2855 10839 2889
rect 10873 2855 10907 2889
rect 10941 2855 10975 2889
rect 11009 2855 11043 2889
rect 11077 2855 11111 2889
rect 11145 2855 11179 2889
rect 11213 2855 11247 2889
rect 11281 2855 11315 2889
rect 11349 2855 11383 2889
rect 11417 2855 11451 2889
rect 11485 2855 11519 2889
rect 11553 2855 11587 2889
rect 11621 2855 11655 2889
rect 11689 2855 11723 2889
rect 11757 2855 11791 2889
rect 11825 2855 11859 2889
rect 11893 2855 11927 2889
rect 11961 2855 11995 2889
rect 12029 2855 12063 2889
rect 12097 2855 12131 2889
rect 12165 2855 12199 2889
rect 12233 2855 12267 2889
rect 12301 2855 12335 2889
rect 12369 2855 12403 2889
rect 12437 2855 12622 2889
rect -362 2822 12622 2855
rect -362 2739 -262 2822
rect -362 2705 -329 2739
rect -295 2705 -262 2739
rect -362 2671 -262 2705
rect -362 2637 -329 2671
rect -295 2637 -262 2671
rect -362 2603 -262 2637
rect -362 2569 -329 2603
rect -295 2569 -262 2603
rect -362 2535 -262 2569
rect -362 2501 -329 2535
rect -295 2501 -262 2535
rect -362 2467 -262 2501
rect -362 2433 -329 2467
rect -295 2433 -262 2467
rect -362 2399 -262 2433
rect -362 2365 -329 2399
rect -295 2365 -262 2399
rect -362 2331 -262 2365
rect -362 2297 -329 2331
rect -295 2297 -262 2331
rect -362 2263 -262 2297
rect -362 2229 -329 2263
rect -295 2229 -262 2263
rect -362 2195 -262 2229
rect -362 2161 -329 2195
rect -295 2161 -262 2195
rect -362 2127 -262 2161
rect -362 2093 -329 2127
rect -295 2093 -262 2127
rect -362 2059 -262 2093
rect -362 2025 -329 2059
rect -295 2025 -262 2059
rect -362 1991 -262 2025
rect -362 1957 -329 1991
rect -295 1957 -262 1991
rect -362 1923 -262 1957
rect -362 1889 -329 1923
rect -295 1889 -262 1923
rect -362 1855 -262 1889
rect -362 1821 -329 1855
rect -295 1821 -262 1855
rect -362 1787 -262 1821
rect -362 1753 -329 1787
rect -295 1753 -262 1787
rect -362 1719 -262 1753
rect -362 1685 -329 1719
rect -295 1685 -262 1719
rect -362 1651 -262 1685
rect -362 1617 -329 1651
rect -295 1617 -262 1651
rect -362 1583 -262 1617
rect -362 1549 -329 1583
rect -295 1549 -262 1583
rect -362 1515 -262 1549
rect -362 1481 -329 1515
rect -295 1481 -262 1515
rect -362 1447 -262 1481
rect -362 1413 -329 1447
rect -295 1413 -262 1447
rect -362 1379 -262 1413
rect -362 1345 -329 1379
rect -295 1345 -262 1379
rect -362 1311 -262 1345
rect -362 1277 -329 1311
rect -295 1277 -262 1311
rect -362 1243 -262 1277
rect -362 1209 -329 1243
rect -295 1209 -262 1243
rect -362 1175 -262 1209
rect -362 1141 -329 1175
rect -295 1141 -262 1175
rect -362 1107 -262 1141
rect -362 1073 -329 1107
rect -295 1073 -262 1107
rect -362 1039 -262 1073
rect -362 1005 -329 1039
rect -295 1005 -262 1039
rect -362 971 -262 1005
rect -362 937 -329 971
rect -295 937 -262 971
rect -362 903 -262 937
rect -362 869 -329 903
rect -295 869 -262 903
rect -362 835 -262 869
rect -362 801 -329 835
rect -295 801 -262 835
rect -362 767 -262 801
rect -362 733 -329 767
rect -295 733 -262 767
rect -362 699 -262 733
rect -362 665 -329 699
rect -295 665 -262 699
rect -362 631 -262 665
rect -362 597 -329 631
rect -295 597 -262 631
rect -362 563 -262 597
rect -362 529 -329 563
rect -295 529 -262 563
rect -362 495 -262 529
rect -362 461 -329 495
rect -295 461 -262 495
rect -362 427 -262 461
rect -362 393 -329 427
rect -295 393 -262 427
rect -362 359 -262 393
rect -362 325 -329 359
rect -295 325 -262 359
rect -362 291 -262 325
rect -362 257 -329 291
rect -295 257 -262 291
rect -362 223 -262 257
rect -362 189 -329 223
rect -295 189 -262 223
rect -362 155 -262 189
rect -362 121 -329 155
rect -295 121 -262 155
rect -362 87 -262 121
rect -362 53 -329 87
rect -295 53 -262 87
rect -362 19 -262 53
rect -362 -15 -329 19
rect -295 -15 -262 19
rect -362 -49 -262 -15
rect -362 -83 -329 -49
rect -295 -83 -262 -49
rect -362 -117 -262 -83
rect -362 -151 -329 -117
rect -295 -151 -262 -117
rect -362 -185 -262 -151
rect -362 -219 -329 -185
rect -295 -219 -262 -185
rect -362 -253 -262 -219
rect -362 -287 -329 -253
rect -295 -287 -262 -253
rect -362 -321 -262 -287
rect -362 -355 -329 -321
rect -295 -355 -262 -321
rect -362 -389 -262 -355
rect -362 -423 -329 -389
rect -295 -423 -262 -389
rect -362 -457 -262 -423
rect -362 -491 -329 -457
rect -295 -491 -262 -457
rect -362 -525 -262 -491
rect -362 -559 -329 -525
rect -295 -559 -262 -525
rect -362 -593 -262 -559
rect -362 -627 -329 -593
rect -295 -627 -262 -593
rect -362 -661 -262 -627
rect -362 -695 -329 -661
rect -295 -695 -262 -661
rect -362 -729 -262 -695
rect -362 -763 -329 -729
rect -295 -763 -262 -729
rect -362 -797 -262 -763
rect -362 -831 -329 -797
rect -295 -831 -262 -797
rect -362 -865 -262 -831
rect -362 -899 -329 -865
rect -295 -899 -262 -865
rect -362 -933 -262 -899
rect -362 -967 -329 -933
rect -295 -967 -262 -933
rect -362 -1001 -262 -967
rect -362 -1035 -329 -1001
rect -295 -1035 -262 -1001
rect -362 -1069 -262 -1035
rect -362 -1103 -329 -1069
rect -295 -1103 -262 -1069
rect -362 -1137 -262 -1103
rect -362 -1171 -329 -1137
rect -295 -1171 -262 -1137
rect -362 -1205 -262 -1171
rect -362 -1239 -329 -1205
rect -295 -1239 -262 -1205
rect -362 -1273 -262 -1239
rect -362 -1307 -329 -1273
rect -295 -1307 -262 -1273
rect -362 -1341 -262 -1307
rect -362 -1375 -329 -1341
rect -295 -1375 -262 -1341
rect -362 -1409 -262 -1375
rect -362 -1443 -329 -1409
rect -295 -1443 -262 -1409
rect -362 -1477 -262 -1443
rect -362 -1511 -329 -1477
rect -295 -1511 -262 -1477
rect -362 -1545 -262 -1511
rect -362 -1579 -329 -1545
rect -295 -1579 -262 -1545
rect -362 -1613 -262 -1579
rect -362 -1647 -329 -1613
rect -295 -1647 -262 -1613
rect -362 -1681 -262 -1647
rect -362 -1715 -329 -1681
rect -295 -1715 -262 -1681
rect -362 -1749 -262 -1715
rect -362 -1783 -329 -1749
rect -295 -1783 -262 -1749
rect -362 -1817 -262 -1783
rect -362 -1851 -329 -1817
rect -295 -1851 -262 -1817
rect -362 -1885 -262 -1851
rect -362 -1919 -329 -1885
rect -295 -1919 -262 -1885
rect -362 -1953 -262 -1919
rect -362 -1987 -329 -1953
rect -295 -1987 -262 -1953
rect -362 -2021 -262 -1987
rect -362 -2055 -329 -2021
rect -295 -2055 -262 -2021
rect -362 -2089 -262 -2055
rect -362 -2123 -329 -2089
rect -295 -2123 -262 -2089
rect -362 -2157 -262 -2123
rect -362 -2191 -329 -2157
rect -295 -2191 -262 -2157
rect -362 -2225 -262 -2191
rect -362 -2259 -329 -2225
rect -295 -2259 -262 -2225
rect -362 -2293 -262 -2259
rect -362 -2327 -329 -2293
rect -295 -2327 -262 -2293
rect -362 -2361 -262 -2327
rect -362 -2395 -329 -2361
rect -295 -2395 -262 -2361
rect -362 -2429 -262 -2395
rect -362 -2463 -329 -2429
rect -295 -2463 -262 -2429
rect -362 -2497 -262 -2463
rect -362 -2531 -329 -2497
rect -295 -2531 -262 -2497
rect -362 -2565 -262 -2531
rect -362 -2599 -329 -2565
rect -295 -2599 -262 -2565
rect -362 -2633 -262 -2599
rect -362 -2667 -329 -2633
rect -295 -2667 -262 -2633
rect -362 -2701 -262 -2667
rect -362 -2735 -329 -2701
rect -295 -2735 -262 -2701
rect -362 -2769 -262 -2735
rect -362 -2803 -329 -2769
rect -295 -2803 -262 -2769
rect -362 -2837 -262 -2803
rect -362 -2871 -329 -2837
rect -295 -2871 -262 -2837
rect -362 -2905 -262 -2871
rect -362 -2939 -329 -2905
rect -295 -2939 -262 -2905
rect -362 -2973 -262 -2939
rect -362 -3007 -329 -2973
rect -295 -3007 -262 -2973
rect -362 -3041 -262 -3007
rect -362 -3075 -329 -3041
rect -295 -3075 -262 -3041
rect -362 -3109 -262 -3075
rect -362 -3143 -329 -3109
rect -295 -3143 -262 -3109
rect -362 -3177 -262 -3143
rect -362 -3211 -329 -3177
rect -295 -3211 -262 -3177
rect -362 -3245 -262 -3211
rect -362 -3279 -329 -3245
rect -295 -3279 -262 -3245
rect -362 -3313 -262 -3279
rect -362 -3347 -329 -3313
rect -295 -3347 -262 -3313
rect -362 -3381 -262 -3347
rect -362 -3415 -329 -3381
rect -295 -3415 -262 -3381
rect -362 -3449 -262 -3415
rect -362 -3483 -329 -3449
rect -295 -3483 -262 -3449
rect -362 -3517 -262 -3483
rect -362 -3551 -329 -3517
rect -295 -3551 -262 -3517
rect -362 -3585 -262 -3551
rect -362 -3619 -329 -3585
rect -295 -3619 -262 -3585
rect -362 -3653 -262 -3619
rect -362 -3687 -329 -3653
rect -295 -3687 -262 -3653
rect -362 -3721 -262 -3687
rect -362 -3755 -329 -3721
rect -295 -3755 -262 -3721
rect -362 -3789 -262 -3755
rect -362 -3823 -329 -3789
rect -295 -3823 -262 -3789
rect -362 -3857 -262 -3823
rect -362 -3891 -329 -3857
rect -295 -3891 -262 -3857
rect -362 -3925 -262 -3891
rect -362 -3959 -329 -3925
rect -295 -3959 -262 -3925
rect -362 -3993 -262 -3959
rect -362 -4027 -329 -3993
rect -295 -4027 -262 -3993
rect -362 -4061 -262 -4027
rect -362 -4095 -329 -4061
rect -295 -4095 -262 -4061
rect -362 -4129 -262 -4095
rect -362 -4163 -329 -4129
rect -295 -4163 -262 -4129
rect -362 -4197 -262 -4163
rect -362 -4231 -329 -4197
rect -295 -4231 -262 -4197
rect -362 -4265 -262 -4231
rect -362 -4299 -329 -4265
rect -295 -4299 -262 -4265
rect -362 -4333 -262 -4299
rect -362 -4367 -329 -4333
rect -295 -4367 -262 -4333
rect -362 -4401 -262 -4367
rect -362 -4435 -329 -4401
rect -295 -4435 -262 -4401
rect -362 -4469 -262 -4435
rect -362 -4503 -329 -4469
rect -295 -4503 -262 -4469
rect -362 -4537 -262 -4503
rect -362 -4571 -329 -4537
rect -295 -4571 -262 -4537
rect -362 -4605 -262 -4571
rect -362 -4639 -329 -4605
rect -295 -4639 -262 -4605
rect -362 -4673 -262 -4639
rect -362 -4707 -329 -4673
rect -295 -4707 -262 -4673
rect -362 -4741 -262 -4707
rect -362 -4775 -329 -4741
rect -295 -4775 -262 -4741
rect -362 -4809 -262 -4775
rect -362 -4843 -329 -4809
rect -295 -4843 -262 -4809
rect -362 -4877 -262 -4843
rect -362 -4911 -329 -4877
rect -295 -4911 -262 -4877
rect -362 -4945 -262 -4911
rect -362 -4979 -329 -4945
rect -295 -4979 -262 -4945
rect -362 -5013 -262 -4979
rect -362 -5047 -329 -5013
rect -295 -5047 -262 -5013
rect -362 -5081 -262 -5047
rect -362 -5115 -329 -5081
rect -295 -5115 -262 -5081
rect -362 -5149 -262 -5115
rect -362 -5183 -329 -5149
rect -295 -5183 -262 -5149
rect -362 -5217 -262 -5183
rect -362 -5251 -329 -5217
rect -295 -5251 -262 -5217
rect -362 -5285 -262 -5251
rect -362 -5319 -329 -5285
rect -295 -5319 -262 -5285
rect -362 -5353 -262 -5319
rect -362 -5387 -329 -5353
rect -295 -5387 -262 -5353
rect -362 -5421 -262 -5387
rect -362 -5455 -329 -5421
rect -295 -5455 -262 -5421
rect -362 -5489 -262 -5455
rect -362 -5523 -329 -5489
rect -295 -5523 -262 -5489
rect -362 -5557 -262 -5523
rect -362 -5591 -329 -5557
rect -295 -5591 -262 -5557
rect -362 -5625 -262 -5591
rect -362 -5659 -329 -5625
rect -295 -5659 -262 -5625
rect -362 -5693 -262 -5659
rect -362 -5727 -329 -5693
rect -295 -5727 -262 -5693
rect -362 -5761 -262 -5727
rect -362 -5795 -329 -5761
rect -295 -5795 -262 -5761
rect -362 -5829 -262 -5795
rect -362 -5863 -329 -5829
rect -295 -5863 -262 -5829
rect -362 -5897 -262 -5863
rect -362 -5931 -329 -5897
rect -295 -5931 -262 -5897
rect -362 -5965 -262 -5931
rect -362 -5999 -329 -5965
rect -295 -5999 -262 -5965
rect -362 -6033 -262 -5999
rect -362 -6067 -329 -6033
rect -295 -6067 -262 -6033
rect -362 -6101 -262 -6067
rect -362 -6135 -329 -6101
rect -295 -6135 -262 -6101
rect -362 -6169 -262 -6135
rect -362 -6203 -329 -6169
rect -295 -6203 -262 -6169
rect -362 -6237 -262 -6203
rect -362 -6271 -329 -6237
rect -295 -6271 -262 -6237
rect -362 -6305 -262 -6271
rect -362 -6339 -329 -6305
rect -295 -6339 -262 -6305
rect -362 -6373 -262 -6339
rect -362 -6407 -329 -6373
rect -295 -6407 -262 -6373
rect -362 -6441 -262 -6407
rect -362 -6475 -329 -6441
rect -295 -6475 -262 -6441
rect -362 -6509 -262 -6475
rect -362 -6543 -329 -6509
rect -295 -6543 -262 -6509
rect -362 -6577 -262 -6543
rect -362 -6611 -329 -6577
rect -295 -6611 -262 -6577
rect -362 -6645 -262 -6611
rect -362 -6679 -329 -6645
rect -295 -6679 -262 -6645
rect -362 -6713 -262 -6679
rect -362 -6747 -329 -6713
rect -295 -6747 -262 -6713
rect -362 -6781 -262 -6747
rect -362 -6815 -329 -6781
rect -295 -6815 -262 -6781
rect -362 -6849 -262 -6815
rect -362 -6883 -329 -6849
rect -295 -6883 -262 -6849
rect -362 -6917 -262 -6883
rect -362 -6951 -329 -6917
rect -295 -6951 -262 -6917
rect -362 -6985 -262 -6951
rect -362 -7019 -329 -6985
rect -295 -7019 -262 -6985
rect -362 -7053 -262 -7019
rect -362 -7087 -329 -7053
rect -295 -7087 -262 -7053
rect -362 -7121 -262 -7087
rect -362 -7155 -329 -7121
rect -295 -7155 -262 -7121
rect -362 -7189 -262 -7155
rect -362 -7223 -329 -7189
rect -295 -7223 -262 -7189
rect -362 -7257 -262 -7223
rect -362 -7291 -329 -7257
rect -295 -7291 -262 -7257
rect -362 -7325 -262 -7291
rect -362 -7359 -329 -7325
rect -295 -7359 -262 -7325
rect -362 -7442 -262 -7359
rect 12522 2739 12622 2822
rect 12522 2705 12555 2739
rect 12589 2705 12622 2739
rect 12522 2671 12622 2705
rect 12522 2637 12555 2671
rect 12589 2637 12622 2671
rect 12522 2603 12622 2637
rect 12522 2569 12555 2603
rect 12589 2569 12622 2603
rect 12522 2535 12622 2569
rect 12522 2501 12555 2535
rect 12589 2501 12622 2535
rect 12522 2467 12622 2501
rect 12522 2433 12555 2467
rect 12589 2433 12622 2467
rect 12522 2399 12622 2433
rect 12522 2365 12555 2399
rect 12589 2365 12622 2399
rect 12522 2331 12622 2365
rect 12522 2297 12555 2331
rect 12589 2297 12622 2331
rect 12522 2263 12622 2297
rect 12522 2229 12555 2263
rect 12589 2229 12622 2263
rect 12522 2195 12622 2229
rect 12522 2161 12555 2195
rect 12589 2161 12622 2195
rect 12522 2127 12622 2161
rect 12522 2093 12555 2127
rect 12589 2093 12622 2127
rect 12522 2059 12622 2093
rect 12522 2025 12555 2059
rect 12589 2025 12622 2059
rect 12522 1991 12622 2025
rect 12522 1957 12555 1991
rect 12589 1957 12622 1991
rect 12522 1923 12622 1957
rect 12522 1889 12555 1923
rect 12589 1889 12622 1923
rect 12522 1855 12622 1889
rect 12522 1821 12555 1855
rect 12589 1821 12622 1855
rect 12522 1787 12622 1821
rect 12522 1753 12555 1787
rect 12589 1753 12622 1787
rect 12522 1719 12622 1753
rect 12522 1685 12555 1719
rect 12589 1685 12622 1719
rect 12522 1651 12622 1685
rect 12522 1617 12555 1651
rect 12589 1617 12622 1651
rect 12522 1583 12622 1617
rect 12522 1549 12555 1583
rect 12589 1549 12622 1583
rect 12522 1515 12622 1549
rect 12522 1481 12555 1515
rect 12589 1481 12622 1515
rect 12522 1447 12622 1481
rect 12522 1413 12555 1447
rect 12589 1413 12622 1447
rect 12522 1379 12622 1413
rect 12522 1345 12555 1379
rect 12589 1345 12622 1379
rect 12522 1311 12622 1345
rect 12522 1277 12555 1311
rect 12589 1277 12622 1311
rect 12522 1243 12622 1277
rect 12522 1209 12555 1243
rect 12589 1209 12622 1243
rect 12522 1175 12622 1209
rect 12522 1141 12555 1175
rect 12589 1141 12622 1175
rect 12522 1107 12622 1141
rect 12522 1073 12555 1107
rect 12589 1073 12622 1107
rect 12522 1039 12622 1073
rect 12522 1005 12555 1039
rect 12589 1005 12622 1039
rect 12522 971 12622 1005
rect 12522 937 12555 971
rect 12589 937 12622 971
rect 12522 903 12622 937
rect 12522 869 12555 903
rect 12589 869 12622 903
rect 12522 835 12622 869
rect 12522 801 12555 835
rect 12589 801 12622 835
rect 12522 767 12622 801
rect 12522 733 12555 767
rect 12589 733 12622 767
rect 12522 699 12622 733
rect 12522 665 12555 699
rect 12589 665 12622 699
rect 12522 631 12622 665
rect 12522 597 12555 631
rect 12589 597 12622 631
rect 12522 563 12622 597
rect 12522 529 12555 563
rect 12589 529 12622 563
rect 12522 495 12622 529
rect 12522 461 12555 495
rect 12589 461 12622 495
rect 12522 427 12622 461
rect 12522 393 12555 427
rect 12589 393 12622 427
rect 12522 359 12622 393
rect 12522 325 12555 359
rect 12589 325 12622 359
rect 12522 291 12622 325
rect 12522 257 12555 291
rect 12589 257 12622 291
rect 12522 223 12622 257
rect 12522 189 12555 223
rect 12589 189 12622 223
rect 12522 155 12622 189
rect 12522 121 12555 155
rect 12589 121 12622 155
rect 12522 87 12622 121
rect 12522 53 12555 87
rect 12589 53 12622 87
rect 12522 19 12622 53
rect 12522 -15 12555 19
rect 12589 -15 12622 19
rect 12522 -49 12622 -15
rect 12522 -83 12555 -49
rect 12589 -83 12622 -49
rect 12522 -117 12622 -83
rect 12522 -151 12555 -117
rect 12589 -151 12622 -117
rect 12522 -185 12622 -151
rect 12522 -219 12555 -185
rect 12589 -219 12622 -185
rect 12522 -253 12622 -219
rect 12522 -287 12555 -253
rect 12589 -287 12622 -253
rect 12522 -321 12622 -287
rect 12522 -355 12555 -321
rect 12589 -355 12622 -321
rect 12522 -389 12622 -355
rect 12522 -423 12555 -389
rect 12589 -423 12622 -389
rect 12522 -457 12622 -423
rect 12522 -491 12555 -457
rect 12589 -491 12622 -457
rect 12522 -525 12622 -491
rect 12522 -559 12555 -525
rect 12589 -559 12622 -525
rect 12522 -593 12622 -559
rect 12522 -627 12555 -593
rect 12589 -627 12622 -593
rect 12522 -661 12622 -627
rect 12522 -695 12555 -661
rect 12589 -695 12622 -661
rect 12522 -729 12622 -695
rect 12522 -763 12555 -729
rect 12589 -763 12622 -729
rect 12522 -797 12622 -763
rect 12522 -831 12555 -797
rect 12589 -831 12622 -797
rect 12522 -865 12622 -831
rect 12522 -899 12555 -865
rect 12589 -899 12622 -865
rect 12522 -933 12622 -899
rect 12522 -967 12555 -933
rect 12589 -967 12622 -933
rect 12522 -1001 12622 -967
rect 12522 -1035 12555 -1001
rect 12589 -1035 12622 -1001
rect 12522 -1069 12622 -1035
rect 12522 -1103 12555 -1069
rect 12589 -1103 12622 -1069
rect 12522 -1137 12622 -1103
rect 12522 -1171 12555 -1137
rect 12589 -1171 12622 -1137
rect 12522 -1205 12622 -1171
rect 12522 -1239 12555 -1205
rect 12589 -1239 12622 -1205
rect 12522 -1273 12622 -1239
rect 12522 -1307 12555 -1273
rect 12589 -1307 12622 -1273
rect 12522 -1341 12622 -1307
rect 12522 -1375 12555 -1341
rect 12589 -1375 12622 -1341
rect 12522 -1409 12622 -1375
rect 12522 -1443 12555 -1409
rect 12589 -1443 12622 -1409
rect 12522 -1477 12622 -1443
rect 12522 -1511 12555 -1477
rect 12589 -1511 12622 -1477
rect 12522 -1545 12622 -1511
rect 12522 -1579 12555 -1545
rect 12589 -1579 12622 -1545
rect 12522 -1613 12622 -1579
rect 12522 -1647 12555 -1613
rect 12589 -1647 12622 -1613
rect 12522 -1681 12622 -1647
rect 12522 -1715 12555 -1681
rect 12589 -1715 12622 -1681
rect 12522 -1749 12622 -1715
rect 12522 -1783 12555 -1749
rect 12589 -1783 12622 -1749
rect 12522 -1817 12622 -1783
rect 12522 -1851 12555 -1817
rect 12589 -1851 12622 -1817
rect 12522 -1885 12622 -1851
rect 12522 -1919 12555 -1885
rect 12589 -1919 12622 -1885
rect 12522 -1953 12622 -1919
rect 12522 -1987 12555 -1953
rect 12589 -1987 12622 -1953
rect 12522 -2021 12622 -1987
rect 12522 -2055 12555 -2021
rect 12589 -2055 12622 -2021
rect 12522 -2089 12622 -2055
rect 12522 -2123 12555 -2089
rect 12589 -2123 12622 -2089
rect 12522 -2157 12622 -2123
rect 12522 -2191 12555 -2157
rect 12589 -2191 12622 -2157
rect 12522 -2225 12622 -2191
rect 12522 -2259 12555 -2225
rect 12589 -2259 12622 -2225
rect 12522 -2293 12622 -2259
rect 12522 -2327 12555 -2293
rect 12589 -2327 12622 -2293
rect 12522 -2361 12622 -2327
rect 12522 -2395 12555 -2361
rect 12589 -2395 12622 -2361
rect 12522 -2429 12622 -2395
rect 12522 -2463 12555 -2429
rect 12589 -2463 12622 -2429
rect 12522 -2497 12622 -2463
rect 12522 -2531 12555 -2497
rect 12589 -2531 12622 -2497
rect 12522 -2565 12622 -2531
rect 12522 -2599 12555 -2565
rect 12589 -2599 12622 -2565
rect 12522 -2633 12622 -2599
rect 12522 -2667 12555 -2633
rect 12589 -2667 12622 -2633
rect 12522 -2701 12622 -2667
rect 12522 -2735 12555 -2701
rect 12589 -2735 12622 -2701
rect 12522 -2769 12622 -2735
rect 12522 -2803 12555 -2769
rect 12589 -2803 12622 -2769
rect 12522 -2837 12622 -2803
rect 12522 -2871 12555 -2837
rect 12589 -2871 12622 -2837
rect 12522 -2905 12622 -2871
rect 12522 -2939 12555 -2905
rect 12589 -2939 12622 -2905
rect 12522 -2973 12622 -2939
rect 12522 -3007 12555 -2973
rect 12589 -3007 12622 -2973
rect 12522 -3041 12622 -3007
rect 12522 -3075 12555 -3041
rect 12589 -3075 12622 -3041
rect 12522 -3109 12622 -3075
rect 12522 -3143 12555 -3109
rect 12589 -3143 12622 -3109
rect 12522 -3177 12622 -3143
rect 12522 -3211 12555 -3177
rect 12589 -3211 12622 -3177
rect 12522 -3245 12622 -3211
rect 12522 -3279 12555 -3245
rect 12589 -3279 12622 -3245
rect 12522 -3313 12622 -3279
rect 12522 -3347 12555 -3313
rect 12589 -3347 12622 -3313
rect 12522 -3381 12622 -3347
rect 12522 -3415 12555 -3381
rect 12589 -3415 12622 -3381
rect 12522 -3449 12622 -3415
rect 12522 -3483 12555 -3449
rect 12589 -3483 12622 -3449
rect 12522 -3517 12622 -3483
rect 12522 -3551 12555 -3517
rect 12589 -3551 12622 -3517
rect 12522 -3585 12622 -3551
rect 12522 -3619 12555 -3585
rect 12589 -3619 12622 -3585
rect 12522 -3653 12622 -3619
rect 12522 -3687 12555 -3653
rect 12589 -3687 12622 -3653
rect 12522 -3721 12622 -3687
rect 12522 -3755 12555 -3721
rect 12589 -3755 12622 -3721
rect 12522 -3789 12622 -3755
rect 12522 -3823 12555 -3789
rect 12589 -3823 12622 -3789
rect 12522 -3857 12622 -3823
rect 12522 -3891 12555 -3857
rect 12589 -3891 12622 -3857
rect 12522 -3925 12622 -3891
rect 12522 -3959 12555 -3925
rect 12589 -3959 12622 -3925
rect 12522 -3993 12622 -3959
rect 12522 -4027 12555 -3993
rect 12589 -4027 12622 -3993
rect 12522 -4061 12622 -4027
rect 12522 -4095 12555 -4061
rect 12589 -4095 12622 -4061
rect 12522 -4129 12622 -4095
rect 12522 -4163 12555 -4129
rect 12589 -4163 12622 -4129
rect 12522 -4197 12622 -4163
rect 12522 -4231 12555 -4197
rect 12589 -4231 12622 -4197
rect 12522 -4265 12622 -4231
rect 12522 -4299 12555 -4265
rect 12589 -4299 12622 -4265
rect 12522 -4333 12622 -4299
rect 12522 -4367 12555 -4333
rect 12589 -4367 12622 -4333
rect 12522 -4401 12622 -4367
rect 12522 -4435 12555 -4401
rect 12589 -4435 12622 -4401
rect 12522 -4469 12622 -4435
rect 12522 -4503 12555 -4469
rect 12589 -4503 12622 -4469
rect 12522 -4537 12622 -4503
rect 12522 -4571 12555 -4537
rect 12589 -4571 12622 -4537
rect 12522 -4605 12622 -4571
rect 12522 -4639 12555 -4605
rect 12589 -4639 12622 -4605
rect 12522 -4673 12622 -4639
rect 12522 -4707 12555 -4673
rect 12589 -4707 12622 -4673
rect 12522 -4741 12622 -4707
rect 12522 -4775 12555 -4741
rect 12589 -4775 12622 -4741
rect 12522 -4809 12622 -4775
rect 12522 -4843 12555 -4809
rect 12589 -4843 12622 -4809
rect 12522 -4877 12622 -4843
rect 12522 -4911 12555 -4877
rect 12589 -4911 12622 -4877
rect 12522 -4945 12622 -4911
rect 12522 -4979 12555 -4945
rect 12589 -4979 12622 -4945
rect 12522 -5013 12622 -4979
rect 12522 -5047 12555 -5013
rect 12589 -5047 12622 -5013
rect 12522 -5081 12622 -5047
rect 12522 -5115 12555 -5081
rect 12589 -5115 12622 -5081
rect 12522 -5149 12622 -5115
rect 12522 -5183 12555 -5149
rect 12589 -5183 12622 -5149
rect 12522 -5217 12622 -5183
rect 12522 -5251 12555 -5217
rect 12589 -5251 12622 -5217
rect 12522 -5285 12622 -5251
rect 12522 -5319 12555 -5285
rect 12589 -5319 12622 -5285
rect 12522 -5353 12622 -5319
rect 12522 -5387 12555 -5353
rect 12589 -5387 12622 -5353
rect 12522 -5421 12622 -5387
rect 12522 -5455 12555 -5421
rect 12589 -5455 12622 -5421
rect 12522 -5489 12622 -5455
rect 12522 -5523 12555 -5489
rect 12589 -5523 12622 -5489
rect 12522 -5557 12622 -5523
rect 12522 -5591 12555 -5557
rect 12589 -5591 12622 -5557
rect 12522 -5625 12622 -5591
rect 12522 -5659 12555 -5625
rect 12589 -5659 12622 -5625
rect 12522 -5693 12622 -5659
rect 12522 -5727 12555 -5693
rect 12589 -5727 12622 -5693
rect 12522 -5761 12622 -5727
rect 12522 -5795 12555 -5761
rect 12589 -5795 12622 -5761
rect 12522 -5829 12622 -5795
rect 12522 -5863 12555 -5829
rect 12589 -5863 12622 -5829
rect 12522 -5897 12622 -5863
rect 12522 -5931 12555 -5897
rect 12589 -5931 12622 -5897
rect 12522 -5965 12622 -5931
rect 12522 -5999 12555 -5965
rect 12589 -5999 12622 -5965
rect 12522 -6033 12622 -5999
rect 12522 -6067 12555 -6033
rect 12589 -6067 12622 -6033
rect 12522 -6101 12622 -6067
rect 12522 -6135 12555 -6101
rect 12589 -6135 12622 -6101
rect 12522 -6169 12622 -6135
rect 12522 -6203 12555 -6169
rect 12589 -6203 12622 -6169
rect 12522 -6237 12622 -6203
rect 12522 -6271 12555 -6237
rect 12589 -6271 12622 -6237
rect 12522 -6305 12622 -6271
rect 12522 -6339 12555 -6305
rect 12589 -6339 12622 -6305
rect 12522 -6373 12622 -6339
rect 12522 -6407 12555 -6373
rect 12589 -6407 12622 -6373
rect 12522 -6441 12622 -6407
rect 12522 -6475 12555 -6441
rect 12589 -6475 12622 -6441
rect 12522 -6509 12622 -6475
rect 12522 -6543 12555 -6509
rect 12589 -6543 12622 -6509
rect 12522 -6577 12622 -6543
rect 12522 -6611 12555 -6577
rect 12589 -6611 12622 -6577
rect 12522 -6645 12622 -6611
rect 12522 -6679 12555 -6645
rect 12589 -6679 12622 -6645
rect 12522 -6713 12622 -6679
rect 12522 -6747 12555 -6713
rect 12589 -6747 12622 -6713
rect 12522 -6781 12622 -6747
rect 12522 -6815 12555 -6781
rect 12589 -6815 12622 -6781
rect 12522 -6849 12622 -6815
rect 12522 -6883 12555 -6849
rect 12589 -6883 12622 -6849
rect 12522 -6917 12622 -6883
rect 12522 -6951 12555 -6917
rect 12589 -6951 12622 -6917
rect 12522 -6985 12622 -6951
rect 12522 -7019 12555 -6985
rect 12589 -7019 12622 -6985
rect 12522 -7053 12622 -7019
rect 12522 -7087 12555 -7053
rect 12589 -7087 12622 -7053
rect 12522 -7121 12622 -7087
rect 12522 -7155 12555 -7121
rect 12589 -7155 12622 -7121
rect 12522 -7189 12622 -7155
rect 12522 -7223 12555 -7189
rect 12589 -7223 12622 -7189
rect 12522 -7257 12622 -7223
rect 12522 -7291 12555 -7257
rect 12589 -7291 12622 -7257
rect 12522 -7325 12622 -7291
rect 12522 -7359 12555 -7325
rect 12589 -7359 12622 -7325
rect 12522 -7442 12622 -7359
rect -362 -7475 12622 -7442
rect -362 -7509 -177 -7475
rect -143 -7509 -109 -7475
rect -75 -7509 -41 -7475
rect -7 -7509 27 -7475
rect 61 -7509 95 -7475
rect 129 -7509 163 -7475
rect 197 -7509 231 -7475
rect 265 -7509 299 -7475
rect 333 -7509 367 -7475
rect 401 -7509 435 -7475
rect 469 -7509 503 -7475
rect 537 -7509 571 -7475
rect 605 -7509 639 -7475
rect 673 -7509 707 -7475
rect 741 -7509 775 -7475
rect 809 -7509 843 -7475
rect 877 -7509 911 -7475
rect 945 -7509 979 -7475
rect 1013 -7509 1047 -7475
rect 1081 -7509 1115 -7475
rect 1149 -7509 1183 -7475
rect 1217 -7509 1251 -7475
rect 1285 -7509 1319 -7475
rect 1353 -7509 1387 -7475
rect 1421 -7509 1455 -7475
rect 1489 -7509 1523 -7475
rect 1557 -7509 1591 -7475
rect 1625 -7509 1659 -7475
rect 1693 -7509 1727 -7475
rect 1761 -7509 1795 -7475
rect 1829 -7509 1863 -7475
rect 1897 -7509 1931 -7475
rect 1965 -7509 1999 -7475
rect 2033 -7509 2067 -7475
rect 2101 -7509 2135 -7475
rect 2169 -7509 2203 -7475
rect 2237 -7509 2271 -7475
rect 2305 -7509 2339 -7475
rect 2373 -7509 2407 -7475
rect 2441 -7509 2475 -7475
rect 2509 -7509 2543 -7475
rect 2577 -7509 2611 -7475
rect 2645 -7509 2679 -7475
rect 2713 -7509 2747 -7475
rect 2781 -7509 2815 -7475
rect 2849 -7509 2883 -7475
rect 2917 -7509 2951 -7475
rect 2985 -7509 3019 -7475
rect 3053 -7509 3087 -7475
rect 3121 -7509 3155 -7475
rect 3189 -7509 3223 -7475
rect 3257 -7509 3291 -7475
rect 3325 -7509 3359 -7475
rect 3393 -7509 3427 -7475
rect 3461 -7509 3495 -7475
rect 3529 -7509 3563 -7475
rect 3597 -7509 3631 -7475
rect 3665 -7509 3699 -7475
rect 3733 -7509 3767 -7475
rect 3801 -7509 3835 -7475
rect 3869 -7509 3903 -7475
rect 3937 -7509 3971 -7475
rect 4005 -7509 4039 -7475
rect 4073 -7509 4107 -7475
rect 4141 -7509 4175 -7475
rect 4209 -7509 4243 -7475
rect 4277 -7509 4311 -7475
rect 4345 -7509 4379 -7475
rect 4413 -7509 4447 -7475
rect 4481 -7509 4515 -7475
rect 4549 -7509 4583 -7475
rect 4617 -7509 4651 -7475
rect 4685 -7509 4719 -7475
rect 4753 -7509 4787 -7475
rect 4821 -7509 4855 -7475
rect 4889 -7509 4923 -7475
rect 4957 -7509 4991 -7475
rect 5025 -7509 5059 -7475
rect 5093 -7509 5127 -7475
rect 5161 -7509 5195 -7475
rect 5229 -7509 5263 -7475
rect 5297 -7509 5331 -7475
rect 5365 -7509 5399 -7475
rect 5433 -7509 5467 -7475
rect 5501 -7509 5535 -7475
rect 5569 -7509 5603 -7475
rect 5637 -7509 5671 -7475
rect 5705 -7509 5739 -7475
rect 5773 -7509 5807 -7475
rect 5841 -7509 5875 -7475
rect 5909 -7509 5943 -7475
rect 5977 -7509 6011 -7475
rect 6045 -7509 6079 -7475
rect 6113 -7509 6147 -7475
rect 6181 -7509 6215 -7475
rect 6249 -7509 6283 -7475
rect 6317 -7509 6351 -7475
rect 6385 -7509 6419 -7475
rect 6453 -7509 6487 -7475
rect 6521 -7509 6555 -7475
rect 6589 -7509 6623 -7475
rect 6657 -7509 6691 -7475
rect 6725 -7509 6759 -7475
rect 6793 -7509 6827 -7475
rect 6861 -7509 6895 -7475
rect 6929 -7509 6963 -7475
rect 6997 -7509 7031 -7475
rect 7065 -7509 7099 -7475
rect 7133 -7509 7167 -7475
rect 7201 -7509 7235 -7475
rect 7269 -7509 7303 -7475
rect 7337 -7509 7371 -7475
rect 7405 -7509 7439 -7475
rect 7473 -7509 7507 -7475
rect 7541 -7509 7575 -7475
rect 7609 -7509 7643 -7475
rect 7677 -7509 7711 -7475
rect 7745 -7509 7779 -7475
rect 7813 -7509 7847 -7475
rect 7881 -7509 7915 -7475
rect 7949 -7509 7983 -7475
rect 8017 -7509 8051 -7475
rect 8085 -7509 8119 -7475
rect 8153 -7509 8187 -7475
rect 8221 -7509 8255 -7475
rect 8289 -7509 8323 -7475
rect 8357 -7509 8391 -7475
rect 8425 -7509 8459 -7475
rect 8493 -7509 8527 -7475
rect 8561 -7509 8595 -7475
rect 8629 -7509 8663 -7475
rect 8697 -7509 8731 -7475
rect 8765 -7509 8799 -7475
rect 8833 -7509 8867 -7475
rect 8901 -7509 8935 -7475
rect 8969 -7509 9003 -7475
rect 9037 -7509 9071 -7475
rect 9105 -7509 9139 -7475
rect 9173 -7509 9207 -7475
rect 9241 -7509 9275 -7475
rect 9309 -7509 9343 -7475
rect 9377 -7509 9411 -7475
rect 9445 -7509 9479 -7475
rect 9513 -7509 9547 -7475
rect 9581 -7509 9615 -7475
rect 9649 -7509 9683 -7475
rect 9717 -7509 9751 -7475
rect 9785 -7509 9819 -7475
rect 9853 -7509 9887 -7475
rect 9921 -7509 9955 -7475
rect 9989 -7509 10023 -7475
rect 10057 -7509 10091 -7475
rect 10125 -7509 10159 -7475
rect 10193 -7509 10227 -7475
rect 10261 -7509 10295 -7475
rect 10329 -7509 10363 -7475
rect 10397 -7509 10431 -7475
rect 10465 -7509 10499 -7475
rect 10533 -7509 10567 -7475
rect 10601 -7509 10635 -7475
rect 10669 -7509 10703 -7475
rect 10737 -7509 10771 -7475
rect 10805 -7509 10839 -7475
rect 10873 -7509 10907 -7475
rect 10941 -7509 10975 -7475
rect 11009 -7509 11043 -7475
rect 11077 -7509 11111 -7475
rect 11145 -7509 11179 -7475
rect 11213 -7509 11247 -7475
rect 11281 -7509 11315 -7475
rect 11349 -7509 11383 -7475
rect 11417 -7509 11451 -7475
rect 11485 -7509 11519 -7475
rect 11553 -7509 11587 -7475
rect 11621 -7509 11655 -7475
rect 11689 -7509 11723 -7475
rect 11757 -7509 11791 -7475
rect 11825 -7509 11859 -7475
rect 11893 -7509 11927 -7475
rect 11961 -7509 11995 -7475
rect 12029 -7509 12063 -7475
rect 12097 -7509 12131 -7475
rect 12165 -7509 12199 -7475
rect 12233 -7509 12267 -7475
rect 12301 -7509 12335 -7475
rect 12369 -7509 12403 -7475
rect 12437 -7509 12622 -7475
rect -362 -7542 12622 -7509
<< psubdiffcont >>
rect -177 -7845 -143 -7811
rect -109 -7845 -75 -7811
rect -41 -7845 -7 -7811
rect 27 -7845 61 -7811
rect 95 -7845 129 -7811
rect 163 -7845 197 -7811
rect 231 -7845 265 -7811
rect 299 -7845 333 -7811
rect 367 -7845 401 -7811
rect 435 -7845 469 -7811
rect 503 -7845 537 -7811
rect 571 -7845 605 -7811
rect 639 -7845 673 -7811
rect 707 -7845 741 -7811
rect 775 -7845 809 -7811
rect 843 -7845 877 -7811
rect 911 -7845 945 -7811
rect 979 -7845 1013 -7811
rect 1047 -7845 1081 -7811
rect 1115 -7845 1149 -7811
rect 1183 -7845 1217 -7811
rect 1251 -7845 1285 -7811
rect 1319 -7845 1353 -7811
rect 1387 -7845 1421 -7811
rect 1455 -7845 1489 -7811
rect 1523 -7845 1557 -7811
rect 1591 -7845 1625 -7811
rect 1659 -7845 1693 -7811
rect 1727 -7845 1761 -7811
rect 1795 -7845 1829 -7811
rect 1863 -7845 1897 -7811
rect 1931 -7845 1965 -7811
rect 1999 -7845 2033 -7811
rect 2067 -7845 2101 -7811
rect 2135 -7845 2169 -7811
rect 2203 -7845 2237 -7811
rect 2271 -7845 2305 -7811
rect 2339 -7845 2373 -7811
rect 2407 -7845 2441 -7811
rect 2475 -7845 2509 -7811
rect 2543 -7845 2577 -7811
rect 2611 -7845 2645 -7811
rect 2679 -7845 2713 -7811
rect 2747 -7845 2781 -7811
rect 2815 -7845 2849 -7811
rect 2883 -7845 2917 -7811
rect 2951 -7845 2985 -7811
rect 3019 -7845 3053 -7811
rect 3087 -7845 3121 -7811
rect 3155 -7845 3189 -7811
rect 3223 -7845 3257 -7811
rect 3291 -7845 3325 -7811
rect 3359 -7845 3393 -7811
rect 3427 -7845 3461 -7811
rect 3495 -7845 3529 -7811
rect 3563 -7845 3597 -7811
rect 3631 -7845 3665 -7811
rect 3699 -7845 3733 -7811
rect 3767 -7845 3801 -7811
rect 3835 -7845 3869 -7811
rect 3903 -7845 3937 -7811
rect 3971 -7845 4005 -7811
rect 4039 -7845 4073 -7811
rect 4107 -7845 4141 -7811
rect 4175 -7845 4209 -7811
rect 4243 -7845 4277 -7811
rect 4311 -7845 4345 -7811
rect 4379 -7845 4413 -7811
rect 4447 -7845 4481 -7811
rect 4515 -7845 4549 -7811
rect 4583 -7845 4617 -7811
rect 4651 -7845 4685 -7811
rect 4719 -7845 4753 -7811
rect 4787 -7845 4821 -7811
rect 4855 -7845 4889 -7811
rect 4923 -7845 4957 -7811
rect 4991 -7845 5025 -7811
rect 5059 -7845 5093 -7811
rect 5127 -7845 5161 -7811
rect 5195 -7845 5229 -7811
rect 5263 -7845 5297 -7811
rect 5331 -7845 5365 -7811
rect 5399 -7845 5433 -7811
rect 5467 -7845 5501 -7811
rect 5535 -7845 5569 -7811
rect 5603 -7845 5637 -7811
rect 5671 -7845 5705 -7811
rect 5739 -7845 5773 -7811
rect 5807 -7845 5841 -7811
rect 5875 -7845 5909 -7811
rect 5943 -7845 5977 -7811
rect 6011 -7845 6045 -7811
rect 6079 -7845 6113 -7811
rect 6147 -7845 6181 -7811
rect 6215 -7845 6249 -7811
rect 6283 -7845 6317 -7811
rect 6351 -7845 6385 -7811
rect 6419 -7845 6453 -7811
rect 6487 -7845 6521 -7811
rect 6555 -7845 6589 -7811
rect 6623 -7845 6657 -7811
rect 6691 -7845 6725 -7811
rect 6759 -7845 6793 -7811
rect 6827 -7845 6861 -7811
rect 6895 -7845 6929 -7811
rect 6963 -7845 6997 -7811
rect 7031 -7845 7065 -7811
rect 7099 -7845 7133 -7811
rect 7167 -7845 7201 -7811
rect 7235 -7845 7269 -7811
rect 7303 -7845 7337 -7811
rect 7371 -7845 7405 -7811
rect 7439 -7845 7473 -7811
rect 7507 -7845 7541 -7811
rect 7575 -7845 7609 -7811
rect 7643 -7845 7677 -7811
rect 7711 -7845 7745 -7811
rect 7779 -7845 7813 -7811
rect 7847 -7845 7881 -7811
rect 7915 -7845 7949 -7811
rect 7983 -7845 8017 -7811
rect 8051 -7845 8085 -7811
rect 8119 -7845 8153 -7811
rect 8187 -7845 8221 -7811
rect 8255 -7845 8289 -7811
rect 8323 -7845 8357 -7811
rect 8391 -7845 8425 -7811
rect 8459 -7845 8493 -7811
rect 8527 -7845 8561 -7811
rect 8595 -7845 8629 -7811
rect 8663 -7845 8697 -7811
rect 8731 -7845 8765 -7811
rect 8799 -7845 8833 -7811
rect 8867 -7845 8901 -7811
rect 8935 -7845 8969 -7811
rect 9003 -7845 9037 -7811
rect 9071 -7845 9105 -7811
rect 9139 -7845 9173 -7811
rect 9207 -7845 9241 -7811
rect 9275 -7845 9309 -7811
rect 9343 -7845 9377 -7811
rect 9411 -7845 9445 -7811
rect 9479 -7845 9513 -7811
rect 9547 -7845 9581 -7811
rect 9615 -7845 9649 -7811
rect 9683 -7845 9717 -7811
rect 9751 -7845 9785 -7811
rect 9819 -7845 9853 -7811
rect 9887 -7845 9921 -7811
rect 9955 -7845 9989 -7811
rect 10023 -7845 10057 -7811
rect 10091 -7845 10125 -7811
rect 10159 -7845 10193 -7811
rect 10227 -7845 10261 -7811
rect 10295 -7845 10329 -7811
rect 10363 -7845 10397 -7811
rect 10431 -7845 10465 -7811
rect 10499 -7845 10533 -7811
rect 10567 -7845 10601 -7811
rect 10635 -7845 10669 -7811
rect 10703 -7845 10737 -7811
rect 10771 -7845 10805 -7811
rect 10839 -7845 10873 -7811
rect 10907 -7845 10941 -7811
rect 10975 -7845 11009 -7811
rect 11043 -7845 11077 -7811
rect 11111 -7845 11145 -7811
rect 11179 -7845 11213 -7811
rect 11247 -7845 11281 -7811
rect 11315 -7845 11349 -7811
rect 11383 -7845 11417 -7811
rect 11451 -7845 11485 -7811
rect 11519 -7845 11553 -7811
rect 11587 -7845 11621 -7811
rect 11655 -7845 11689 -7811
rect 11723 -7845 11757 -7811
rect 11791 -7845 11825 -7811
rect 11859 -7845 11893 -7811
rect 11927 -7845 11961 -7811
rect 11995 -7845 12029 -7811
rect 12063 -7845 12097 -7811
rect 12131 -7845 12165 -7811
rect 12199 -7845 12233 -7811
rect 12267 -7845 12301 -7811
rect 12335 -7845 12369 -7811
rect 12403 -7845 12437 -7811
rect -329 -7991 -295 -7957
rect -329 -8059 -295 -8025
rect -329 -8127 -295 -8093
rect -329 -8195 -295 -8161
rect -329 -8263 -295 -8229
rect -329 -8331 -295 -8297
rect -329 -8399 -295 -8365
rect -329 -8467 -295 -8433
rect -329 -8535 -295 -8501
rect -329 -8603 -295 -8569
rect -329 -8671 -295 -8637
rect -329 -8739 -295 -8705
rect -329 -8807 -295 -8773
rect -329 -8875 -295 -8841
rect -329 -8943 -295 -8909
rect -329 -9011 -295 -8977
rect -329 -9079 -295 -9045
rect -329 -9147 -295 -9113
rect -329 -9215 -295 -9181
rect -329 -9283 -295 -9249
rect -329 -9351 -295 -9317
rect -329 -9419 -295 -9385
rect -329 -9487 -295 -9453
rect -329 -9555 -295 -9521
rect -329 -9623 -295 -9589
rect -329 -9691 -295 -9657
rect -329 -9759 -295 -9725
rect -329 -9827 -295 -9793
rect -329 -9895 -295 -9861
rect -329 -9963 -295 -9929
rect -329 -10031 -295 -9997
rect -329 -10099 -295 -10065
rect -329 -10167 -295 -10133
rect -329 -10235 -295 -10201
rect -329 -10303 -295 -10269
rect -329 -10371 -295 -10337
rect -329 -10439 -295 -10405
rect -329 -10507 -295 -10473
rect -329 -10575 -295 -10541
rect -329 -10643 -295 -10609
rect 12555 -7991 12589 -7957
rect 12555 -8059 12589 -8025
rect 12555 -8127 12589 -8093
rect 12555 -8195 12589 -8161
rect 12555 -8263 12589 -8229
rect 12555 -8331 12589 -8297
rect 12555 -8399 12589 -8365
rect 12555 -8467 12589 -8433
rect 12555 -8535 12589 -8501
rect 12555 -8603 12589 -8569
rect 12555 -8671 12589 -8637
rect 12555 -8739 12589 -8705
rect 12555 -8807 12589 -8773
rect 12555 -8875 12589 -8841
rect 12555 -8943 12589 -8909
rect 12555 -9011 12589 -8977
rect 12555 -9079 12589 -9045
rect 12555 -9147 12589 -9113
rect 12555 -9215 12589 -9181
rect 12555 -9283 12589 -9249
rect 12555 -9351 12589 -9317
rect 12555 -9419 12589 -9385
rect 12555 -9487 12589 -9453
rect 12555 -9555 12589 -9521
rect 12555 -9623 12589 -9589
rect 12555 -9691 12589 -9657
rect 12555 -9759 12589 -9725
rect 12555 -9827 12589 -9793
rect 12555 -9895 12589 -9861
rect 12555 -9963 12589 -9929
rect 12555 -10031 12589 -9997
rect 12555 -10099 12589 -10065
rect 12555 -10167 12589 -10133
rect 12555 -10235 12589 -10201
rect 12555 -10303 12589 -10269
rect 12555 -10371 12589 -10337
rect 12555 -10439 12589 -10405
rect 12555 -10507 12589 -10473
rect 12555 -10575 12589 -10541
rect 12555 -10643 12589 -10609
rect -177 -10789 -143 -10755
rect -109 -10789 -75 -10755
rect -41 -10789 -7 -10755
rect 27 -10789 61 -10755
rect 95 -10789 129 -10755
rect 163 -10789 197 -10755
rect 231 -10789 265 -10755
rect 299 -10789 333 -10755
rect 367 -10789 401 -10755
rect 435 -10789 469 -10755
rect 503 -10789 537 -10755
rect 571 -10789 605 -10755
rect 639 -10789 673 -10755
rect 707 -10789 741 -10755
rect 775 -10789 809 -10755
rect 843 -10789 877 -10755
rect 911 -10789 945 -10755
rect 979 -10789 1013 -10755
rect 1047 -10789 1081 -10755
rect 1115 -10789 1149 -10755
rect 1183 -10789 1217 -10755
rect 1251 -10789 1285 -10755
rect 1319 -10789 1353 -10755
rect 1387 -10789 1421 -10755
rect 1455 -10789 1489 -10755
rect 1523 -10789 1557 -10755
rect 1591 -10789 1625 -10755
rect 1659 -10789 1693 -10755
rect 1727 -10789 1761 -10755
rect 1795 -10789 1829 -10755
rect 1863 -10789 1897 -10755
rect 1931 -10789 1965 -10755
rect 1999 -10789 2033 -10755
rect 2067 -10789 2101 -10755
rect 2135 -10789 2169 -10755
rect 2203 -10789 2237 -10755
rect 2271 -10789 2305 -10755
rect 2339 -10789 2373 -10755
rect 2407 -10789 2441 -10755
rect 2475 -10789 2509 -10755
rect 2543 -10789 2577 -10755
rect 2611 -10789 2645 -10755
rect 2679 -10789 2713 -10755
rect 2747 -10789 2781 -10755
rect 2815 -10789 2849 -10755
rect 2883 -10789 2917 -10755
rect 2951 -10789 2985 -10755
rect 3019 -10789 3053 -10755
rect 3087 -10789 3121 -10755
rect 3155 -10789 3189 -10755
rect 3223 -10789 3257 -10755
rect 3291 -10789 3325 -10755
rect 3359 -10789 3393 -10755
rect 3427 -10789 3461 -10755
rect 3495 -10789 3529 -10755
rect 3563 -10789 3597 -10755
rect 3631 -10789 3665 -10755
rect 3699 -10789 3733 -10755
rect 3767 -10789 3801 -10755
rect 3835 -10789 3869 -10755
rect 3903 -10789 3937 -10755
rect 3971 -10789 4005 -10755
rect 4039 -10789 4073 -10755
rect 4107 -10789 4141 -10755
rect 4175 -10789 4209 -10755
rect 4243 -10789 4277 -10755
rect 4311 -10789 4345 -10755
rect 4379 -10789 4413 -10755
rect 4447 -10789 4481 -10755
rect 4515 -10789 4549 -10755
rect 4583 -10789 4617 -10755
rect 4651 -10789 4685 -10755
rect 4719 -10789 4753 -10755
rect 4787 -10789 4821 -10755
rect 4855 -10789 4889 -10755
rect 4923 -10789 4957 -10755
rect 4991 -10789 5025 -10755
rect 5059 -10789 5093 -10755
rect 5127 -10789 5161 -10755
rect 5195 -10789 5229 -10755
rect 5263 -10789 5297 -10755
rect 5331 -10789 5365 -10755
rect 5399 -10789 5433 -10755
rect 5467 -10789 5501 -10755
rect 5535 -10789 5569 -10755
rect 5603 -10789 5637 -10755
rect 5671 -10789 5705 -10755
rect 5739 -10789 5773 -10755
rect 5807 -10789 5841 -10755
rect 5875 -10789 5909 -10755
rect 5943 -10789 5977 -10755
rect 6011 -10789 6045 -10755
rect 6079 -10789 6113 -10755
rect 6147 -10789 6181 -10755
rect 6215 -10789 6249 -10755
rect 6283 -10789 6317 -10755
rect 6351 -10789 6385 -10755
rect 6419 -10789 6453 -10755
rect 6487 -10789 6521 -10755
rect 6555 -10789 6589 -10755
rect 6623 -10789 6657 -10755
rect 6691 -10789 6725 -10755
rect 6759 -10789 6793 -10755
rect 6827 -10789 6861 -10755
rect 6895 -10789 6929 -10755
rect 6963 -10789 6997 -10755
rect 7031 -10789 7065 -10755
rect 7099 -10789 7133 -10755
rect 7167 -10789 7201 -10755
rect 7235 -10789 7269 -10755
rect 7303 -10789 7337 -10755
rect 7371 -10789 7405 -10755
rect 7439 -10789 7473 -10755
rect 7507 -10789 7541 -10755
rect 7575 -10789 7609 -10755
rect 7643 -10789 7677 -10755
rect 7711 -10789 7745 -10755
rect 7779 -10789 7813 -10755
rect 7847 -10789 7881 -10755
rect 7915 -10789 7949 -10755
rect 7983 -10789 8017 -10755
rect 8051 -10789 8085 -10755
rect 8119 -10789 8153 -10755
rect 8187 -10789 8221 -10755
rect 8255 -10789 8289 -10755
rect 8323 -10789 8357 -10755
rect 8391 -10789 8425 -10755
rect 8459 -10789 8493 -10755
rect 8527 -10789 8561 -10755
rect 8595 -10789 8629 -10755
rect 8663 -10789 8697 -10755
rect 8731 -10789 8765 -10755
rect 8799 -10789 8833 -10755
rect 8867 -10789 8901 -10755
rect 8935 -10789 8969 -10755
rect 9003 -10789 9037 -10755
rect 9071 -10789 9105 -10755
rect 9139 -10789 9173 -10755
rect 9207 -10789 9241 -10755
rect 9275 -10789 9309 -10755
rect 9343 -10789 9377 -10755
rect 9411 -10789 9445 -10755
rect 9479 -10789 9513 -10755
rect 9547 -10789 9581 -10755
rect 9615 -10789 9649 -10755
rect 9683 -10789 9717 -10755
rect 9751 -10789 9785 -10755
rect 9819 -10789 9853 -10755
rect 9887 -10789 9921 -10755
rect 9955 -10789 9989 -10755
rect 10023 -10789 10057 -10755
rect 10091 -10789 10125 -10755
rect 10159 -10789 10193 -10755
rect 10227 -10789 10261 -10755
rect 10295 -10789 10329 -10755
rect 10363 -10789 10397 -10755
rect 10431 -10789 10465 -10755
rect 10499 -10789 10533 -10755
rect 10567 -10789 10601 -10755
rect 10635 -10789 10669 -10755
rect 10703 -10789 10737 -10755
rect 10771 -10789 10805 -10755
rect 10839 -10789 10873 -10755
rect 10907 -10789 10941 -10755
rect 10975 -10789 11009 -10755
rect 11043 -10789 11077 -10755
rect 11111 -10789 11145 -10755
rect 11179 -10789 11213 -10755
rect 11247 -10789 11281 -10755
rect 11315 -10789 11349 -10755
rect 11383 -10789 11417 -10755
rect 11451 -10789 11485 -10755
rect 11519 -10789 11553 -10755
rect 11587 -10789 11621 -10755
rect 11655 -10789 11689 -10755
rect 11723 -10789 11757 -10755
rect 11791 -10789 11825 -10755
rect 11859 -10789 11893 -10755
rect 11927 -10789 11961 -10755
rect 11995 -10789 12029 -10755
rect 12063 -10789 12097 -10755
rect 12131 -10789 12165 -10755
rect 12199 -10789 12233 -10755
rect 12267 -10789 12301 -10755
rect 12335 -10789 12369 -10755
rect 12403 -10789 12437 -10755
<< nsubdiffcont >>
rect -177 2855 -143 2889
rect -109 2855 -75 2889
rect -41 2855 -7 2889
rect 27 2855 61 2889
rect 95 2855 129 2889
rect 163 2855 197 2889
rect 231 2855 265 2889
rect 299 2855 333 2889
rect 367 2855 401 2889
rect 435 2855 469 2889
rect 503 2855 537 2889
rect 571 2855 605 2889
rect 639 2855 673 2889
rect 707 2855 741 2889
rect 775 2855 809 2889
rect 843 2855 877 2889
rect 911 2855 945 2889
rect 979 2855 1013 2889
rect 1047 2855 1081 2889
rect 1115 2855 1149 2889
rect 1183 2855 1217 2889
rect 1251 2855 1285 2889
rect 1319 2855 1353 2889
rect 1387 2855 1421 2889
rect 1455 2855 1489 2889
rect 1523 2855 1557 2889
rect 1591 2855 1625 2889
rect 1659 2855 1693 2889
rect 1727 2855 1761 2889
rect 1795 2855 1829 2889
rect 1863 2855 1897 2889
rect 1931 2855 1965 2889
rect 1999 2855 2033 2889
rect 2067 2855 2101 2889
rect 2135 2855 2169 2889
rect 2203 2855 2237 2889
rect 2271 2855 2305 2889
rect 2339 2855 2373 2889
rect 2407 2855 2441 2889
rect 2475 2855 2509 2889
rect 2543 2855 2577 2889
rect 2611 2855 2645 2889
rect 2679 2855 2713 2889
rect 2747 2855 2781 2889
rect 2815 2855 2849 2889
rect 2883 2855 2917 2889
rect 2951 2855 2985 2889
rect 3019 2855 3053 2889
rect 3087 2855 3121 2889
rect 3155 2855 3189 2889
rect 3223 2855 3257 2889
rect 3291 2855 3325 2889
rect 3359 2855 3393 2889
rect 3427 2855 3461 2889
rect 3495 2855 3529 2889
rect 3563 2855 3597 2889
rect 3631 2855 3665 2889
rect 3699 2855 3733 2889
rect 3767 2855 3801 2889
rect 3835 2855 3869 2889
rect 3903 2855 3937 2889
rect 3971 2855 4005 2889
rect 4039 2855 4073 2889
rect 4107 2855 4141 2889
rect 4175 2855 4209 2889
rect 4243 2855 4277 2889
rect 4311 2855 4345 2889
rect 4379 2855 4413 2889
rect 4447 2855 4481 2889
rect 4515 2855 4549 2889
rect 4583 2855 4617 2889
rect 4651 2855 4685 2889
rect 4719 2855 4753 2889
rect 4787 2855 4821 2889
rect 4855 2855 4889 2889
rect 4923 2855 4957 2889
rect 4991 2855 5025 2889
rect 5059 2855 5093 2889
rect 5127 2855 5161 2889
rect 5195 2855 5229 2889
rect 5263 2855 5297 2889
rect 5331 2855 5365 2889
rect 5399 2855 5433 2889
rect 5467 2855 5501 2889
rect 5535 2855 5569 2889
rect 5603 2855 5637 2889
rect 5671 2855 5705 2889
rect 5739 2855 5773 2889
rect 5807 2855 5841 2889
rect 5875 2855 5909 2889
rect 5943 2855 5977 2889
rect 6011 2855 6045 2889
rect 6079 2855 6113 2889
rect 6147 2855 6181 2889
rect 6215 2855 6249 2889
rect 6283 2855 6317 2889
rect 6351 2855 6385 2889
rect 6419 2855 6453 2889
rect 6487 2855 6521 2889
rect 6555 2855 6589 2889
rect 6623 2855 6657 2889
rect 6691 2855 6725 2889
rect 6759 2855 6793 2889
rect 6827 2855 6861 2889
rect 6895 2855 6929 2889
rect 6963 2855 6997 2889
rect 7031 2855 7065 2889
rect 7099 2855 7133 2889
rect 7167 2855 7201 2889
rect 7235 2855 7269 2889
rect 7303 2855 7337 2889
rect 7371 2855 7405 2889
rect 7439 2855 7473 2889
rect 7507 2855 7541 2889
rect 7575 2855 7609 2889
rect 7643 2855 7677 2889
rect 7711 2855 7745 2889
rect 7779 2855 7813 2889
rect 7847 2855 7881 2889
rect 7915 2855 7949 2889
rect 7983 2855 8017 2889
rect 8051 2855 8085 2889
rect 8119 2855 8153 2889
rect 8187 2855 8221 2889
rect 8255 2855 8289 2889
rect 8323 2855 8357 2889
rect 8391 2855 8425 2889
rect 8459 2855 8493 2889
rect 8527 2855 8561 2889
rect 8595 2855 8629 2889
rect 8663 2855 8697 2889
rect 8731 2855 8765 2889
rect 8799 2855 8833 2889
rect 8867 2855 8901 2889
rect 8935 2855 8969 2889
rect 9003 2855 9037 2889
rect 9071 2855 9105 2889
rect 9139 2855 9173 2889
rect 9207 2855 9241 2889
rect 9275 2855 9309 2889
rect 9343 2855 9377 2889
rect 9411 2855 9445 2889
rect 9479 2855 9513 2889
rect 9547 2855 9581 2889
rect 9615 2855 9649 2889
rect 9683 2855 9717 2889
rect 9751 2855 9785 2889
rect 9819 2855 9853 2889
rect 9887 2855 9921 2889
rect 9955 2855 9989 2889
rect 10023 2855 10057 2889
rect 10091 2855 10125 2889
rect 10159 2855 10193 2889
rect 10227 2855 10261 2889
rect 10295 2855 10329 2889
rect 10363 2855 10397 2889
rect 10431 2855 10465 2889
rect 10499 2855 10533 2889
rect 10567 2855 10601 2889
rect 10635 2855 10669 2889
rect 10703 2855 10737 2889
rect 10771 2855 10805 2889
rect 10839 2855 10873 2889
rect 10907 2855 10941 2889
rect 10975 2855 11009 2889
rect 11043 2855 11077 2889
rect 11111 2855 11145 2889
rect 11179 2855 11213 2889
rect 11247 2855 11281 2889
rect 11315 2855 11349 2889
rect 11383 2855 11417 2889
rect 11451 2855 11485 2889
rect 11519 2855 11553 2889
rect 11587 2855 11621 2889
rect 11655 2855 11689 2889
rect 11723 2855 11757 2889
rect 11791 2855 11825 2889
rect 11859 2855 11893 2889
rect 11927 2855 11961 2889
rect 11995 2855 12029 2889
rect 12063 2855 12097 2889
rect 12131 2855 12165 2889
rect 12199 2855 12233 2889
rect 12267 2855 12301 2889
rect 12335 2855 12369 2889
rect 12403 2855 12437 2889
rect -329 2705 -295 2739
rect -329 2637 -295 2671
rect -329 2569 -295 2603
rect -329 2501 -295 2535
rect -329 2433 -295 2467
rect -329 2365 -295 2399
rect -329 2297 -295 2331
rect -329 2229 -295 2263
rect -329 2161 -295 2195
rect -329 2093 -295 2127
rect -329 2025 -295 2059
rect -329 1957 -295 1991
rect -329 1889 -295 1923
rect -329 1821 -295 1855
rect -329 1753 -295 1787
rect -329 1685 -295 1719
rect -329 1617 -295 1651
rect -329 1549 -295 1583
rect -329 1481 -295 1515
rect -329 1413 -295 1447
rect -329 1345 -295 1379
rect -329 1277 -295 1311
rect -329 1209 -295 1243
rect -329 1141 -295 1175
rect -329 1073 -295 1107
rect -329 1005 -295 1039
rect -329 937 -295 971
rect -329 869 -295 903
rect -329 801 -295 835
rect -329 733 -295 767
rect -329 665 -295 699
rect -329 597 -295 631
rect -329 529 -295 563
rect -329 461 -295 495
rect -329 393 -295 427
rect -329 325 -295 359
rect -329 257 -295 291
rect -329 189 -295 223
rect -329 121 -295 155
rect -329 53 -295 87
rect -329 -15 -295 19
rect -329 -83 -295 -49
rect -329 -151 -295 -117
rect -329 -219 -295 -185
rect -329 -287 -295 -253
rect -329 -355 -295 -321
rect -329 -423 -295 -389
rect -329 -491 -295 -457
rect -329 -559 -295 -525
rect -329 -627 -295 -593
rect -329 -695 -295 -661
rect -329 -763 -295 -729
rect -329 -831 -295 -797
rect -329 -899 -295 -865
rect -329 -967 -295 -933
rect -329 -1035 -295 -1001
rect -329 -1103 -295 -1069
rect -329 -1171 -295 -1137
rect -329 -1239 -295 -1205
rect -329 -1307 -295 -1273
rect -329 -1375 -295 -1341
rect -329 -1443 -295 -1409
rect -329 -1511 -295 -1477
rect -329 -1579 -295 -1545
rect -329 -1647 -295 -1613
rect -329 -1715 -295 -1681
rect -329 -1783 -295 -1749
rect -329 -1851 -295 -1817
rect -329 -1919 -295 -1885
rect -329 -1987 -295 -1953
rect -329 -2055 -295 -2021
rect -329 -2123 -295 -2089
rect -329 -2191 -295 -2157
rect -329 -2259 -295 -2225
rect -329 -2327 -295 -2293
rect -329 -2395 -295 -2361
rect -329 -2463 -295 -2429
rect -329 -2531 -295 -2497
rect -329 -2599 -295 -2565
rect -329 -2667 -295 -2633
rect -329 -2735 -295 -2701
rect -329 -2803 -295 -2769
rect -329 -2871 -295 -2837
rect -329 -2939 -295 -2905
rect -329 -3007 -295 -2973
rect -329 -3075 -295 -3041
rect -329 -3143 -295 -3109
rect -329 -3211 -295 -3177
rect -329 -3279 -295 -3245
rect -329 -3347 -295 -3313
rect -329 -3415 -295 -3381
rect -329 -3483 -295 -3449
rect -329 -3551 -295 -3517
rect -329 -3619 -295 -3585
rect -329 -3687 -295 -3653
rect -329 -3755 -295 -3721
rect -329 -3823 -295 -3789
rect -329 -3891 -295 -3857
rect -329 -3959 -295 -3925
rect -329 -4027 -295 -3993
rect -329 -4095 -295 -4061
rect -329 -4163 -295 -4129
rect -329 -4231 -295 -4197
rect -329 -4299 -295 -4265
rect -329 -4367 -295 -4333
rect -329 -4435 -295 -4401
rect -329 -4503 -295 -4469
rect -329 -4571 -295 -4537
rect -329 -4639 -295 -4605
rect -329 -4707 -295 -4673
rect -329 -4775 -295 -4741
rect -329 -4843 -295 -4809
rect -329 -4911 -295 -4877
rect -329 -4979 -295 -4945
rect -329 -5047 -295 -5013
rect -329 -5115 -295 -5081
rect -329 -5183 -295 -5149
rect -329 -5251 -295 -5217
rect -329 -5319 -295 -5285
rect -329 -5387 -295 -5353
rect -329 -5455 -295 -5421
rect -329 -5523 -295 -5489
rect -329 -5591 -295 -5557
rect -329 -5659 -295 -5625
rect -329 -5727 -295 -5693
rect -329 -5795 -295 -5761
rect -329 -5863 -295 -5829
rect -329 -5931 -295 -5897
rect -329 -5999 -295 -5965
rect -329 -6067 -295 -6033
rect -329 -6135 -295 -6101
rect -329 -6203 -295 -6169
rect -329 -6271 -295 -6237
rect -329 -6339 -295 -6305
rect -329 -6407 -295 -6373
rect -329 -6475 -295 -6441
rect -329 -6543 -295 -6509
rect -329 -6611 -295 -6577
rect -329 -6679 -295 -6645
rect -329 -6747 -295 -6713
rect -329 -6815 -295 -6781
rect -329 -6883 -295 -6849
rect -329 -6951 -295 -6917
rect -329 -7019 -295 -6985
rect -329 -7087 -295 -7053
rect -329 -7155 -295 -7121
rect -329 -7223 -295 -7189
rect -329 -7291 -295 -7257
rect -329 -7359 -295 -7325
rect 12555 2705 12589 2739
rect 12555 2637 12589 2671
rect 12555 2569 12589 2603
rect 12555 2501 12589 2535
rect 12555 2433 12589 2467
rect 12555 2365 12589 2399
rect 12555 2297 12589 2331
rect 12555 2229 12589 2263
rect 12555 2161 12589 2195
rect 12555 2093 12589 2127
rect 12555 2025 12589 2059
rect 12555 1957 12589 1991
rect 12555 1889 12589 1923
rect 12555 1821 12589 1855
rect 12555 1753 12589 1787
rect 12555 1685 12589 1719
rect 12555 1617 12589 1651
rect 12555 1549 12589 1583
rect 12555 1481 12589 1515
rect 12555 1413 12589 1447
rect 12555 1345 12589 1379
rect 12555 1277 12589 1311
rect 12555 1209 12589 1243
rect 12555 1141 12589 1175
rect 12555 1073 12589 1107
rect 12555 1005 12589 1039
rect 12555 937 12589 971
rect 12555 869 12589 903
rect 12555 801 12589 835
rect 12555 733 12589 767
rect 12555 665 12589 699
rect 12555 597 12589 631
rect 12555 529 12589 563
rect 12555 461 12589 495
rect 12555 393 12589 427
rect 12555 325 12589 359
rect 12555 257 12589 291
rect 12555 189 12589 223
rect 12555 121 12589 155
rect 12555 53 12589 87
rect 12555 -15 12589 19
rect 12555 -83 12589 -49
rect 12555 -151 12589 -117
rect 12555 -219 12589 -185
rect 12555 -287 12589 -253
rect 12555 -355 12589 -321
rect 12555 -423 12589 -389
rect 12555 -491 12589 -457
rect 12555 -559 12589 -525
rect 12555 -627 12589 -593
rect 12555 -695 12589 -661
rect 12555 -763 12589 -729
rect 12555 -831 12589 -797
rect 12555 -899 12589 -865
rect 12555 -967 12589 -933
rect 12555 -1035 12589 -1001
rect 12555 -1103 12589 -1069
rect 12555 -1171 12589 -1137
rect 12555 -1239 12589 -1205
rect 12555 -1307 12589 -1273
rect 12555 -1375 12589 -1341
rect 12555 -1443 12589 -1409
rect 12555 -1511 12589 -1477
rect 12555 -1579 12589 -1545
rect 12555 -1647 12589 -1613
rect 12555 -1715 12589 -1681
rect 12555 -1783 12589 -1749
rect 12555 -1851 12589 -1817
rect 12555 -1919 12589 -1885
rect 12555 -1987 12589 -1953
rect 12555 -2055 12589 -2021
rect 12555 -2123 12589 -2089
rect 12555 -2191 12589 -2157
rect 12555 -2259 12589 -2225
rect 12555 -2327 12589 -2293
rect 12555 -2395 12589 -2361
rect 12555 -2463 12589 -2429
rect 12555 -2531 12589 -2497
rect 12555 -2599 12589 -2565
rect 12555 -2667 12589 -2633
rect 12555 -2735 12589 -2701
rect 12555 -2803 12589 -2769
rect 12555 -2871 12589 -2837
rect 12555 -2939 12589 -2905
rect 12555 -3007 12589 -2973
rect 12555 -3075 12589 -3041
rect 12555 -3143 12589 -3109
rect 12555 -3211 12589 -3177
rect 12555 -3279 12589 -3245
rect 12555 -3347 12589 -3313
rect 12555 -3415 12589 -3381
rect 12555 -3483 12589 -3449
rect 12555 -3551 12589 -3517
rect 12555 -3619 12589 -3585
rect 12555 -3687 12589 -3653
rect 12555 -3755 12589 -3721
rect 12555 -3823 12589 -3789
rect 12555 -3891 12589 -3857
rect 12555 -3959 12589 -3925
rect 12555 -4027 12589 -3993
rect 12555 -4095 12589 -4061
rect 12555 -4163 12589 -4129
rect 12555 -4231 12589 -4197
rect 12555 -4299 12589 -4265
rect 12555 -4367 12589 -4333
rect 12555 -4435 12589 -4401
rect 12555 -4503 12589 -4469
rect 12555 -4571 12589 -4537
rect 12555 -4639 12589 -4605
rect 12555 -4707 12589 -4673
rect 12555 -4775 12589 -4741
rect 12555 -4843 12589 -4809
rect 12555 -4911 12589 -4877
rect 12555 -4979 12589 -4945
rect 12555 -5047 12589 -5013
rect 12555 -5115 12589 -5081
rect 12555 -5183 12589 -5149
rect 12555 -5251 12589 -5217
rect 12555 -5319 12589 -5285
rect 12555 -5387 12589 -5353
rect 12555 -5455 12589 -5421
rect 12555 -5523 12589 -5489
rect 12555 -5591 12589 -5557
rect 12555 -5659 12589 -5625
rect 12555 -5727 12589 -5693
rect 12555 -5795 12589 -5761
rect 12555 -5863 12589 -5829
rect 12555 -5931 12589 -5897
rect 12555 -5999 12589 -5965
rect 12555 -6067 12589 -6033
rect 12555 -6135 12589 -6101
rect 12555 -6203 12589 -6169
rect 12555 -6271 12589 -6237
rect 12555 -6339 12589 -6305
rect 12555 -6407 12589 -6373
rect 12555 -6475 12589 -6441
rect 12555 -6543 12589 -6509
rect 12555 -6611 12589 -6577
rect 12555 -6679 12589 -6645
rect 12555 -6747 12589 -6713
rect 12555 -6815 12589 -6781
rect 12555 -6883 12589 -6849
rect 12555 -6951 12589 -6917
rect 12555 -7019 12589 -6985
rect 12555 -7087 12589 -7053
rect 12555 -7155 12589 -7121
rect 12555 -7223 12589 -7189
rect 12555 -7291 12589 -7257
rect 12555 -7359 12589 -7325
rect -177 -7509 -143 -7475
rect -109 -7509 -75 -7475
rect -41 -7509 -7 -7475
rect 27 -7509 61 -7475
rect 95 -7509 129 -7475
rect 163 -7509 197 -7475
rect 231 -7509 265 -7475
rect 299 -7509 333 -7475
rect 367 -7509 401 -7475
rect 435 -7509 469 -7475
rect 503 -7509 537 -7475
rect 571 -7509 605 -7475
rect 639 -7509 673 -7475
rect 707 -7509 741 -7475
rect 775 -7509 809 -7475
rect 843 -7509 877 -7475
rect 911 -7509 945 -7475
rect 979 -7509 1013 -7475
rect 1047 -7509 1081 -7475
rect 1115 -7509 1149 -7475
rect 1183 -7509 1217 -7475
rect 1251 -7509 1285 -7475
rect 1319 -7509 1353 -7475
rect 1387 -7509 1421 -7475
rect 1455 -7509 1489 -7475
rect 1523 -7509 1557 -7475
rect 1591 -7509 1625 -7475
rect 1659 -7509 1693 -7475
rect 1727 -7509 1761 -7475
rect 1795 -7509 1829 -7475
rect 1863 -7509 1897 -7475
rect 1931 -7509 1965 -7475
rect 1999 -7509 2033 -7475
rect 2067 -7509 2101 -7475
rect 2135 -7509 2169 -7475
rect 2203 -7509 2237 -7475
rect 2271 -7509 2305 -7475
rect 2339 -7509 2373 -7475
rect 2407 -7509 2441 -7475
rect 2475 -7509 2509 -7475
rect 2543 -7509 2577 -7475
rect 2611 -7509 2645 -7475
rect 2679 -7509 2713 -7475
rect 2747 -7509 2781 -7475
rect 2815 -7509 2849 -7475
rect 2883 -7509 2917 -7475
rect 2951 -7509 2985 -7475
rect 3019 -7509 3053 -7475
rect 3087 -7509 3121 -7475
rect 3155 -7509 3189 -7475
rect 3223 -7509 3257 -7475
rect 3291 -7509 3325 -7475
rect 3359 -7509 3393 -7475
rect 3427 -7509 3461 -7475
rect 3495 -7509 3529 -7475
rect 3563 -7509 3597 -7475
rect 3631 -7509 3665 -7475
rect 3699 -7509 3733 -7475
rect 3767 -7509 3801 -7475
rect 3835 -7509 3869 -7475
rect 3903 -7509 3937 -7475
rect 3971 -7509 4005 -7475
rect 4039 -7509 4073 -7475
rect 4107 -7509 4141 -7475
rect 4175 -7509 4209 -7475
rect 4243 -7509 4277 -7475
rect 4311 -7509 4345 -7475
rect 4379 -7509 4413 -7475
rect 4447 -7509 4481 -7475
rect 4515 -7509 4549 -7475
rect 4583 -7509 4617 -7475
rect 4651 -7509 4685 -7475
rect 4719 -7509 4753 -7475
rect 4787 -7509 4821 -7475
rect 4855 -7509 4889 -7475
rect 4923 -7509 4957 -7475
rect 4991 -7509 5025 -7475
rect 5059 -7509 5093 -7475
rect 5127 -7509 5161 -7475
rect 5195 -7509 5229 -7475
rect 5263 -7509 5297 -7475
rect 5331 -7509 5365 -7475
rect 5399 -7509 5433 -7475
rect 5467 -7509 5501 -7475
rect 5535 -7509 5569 -7475
rect 5603 -7509 5637 -7475
rect 5671 -7509 5705 -7475
rect 5739 -7509 5773 -7475
rect 5807 -7509 5841 -7475
rect 5875 -7509 5909 -7475
rect 5943 -7509 5977 -7475
rect 6011 -7509 6045 -7475
rect 6079 -7509 6113 -7475
rect 6147 -7509 6181 -7475
rect 6215 -7509 6249 -7475
rect 6283 -7509 6317 -7475
rect 6351 -7509 6385 -7475
rect 6419 -7509 6453 -7475
rect 6487 -7509 6521 -7475
rect 6555 -7509 6589 -7475
rect 6623 -7509 6657 -7475
rect 6691 -7509 6725 -7475
rect 6759 -7509 6793 -7475
rect 6827 -7509 6861 -7475
rect 6895 -7509 6929 -7475
rect 6963 -7509 6997 -7475
rect 7031 -7509 7065 -7475
rect 7099 -7509 7133 -7475
rect 7167 -7509 7201 -7475
rect 7235 -7509 7269 -7475
rect 7303 -7509 7337 -7475
rect 7371 -7509 7405 -7475
rect 7439 -7509 7473 -7475
rect 7507 -7509 7541 -7475
rect 7575 -7509 7609 -7475
rect 7643 -7509 7677 -7475
rect 7711 -7509 7745 -7475
rect 7779 -7509 7813 -7475
rect 7847 -7509 7881 -7475
rect 7915 -7509 7949 -7475
rect 7983 -7509 8017 -7475
rect 8051 -7509 8085 -7475
rect 8119 -7509 8153 -7475
rect 8187 -7509 8221 -7475
rect 8255 -7509 8289 -7475
rect 8323 -7509 8357 -7475
rect 8391 -7509 8425 -7475
rect 8459 -7509 8493 -7475
rect 8527 -7509 8561 -7475
rect 8595 -7509 8629 -7475
rect 8663 -7509 8697 -7475
rect 8731 -7509 8765 -7475
rect 8799 -7509 8833 -7475
rect 8867 -7509 8901 -7475
rect 8935 -7509 8969 -7475
rect 9003 -7509 9037 -7475
rect 9071 -7509 9105 -7475
rect 9139 -7509 9173 -7475
rect 9207 -7509 9241 -7475
rect 9275 -7509 9309 -7475
rect 9343 -7509 9377 -7475
rect 9411 -7509 9445 -7475
rect 9479 -7509 9513 -7475
rect 9547 -7509 9581 -7475
rect 9615 -7509 9649 -7475
rect 9683 -7509 9717 -7475
rect 9751 -7509 9785 -7475
rect 9819 -7509 9853 -7475
rect 9887 -7509 9921 -7475
rect 9955 -7509 9989 -7475
rect 10023 -7509 10057 -7475
rect 10091 -7509 10125 -7475
rect 10159 -7509 10193 -7475
rect 10227 -7509 10261 -7475
rect 10295 -7509 10329 -7475
rect 10363 -7509 10397 -7475
rect 10431 -7509 10465 -7475
rect 10499 -7509 10533 -7475
rect 10567 -7509 10601 -7475
rect 10635 -7509 10669 -7475
rect 10703 -7509 10737 -7475
rect 10771 -7509 10805 -7475
rect 10839 -7509 10873 -7475
rect 10907 -7509 10941 -7475
rect 10975 -7509 11009 -7475
rect 11043 -7509 11077 -7475
rect 11111 -7509 11145 -7475
rect 11179 -7509 11213 -7475
rect 11247 -7509 11281 -7475
rect 11315 -7509 11349 -7475
rect 11383 -7509 11417 -7475
rect 11451 -7509 11485 -7475
rect 11519 -7509 11553 -7475
rect 11587 -7509 11621 -7475
rect 11655 -7509 11689 -7475
rect 11723 -7509 11757 -7475
rect 11791 -7509 11825 -7475
rect 11859 -7509 11893 -7475
rect 11927 -7509 11961 -7475
rect 11995 -7509 12029 -7475
rect 12063 -7509 12097 -7475
rect 12131 -7509 12165 -7475
rect 12199 -7509 12233 -7475
rect 12267 -7509 12301 -7475
rect 12335 -7509 12369 -7475
rect 12403 -7509 12437 -7475
<< locali >>
rect -362 2889 12622 2922
rect -362 2855 -259 2889
rect -225 2855 -187 2889
rect -143 2855 -115 2889
rect -75 2855 -43 2889
rect -7 2855 27 2889
rect 63 2855 95 2889
rect 135 2855 163 2889
rect 207 2855 231 2889
rect 279 2855 299 2889
rect 351 2855 367 2889
rect 423 2855 435 2889
rect 495 2855 503 2889
rect 567 2855 571 2889
rect 673 2855 677 2889
rect 741 2855 749 2889
rect 809 2855 821 2889
rect 877 2855 893 2889
rect 945 2855 965 2889
rect 1013 2855 1037 2889
rect 1081 2855 1109 2889
rect 1149 2855 1181 2889
rect 1217 2855 1251 2889
rect 1287 2855 1319 2889
rect 1359 2855 1387 2889
rect 1431 2855 1455 2889
rect 1503 2855 1523 2889
rect 1575 2855 1591 2889
rect 1647 2855 1659 2889
rect 1719 2855 1727 2889
rect 1791 2855 1795 2889
rect 1897 2855 1901 2889
rect 1965 2855 1973 2889
rect 2033 2855 2045 2889
rect 2101 2855 2117 2889
rect 2169 2855 2189 2889
rect 2237 2855 2261 2889
rect 2305 2855 2333 2889
rect 2373 2855 2405 2889
rect 2441 2855 2475 2889
rect 2511 2855 2543 2889
rect 2583 2855 2611 2889
rect 2655 2855 2679 2889
rect 2727 2855 2747 2889
rect 2799 2855 2815 2889
rect 2871 2855 2883 2889
rect 2943 2855 2951 2889
rect 3015 2855 3019 2889
rect 3121 2855 3125 2889
rect 3189 2855 3197 2889
rect 3257 2855 3269 2889
rect 3325 2855 3341 2889
rect 3393 2855 3413 2889
rect 3461 2855 3485 2889
rect 3529 2855 3557 2889
rect 3597 2855 3629 2889
rect 3665 2855 3699 2889
rect 3735 2855 3767 2889
rect 3807 2855 3835 2889
rect 3879 2855 3903 2889
rect 3951 2855 3971 2889
rect 4023 2855 4039 2889
rect 4095 2855 4107 2889
rect 4167 2855 4175 2889
rect 4239 2855 4243 2889
rect 4345 2855 4349 2889
rect 4413 2855 4421 2889
rect 4481 2855 4493 2889
rect 4549 2855 4565 2889
rect 4617 2855 4637 2889
rect 4685 2855 4709 2889
rect 4753 2855 4781 2889
rect 4821 2855 4853 2889
rect 4889 2855 4923 2889
rect 4959 2855 4991 2889
rect 5031 2855 5059 2889
rect 5103 2855 5127 2889
rect 5175 2855 5195 2889
rect 5247 2855 5263 2889
rect 5319 2855 5331 2889
rect 5391 2855 5399 2889
rect 5463 2855 5467 2889
rect 5569 2855 5573 2889
rect 5637 2855 5645 2889
rect 5705 2855 5717 2889
rect 5773 2855 5789 2889
rect 5841 2855 5861 2889
rect 5909 2855 5933 2889
rect 5977 2855 6005 2889
rect 6045 2855 6077 2889
rect 6113 2855 6147 2889
rect 6183 2855 6215 2889
rect 6255 2855 6283 2889
rect 6327 2855 6351 2889
rect 6399 2855 6419 2889
rect 6471 2855 6487 2889
rect 6543 2855 6555 2889
rect 6615 2855 6623 2889
rect 6687 2855 6691 2889
rect 6793 2855 6797 2889
rect 6861 2855 6869 2889
rect 6929 2855 6941 2889
rect 6997 2855 7013 2889
rect 7065 2855 7085 2889
rect 7133 2855 7157 2889
rect 7201 2855 7229 2889
rect 7269 2855 7301 2889
rect 7337 2855 7371 2889
rect 7407 2855 7439 2889
rect 7479 2855 7507 2889
rect 7551 2855 7575 2889
rect 7623 2855 7643 2889
rect 7695 2855 7711 2889
rect 7767 2855 7779 2889
rect 7839 2855 7847 2889
rect 7911 2855 7915 2889
rect 8017 2855 8021 2889
rect 8085 2855 8093 2889
rect 8153 2855 8165 2889
rect 8221 2855 8237 2889
rect 8289 2855 8309 2889
rect 8357 2855 8381 2889
rect 8425 2855 8453 2889
rect 8493 2855 8525 2889
rect 8561 2855 8595 2889
rect 8631 2855 8663 2889
rect 8703 2855 8731 2889
rect 8775 2855 8799 2889
rect 8847 2855 8867 2889
rect 8919 2855 8935 2889
rect 8991 2855 9003 2889
rect 9063 2855 9071 2889
rect 9135 2855 9139 2889
rect 9241 2855 9245 2889
rect 9309 2855 9317 2889
rect 9377 2855 9389 2889
rect 9445 2855 9461 2889
rect 9513 2855 9533 2889
rect 9581 2855 9605 2889
rect 9649 2855 9677 2889
rect 9717 2855 9749 2889
rect 9785 2855 9819 2889
rect 9855 2855 9887 2889
rect 9927 2855 9955 2889
rect 9999 2855 10023 2889
rect 10071 2855 10091 2889
rect 10143 2855 10159 2889
rect 10215 2855 10227 2889
rect 10287 2855 10295 2889
rect 10359 2855 10363 2889
rect 10465 2855 10469 2889
rect 10533 2855 10541 2889
rect 10601 2855 10613 2889
rect 10669 2855 10685 2889
rect 10737 2855 10757 2889
rect 10805 2855 10829 2889
rect 10873 2855 10901 2889
rect 10941 2855 10973 2889
rect 11009 2855 11043 2889
rect 11079 2855 11111 2889
rect 11151 2855 11179 2889
rect 11223 2855 11247 2889
rect 11295 2855 11315 2889
rect 11367 2855 11383 2889
rect 11439 2855 11451 2889
rect 11511 2855 11519 2889
rect 11583 2855 11587 2889
rect 11689 2855 11693 2889
rect 11757 2855 11765 2889
rect 11825 2855 11837 2889
rect 11893 2855 11909 2889
rect 11961 2855 11981 2889
rect 12029 2855 12053 2889
rect 12097 2855 12125 2889
rect 12165 2855 12197 2889
rect 12233 2855 12267 2889
rect 12303 2855 12335 2889
rect 12375 2855 12403 2889
rect 12447 2855 12485 2889
rect 12519 2855 12622 2889
rect -362 2822 12622 2855
rect -362 2739 -262 2822
rect -362 2705 -329 2739
rect -295 2705 -262 2739
rect -362 2671 -262 2705
rect -362 2637 -329 2671
rect -295 2637 -262 2671
rect -362 2603 -262 2637
rect -362 2569 -329 2603
rect -295 2569 -262 2603
rect -362 2535 -262 2569
rect -362 2501 -329 2535
rect -295 2501 -262 2535
rect -362 2467 -262 2501
rect -362 2433 -329 2467
rect -295 2433 -262 2467
rect -362 2399 -262 2433
rect -362 2365 -329 2399
rect -295 2365 -262 2399
rect -362 2331 -262 2365
rect -362 2297 -329 2331
rect -295 2297 -262 2331
rect -362 2287 -262 2297
rect -362 2229 -329 2287
rect -295 2229 -262 2287
rect -362 2215 -262 2229
rect -362 2161 -329 2215
rect -295 2161 -262 2215
rect -362 2143 -262 2161
rect -362 2093 -329 2143
rect -295 2093 -262 2143
rect -362 2071 -262 2093
rect -362 2025 -329 2071
rect -295 2025 -262 2071
rect -362 1999 -262 2025
rect -362 1957 -329 1999
rect -295 1957 -262 1999
rect -362 1927 -262 1957
rect -362 1889 -329 1927
rect -295 1889 -262 1927
rect -362 1855 -262 1889
rect -362 1821 -329 1855
rect -295 1821 -262 1855
rect -362 1787 -262 1821
rect -362 1749 -329 1787
rect -295 1749 -262 1787
rect -362 1719 -262 1749
rect -362 1677 -329 1719
rect -295 1677 -262 1719
rect -362 1651 -262 1677
rect -362 1605 -329 1651
rect -295 1605 -262 1651
rect -362 1583 -262 1605
rect -362 1533 -329 1583
rect -295 1533 -262 1583
rect -362 1515 -262 1533
rect -362 1461 -329 1515
rect -295 1461 -262 1515
rect -362 1447 -262 1461
rect -362 1389 -329 1447
rect -295 1389 -262 1447
rect -362 1379 -262 1389
rect -362 1317 -329 1379
rect -295 1317 -262 1379
rect -362 1311 -262 1317
rect -362 1245 -329 1311
rect -295 1245 -262 1311
rect -362 1243 -262 1245
rect -362 1209 -329 1243
rect -295 1209 -262 1243
rect -362 1207 -262 1209
rect -362 1141 -329 1207
rect -295 1141 -262 1207
rect -362 1135 -262 1141
rect -362 1073 -329 1135
rect -295 1073 -262 1135
rect -362 1063 -262 1073
rect -362 1005 -329 1063
rect -295 1005 -262 1063
rect -362 991 -262 1005
rect -362 937 -329 991
rect -295 937 -262 991
rect -362 919 -262 937
rect -362 869 -329 919
rect -295 869 -262 919
rect -362 847 -262 869
rect -362 801 -329 847
rect -295 801 -262 847
rect -362 775 -262 801
rect -362 733 -329 775
rect -295 733 -262 775
rect -362 703 -262 733
rect -362 665 -329 703
rect -295 665 -262 703
rect -362 631 -262 665
rect -362 597 -329 631
rect -295 597 -262 631
rect -362 563 -262 597
rect -362 525 -329 563
rect -295 525 -262 563
rect -362 495 -262 525
rect -362 453 -329 495
rect -295 453 -262 495
rect -362 427 -262 453
rect -362 381 -329 427
rect -295 381 -262 427
rect -362 359 -262 381
rect -362 309 -329 359
rect -295 309 -262 359
rect -362 291 -262 309
rect -362 237 -329 291
rect -295 237 -262 291
rect -362 223 -262 237
rect -362 165 -329 223
rect -295 165 -262 223
rect -362 155 -262 165
rect -362 93 -329 155
rect -295 93 -262 155
rect -362 87 -262 93
rect -362 21 -329 87
rect -295 21 -262 87
rect -362 19 -262 21
rect -362 -15 -329 19
rect -295 -15 -262 19
rect -362 -17 -262 -15
rect -362 -83 -329 -17
rect -295 -83 -262 -17
rect -362 -89 -262 -83
rect -362 -151 -329 -89
rect -295 -151 -262 -89
rect -362 -161 -262 -151
rect -362 -219 -329 -161
rect -295 -219 -262 -161
rect -362 -233 -262 -219
rect -362 -287 -329 -233
rect -295 -287 -262 -233
rect -362 -305 -262 -287
rect -362 -355 -329 -305
rect -295 -355 -262 -305
rect -362 -377 -262 -355
rect -362 -423 -329 -377
rect -295 -423 -262 -377
rect -362 -449 -262 -423
rect -362 -491 -329 -449
rect -295 -491 -262 -449
rect -362 -521 -262 -491
rect -362 -559 -329 -521
rect -295 -559 -262 -521
rect -362 -593 -262 -559
rect -362 -627 -329 -593
rect -295 -627 -262 -593
rect -362 -661 -262 -627
rect -362 -699 -329 -661
rect -295 -699 -262 -661
rect -362 -729 -262 -699
rect -362 -771 -329 -729
rect -295 -771 -262 -729
rect -362 -797 -262 -771
rect -362 -843 -329 -797
rect -295 -843 -262 -797
rect -362 -865 -262 -843
rect -362 -915 -329 -865
rect -295 -915 -262 -865
rect -362 -933 -262 -915
rect -362 -987 -329 -933
rect -295 -987 -262 -933
rect -362 -1001 -262 -987
rect -362 -1059 -329 -1001
rect -295 -1059 -262 -1001
rect -362 -1069 -262 -1059
rect -362 -1131 -329 -1069
rect -295 -1131 -262 -1069
rect -362 -1137 -262 -1131
rect -362 -1203 -329 -1137
rect -295 -1203 -262 -1137
rect -362 -1205 -262 -1203
rect -362 -1239 -329 -1205
rect -295 -1239 -262 -1205
rect -362 -1241 -262 -1239
rect -362 -1307 -329 -1241
rect -295 -1307 -262 -1241
rect -362 -1313 -262 -1307
rect -362 -1375 -329 -1313
rect -295 -1375 -262 -1313
rect -362 -1385 -262 -1375
rect -362 -1443 -329 -1385
rect -295 -1443 -262 -1385
rect -362 -1457 -262 -1443
rect -362 -1511 -329 -1457
rect -295 -1511 -262 -1457
rect -362 -1529 -262 -1511
rect -362 -1579 -329 -1529
rect -295 -1579 -262 -1529
rect -362 -1601 -262 -1579
rect -362 -1647 -329 -1601
rect -295 -1647 -262 -1601
rect -362 -1673 -262 -1647
rect -362 -1715 -329 -1673
rect -295 -1715 -262 -1673
rect -362 -1745 -262 -1715
rect -362 -1783 -329 -1745
rect -295 -1783 -262 -1745
rect -362 -1817 -262 -1783
rect -362 -1851 -329 -1817
rect -295 -1851 -262 -1817
rect -362 -1885 -262 -1851
rect -362 -1923 -329 -1885
rect -295 -1923 -262 -1885
rect -362 -1953 -262 -1923
rect -362 -1995 -329 -1953
rect -295 -1995 -262 -1953
rect -362 -2021 -262 -1995
rect -362 -2067 -329 -2021
rect -295 -2067 -262 -2021
rect -362 -2089 -262 -2067
rect -362 -2139 -329 -2089
rect -295 -2139 -262 -2089
rect -362 -2157 -262 -2139
rect -362 -2211 -329 -2157
rect -295 -2211 -262 -2157
rect -362 -2225 -262 -2211
rect -362 -2283 -329 -2225
rect -295 -2283 -262 -2225
rect -362 -2293 -262 -2283
rect -362 -2355 -329 -2293
rect -295 -2355 -262 -2293
rect -362 -2361 -262 -2355
rect -362 -2427 -329 -2361
rect -295 -2427 -262 -2361
rect -362 -2429 -262 -2427
rect -362 -2463 -329 -2429
rect -295 -2463 -262 -2429
rect -362 -2465 -262 -2463
rect -362 -2531 -329 -2465
rect -295 -2531 -262 -2465
rect -362 -2537 -262 -2531
rect -362 -2599 -329 -2537
rect -295 -2599 -262 -2537
rect -362 -2609 -262 -2599
rect -362 -2667 -329 -2609
rect -295 -2667 -262 -2609
rect -362 -2681 -262 -2667
rect -362 -2735 -329 -2681
rect -295 -2735 -262 -2681
rect -362 -2753 -262 -2735
rect -362 -2803 -329 -2753
rect -295 -2803 -262 -2753
rect -362 -2825 -262 -2803
rect -362 -2871 -329 -2825
rect -295 -2871 -262 -2825
rect -362 -2897 -262 -2871
rect -362 -2939 -329 -2897
rect -295 -2939 -262 -2897
rect -362 -2969 -262 -2939
rect -362 -3007 -329 -2969
rect -295 -3007 -262 -2969
rect -362 -3041 -262 -3007
rect -362 -3075 -329 -3041
rect -295 -3075 -262 -3041
rect -362 -3109 -262 -3075
rect -362 -3147 -329 -3109
rect -295 -3147 -262 -3109
rect -362 -3177 -262 -3147
rect -362 -3219 -329 -3177
rect -295 -3219 -262 -3177
rect -362 -3245 -262 -3219
rect -362 -3291 -329 -3245
rect -295 -3291 -262 -3245
rect -362 -3313 -262 -3291
rect -362 -3363 -329 -3313
rect -295 -3363 -262 -3313
rect -362 -3381 -262 -3363
rect -362 -3435 -329 -3381
rect -295 -3435 -262 -3381
rect -362 -3449 -262 -3435
rect -362 -3507 -329 -3449
rect -295 -3507 -262 -3449
rect -362 -3517 -262 -3507
rect -362 -3579 -329 -3517
rect -295 -3579 -262 -3517
rect -362 -3585 -262 -3579
rect -362 -3651 -329 -3585
rect -295 -3651 -262 -3585
rect -362 -3653 -262 -3651
rect -362 -3687 -329 -3653
rect -295 -3687 -262 -3653
rect -362 -3689 -262 -3687
rect -362 -3755 -329 -3689
rect -295 -3755 -262 -3689
rect -362 -3761 -262 -3755
rect -362 -3823 -329 -3761
rect -295 -3823 -262 -3761
rect -362 -3833 -262 -3823
rect -362 -3891 -329 -3833
rect -295 -3891 -262 -3833
rect -362 -3905 -262 -3891
rect -362 -3959 -329 -3905
rect -295 -3959 -262 -3905
rect -362 -3977 -262 -3959
rect -362 -4027 -329 -3977
rect -295 -4027 -262 -3977
rect -362 -4049 -262 -4027
rect -362 -4095 -329 -4049
rect -295 -4095 -262 -4049
rect -362 -4121 -262 -4095
rect -362 -4163 -329 -4121
rect -295 -4163 -262 -4121
rect -362 -4193 -262 -4163
rect -362 -4231 -329 -4193
rect -295 -4231 -262 -4193
rect -362 -4265 -262 -4231
rect -362 -4299 -329 -4265
rect -295 -4299 -262 -4265
rect -362 -4333 -262 -4299
rect -362 -4371 -329 -4333
rect -295 -4371 -262 -4333
rect -362 -4401 -262 -4371
rect -362 -4443 -329 -4401
rect -295 -4443 -262 -4401
rect -362 -4469 -262 -4443
rect -362 -4515 -329 -4469
rect -295 -4515 -262 -4469
rect -362 -4537 -262 -4515
rect -362 -4587 -329 -4537
rect -295 -4587 -262 -4537
rect -362 -4605 -262 -4587
rect -362 -4659 -329 -4605
rect -295 -4659 -262 -4605
rect -362 -4673 -262 -4659
rect -362 -4731 -329 -4673
rect -295 -4731 -262 -4673
rect -362 -4741 -262 -4731
rect -362 -4803 -329 -4741
rect -295 -4803 -262 -4741
rect -362 -4809 -262 -4803
rect -362 -4875 -329 -4809
rect -295 -4875 -262 -4809
rect -362 -4877 -262 -4875
rect -362 -4911 -329 -4877
rect -295 -4911 -262 -4877
rect -362 -4913 -262 -4911
rect -362 -4979 -329 -4913
rect -295 -4979 -262 -4913
rect -362 -4985 -262 -4979
rect -362 -5047 -329 -4985
rect -295 -5047 -262 -4985
rect -362 -5057 -262 -5047
rect -362 -5115 -329 -5057
rect -295 -5115 -262 -5057
rect -362 -5129 -262 -5115
rect -362 -5183 -329 -5129
rect -295 -5183 -262 -5129
rect -362 -5201 -262 -5183
rect -362 -5251 -329 -5201
rect -295 -5251 -262 -5201
rect -362 -5273 -262 -5251
rect -362 -5319 -329 -5273
rect -295 -5319 -262 -5273
rect -362 -5345 -262 -5319
rect -362 -5387 -329 -5345
rect -295 -5387 -262 -5345
rect -362 -5417 -262 -5387
rect -362 -5455 -329 -5417
rect -295 -5455 -262 -5417
rect -362 -5489 -262 -5455
rect -362 -5523 -329 -5489
rect -295 -5523 -262 -5489
rect -362 -5557 -262 -5523
rect -362 -5595 -329 -5557
rect -295 -5595 -262 -5557
rect -362 -5625 -262 -5595
rect -362 -5667 -329 -5625
rect -295 -5667 -262 -5625
rect -362 -5693 -262 -5667
rect -362 -5739 -329 -5693
rect -295 -5739 -262 -5693
rect -362 -5761 -262 -5739
rect -362 -5811 -329 -5761
rect -295 -5811 -262 -5761
rect -362 -5829 -262 -5811
rect -362 -5883 -329 -5829
rect -295 -5883 -262 -5829
rect -362 -5897 -262 -5883
rect -362 -5955 -329 -5897
rect -295 -5955 -262 -5897
rect -362 -5965 -262 -5955
rect -362 -6027 -329 -5965
rect -295 -6027 -262 -5965
rect -362 -6033 -262 -6027
rect -362 -6099 -329 -6033
rect -295 -6099 -262 -6033
rect -362 -6101 -262 -6099
rect -362 -6135 -329 -6101
rect -295 -6135 -262 -6101
rect -362 -6137 -262 -6135
rect -362 -6203 -329 -6137
rect -295 -6203 -262 -6137
rect -362 -6209 -262 -6203
rect -362 -6271 -329 -6209
rect -295 -6271 -262 -6209
rect -362 -6281 -262 -6271
rect -362 -6339 -329 -6281
rect -295 -6339 -262 -6281
rect -362 -6353 -262 -6339
rect -362 -6407 -329 -6353
rect -295 -6407 -262 -6353
rect -362 -6425 -262 -6407
rect -362 -6475 -329 -6425
rect -295 -6475 -262 -6425
rect -362 -6497 -262 -6475
rect -362 -6543 -329 -6497
rect -295 -6543 -262 -6497
rect -362 -6569 -262 -6543
rect -362 -6611 -329 -6569
rect -295 -6611 -262 -6569
rect -362 -6641 -262 -6611
rect -362 -6679 -329 -6641
rect -295 -6679 -262 -6641
rect -362 -6713 -262 -6679
rect -362 -6747 -329 -6713
rect -295 -6747 -262 -6713
rect -362 -6781 -262 -6747
rect -362 -6819 -329 -6781
rect -295 -6819 -262 -6781
rect -362 -6849 -262 -6819
rect -362 -6891 -329 -6849
rect -295 -6891 -262 -6849
rect -362 -6917 -262 -6891
rect -362 -6963 -329 -6917
rect -295 -6963 -262 -6917
rect -362 -6985 -262 -6963
rect -362 -7035 -329 -6985
rect -295 -7035 -262 -6985
rect -362 -7053 -262 -7035
rect -362 -7107 -329 -7053
rect -295 -7107 -262 -7053
rect -362 -7121 -262 -7107
rect -362 -7155 -329 -7121
rect -295 -7155 -262 -7121
rect -362 -7189 -262 -7155
rect -362 -7223 -329 -7189
rect -295 -7223 -262 -7189
rect -362 -7257 -262 -7223
rect -362 -7291 -329 -7257
rect -295 -7291 -262 -7257
rect -362 -7325 -262 -7291
rect -362 -7359 -329 -7325
rect -295 -7359 -262 -7325
rect -362 -7442 -262 -7359
rect 12522 2739 12622 2822
rect 12522 2705 12555 2739
rect 12589 2705 12622 2739
rect 12522 2671 12622 2705
rect 12522 2637 12555 2671
rect 12589 2637 12622 2671
rect 12522 2603 12622 2637
rect 12522 2569 12555 2603
rect 12589 2569 12622 2603
rect 12522 2535 12622 2569
rect 12522 2501 12555 2535
rect 12589 2501 12622 2535
rect 12522 2467 12622 2501
rect 12522 2433 12555 2467
rect 12589 2433 12622 2467
rect 12522 2399 12622 2433
rect 12522 2365 12555 2399
rect 12589 2365 12622 2399
rect 12522 2331 12622 2365
rect 12522 2297 12555 2331
rect 12589 2297 12622 2331
rect 12522 2287 12622 2297
rect 12522 2229 12555 2287
rect 12589 2229 12622 2287
rect 12522 2215 12622 2229
rect 12522 2161 12555 2215
rect 12589 2161 12622 2215
rect 12522 2143 12622 2161
rect 12522 2093 12555 2143
rect 12589 2093 12622 2143
rect 12522 2071 12622 2093
rect 12522 2025 12555 2071
rect 12589 2025 12622 2071
rect 12522 1999 12622 2025
rect 12522 1957 12555 1999
rect 12589 1957 12622 1999
rect 12522 1927 12622 1957
rect 12522 1889 12555 1927
rect 12589 1889 12622 1927
rect 12522 1855 12622 1889
rect 12522 1821 12555 1855
rect 12589 1821 12622 1855
rect 12522 1787 12622 1821
rect 12522 1749 12555 1787
rect 12589 1749 12622 1787
rect 12522 1719 12622 1749
rect 12522 1677 12555 1719
rect 12589 1677 12622 1719
rect 12522 1651 12622 1677
rect 12522 1605 12555 1651
rect 12589 1605 12622 1651
rect 12522 1583 12622 1605
rect 12522 1533 12555 1583
rect 12589 1533 12622 1583
rect 12522 1515 12622 1533
rect 12522 1461 12555 1515
rect 12589 1461 12622 1515
rect 12522 1447 12622 1461
rect 12522 1389 12555 1447
rect 12589 1389 12622 1447
rect 12522 1379 12622 1389
rect 12522 1317 12555 1379
rect 12589 1317 12622 1379
rect 12522 1311 12622 1317
rect 12522 1245 12555 1311
rect 12589 1245 12622 1311
rect 12522 1243 12622 1245
rect 12522 1209 12555 1243
rect 12589 1209 12622 1243
rect 12522 1207 12622 1209
rect 12522 1141 12555 1207
rect 12589 1141 12622 1207
rect 12522 1135 12622 1141
rect 12522 1073 12555 1135
rect 12589 1073 12622 1135
rect 12522 1063 12622 1073
rect 12522 1005 12555 1063
rect 12589 1005 12622 1063
rect 12522 991 12622 1005
rect 12522 937 12555 991
rect 12589 937 12622 991
rect 12522 919 12622 937
rect 12522 869 12555 919
rect 12589 869 12622 919
rect 12522 847 12622 869
rect 12522 801 12555 847
rect 12589 801 12622 847
rect 12522 775 12622 801
rect 12522 733 12555 775
rect 12589 733 12622 775
rect 12522 703 12622 733
rect 12522 665 12555 703
rect 12589 665 12622 703
rect 12522 631 12622 665
rect 12522 597 12555 631
rect 12589 597 12622 631
rect 12522 563 12622 597
rect 12522 525 12555 563
rect 12589 525 12622 563
rect 12522 495 12622 525
rect 12522 453 12555 495
rect 12589 453 12622 495
rect 12522 427 12622 453
rect 12522 381 12555 427
rect 12589 381 12622 427
rect 12522 359 12622 381
rect 12522 309 12555 359
rect 12589 309 12622 359
rect 12522 291 12622 309
rect 12522 237 12555 291
rect 12589 237 12622 291
rect 12522 223 12622 237
rect 12522 165 12555 223
rect 12589 165 12622 223
rect 12522 155 12622 165
rect 12522 93 12555 155
rect 12589 93 12622 155
rect 12522 87 12622 93
rect 12522 21 12555 87
rect 12589 21 12622 87
rect 12522 19 12622 21
rect 12522 -15 12555 19
rect 12589 -15 12622 19
rect 12522 -17 12622 -15
rect 12522 -83 12555 -17
rect 12589 -83 12622 -17
rect 12522 -89 12622 -83
rect 12522 -151 12555 -89
rect 12589 -151 12622 -89
rect 12522 -161 12622 -151
rect 12522 -219 12555 -161
rect 12589 -219 12622 -161
rect 12522 -233 12622 -219
rect 12522 -287 12555 -233
rect 12589 -287 12622 -233
rect 12522 -305 12622 -287
rect 12522 -355 12555 -305
rect 12589 -355 12622 -305
rect 12522 -377 12622 -355
rect 12522 -423 12555 -377
rect 12589 -423 12622 -377
rect 12522 -449 12622 -423
rect 12522 -491 12555 -449
rect 12589 -491 12622 -449
rect 12522 -521 12622 -491
rect 12522 -559 12555 -521
rect 12589 -559 12622 -521
rect 12522 -593 12622 -559
rect 12522 -627 12555 -593
rect 12589 -627 12622 -593
rect 12522 -661 12622 -627
rect 12522 -699 12555 -661
rect 12589 -699 12622 -661
rect 12522 -729 12622 -699
rect 12522 -771 12555 -729
rect 12589 -771 12622 -729
rect 12522 -797 12622 -771
rect 12522 -843 12555 -797
rect 12589 -843 12622 -797
rect 12522 -865 12622 -843
rect 12522 -915 12555 -865
rect 12589 -915 12622 -865
rect 12522 -933 12622 -915
rect 12522 -987 12555 -933
rect 12589 -987 12622 -933
rect 12522 -1001 12622 -987
rect 12522 -1059 12555 -1001
rect 12589 -1059 12622 -1001
rect 12522 -1069 12622 -1059
rect 12522 -1131 12555 -1069
rect 12589 -1131 12622 -1069
rect 12522 -1137 12622 -1131
rect 12522 -1203 12555 -1137
rect 12589 -1203 12622 -1137
rect 12522 -1205 12622 -1203
rect 12522 -1239 12555 -1205
rect 12589 -1239 12622 -1205
rect 12522 -1241 12622 -1239
rect 12522 -1307 12555 -1241
rect 12589 -1307 12622 -1241
rect 12522 -1313 12622 -1307
rect 12522 -1375 12555 -1313
rect 12589 -1375 12622 -1313
rect 12522 -1385 12622 -1375
rect 12522 -1443 12555 -1385
rect 12589 -1443 12622 -1385
rect 12522 -1457 12622 -1443
rect 12522 -1511 12555 -1457
rect 12589 -1511 12622 -1457
rect 12522 -1529 12622 -1511
rect 12522 -1579 12555 -1529
rect 12589 -1579 12622 -1529
rect 12522 -1601 12622 -1579
rect 12522 -1647 12555 -1601
rect 12589 -1647 12622 -1601
rect 12522 -1673 12622 -1647
rect 12522 -1715 12555 -1673
rect 12589 -1715 12622 -1673
rect 12522 -1745 12622 -1715
rect 12522 -1783 12555 -1745
rect 12589 -1783 12622 -1745
rect 12522 -1817 12622 -1783
rect 12522 -1851 12555 -1817
rect 12589 -1851 12622 -1817
rect 12522 -1885 12622 -1851
rect 12522 -1923 12555 -1885
rect 12589 -1923 12622 -1885
rect 12522 -1953 12622 -1923
rect 12522 -1995 12555 -1953
rect 12589 -1995 12622 -1953
rect 12522 -2021 12622 -1995
rect 12522 -2067 12555 -2021
rect 12589 -2067 12622 -2021
rect 12522 -2089 12622 -2067
rect 12522 -2139 12555 -2089
rect 12589 -2139 12622 -2089
rect 12522 -2157 12622 -2139
rect 12522 -2211 12555 -2157
rect 12589 -2211 12622 -2157
rect 12522 -2225 12622 -2211
rect 12522 -2283 12555 -2225
rect 12589 -2283 12622 -2225
rect 12522 -2293 12622 -2283
rect 12522 -2355 12555 -2293
rect 12589 -2355 12622 -2293
rect 12522 -2361 12622 -2355
rect 12522 -2427 12555 -2361
rect 12589 -2427 12622 -2361
rect 12522 -2429 12622 -2427
rect 12522 -2463 12555 -2429
rect 12589 -2463 12622 -2429
rect 12522 -2465 12622 -2463
rect 12522 -2531 12555 -2465
rect 12589 -2531 12622 -2465
rect 12522 -2537 12622 -2531
rect 12522 -2599 12555 -2537
rect 12589 -2599 12622 -2537
rect 12522 -2609 12622 -2599
rect 12522 -2667 12555 -2609
rect 12589 -2667 12622 -2609
rect 12522 -2681 12622 -2667
rect 12522 -2735 12555 -2681
rect 12589 -2735 12622 -2681
rect 12522 -2753 12622 -2735
rect 12522 -2803 12555 -2753
rect 12589 -2803 12622 -2753
rect 12522 -2825 12622 -2803
rect 12522 -2871 12555 -2825
rect 12589 -2871 12622 -2825
rect 12522 -2897 12622 -2871
rect 12522 -2939 12555 -2897
rect 12589 -2939 12622 -2897
rect 12522 -2969 12622 -2939
rect 12522 -3007 12555 -2969
rect 12589 -3007 12622 -2969
rect 12522 -3041 12622 -3007
rect 12522 -3075 12555 -3041
rect 12589 -3075 12622 -3041
rect 12522 -3109 12622 -3075
rect 12522 -3147 12555 -3109
rect 12589 -3147 12622 -3109
rect 12522 -3177 12622 -3147
rect 12522 -3219 12555 -3177
rect 12589 -3219 12622 -3177
rect 12522 -3245 12622 -3219
rect 12522 -3291 12555 -3245
rect 12589 -3291 12622 -3245
rect 12522 -3313 12622 -3291
rect 12522 -3363 12555 -3313
rect 12589 -3363 12622 -3313
rect 12522 -3381 12622 -3363
rect 12522 -3435 12555 -3381
rect 12589 -3435 12622 -3381
rect 12522 -3449 12622 -3435
rect 12522 -3507 12555 -3449
rect 12589 -3507 12622 -3449
rect 12522 -3517 12622 -3507
rect 12522 -3579 12555 -3517
rect 12589 -3579 12622 -3517
rect 12522 -3585 12622 -3579
rect 12522 -3651 12555 -3585
rect 12589 -3651 12622 -3585
rect 12522 -3653 12622 -3651
rect 12522 -3687 12555 -3653
rect 12589 -3687 12622 -3653
rect 12522 -3689 12622 -3687
rect 12522 -3755 12555 -3689
rect 12589 -3755 12622 -3689
rect 12522 -3761 12622 -3755
rect 12522 -3823 12555 -3761
rect 12589 -3823 12622 -3761
rect 12522 -3833 12622 -3823
rect 12522 -3891 12555 -3833
rect 12589 -3891 12622 -3833
rect 12522 -3905 12622 -3891
rect 12522 -3959 12555 -3905
rect 12589 -3959 12622 -3905
rect 12522 -3977 12622 -3959
rect 12522 -4027 12555 -3977
rect 12589 -4027 12622 -3977
rect 12522 -4049 12622 -4027
rect 12522 -4095 12555 -4049
rect 12589 -4095 12622 -4049
rect 12522 -4121 12622 -4095
rect 12522 -4163 12555 -4121
rect 12589 -4163 12622 -4121
rect 12522 -4193 12622 -4163
rect 12522 -4231 12555 -4193
rect 12589 -4231 12622 -4193
rect 12522 -4265 12622 -4231
rect 12522 -4299 12555 -4265
rect 12589 -4299 12622 -4265
rect 12522 -4333 12622 -4299
rect 12522 -4371 12555 -4333
rect 12589 -4371 12622 -4333
rect 12522 -4401 12622 -4371
rect 12522 -4443 12555 -4401
rect 12589 -4443 12622 -4401
rect 12522 -4469 12622 -4443
rect 12522 -4515 12555 -4469
rect 12589 -4515 12622 -4469
rect 12522 -4537 12622 -4515
rect 12522 -4587 12555 -4537
rect 12589 -4587 12622 -4537
rect 12522 -4605 12622 -4587
rect 12522 -4659 12555 -4605
rect 12589 -4659 12622 -4605
rect 12522 -4673 12622 -4659
rect 12522 -4731 12555 -4673
rect 12589 -4731 12622 -4673
rect 12522 -4741 12622 -4731
rect 12522 -4803 12555 -4741
rect 12589 -4803 12622 -4741
rect 12522 -4809 12622 -4803
rect 12522 -4875 12555 -4809
rect 12589 -4875 12622 -4809
rect 12522 -4877 12622 -4875
rect 12522 -4911 12555 -4877
rect 12589 -4911 12622 -4877
rect 12522 -4913 12622 -4911
rect 12522 -4979 12555 -4913
rect 12589 -4979 12622 -4913
rect 12522 -4985 12622 -4979
rect 12522 -5047 12555 -4985
rect 12589 -5047 12622 -4985
rect 12522 -5057 12622 -5047
rect 12522 -5115 12555 -5057
rect 12589 -5115 12622 -5057
rect 12522 -5129 12622 -5115
rect 12522 -5183 12555 -5129
rect 12589 -5183 12622 -5129
rect 12522 -5201 12622 -5183
rect 12522 -5251 12555 -5201
rect 12589 -5251 12622 -5201
rect 12522 -5273 12622 -5251
rect 12522 -5319 12555 -5273
rect 12589 -5319 12622 -5273
rect 12522 -5345 12622 -5319
rect 12522 -5387 12555 -5345
rect 12589 -5387 12622 -5345
rect 12522 -5417 12622 -5387
rect 12522 -5455 12555 -5417
rect 12589 -5455 12622 -5417
rect 12522 -5489 12622 -5455
rect 12522 -5523 12555 -5489
rect 12589 -5523 12622 -5489
rect 12522 -5557 12622 -5523
rect 12522 -5595 12555 -5557
rect 12589 -5595 12622 -5557
rect 12522 -5625 12622 -5595
rect 12522 -5667 12555 -5625
rect 12589 -5667 12622 -5625
rect 12522 -5693 12622 -5667
rect 12522 -5739 12555 -5693
rect 12589 -5739 12622 -5693
rect 12522 -5761 12622 -5739
rect 12522 -5811 12555 -5761
rect 12589 -5811 12622 -5761
rect 12522 -5829 12622 -5811
rect 12522 -5883 12555 -5829
rect 12589 -5883 12622 -5829
rect 12522 -5897 12622 -5883
rect 12522 -5955 12555 -5897
rect 12589 -5955 12622 -5897
rect 12522 -5965 12622 -5955
rect 12522 -6027 12555 -5965
rect 12589 -6027 12622 -5965
rect 12522 -6033 12622 -6027
rect 12522 -6099 12555 -6033
rect 12589 -6099 12622 -6033
rect 12522 -6101 12622 -6099
rect 12522 -6135 12555 -6101
rect 12589 -6135 12622 -6101
rect 12522 -6137 12622 -6135
rect 12522 -6203 12555 -6137
rect 12589 -6203 12622 -6137
rect 12522 -6209 12622 -6203
rect 12522 -6271 12555 -6209
rect 12589 -6271 12622 -6209
rect 12522 -6281 12622 -6271
rect 12522 -6339 12555 -6281
rect 12589 -6339 12622 -6281
rect 12522 -6353 12622 -6339
rect 12522 -6407 12555 -6353
rect 12589 -6407 12622 -6353
rect 12522 -6425 12622 -6407
rect 12522 -6475 12555 -6425
rect 12589 -6475 12622 -6425
rect 12522 -6497 12622 -6475
rect 12522 -6543 12555 -6497
rect 12589 -6543 12622 -6497
rect 12522 -6569 12622 -6543
rect 12522 -6611 12555 -6569
rect 12589 -6611 12622 -6569
rect 12522 -6641 12622 -6611
rect 12522 -6679 12555 -6641
rect 12589 -6679 12622 -6641
rect 12522 -6713 12622 -6679
rect 12522 -6747 12555 -6713
rect 12589 -6747 12622 -6713
rect 12522 -6781 12622 -6747
rect 12522 -6819 12555 -6781
rect 12589 -6819 12622 -6781
rect 12522 -6849 12622 -6819
rect 12522 -6891 12555 -6849
rect 12589 -6891 12622 -6849
rect 12522 -6917 12622 -6891
rect 12522 -6963 12555 -6917
rect 12589 -6963 12622 -6917
rect 12522 -6985 12622 -6963
rect 12522 -7035 12555 -6985
rect 12589 -7035 12622 -6985
rect 12522 -7053 12622 -7035
rect 12522 -7107 12555 -7053
rect 12589 -7107 12622 -7053
rect 12522 -7121 12622 -7107
rect 12522 -7155 12555 -7121
rect 12589 -7155 12622 -7121
rect 12522 -7189 12622 -7155
rect 12522 -7223 12555 -7189
rect 12589 -7223 12622 -7189
rect 12522 -7257 12622 -7223
rect 12522 -7291 12555 -7257
rect 12589 -7291 12622 -7257
rect 12522 -7325 12622 -7291
rect 12522 -7359 12555 -7325
rect 12589 -7359 12622 -7325
rect 12522 -7442 12622 -7359
rect -362 -7475 12622 -7442
rect -362 -7509 -259 -7475
rect -225 -7509 -187 -7475
rect -143 -7509 -115 -7475
rect -75 -7509 -43 -7475
rect -7 -7509 27 -7475
rect 63 -7509 95 -7475
rect 135 -7509 163 -7475
rect 207 -7509 231 -7475
rect 279 -7509 299 -7475
rect 351 -7509 367 -7475
rect 423 -7509 435 -7475
rect 495 -7509 503 -7475
rect 567 -7509 571 -7475
rect 673 -7509 677 -7475
rect 741 -7509 749 -7475
rect 809 -7509 821 -7475
rect 877 -7509 893 -7475
rect 945 -7509 965 -7475
rect 1013 -7509 1037 -7475
rect 1081 -7509 1109 -7475
rect 1149 -7509 1181 -7475
rect 1217 -7509 1251 -7475
rect 1287 -7509 1319 -7475
rect 1359 -7509 1387 -7475
rect 1431 -7509 1455 -7475
rect 1503 -7509 1523 -7475
rect 1575 -7509 1591 -7475
rect 1647 -7509 1659 -7475
rect 1719 -7509 1727 -7475
rect 1791 -7509 1795 -7475
rect 1897 -7509 1901 -7475
rect 1965 -7509 1973 -7475
rect 2033 -7509 2045 -7475
rect 2101 -7509 2117 -7475
rect 2169 -7509 2189 -7475
rect 2237 -7509 2261 -7475
rect 2305 -7509 2333 -7475
rect 2373 -7509 2405 -7475
rect 2441 -7509 2475 -7475
rect 2511 -7509 2543 -7475
rect 2583 -7509 2611 -7475
rect 2655 -7509 2679 -7475
rect 2727 -7509 2747 -7475
rect 2799 -7509 2815 -7475
rect 2871 -7509 2883 -7475
rect 2943 -7509 2951 -7475
rect 3015 -7509 3019 -7475
rect 3121 -7509 3125 -7475
rect 3189 -7509 3197 -7475
rect 3257 -7509 3269 -7475
rect 3325 -7509 3341 -7475
rect 3393 -7509 3413 -7475
rect 3461 -7509 3485 -7475
rect 3529 -7509 3557 -7475
rect 3597 -7509 3629 -7475
rect 3665 -7509 3699 -7475
rect 3735 -7509 3767 -7475
rect 3807 -7509 3835 -7475
rect 3879 -7509 3903 -7475
rect 3951 -7509 3971 -7475
rect 4023 -7509 4039 -7475
rect 4095 -7509 4107 -7475
rect 4167 -7509 4175 -7475
rect 4239 -7509 4243 -7475
rect 4345 -7509 4349 -7475
rect 4413 -7509 4421 -7475
rect 4481 -7509 4493 -7475
rect 4549 -7509 4565 -7475
rect 4617 -7509 4637 -7475
rect 4685 -7509 4709 -7475
rect 4753 -7509 4781 -7475
rect 4821 -7509 4853 -7475
rect 4889 -7509 4923 -7475
rect 4959 -7509 4991 -7475
rect 5031 -7509 5059 -7475
rect 5103 -7509 5127 -7475
rect 5175 -7509 5195 -7475
rect 5247 -7509 5263 -7475
rect 5319 -7509 5331 -7475
rect 5391 -7509 5399 -7475
rect 5463 -7509 5467 -7475
rect 5569 -7509 5573 -7475
rect 5637 -7509 5645 -7475
rect 5705 -7509 5717 -7475
rect 5773 -7509 5789 -7475
rect 5841 -7509 5861 -7475
rect 5909 -7509 5933 -7475
rect 5977 -7509 6005 -7475
rect 6045 -7509 6077 -7475
rect 6113 -7509 6147 -7475
rect 6183 -7509 6215 -7475
rect 6255 -7509 6283 -7475
rect 6327 -7509 6351 -7475
rect 6399 -7509 6419 -7475
rect 6471 -7509 6487 -7475
rect 6543 -7509 6555 -7475
rect 6615 -7509 6623 -7475
rect 6687 -7509 6691 -7475
rect 6793 -7509 6797 -7475
rect 6861 -7509 6869 -7475
rect 6929 -7509 6941 -7475
rect 6997 -7509 7013 -7475
rect 7065 -7509 7085 -7475
rect 7133 -7509 7157 -7475
rect 7201 -7509 7229 -7475
rect 7269 -7509 7301 -7475
rect 7337 -7509 7371 -7475
rect 7407 -7509 7439 -7475
rect 7479 -7509 7507 -7475
rect 7551 -7509 7575 -7475
rect 7623 -7509 7643 -7475
rect 7695 -7509 7711 -7475
rect 7767 -7509 7779 -7475
rect 7839 -7509 7847 -7475
rect 7911 -7509 7915 -7475
rect 8017 -7509 8021 -7475
rect 8085 -7509 8093 -7475
rect 8153 -7509 8165 -7475
rect 8221 -7509 8237 -7475
rect 8289 -7509 8309 -7475
rect 8357 -7509 8381 -7475
rect 8425 -7509 8453 -7475
rect 8493 -7509 8525 -7475
rect 8561 -7509 8595 -7475
rect 8631 -7509 8663 -7475
rect 8703 -7509 8731 -7475
rect 8775 -7509 8799 -7475
rect 8847 -7509 8867 -7475
rect 8919 -7509 8935 -7475
rect 8991 -7509 9003 -7475
rect 9063 -7509 9071 -7475
rect 9135 -7509 9139 -7475
rect 9241 -7509 9245 -7475
rect 9309 -7509 9317 -7475
rect 9377 -7509 9389 -7475
rect 9445 -7509 9461 -7475
rect 9513 -7509 9533 -7475
rect 9581 -7509 9605 -7475
rect 9649 -7509 9677 -7475
rect 9717 -7509 9749 -7475
rect 9785 -7509 9819 -7475
rect 9855 -7509 9887 -7475
rect 9927 -7509 9955 -7475
rect 9999 -7509 10023 -7475
rect 10071 -7509 10091 -7475
rect 10143 -7509 10159 -7475
rect 10215 -7509 10227 -7475
rect 10287 -7509 10295 -7475
rect 10359 -7509 10363 -7475
rect 10465 -7509 10469 -7475
rect 10533 -7509 10541 -7475
rect 10601 -7509 10613 -7475
rect 10669 -7509 10685 -7475
rect 10737 -7509 10757 -7475
rect 10805 -7509 10829 -7475
rect 10873 -7509 10901 -7475
rect 10941 -7509 10973 -7475
rect 11009 -7509 11043 -7475
rect 11079 -7509 11111 -7475
rect 11151 -7509 11179 -7475
rect 11223 -7509 11247 -7475
rect 11295 -7509 11315 -7475
rect 11367 -7509 11383 -7475
rect 11439 -7509 11451 -7475
rect 11511 -7509 11519 -7475
rect 11583 -7509 11587 -7475
rect 11689 -7509 11693 -7475
rect 11757 -7509 11765 -7475
rect 11825 -7509 11837 -7475
rect 11893 -7509 11909 -7475
rect 11961 -7509 11981 -7475
rect 12029 -7509 12053 -7475
rect 12097 -7509 12125 -7475
rect 12165 -7509 12197 -7475
rect 12233 -7509 12267 -7475
rect 12303 -7509 12335 -7475
rect 12375 -7509 12403 -7475
rect 12447 -7509 12485 -7475
rect 12519 -7509 12622 -7475
rect -362 -7542 12622 -7509
rect -362 -7811 12622 -7778
rect -362 -7845 -259 -7811
rect -225 -7845 -187 -7811
rect -143 -7845 -115 -7811
rect -75 -7845 -43 -7811
rect -7 -7845 27 -7811
rect 63 -7845 95 -7811
rect 135 -7845 163 -7811
rect 207 -7845 231 -7811
rect 279 -7845 299 -7811
rect 351 -7845 367 -7811
rect 423 -7845 435 -7811
rect 495 -7845 503 -7811
rect 567 -7845 571 -7811
rect 673 -7845 677 -7811
rect 741 -7845 749 -7811
rect 809 -7845 821 -7811
rect 877 -7845 893 -7811
rect 945 -7845 965 -7811
rect 1013 -7845 1037 -7811
rect 1081 -7845 1109 -7811
rect 1149 -7845 1181 -7811
rect 1217 -7845 1251 -7811
rect 1287 -7845 1319 -7811
rect 1359 -7845 1387 -7811
rect 1431 -7845 1455 -7811
rect 1503 -7845 1523 -7811
rect 1575 -7845 1591 -7811
rect 1647 -7845 1659 -7811
rect 1719 -7845 1727 -7811
rect 1791 -7845 1795 -7811
rect 1897 -7845 1901 -7811
rect 1965 -7845 1973 -7811
rect 2033 -7845 2045 -7811
rect 2101 -7845 2117 -7811
rect 2169 -7845 2189 -7811
rect 2237 -7845 2261 -7811
rect 2305 -7845 2333 -7811
rect 2373 -7845 2405 -7811
rect 2441 -7845 2475 -7811
rect 2511 -7845 2543 -7811
rect 2583 -7845 2611 -7811
rect 2655 -7845 2679 -7811
rect 2727 -7845 2747 -7811
rect 2799 -7845 2815 -7811
rect 2871 -7845 2883 -7811
rect 2943 -7845 2951 -7811
rect 3015 -7845 3019 -7811
rect 3121 -7845 3125 -7811
rect 3189 -7845 3197 -7811
rect 3257 -7845 3269 -7811
rect 3325 -7845 3341 -7811
rect 3393 -7845 3413 -7811
rect 3461 -7845 3485 -7811
rect 3529 -7845 3557 -7811
rect 3597 -7845 3629 -7811
rect 3665 -7845 3699 -7811
rect 3735 -7845 3767 -7811
rect 3807 -7845 3835 -7811
rect 3879 -7845 3903 -7811
rect 3951 -7845 3971 -7811
rect 4023 -7845 4039 -7811
rect 4095 -7845 4107 -7811
rect 4167 -7845 4175 -7811
rect 4239 -7845 4243 -7811
rect 4345 -7845 4349 -7811
rect 4413 -7845 4421 -7811
rect 4481 -7845 4493 -7811
rect 4549 -7845 4565 -7811
rect 4617 -7845 4637 -7811
rect 4685 -7845 4709 -7811
rect 4753 -7845 4781 -7811
rect 4821 -7845 4853 -7811
rect 4889 -7845 4923 -7811
rect 4959 -7845 4991 -7811
rect 5031 -7845 5059 -7811
rect 5103 -7845 5127 -7811
rect 5175 -7845 5195 -7811
rect 5247 -7845 5263 -7811
rect 5319 -7845 5331 -7811
rect 5391 -7845 5399 -7811
rect 5463 -7845 5467 -7811
rect 5569 -7845 5573 -7811
rect 5637 -7845 5645 -7811
rect 5705 -7845 5717 -7811
rect 5773 -7845 5789 -7811
rect 5841 -7845 5861 -7811
rect 5909 -7845 5933 -7811
rect 5977 -7845 6005 -7811
rect 6045 -7845 6077 -7811
rect 6113 -7845 6147 -7811
rect 6183 -7845 6215 -7811
rect 6255 -7845 6283 -7811
rect 6327 -7845 6351 -7811
rect 6399 -7845 6419 -7811
rect 6471 -7845 6487 -7811
rect 6543 -7845 6555 -7811
rect 6615 -7845 6623 -7811
rect 6687 -7845 6691 -7811
rect 6793 -7845 6797 -7811
rect 6861 -7845 6869 -7811
rect 6929 -7845 6941 -7811
rect 6997 -7845 7013 -7811
rect 7065 -7845 7085 -7811
rect 7133 -7845 7157 -7811
rect 7201 -7845 7229 -7811
rect 7269 -7845 7301 -7811
rect 7337 -7845 7371 -7811
rect 7407 -7845 7439 -7811
rect 7479 -7845 7507 -7811
rect 7551 -7845 7575 -7811
rect 7623 -7845 7643 -7811
rect 7695 -7845 7711 -7811
rect 7767 -7845 7779 -7811
rect 7839 -7845 7847 -7811
rect 7911 -7845 7915 -7811
rect 8017 -7845 8021 -7811
rect 8085 -7845 8093 -7811
rect 8153 -7845 8165 -7811
rect 8221 -7845 8237 -7811
rect 8289 -7845 8309 -7811
rect 8357 -7845 8381 -7811
rect 8425 -7845 8453 -7811
rect 8493 -7845 8525 -7811
rect 8561 -7845 8595 -7811
rect 8631 -7845 8663 -7811
rect 8703 -7845 8731 -7811
rect 8775 -7845 8799 -7811
rect 8847 -7845 8867 -7811
rect 8919 -7845 8935 -7811
rect 8991 -7845 9003 -7811
rect 9063 -7845 9071 -7811
rect 9135 -7845 9139 -7811
rect 9241 -7845 9245 -7811
rect 9309 -7845 9317 -7811
rect 9377 -7845 9389 -7811
rect 9445 -7845 9461 -7811
rect 9513 -7845 9533 -7811
rect 9581 -7845 9605 -7811
rect 9649 -7845 9677 -7811
rect 9717 -7845 9749 -7811
rect 9785 -7845 9819 -7811
rect 9855 -7845 9887 -7811
rect 9927 -7845 9955 -7811
rect 9999 -7845 10023 -7811
rect 10071 -7845 10091 -7811
rect 10143 -7845 10159 -7811
rect 10215 -7845 10227 -7811
rect 10287 -7845 10295 -7811
rect 10359 -7845 10363 -7811
rect 10465 -7845 10469 -7811
rect 10533 -7845 10541 -7811
rect 10601 -7845 10613 -7811
rect 10669 -7845 10685 -7811
rect 10737 -7845 10757 -7811
rect 10805 -7845 10829 -7811
rect 10873 -7845 10901 -7811
rect 10941 -7845 10973 -7811
rect 11009 -7845 11043 -7811
rect 11079 -7845 11111 -7811
rect 11151 -7845 11179 -7811
rect 11223 -7845 11247 -7811
rect 11295 -7845 11315 -7811
rect 11367 -7845 11383 -7811
rect 11439 -7845 11451 -7811
rect 11511 -7845 11519 -7811
rect 11583 -7845 11587 -7811
rect 11689 -7845 11693 -7811
rect 11757 -7845 11765 -7811
rect 11825 -7845 11837 -7811
rect 11893 -7845 11909 -7811
rect 11961 -7845 11981 -7811
rect 12029 -7845 12053 -7811
rect 12097 -7845 12125 -7811
rect 12165 -7845 12197 -7811
rect 12233 -7845 12267 -7811
rect 12303 -7845 12335 -7811
rect 12375 -7845 12403 -7811
rect 12447 -7845 12485 -7811
rect 12519 -7845 12622 -7811
rect -362 -7878 12622 -7845
rect -362 -7957 -262 -7878
rect -362 -7991 -329 -7957
rect -295 -7991 -262 -7957
rect -362 -7999 -262 -7991
rect -362 -8059 -329 -7999
rect -295 -8059 -262 -7999
rect -362 -8071 -262 -8059
rect -362 -8127 -329 -8071
rect -295 -8127 -262 -8071
rect -362 -8143 -262 -8127
rect -362 -8195 -329 -8143
rect -295 -8195 -262 -8143
rect -362 -8215 -262 -8195
rect -362 -8263 -329 -8215
rect -295 -8263 -262 -8215
rect -362 -8287 -262 -8263
rect -362 -8331 -329 -8287
rect -295 -8331 -262 -8287
rect -362 -8359 -262 -8331
rect -362 -8399 -329 -8359
rect -295 -8399 -262 -8359
rect -362 -8431 -262 -8399
rect -362 -8467 -329 -8431
rect -295 -8467 -262 -8431
rect -362 -8501 -262 -8467
rect -362 -8537 -329 -8501
rect -295 -8537 -262 -8501
rect -362 -8569 -262 -8537
rect -362 -8609 -329 -8569
rect -295 -8609 -262 -8569
rect -362 -8637 -262 -8609
rect -362 -8681 -329 -8637
rect -295 -8681 -262 -8637
rect -362 -8705 -262 -8681
rect -362 -8753 -329 -8705
rect -295 -8753 -262 -8705
rect -362 -8773 -262 -8753
rect -362 -8825 -329 -8773
rect -295 -8825 -262 -8773
rect -362 -8841 -262 -8825
rect -362 -8897 -329 -8841
rect -295 -8897 -262 -8841
rect -362 -8909 -262 -8897
rect -362 -8969 -329 -8909
rect -295 -8969 -262 -8909
rect -362 -8977 -262 -8969
rect -362 -9041 -329 -8977
rect -295 -9041 -262 -8977
rect -362 -9045 -262 -9041
rect -362 -9147 -329 -9045
rect -295 -9147 -262 -9045
rect -362 -9151 -262 -9147
rect -362 -9215 -329 -9151
rect -295 -9215 -262 -9151
rect -362 -9223 -262 -9215
rect -362 -9283 -329 -9223
rect -295 -9283 -262 -9223
rect -362 -9295 -262 -9283
rect -362 -9351 -329 -9295
rect -295 -9351 -262 -9295
rect -362 -9367 -262 -9351
rect -362 -9419 -329 -9367
rect -295 -9419 -262 -9367
rect -362 -9439 -262 -9419
rect -362 -9487 -329 -9439
rect -295 -9487 -262 -9439
rect -362 -9511 -262 -9487
rect -362 -9555 -329 -9511
rect -295 -9555 -262 -9511
rect -362 -9583 -262 -9555
rect -362 -9623 -329 -9583
rect -295 -9623 -262 -9583
rect -362 -9655 -262 -9623
rect -362 -9691 -329 -9655
rect -295 -9691 -262 -9655
rect -362 -9725 -262 -9691
rect -362 -9761 -329 -9725
rect -295 -9761 -262 -9725
rect -362 -9793 -262 -9761
rect -362 -9833 -329 -9793
rect -295 -9833 -262 -9793
rect -362 -9861 -262 -9833
rect -362 -9905 -329 -9861
rect -295 -9905 -262 -9861
rect -362 -9929 -262 -9905
rect -362 -9977 -329 -9929
rect -295 -9977 -262 -9929
rect -362 -9997 -262 -9977
rect -362 -10049 -329 -9997
rect -295 -10049 -262 -9997
rect -362 -10065 -262 -10049
rect -362 -10121 -329 -10065
rect -295 -10121 -262 -10065
rect -362 -10133 -262 -10121
rect -362 -10193 -329 -10133
rect -295 -10193 -262 -10133
rect -362 -10201 -262 -10193
rect -362 -10265 -329 -10201
rect -295 -10265 -262 -10201
rect -362 -10269 -262 -10265
rect -362 -10371 -329 -10269
rect -295 -10371 -262 -10269
rect -362 -10375 -262 -10371
rect -362 -10439 -329 -10375
rect -295 -10439 -262 -10375
rect -362 -10447 -262 -10439
rect -362 -10507 -329 -10447
rect -295 -10507 -262 -10447
rect -362 -10519 -262 -10507
rect -362 -10575 -329 -10519
rect -295 -10575 -262 -10519
rect -362 -10609 -262 -10575
rect -362 -10643 -329 -10609
rect -295 -10643 -262 -10609
rect -362 -10722 -262 -10643
rect 12522 -7957 12622 -7878
rect 12522 -7991 12555 -7957
rect 12589 -7991 12622 -7957
rect 12522 -7999 12622 -7991
rect 12522 -8059 12555 -7999
rect 12589 -8059 12622 -7999
rect 12522 -8071 12622 -8059
rect 12522 -8127 12555 -8071
rect 12589 -8127 12622 -8071
rect 12522 -8143 12622 -8127
rect 12522 -8195 12555 -8143
rect 12589 -8195 12622 -8143
rect 12522 -8215 12622 -8195
rect 12522 -8263 12555 -8215
rect 12589 -8263 12622 -8215
rect 12522 -8287 12622 -8263
rect 12522 -8331 12555 -8287
rect 12589 -8331 12622 -8287
rect 12522 -8359 12622 -8331
rect 12522 -8399 12555 -8359
rect 12589 -8399 12622 -8359
rect 12522 -8431 12622 -8399
rect 12522 -8467 12555 -8431
rect 12589 -8467 12622 -8431
rect 12522 -8501 12622 -8467
rect 12522 -8537 12555 -8501
rect 12589 -8537 12622 -8501
rect 12522 -8569 12622 -8537
rect 12522 -8609 12555 -8569
rect 12589 -8609 12622 -8569
rect 12522 -8637 12622 -8609
rect 12522 -8681 12555 -8637
rect 12589 -8681 12622 -8637
rect 12522 -8705 12622 -8681
rect 12522 -8753 12555 -8705
rect 12589 -8753 12622 -8705
rect 12522 -8773 12622 -8753
rect 12522 -8825 12555 -8773
rect 12589 -8825 12622 -8773
rect 12522 -8841 12622 -8825
rect 12522 -8897 12555 -8841
rect 12589 -8897 12622 -8841
rect 12522 -8909 12622 -8897
rect 12522 -8969 12555 -8909
rect 12589 -8969 12622 -8909
rect 12522 -8977 12622 -8969
rect 12522 -9041 12555 -8977
rect 12589 -9041 12622 -8977
rect 12522 -9045 12622 -9041
rect 12522 -9147 12555 -9045
rect 12589 -9147 12622 -9045
rect 12522 -9151 12622 -9147
rect 12522 -9215 12555 -9151
rect 12589 -9215 12622 -9151
rect 12522 -9223 12622 -9215
rect 12522 -9283 12555 -9223
rect 12589 -9283 12622 -9223
rect 12522 -9295 12622 -9283
rect 12522 -9351 12555 -9295
rect 12589 -9351 12622 -9295
rect 12522 -9367 12622 -9351
rect 12522 -9419 12555 -9367
rect 12589 -9419 12622 -9367
rect 12522 -9439 12622 -9419
rect 12522 -9487 12555 -9439
rect 12589 -9487 12622 -9439
rect 12522 -9511 12622 -9487
rect 12522 -9555 12555 -9511
rect 12589 -9555 12622 -9511
rect 12522 -9583 12622 -9555
rect 12522 -9623 12555 -9583
rect 12589 -9623 12622 -9583
rect 12522 -9655 12622 -9623
rect 12522 -9691 12555 -9655
rect 12589 -9691 12622 -9655
rect 12522 -9725 12622 -9691
rect 12522 -9761 12555 -9725
rect 12589 -9761 12622 -9725
rect 12522 -9793 12622 -9761
rect 12522 -9833 12555 -9793
rect 12589 -9833 12622 -9793
rect 12522 -9861 12622 -9833
rect 12522 -9905 12555 -9861
rect 12589 -9905 12622 -9861
rect 12522 -9929 12622 -9905
rect 12522 -9977 12555 -9929
rect 12589 -9977 12622 -9929
rect 12522 -9997 12622 -9977
rect 12522 -10049 12555 -9997
rect 12589 -10049 12622 -9997
rect 12522 -10065 12622 -10049
rect 12522 -10121 12555 -10065
rect 12589 -10121 12622 -10065
rect 12522 -10133 12622 -10121
rect 12522 -10193 12555 -10133
rect 12589 -10193 12622 -10133
rect 12522 -10201 12622 -10193
rect 12522 -10265 12555 -10201
rect 12589 -10265 12622 -10201
rect 12522 -10269 12622 -10265
rect 12522 -10371 12555 -10269
rect 12589 -10371 12622 -10269
rect 12522 -10375 12622 -10371
rect 12522 -10439 12555 -10375
rect 12589 -10439 12622 -10375
rect 12522 -10447 12622 -10439
rect 12522 -10507 12555 -10447
rect 12589 -10507 12622 -10447
rect 12522 -10519 12622 -10507
rect 12522 -10575 12555 -10519
rect 12589 -10575 12622 -10519
rect 12522 -10609 12622 -10575
rect 12522 -10643 12555 -10609
rect 12589 -10643 12622 -10609
rect 12522 -10722 12622 -10643
rect -362 -10755 12622 -10722
rect -362 -10789 -259 -10755
rect -225 -10789 -187 -10755
rect -143 -10789 -115 -10755
rect -75 -10789 -43 -10755
rect -7 -10789 27 -10755
rect 63 -10789 95 -10755
rect 135 -10789 163 -10755
rect 207 -10789 231 -10755
rect 279 -10789 299 -10755
rect 351 -10789 367 -10755
rect 423 -10789 435 -10755
rect 495 -10789 503 -10755
rect 567 -10789 571 -10755
rect 673 -10789 677 -10755
rect 741 -10789 749 -10755
rect 809 -10789 821 -10755
rect 877 -10789 893 -10755
rect 945 -10789 965 -10755
rect 1013 -10789 1037 -10755
rect 1081 -10789 1109 -10755
rect 1149 -10789 1181 -10755
rect 1217 -10789 1251 -10755
rect 1287 -10789 1319 -10755
rect 1359 -10789 1387 -10755
rect 1431 -10789 1455 -10755
rect 1503 -10789 1523 -10755
rect 1575 -10789 1591 -10755
rect 1647 -10789 1659 -10755
rect 1719 -10789 1727 -10755
rect 1791 -10789 1795 -10755
rect 1897 -10789 1901 -10755
rect 1965 -10789 1973 -10755
rect 2033 -10789 2045 -10755
rect 2101 -10789 2117 -10755
rect 2169 -10789 2189 -10755
rect 2237 -10789 2261 -10755
rect 2305 -10789 2333 -10755
rect 2373 -10789 2405 -10755
rect 2441 -10789 2475 -10755
rect 2511 -10789 2543 -10755
rect 2583 -10789 2611 -10755
rect 2655 -10789 2679 -10755
rect 2727 -10789 2747 -10755
rect 2799 -10789 2815 -10755
rect 2871 -10789 2883 -10755
rect 2943 -10789 2951 -10755
rect 3015 -10789 3019 -10755
rect 3121 -10789 3125 -10755
rect 3189 -10789 3197 -10755
rect 3257 -10789 3269 -10755
rect 3325 -10789 3341 -10755
rect 3393 -10789 3413 -10755
rect 3461 -10789 3485 -10755
rect 3529 -10789 3557 -10755
rect 3597 -10789 3629 -10755
rect 3665 -10789 3699 -10755
rect 3735 -10789 3767 -10755
rect 3807 -10789 3835 -10755
rect 3879 -10789 3903 -10755
rect 3951 -10789 3971 -10755
rect 4023 -10789 4039 -10755
rect 4095 -10789 4107 -10755
rect 4167 -10789 4175 -10755
rect 4239 -10789 4243 -10755
rect 4345 -10789 4349 -10755
rect 4413 -10789 4421 -10755
rect 4481 -10789 4493 -10755
rect 4549 -10789 4565 -10755
rect 4617 -10789 4637 -10755
rect 4685 -10789 4709 -10755
rect 4753 -10789 4781 -10755
rect 4821 -10789 4853 -10755
rect 4889 -10789 4923 -10755
rect 4959 -10789 4991 -10755
rect 5031 -10789 5059 -10755
rect 5103 -10789 5127 -10755
rect 5175 -10789 5195 -10755
rect 5247 -10789 5263 -10755
rect 5319 -10789 5331 -10755
rect 5391 -10789 5399 -10755
rect 5463 -10789 5467 -10755
rect 5569 -10789 5573 -10755
rect 5637 -10789 5645 -10755
rect 5705 -10789 5717 -10755
rect 5773 -10789 5789 -10755
rect 5841 -10789 5861 -10755
rect 5909 -10789 5933 -10755
rect 5977 -10789 6005 -10755
rect 6045 -10789 6077 -10755
rect 6113 -10789 6147 -10755
rect 6183 -10789 6215 -10755
rect 6255 -10789 6283 -10755
rect 6327 -10789 6351 -10755
rect 6399 -10789 6419 -10755
rect 6471 -10789 6487 -10755
rect 6543 -10789 6555 -10755
rect 6615 -10789 6623 -10755
rect 6687 -10789 6691 -10755
rect 6793 -10789 6797 -10755
rect 6861 -10789 6869 -10755
rect 6929 -10789 6941 -10755
rect 6997 -10789 7013 -10755
rect 7065 -10789 7085 -10755
rect 7133 -10789 7157 -10755
rect 7201 -10789 7229 -10755
rect 7269 -10789 7301 -10755
rect 7337 -10789 7371 -10755
rect 7407 -10789 7439 -10755
rect 7479 -10789 7507 -10755
rect 7551 -10789 7575 -10755
rect 7623 -10789 7643 -10755
rect 7695 -10789 7711 -10755
rect 7767 -10789 7779 -10755
rect 7839 -10789 7847 -10755
rect 7911 -10789 7915 -10755
rect 8017 -10789 8021 -10755
rect 8085 -10789 8093 -10755
rect 8153 -10789 8165 -10755
rect 8221 -10789 8237 -10755
rect 8289 -10789 8309 -10755
rect 8357 -10789 8381 -10755
rect 8425 -10789 8453 -10755
rect 8493 -10789 8525 -10755
rect 8561 -10789 8595 -10755
rect 8631 -10789 8663 -10755
rect 8703 -10789 8731 -10755
rect 8775 -10789 8799 -10755
rect 8847 -10789 8867 -10755
rect 8919 -10789 8935 -10755
rect 8991 -10789 9003 -10755
rect 9063 -10789 9071 -10755
rect 9135 -10789 9139 -10755
rect 9241 -10789 9245 -10755
rect 9309 -10789 9317 -10755
rect 9377 -10789 9389 -10755
rect 9445 -10789 9461 -10755
rect 9513 -10789 9533 -10755
rect 9581 -10789 9605 -10755
rect 9649 -10789 9677 -10755
rect 9717 -10789 9749 -10755
rect 9785 -10789 9819 -10755
rect 9855 -10789 9887 -10755
rect 9927 -10789 9955 -10755
rect 9999 -10789 10023 -10755
rect 10071 -10789 10091 -10755
rect 10143 -10789 10159 -10755
rect 10215 -10789 10227 -10755
rect 10287 -10789 10295 -10755
rect 10359 -10789 10363 -10755
rect 10465 -10789 10469 -10755
rect 10533 -10789 10541 -10755
rect 10601 -10789 10613 -10755
rect 10669 -10789 10685 -10755
rect 10737 -10789 10757 -10755
rect 10805 -10789 10829 -10755
rect 10873 -10789 10901 -10755
rect 10941 -10789 10973 -10755
rect 11009 -10789 11043 -10755
rect 11079 -10789 11111 -10755
rect 11151 -10789 11179 -10755
rect 11223 -10789 11247 -10755
rect 11295 -10789 11315 -10755
rect 11367 -10789 11383 -10755
rect 11439 -10789 11451 -10755
rect 11511 -10789 11519 -10755
rect 11583 -10789 11587 -10755
rect 11689 -10789 11693 -10755
rect 11757 -10789 11765 -10755
rect 11825 -10789 11837 -10755
rect 11893 -10789 11909 -10755
rect 11961 -10789 11981 -10755
rect 12029 -10789 12053 -10755
rect 12097 -10789 12125 -10755
rect 12165 -10789 12197 -10755
rect 12233 -10789 12267 -10755
rect 12303 -10789 12335 -10755
rect 12375 -10789 12403 -10755
rect 12447 -10789 12485 -10755
rect 12519 -10789 12622 -10755
rect -362 -10822 12622 -10789
<< viali >>
rect -259 2855 -225 2889
rect -187 2855 -177 2889
rect -177 2855 -153 2889
rect -115 2855 -109 2889
rect -109 2855 -81 2889
rect -43 2855 -41 2889
rect -41 2855 -9 2889
rect 29 2855 61 2889
rect 61 2855 63 2889
rect 101 2855 129 2889
rect 129 2855 135 2889
rect 173 2855 197 2889
rect 197 2855 207 2889
rect 245 2855 265 2889
rect 265 2855 279 2889
rect 317 2855 333 2889
rect 333 2855 351 2889
rect 389 2855 401 2889
rect 401 2855 423 2889
rect 461 2855 469 2889
rect 469 2855 495 2889
rect 533 2855 537 2889
rect 537 2855 567 2889
rect 605 2855 639 2889
rect 677 2855 707 2889
rect 707 2855 711 2889
rect 749 2855 775 2889
rect 775 2855 783 2889
rect 821 2855 843 2889
rect 843 2855 855 2889
rect 893 2855 911 2889
rect 911 2855 927 2889
rect 965 2855 979 2889
rect 979 2855 999 2889
rect 1037 2855 1047 2889
rect 1047 2855 1071 2889
rect 1109 2855 1115 2889
rect 1115 2855 1143 2889
rect 1181 2855 1183 2889
rect 1183 2855 1215 2889
rect 1253 2855 1285 2889
rect 1285 2855 1287 2889
rect 1325 2855 1353 2889
rect 1353 2855 1359 2889
rect 1397 2855 1421 2889
rect 1421 2855 1431 2889
rect 1469 2855 1489 2889
rect 1489 2855 1503 2889
rect 1541 2855 1557 2889
rect 1557 2855 1575 2889
rect 1613 2855 1625 2889
rect 1625 2855 1647 2889
rect 1685 2855 1693 2889
rect 1693 2855 1719 2889
rect 1757 2855 1761 2889
rect 1761 2855 1791 2889
rect 1829 2855 1863 2889
rect 1901 2855 1931 2889
rect 1931 2855 1935 2889
rect 1973 2855 1999 2889
rect 1999 2855 2007 2889
rect 2045 2855 2067 2889
rect 2067 2855 2079 2889
rect 2117 2855 2135 2889
rect 2135 2855 2151 2889
rect 2189 2855 2203 2889
rect 2203 2855 2223 2889
rect 2261 2855 2271 2889
rect 2271 2855 2295 2889
rect 2333 2855 2339 2889
rect 2339 2855 2367 2889
rect 2405 2855 2407 2889
rect 2407 2855 2439 2889
rect 2477 2855 2509 2889
rect 2509 2855 2511 2889
rect 2549 2855 2577 2889
rect 2577 2855 2583 2889
rect 2621 2855 2645 2889
rect 2645 2855 2655 2889
rect 2693 2855 2713 2889
rect 2713 2855 2727 2889
rect 2765 2855 2781 2889
rect 2781 2855 2799 2889
rect 2837 2855 2849 2889
rect 2849 2855 2871 2889
rect 2909 2855 2917 2889
rect 2917 2855 2943 2889
rect 2981 2855 2985 2889
rect 2985 2855 3015 2889
rect 3053 2855 3087 2889
rect 3125 2855 3155 2889
rect 3155 2855 3159 2889
rect 3197 2855 3223 2889
rect 3223 2855 3231 2889
rect 3269 2855 3291 2889
rect 3291 2855 3303 2889
rect 3341 2855 3359 2889
rect 3359 2855 3375 2889
rect 3413 2855 3427 2889
rect 3427 2855 3447 2889
rect 3485 2855 3495 2889
rect 3495 2855 3519 2889
rect 3557 2855 3563 2889
rect 3563 2855 3591 2889
rect 3629 2855 3631 2889
rect 3631 2855 3663 2889
rect 3701 2855 3733 2889
rect 3733 2855 3735 2889
rect 3773 2855 3801 2889
rect 3801 2855 3807 2889
rect 3845 2855 3869 2889
rect 3869 2855 3879 2889
rect 3917 2855 3937 2889
rect 3937 2855 3951 2889
rect 3989 2855 4005 2889
rect 4005 2855 4023 2889
rect 4061 2855 4073 2889
rect 4073 2855 4095 2889
rect 4133 2855 4141 2889
rect 4141 2855 4167 2889
rect 4205 2855 4209 2889
rect 4209 2855 4239 2889
rect 4277 2855 4311 2889
rect 4349 2855 4379 2889
rect 4379 2855 4383 2889
rect 4421 2855 4447 2889
rect 4447 2855 4455 2889
rect 4493 2855 4515 2889
rect 4515 2855 4527 2889
rect 4565 2855 4583 2889
rect 4583 2855 4599 2889
rect 4637 2855 4651 2889
rect 4651 2855 4671 2889
rect 4709 2855 4719 2889
rect 4719 2855 4743 2889
rect 4781 2855 4787 2889
rect 4787 2855 4815 2889
rect 4853 2855 4855 2889
rect 4855 2855 4887 2889
rect 4925 2855 4957 2889
rect 4957 2855 4959 2889
rect 4997 2855 5025 2889
rect 5025 2855 5031 2889
rect 5069 2855 5093 2889
rect 5093 2855 5103 2889
rect 5141 2855 5161 2889
rect 5161 2855 5175 2889
rect 5213 2855 5229 2889
rect 5229 2855 5247 2889
rect 5285 2855 5297 2889
rect 5297 2855 5319 2889
rect 5357 2855 5365 2889
rect 5365 2855 5391 2889
rect 5429 2855 5433 2889
rect 5433 2855 5463 2889
rect 5501 2855 5535 2889
rect 5573 2855 5603 2889
rect 5603 2855 5607 2889
rect 5645 2855 5671 2889
rect 5671 2855 5679 2889
rect 5717 2855 5739 2889
rect 5739 2855 5751 2889
rect 5789 2855 5807 2889
rect 5807 2855 5823 2889
rect 5861 2855 5875 2889
rect 5875 2855 5895 2889
rect 5933 2855 5943 2889
rect 5943 2855 5967 2889
rect 6005 2855 6011 2889
rect 6011 2855 6039 2889
rect 6077 2855 6079 2889
rect 6079 2855 6111 2889
rect 6149 2855 6181 2889
rect 6181 2855 6183 2889
rect 6221 2855 6249 2889
rect 6249 2855 6255 2889
rect 6293 2855 6317 2889
rect 6317 2855 6327 2889
rect 6365 2855 6385 2889
rect 6385 2855 6399 2889
rect 6437 2855 6453 2889
rect 6453 2855 6471 2889
rect 6509 2855 6521 2889
rect 6521 2855 6543 2889
rect 6581 2855 6589 2889
rect 6589 2855 6615 2889
rect 6653 2855 6657 2889
rect 6657 2855 6687 2889
rect 6725 2855 6759 2889
rect 6797 2855 6827 2889
rect 6827 2855 6831 2889
rect 6869 2855 6895 2889
rect 6895 2855 6903 2889
rect 6941 2855 6963 2889
rect 6963 2855 6975 2889
rect 7013 2855 7031 2889
rect 7031 2855 7047 2889
rect 7085 2855 7099 2889
rect 7099 2855 7119 2889
rect 7157 2855 7167 2889
rect 7167 2855 7191 2889
rect 7229 2855 7235 2889
rect 7235 2855 7263 2889
rect 7301 2855 7303 2889
rect 7303 2855 7335 2889
rect 7373 2855 7405 2889
rect 7405 2855 7407 2889
rect 7445 2855 7473 2889
rect 7473 2855 7479 2889
rect 7517 2855 7541 2889
rect 7541 2855 7551 2889
rect 7589 2855 7609 2889
rect 7609 2855 7623 2889
rect 7661 2855 7677 2889
rect 7677 2855 7695 2889
rect 7733 2855 7745 2889
rect 7745 2855 7767 2889
rect 7805 2855 7813 2889
rect 7813 2855 7839 2889
rect 7877 2855 7881 2889
rect 7881 2855 7911 2889
rect 7949 2855 7983 2889
rect 8021 2855 8051 2889
rect 8051 2855 8055 2889
rect 8093 2855 8119 2889
rect 8119 2855 8127 2889
rect 8165 2855 8187 2889
rect 8187 2855 8199 2889
rect 8237 2855 8255 2889
rect 8255 2855 8271 2889
rect 8309 2855 8323 2889
rect 8323 2855 8343 2889
rect 8381 2855 8391 2889
rect 8391 2855 8415 2889
rect 8453 2855 8459 2889
rect 8459 2855 8487 2889
rect 8525 2855 8527 2889
rect 8527 2855 8559 2889
rect 8597 2855 8629 2889
rect 8629 2855 8631 2889
rect 8669 2855 8697 2889
rect 8697 2855 8703 2889
rect 8741 2855 8765 2889
rect 8765 2855 8775 2889
rect 8813 2855 8833 2889
rect 8833 2855 8847 2889
rect 8885 2855 8901 2889
rect 8901 2855 8919 2889
rect 8957 2855 8969 2889
rect 8969 2855 8991 2889
rect 9029 2855 9037 2889
rect 9037 2855 9063 2889
rect 9101 2855 9105 2889
rect 9105 2855 9135 2889
rect 9173 2855 9207 2889
rect 9245 2855 9275 2889
rect 9275 2855 9279 2889
rect 9317 2855 9343 2889
rect 9343 2855 9351 2889
rect 9389 2855 9411 2889
rect 9411 2855 9423 2889
rect 9461 2855 9479 2889
rect 9479 2855 9495 2889
rect 9533 2855 9547 2889
rect 9547 2855 9567 2889
rect 9605 2855 9615 2889
rect 9615 2855 9639 2889
rect 9677 2855 9683 2889
rect 9683 2855 9711 2889
rect 9749 2855 9751 2889
rect 9751 2855 9783 2889
rect 9821 2855 9853 2889
rect 9853 2855 9855 2889
rect 9893 2855 9921 2889
rect 9921 2855 9927 2889
rect 9965 2855 9989 2889
rect 9989 2855 9999 2889
rect 10037 2855 10057 2889
rect 10057 2855 10071 2889
rect 10109 2855 10125 2889
rect 10125 2855 10143 2889
rect 10181 2855 10193 2889
rect 10193 2855 10215 2889
rect 10253 2855 10261 2889
rect 10261 2855 10287 2889
rect 10325 2855 10329 2889
rect 10329 2855 10359 2889
rect 10397 2855 10431 2889
rect 10469 2855 10499 2889
rect 10499 2855 10503 2889
rect 10541 2855 10567 2889
rect 10567 2855 10575 2889
rect 10613 2855 10635 2889
rect 10635 2855 10647 2889
rect 10685 2855 10703 2889
rect 10703 2855 10719 2889
rect 10757 2855 10771 2889
rect 10771 2855 10791 2889
rect 10829 2855 10839 2889
rect 10839 2855 10863 2889
rect 10901 2855 10907 2889
rect 10907 2855 10935 2889
rect 10973 2855 10975 2889
rect 10975 2855 11007 2889
rect 11045 2855 11077 2889
rect 11077 2855 11079 2889
rect 11117 2855 11145 2889
rect 11145 2855 11151 2889
rect 11189 2855 11213 2889
rect 11213 2855 11223 2889
rect 11261 2855 11281 2889
rect 11281 2855 11295 2889
rect 11333 2855 11349 2889
rect 11349 2855 11367 2889
rect 11405 2855 11417 2889
rect 11417 2855 11439 2889
rect 11477 2855 11485 2889
rect 11485 2855 11511 2889
rect 11549 2855 11553 2889
rect 11553 2855 11583 2889
rect 11621 2855 11655 2889
rect 11693 2855 11723 2889
rect 11723 2855 11727 2889
rect 11765 2855 11791 2889
rect 11791 2855 11799 2889
rect 11837 2855 11859 2889
rect 11859 2855 11871 2889
rect 11909 2855 11927 2889
rect 11927 2855 11943 2889
rect 11981 2855 11995 2889
rect 11995 2855 12015 2889
rect 12053 2855 12063 2889
rect 12063 2855 12087 2889
rect 12125 2855 12131 2889
rect 12131 2855 12159 2889
rect 12197 2855 12199 2889
rect 12199 2855 12231 2889
rect 12269 2855 12301 2889
rect 12301 2855 12303 2889
rect 12341 2855 12369 2889
rect 12369 2855 12375 2889
rect 12413 2855 12437 2889
rect 12437 2855 12447 2889
rect 12485 2855 12519 2889
rect -329 2263 -295 2287
rect -329 2253 -295 2263
rect -329 2195 -295 2215
rect -329 2181 -295 2195
rect -329 2127 -295 2143
rect -329 2109 -295 2127
rect -329 2059 -295 2071
rect -329 2037 -295 2059
rect -329 1991 -295 1999
rect -329 1965 -295 1991
rect -329 1923 -295 1927
rect -329 1893 -295 1923
rect -329 1821 -295 1855
rect -329 1753 -295 1783
rect -329 1749 -295 1753
rect -329 1685 -295 1711
rect -329 1677 -295 1685
rect -329 1617 -295 1639
rect -329 1605 -295 1617
rect -329 1549 -295 1567
rect -329 1533 -295 1549
rect -329 1481 -295 1495
rect -329 1461 -295 1481
rect -329 1413 -295 1423
rect -329 1389 -295 1413
rect -329 1345 -295 1351
rect -329 1317 -295 1345
rect -329 1277 -295 1279
rect -329 1245 -295 1277
rect -329 1175 -295 1207
rect -329 1173 -295 1175
rect -329 1107 -295 1135
rect -329 1101 -295 1107
rect -329 1039 -295 1063
rect -329 1029 -295 1039
rect -329 971 -295 991
rect -329 957 -295 971
rect -329 903 -295 919
rect -329 885 -295 903
rect -329 835 -295 847
rect -329 813 -295 835
rect -329 767 -295 775
rect -329 741 -295 767
rect -329 699 -295 703
rect -329 669 -295 699
rect -329 597 -295 631
rect -329 529 -295 559
rect -329 525 -295 529
rect -329 461 -295 487
rect -329 453 -295 461
rect -329 393 -295 415
rect -329 381 -295 393
rect -329 325 -295 343
rect -329 309 -295 325
rect -329 257 -295 271
rect -329 237 -295 257
rect -329 189 -295 199
rect -329 165 -295 189
rect -329 121 -295 127
rect -329 93 -295 121
rect -329 53 -295 55
rect -329 21 -295 53
rect -329 -49 -295 -17
rect -329 -51 -295 -49
rect -329 -117 -295 -89
rect -329 -123 -295 -117
rect -329 -185 -295 -161
rect -329 -195 -295 -185
rect -329 -253 -295 -233
rect -329 -267 -295 -253
rect -329 -321 -295 -305
rect -329 -339 -295 -321
rect -329 -389 -295 -377
rect -329 -411 -295 -389
rect -329 -457 -295 -449
rect -329 -483 -295 -457
rect -329 -525 -295 -521
rect -329 -555 -295 -525
rect -329 -627 -295 -593
rect -329 -695 -295 -665
rect -329 -699 -295 -695
rect -329 -763 -295 -737
rect -329 -771 -295 -763
rect -329 -831 -295 -809
rect -329 -843 -295 -831
rect -329 -899 -295 -881
rect -329 -915 -295 -899
rect -329 -967 -295 -953
rect -329 -987 -295 -967
rect -329 -1035 -295 -1025
rect -329 -1059 -295 -1035
rect -329 -1103 -295 -1097
rect -329 -1131 -295 -1103
rect -329 -1171 -295 -1169
rect -329 -1203 -295 -1171
rect -329 -1273 -295 -1241
rect -329 -1275 -295 -1273
rect -329 -1341 -295 -1313
rect -329 -1347 -295 -1341
rect -329 -1409 -295 -1385
rect -329 -1419 -295 -1409
rect -329 -1477 -295 -1457
rect -329 -1491 -295 -1477
rect -329 -1545 -295 -1529
rect -329 -1563 -295 -1545
rect -329 -1613 -295 -1601
rect -329 -1635 -295 -1613
rect -329 -1681 -295 -1673
rect -329 -1707 -295 -1681
rect -329 -1749 -295 -1745
rect -329 -1779 -295 -1749
rect -329 -1851 -295 -1817
rect -329 -1919 -295 -1889
rect -329 -1923 -295 -1919
rect -329 -1987 -295 -1961
rect -329 -1995 -295 -1987
rect -329 -2055 -295 -2033
rect -329 -2067 -295 -2055
rect -329 -2123 -295 -2105
rect -329 -2139 -295 -2123
rect -329 -2191 -295 -2177
rect -329 -2211 -295 -2191
rect -329 -2259 -295 -2249
rect -329 -2283 -295 -2259
rect -329 -2327 -295 -2321
rect -329 -2355 -295 -2327
rect -329 -2395 -295 -2393
rect -329 -2427 -295 -2395
rect -329 -2497 -295 -2465
rect -329 -2499 -295 -2497
rect -329 -2565 -295 -2537
rect -329 -2571 -295 -2565
rect -329 -2633 -295 -2609
rect -329 -2643 -295 -2633
rect -329 -2701 -295 -2681
rect -329 -2715 -295 -2701
rect -329 -2769 -295 -2753
rect -329 -2787 -295 -2769
rect -329 -2837 -295 -2825
rect -329 -2859 -295 -2837
rect -329 -2905 -295 -2897
rect -329 -2931 -295 -2905
rect -329 -2973 -295 -2969
rect -329 -3003 -295 -2973
rect -329 -3075 -295 -3041
rect -329 -3143 -295 -3113
rect -329 -3147 -295 -3143
rect -329 -3211 -295 -3185
rect -329 -3219 -295 -3211
rect -329 -3279 -295 -3257
rect -329 -3291 -295 -3279
rect -329 -3347 -295 -3329
rect -329 -3363 -295 -3347
rect -329 -3415 -295 -3401
rect -329 -3435 -295 -3415
rect -329 -3483 -295 -3473
rect -329 -3507 -295 -3483
rect -329 -3551 -295 -3545
rect -329 -3579 -295 -3551
rect -329 -3619 -295 -3617
rect -329 -3651 -295 -3619
rect -329 -3721 -295 -3689
rect -329 -3723 -295 -3721
rect -329 -3789 -295 -3761
rect -329 -3795 -295 -3789
rect -329 -3857 -295 -3833
rect -329 -3867 -295 -3857
rect -329 -3925 -295 -3905
rect -329 -3939 -295 -3925
rect -329 -3993 -295 -3977
rect -329 -4011 -295 -3993
rect -329 -4061 -295 -4049
rect -329 -4083 -295 -4061
rect -329 -4129 -295 -4121
rect -329 -4155 -295 -4129
rect -329 -4197 -295 -4193
rect -329 -4227 -295 -4197
rect -329 -4299 -295 -4265
rect -329 -4367 -295 -4337
rect -329 -4371 -295 -4367
rect -329 -4435 -295 -4409
rect -329 -4443 -295 -4435
rect -329 -4503 -295 -4481
rect -329 -4515 -295 -4503
rect -329 -4571 -295 -4553
rect -329 -4587 -295 -4571
rect -329 -4639 -295 -4625
rect -329 -4659 -295 -4639
rect -329 -4707 -295 -4697
rect -329 -4731 -295 -4707
rect -329 -4775 -295 -4769
rect -329 -4803 -295 -4775
rect -329 -4843 -295 -4841
rect -329 -4875 -295 -4843
rect -329 -4945 -295 -4913
rect -329 -4947 -295 -4945
rect -329 -5013 -295 -4985
rect -329 -5019 -295 -5013
rect -329 -5081 -295 -5057
rect -329 -5091 -295 -5081
rect -329 -5149 -295 -5129
rect -329 -5163 -295 -5149
rect -329 -5217 -295 -5201
rect -329 -5235 -295 -5217
rect -329 -5285 -295 -5273
rect -329 -5307 -295 -5285
rect -329 -5353 -295 -5345
rect -329 -5379 -295 -5353
rect -329 -5421 -295 -5417
rect -329 -5451 -295 -5421
rect -329 -5523 -295 -5489
rect -329 -5591 -295 -5561
rect -329 -5595 -295 -5591
rect -329 -5659 -295 -5633
rect -329 -5667 -295 -5659
rect -329 -5727 -295 -5705
rect -329 -5739 -295 -5727
rect -329 -5795 -295 -5777
rect -329 -5811 -295 -5795
rect -329 -5863 -295 -5849
rect -329 -5883 -295 -5863
rect -329 -5931 -295 -5921
rect -329 -5955 -295 -5931
rect -329 -5999 -295 -5993
rect -329 -6027 -295 -5999
rect -329 -6067 -295 -6065
rect -329 -6099 -295 -6067
rect -329 -6169 -295 -6137
rect -329 -6171 -295 -6169
rect -329 -6237 -295 -6209
rect -329 -6243 -295 -6237
rect -329 -6305 -295 -6281
rect -329 -6315 -295 -6305
rect -329 -6373 -295 -6353
rect -329 -6387 -295 -6373
rect -329 -6441 -295 -6425
rect -329 -6459 -295 -6441
rect -329 -6509 -295 -6497
rect -329 -6531 -295 -6509
rect -329 -6577 -295 -6569
rect -329 -6603 -295 -6577
rect -329 -6645 -295 -6641
rect -329 -6675 -295 -6645
rect -329 -6747 -295 -6713
rect -329 -6815 -295 -6785
rect -329 -6819 -295 -6815
rect -329 -6883 -295 -6857
rect -329 -6891 -295 -6883
rect -329 -6951 -295 -6929
rect -329 -6963 -295 -6951
rect -329 -7019 -295 -7001
rect -329 -7035 -295 -7019
rect -329 -7087 -295 -7073
rect -329 -7107 -295 -7087
rect 12555 2263 12589 2287
rect 12555 2253 12589 2263
rect 12555 2195 12589 2215
rect 12555 2181 12589 2195
rect 12555 2127 12589 2143
rect 12555 2109 12589 2127
rect 12555 2059 12589 2071
rect 12555 2037 12589 2059
rect 12555 1991 12589 1999
rect 12555 1965 12589 1991
rect 12555 1923 12589 1927
rect 12555 1893 12589 1923
rect 12555 1821 12589 1855
rect 12555 1753 12589 1783
rect 12555 1749 12589 1753
rect 12555 1685 12589 1711
rect 12555 1677 12589 1685
rect 12555 1617 12589 1639
rect 12555 1605 12589 1617
rect 12555 1549 12589 1567
rect 12555 1533 12589 1549
rect 12555 1481 12589 1495
rect 12555 1461 12589 1481
rect 12555 1413 12589 1423
rect 12555 1389 12589 1413
rect 12555 1345 12589 1351
rect 12555 1317 12589 1345
rect 12555 1277 12589 1279
rect 12555 1245 12589 1277
rect 12555 1175 12589 1207
rect 12555 1173 12589 1175
rect 12555 1107 12589 1135
rect 12555 1101 12589 1107
rect 12555 1039 12589 1063
rect 12555 1029 12589 1039
rect 12555 971 12589 991
rect 12555 957 12589 971
rect 12555 903 12589 919
rect 12555 885 12589 903
rect 12555 835 12589 847
rect 12555 813 12589 835
rect 12555 767 12589 775
rect 12555 741 12589 767
rect 12555 699 12589 703
rect 12555 669 12589 699
rect 12555 597 12589 631
rect 12555 529 12589 559
rect 12555 525 12589 529
rect 12555 461 12589 487
rect 12555 453 12589 461
rect 12555 393 12589 415
rect 12555 381 12589 393
rect 12555 325 12589 343
rect 12555 309 12589 325
rect 12555 257 12589 271
rect 12555 237 12589 257
rect 12555 189 12589 199
rect 12555 165 12589 189
rect 12555 121 12589 127
rect 12555 93 12589 121
rect 12555 53 12589 55
rect 12555 21 12589 53
rect 12555 -49 12589 -17
rect 12555 -51 12589 -49
rect 12555 -117 12589 -89
rect 12555 -123 12589 -117
rect 12555 -185 12589 -161
rect 12555 -195 12589 -185
rect 12555 -253 12589 -233
rect 12555 -267 12589 -253
rect 12555 -321 12589 -305
rect 12555 -339 12589 -321
rect 12555 -389 12589 -377
rect 12555 -411 12589 -389
rect 12555 -457 12589 -449
rect 12555 -483 12589 -457
rect 12555 -525 12589 -521
rect 12555 -555 12589 -525
rect 12555 -627 12589 -593
rect 12555 -695 12589 -665
rect 12555 -699 12589 -695
rect 12555 -763 12589 -737
rect 12555 -771 12589 -763
rect 12555 -831 12589 -809
rect 12555 -843 12589 -831
rect 12555 -899 12589 -881
rect 12555 -915 12589 -899
rect 12555 -967 12589 -953
rect 12555 -987 12589 -967
rect 12555 -1035 12589 -1025
rect 12555 -1059 12589 -1035
rect 12555 -1103 12589 -1097
rect 12555 -1131 12589 -1103
rect 12555 -1171 12589 -1169
rect 12555 -1203 12589 -1171
rect 12555 -1273 12589 -1241
rect 12555 -1275 12589 -1273
rect 12555 -1341 12589 -1313
rect 12555 -1347 12589 -1341
rect 12555 -1409 12589 -1385
rect 12555 -1419 12589 -1409
rect 12555 -1477 12589 -1457
rect 12555 -1491 12589 -1477
rect 12555 -1545 12589 -1529
rect 12555 -1563 12589 -1545
rect 12555 -1613 12589 -1601
rect 12555 -1635 12589 -1613
rect 12555 -1681 12589 -1673
rect 12555 -1707 12589 -1681
rect 12555 -1749 12589 -1745
rect 12555 -1779 12589 -1749
rect 12555 -1851 12589 -1817
rect 12555 -1919 12589 -1889
rect 12555 -1923 12589 -1919
rect 12555 -1987 12589 -1961
rect 12555 -1995 12589 -1987
rect 12555 -2055 12589 -2033
rect 12555 -2067 12589 -2055
rect 12555 -2123 12589 -2105
rect 12555 -2139 12589 -2123
rect 12555 -2191 12589 -2177
rect 12555 -2211 12589 -2191
rect 12555 -2259 12589 -2249
rect 12555 -2283 12589 -2259
rect 12555 -2327 12589 -2321
rect 12555 -2355 12589 -2327
rect 12555 -2395 12589 -2393
rect 12555 -2427 12589 -2395
rect 12555 -2497 12589 -2465
rect 12555 -2499 12589 -2497
rect 12555 -2565 12589 -2537
rect 12555 -2571 12589 -2565
rect 12555 -2633 12589 -2609
rect 12555 -2643 12589 -2633
rect 12555 -2701 12589 -2681
rect 12555 -2715 12589 -2701
rect 12555 -2769 12589 -2753
rect 12555 -2787 12589 -2769
rect 12555 -2837 12589 -2825
rect 12555 -2859 12589 -2837
rect 12555 -2905 12589 -2897
rect 12555 -2931 12589 -2905
rect 12555 -2973 12589 -2969
rect 12555 -3003 12589 -2973
rect 12555 -3075 12589 -3041
rect 12555 -3143 12589 -3113
rect 12555 -3147 12589 -3143
rect 12555 -3211 12589 -3185
rect 12555 -3219 12589 -3211
rect 12555 -3279 12589 -3257
rect 12555 -3291 12589 -3279
rect 12555 -3347 12589 -3329
rect 12555 -3363 12589 -3347
rect 12555 -3415 12589 -3401
rect 12555 -3435 12589 -3415
rect 12555 -3483 12589 -3473
rect 12555 -3507 12589 -3483
rect 12555 -3551 12589 -3545
rect 12555 -3579 12589 -3551
rect 12555 -3619 12589 -3617
rect 12555 -3651 12589 -3619
rect 12555 -3721 12589 -3689
rect 12555 -3723 12589 -3721
rect 12555 -3789 12589 -3761
rect 12555 -3795 12589 -3789
rect 12555 -3857 12589 -3833
rect 12555 -3867 12589 -3857
rect 12555 -3925 12589 -3905
rect 12555 -3939 12589 -3925
rect 12555 -3993 12589 -3977
rect 12555 -4011 12589 -3993
rect 12555 -4061 12589 -4049
rect 12555 -4083 12589 -4061
rect 12555 -4129 12589 -4121
rect 12555 -4155 12589 -4129
rect 12555 -4197 12589 -4193
rect 12555 -4227 12589 -4197
rect 12555 -4299 12589 -4265
rect 12555 -4367 12589 -4337
rect 12555 -4371 12589 -4367
rect 12555 -4435 12589 -4409
rect 12555 -4443 12589 -4435
rect 12555 -4503 12589 -4481
rect 12555 -4515 12589 -4503
rect 12555 -4571 12589 -4553
rect 12555 -4587 12589 -4571
rect 12555 -4639 12589 -4625
rect 12555 -4659 12589 -4639
rect 12555 -4707 12589 -4697
rect 12555 -4731 12589 -4707
rect 12555 -4775 12589 -4769
rect 12555 -4803 12589 -4775
rect 12555 -4843 12589 -4841
rect 12555 -4875 12589 -4843
rect 12555 -4945 12589 -4913
rect 12555 -4947 12589 -4945
rect 12555 -5013 12589 -4985
rect 12555 -5019 12589 -5013
rect 12555 -5081 12589 -5057
rect 12555 -5091 12589 -5081
rect 12555 -5149 12589 -5129
rect 12555 -5163 12589 -5149
rect 12555 -5217 12589 -5201
rect 12555 -5235 12589 -5217
rect 12555 -5285 12589 -5273
rect 12555 -5307 12589 -5285
rect 12555 -5353 12589 -5345
rect 12555 -5379 12589 -5353
rect 12555 -5421 12589 -5417
rect 12555 -5451 12589 -5421
rect 12555 -5523 12589 -5489
rect 12555 -5591 12589 -5561
rect 12555 -5595 12589 -5591
rect 12555 -5659 12589 -5633
rect 12555 -5667 12589 -5659
rect 12555 -5727 12589 -5705
rect 12555 -5739 12589 -5727
rect 12555 -5795 12589 -5777
rect 12555 -5811 12589 -5795
rect 12555 -5863 12589 -5849
rect 12555 -5883 12589 -5863
rect 12555 -5931 12589 -5921
rect 12555 -5955 12589 -5931
rect 12555 -5999 12589 -5993
rect 12555 -6027 12589 -5999
rect 12555 -6067 12589 -6065
rect 12555 -6099 12589 -6067
rect 12555 -6169 12589 -6137
rect 12555 -6171 12589 -6169
rect 12555 -6237 12589 -6209
rect 12555 -6243 12589 -6237
rect 12555 -6305 12589 -6281
rect 12555 -6315 12589 -6305
rect 12555 -6373 12589 -6353
rect 12555 -6387 12589 -6373
rect 12555 -6441 12589 -6425
rect 12555 -6459 12589 -6441
rect 12555 -6509 12589 -6497
rect 12555 -6531 12589 -6509
rect 12555 -6577 12589 -6569
rect 12555 -6603 12589 -6577
rect 12555 -6645 12589 -6641
rect 12555 -6675 12589 -6645
rect 12555 -6747 12589 -6713
rect 12555 -6815 12589 -6785
rect 12555 -6819 12589 -6815
rect 12555 -6883 12589 -6857
rect 12555 -6891 12589 -6883
rect 12555 -6951 12589 -6929
rect 12555 -6963 12589 -6951
rect 12555 -7019 12589 -7001
rect 12555 -7035 12589 -7019
rect 12555 -7087 12589 -7073
rect 12555 -7107 12589 -7087
rect -259 -7509 -225 -7475
rect -187 -7509 -177 -7475
rect -177 -7509 -153 -7475
rect -115 -7509 -109 -7475
rect -109 -7509 -81 -7475
rect -43 -7509 -41 -7475
rect -41 -7509 -9 -7475
rect 29 -7509 61 -7475
rect 61 -7509 63 -7475
rect 101 -7509 129 -7475
rect 129 -7509 135 -7475
rect 173 -7509 197 -7475
rect 197 -7509 207 -7475
rect 245 -7509 265 -7475
rect 265 -7509 279 -7475
rect 317 -7509 333 -7475
rect 333 -7509 351 -7475
rect 389 -7509 401 -7475
rect 401 -7509 423 -7475
rect 461 -7509 469 -7475
rect 469 -7509 495 -7475
rect 533 -7509 537 -7475
rect 537 -7509 567 -7475
rect 605 -7509 639 -7475
rect 677 -7509 707 -7475
rect 707 -7509 711 -7475
rect 749 -7509 775 -7475
rect 775 -7509 783 -7475
rect 821 -7509 843 -7475
rect 843 -7509 855 -7475
rect 893 -7509 911 -7475
rect 911 -7509 927 -7475
rect 965 -7509 979 -7475
rect 979 -7509 999 -7475
rect 1037 -7509 1047 -7475
rect 1047 -7509 1071 -7475
rect 1109 -7509 1115 -7475
rect 1115 -7509 1143 -7475
rect 1181 -7509 1183 -7475
rect 1183 -7509 1215 -7475
rect 1253 -7509 1285 -7475
rect 1285 -7509 1287 -7475
rect 1325 -7509 1353 -7475
rect 1353 -7509 1359 -7475
rect 1397 -7509 1421 -7475
rect 1421 -7509 1431 -7475
rect 1469 -7509 1489 -7475
rect 1489 -7509 1503 -7475
rect 1541 -7509 1557 -7475
rect 1557 -7509 1575 -7475
rect 1613 -7509 1625 -7475
rect 1625 -7509 1647 -7475
rect 1685 -7509 1693 -7475
rect 1693 -7509 1719 -7475
rect 1757 -7509 1761 -7475
rect 1761 -7509 1791 -7475
rect 1829 -7509 1863 -7475
rect 1901 -7509 1931 -7475
rect 1931 -7509 1935 -7475
rect 1973 -7509 1999 -7475
rect 1999 -7509 2007 -7475
rect 2045 -7509 2067 -7475
rect 2067 -7509 2079 -7475
rect 2117 -7509 2135 -7475
rect 2135 -7509 2151 -7475
rect 2189 -7509 2203 -7475
rect 2203 -7509 2223 -7475
rect 2261 -7509 2271 -7475
rect 2271 -7509 2295 -7475
rect 2333 -7509 2339 -7475
rect 2339 -7509 2367 -7475
rect 2405 -7509 2407 -7475
rect 2407 -7509 2439 -7475
rect 2477 -7509 2509 -7475
rect 2509 -7509 2511 -7475
rect 2549 -7509 2577 -7475
rect 2577 -7509 2583 -7475
rect 2621 -7509 2645 -7475
rect 2645 -7509 2655 -7475
rect 2693 -7509 2713 -7475
rect 2713 -7509 2727 -7475
rect 2765 -7509 2781 -7475
rect 2781 -7509 2799 -7475
rect 2837 -7509 2849 -7475
rect 2849 -7509 2871 -7475
rect 2909 -7509 2917 -7475
rect 2917 -7509 2943 -7475
rect 2981 -7509 2985 -7475
rect 2985 -7509 3015 -7475
rect 3053 -7509 3087 -7475
rect 3125 -7509 3155 -7475
rect 3155 -7509 3159 -7475
rect 3197 -7509 3223 -7475
rect 3223 -7509 3231 -7475
rect 3269 -7509 3291 -7475
rect 3291 -7509 3303 -7475
rect 3341 -7509 3359 -7475
rect 3359 -7509 3375 -7475
rect 3413 -7509 3427 -7475
rect 3427 -7509 3447 -7475
rect 3485 -7509 3495 -7475
rect 3495 -7509 3519 -7475
rect 3557 -7509 3563 -7475
rect 3563 -7509 3591 -7475
rect 3629 -7509 3631 -7475
rect 3631 -7509 3663 -7475
rect 3701 -7509 3733 -7475
rect 3733 -7509 3735 -7475
rect 3773 -7509 3801 -7475
rect 3801 -7509 3807 -7475
rect 3845 -7509 3869 -7475
rect 3869 -7509 3879 -7475
rect 3917 -7509 3937 -7475
rect 3937 -7509 3951 -7475
rect 3989 -7509 4005 -7475
rect 4005 -7509 4023 -7475
rect 4061 -7509 4073 -7475
rect 4073 -7509 4095 -7475
rect 4133 -7509 4141 -7475
rect 4141 -7509 4167 -7475
rect 4205 -7509 4209 -7475
rect 4209 -7509 4239 -7475
rect 4277 -7509 4311 -7475
rect 4349 -7509 4379 -7475
rect 4379 -7509 4383 -7475
rect 4421 -7509 4447 -7475
rect 4447 -7509 4455 -7475
rect 4493 -7509 4515 -7475
rect 4515 -7509 4527 -7475
rect 4565 -7509 4583 -7475
rect 4583 -7509 4599 -7475
rect 4637 -7509 4651 -7475
rect 4651 -7509 4671 -7475
rect 4709 -7509 4719 -7475
rect 4719 -7509 4743 -7475
rect 4781 -7509 4787 -7475
rect 4787 -7509 4815 -7475
rect 4853 -7509 4855 -7475
rect 4855 -7509 4887 -7475
rect 4925 -7509 4957 -7475
rect 4957 -7509 4959 -7475
rect 4997 -7509 5025 -7475
rect 5025 -7509 5031 -7475
rect 5069 -7509 5093 -7475
rect 5093 -7509 5103 -7475
rect 5141 -7509 5161 -7475
rect 5161 -7509 5175 -7475
rect 5213 -7509 5229 -7475
rect 5229 -7509 5247 -7475
rect 5285 -7509 5297 -7475
rect 5297 -7509 5319 -7475
rect 5357 -7509 5365 -7475
rect 5365 -7509 5391 -7475
rect 5429 -7509 5433 -7475
rect 5433 -7509 5463 -7475
rect 5501 -7509 5535 -7475
rect 5573 -7509 5603 -7475
rect 5603 -7509 5607 -7475
rect 5645 -7509 5671 -7475
rect 5671 -7509 5679 -7475
rect 5717 -7509 5739 -7475
rect 5739 -7509 5751 -7475
rect 5789 -7509 5807 -7475
rect 5807 -7509 5823 -7475
rect 5861 -7509 5875 -7475
rect 5875 -7509 5895 -7475
rect 5933 -7509 5943 -7475
rect 5943 -7509 5967 -7475
rect 6005 -7509 6011 -7475
rect 6011 -7509 6039 -7475
rect 6077 -7509 6079 -7475
rect 6079 -7509 6111 -7475
rect 6149 -7509 6181 -7475
rect 6181 -7509 6183 -7475
rect 6221 -7509 6249 -7475
rect 6249 -7509 6255 -7475
rect 6293 -7509 6317 -7475
rect 6317 -7509 6327 -7475
rect 6365 -7509 6385 -7475
rect 6385 -7509 6399 -7475
rect 6437 -7509 6453 -7475
rect 6453 -7509 6471 -7475
rect 6509 -7509 6521 -7475
rect 6521 -7509 6543 -7475
rect 6581 -7509 6589 -7475
rect 6589 -7509 6615 -7475
rect 6653 -7509 6657 -7475
rect 6657 -7509 6687 -7475
rect 6725 -7509 6759 -7475
rect 6797 -7509 6827 -7475
rect 6827 -7509 6831 -7475
rect 6869 -7509 6895 -7475
rect 6895 -7509 6903 -7475
rect 6941 -7509 6963 -7475
rect 6963 -7509 6975 -7475
rect 7013 -7509 7031 -7475
rect 7031 -7509 7047 -7475
rect 7085 -7509 7099 -7475
rect 7099 -7509 7119 -7475
rect 7157 -7509 7167 -7475
rect 7167 -7509 7191 -7475
rect 7229 -7509 7235 -7475
rect 7235 -7509 7263 -7475
rect 7301 -7509 7303 -7475
rect 7303 -7509 7335 -7475
rect 7373 -7509 7405 -7475
rect 7405 -7509 7407 -7475
rect 7445 -7509 7473 -7475
rect 7473 -7509 7479 -7475
rect 7517 -7509 7541 -7475
rect 7541 -7509 7551 -7475
rect 7589 -7509 7609 -7475
rect 7609 -7509 7623 -7475
rect 7661 -7509 7677 -7475
rect 7677 -7509 7695 -7475
rect 7733 -7509 7745 -7475
rect 7745 -7509 7767 -7475
rect 7805 -7509 7813 -7475
rect 7813 -7509 7839 -7475
rect 7877 -7509 7881 -7475
rect 7881 -7509 7911 -7475
rect 7949 -7509 7983 -7475
rect 8021 -7509 8051 -7475
rect 8051 -7509 8055 -7475
rect 8093 -7509 8119 -7475
rect 8119 -7509 8127 -7475
rect 8165 -7509 8187 -7475
rect 8187 -7509 8199 -7475
rect 8237 -7509 8255 -7475
rect 8255 -7509 8271 -7475
rect 8309 -7509 8323 -7475
rect 8323 -7509 8343 -7475
rect 8381 -7509 8391 -7475
rect 8391 -7509 8415 -7475
rect 8453 -7509 8459 -7475
rect 8459 -7509 8487 -7475
rect 8525 -7509 8527 -7475
rect 8527 -7509 8559 -7475
rect 8597 -7509 8629 -7475
rect 8629 -7509 8631 -7475
rect 8669 -7509 8697 -7475
rect 8697 -7509 8703 -7475
rect 8741 -7509 8765 -7475
rect 8765 -7509 8775 -7475
rect 8813 -7509 8833 -7475
rect 8833 -7509 8847 -7475
rect 8885 -7509 8901 -7475
rect 8901 -7509 8919 -7475
rect 8957 -7509 8969 -7475
rect 8969 -7509 8991 -7475
rect 9029 -7509 9037 -7475
rect 9037 -7509 9063 -7475
rect 9101 -7509 9105 -7475
rect 9105 -7509 9135 -7475
rect 9173 -7509 9207 -7475
rect 9245 -7509 9275 -7475
rect 9275 -7509 9279 -7475
rect 9317 -7509 9343 -7475
rect 9343 -7509 9351 -7475
rect 9389 -7509 9411 -7475
rect 9411 -7509 9423 -7475
rect 9461 -7509 9479 -7475
rect 9479 -7509 9495 -7475
rect 9533 -7509 9547 -7475
rect 9547 -7509 9567 -7475
rect 9605 -7509 9615 -7475
rect 9615 -7509 9639 -7475
rect 9677 -7509 9683 -7475
rect 9683 -7509 9711 -7475
rect 9749 -7509 9751 -7475
rect 9751 -7509 9783 -7475
rect 9821 -7509 9853 -7475
rect 9853 -7509 9855 -7475
rect 9893 -7509 9921 -7475
rect 9921 -7509 9927 -7475
rect 9965 -7509 9989 -7475
rect 9989 -7509 9999 -7475
rect 10037 -7509 10057 -7475
rect 10057 -7509 10071 -7475
rect 10109 -7509 10125 -7475
rect 10125 -7509 10143 -7475
rect 10181 -7509 10193 -7475
rect 10193 -7509 10215 -7475
rect 10253 -7509 10261 -7475
rect 10261 -7509 10287 -7475
rect 10325 -7509 10329 -7475
rect 10329 -7509 10359 -7475
rect 10397 -7509 10431 -7475
rect 10469 -7509 10499 -7475
rect 10499 -7509 10503 -7475
rect 10541 -7509 10567 -7475
rect 10567 -7509 10575 -7475
rect 10613 -7509 10635 -7475
rect 10635 -7509 10647 -7475
rect 10685 -7509 10703 -7475
rect 10703 -7509 10719 -7475
rect 10757 -7509 10771 -7475
rect 10771 -7509 10791 -7475
rect 10829 -7509 10839 -7475
rect 10839 -7509 10863 -7475
rect 10901 -7509 10907 -7475
rect 10907 -7509 10935 -7475
rect 10973 -7509 10975 -7475
rect 10975 -7509 11007 -7475
rect 11045 -7509 11077 -7475
rect 11077 -7509 11079 -7475
rect 11117 -7509 11145 -7475
rect 11145 -7509 11151 -7475
rect 11189 -7509 11213 -7475
rect 11213 -7509 11223 -7475
rect 11261 -7509 11281 -7475
rect 11281 -7509 11295 -7475
rect 11333 -7509 11349 -7475
rect 11349 -7509 11367 -7475
rect 11405 -7509 11417 -7475
rect 11417 -7509 11439 -7475
rect 11477 -7509 11485 -7475
rect 11485 -7509 11511 -7475
rect 11549 -7509 11553 -7475
rect 11553 -7509 11583 -7475
rect 11621 -7509 11655 -7475
rect 11693 -7509 11723 -7475
rect 11723 -7509 11727 -7475
rect 11765 -7509 11791 -7475
rect 11791 -7509 11799 -7475
rect 11837 -7509 11859 -7475
rect 11859 -7509 11871 -7475
rect 11909 -7509 11927 -7475
rect 11927 -7509 11943 -7475
rect 11981 -7509 11995 -7475
rect 11995 -7509 12015 -7475
rect 12053 -7509 12063 -7475
rect 12063 -7509 12087 -7475
rect 12125 -7509 12131 -7475
rect 12131 -7509 12159 -7475
rect 12197 -7509 12199 -7475
rect 12199 -7509 12231 -7475
rect 12269 -7509 12301 -7475
rect 12301 -7509 12303 -7475
rect 12341 -7509 12369 -7475
rect 12369 -7509 12375 -7475
rect 12413 -7509 12437 -7475
rect 12437 -7509 12447 -7475
rect 12485 -7509 12519 -7475
rect -259 -7845 -225 -7811
rect -187 -7845 -177 -7811
rect -177 -7845 -153 -7811
rect -115 -7845 -109 -7811
rect -109 -7845 -81 -7811
rect -43 -7845 -41 -7811
rect -41 -7845 -9 -7811
rect 29 -7845 61 -7811
rect 61 -7845 63 -7811
rect 101 -7845 129 -7811
rect 129 -7845 135 -7811
rect 173 -7845 197 -7811
rect 197 -7845 207 -7811
rect 245 -7845 265 -7811
rect 265 -7845 279 -7811
rect 317 -7845 333 -7811
rect 333 -7845 351 -7811
rect 389 -7845 401 -7811
rect 401 -7845 423 -7811
rect 461 -7845 469 -7811
rect 469 -7845 495 -7811
rect 533 -7845 537 -7811
rect 537 -7845 567 -7811
rect 605 -7845 639 -7811
rect 677 -7845 707 -7811
rect 707 -7845 711 -7811
rect 749 -7845 775 -7811
rect 775 -7845 783 -7811
rect 821 -7845 843 -7811
rect 843 -7845 855 -7811
rect 893 -7845 911 -7811
rect 911 -7845 927 -7811
rect 965 -7845 979 -7811
rect 979 -7845 999 -7811
rect 1037 -7845 1047 -7811
rect 1047 -7845 1071 -7811
rect 1109 -7845 1115 -7811
rect 1115 -7845 1143 -7811
rect 1181 -7845 1183 -7811
rect 1183 -7845 1215 -7811
rect 1253 -7845 1285 -7811
rect 1285 -7845 1287 -7811
rect 1325 -7845 1353 -7811
rect 1353 -7845 1359 -7811
rect 1397 -7845 1421 -7811
rect 1421 -7845 1431 -7811
rect 1469 -7845 1489 -7811
rect 1489 -7845 1503 -7811
rect 1541 -7845 1557 -7811
rect 1557 -7845 1575 -7811
rect 1613 -7845 1625 -7811
rect 1625 -7845 1647 -7811
rect 1685 -7845 1693 -7811
rect 1693 -7845 1719 -7811
rect 1757 -7845 1761 -7811
rect 1761 -7845 1791 -7811
rect 1829 -7845 1863 -7811
rect 1901 -7845 1931 -7811
rect 1931 -7845 1935 -7811
rect 1973 -7845 1999 -7811
rect 1999 -7845 2007 -7811
rect 2045 -7845 2067 -7811
rect 2067 -7845 2079 -7811
rect 2117 -7845 2135 -7811
rect 2135 -7845 2151 -7811
rect 2189 -7845 2203 -7811
rect 2203 -7845 2223 -7811
rect 2261 -7845 2271 -7811
rect 2271 -7845 2295 -7811
rect 2333 -7845 2339 -7811
rect 2339 -7845 2367 -7811
rect 2405 -7845 2407 -7811
rect 2407 -7845 2439 -7811
rect 2477 -7845 2509 -7811
rect 2509 -7845 2511 -7811
rect 2549 -7845 2577 -7811
rect 2577 -7845 2583 -7811
rect 2621 -7845 2645 -7811
rect 2645 -7845 2655 -7811
rect 2693 -7845 2713 -7811
rect 2713 -7845 2727 -7811
rect 2765 -7845 2781 -7811
rect 2781 -7845 2799 -7811
rect 2837 -7845 2849 -7811
rect 2849 -7845 2871 -7811
rect 2909 -7845 2917 -7811
rect 2917 -7845 2943 -7811
rect 2981 -7845 2985 -7811
rect 2985 -7845 3015 -7811
rect 3053 -7845 3087 -7811
rect 3125 -7845 3155 -7811
rect 3155 -7845 3159 -7811
rect 3197 -7845 3223 -7811
rect 3223 -7845 3231 -7811
rect 3269 -7845 3291 -7811
rect 3291 -7845 3303 -7811
rect 3341 -7845 3359 -7811
rect 3359 -7845 3375 -7811
rect 3413 -7845 3427 -7811
rect 3427 -7845 3447 -7811
rect 3485 -7845 3495 -7811
rect 3495 -7845 3519 -7811
rect 3557 -7845 3563 -7811
rect 3563 -7845 3591 -7811
rect 3629 -7845 3631 -7811
rect 3631 -7845 3663 -7811
rect 3701 -7845 3733 -7811
rect 3733 -7845 3735 -7811
rect 3773 -7845 3801 -7811
rect 3801 -7845 3807 -7811
rect 3845 -7845 3869 -7811
rect 3869 -7845 3879 -7811
rect 3917 -7845 3937 -7811
rect 3937 -7845 3951 -7811
rect 3989 -7845 4005 -7811
rect 4005 -7845 4023 -7811
rect 4061 -7845 4073 -7811
rect 4073 -7845 4095 -7811
rect 4133 -7845 4141 -7811
rect 4141 -7845 4167 -7811
rect 4205 -7845 4209 -7811
rect 4209 -7845 4239 -7811
rect 4277 -7845 4311 -7811
rect 4349 -7845 4379 -7811
rect 4379 -7845 4383 -7811
rect 4421 -7845 4447 -7811
rect 4447 -7845 4455 -7811
rect 4493 -7845 4515 -7811
rect 4515 -7845 4527 -7811
rect 4565 -7845 4583 -7811
rect 4583 -7845 4599 -7811
rect 4637 -7845 4651 -7811
rect 4651 -7845 4671 -7811
rect 4709 -7845 4719 -7811
rect 4719 -7845 4743 -7811
rect 4781 -7845 4787 -7811
rect 4787 -7845 4815 -7811
rect 4853 -7845 4855 -7811
rect 4855 -7845 4887 -7811
rect 4925 -7845 4957 -7811
rect 4957 -7845 4959 -7811
rect 4997 -7845 5025 -7811
rect 5025 -7845 5031 -7811
rect 5069 -7845 5093 -7811
rect 5093 -7845 5103 -7811
rect 5141 -7845 5161 -7811
rect 5161 -7845 5175 -7811
rect 5213 -7845 5229 -7811
rect 5229 -7845 5247 -7811
rect 5285 -7845 5297 -7811
rect 5297 -7845 5319 -7811
rect 5357 -7845 5365 -7811
rect 5365 -7845 5391 -7811
rect 5429 -7845 5433 -7811
rect 5433 -7845 5463 -7811
rect 5501 -7845 5535 -7811
rect 5573 -7845 5603 -7811
rect 5603 -7845 5607 -7811
rect 5645 -7845 5671 -7811
rect 5671 -7845 5679 -7811
rect 5717 -7845 5739 -7811
rect 5739 -7845 5751 -7811
rect 5789 -7845 5807 -7811
rect 5807 -7845 5823 -7811
rect 5861 -7845 5875 -7811
rect 5875 -7845 5895 -7811
rect 5933 -7845 5943 -7811
rect 5943 -7845 5967 -7811
rect 6005 -7845 6011 -7811
rect 6011 -7845 6039 -7811
rect 6077 -7845 6079 -7811
rect 6079 -7845 6111 -7811
rect 6149 -7845 6181 -7811
rect 6181 -7845 6183 -7811
rect 6221 -7845 6249 -7811
rect 6249 -7845 6255 -7811
rect 6293 -7845 6317 -7811
rect 6317 -7845 6327 -7811
rect 6365 -7845 6385 -7811
rect 6385 -7845 6399 -7811
rect 6437 -7845 6453 -7811
rect 6453 -7845 6471 -7811
rect 6509 -7845 6521 -7811
rect 6521 -7845 6543 -7811
rect 6581 -7845 6589 -7811
rect 6589 -7845 6615 -7811
rect 6653 -7845 6657 -7811
rect 6657 -7845 6687 -7811
rect 6725 -7845 6759 -7811
rect 6797 -7845 6827 -7811
rect 6827 -7845 6831 -7811
rect 6869 -7845 6895 -7811
rect 6895 -7845 6903 -7811
rect 6941 -7845 6963 -7811
rect 6963 -7845 6975 -7811
rect 7013 -7845 7031 -7811
rect 7031 -7845 7047 -7811
rect 7085 -7845 7099 -7811
rect 7099 -7845 7119 -7811
rect 7157 -7845 7167 -7811
rect 7167 -7845 7191 -7811
rect 7229 -7845 7235 -7811
rect 7235 -7845 7263 -7811
rect 7301 -7845 7303 -7811
rect 7303 -7845 7335 -7811
rect 7373 -7845 7405 -7811
rect 7405 -7845 7407 -7811
rect 7445 -7845 7473 -7811
rect 7473 -7845 7479 -7811
rect 7517 -7845 7541 -7811
rect 7541 -7845 7551 -7811
rect 7589 -7845 7609 -7811
rect 7609 -7845 7623 -7811
rect 7661 -7845 7677 -7811
rect 7677 -7845 7695 -7811
rect 7733 -7845 7745 -7811
rect 7745 -7845 7767 -7811
rect 7805 -7845 7813 -7811
rect 7813 -7845 7839 -7811
rect 7877 -7845 7881 -7811
rect 7881 -7845 7911 -7811
rect 7949 -7845 7983 -7811
rect 8021 -7845 8051 -7811
rect 8051 -7845 8055 -7811
rect 8093 -7845 8119 -7811
rect 8119 -7845 8127 -7811
rect 8165 -7845 8187 -7811
rect 8187 -7845 8199 -7811
rect 8237 -7845 8255 -7811
rect 8255 -7845 8271 -7811
rect 8309 -7845 8323 -7811
rect 8323 -7845 8343 -7811
rect 8381 -7845 8391 -7811
rect 8391 -7845 8415 -7811
rect 8453 -7845 8459 -7811
rect 8459 -7845 8487 -7811
rect 8525 -7845 8527 -7811
rect 8527 -7845 8559 -7811
rect 8597 -7845 8629 -7811
rect 8629 -7845 8631 -7811
rect 8669 -7845 8697 -7811
rect 8697 -7845 8703 -7811
rect 8741 -7845 8765 -7811
rect 8765 -7845 8775 -7811
rect 8813 -7845 8833 -7811
rect 8833 -7845 8847 -7811
rect 8885 -7845 8901 -7811
rect 8901 -7845 8919 -7811
rect 8957 -7845 8969 -7811
rect 8969 -7845 8991 -7811
rect 9029 -7845 9037 -7811
rect 9037 -7845 9063 -7811
rect 9101 -7845 9105 -7811
rect 9105 -7845 9135 -7811
rect 9173 -7845 9207 -7811
rect 9245 -7845 9275 -7811
rect 9275 -7845 9279 -7811
rect 9317 -7845 9343 -7811
rect 9343 -7845 9351 -7811
rect 9389 -7845 9411 -7811
rect 9411 -7845 9423 -7811
rect 9461 -7845 9479 -7811
rect 9479 -7845 9495 -7811
rect 9533 -7845 9547 -7811
rect 9547 -7845 9567 -7811
rect 9605 -7845 9615 -7811
rect 9615 -7845 9639 -7811
rect 9677 -7845 9683 -7811
rect 9683 -7845 9711 -7811
rect 9749 -7845 9751 -7811
rect 9751 -7845 9783 -7811
rect 9821 -7845 9853 -7811
rect 9853 -7845 9855 -7811
rect 9893 -7845 9921 -7811
rect 9921 -7845 9927 -7811
rect 9965 -7845 9989 -7811
rect 9989 -7845 9999 -7811
rect 10037 -7845 10057 -7811
rect 10057 -7845 10071 -7811
rect 10109 -7845 10125 -7811
rect 10125 -7845 10143 -7811
rect 10181 -7845 10193 -7811
rect 10193 -7845 10215 -7811
rect 10253 -7845 10261 -7811
rect 10261 -7845 10287 -7811
rect 10325 -7845 10329 -7811
rect 10329 -7845 10359 -7811
rect 10397 -7845 10431 -7811
rect 10469 -7845 10499 -7811
rect 10499 -7845 10503 -7811
rect 10541 -7845 10567 -7811
rect 10567 -7845 10575 -7811
rect 10613 -7845 10635 -7811
rect 10635 -7845 10647 -7811
rect 10685 -7845 10703 -7811
rect 10703 -7845 10719 -7811
rect 10757 -7845 10771 -7811
rect 10771 -7845 10791 -7811
rect 10829 -7845 10839 -7811
rect 10839 -7845 10863 -7811
rect 10901 -7845 10907 -7811
rect 10907 -7845 10935 -7811
rect 10973 -7845 10975 -7811
rect 10975 -7845 11007 -7811
rect 11045 -7845 11077 -7811
rect 11077 -7845 11079 -7811
rect 11117 -7845 11145 -7811
rect 11145 -7845 11151 -7811
rect 11189 -7845 11213 -7811
rect 11213 -7845 11223 -7811
rect 11261 -7845 11281 -7811
rect 11281 -7845 11295 -7811
rect 11333 -7845 11349 -7811
rect 11349 -7845 11367 -7811
rect 11405 -7845 11417 -7811
rect 11417 -7845 11439 -7811
rect 11477 -7845 11485 -7811
rect 11485 -7845 11511 -7811
rect 11549 -7845 11553 -7811
rect 11553 -7845 11583 -7811
rect 11621 -7845 11655 -7811
rect 11693 -7845 11723 -7811
rect 11723 -7845 11727 -7811
rect 11765 -7845 11791 -7811
rect 11791 -7845 11799 -7811
rect 11837 -7845 11859 -7811
rect 11859 -7845 11871 -7811
rect 11909 -7845 11927 -7811
rect 11927 -7845 11943 -7811
rect 11981 -7845 11995 -7811
rect 11995 -7845 12015 -7811
rect 12053 -7845 12063 -7811
rect 12063 -7845 12087 -7811
rect 12125 -7845 12131 -7811
rect 12131 -7845 12159 -7811
rect 12197 -7845 12199 -7811
rect 12199 -7845 12231 -7811
rect 12269 -7845 12301 -7811
rect 12301 -7845 12303 -7811
rect 12341 -7845 12369 -7811
rect 12369 -7845 12375 -7811
rect 12413 -7845 12437 -7811
rect 12437 -7845 12447 -7811
rect 12485 -7845 12519 -7811
rect -329 -8025 -295 -7999
rect -329 -8033 -295 -8025
rect -329 -8093 -295 -8071
rect -329 -8105 -295 -8093
rect -329 -8161 -295 -8143
rect -329 -8177 -295 -8161
rect -329 -8229 -295 -8215
rect -329 -8249 -295 -8229
rect -329 -8297 -295 -8287
rect -329 -8321 -295 -8297
rect -329 -8365 -295 -8359
rect -329 -8393 -295 -8365
rect -329 -8433 -295 -8431
rect -329 -8465 -295 -8433
rect -329 -8535 -295 -8503
rect -329 -8537 -295 -8535
rect -329 -8603 -295 -8575
rect -329 -8609 -295 -8603
rect -329 -8671 -295 -8647
rect -329 -8681 -295 -8671
rect -329 -8739 -295 -8719
rect -329 -8753 -295 -8739
rect -329 -8807 -295 -8791
rect -329 -8825 -295 -8807
rect -329 -8875 -295 -8863
rect -329 -8897 -295 -8875
rect -329 -8943 -295 -8935
rect -329 -8969 -295 -8943
rect -329 -9011 -295 -9007
rect -329 -9041 -295 -9011
rect -329 -9113 -295 -9079
rect -329 -9181 -295 -9151
rect -329 -9185 -295 -9181
rect -329 -9249 -295 -9223
rect -329 -9257 -295 -9249
rect -329 -9317 -295 -9295
rect -329 -9329 -295 -9317
rect -329 -9385 -295 -9367
rect -329 -9401 -295 -9385
rect -329 -9453 -295 -9439
rect -329 -9473 -295 -9453
rect -329 -9521 -295 -9511
rect -329 -9545 -295 -9521
rect -329 -9589 -295 -9583
rect -329 -9617 -295 -9589
rect -329 -9657 -295 -9655
rect -329 -9689 -295 -9657
rect -329 -9759 -295 -9727
rect -329 -9761 -295 -9759
rect -329 -9827 -295 -9799
rect -329 -9833 -295 -9827
rect -329 -9895 -295 -9871
rect -329 -9905 -295 -9895
rect -329 -9963 -295 -9943
rect -329 -9977 -295 -9963
rect -329 -10031 -295 -10015
rect -329 -10049 -295 -10031
rect -329 -10099 -295 -10087
rect -329 -10121 -295 -10099
rect -329 -10167 -295 -10159
rect -329 -10193 -295 -10167
rect -329 -10235 -295 -10231
rect -329 -10265 -295 -10235
rect -329 -10337 -295 -10303
rect -329 -10405 -295 -10375
rect -329 -10409 -295 -10405
rect -329 -10473 -295 -10447
rect -329 -10481 -295 -10473
rect -329 -10541 -295 -10519
rect -329 -10553 -295 -10541
rect 12555 -8025 12589 -7999
rect 12555 -8033 12589 -8025
rect 12555 -8093 12589 -8071
rect 12555 -8105 12589 -8093
rect 12555 -8161 12589 -8143
rect 12555 -8177 12589 -8161
rect 12555 -8229 12589 -8215
rect 12555 -8249 12589 -8229
rect 12555 -8297 12589 -8287
rect 12555 -8321 12589 -8297
rect 12555 -8365 12589 -8359
rect 12555 -8393 12589 -8365
rect 12555 -8433 12589 -8431
rect 12555 -8465 12589 -8433
rect 12555 -8535 12589 -8503
rect 12555 -8537 12589 -8535
rect 12555 -8603 12589 -8575
rect 12555 -8609 12589 -8603
rect 12555 -8671 12589 -8647
rect 12555 -8681 12589 -8671
rect 12555 -8739 12589 -8719
rect 12555 -8753 12589 -8739
rect 12555 -8807 12589 -8791
rect 12555 -8825 12589 -8807
rect 12555 -8875 12589 -8863
rect 12555 -8897 12589 -8875
rect 12555 -8943 12589 -8935
rect 12555 -8969 12589 -8943
rect 12555 -9011 12589 -9007
rect 12555 -9041 12589 -9011
rect 12555 -9113 12589 -9079
rect 12555 -9181 12589 -9151
rect 12555 -9185 12589 -9181
rect 12555 -9249 12589 -9223
rect 12555 -9257 12589 -9249
rect 12555 -9317 12589 -9295
rect 12555 -9329 12589 -9317
rect 12555 -9385 12589 -9367
rect 12555 -9401 12589 -9385
rect 12555 -9453 12589 -9439
rect 12555 -9473 12589 -9453
rect 12555 -9521 12589 -9511
rect 12555 -9545 12589 -9521
rect 12555 -9589 12589 -9583
rect 12555 -9617 12589 -9589
rect 12555 -9657 12589 -9655
rect 12555 -9689 12589 -9657
rect 12555 -9759 12589 -9727
rect 12555 -9761 12589 -9759
rect 12555 -9827 12589 -9799
rect 12555 -9833 12589 -9827
rect 12555 -9895 12589 -9871
rect 12555 -9905 12589 -9895
rect 12555 -9963 12589 -9943
rect 12555 -9977 12589 -9963
rect 12555 -10031 12589 -10015
rect 12555 -10049 12589 -10031
rect 12555 -10099 12589 -10087
rect 12555 -10121 12589 -10099
rect 12555 -10167 12589 -10159
rect 12555 -10193 12589 -10167
rect 12555 -10235 12589 -10231
rect 12555 -10265 12589 -10235
rect 12555 -10337 12589 -10303
rect 12555 -10405 12589 -10375
rect 12555 -10409 12589 -10405
rect 12555 -10473 12589 -10447
rect 12555 -10481 12589 -10473
rect 12555 -10541 12589 -10519
rect 12555 -10553 12589 -10541
rect -259 -10789 -225 -10755
rect -187 -10789 -177 -10755
rect -177 -10789 -153 -10755
rect -115 -10789 -109 -10755
rect -109 -10789 -81 -10755
rect -43 -10789 -41 -10755
rect -41 -10789 -9 -10755
rect 29 -10789 61 -10755
rect 61 -10789 63 -10755
rect 101 -10789 129 -10755
rect 129 -10789 135 -10755
rect 173 -10789 197 -10755
rect 197 -10789 207 -10755
rect 245 -10789 265 -10755
rect 265 -10789 279 -10755
rect 317 -10789 333 -10755
rect 333 -10789 351 -10755
rect 389 -10789 401 -10755
rect 401 -10789 423 -10755
rect 461 -10789 469 -10755
rect 469 -10789 495 -10755
rect 533 -10789 537 -10755
rect 537 -10789 567 -10755
rect 605 -10789 639 -10755
rect 677 -10789 707 -10755
rect 707 -10789 711 -10755
rect 749 -10789 775 -10755
rect 775 -10789 783 -10755
rect 821 -10789 843 -10755
rect 843 -10789 855 -10755
rect 893 -10789 911 -10755
rect 911 -10789 927 -10755
rect 965 -10789 979 -10755
rect 979 -10789 999 -10755
rect 1037 -10789 1047 -10755
rect 1047 -10789 1071 -10755
rect 1109 -10789 1115 -10755
rect 1115 -10789 1143 -10755
rect 1181 -10789 1183 -10755
rect 1183 -10789 1215 -10755
rect 1253 -10789 1285 -10755
rect 1285 -10789 1287 -10755
rect 1325 -10789 1353 -10755
rect 1353 -10789 1359 -10755
rect 1397 -10789 1421 -10755
rect 1421 -10789 1431 -10755
rect 1469 -10789 1489 -10755
rect 1489 -10789 1503 -10755
rect 1541 -10789 1557 -10755
rect 1557 -10789 1575 -10755
rect 1613 -10789 1625 -10755
rect 1625 -10789 1647 -10755
rect 1685 -10789 1693 -10755
rect 1693 -10789 1719 -10755
rect 1757 -10789 1761 -10755
rect 1761 -10789 1791 -10755
rect 1829 -10789 1863 -10755
rect 1901 -10789 1931 -10755
rect 1931 -10789 1935 -10755
rect 1973 -10789 1999 -10755
rect 1999 -10789 2007 -10755
rect 2045 -10789 2067 -10755
rect 2067 -10789 2079 -10755
rect 2117 -10789 2135 -10755
rect 2135 -10789 2151 -10755
rect 2189 -10789 2203 -10755
rect 2203 -10789 2223 -10755
rect 2261 -10789 2271 -10755
rect 2271 -10789 2295 -10755
rect 2333 -10789 2339 -10755
rect 2339 -10789 2367 -10755
rect 2405 -10789 2407 -10755
rect 2407 -10789 2439 -10755
rect 2477 -10789 2509 -10755
rect 2509 -10789 2511 -10755
rect 2549 -10789 2577 -10755
rect 2577 -10789 2583 -10755
rect 2621 -10789 2645 -10755
rect 2645 -10789 2655 -10755
rect 2693 -10789 2713 -10755
rect 2713 -10789 2727 -10755
rect 2765 -10789 2781 -10755
rect 2781 -10789 2799 -10755
rect 2837 -10789 2849 -10755
rect 2849 -10789 2871 -10755
rect 2909 -10789 2917 -10755
rect 2917 -10789 2943 -10755
rect 2981 -10789 2985 -10755
rect 2985 -10789 3015 -10755
rect 3053 -10789 3087 -10755
rect 3125 -10789 3155 -10755
rect 3155 -10789 3159 -10755
rect 3197 -10789 3223 -10755
rect 3223 -10789 3231 -10755
rect 3269 -10789 3291 -10755
rect 3291 -10789 3303 -10755
rect 3341 -10789 3359 -10755
rect 3359 -10789 3375 -10755
rect 3413 -10789 3427 -10755
rect 3427 -10789 3447 -10755
rect 3485 -10789 3495 -10755
rect 3495 -10789 3519 -10755
rect 3557 -10789 3563 -10755
rect 3563 -10789 3591 -10755
rect 3629 -10789 3631 -10755
rect 3631 -10789 3663 -10755
rect 3701 -10789 3733 -10755
rect 3733 -10789 3735 -10755
rect 3773 -10789 3801 -10755
rect 3801 -10789 3807 -10755
rect 3845 -10789 3869 -10755
rect 3869 -10789 3879 -10755
rect 3917 -10789 3937 -10755
rect 3937 -10789 3951 -10755
rect 3989 -10789 4005 -10755
rect 4005 -10789 4023 -10755
rect 4061 -10789 4073 -10755
rect 4073 -10789 4095 -10755
rect 4133 -10789 4141 -10755
rect 4141 -10789 4167 -10755
rect 4205 -10789 4209 -10755
rect 4209 -10789 4239 -10755
rect 4277 -10789 4311 -10755
rect 4349 -10789 4379 -10755
rect 4379 -10789 4383 -10755
rect 4421 -10789 4447 -10755
rect 4447 -10789 4455 -10755
rect 4493 -10789 4515 -10755
rect 4515 -10789 4527 -10755
rect 4565 -10789 4583 -10755
rect 4583 -10789 4599 -10755
rect 4637 -10789 4651 -10755
rect 4651 -10789 4671 -10755
rect 4709 -10789 4719 -10755
rect 4719 -10789 4743 -10755
rect 4781 -10789 4787 -10755
rect 4787 -10789 4815 -10755
rect 4853 -10789 4855 -10755
rect 4855 -10789 4887 -10755
rect 4925 -10789 4957 -10755
rect 4957 -10789 4959 -10755
rect 4997 -10789 5025 -10755
rect 5025 -10789 5031 -10755
rect 5069 -10789 5093 -10755
rect 5093 -10789 5103 -10755
rect 5141 -10789 5161 -10755
rect 5161 -10789 5175 -10755
rect 5213 -10789 5229 -10755
rect 5229 -10789 5247 -10755
rect 5285 -10789 5297 -10755
rect 5297 -10789 5319 -10755
rect 5357 -10789 5365 -10755
rect 5365 -10789 5391 -10755
rect 5429 -10789 5433 -10755
rect 5433 -10789 5463 -10755
rect 5501 -10789 5535 -10755
rect 5573 -10789 5603 -10755
rect 5603 -10789 5607 -10755
rect 5645 -10789 5671 -10755
rect 5671 -10789 5679 -10755
rect 5717 -10789 5739 -10755
rect 5739 -10789 5751 -10755
rect 5789 -10789 5807 -10755
rect 5807 -10789 5823 -10755
rect 5861 -10789 5875 -10755
rect 5875 -10789 5895 -10755
rect 5933 -10789 5943 -10755
rect 5943 -10789 5967 -10755
rect 6005 -10789 6011 -10755
rect 6011 -10789 6039 -10755
rect 6077 -10789 6079 -10755
rect 6079 -10789 6111 -10755
rect 6149 -10789 6181 -10755
rect 6181 -10789 6183 -10755
rect 6221 -10789 6249 -10755
rect 6249 -10789 6255 -10755
rect 6293 -10789 6317 -10755
rect 6317 -10789 6327 -10755
rect 6365 -10789 6385 -10755
rect 6385 -10789 6399 -10755
rect 6437 -10789 6453 -10755
rect 6453 -10789 6471 -10755
rect 6509 -10789 6521 -10755
rect 6521 -10789 6543 -10755
rect 6581 -10789 6589 -10755
rect 6589 -10789 6615 -10755
rect 6653 -10789 6657 -10755
rect 6657 -10789 6687 -10755
rect 6725 -10789 6759 -10755
rect 6797 -10789 6827 -10755
rect 6827 -10789 6831 -10755
rect 6869 -10789 6895 -10755
rect 6895 -10789 6903 -10755
rect 6941 -10789 6963 -10755
rect 6963 -10789 6975 -10755
rect 7013 -10789 7031 -10755
rect 7031 -10789 7047 -10755
rect 7085 -10789 7099 -10755
rect 7099 -10789 7119 -10755
rect 7157 -10789 7167 -10755
rect 7167 -10789 7191 -10755
rect 7229 -10789 7235 -10755
rect 7235 -10789 7263 -10755
rect 7301 -10789 7303 -10755
rect 7303 -10789 7335 -10755
rect 7373 -10789 7405 -10755
rect 7405 -10789 7407 -10755
rect 7445 -10789 7473 -10755
rect 7473 -10789 7479 -10755
rect 7517 -10789 7541 -10755
rect 7541 -10789 7551 -10755
rect 7589 -10789 7609 -10755
rect 7609 -10789 7623 -10755
rect 7661 -10789 7677 -10755
rect 7677 -10789 7695 -10755
rect 7733 -10789 7745 -10755
rect 7745 -10789 7767 -10755
rect 7805 -10789 7813 -10755
rect 7813 -10789 7839 -10755
rect 7877 -10789 7881 -10755
rect 7881 -10789 7911 -10755
rect 7949 -10789 7983 -10755
rect 8021 -10789 8051 -10755
rect 8051 -10789 8055 -10755
rect 8093 -10789 8119 -10755
rect 8119 -10789 8127 -10755
rect 8165 -10789 8187 -10755
rect 8187 -10789 8199 -10755
rect 8237 -10789 8255 -10755
rect 8255 -10789 8271 -10755
rect 8309 -10789 8323 -10755
rect 8323 -10789 8343 -10755
rect 8381 -10789 8391 -10755
rect 8391 -10789 8415 -10755
rect 8453 -10789 8459 -10755
rect 8459 -10789 8487 -10755
rect 8525 -10789 8527 -10755
rect 8527 -10789 8559 -10755
rect 8597 -10789 8629 -10755
rect 8629 -10789 8631 -10755
rect 8669 -10789 8697 -10755
rect 8697 -10789 8703 -10755
rect 8741 -10789 8765 -10755
rect 8765 -10789 8775 -10755
rect 8813 -10789 8833 -10755
rect 8833 -10789 8847 -10755
rect 8885 -10789 8901 -10755
rect 8901 -10789 8919 -10755
rect 8957 -10789 8969 -10755
rect 8969 -10789 8991 -10755
rect 9029 -10789 9037 -10755
rect 9037 -10789 9063 -10755
rect 9101 -10789 9105 -10755
rect 9105 -10789 9135 -10755
rect 9173 -10789 9207 -10755
rect 9245 -10789 9275 -10755
rect 9275 -10789 9279 -10755
rect 9317 -10789 9343 -10755
rect 9343 -10789 9351 -10755
rect 9389 -10789 9411 -10755
rect 9411 -10789 9423 -10755
rect 9461 -10789 9479 -10755
rect 9479 -10789 9495 -10755
rect 9533 -10789 9547 -10755
rect 9547 -10789 9567 -10755
rect 9605 -10789 9615 -10755
rect 9615 -10789 9639 -10755
rect 9677 -10789 9683 -10755
rect 9683 -10789 9711 -10755
rect 9749 -10789 9751 -10755
rect 9751 -10789 9783 -10755
rect 9821 -10789 9853 -10755
rect 9853 -10789 9855 -10755
rect 9893 -10789 9921 -10755
rect 9921 -10789 9927 -10755
rect 9965 -10789 9989 -10755
rect 9989 -10789 9999 -10755
rect 10037 -10789 10057 -10755
rect 10057 -10789 10071 -10755
rect 10109 -10789 10125 -10755
rect 10125 -10789 10143 -10755
rect 10181 -10789 10193 -10755
rect 10193 -10789 10215 -10755
rect 10253 -10789 10261 -10755
rect 10261 -10789 10287 -10755
rect 10325 -10789 10329 -10755
rect 10329 -10789 10359 -10755
rect 10397 -10789 10431 -10755
rect 10469 -10789 10499 -10755
rect 10499 -10789 10503 -10755
rect 10541 -10789 10567 -10755
rect 10567 -10789 10575 -10755
rect 10613 -10789 10635 -10755
rect 10635 -10789 10647 -10755
rect 10685 -10789 10703 -10755
rect 10703 -10789 10719 -10755
rect 10757 -10789 10771 -10755
rect 10771 -10789 10791 -10755
rect 10829 -10789 10839 -10755
rect 10839 -10789 10863 -10755
rect 10901 -10789 10907 -10755
rect 10907 -10789 10935 -10755
rect 10973 -10789 10975 -10755
rect 10975 -10789 11007 -10755
rect 11045 -10789 11077 -10755
rect 11077 -10789 11079 -10755
rect 11117 -10789 11145 -10755
rect 11145 -10789 11151 -10755
rect 11189 -10789 11213 -10755
rect 11213 -10789 11223 -10755
rect 11261 -10789 11281 -10755
rect 11281 -10789 11295 -10755
rect 11333 -10789 11349 -10755
rect 11349 -10789 11367 -10755
rect 11405 -10789 11417 -10755
rect 11417 -10789 11439 -10755
rect 11477 -10789 11485 -10755
rect 11485 -10789 11511 -10755
rect 11549 -10789 11553 -10755
rect 11553 -10789 11583 -10755
rect 11621 -10789 11655 -10755
rect 11693 -10789 11723 -10755
rect 11723 -10789 11727 -10755
rect 11765 -10789 11791 -10755
rect 11791 -10789 11799 -10755
rect 11837 -10789 11859 -10755
rect 11859 -10789 11871 -10755
rect 11909 -10789 11927 -10755
rect 11927 -10789 11943 -10755
rect 11981 -10789 11995 -10755
rect 11995 -10789 12015 -10755
rect 12053 -10789 12063 -10755
rect 12063 -10789 12087 -10755
rect 12125 -10789 12131 -10755
rect 12131 -10789 12159 -10755
rect 12197 -10789 12199 -10755
rect 12199 -10789 12231 -10755
rect 12269 -10789 12301 -10755
rect 12301 -10789 12303 -10755
rect 12341 -10789 12369 -10755
rect 12369 -10789 12375 -10755
rect 12413 -10789 12437 -10755
rect 12437 -10789 12447 -10755
rect 12485 -10789 12519 -10755
<< metal1 >>
rect -368 2889 12628 2928
rect -368 2855 -259 2889
rect -225 2855 -187 2889
rect -153 2855 -115 2889
rect -81 2855 -43 2889
rect -9 2855 29 2889
rect 63 2855 101 2889
rect 135 2855 173 2889
rect 207 2855 245 2889
rect 279 2855 317 2889
rect 351 2855 389 2889
rect 423 2855 461 2889
rect 495 2855 533 2889
rect 567 2855 605 2889
rect 639 2855 677 2889
rect 711 2855 749 2889
rect 783 2855 821 2889
rect 855 2855 893 2889
rect 927 2855 965 2889
rect 999 2855 1037 2889
rect 1071 2855 1109 2889
rect 1143 2855 1181 2889
rect 1215 2855 1253 2889
rect 1287 2855 1325 2889
rect 1359 2855 1397 2889
rect 1431 2855 1469 2889
rect 1503 2855 1541 2889
rect 1575 2855 1613 2889
rect 1647 2855 1685 2889
rect 1719 2855 1757 2889
rect 1791 2855 1829 2889
rect 1863 2855 1901 2889
rect 1935 2855 1973 2889
rect 2007 2855 2045 2889
rect 2079 2855 2117 2889
rect 2151 2855 2189 2889
rect 2223 2855 2261 2889
rect 2295 2855 2333 2889
rect 2367 2855 2405 2889
rect 2439 2855 2477 2889
rect 2511 2855 2549 2889
rect 2583 2855 2621 2889
rect 2655 2855 2693 2889
rect 2727 2855 2765 2889
rect 2799 2855 2837 2889
rect 2871 2855 2909 2889
rect 2943 2855 2981 2889
rect 3015 2855 3053 2889
rect 3087 2855 3125 2889
rect 3159 2855 3197 2889
rect 3231 2855 3269 2889
rect 3303 2855 3341 2889
rect 3375 2855 3413 2889
rect 3447 2855 3485 2889
rect 3519 2855 3557 2889
rect 3591 2855 3629 2889
rect 3663 2855 3701 2889
rect 3735 2855 3773 2889
rect 3807 2855 3845 2889
rect 3879 2855 3917 2889
rect 3951 2855 3989 2889
rect 4023 2855 4061 2889
rect 4095 2855 4133 2889
rect 4167 2855 4205 2889
rect 4239 2855 4277 2889
rect 4311 2855 4349 2889
rect 4383 2855 4421 2889
rect 4455 2855 4493 2889
rect 4527 2855 4565 2889
rect 4599 2855 4637 2889
rect 4671 2855 4709 2889
rect 4743 2855 4781 2889
rect 4815 2855 4853 2889
rect 4887 2855 4925 2889
rect 4959 2855 4997 2889
rect 5031 2855 5069 2889
rect 5103 2855 5141 2889
rect 5175 2855 5213 2889
rect 5247 2855 5285 2889
rect 5319 2855 5357 2889
rect 5391 2855 5429 2889
rect 5463 2855 5501 2889
rect 5535 2855 5573 2889
rect 5607 2855 5645 2889
rect 5679 2855 5717 2889
rect 5751 2855 5789 2889
rect 5823 2855 5861 2889
rect 5895 2855 5933 2889
rect 5967 2855 6005 2889
rect 6039 2855 6077 2889
rect 6111 2855 6149 2889
rect 6183 2855 6221 2889
rect 6255 2855 6293 2889
rect 6327 2855 6365 2889
rect 6399 2855 6437 2889
rect 6471 2855 6509 2889
rect 6543 2855 6581 2889
rect 6615 2855 6653 2889
rect 6687 2855 6725 2889
rect 6759 2855 6797 2889
rect 6831 2855 6869 2889
rect 6903 2855 6941 2889
rect 6975 2855 7013 2889
rect 7047 2855 7085 2889
rect 7119 2855 7157 2889
rect 7191 2855 7229 2889
rect 7263 2855 7301 2889
rect 7335 2855 7373 2889
rect 7407 2855 7445 2889
rect 7479 2855 7517 2889
rect 7551 2855 7589 2889
rect 7623 2855 7661 2889
rect 7695 2855 7733 2889
rect 7767 2855 7805 2889
rect 7839 2855 7877 2889
rect 7911 2855 7949 2889
rect 7983 2855 8021 2889
rect 8055 2855 8093 2889
rect 8127 2855 8165 2889
rect 8199 2855 8237 2889
rect 8271 2855 8309 2889
rect 8343 2855 8381 2889
rect 8415 2855 8453 2889
rect 8487 2855 8525 2889
rect 8559 2855 8597 2889
rect 8631 2855 8669 2889
rect 8703 2855 8741 2889
rect 8775 2855 8813 2889
rect 8847 2855 8885 2889
rect 8919 2855 8957 2889
rect 8991 2855 9029 2889
rect 9063 2855 9101 2889
rect 9135 2855 9173 2889
rect 9207 2855 9245 2889
rect 9279 2855 9317 2889
rect 9351 2855 9389 2889
rect 9423 2855 9461 2889
rect 9495 2855 9533 2889
rect 9567 2855 9605 2889
rect 9639 2855 9677 2889
rect 9711 2855 9749 2889
rect 9783 2855 9821 2889
rect 9855 2855 9893 2889
rect 9927 2855 9965 2889
rect 9999 2855 10037 2889
rect 10071 2855 10109 2889
rect 10143 2855 10181 2889
rect 10215 2855 10253 2889
rect 10287 2855 10325 2889
rect 10359 2855 10397 2889
rect 10431 2855 10469 2889
rect 10503 2855 10541 2889
rect 10575 2855 10613 2889
rect 10647 2855 10685 2889
rect 10719 2855 10757 2889
rect 10791 2855 10829 2889
rect 10863 2855 10901 2889
rect 10935 2855 10973 2889
rect 11007 2855 11045 2889
rect 11079 2855 11117 2889
rect 11151 2855 11189 2889
rect 11223 2855 11261 2889
rect 11295 2855 11333 2889
rect 11367 2855 11405 2889
rect 11439 2855 11477 2889
rect 11511 2855 11549 2889
rect 11583 2855 11621 2889
rect 11655 2855 11693 2889
rect 11727 2855 11765 2889
rect 11799 2855 11837 2889
rect 11871 2855 11909 2889
rect 11943 2855 11981 2889
rect 12015 2855 12053 2889
rect 12087 2855 12125 2889
rect 12159 2855 12197 2889
rect 12231 2855 12269 2889
rect 12303 2855 12341 2889
rect 12375 2855 12413 2889
rect 12447 2855 12485 2889
rect 12519 2855 12628 2889
rect -368 2816 12628 2855
rect -368 2788 354 2816
rect -368 2544 -238 2788
rect 326 2544 354 2788
rect -368 2516 354 2544
rect 11906 2788 12628 2816
rect 11906 2544 11934 2788
rect 12498 2544 12628 2788
rect 11906 2516 12628 2544
rect -368 2287 -256 2516
rect -368 2253 -329 2287
rect -295 2253 -256 2287
rect -368 2215 -256 2253
rect -368 2181 -329 2215
rect -295 2181 -256 2215
rect 110 2372 12310 2438
rect 110 2256 171 2372
rect 12255 2256 12310 2372
rect 110 2192 12310 2256
rect 12516 2287 12628 2516
rect 12516 2253 12555 2287
rect 12589 2253 12628 2287
rect 12516 2215 12628 2253
rect -368 2143 -256 2181
rect -368 2109 -329 2143
rect -295 2109 -256 2143
rect 172 2110 232 2192
rect 596 2110 656 2192
rect 1032 2110 1092 2192
rect 2746 2110 2806 2192
rect 4466 2110 4526 2192
rect 6174 2110 6234 2192
rect 7894 2110 7954 2192
rect 9608 2110 9668 2192
rect 11326 2110 11386 2192
rect 11754 2110 11814 2192
rect 12186 2110 12246 2192
rect 12516 2181 12555 2215
rect 12589 2181 12628 2215
rect 12516 2143 12628 2181
rect -368 2108 -256 2109
rect 166 2108 238 2110
rect -368 2106 238 2108
rect -368 2071 176 2106
rect -368 2037 -329 2071
rect -295 2054 176 2071
rect 228 2054 238 2106
rect -295 2050 238 2054
rect 590 2106 662 2110
rect 590 2054 600 2106
rect 652 2054 662 2106
rect 590 2050 662 2054
rect 1026 2106 1098 2110
rect 1026 2054 1036 2106
rect 1088 2054 1098 2106
rect 1026 2050 1098 2054
rect 2740 2106 2812 2110
rect 2740 2054 2750 2106
rect 2802 2054 2812 2106
rect 2740 2050 2812 2054
rect 4460 2106 4532 2110
rect 4460 2054 4470 2106
rect 4522 2054 4532 2106
rect 4460 2050 4532 2054
rect 6168 2106 6240 2110
rect 6168 2054 6178 2106
rect 6230 2054 6240 2106
rect 6168 2050 6240 2054
rect 7888 2106 7960 2110
rect 7888 2054 7898 2106
rect 7950 2054 7960 2106
rect 7888 2050 7960 2054
rect 9602 2106 9674 2110
rect 9602 2054 9612 2106
rect 9664 2054 9674 2106
rect 9602 2050 9674 2054
rect 11320 2106 11392 2110
rect 11320 2054 11330 2106
rect 11382 2054 11392 2106
rect 11320 2050 11392 2054
rect 11748 2106 11820 2110
rect 11748 2054 11758 2106
rect 11810 2054 11820 2106
rect 11748 2050 11820 2054
rect 12180 2108 12252 2110
rect 12516 2109 12555 2143
rect 12589 2109 12628 2143
rect 12516 2108 12628 2109
rect 12180 2106 12628 2108
rect 12180 2054 12190 2106
rect 12242 2071 12628 2106
rect 12242 2054 12555 2071
rect 12180 2050 12555 2054
rect -295 2048 232 2050
rect -295 2037 -256 2048
rect -368 1999 -256 2037
rect -368 1965 -329 1999
rect -295 1965 -256 1999
rect -368 1927 -256 1965
rect -368 1893 -329 1927
rect -295 1893 -256 1927
rect -368 1855 -256 1893
rect -368 1821 -329 1855
rect -295 1821 -256 1855
rect -368 1783 -256 1821
rect -98 1842 -26 1846
rect -98 1790 -88 1842
rect -36 1790 -26 1842
rect -98 1786 -26 1790
rect -368 1749 -329 1783
rect -295 1749 -256 1783
rect -368 1711 -256 1749
rect -368 1677 -329 1711
rect -295 1677 -256 1711
rect -368 1639 -256 1677
rect -368 1605 -329 1639
rect -295 1605 -256 1639
rect -368 1567 -256 1605
rect -368 1533 -329 1567
rect -295 1533 -256 1567
rect -368 1495 -256 1533
rect -368 1461 -329 1495
rect -295 1461 -256 1495
rect -368 1423 -256 1461
rect -368 1389 -329 1423
rect -295 1389 -256 1423
rect -368 1351 -256 1389
rect -368 1317 -329 1351
rect -295 1317 -256 1351
rect -368 1279 -256 1317
rect -368 1245 -329 1279
rect -295 1245 -256 1279
rect -368 1207 -256 1245
rect -368 1173 -329 1207
rect -295 1173 -256 1207
rect -368 1135 -256 1173
rect -368 1101 -329 1135
rect -295 1101 -256 1135
rect -368 1063 -256 1101
rect -368 1029 -329 1063
rect -295 1029 -256 1063
rect -368 991 -256 1029
rect -368 957 -329 991
rect -295 957 -256 991
rect -368 919 -256 957
rect -368 885 -329 919
rect -295 885 -256 919
rect -368 847 -256 885
rect -368 813 -329 847
rect -295 813 -256 847
rect -368 775 -256 813
rect -368 741 -329 775
rect -295 741 -256 775
rect -368 703 -256 741
rect -368 669 -329 703
rect -295 669 -256 703
rect -368 631 -256 669
rect -368 597 -329 631
rect -295 597 -256 631
rect -368 559 -256 597
rect -368 525 -329 559
rect -295 525 -256 559
rect -368 487 -256 525
rect -368 453 -329 487
rect -295 453 -256 487
rect -368 415 -256 453
rect -368 381 -329 415
rect -295 381 -256 415
rect -368 343 -256 381
rect -368 309 -329 343
rect -295 309 -256 343
rect -368 271 -256 309
rect -368 237 -329 271
rect -295 237 -256 271
rect -368 199 -256 237
rect -368 165 -329 199
rect -295 165 -256 199
rect -368 127 -256 165
rect -368 93 -329 127
rect -295 93 -256 127
rect -368 55 -256 93
rect -368 21 -329 55
rect -295 21 -256 55
rect -368 -17 -256 21
rect -368 -51 -329 -17
rect -295 -51 -256 -17
rect -92 -50 -32 1786
rect 44 1714 116 1718
rect 44 1662 54 1714
rect 106 1662 116 1714
rect 44 1658 116 1662
rect 50 56 110 1658
rect 172 1414 232 2048
rect 596 1550 656 2050
rect 1032 1414 1092 2050
rect 1452 1978 1524 1982
rect 1452 1926 1462 1978
rect 1514 1926 1524 1978
rect 1452 1922 1524 1926
rect 2306 1978 2378 1982
rect 2306 1926 2316 1978
rect 2368 1926 2378 1978
rect 2306 1922 2378 1926
rect 1458 1550 1518 1922
rect 2312 1556 2372 1922
rect 2746 1422 2806 2050
rect 3166 1978 3238 1982
rect 3166 1926 3176 1978
rect 3228 1926 3238 1978
rect 3166 1922 3238 1926
rect 4026 1978 4098 1982
rect 4026 1926 4036 1978
rect 4088 1926 4098 1978
rect 4026 1922 4098 1926
rect 3172 1556 3232 1922
rect 4032 1556 4092 1922
rect 4466 1436 4526 2050
rect 4886 1978 4958 1982
rect 4886 1926 4896 1978
rect 4948 1926 4958 1978
rect 4886 1922 4958 1926
rect 5746 1978 5818 1982
rect 5746 1926 5756 1978
rect 5808 1926 5818 1978
rect 5746 1922 5818 1926
rect 4892 1556 4952 1922
rect 5752 1556 5812 1922
rect 6174 1436 6234 2050
rect 6606 1978 6678 1982
rect 6606 1926 6616 1978
rect 6668 1926 6678 1978
rect 6606 1922 6678 1926
rect 7466 1978 7538 1982
rect 7466 1926 7476 1978
rect 7528 1926 7538 1978
rect 7466 1922 7538 1926
rect 6612 1556 6672 1922
rect 7472 1556 7532 1922
rect 7894 1416 7954 2050
rect 8326 1978 8398 1982
rect 8326 1926 8336 1978
rect 8388 1926 8398 1978
rect 8326 1922 8398 1926
rect 9166 1978 9238 1982
rect 9166 1926 9176 1978
rect 9228 1926 9238 1978
rect 9166 1922 9238 1926
rect 8332 1556 8392 1922
rect 8746 1714 8818 1718
rect 8746 1662 8756 1714
rect 8808 1662 8818 1714
rect 8746 1658 8818 1662
rect 8752 1342 8812 1658
rect 9172 1556 9232 1922
rect 9608 1414 9668 2050
rect 10024 1978 10096 1982
rect 10024 1926 10034 1978
rect 10086 1926 10096 1978
rect 10024 1922 10096 1926
rect 10886 1978 10958 1982
rect 10886 1926 10896 1978
rect 10948 1926 10958 1978
rect 10886 1922 10958 1926
rect 10030 1548 10090 1922
rect 10462 1842 10534 1846
rect 10462 1790 10472 1842
rect 10524 1790 10534 1842
rect 10462 1786 10534 1790
rect 10468 1356 10528 1786
rect 10892 1548 10952 1922
rect 11326 1432 11386 2050
rect 11754 1544 11814 2050
rect 12186 2048 12555 2050
rect 12186 1418 12246 2048
rect 12516 2037 12555 2048
rect 12589 2037 12628 2071
rect 12516 1999 12628 2037
rect 12516 1965 12555 1999
rect 12589 1965 12628 1999
rect 12516 1927 12628 1965
rect 12516 1893 12555 1927
rect 12589 1893 12628 1927
rect 12516 1855 12628 1893
rect 12516 1821 12555 1855
rect 12589 1821 12628 1855
rect 12516 1783 12628 1821
rect 12516 1749 12555 1783
rect 12589 1749 12628 1783
rect 12516 1711 12628 1749
rect 12516 1677 12555 1711
rect 12589 1677 12628 1711
rect 12516 1639 12628 1677
rect 12516 1605 12555 1639
rect 12589 1605 12628 1639
rect 12516 1567 12628 1605
rect 12516 1533 12555 1567
rect 12589 1533 12628 1567
rect 12516 1495 12628 1533
rect 12516 1461 12555 1495
rect 12589 1461 12628 1495
rect 12516 1423 12628 1461
rect 12516 1389 12555 1423
rect 12589 1389 12628 1423
rect 12516 1351 12628 1389
rect 12516 1317 12555 1351
rect 12589 1317 12628 1351
rect 12516 1279 12628 1317
rect 12516 1245 12555 1279
rect 12589 1245 12628 1279
rect 12516 1207 12628 1245
rect 12516 1173 12555 1207
rect 12589 1173 12628 1207
rect 12516 1135 12628 1173
rect 12516 1101 12555 1135
rect 12589 1101 12628 1135
rect 12516 1063 12628 1101
rect 12516 1029 12555 1063
rect 12589 1029 12628 1063
rect 12516 991 12628 1029
rect 12516 957 12555 991
rect 12589 957 12628 991
rect 12516 919 12628 957
rect 12516 885 12555 919
rect 12589 885 12628 919
rect 12516 847 12628 885
rect 12516 813 12555 847
rect 12589 813 12628 847
rect 12516 775 12628 813
rect 12516 741 12555 775
rect 12589 741 12628 775
rect 12516 703 12628 741
rect 12516 669 12555 703
rect 12589 669 12628 703
rect 12516 631 12628 669
rect 12516 597 12555 631
rect 12589 597 12628 631
rect 12516 559 12628 597
rect 12516 525 12555 559
rect 12589 525 12628 559
rect 12516 487 12628 525
rect 170 62 230 394
rect 600 62 660 252
rect 1030 62 1090 396
rect 44 52 116 56
rect 44 0 54 52
rect 106 0 116 52
rect 44 -4 116 0
rect 170 -6 1090 62
rect -368 -89 -256 -51
rect -368 -123 -329 -89
rect -295 -123 -256 -89
rect -98 -54 -26 -50
rect -98 -106 -88 -54
rect -36 -106 -26 -54
rect -98 -110 -26 -106
rect -368 -161 -256 -123
rect -368 -195 -329 -161
rect -295 -195 -256 -161
rect -368 -233 -256 -195
rect -368 -267 -329 -233
rect -295 -267 -256 -233
rect -368 -305 -256 -267
rect -368 -339 -329 -305
rect -295 -339 -256 -305
rect -368 -377 -256 -339
rect -368 -411 -329 -377
rect -295 -411 -256 -377
rect -368 -449 -256 -411
rect -368 -483 -329 -449
rect -295 -483 -256 -449
rect -368 -521 -256 -483
rect -368 -555 -329 -521
rect -295 -555 -256 -521
rect -368 -593 -256 -555
rect -368 -627 -329 -593
rect -295 -627 -256 -593
rect -368 -665 -256 -627
rect -368 -699 -329 -665
rect -295 -699 -256 -665
rect -368 -737 -256 -699
rect -368 -771 -329 -737
rect -295 -771 -256 -737
rect -368 -809 -256 -771
rect -368 -843 -329 -809
rect -295 -843 -256 -809
rect -368 -881 -256 -843
rect -368 -915 -329 -881
rect -295 -915 -256 -881
rect -368 -953 -256 -915
rect -368 -987 -329 -953
rect -295 -987 -256 -953
rect -368 -1025 -256 -987
rect -368 -1059 -329 -1025
rect -295 -1059 -256 -1025
rect -368 -1097 -256 -1059
rect -368 -1131 -329 -1097
rect -295 -1131 -256 -1097
rect -368 -1169 -256 -1131
rect -368 -1203 -329 -1169
rect -295 -1203 -256 -1169
rect -368 -1241 -256 -1203
rect -368 -1275 -329 -1241
rect -295 -1275 -256 -1241
rect -368 -1313 -256 -1275
rect -368 -1347 -329 -1313
rect -295 -1347 -256 -1313
rect -368 -1385 -256 -1347
rect -368 -1419 -329 -1385
rect -295 -1419 -256 -1385
rect -368 -1457 -256 -1419
rect -368 -1491 -329 -1457
rect -295 -1491 -256 -1457
rect -368 -1529 -256 -1491
rect -368 -1563 -329 -1529
rect -295 -1563 -256 -1529
rect -368 -1601 -256 -1563
rect -368 -1635 -329 -1601
rect -295 -1635 -256 -1601
rect -368 -1673 -256 -1635
rect -98 -1584 -26 -1580
rect -98 -1636 -88 -1584
rect -36 -1636 -26 -1584
rect -98 -1640 -26 -1636
rect -368 -1707 -329 -1673
rect -295 -1707 -256 -1673
rect -368 -1745 -256 -1707
rect -368 -1779 -329 -1745
rect -295 -1779 -256 -1745
rect -368 -1817 -256 -1779
rect -368 -1851 -329 -1817
rect -295 -1851 -256 -1817
rect -368 -1889 -256 -1851
rect -368 -1923 -329 -1889
rect -295 -1923 -256 -1889
rect -368 -1961 -256 -1923
rect -368 -1995 -329 -1961
rect -295 -1995 -256 -1961
rect -368 -2033 -256 -1995
rect -368 -2067 -329 -2033
rect -295 -2067 -256 -2033
rect -368 -2105 -256 -2067
rect -368 -2139 -329 -2105
rect -295 -2139 -256 -2105
rect -368 -2177 -256 -2139
rect -368 -2211 -329 -2177
rect -295 -2211 -256 -2177
rect -368 -2249 -256 -2211
rect -368 -2283 -329 -2249
rect -295 -2283 -256 -2249
rect -368 -2321 -256 -2283
rect -368 -2355 -329 -2321
rect -295 -2355 -256 -2321
rect -368 -2393 -256 -2355
rect -368 -2427 -329 -2393
rect -295 -2427 -256 -2393
rect -368 -2465 -256 -2427
rect -368 -2499 -329 -2465
rect -295 -2499 -256 -2465
rect -368 -2537 -256 -2499
rect -368 -2571 -329 -2537
rect -295 -2571 -256 -2537
rect -368 -2609 -256 -2571
rect -368 -2643 -329 -2609
rect -295 -2643 -256 -2609
rect -368 -2681 -256 -2643
rect -368 -2715 -329 -2681
rect -295 -2715 -256 -2681
rect -368 -2753 -256 -2715
rect -368 -2787 -329 -2753
rect -295 -2787 -256 -2753
rect -368 -2825 -256 -2787
rect -368 -2859 -329 -2825
rect -295 -2859 -256 -2825
rect -368 -2897 -256 -2859
rect -368 -2931 -329 -2897
rect -295 -2931 -256 -2897
rect -368 -2969 -256 -2931
rect -368 -3003 -329 -2969
rect -295 -3003 -256 -2969
rect -368 -3041 -256 -3003
rect -368 -3075 -329 -3041
rect -295 -3075 -256 -3041
rect -368 -3113 -256 -3075
rect -368 -3147 -329 -3113
rect -295 -3147 -256 -3113
rect -368 -3185 -256 -3147
rect -368 -3219 -329 -3185
rect -295 -3219 -256 -3185
rect -368 -3257 -256 -3219
rect -368 -3291 -329 -3257
rect -295 -3291 -256 -3257
rect -368 -3329 -256 -3291
rect -368 -3363 -329 -3329
rect -295 -3363 -256 -3329
rect -368 -3401 -256 -3363
rect -368 -3435 -329 -3401
rect -295 -3435 -256 -3401
rect -368 -3473 -256 -3435
rect -368 -3507 -329 -3473
rect -295 -3507 -256 -3473
rect -368 -3545 -256 -3507
rect -92 -3530 -32 -1640
rect 170 -1682 230 -6
rect 600 -195 660 -6
rect 600 -1682 660 -1482
rect 1030 -1682 1090 -6
rect 1460 -195 1520 252
rect 1888 156 1948 454
rect 12516 453 12555 487
rect 12589 453 12628 487
rect 1882 152 1954 156
rect 1882 100 1892 152
rect 1944 100 1954 152
rect 1882 96 1954 100
rect 1884 -54 1956 -50
rect 1884 -106 1894 -54
rect 1946 -106 1956 -54
rect 1884 -110 1956 -106
rect 1890 -298 1950 -110
rect 2320 -195 2380 252
rect 1460 -1678 1520 -1482
rect 170 -1742 1090 -1682
rect 44 -1790 116 -1786
rect 44 -1842 54 -1790
rect 106 -1842 116 -1790
rect 44 -1846 116 -1842
rect 50 -3424 110 -1846
rect 170 -3424 230 -1742
rect 600 -1929 660 -1742
rect 600 -3424 660 -3222
rect 1030 -3424 1090 -1742
rect 1458 -1688 1520 -1678
rect 1458 -1740 1462 -1688
rect 1514 -1740 1520 -1688
rect 1458 -1750 1520 -1740
rect 1460 -1929 1520 -1750
rect 2320 -1688 2380 -1482
rect 2320 -1740 2324 -1688
rect 2376 -1740 2380 -1688
rect 2320 -1929 2380 -1740
rect 44 -3428 116 -3424
rect 44 -3480 54 -3428
rect 106 -3480 116 -3428
rect 44 -3484 116 -3480
rect 170 -3484 1090 -3424
rect -368 -3579 -329 -3545
rect -295 -3579 -256 -3545
rect -368 -3617 -256 -3579
rect -98 -3534 -26 -3530
rect -98 -3586 -88 -3534
rect -36 -3586 -26 -3534
rect -98 -3590 -26 -3586
rect -368 -3651 -329 -3617
rect -295 -3651 -256 -3617
rect -368 -3689 -256 -3651
rect -368 -3723 -329 -3689
rect -295 -3723 -256 -3689
rect -368 -3761 -256 -3723
rect -368 -3795 -329 -3761
rect -295 -3795 -256 -3761
rect -368 -3833 -256 -3795
rect -368 -3867 -329 -3833
rect -295 -3867 -256 -3833
rect -368 -3905 -256 -3867
rect -368 -3939 -329 -3905
rect -295 -3939 -256 -3905
rect -368 -3977 -256 -3939
rect -368 -4011 -329 -3977
rect -295 -4011 -256 -3977
rect -368 -4049 -256 -4011
rect -368 -4083 -329 -4049
rect -295 -4083 -256 -4049
rect -368 -4121 -256 -4083
rect -368 -4155 -329 -4121
rect -295 -4155 -256 -4121
rect -368 -4193 -256 -4155
rect -368 -4227 -329 -4193
rect -295 -4227 -256 -4193
rect -368 -4265 -256 -4227
rect -368 -4299 -329 -4265
rect -295 -4299 -256 -4265
rect -368 -4337 -256 -4299
rect -368 -4371 -329 -4337
rect -295 -4371 -256 -4337
rect -368 -4409 -256 -4371
rect -368 -4443 -329 -4409
rect -295 -4443 -256 -4409
rect -368 -4481 -256 -4443
rect -368 -4515 -329 -4481
rect -295 -4515 -256 -4481
rect -368 -4553 -256 -4515
rect -368 -4587 -329 -4553
rect -295 -4587 -256 -4553
rect -368 -4625 -256 -4587
rect -368 -4659 -329 -4625
rect -295 -4659 -256 -4625
rect -368 -4697 -256 -4659
rect -368 -4731 -329 -4697
rect -295 -4731 -256 -4697
rect -368 -4769 -256 -4731
rect -368 -4803 -329 -4769
rect -295 -4803 -256 -4769
rect -368 -4841 -256 -4803
rect -368 -4875 -329 -4841
rect -295 -4875 -256 -4841
rect -368 -4913 -256 -4875
rect -368 -4947 -329 -4913
rect -295 -4947 -256 -4913
rect -368 -4985 -256 -4947
rect -368 -5019 -329 -4985
rect -295 -5019 -256 -4985
rect -368 -5057 -256 -5019
rect -368 -5091 -329 -5057
rect -295 -5091 -256 -5057
rect -368 -5129 -256 -5091
rect -368 -5163 -329 -5129
rect -295 -5150 -256 -5129
rect 170 -5150 230 -3484
rect 600 -3669 660 -3484
rect 600 -5150 660 -4964
rect 1030 -5150 1090 -3484
rect 1460 -3669 1520 -3222
rect 1888 -3324 1948 -3026
rect 1882 -3328 1954 -3324
rect 1882 -3380 1892 -3328
rect 1944 -3380 1954 -3328
rect 1882 -3384 1954 -3380
rect 1884 -3534 1956 -3530
rect 1884 -3586 1894 -3534
rect 1946 -3586 1956 -3534
rect 1884 -3590 1956 -3586
rect 1890 -3778 1950 -3590
rect 2320 -3669 2380 -3222
rect 1460 -5050 1520 -4964
rect 1454 -5054 1526 -5050
rect 1454 -5106 1464 -5054
rect 1516 -5106 1526 -5054
rect 1454 -5110 1526 -5106
rect 2320 -5054 2380 -4964
rect 2320 -5106 2324 -5054
rect 2376 -5106 2380 -5054
rect -295 -5163 1090 -5150
rect -368 -5201 1090 -5163
rect -368 -5235 -329 -5201
rect -295 -5210 1090 -5201
rect -295 -5235 -256 -5210
rect -368 -5273 -256 -5235
rect -368 -5307 -329 -5273
rect -295 -5307 -256 -5273
rect -368 -5345 -256 -5307
rect -368 -5379 -329 -5345
rect -295 -5379 -256 -5345
rect -368 -5417 -256 -5379
rect -368 -5451 -329 -5417
rect -295 -5451 -256 -5417
rect -368 -5489 -256 -5451
rect -368 -5523 -329 -5489
rect -295 -5523 -256 -5489
rect -368 -5561 -256 -5523
rect -368 -5595 -329 -5561
rect -295 -5595 -256 -5561
rect -368 -5633 -256 -5595
rect -368 -5667 -329 -5633
rect -295 -5667 -256 -5633
rect -368 -5705 -256 -5667
rect -368 -5739 -329 -5705
rect -295 -5739 -256 -5705
rect -368 -5777 -256 -5739
rect -368 -5811 -329 -5777
rect -295 -5811 -256 -5777
rect -368 -5849 -256 -5811
rect -368 -5883 -329 -5849
rect -295 -5883 -256 -5849
rect -368 -5921 -256 -5883
rect -368 -5955 -329 -5921
rect -295 -5955 -256 -5921
rect -368 -5993 -256 -5955
rect -368 -6027 -329 -5993
rect -295 -6027 -256 -5993
rect -368 -6065 -256 -6027
rect -368 -6099 -329 -6065
rect -295 -6099 -256 -6065
rect -368 -6137 -256 -6099
rect -368 -6171 -329 -6137
rect -295 -6171 -256 -6137
rect -368 -6209 -256 -6171
rect -368 -6243 -329 -6209
rect -295 -6243 -256 -6209
rect -368 -6281 -256 -6243
rect -368 -6315 -329 -6281
rect -295 -6315 -256 -6281
rect -368 -6353 -256 -6315
rect -368 -6387 -329 -6353
rect -295 -6387 -256 -6353
rect -368 -6425 -256 -6387
rect -368 -6459 -329 -6425
rect -295 -6459 -256 -6425
rect -368 -6497 -256 -6459
rect -368 -6531 -329 -6497
rect -295 -6531 -256 -6497
rect -368 -6569 -256 -6531
rect -368 -6603 -329 -6569
rect -295 -6603 -256 -6569
rect -368 -6641 -256 -6603
rect -368 -6675 -329 -6641
rect -295 -6675 -256 -6641
rect -368 -6713 -256 -6675
rect -368 -6747 -329 -6713
rect -295 -6747 -256 -6713
rect -368 -6785 -256 -6747
rect -368 -6819 -329 -6785
rect -295 -6819 -256 -6785
rect -368 -6857 -256 -6819
rect -368 -6891 -329 -6857
rect -295 -6891 -256 -6857
rect -368 -6929 -256 -6891
rect -368 -6963 -329 -6929
rect -295 -6963 -256 -6929
rect -368 -7001 -256 -6963
rect -368 -7035 -329 -7001
rect -295 -7035 -256 -7001
rect -368 -7073 -256 -7035
rect 170 -7070 230 -5210
rect 600 -5411 660 -5210
rect 1030 -5542 1090 -5210
rect 1460 -5411 1520 -5110
rect 1882 -5272 1954 -5268
rect 1882 -5324 1892 -5272
rect 1944 -5324 1954 -5272
rect 1882 -5328 1954 -5324
rect 1888 -5580 1948 -5328
rect 2320 -5411 2380 -5106
rect 590 -7070 650 -6700
rect 1030 -7070 1090 -6548
rect 1456 -6926 1516 -6700
rect 2326 -6926 2386 -6697
rect 1450 -6930 1522 -6926
rect 1450 -6982 1460 -6930
rect 1512 -6982 1522 -6930
rect 1450 -6986 1522 -6982
rect 2320 -6930 2392 -6926
rect 2320 -6982 2330 -6930
rect 2382 -6982 2392 -6930
rect 2320 -6986 2392 -6982
rect 2748 -7070 2808 388
rect 3180 -195 3240 252
rect 3464 52 3536 56
rect 3604 54 3664 360
rect 3464 0 3474 52
rect 3526 0 3536 52
rect 3464 -4 3536 0
rect 3598 50 3670 54
rect 3598 -2 3608 50
rect 3660 -2 3670 50
rect 3470 -48 3530 -4
rect 3598 -6 3670 -2
rect 3470 -108 3664 -48
rect 3604 -312 3664 -108
rect 4040 -195 4100 252
rect 3180 -1678 3240 -1482
rect 3180 -1688 3242 -1678
rect 3180 -1740 3186 -1688
rect 3238 -1740 3242 -1688
rect 3180 -1750 3242 -1740
rect 4040 -1688 4100 -1482
rect 4040 -1740 4044 -1688
rect 4096 -1740 4100 -1688
rect 3180 -1929 3240 -1750
rect 4040 -1929 4100 -1740
rect 3180 -3669 3240 -3222
rect 3464 -3428 3536 -3424
rect 3604 -3426 3664 -3120
rect 3464 -3480 3474 -3428
rect 3526 -3480 3536 -3428
rect 3464 -3484 3536 -3480
rect 3598 -3430 3670 -3426
rect 3598 -3482 3608 -3430
rect 3660 -3482 3670 -3430
rect 3470 -3528 3530 -3484
rect 3598 -3486 3670 -3482
rect 3470 -3588 3664 -3528
rect 3604 -3792 3664 -3588
rect 4040 -3669 4100 -3222
rect 4462 -3536 4522 386
rect 4900 -195 4960 252
rect 5318 54 5378 420
rect 12516 415 12628 453
rect 7038 156 7098 368
rect 7038 96 7226 156
rect 5318 -6 7096 54
rect 5314 -54 5386 -50
rect 5314 -106 5324 -54
rect 5376 -106 5386 -54
rect 5314 -110 5386 -106
rect 5320 -406 5380 -110
rect 7036 -112 7096 -6
rect 7166 -50 7226 96
rect 7160 -54 7232 -50
rect 7160 -106 7170 -54
rect 7222 -106 7232 -54
rect 7160 -110 7232 -106
rect 7036 -280 7098 -112
rect 7480 -195 7540 252
rect 7038 -294 7098 -280
rect 4900 -1688 4960 -1482
rect 4900 -1740 4904 -1688
rect 4956 -1740 4960 -1688
rect 4900 -1929 4960 -1740
rect 5744 -1688 5804 -1485
rect 5744 -1740 5748 -1688
rect 5800 -1740 5804 -1688
rect 5744 -1936 5804 -1740
rect 4462 -3588 4466 -3536
rect 4518 -3588 4522 -3536
rect 3180 -5044 3240 -4964
rect 3176 -5054 3240 -5044
rect 3176 -5106 3180 -5054
rect 3232 -5106 3240 -5054
rect 3176 -5116 3240 -5106
rect 3180 -5411 3240 -5116
rect 4040 -5044 4100 -4964
rect 4040 -5054 4102 -5044
rect 4040 -5106 4046 -5054
rect 4098 -5106 4102 -5054
rect 4040 -5116 4102 -5106
rect 3600 -5158 3672 -5154
rect 3600 -5210 3610 -5158
rect 3662 -5210 3672 -5158
rect 3600 -5214 3672 -5210
rect 3606 -5520 3666 -5214
rect 4040 -5411 4100 -5116
rect 3184 -6926 3244 -6697
rect 4042 -6926 4102 -6697
rect 3178 -6930 3250 -6926
rect 3178 -6982 3188 -6930
rect 3240 -6982 3250 -6930
rect 3178 -6986 3250 -6982
rect 4036 -6930 4108 -6926
rect 4036 -6982 4046 -6930
rect 4098 -6982 4108 -6930
rect 4036 -6986 4108 -6982
rect 4462 -7070 4522 -3588
rect 4900 -3669 4960 -3222
rect 5318 -3426 5378 -3060
rect 6180 -3200 6240 -332
rect 6614 -1688 6674 -1481
rect 6614 -1740 6618 -1688
rect 6670 -1740 6674 -1688
rect 6614 -1932 6674 -1740
rect 7480 -1688 7540 -1482
rect 7480 -1740 7484 -1688
rect 7536 -1740 7540 -1688
rect 7480 -1929 7540 -1740
rect 6180 -3252 6184 -3200
rect 6236 -3252 6240 -3200
rect 6180 -3262 6240 -3252
rect 7038 -3324 7098 -3112
rect 7038 -3384 7226 -3324
rect 5318 -3486 7096 -3426
rect 5314 -3534 5386 -3530
rect 5314 -3586 5324 -3534
rect 5376 -3586 5386 -3534
rect 5314 -3590 5386 -3586
rect 5320 -3886 5380 -3590
rect 7036 -3592 7096 -3486
rect 7166 -3530 7226 -3384
rect 7160 -3534 7232 -3530
rect 7160 -3586 7170 -3534
rect 7222 -3586 7232 -3534
rect 7160 -3590 7232 -3586
rect 7036 -3760 7098 -3592
rect 7480 -3669 7540 -3222
rect 7894 -3534 7954 384
rect 8336 -195 8396 252
rect 8750 50 8822 54
rect 8750 -2 8760 50
rect 8812 -2 8822 50
rect 8750 -6 8822 -2
rect 8756 -340 8816 -6
rect 9192 -195 9252 252
rect 8336 -1688 8396 -1482
rect 8336 -1740 8340 -1688
rect 8392 -1740 8396 -1688
rect 8336 -1929 8396 -1740
rect 9192 -1688 9252 -1482
rect 9192 -1740 9196 -1688
rect 9248 -1740 9252 -1688
rect 8746 -1790 8818 -1786
rect 8746 -1842 8756 -1790
rect 8808 -1842 8818 -1790
rect 8746 -1846 8818 -1842
rect 8752 -2138 8812 -1846
rect 9192 -1929 9252 -1740
rect 7894 -3586 7898 -3534
rect 7950 -3586 7954 -3534
rect 7038 -3774 7098 -3760
rect 4900 -5044 4960 -4964
rect 4898 -5054 4960 -5044
rect 4898 -5106 4902 -5054
rect 4954 -5106 4960 -5054
rect 4898 -5116 4960 -5106
rect 4900 -5411 4960 -5116
rect 5742 -5044 5802 -4967
rect 5742 -5054 5806 -5044
rect 5742 -5106 5750 -5054
rect 5802 -5106 5806 -5054
rect 5742 -5116 5806 -5106
rect 5742 -5418 5802 -5116
rect 4900 -6926 4960 -6697
rect 5320 -6800 5380 -6540
rect 5314 -6804 5386 -6800
rect 5314 -6856 5324 -6804
rect 5376 -6856 5386 -6804
rect 5314 -6860 5386 -6856
rect 5758 -6926 5818 -6697
rect 4894 -6930 4966 -6926
rect 4894 -6982 4904 -6930
rect 4956 -6982 4966 -6930
rect 4894 -6986 4966 -6982
rect 5752 -6930 5824 -6926
rect 5752 -6982 5762 -6930
rect 5814 -6982 5824 -6930
rect 5752 -6986 5824 -6982
rect 6180 -7070 6240 -3788
rect 6602 -5044 6662 -4959
rect 6600 -5054 6662 -5044
rect 6600 -5106 6604 -5054
rect 6656 -5106 6662 -5054
rect 6600 -5116 6662 -5106
rect 6602 -5410 6662 -5116
rect 7480 -5054 7540 -4964
rect 7480 -5106 7484 -5054
rect 7536 -5106 7540 -5054
rect 7480 -5411 7540 -5106
rect 6616 -6926 6676 -6697
rect 7038 -6800 7098 -6602
rect 7032 -6804 7104 -6800
rect 7032 -6856 7042 -6804
rect 7094 -6856 7104 -6804
rect 7032 -6860 7104 -6856
rect 7474 -6926 7534 -6697
rect 6610 -6930 6682 -6926
rect 6610 -6982 6620 -6930
rect 6672 -6982 6682 -6930
rect 6610 -6986 6682 -6982
rect 7468 -6930 7540 -6926
rect 7468 -6982 7478 -6930
rect 7530 -6982 7540 -6930
rect 7468 -6986 7540 -6982
rect 7894 -7070 7954 -3586
rect 8336 -3669 8396 -3222
rect 8750 -3430 8822 -3426
rect 8750 -3482 8760 -3430
rect 8812 -3482 8822 -3430
rect 8750 -3486 8822 -3482
rect 8756 -3820 8816 -3486
rect 9192 -3669 9252 -3222
rect 8336 -5044 8396 -4964
rect 8334 -5054 8396 -5044
rect 8334 -5106 8338 -5054
rect 8390 -5106 8396 -5054
rect 8334 -5116 8396 -5106
rect 8336 -5411 8396 -5116
rect 9192 -5058 9252 -4964
rect 9192 -5110 9196 -5058
rect 9248 -5110 9252 -5058
rect 8746 -5158 8818 -5154
rect 8746 -5210 8756 -5158
rect 8808 -5210 8818 -5158
rect 8746 -5214 8818 -5210
rect 8752 -5518 8812 -5214
rect 9192 -5411 9252 -5110
rect 8332 -6926 8392 -6697
rect 9190 -6926 9250 -6697
rect 8326 -6930 8398 -6926
rect 8326 -6982 8336 -6930
rect 8388 -6982 8398 -6930
rect 8326 -6986 8398 -6982
rect 9184 -6930 9256 -6926
rect 9184 -6982 9194 -6930
rect 9246 -6982 9256 -6930
rect 9184 -6986 9256 -6982
rect 9608 -7070 9668 390
rect 10048 -195 10108 252
rect 10464 152 10536 156
rect 10464 100 10474 152
rect 10526 100 10536 152
rect 10464 96 10536 100
rect 10470 -304 10530 96
rect 10904 -190 10964 252
rect 11326 66 11386 406
rect 11750 66 11810 255
rect 12184 66 12244 394
rect 12516 381 12555 415
rect 12589 381 12628 415
rect 12516 343 12628 381
rect 12516 309 12555 343
rect 12589 309 12628 343
rect 12516 271 12628 309
rect 12516 237 12555 271
rect 12589 237 12628 271
rect 12516 199 12628 237
rect 12516 165 12555 199
rect 12589 165 12628 199
rect 12516 127 12628 165
rect 12516 93 12555 127
rect 12589 93 12628 127
rect 12516 66 12628 93
rect 11326 55 12628 66
rect 11326 21 12555 55
rect 12589 21 12628 55
rect 11326 6 12628 21
rect 10048 -1678 10108 -1482
rect 10462 -1584 10534 -1580
rect 10462 -1636 10472 -1584
rect 10524 -1636 10534 -1584
rect 10462 -1640 10534 -1636
rect 10046 -1688 10108 -1678
rect 10046 -1740 10050 -1688
rect 10102 -1740 10108 -1688
rect 10046 -1750 10108 -1740
rect 10048 -1929 10108 -1750
rect 10468 -2124 10528 -1640
rect 10904 -1684 10964 -1482
rect 11326 -1680 11386 6
rect 11750 -196 11810 6
rect 11754 -1680 11814 -1481
rect 12184 -1680 12244 6
rect 12516 -17 12628 6
rect 12516 -51 12555 -17
rect 12589 -51 12628 -17
rect 12516 -89 12628 -51
rect 12516 -123 12555 -89
rect 12589 -123 12628 -89
rect 12516 -161 12628 -123
rect 12516 -195 12555 -161
rect 12589 -195 12628 -161
rect 12516 -233 12628 -195
rect 12516 -267 12555 -233
rect 12589 -267 12628 -233
rect 12516 -305 12628 -267
rect 12516 -339 12555 -305
rect 12589 -339 12628 -305
rect 12516 -377 12628 -339
rect 12516 -411 12555 -377
rect 12589 -411 12628 -377
rect 12516 -449 12628 -411
rect 12516 -483 12555 -449
rect 12589 -483 12628 -449
rect 12516 -521 12628 -483
rect 12516 -555 12555 -521
rect 12589 -555 12628 -521
rect 12516 -593 12628 -555
rect 12516 -627 12555 -593
rect 12589 -627 12628 -593
rect 12516 -665 12628 -627
rect 12516 -699 12555 -665
rect 12589 -699 12628 -665
rect 12516 -737 12628 -699
rect 12516 -771 12555 -737
rect 12589 -771 12628 -737
rect 12516 -809 12628 -771
rect 12516 -843 12555 -809
rect 12589 -843 12628 -809
rect 12516 -881 12628 -843
rect 12516 -915 12555 -881
rect 12589 -915 12628 -881
rect 12516 -953 12628 -915
rect 12516 -987 12555 -953
rect 12589 -987 12628 -953
rect 12516 -1025 12628 -987
rect 12516 -1059 12555 -1025
rect 12589 -1059 12628 -1025
rect 12516 -1097 12628 -1059
rect 12516 -1131 12555 -1097
rect 12589 -1131 12628 -1097
rect 12516 -1169 12628 -1131
rect 12516 -1203 12555 -1169
rect 12589 -1203 12628 -1169
rect 12516 -1241 12628 -1203
rect 12516 -1275 12555 -1241
rect 12589 -1275 12628 -1241
rect 12516 -1313 12628 -1275
rect 12516 -1347 12555 -1313
rect 12589 -1347 12628 -1313
rect 12516 -1385 12628 -1347
rect 12516 -1419 12555 -1385
rect 12589 -1419 12628 -1385
rect 12516 -1457 12628 -1419
rect 12516 -1491 12555 -1457
rect 12589 -1491 12628 -1457
rect 12516 -1529 12628 -1491
rect 12516 -1563 12555 -1529
rect 12589 -1563 12628 -1529
rect 12516 -1601 12628 -1563
rect 12516 -1635 12555 -1601
rect 12589 -1635 12628 -1601
rect 12516 -1673 12628 -1635
rect 12516 -1680 12555 -1673
rect 10898 -1688 10970 -1684
rect 10898 -1740 10908 -1688
rect 10960 -1740 10970 -1688
rect 10898 -1744 10970 -1740
rect 11326 -1707 12555 -1680
rect 12589 -1707 12628 -1673
rect 11326 -1740 12628 -1707
rect 10904 -1929 10964 -1744
rect 10048 -3669 10108 -3222
rect 10464 -3328 10536 -3324
rect 10464 -3380 10474 -3328
rect 10526 -3380 10536 -3328
rect 10464 -3384 10536 -3380
rect 10470 -3784 10530 -3384
rect 10904 -3669 10964 -3222
rect 11326 -3412 11386 -1740
rect 11754 -1932 11814 -1740
rect 11750 -3412 11810 -3223
rect 12184 -3412 12244 -1740
rect 12516 -1745 12628 -1740
rect 12516 -1779 12555 -1745
rect 12589 -1779 12628 -1745
rect 12516 -1817 12628 -1779
rect 12516 -1851 12555 -1817
rect 12589 -1851 12628 -1817
rect 12516 -1889 12628 -1851
rect 12516 -1923 12555 -1889
rect 12589 -1923 12628 -1889
rect 12516 -1961 12628 -1923
rect 12516 -1995 12555 -1961
rect 12589 -1995 12628 -1961
rect 12516 -2033 12628 -1995
rect 12516 -2067 12555 -2033
rect 12589 -2067 12628 -2033
rect 12516 -2105 12628 -2067
rect 12516 -2139 12555 -2105
rect 12589 -2139 12628 -2105
rect 12516 -2177 12628 -2139
rect 12516 -2211 12555 -2177
rect 12589 -2211 12628 -2177
rect 12516 -2249 12628 -2211
rect 12516 -2283 12555 -2249
rect 12589 -2283 12628 -2249
rect 12516 -2321 12628 -2283
rect 12516 -2355 12555 -2321
rect 12589 -2355 12628 -2321
rect 12516 -2393 12628 -2355
rect 12516 -2427 12555 -2393
rect 12589 -2427 12628 -2393
rect 12516 -2465 12628 -2427
rect 12516 -2499 12555 -2465
rect 12589 -2499 12628 -2465
rect 12516 -2537 12628 -2499
rect 12516 -2571 12555 -2537
rect 12589 -2571 12628 -2537
rect 12516 -2609 12628 -2571
rect 12516 -2643 12555 -2609
rect 12589 -2643 12628 -2609
rect 12516 -2681 12628 -2643
rect 12516 -2715 12555 -2681
rect 12589 -2715 12628 -2681
rect 12516 -2753 12628 -2715
rect 12516 -2787 12555 -2753
rect 12589 -2787 12628 -2753
rect 12516 -2825 12628 -2787
rect 12516 -2859 12555 -2825
rect 12589 -2859 12628 -2825
rect 12516 -2897 12628 -2859
rect 12516 -2931 12555 -2897
rect 12589 -2931 12628 -2897
rect 12516 -2969 12628 -2931
rect 12516 -3003 12555 -2969
rect 12589 -3003 12628 -2969
rect 12516 -3041 12628 -3003
rect 12516 -3075 12555 -3041
rect 12589 -3075 12628 -3041
rect 12516 -3113 12628 -3075
rect 12516 -3147 12555 -3113
rect 12589 -3147 12628 -3113
rect 12516 -3185 12628 -3147
rect 12516 -3219 12555 -3185
rect 12589 -3219 12628 -3185
rect 12516 -3257 12628 -3219
rect 12516 -3291 12555 -3257
rect 12589 -3291 12628 -3257
rect 12516 -3329 12628 -3291
rect 12516 -3363 12555 -3329
rect 12589 -3363 12628 -3329
rect 12516 -3401 12628 -3363
rect 12516 -3412 12555 -3401
rect 11326 -3435 12555 -3412
rect 12589 -3435 12628 -3401
rect 11326 -3472 12628 -3435
rect 10048 -5054 10108 -4964
rect 10048 -5106 10052 -5054
rect 10104 -5106 10108 -5054
rect 10048 -5411 10108 -5106
rect 10904 -5044 10964 -4964
rect 10904 -5054 10966 -5044
rect 10904 -5106 10910 -5054
rect 10962 -5106 10966 -5054
rect 10904 -5116 10966 -5106
rect 10464 -5272 10536 -5268
rect 10464 -5324 10474 -5272
rect 10526 -5324 10536 -5272
rect 10464 -5328 10536 -5324
rect 10470 -5518 10530 -5328
rect 10904 -5411 10964 -5116
rect 11326 -5154 11386 -3472
rect 11750 -3674 11810 -3472
rect 11754 -5154 11814 -4959
rect 12184 -5154 12244 -3472
rect 12516 -3473 12628 -3472
rect 12516 -3507 12555 -3473
rect 12589 -3507 12628 -3473
rect 12516 -3545 12628 -3507
rect 12516 -3579 12555 -3545
rect 12589 -3579 12628 -3545
rect 12516 -3617 12628 -3579
rect 12516 -3651 12555 -3617
rect 12589 -3651 12628 -3617
rect 12516 -3689 12628 -3651
rect 12516 -3723 12555 -3689
rect 12589 -3723 12628 -3689
rect 12516 -3761 12628 -3723
rect 12516 -3795 12555 -3761
rect 12589 -3795 12628 -3761
rect 12516 -3833 12628 -3795
rect 12516 -3867 12555 -3833
rect 12589 -3867 12628 -3833
rect 12516 -3905 12628 -3867
rect 12516 -3939 12555 -3905
rect 12589 -3939 12628 -3905
rect 12516 -3977 12628 -3939
rect 12516 -4011 12555 -3977
rect 12589 -4011 12628 -3977
rect 12516 -4049 12628 -4011
rect 12516 -4083 12555 -4049
rect 12589 -4083 12628 -4049
rect 12516 -4121 12628 -4083
rect 12516 -4155 12555 -4121
rect 12589 -4155 12628 -4121
rect 12516 -4193 12628 -4155
rect 12516 -4227 12555 -4193
rect 12589 -4227 12628 -4193
rect 12516 -4265 12628 -4227
rect 12516 -4299 12555 -4265
rect 12589 -4299 12628 -4265
rect 12516 -4337 12628 -4299
rect 12516 -4371 12555 -4337
rect 12589 -4371 12628 -4337
rect 12516 -4409 12628 -4371
rect 12516 -4443 12555 -4409
rect 12589 -4443 12628 -4409
rect 12516 -4481 12628 -4443
rect 12516 -4515 12555 -4481
rect 12589 -4515 12628 -4481
rect 12516 -4553 12628 -4515
rect 12516 -4587 12555 -4553
rect 12589 -4587 12628 -4553
rect 12516 -4625 12628 -4587
rect 12516 -4659 12555 -4625
rect 12589 -4659 12628 -4625
rect 12516 -4697 12628 -4659
rect 12516 -4731 12555 -4697
rect 12589 -4731 12628 -4697
rect 12516 -4769 12628 -4731
rect 12516 -4803 12555 -4769
rect 12589 -4803 12628 -4769
rect 12516 -4841 12628 -4803
rect 12516 -4875 12555 -4841
rect 12589 -4875 12628 -4841
rect 12516 -4913 12628 -4875
rect 12516 -4947 12555 -4913
rect 12589 -4947 12628 -4913
rect 12516 -4985 12628 -4947
rect 12516 -5019 12555 -4985
rect 12589 -5019 12628 -4985
rect 12516 -5057 12628 -5019
rect 12516 -5091 12555 -5057
rect 12589 -5091 12628 -5057
rect 12516 -5129 12628 -5091
rect 12516 -5154 12555 -5129
rect 11326 -5163 12555 -5154
rect 12589 -5163 12628 -5129
rect 11326 -5201 12628 -5163
rect 11326 -5214 12555 -5201
rect 11326 -5572 11386 -5214
rect 11754 -5410 11814 -5214
rect 12184 -5568 12244 -5214
rect 12516 -5235 12555 -5214
rect 12589 -5235 12628 -5201
rect 12516 -5273 12628 -5235
rect 12516 -5307 12555 -5273
rect 12589 -5307 12628 -5273
rect 12516 -5345 12628 -5307
rect 12516 -5379 12555 -5345
rect 12589 -5379 12628 -5345
rect 12516 -5417 12628 -5379
rect 12516 -5451 12555 -5417
rect 12589 -5451 12628 -5417
rect 12516 -5489 12628 -5451
rect 12516 -5523 12555 -5489
rect 12589 -5523 12628 -5489
rect 12516 -5561 12628 -5523
rect 12516 -5595 12555 -5561
rect 12589 -5595 12628 -5561
rect 12516 -5633 12628 -5595
rect 12516 -5667 12555 -5633
rect 12589 -5667 12628 -5633
rect 12516 -5705 12628 -5667
rect 12516 -5739 12555 -5705
rect 12589 -5739 12628 -5705
rect 12516 -5777 12628 -5739
rect 12516 -5811 12555 -5777
rect 12589 -5811 12628 -5777
rect 12516 -5849 12628 -5811
rect 12516 -5883 12555 -5849
rect 12589 -5883 12628 -5849
rect 12516 -5921 12628 -5883
rect 12516 -5955 12555 -5921
rect 12589 -5955 12628 -5921
rect 12516 -5993 12628 -5955
rect 12516 -6027 12555 -5993
rect 12589 -6027 12628 -5993
rect 12516 -6065 12628 -6027
rect 12516 -6099 12555 -6065
rect 12589 -6099 12628 -6065
rect 12516 -6137 12628 -6099
rect 12516 -6171 12555 -6137
rect 12589 -6171 12628 -6137
rect 12516 -6209 12628 -6171
rect 12516 -6243 12555 -6209
rect 12589 -6243 12628 -6209
rect 12516 -6281 12628 -6243
rect 12516 -6315 12555 -6281
rect 12589 -6315 12628 -6281
rect 12516 -6353 12628 -6315
rect 12516 -6387 12555 -6353
rect 12589 -6387 12628 -6353
rect 12516 -6425 12628 -6387
rect 12516 -6459 12555 -6425
rect 12589 -6459 12628 -6425
rect 12516 -6497 12628 -6459
rect 12516 -6531 12555 -6497
rect 12589 -6531 12628 -6497
rect 12516 -6569 12628 -6531
rect 10048 -6926 10108 -6697
rect 10904 -6926 10964 -6700
rect 10042 -6930 10114 -6926
rect 10042 -6982 10052 -6930
rect 10104 -6982 10114 -6930
rect 10042 -6986 10114 -6982
rect 10898 -6930 10970 -6926
rect 10898 -6982 10908 -6930
rect 10960 -6982 10970 -6930
rect 10898 -6986 10970 -6982
rect 11324 -7070 11384 -6594
rect 11750 -7070 11810 -6704
rect 12184 -7070 12244 -6588
rect 12516 -6603 12555 -6569
rect 12589 -6603 12628 -6569
rect 12516 -6641 12628 -6603
rect 12516 -6675 12555 -6641
rect 12589 -6675 12628 -6641
rect 12516 -6713 12628 -6675
rect 12516 -6747 12555 -6713
rect 12589 -6747 12628 -6713
rect 12516 -6785 12628 -6747
rect 12516 -6819 12555 -6785
rect 12589 -6819 12628 -6785
rect 12516 -6857 12628 -6819
rect 12516 -6891 12555 -6857
rect 12589 -6891 12628 -6857
rect 12516 -6929 12628 -6891
rect 12516 -6963 12555 -6929
rect 12589 -6963 12628 -6929
rect 12516 -7001 12628 -6963
rect 12516 -7035 12555 -7001
rect 12589 -7035 12628 -7001
rect -368 -7107 -329 -7073
rect -295 -7076 -256 -7073
rect 164 -7074 236 -7070
rect 164 -7076 174 -7074
rect -295 -7107 174 -7076
rect -368 -7126 174 -7107
rect 226 -7126 236 -7074
rect -368 -7130 236 -7126
rect 584 -7074 656 -7070
rect 584 -7126 594 -7074
rect 646 -7126 656 -7074
rect 584 -7130 656 -7126
rect 1024 -7074 1096 -7070
rect 1024 -7126 1034 -7074
rect 1086 -7126 1096 -7074
rect 1024 -7130 1096 -7126
rect 2742 -7074 2814 -7070
rect 2742 -7126 2752 -7074
rect 2804 -7126 2814 -7074
rect 2742 -7130 2814 -7126
rect 4456 -7074 4528 -7070
rect 4456 -7126 4466 -7074
rect 4518 -7126 4528 -7074
rect 4456 -7130 4528 -7126
rect 6174 -7074 6246 -7070
rect 6174 -7126 6184 -7074
rect 6236 -7126 6246 -7074
rect 6174 -7130 6246 -7126
rect 7888 -7074 7960 -7070
rect 7888 -7126 7898 -7074
rect 7950 -7126 7960 -7074
rect 7888 -7130 7960 -7126
rect 9602 -7074 9674 -7070
rect 9602 -7126 9612 -7074
rect 9664 -7126 9674 -7074
rect 9602 -7130 9674 -7126
rect 11318 -7074 11390 -7070
rect 11318 -7126 11328 -7074
rect 11380 -7126 11390 -7074
rect 11318 -7130 11390 -7126
rect 11744 -7074 11816 -7070
rect 11744 -7126 11754 -7074
rect 11806 -7126 11816 -7074
rect 11744 -7130 11816 -7126
rect 12178 -7072 12250 -7070
rect 12516 -7072 12628 -7035
rect 12178 -7073 12628 -7072
rect 12178 -7074 12555 -7073
rect 12178 -7126 12188 -7074
rect 12240 -7107 12555 -7074
rect 12589 -7107 12628 -7073
rect 12240 -7126 12628 -7107
rect 12178 -7130 12628 -7126
rect -368 -7136 230 -7130
rect -368 -7436 -256 -7136
rect 170 -7436 230 -7136
rect 590 -7436 650 -7130
rect 1030 -7436 1090 -7130
rect 2748 -7436 2808 -7130
rect 4462 -7436 4522 -7130
rect 6180 -7436 6240 -7130
rect 7894 -7436 7954 -7130
rect 9608 -7436 9668 -7130
rect 11324 -7436 11384 -7130
rect 11750 -7436 11810 -7130
rect 12184 -7132 12628 -7130
rect 12184 -7436 12244 -7132
rect 12516 -7436 12628 -7132
rect -368 -7475 12628 -7436
rect -368 -7509 -259 -7475
rect -225 -7509 -187 -7475
rect -153 -7509 -115 -7475
rect -81 -7509 -43 -7475
rect -9 -7509 29 -7475
rect 63 -7509 101 -7475
rect 135 -7509 173 -7475
rect 207 -7509 245 -7475
rect 279 -7509 317 -7475
rect 351 -7509 389 -7475
rect 423 -7509 461 -7475
rect 495 -7509 533 -7475
rect 567 -7509 605 -7475
rect 639 -7509 677 -7475
rect 711 -7509 749 -7475
rect 783 -7509 821 -7475
rect 855 -7509 893 -7475
rect 927 -7509 965 -7475
rect 999 -7509 1037 -7475
rect 1071 -7509 1109 -7475
rect 1143 -7509 1181 -7475
rect 1215 -7509 1253 -7475
rect 1287 -7509 1325 -7475
rect 1359 -7509 1397 -7475
rect 1431 -7509 1469 -7475
rect 1503 -7509 1541 -7475
rect 1575 -7509 1613 -7475
rect 1647 -7509 1685 -7475
rect 1719 -7509 1757 -7475
rect 1791 -7509 1829 -7475
rect 1863 -7509 1901 -7475
rect 1935 -7509 1973 -7475
rect 2007 -7509 2045 -7475
rect 2079 -7509 2117 -7475
rect 2151 -7509 2189 -7475
rect 2223 -7509 2261 -7475
rect 2295 -7509 2333 -7475
rect 2367 -7509 2405 -7475
rect 2439 -7509 2477 -7475
rect 2511 -7509 2549 -7475
rect 2583 -7509 2621 -7475
rect 2655 -7509 2693 -7475
rect 2727 -7509 2765 -7475
rect 2799 -7509 2837 -7475
rect 2871 -7509 2909 -7475
rect 2943 -7509 2981 -7475
rect 3015 -7509 3053 -7475
rect 3087 -7509 3125 -7475
rect 3159 -7509 3197 -7475
rect 3231 -7509 3269 -7475
rect 3303 -7509 3341 -7475
rect 3375 -7509 3413 -7475
rect 3447 -7509 3485 -7475
rect 3519 -7509 3557 -7475
rect 3591 -7509 3629 -7475
rect 3663 -7509 3701 -7475
rect 3735 -7509 3773 -7475
rect 3807 -7509 3845 -7475
rect 3879 -7509 3917 -7475
rect 3951 -7509 3989 -7475
rect 4023 -7509 4061 -7475
rect 4095 -7509 4133 -7475
rect 4167 -7509 4205 -7475
rect 4239 -7509 4277 -7475
rect 4311 -7509 4349 -7475
rect 4383 -7509 4421 -7475
rect 4455 -7509 4493 -7475
rect 4527 -7509 4565 -7475
rect 4599 -7509 4637 -7475
rect 4671 -7509 4709 -7475
rect 4743 -7509 4781 -7475
rect 4815 -7509 4853 -7475
rect 4887 -7509 4925 -7475
rect 4959 -7509 4997 -7475
rect 5031 -7509 5069 -7475
rect 5103 -7509 5141 -7475
rect 5175 -7509 5213 -7475
rect 5247 -7509 5285 -7475
rect 5319 -7509 5357 -7475
rect 5391 -7509 5429 -7475
rect 5463 -7509 5501 -7475
rect 5535 -7509 5573 -7475
rect 5607 -7509 5645 -7475
rect 5679 -7509 5717 -7475
rect 5751 -7509 5789 -7475
rect 5823 -7509 5861 -7475
rect 5895 -7509 5933 -7475
rect 5967 -7509 6005 -7475
rect 6039 -7509 6077 -7475
rect 6111 -7509 6149 -7475
rect 6183 -7509 6221 -7475
rect 6255 -7509 6293 -7475
rect 6327 -7509 6365 -7475
rect 6399 -7509 6437 -7475
rect 6471 -7509 6509 -7475
rect 6543 -7509 6581 -7475
rect 6615 -7509 6653 -7475
rect 6687 -7509 6725 -7475
rect 6759 -7509 6797 -7475
rect 6831 -7509 6869 -7475
rect 6903 -7509 6941 -7475
rect 6975 -7509 7013 -7475
rect 7047 -7509 7085 -7475
rect 7119 -7509 7157 -7475
rect 7191 -7509 7229 -7475
rect 7263 -7509 7301 -7475
rect 7335 -7509 7373 -7475
rect 7407 -7509 7445 -7475
rect 7479 -7509 7517 -7475
rect 7551 -7509 7589 -7475
rect 7623 -7509 7661 -7475
rect 7695 -7509 7733 -7475
rect 7767 -7509 7805 -7475
rect 7839 -7509 7877 -7475
rect 7911 -7509 7949 -7475
rect 7983 -7509 8021 -7475
rect 8055 -7509 8093 -7475
rect 8127 -7509 8165 -7475
rect 8199 -7509 8237 -7475
rect 8271 -7509 8309 -7475
rect 8343 -7509 8381 -7475
rect 8415 -7509 8453 -7475
rect 8487 -7509 8525 -7475
rect 8559 -7509 8597 -7475
rect 8631 -7509 8669 -7475
rect 8703 -7509 8741 -7475
rect 8775 -7509 8813 -7475
rect 8847 -7509 8885 -7475
rect 8919 -7509 8957 -7475
rect 8991 -7509 9029 -7475
rect 9063 -7509 9101 -7475
rect 9135 -7509 9173 -7475
rect 9207 -7509 9245 -7475
rect 9279 -7509 9317 -7475
rect 9351 -7509 9389 -7475
rect 9423 -7509 9461 -7475
rect 9495 -7509 9533 -7475
rect 9567 -7509 9605 -7475
rect 9639 -7509 9677 -7475
rect 9711 -7509 9749 -7475
rect 9783 -7509 9821 -7475
rect 9855 -7509 9893 -7475
rect 9927 -7509 9965 -7475
rect 9999 -7509 10037 -7475
rect 10071 -7509 10109 -7475
rect 10143 -7509 10181 -7475
rect 10215 -7509 10253 -7475
rect 10287 -7509 10325 -7475
rect 10359 -7509 10397 -7475
rect 10431 -7509 10469 -7475
rect 10503 -7509 10541 -7475
rect 10575 -7509 10613 -7475
rect 10647 -7509 10685 -7475
rect 10719 -7509 10757 -7475
rect 10791 -7509 10829 -7475
rect 10863 -7509 10901 -7475
rect 10935 -7509 10973 -7475
rect 11007 -7509 11045 -7475
rect 11079 -7509 11117 -7475
rect 11151 -7509 11189 -7475
rect 11223 -7509 11261 -7475
rect 11295 -7509 11333 -7475
rect 11367 -7509 11405 -7475
rect 11439 -7509 11477 -7475
rect 11511 -7509 11549 -7475
rect 11583 -7509 11621 -7475
rect 11655 -7509 11693 -7475
rect 11727 -7509 11765 -7475
rect 11799 -7509 11837 -7475
rect 11871 -7509 11909 -7475
rect 11943 -7509 11981 -7475
rect 12015 -7509 12053 -7475
rect 12087 -7509 12125 -7475
rect 12159 -7509 12197 -7475
rect 12231 -7509 12269 -7475
rect 12303 -7509 12341 -7475
rect 12375 -7509 12413 -7475
rect 12447 -7509 12485 -7475
rect 12519 -7509 12628 -7475
rect -368 -7548 12628 -7509
rect -368 -7811 12628 -7772
rect -368 -7845 -259 -7811
rect -225 -7845 -187 -7811
rect -153 -7845 -115 -7811
rect -81 -7845 -43 -7811
rect -9 -7845 29 -7811
rect 63 -7845 101 -7811
rect 135 -7845 173 -7811
rect 207 -7845 245 -7811
rect 279 -7845 317 -7811
rect 351 -7845 389 -7811
rect 423 -7845 461 -7811
rect 495 -7845 533 -7811
rect 567 -7845 605 -7811
rect 639 -7845 677 -7811
rect 711 -7845 749 -7811
rect 783 -7845 821 -7811
rect 855 -7845 893 -7811
rect 927 -7845 965 -7811
rect 999 -7845 1037 -7811
rect 1071 -7845 1109 -7811
rect 1143 -7845 1181 -7811
rect 1215 -7845 1253 -7811
rect 1287 -7845 1325 -7811
rect 1359 -7845 1397 -7811
rect 1431 -7845 1469 -7811
rect 1503 -7845 1541 -7811
rect 1575 -7845 1613 -7811
rect 1647 -7845 1685 -7811
rect 1719 -7845 1757 -7811
rect 1791 -7845 1829 -7811
rect 1863 -7845 1901 -7811
rect 1935 -7845 1973 -7811
rect 2007 -7845 2045 -7811
rect 2079 -7845 2117 -7811
rect 2151 -7845 2189 -7811
rect 2223 -7845 2261 -7811
rect 2295 -7845 2333 -7811
rect 2367 -7845 2405 -7811
rect 2439 -7845 2477 -7811
rect 2511 -7845 2549 -7811
rect 2583 -7845 2621 -7811
rect 2655 -7845 2693 -7811
rect 2727 -7845 2765 -7811
rect 2799 -7845 2837 -7811
rect 2871 -7845 2909 -7811
rect 2943 -7845 2981 -7811
rect 3015 -7845 3053 -7811
rect 3087 -7845 3125 -7811
rect 3159 -7845 3197 -7811
rect 3231 -7845 3269 -7811
rect 3303 -7845 3341 -7811
rect 3375 -7845 3413 -7811
rect 3447 -7845 3485 -7811
rect 3519 -7845 3557 -7811
rect 3591 -7845 3629 -7811
rect 3663 -7845 3701 -7811
rect 3735 -7845 3773 -7811
rect 3807 -7845 3845 -7811
rect 3879 -7845 3917 -7811
rect 3951 -7845 3989 -7811
rect 4023 -7845 4061 -7811
rect 4095 -7845 4133 -7811
rect 4167 -7845 4205 -7811
rect 4239 -7845 4277 -7811
rect 4311 -7845 4349 -7811
rect 4383 -7845 4421 -7811
rect 4455 -7845 4493 -7811
rect 4527 -7845 4565 -7811
rect 4599 -7845 4637 -7811
rect 4671 -7845 4709 -7811
rect 4743 -7845 4781 -7811
rect 4815 -7845 4853 -7811
rect 4887 -7845 4925 -7811
rect 4959 -7845 4997 -7811
rect 5031 -7845 5069 -7811
rect 5103 -7845 5141 -7811
rect 5175 -7845 5213 -7811
rect 5247 -7845 5285 -7811
rect 5319 -7845 5357 -7811
rect 5391 -7845 5429 -7811
rect 5463 -7845 5501 -7811
rect 5535 -7845 5573 -7811
rect 5607 -7845 5645 -7811
rect 5679 -7845 5717 -7811
rect 5751 -7845 5789 -7811
rect 5823 -7845 5861 -7811
rect 5895 -7845 5933 -7811
rect 5967 -7845 6005 -7811
rect 6039 -7845 6077 -7811
rect 6111 -7845 6149 -7811
rect 6183 -7845 6221 -7811
rect 6255 -7845 6293 -7811
rect 6327 -7845 6365 -7811
rect 6399 -7845 6437 -7811
rect 6471 -7845 6509 -7811
rect 6543 -7845 6581 -7811
rect 6615 -7845 6653 -7811
rect 6687 -7845 6725 -7811
rect 6759 -7845 6797 -7811
rect 6831 -7845 6869 -7811
rect 6903 -7845 6941 -7811
rect 6975 -7845 7013 -7811
rect 7047 -7845 7085 -7811
rect 7119 -7845 7157 -7811
rect 7191 -7845 7229 -7811
rect 7263 -7845 7301 -7811
rect 7335 -7845 7373 -7811
rect 7407 -7845 7445 -7811
rect 7479 -7845 7517 -7811
rect 7551 -7845 7589 -7811
rect 7623 -7845 7661 -7811
rect 7695 -7845 7733 -7811
rect 7767 -7845 7805 -7811
rect 7839 -7845 7877 -7811
rect 7911 -7845 7949 -7811
rect 7983 -7845 8021 -7811
rect 8055 -7845 8093 -7811
rect 8127 -7845 8165 -7811
rect 8199 -7845 8237 -7811
rect 8271 -7845 8309 -7811
rect 8343 -7845 8381 -7811
rect 8415 -7845 8453 -7811
rect 8487 -7845 8525 -7811
rect 8559 -7845 8597 -7811
rect 8631 -7845 8669 -7811
rect 8703 -7845 8741 -7811
rect 8775 -7845 8813 -7811
rect 8847 -7845 8885 -7811
rect 8919 -7845 8957 -7811
rect 8991 -7845 9029 -7811
rect 9063 -7845 9101 -7811
rect 9135 -7845 9173 -7811
rect 9207 -7845 9245 -7811
rect 9279 -7845 9317 -7811
rect 9351 -7845 9389 -7811
rect 9423 -7845 9461 -7811
rect 9495 -7845 9533 -7811
rect 9567 -7845 9605 -7811
rect 9639 -7845 9677 -7811
rect 9711 -7845 9749 -7811
rect 9783 -7845 9821 -7811
rect 9855 -7845 9893 -7811
rect 9927 -7845 9965 -7811
rect 9999 -7845 10037 -7811
rect 10071 -7845 10109 -7811
rect 10143 -7845 10181 -7811
rect 10215 -7845 10253 -7811
rect 10287 -7845 10325 -7811
rect 10359 -7845 10397 -7811
rect 10431 -7845 10469 -7811
rect 10503 -7845 10541 -7811
rect 10575 -7845 10613 -7811
rect 10647 -7845 10685 -7811
rect 10719 -7845 10757 -7811
rect 10791 -7845 10829 -7811
rect 10863 -7845 10901 -7811
rect 10935 -7845 10973 -7811
rect 11007 -7845 11045 -7811
rect 11079 -7845 11117 -7811
rect 11151 -7845 11189 -7811
rect 11223 -7845 11261 -7811
rect 11295 -7845 11333 -7811
rect 11367 -7845 11405 -7811
rect 11439 -7845 11477 -7811
rect 11511 -7845 11549 -7811
rect 11583 -7845 11621 -7811
rect 11655 -7845 11693 -7811
rect 11727 -7845 11765 -7811
rect 11799 -7845 11837 -7811
rect 11871 -7845 11909 -7811
rect 11943 -7845 11981 -7811
rect 12015 -7845 12053 -7811
rect 12087 -7845 12125 -7811
rect 12159 -7845 12197 -7811
rect 12231 -7845 12269 -7811
rect 12303 -7845 12341 -7811
rect 12375 -7845 12413 -7811
rect 12447 -7845 12485 -7811
rect 12519 -7845 12628 -7811
rect -368 -7884 12628 -7845
rect -368 -7999 -256 -7884
rect -368 -8033 -329 -7999
rect -295 -8033 -256 -7999
rect -368 -8071 -256 -8033
rect -368 -8105 -329 -8071
rect -295 -8105 -256 -8071
rect -368 -8143 -256 -8105
rect -368 -8177 -329 -8143
rect -295 -8177 -256 -8143
rect -368 -8215 -256 -8177
rect -368 -8249 -329 -8215
rect -295 -8249 -256 -8215
rect 4792 -8166 4864 -8162
rect 4792 -8218 4802 -8166
rect 4854 -8218 4864 -8166
rect 4792 -8222 4864 -8218
rect -368 -8287 -256 -8249
rect -368 -8321 -329 -8287
rect -295 -8321 -256 -8287
rect -368 -8359 -256 -8321
rect -368 -8393 -329 -8359
rect -295 -8393 -256 -8359
rect -368 -8431 -256 -8393
rect -368 -8465 -329 -8431
rect -295 -8465 -256 -8431
rect -368 -8503 -256 -8465
rect -368 -8537 -329 -8503
rect -295 -8537 -256 -8503
rect -368 -8575 -256 -8537
rect -368 -8609 -329 -8575
rect -295 -8609 -256 -8575
rect -368 -8647 -256 -8609
rect -368 -8681 -329 -8647
rect -295 -8681 -256 -8647
rect -368 -8719 -256 -8681
rect -368 -8753 -329 -8719
rect -295 -8753 -256 -8719
rect -368 -8791 -256 -8753
rect -368 -8825 -329 -8791
rect -295 -8825 -256 -8791
rect -368 -8863 -256 -8825
rect -368 -8897 -329 -8863
rect -295 -8897 -256 -8863
rect -368 -8935 -256 -8897
rect -368 -8969 -329 -8935
rect -295 -8969 -256 -8935
rect -368 -9007 -256 -8969
rect -368 -9041 -329 -9007
rect -295 -9041 -256 -9007
rect -368 -9079 -256 -9041
rect -368 -9113 -329 -9079
rect -295 -9113 -256 -9079
rect 4798 -9092 4858 -8222
rect 4896 -8272 4956 -7884
rect 5124 -8272 5184 -7884
rect 4896 -8332 5184 -8272
rect 5576 -8274 5648 -8270
rect 5576 -8326 5586 -8274
rect 5638 -8326 5648 -8274
rect 5576 -8330 5648 -8326
rect 4896 -9032 4956 -8332
rect 5124 -8420 5184 -8332
rect 5582 -8424 5642 -8330
rect 5124 -9032 5184 -8892
rect 5356 -8978 5416 -8826
rect 4896 -9092 5184 -9032
rect 5350 -8982 5422 -8978
rect 5350 -9034 5360 -8982
rect 5412 -9034 5422 -8982
rect 5350 -9038 5422 -9034
rect -368 -9151 -256 -9113
rect -368 -9185 -329 -9151
rect -295 -9185 -256 -9151
rect 4792 -9096 4864 -9092
rect 4792 -9148 4802 -9096
rect 4854 -9148 4864 -9096
rect 4792 -9152 4864 -9148
rect -368 -9223 -256 -9185
rect -368 -9257 -329 -9223
rect -295 -9257 -256 -9223
rect -368 -9295 -256 -9257
rect -368 -9329 -329 -9295
rect -295 -9329 -256 -9295
rect -368 -9367 -256 -9329
rect -368 -9401 -329 -9367
rect -295 -9401 -256 -9367
rect -368 -9439 -256 -9401
rect -368 -9473 -329 -9439
rect -295 -9473 -256 -9439
rect -368 -9511 -256 -9473
rect -368 -9545 -329 -9511
rect -295 -9545 -256 -9511
rect -368 -9583 -256 -9545
rect -368 -9617 -329 -9583
rect -295 -9617 -256 -9583
rect -368 -9655 -256 -9617
rect -368 -9689 -329 -9655
rect -295 -9689 -256 -9655
rect -368 -9727 -256 -9689
rect -368 -9761 -329 -9727
rect -295 -9761 -256 -9727
rect -368 -9799 -256 -9761
rect -368 -9833 -329 -9799
rect -295 -9833 -256 -9799
rect -368 -9871 -256 -9833
rect -368 -9905 -329 -9871
rect -295 -9905 -256 -9871
rect -368 -9943 -256 -9905
rect -368 -9977 -329 -9943
rect -295 -9977 -256 -9943
rect -368 -10015 -256 -9977
rect -368 -10049 -329 -10015
rect -295 -10049 -256 -10015
rect -368 -10087 -256 -10049
rect -368 -10121 -329 -10087
rect -295 -10121 -256 -10087
rect 4896 -9794 4956 -9092
rect 5124 -9228 5184 -9092
rect 5350 -9096 5422 -9092
rect 5350 -9148 5360 -9096
rect 5412 -9148 5422 -9096
rect 5350 -9152 5422 -9148
rect 5356 -9316 5416 -9152
rect 5584 -9224 5644 -8898
rect 5124 -9794 5184 -9696
rect 5584 -9792 5644 -9690
rect 4896 -9854 5184 -9794
rect 5578 -9796 5650 -9792
rect 5578 -9848 5588 -9796
rect 5640 -9848 5650 -9796
rect 5578 -9852 5650 -9848
rect 4896 -10100 4956 -9854
rect 5124 -10100 5184 -9854
rect 5814 -9918 5874 -7884
rect 6264 -8166 6336 -8162
rect 6264 -8218 6274 -8166
rect 6326 -8218 6336 -8166
rect 6264 -8222 6336 -8218
rect 6036 -8274 6108 -8270
rect 6036 -8326 6046 -8274
rect 6098 -8326 6108 -8274
rect 6036 -8330 6108 -8326
rect 6042 -8424 6102 -8330
rect 6270 -8494 6330 -8222
rect 6498 -8274 6570 -8270
rect 6498 -8326 6508 -8274
rect 6560 -8326 6570 -8274
rect 6498 -8330 6570 -8326
rect 6504 -8424 6564 -8330
rect 6044 -9228 6104 -8892
rect 6264 -8982 6336 -8978
rect 6264 -9034 6274 -8982
rect 6326 -9034 6336 -8982
rect 6264 -9038 6336 -9034
rect 6270 -9324 6330 -9038
rect 6504 -9228 6564 -8892
rect 6044 -9792 6104 -9698
rect 6504 -9792 6564 -9696
rect 6038 -9796 6110 -9792
rect 6038 -9848 6048 -9796
rect 6100 -9848 6110 -9796
rect 6038 -9852 6110 -9848
rect 6498 -9796 6570 -9792
rect 6498 -9848 6508 -9796
rect 6560 -9848 6570 -9796
rect 6498 -9852 6570 -9848
rect 6728 -9918 6788 -7884
rect 7422 -8268 7482 -7884
rect 7646 -8268 7706 -7884
rect 6954 -8274 7026 -8270
rect 6954 -8326 6964 -8274
rect 7016 -8326 7026 -8274
rect 6954 -8330 7026 -8326
rect 7422 -8328 7706 -8268
rect 6960 -8424 7020 -8330
rect 7422 -8416 7482 -8328
rect 6964 -9228 7024 -8892
rect 7186 -8978 7246 -8804
rect 7180 -8982 7252 -8978
rect 7180 -9034 7190 -8982
rect 7242 -9034 7252 -8982
rect 7180 -9038 7252 -9034
rect 7424 -9034 7484 -8892
rect 7646 -9034 7706 -8328
rect 7180 -9096 7252 -9092
rect 7180 -9148 7190 -9096
rect 7242 -9148 7252 -9096
rect 7180 -9152 7252 -9148
rect 7424 -9094 7706 -9034
rect 7186 -9314 7246 -9152
rect 7424 -9228 7484 -9094
rect 6958 -9792 7018 -9694
rect 7422 -9790 7482 -9698
rect 7646 -9790 7706 -9094
rect 6952 -9796 7024 -9792
rect 6952 -9848 6962 -9796
rect 7014 -9848 7024 -9796
rect 6952 -9852 7024 -9848
rect 7422 -9850 7706 -9790
rect 5808 -9922 5880 -9918
rect 5808 -9974 5818 -9922
rect 5870 -9974 5880 -9922
rect 5808 -9978 5880 -9974
rect 6722 -9922 6794 -9918
rect 6722 -9974 6732 -9922
rect 6784 -9974 6794 -9922
rect 6722 -9978 6794 -9974
rect 5814 -10100 5874 -9978
rect 6728 -10100 6788 -9978
rect 7422 -10100 7482 -9850
rect 7646 -10100 7706 -9850
rect 12516 -7999 12628 -7884
rect 12516 -8033 12555 -7999
rect 12589 -8033 12628 -7999
rect 12516 -8071 12628 -8033
rect 12516 -8105 12555 -8071
rect 12589 -8105 12628 -8071
rect 12516 -8143 12628 -8105
rect 12516 -8177 12555 -8143
rect 12589 -8177 12628 -8143
rect 12516 -8215 12628 -8177
rect 12516 -8249 12555 -8215
rect 12589 -8249 12628 -8215
rect 12516 -8287 12628 -8249
rect 12516 -8321 12555 -8287
rect 12589 -8321 12628 -8287
rect 12516 -8359 12628 -8321
rect 12516 -8393 12555 -8359
rect 12589 -8393 12628 -8359
rect 12516 -8431 12628 -8393
rect 12516 -8465 12555 -8431
rect 12589 -8465 12628 -8431
rect 12516 -8503 12628 -8465
rect 12516 -8537 12555 -8503
rect 12589 -8537 12628 -8503
rect 12516 -8575 12628 -8537
rect 12516 -8609 12555 -8575
rect 12589 -8609 12628 -8575
rect 12516 -8647 12628 -8609
rect 12516 -8681 12555 -8647
rect 12589 -8681 12628 -8647
rect 12516 -8719 12628 -8681
rect 12516 -8753 12555 -8719
rect 12589 -8753 12628 -8719
rect 12516 -8791 12628 -8753
rect 12516 -8825 12555 -8791
rect 12589 -8825 12628 -8791
rect 12516 -8863 12628 -8825
rect 12516 -8897 12555 -8863
rect 12589 -8897 12628 -8863
rect 12516 -8935 12628 -8897
rect 12516 -8969 12555 -8935
rect 12589 -8969 12628 -8935
rect 12516 -9007 12628 -8969
rect 12516 -9041 12555 -9007
rect 12589 -9041 12628 -9007
rect 12516 -9079 12628 -9041
rect 12516 -9113 12555 -9079
rect 12589 -9113 12628 -9079
rect 12516 -9151 12628 -9113
rect 12516 -9185 12555 -9151
rect 12589 -9185 12628 -9151
rect 12516 -9223 12628 -9185
rect 12516 -9257 12555 -9223
rect 12589 -9257 12628 -9223
rect 12516 -9295 12628 -9257
rect 12516 -9329 12555 -9295
rect 12589 -9329 12628 -9295
rect 12516 -9367 12628 -9329
rect 12516 -9401 12555 -9367
rect 12589 -9401 12628 -9367
rect 12516 -9439 12628 -9401
rect 12516 -9473 12555 -9439
rect 12589 -9473 12628 -9439
rect 12516 -9511 12628 -9473
rect 12516 -9545 12555 -9511
rect 12589 -9545 12628 -9511
rect 12516 -9583 12628 -9545
rect 12516 -9617 12555 -9583
rect 12589 -9617 12628 -9583
rect 12516 -9655 12628 -9617
rect 12516 -9689 12555 -9655
rect 12589 -9689 12628 -9655
rect 12516 -9727 12628 -9689
rect 12516 -9761 12555 -9727
rect 12589 -9761 12628 -9727
rect 12516 -9799 12628 -9761
rect 12516 -9833 12555 -9799
rect 12589 -9833 12628 -9799
rect 12516 -9871 12628 -9833
rect 12516 -9905 12555 -9871
rect 12589 -9905 12628 -9871
rect 12516 -9943 12628 -9905
rect 12516 -9977 12555 -9943
rect 12589 -9977 12628 -9943
rect 12516 -10015 12628 -9977
rect 12516 -10049 12555 -10015
rect 12589 -10049 12628 -10015
rect 12516 -10087 12628 -10049
rect -368 -10159 -256 -10121
rect -368 -10193 -329 -10159
rect -295 -10193 -256 -10159
rect -368 -10231 -256 -10193
rect -368 -10265 -329 -10231
rect -295 -10265 -256 -10231
rect -368 -10303 -256 -10265
rect -368 -10337 -329 -10303
rect -295 -10337 -256 -10303
rect -368 -10375 -256 -10337
rect -368 -10409 -329 -10375
rect -295 -10409 -256 -10375
rect -368 -10416 -256 -10409
rect 4664 -10195 7854 -10100
rect -368 -10444 354 -10416
rect -368 -10447 -238 -10444
rect -368 -10481 -329 -10447
rect -295 -10481 -238 -10447
rect -368 -10519 -238 -10481
rect -368 -10553 -329 -10519
rect -295 -10553 -238 -10519
rect -368 -10688 -238 -10553
rect 326 -10688 354 -10444
rect 4664 -10567 4736 -10195
rect 7796 -10567 7854 -10195
rect 12516 -10121 12555 -10087
rect 12589 -10121 12628 -10087
rect 12516 -10159 12628 -10121
rect 12516 -10193 12555 -10159
rect 12589 -10193 12628 -10159
rect 12516 -10231 12628 -10193
rect 12516 -10265 12555 -10231
rect 12589 -10265 12628 -10231
rect 12516 -10303 12628 -10265
rect 12516 -10337 12555 -10303
rect 12589 -10337 12628 -10303
rect 12516 -10375 12628 -10337
rect 12516 -10409 12555 -10375
rect 12589 -10409 12628 -10375
rect 12516 -10416 12628 -10409
rect 4664 -10646 7854 -10567
rect 11906 -10444 12628 -10416
rect -368 -10716 354 -10688
rect 11906 -10688 11934 -10444
rect 12498 -10447 12628 -10444
rect 12498 -10481 12555 -10447
rect 12589 -10481 12628 -10447
rect 12498 -10519 12628 -10481
rect 12498 -10553 12555 -10519
rect 12589 -10553 12628 -10519
rect 12498 -10688 12628 -10553
rect 11906 -10716 12628 -10688
rect -368 -10755 12628 -10716
rect -368 -10789 -259 -10755
rect -225 -10789 -187 -10755
rect -153 -10789 -115 -10755
rect -81 -10789 -43 -10755
rect -9 -10789 29 -10755
rect 63 -10789 101 -10755
rect 135 -10789 173 -10755
rect 207 -10789 245 -10755
rect 279 -10789 317 -10755
rect 351 -10789 389 -10755
rect 423 -10789 461 -10755
rect 495 -10789 533 -10755
rect 567 -10789 605 -10755
rect 639 -10789 677 -10755
rect 711 -10789 749 -10755
rect 783 -10789 821 -10755
rect 855 -10789 893 -10755
rect 927 -10789 965 -10755
rect 999 -10789 1037 -10755
rect 1071 -10789 1109 -10755
rect 1143 -10789 1181 -10755
rect 1215 -10789 1253 -10755
rect 1287 -10789 1325 -10755
rect 1359 -10789 1397 -10755
rect 1431 -10789 1469 -10755
rect 1503 -10789 1541 -10755
rect 1575 -10789 1613 -10755
rect 1647 -10789 1685 -10755
rect 1719 -10789 1757 -10755
rect 1791 -10789 1829 -10755
rect 1863 -10789 1901 -10755
rect 1935 -10789 1973 -10755
rect 2007 -10789 2045 -10755
rect 2079 -10789 2117 -10755
rect 2151 -10789 2189 -10755
rect 2223 -10789 2261 -10755
rect 2295 -10789 2333 -10755
rect 2367 -10789 2405 -10755
rect 2439 -10789 2477 -10755
rect 2511 -10789 2549 -10755
rect 2583 -10789 2621 -10755
rect 2655 -10789 2693 -10755
rect 2727 -10789 2765 -10755
rect 2799 -10789 2837 -10755
rect 2871 -10789 2909 -10755
rect 2943 -10789 2981 -10755
rect 3015 -10789 3053 -10755
rect 3087 -10789 3125 -10755
rect 3159 -10789 3197 -10755
rect 3231 -10789 3269 -10755
rect 3303 -10789 3341 -10755
rect 3375 -10789 3413 -10755
rect 3447 -10789 3485 -10755
rect 3519 -10789 3557 -10755
rect 3591 -10789 3629 -10755
rect 3663 -10789 3701 -10755
rect 3735 -10789 3773 -10755
rect 3807 -10789 3845 -10755
rect 3879 -10789 3917 -10755
rect 3951 -10789 3989 -10755
rect 4023 -10789 4061 -10755
rect 4095 -10789 4133 -10755
rect 4167 -10789 4205 -10755
rect 4239 -10789 4277 -10755
rect 4311 -10789 4349 -10755
rect 4383 -10789 4421 -10755
rect 4455 -10789 4493 -10755
rect 4527 -10789 4565 -10755
rect 4599 -10789 4637 -10755
rect 4671 -10789 4709 -10755
rect 4743 -10789 4781 -10755
rect 4815 -10789 4853 -10755
rect 4887 -10789 4925 -10755
rect 4959 -10789 4997 -10755
rect 5031 -10789 5069 -10755
rect 5103 -10789 5141 -10755
rect 5175 -10789 5213 -10755
rect 5247 -10789 5285 -10755
rect 5319 -10789 5357 -10755
rect 5391 -10789 5429 -10755
rect 5463 -10789 5501 -10755
rect 5535 -10789 5573 -10755
rect 5607 -10789 5645 -10755
rect 5679 -10789 5717 -10755
rect 5751 -10789 5789 -10755
rect 5823 -10789 5861 -10755
rect 5895 -10789 5933 -10755
rect 5967 -10789 6005 -10755
rect 6039 -10789 6077 -10755
rect 6111 -10789 6149 -10755
rect 6183 -10789 6221 -10755
rect 6255 -10789 6293 -10755
rect 6327 -10789 6365 -10755
rect 6399 -10789 6437 -10755
rect 6471 -10789 6509 -10755
rect 6543 -10789 6581 -10755
rect 6615 -10789 6653 -10755
rect 6687 -10789 6725 -10755
rect 6759 -10789 6797 -10755
rect 6831 -10789 6869 -10755
rect 6903 -10789 6941 -10755
rect 6975 -10789 7013 -10755
rect 7047 -10789 7085 -10755
rect 7119 -10789 7157 -10755
rect 7191 -10789 7229 -10755
rect 7263 -10789 7301 -10755
rect 7335 -10789 7373 -10755
rect 7407 -10789 7445 -10755
rect 7479 -10789 7517 -10755
rect 7551 -10789 7589 -10755
rect 7623 -10789 7661 -10755
rect 7695 -10789 7733 -10755
rect 7767 -10789 7805 -10755
rect 7839 -10789 7877 -10755
rect 7911 -10789 7949 -10755
rect 7983 -10789 8021 -10755
rect 8055 -10789 8093 -10755
rect 8127 -10789 8165 -10755
rect 8199 -10789 8237 -10755
rect 8271 -10789 8309 -10755
rect 8343 -10789 8381 -10755
rect 8415 -10789 8453 -10755
rect 8487 -10789 8525 -10755
rect 8559 -10789 8597 -10755
rect 8631 -10789 8669 -10755
rect 8703 -10789 8741 -10755
rect 8775 -10789 8813 -10755
rect 8847 -10789 8885 -10755
rect 8919 -10789 8957 -10755
rect 8991 -10789 9029 -10755
rect 9063 -10789 9101 -10755
rect 9135 -10789 9173 -10755
rect 9207 -10789 9245 -10755
rect 9279 -10789 9317 -10755
rect 9351 -10789 9389 -10755
rect 9423 -10789 9461 -10755
rect 9495 -10789 9533 -10755
rect 9567 -10789 9605 -10755
rect 9639 -10789 9677 -10755
rect 9711 -10789 9749 -10755
rect 9783 -10789 9821 -10755
rect 9855 -10789 9893 -10755
rect 9927 -10789 9965 -10755
rect 9999 -10789 10037 -10755
rect 10071 -10789 10109 -10755
rect 10143 -10789 10181 -10755
rect 10215 -10789 10253 -10755
rect 10287 -10789 10325 -10755
rect 10359 -10789 10397 -10755
rect 10431 -10789 10469 -10755
rect 10503 -10789 10541 -10755
rect 10575 -10789 10613 -10755
rect 10647 -10789 10685 -10755
rect 10719 -10789 10757 -10755
rect 10791 -10789 10829 -10755
rect 10863 -10789 10901 -10755
rect 10935 -10789 10973 -10755
rect 11007 -10789 11045 -10755
rect 11079 -10789 11117 -10755
rect 11151 -10789 11189 -10755
rect 11223 -10789 11261 -10755
rect 11295 -10789 11333 -10755
rect 11367 -10789 11405 -10755
rect 11439 -10789 11477 -10755
rect 11511 -10789 11549 -10755
rect 11583 -10789 11621 -10755
rect 11655 -10789 11693 -10755
rect 11727 -10789 11765 -10755
rect 11799 -10789 11837 -10755
rect 11871 -10789 11909 -10755
rect 11943 -10789 11981 -10755
rect 12015 -10789 12053 -10755
rect 12087 -10789 12125 -10755
rect 12159 -10789 12197 -10755
rect 12231 -10789 12269 -10755
rect 12303 -10789 12341 -10755
rect 12375 -10789 12413 -10755
rect 12447 -10789 12485 -10755
rect 12519 -10789 12628 -10755
rect -368 -10828 12628 -10789
<< via1 >>
rect -238 2544 326 2788
rect 11934 2544 12498 2788
rect 171 2256 12255 2372
rect 176 2054 228 2106
rect 600 2054 652 2106
rect 1036 2054 1088 2106
rect 2750 2054 2802 2106
rect 4470 2054 4522 2106
rect 6178 2054 6230 2106
rect 7898 2054 7950 2106
rect 9612 2054 9664 2106
rect 11330 2054 11382 2106
rect 11758 2054 11810 2106
rect 12190 2054 12242 2106
rect -88 1790 -36 1842
rect 54 1662 106 1714
rect 1462 1926 1514 1978
rect 2316 1926 2368 1978
rect 3176 1926 3228 1978
rect 4036 1926 4088 1978
rect 4896 1926 4948 1978
rect 5756 1926 5808 1978
rect 6616 1926 6668 1978
rect 7476 1926 7528 1978
rect 8336 1926 8388 1978
rect 9176 1926 9228 1978
rect 8756 1662 8808 1714
rect 10034 1926 10086 1978
rect 10896 1926 10948 1978
rect 10472 1790 10524 1842
rect 54 0 106 52
rect -88 -106 -36 -54
rect -88 -1636 -36 -1584
rect 1892 100 1944 152
rect 1894 -106 1946 -54
rect 54 -1842 106 -1790
rect 1462 -1740 1514 -1688
rect 2324 -1740 2376 -1688
rect 54 -3480 106 -3428
rect -88 -3586 -36 -3534
rect 1892 -3380 1944 -3328
rect 1894 -3586 1946 -3534
rect 1464 -5106 1516 -5054
rect 2324 -5106 2376 -5054
rect 1892 -5324 1944 -5272
rect 1460 -6982 1512 -6930
rect 2330 -6982 2382 -6930
rect 3474 0 3526 52
rect 3608 -2 3660 50
rect 3186 -1740 3238 -1688
rect 4044 -1740 4096 -1688
rect 3474 -3480 3526 -3428
rect 3608 -3482 3660 -3430
rect 5324 -106 5376 -54
rect 7170 -106 7222 -54
rect 4904 -1740 4956 -1688
rect 5748 -1740 5800 -1688
rect 4466 -3588 4518 -3536
rect 3180 -5106 3232 -5054
rect 4046 -5106 4098 -5054
rect 3610 -5210 3662 -5158
rect 3188 -6982 3240 -6930
rect 4046 -6982 4098 -6930
rect 6618 -1740 6670 -1688
rect 7484 -1740 7536 -1688
rect 6184 -3252 6236 -3200
rect 5324 -3586 5376 -3534
rect 7170 -3586 7222 -3534
rect 8760 -2 8812 50
rect 8340 -1740 8392 -1688
rect 9196 -1740 9248 -1688
rect 8756 -1842 8808 -1790
rect 7898 -3586 7950 -3534
rect 4902 -5106 4954 -5054
rect 5750 -5106 5802 -5054
rect 5324 -6856 5376 -6804
rect 4904 -6982 4956 -6930
rect 5762 -6982 5814 -6930
rect 6604 -5106 6656 -5054
rect 7484 -5106 7536 -5054
rect 7042 -6856 7094 -6804
rect 6620 -6982 6672 -6930
rect 7478 -6982 7530 -6930
rect 8760 -3482 8812 -3430
rect 8338 -5106 8390 -5054
rect 9196 -5110 9248 -5058
rect 8756 -5210 8808 -5158
rect 8336 -6982 8388 -6930
rect 9194 -6982 9246 -6930
rect 10474 100 10526 152
rect 10472 -1636 10524 -1584
rect 10050 -1740 10102 -1688
rect 10908 -1740 10960 -1688
rect 10474 -3380 10526 -3328
rect 10052 -5106 10104 -5054
rect 10910 -5106 10962 -5054
rect 10474 -5324 10526 -5272
rect 10052 -6982 10104 -6930
rect 10908 -6982 10960 -6930
rect 174 -7126 226 -7074
rect 594 -7126 646 -7074
rect 1034 -7126 1086 -7074
rect 2752 -7126 2804 -7074
rect 4466 -7126 4518 -7074
rect 6184 -7126 6236 -7074
rect 7898 -7126 7950 -7074
rect 9612 -7126 9664 -7074
rect 11328 -7126 11380 -7074
rect 11754 -7126 11806 -7074
rect 12188 -7126 12240 -7074
rect 4802 -8218 4854 -8166
rect 5586 -8326 5638 -8274
rect 5360 -9034 5412 -8982
rect 4802 -9148 4854 -9096
rect 5360 -9148 5412 -9096
rect 5588 -9848 5640 -9796
rect 6274 -8218 6326 -8166
rect 6046 -8326 6098 -8274
rect 6508 -8326 6560 -8274
rect 6274 -9034 6326 -8982
rect 6048 -9848 6100 -9796
rect 6508 -9848 6560 -9796
rect 6964 -8326 7016 -8274
rect 7190 -9034 7242 -8982
rect 7190 -9148 7242 -9096
rect 6962 -9848 7014 -9796
rect 5818 -9974 5870 -9922
rect 6732 -9974 6784 -9922
rect -238 -10688 326 -10444
rect 4736 -10567 7796 -10195
rect 11934 -10688 12498 -10444
<< metal2 >>
rect -256 2814 344 2826
rect -256 2788 -224 2814
rect 312 2788 344 2814
rect -256 2544 -238 2788
rect 326 2544 344 2788
rect -256 2518 -224 2544
rect 312 2518 344 2544
rect -256 2506 344 2518
rect 11916 2814 12516 2826
rect 11916 2788 11948 2814
rect 12484 2788 12516 2814
rect 11916 2544 11934 2788
rect 12498 2544 12516 2788
rect 11916 2518 11948 2544
rect 12484 2518 12516 2544
rect 11916 2506 12516 2518
rect 110 2382 12310 2438
rect 110 2372 185 2382
rect 12241 2372 12310 2382
rect 110 2256 171 2372
rect 12255 2256 12310 2372
rect 110 2246 185 2256
rect 12241 2246 12310 2256
rect 110 2192 12310 2246
rect 172 2110 232 2116
rect 596 2110 656 2116
rect 1032 2110 1092 2116
rect 2746 2110 2806 2116
rect 4466 2110 4526 2116
rect 6174 2110 6234 2116
rect 7894 2110 7954 2116
rect 9608 2110 9668 2116
rect 11326 2110 11386 2116
rect 11754 2110 11814 2116
rect 12186 2110 12246 2116
rect 172 2106 12246 2110
rect 172 2054 176 2106
rect 228 2054 600 2106
rect 652 2054 1036 2106
rect 1088 2054 2750 2106
rect 2802 2054 4470 2106
rect 4522 2054 6178 2106
rect 6230 2054 7898 2106
rect 7950 2054 9612 2106
rect 9664 2054 11330 2106
rect 11382 2054 11758 2106
rect 11810 2054 12190 2106
rect 12242 2054 12246 2106
rect 172 2050 12246 2054
rect 172 2044 232 2050
rect 596 2044 656 2050
rect 1032 2044 1092 2050
rect 2746 2044 2806 2050
rect 4466 2044 4526 2050
rect 6174 2044 6234 2050
rect 7894 2044 7954 2050
rect 9608 2044 9668 2050
rect 11326 2044 11386 2050
rect 11754 2044 11814 2050
rect 12186 2044 12246 2050
rect 1458 1982 1518 1988
rect 2312 1982 2372 1988
rect 3172 1982 3232 1988
rect 4032 1982 4092 1988
rect 4892 1982 4952 1988
rect 5752 1982 5812 1988
rect 6612 1982 6672 1988
rect 7472 1982 7532 1988
rect 8332 1982 8392 1988
rect 9172 1982 9232 1988
rect 10030 1982 10090 1988
rect 10892 1982 10952 1988
rect 1458 1978 10952 1982
rect 1458 1926 1462 1978
rect 1514 1926 2316 1978
rect 2368 1926 3176 1978
rect 3228 1926 4036 1978
rect 4088 1926 4896 1978
rect 4948 1926 5756 1978
rect 5808 1926 6616 1978
rect 6668 1926 7476 1978
rect 7528 1926 8336 1978
rect 8388 1926 9176 1978
rect 9228 1926 10034 1978
rect 10086 1926 10896 1978
rect 10948 1926 10952 1978
rect 1458 1922 10952 1926
rect 1458 1916 1518 1922
rect 2312 1916 2372 1922
rect 3172 1916 3232 1922
rect 4032 1916 4092 1922
rect 4892 1916 4952 1922
rect 5752 1916 5812 1922
rect 6612 1916 6672 1922
rect 7472 1916 7532 1922
rect 8332 1916 8392 1922
rect 9172 1916 9232 1922
rect 10030 1916 10090 1922
rect 10892 1916 10952 1922
rect -92 1846 -32 1852
rect 10468 1846 10528 1852
rect -92 1842 10528 1846
rect -92 1790 -88 1842
rect -36 1790 10472 1842
rect 10524 1790 10528 1842
rect -92 1786 10528 1790
rect -92 1780 -32 1786
rect 10468 1780 10528 1786
rect 50 1718 110 1724
rect 8752 1718 8812 1724
rect 50 1714 8812 1718
rect 50 1662 54 1714
rect 106 1662 8756 1714
rect 8808 1662 8812 1714
rect 50 1658 8812 1662
rect 50 1652 110 1658
rect 8752 1652 8812 1658
rect 1888 156 1948 162
rect 10470 156 10530 162
rect 1888 152 10530 156
rect 1888 100 1892 152
rect 1944 100 10474 152
rect 10526 100 10530 152
rect 1888 96 10530 100
rect 1888 90 1948 96
rect 10470 90 10530 96
rect 50 56 110 62
rect 3470 56 3530 62
rect 50 52 3530 56
rect 50 0 54 52
rect 106 0 3474 52
rect 3526 0 3530 52
rect 50 -4 3530 0
rect 50 -10 110 -4
rect 3470 -10 3530 -4
rect 3604 54 3664 60
rect 8756 54 8816 60
rect 3604 50 8816 54
rect 3604 -2 3608 50
rect 3660 -2 8760 50
rect 8812 -2 8816 50
rect 3604 -6 8816 -2
rect 3604 -12 3664 -6
rect 8756 -12 8816 -6
rect -92 -50 -32 -44
rect 1890 -50 1950 -44
rect -92 -54 1950 -50
rect -92 -106 -88 -54
rect -36 -106 1894 -54
rect 1946 -106 1950 -54
rect -92 -110 1950 -106
rect -92 -116 -32 -110
rect 1890 -116 1950 -110
rect 5320 -50 5380 -44
rect 7166 -50 7226 -44
rect 5320 -54 7226 -50
rect 5320 -106 5324 -54
rect 5376 -106 7170 -54
rect 7222 -106 7226 -54
rect 5320 -110 7226 -106
rect 5320 -116 5380 -110
rect 7166 -116 7226 -110
rect -92 -1580 -32 -1574
rect 10468 -1580 10528 -1574
rect -92 -1584 10528 -1580
rect -92 -1636 -88 -1584
rect -36 -1636 10472 -1584
rect 10524 -1636 10528 -1584
rect -92 -1640 10528 -1636
rect -92 -1646 -32 -1640
rect 10468 -1646 10528 -1640
rect 10904 -1684 10964 -1678
rect 1452 -1688 10964 -1684
rect 1452 -1740 1462 -1688
rect 1514 -1740 2324 -1688
rect 2376 -1740 3186 -1688
rect 3238 -1740 4044 -1688
rect 4096 -1740 4904 -1688
rect 4956 -1740 5748 -1688
rect 5800 -1740 6618 -1688
rect 6670 -1740 7484 -1688
rect 7536 -1740 8340 -1688
rect 8392 -1740 9196 -1688
rect 9248 -1740 10050 -1688
rect 10102 -1740 10908 -1688
rect 10960 -1740 10964 -1688
rect 1452 -1744 10964 -1740
rect 10904 -1750 10964 -1744
rect 50 -1786 110 -1780
rect 8752 -1786 8812 -1780
rect 50 -1790 8812 -1786
rect 50 -1842 54 -1790
rect 106 -1842 8756 -1790
rect 8808 -1842 8812 -1790
rect 50 -1846 8812 -1842
rect 50 -1852 110 -1846
rect 8752 -1852 8812 -1846
rect 6180 -3196 6240 -3187
rect 6174 -3198 6246 -3196
rect 6174 -3254 6182 -3198
rect 6238 -3254 6246 -3198
rect 6174 -3256 6246 -3254
rect 6180 -3265 6240 -3256
rect 1888 -3324 1948 -3318
rect 10470 -3324 10530 -3318
rect 1888 -3328 10530 -3324
rect 1888 -3380 1892 -3328
rect 1944 -3380 10474 -3328
rect 10526 -3380 10530 -3328
rect 1888 -3384 10530 -3380
rect 1888 -3390 1948 -3384
rect 10470 -3390 10530 -3384
rect 50 -3424 110 -3418
rect 3470 -3424 3530 -3418
rect 50 -3428 3530 -3424
rect 50 -3480 54 -3428
rect 106 -3480 3474 -3428
rect 3526 -3480 3530 -3428
rect 50 -3484 3530 -3480
rect 50 -3490 110 -3484
rect 3470 -3490 3530 -3484
rect 3604 -3426 3664 -3420
rect 8756 -3426 8816 -3420
rect 3604 -3430 8816 -3426
rect 3604 -3482 3608 -3430
rect 3660 -3482 8760 -3430
rect 8812 -3482 8816 -3430
rect 3604 -3486 8816 -3482
rect 3604 -3492 3664 -3486
rect 8756 -3492 8816 -3486
rect -92 -3530 -32 -3524
rect 1890 -3530 1950 -3524
rect -92 -3534 1950 -3530
rect 4462 -3532 4522 -3523
rect 5320 -3530 5380 -3524
rect 7166 -3530 7226 -3524
rect 7894 -3530 7954 -3521
rect -92 -3586 -88 -3534
rect -36 -3586 1894 -3534
rect 1946 -3586 1950 -3534
rect -92 -3590 1950 -3586
rect -92 -3596 -32 -3590
rect 1890 -3596 1950 -3590
rect 4456 -3534 4528 -3532
rect 4456 -3590 4464 -3534
rect 4520 -3590 4528 -3534
rect 4456 -3592 4528 -3590
rect 5320 -3534 7226 -3530
rect 5320 -3586 5324 -3534
rect 5376 -3586 7170 -3534
rect 7222 -3586 7226 -3534
rect 5320 -3590 7226 -3586
rect 7888 -3532 7960 -3530
rect 7888 -3588 7896 -3532
rect 7952 -3588 7960 -3532
rect 7888 -3590 7960 -3588
rect 4462 -3601 4522 -3592
rect 5320 -3596 5380 -3590
rect 7166 -3596 7226 -3590
rect 7894 -3599 7954 -3590
rect 1460 -5050 1520 -5044
rect 1460 -5054 10972 -5050
rect 1460 -5106 1464 -5054
rect 1516 -5106 2324 -5054
rect 2376 -5106 3180 -5054
rect 3232 -5106 4046 -5054
rect 4098 -5106 4902 -5054
rect 4954 -5106 5750 -5054
rect 5802 -5106 6604 -5054
rect 6656 -5106 7484 -5054
rect 7536 -5106 8338 -5054
rect 8390 -5058 10052 -5054
rect 8390 -5106 9196 -5058
rect 1460 -5110 9196 -5106
rect 9248 -5106 10052 -5058
rect 10104 -5106 10910 -5054
rect 10962 -5106 10972 -5054
rect 9248 -5110 10972 -5106
rect 1460 -5116 1520 -5110
rect 9186 -5114 9258 -5110
rect 3606 -5154 3666 -5148
rect 8752 -5154 8812 -5148
rect 3606 -5158 8812 -5154
rect 3606 -5210 3610 -5158
rect 3662 -5210 8756 -5158
rect 8808 -5210 8812 -5158
rect 3606 -5214 8812 -5210
rect 3606 -5220 3666 -5214
rect 8752 -5220 8812 -5214
rect 1888 -5268 1948 -5262
rect 10470 -5268 10530 -5262
rect 1888 -5272 10530 -5268
rect 1888 -5324 1892 -5272
rect 1944 -5324 10474 -5272
rect 10526 -5324 10530 -5272
rect 1888 -5328 10530 -5324
rect 1888 -5334 1948 -5328
rect 10470 -5334 10530 -5328
rect 5320 -6800 5380 -6794
rect 7038 -6800 7098 -6794
rect 5320 -6804 7098 -6800
rect 5320 -6856 5324 -6804
rect 5376 -6856 7042 -6804
rect 7094 -6856 7098 -6804
rect 5320 -6860 7098 -6856
rect 5320 -6866 5380 -6860
rect 7038 -6866 7098 -6860
rect 1456 -6926 1516 -6920
rect 2326 -6926 2386 -6920
rect 3184 -6926 3244 -6920
rect 4042 -6926 4102 -6920
rect 4900 -6926 4960 -6920
rect 5758 -6926 5818 -6920
rect 6616 -6926 6676 -6920
rect 7474 -6926 7534 -6920
rect 8332 -6926 8392 -6920
rect 9190 -6926 9250 -6920
rect 10048 -6926 10108 -6920
rect 10904 -6926 10964 -6920
rect 1456 -6930 10964 -6926
rect 1456 -6982 1460 -6930
rect 1512 -6982 2330 -6930
rect 2382 -6982 3188 -6930
rect 3240 -6982 4046 -6930
rect 4098 -6982 4904 -6930
rect 4956 -6982 5762 -6930
rect 5814 -6982 6620 -6930
rect 6672 -6982 7478 -6930
rect 7530 -6982 8336 -6930
rect 8388 -6982 9194 -6930
rect 9246 -6982 10052 -6930
rect 10104 -6982 10908 -6930
rect 10960 -6982 10964 -6930
rect 1456 -6986 10964 -6982
rect 1456 -6992 1516 -6986
rect 2326 -6992 2386 -6986
rect 3184 -6992 3244 -6986
rect 4042 -6992 4102 -6986
rect 4900 -6992 4960 -6986
rect 5758 -6992 5818 -6986
rect 6616 -6992 6676 -6986
rect 7474 -6992 7534 -6986
rect 8332 -6992 8392 -6986
rect 9190 -6992 9250 -6986
rect 10048 -6992 10108 -6986
rect 10904 -6992 10964 -6986
rect 170 -7070 230 -7064
rect 590 -7070 650 -7064
rect 1030 -7070 1090 -7064
rect 2748 -7070 2808 -7064
rect 4462 -7070 4522 -7064
rect 6180 -7070 6240 -7064
rect 7894 -7070 7954 -7064
rect 9608 -7070 9668 -7064
rect 11324 -7070 11384 -7064
rect 11750 -7070 11810 -7064
rect 12184 -7070 12244 -7064
rect 170 -7074 12244 -7070
rect 170 -7126 174 -7074
rect 226 -7126 594 -7074
rect 646 -7126 1034 -7074
rect 1086 -7126 2752 -7074
rect 2804 -7126 4466 -7074
rect 4518 -7126 6184 -7074
rect 6236 -7126 7898 -7074
rect 7950 -7126 9612 -7074
rect 9664 -7126 11328 -7074
rect 11380 -7126 11754 -7074
rect 11806 -7126 12188 -7074
rect 12240 -7126 12244 -7074
rect 170 -7130 12244 -7126
rect 170 -7136 230 -7130
rect 590 -7136 650 -7130
rect 1030 -7136 1090 -7130
rect 2748 -7136 2808 -7130
rect 4462 -7136 4522 -7130
rect 6180 -7136 6240 -7130
rect 7894 -7136 7954 -7130
rect 9608 -7136 9668 -7130
rect 11324 -7136 11384 -7130
rect 11750 -7136 11810 -7130
rect 12184 -7136 12244 -7130
rect 4798 -8162 4858 -8156
rect 6270 -8162 6330 -8156
rect 4798 -8166 6330 -8162
rect 4798 -8218 4802 -8166
rect 4854 -8218 6274 -8166
rect 6326 -8218 6330 -8166
rect 4798 -8222 6330 -8218
rect 4798 -8228 4858 -8222
rect 6270 -8228 6330 -8222
rect 5582 -8270 5642 -8264
rect 6042 -8270 6102 -8264
rect 6504 -8270 6564 -8264
rect 6960 -8270 7020 -8264
rect 5582 -8274 7020 -8270
rect 5582 -8326 5586 -8274
rect 5638 -8326 6046 -8274
rect 6098 -8326 6508 -8274
rect 6560 -8326 6964 -8274
rect 7016 -8326 7020 -8274
rect 5582 -8330 7020 -8326
rect 5582 -8336 5642 -8330
rect 6042 -8336 6102 -8330
rect 6504 -8336 6564 -8330
rect 6960 -8336 7020 -8330
rect 5356 -8978 5416 -8972
rect 6270 -8978 6330 -8972
rect 7186 -8978 7246 -8972
rect 5356 -8982 7246 -8978
rect 5356 -9034 5360 -8982
rect 5412 -9034 6274 -8982
rect 6326 -9034 7190 -8982
rect 7242 -9034 7246 -8982
rect 5356 -9038 7246 -9034
rect 5356 -9044 5416 -9038
rect 6270 -9044 6330 -9038
rect 7186 -9044 7246 -9038
rect 4798 -9092 4858 -9086
rect 5356 -9092 5416 -9086
rect 7186 -9092 7246 -9086
rect 4798 -9096 7246 -9092
rect 4798 -9148 4802 -9096
rect 4854 -9148 5360 -9096
rect 5412 -9148 7190 -9096
rect 7242 -9148 7246 -9096
rect 4798 -9152 7246 -9148
rect 4798 -9158 4858 -9152
rect 5356 -9158 5416 -9152
rect 7186 -9158 7246 -9152
rect 5584 -9792 5644 -9786
rect 6044 -9792 6104 -9786
rect 6504 -9792 6564 -9786
rect 6958 -9792 7018 -9786
rect 5584 -9796 7018 -9792
rect 5584 -9848 5588 -9796
rect 5640 -9848 6048 -9796
rect 6100 -9848 6508 -9796
rect 6560 -9848 6962 -9796
rect 7014 -9848 7018 -9796
rect 5584 -9852 7018 -9848
rect 5584 -9858 5644 -9852
rect 6044 -9858 6104 -9852
rect 6504 -9858 6564 -9852
rect 6958 -9858 7018 -9852
rect 5814 -9918 5874 -9912
rect 6728 -9918 6788 -9912
rect 5814 -9922 6788 -9918
rect 5814 -9974 5818 -9922
rect 5870 -9974 6732 -9922
rect 6784 -9974 6788 -9922
rect 5814 -9978 6788 -9974
rect 5814 -9984 5874 -9978
rect 6728 -9984 6788 -9978
rect 4664 -10193 7854 -10100
rect 4664 -10195 4758 -10193
rect 7774 -10195 7854 -10193
rect -256 -10418 344 -10406
rect -256 -10444 -224 -10418
rect 312 -10444 344 -10418
rect -256 -10688 -238 -10444
rect 326 -10688 344 -10444
rect 4664 -10567 4736 -10195
rect 7796 -10567 7854 -10195
rect 4664 -10569 4758 -10567
rect 7774 -10569 7854 -10567
rect 4664 -10646 7854 -10569
rect 11916 -10418 12516 -10406
rect 11916 -10444 11948 -10418
rect 12484 -10444 12516 -10418
rect -256 -10714 -224 -10688
rect 312 -10714 344 -10688
rect -256 -10726 344 -10714
rect 11916 -10688 11934 -10444
rect 12498 -10688 12516 -10444
rect 11916 -10714 11948 -10688
rect 12484 -10714 12516 -10688
rect 11916 -10726 12516 -10714
<< via2 >>
rect -224 2788 312 2814
rect -224 2544 312 2788
rect -224 2518 312 2544
rect 11948 2788 12484 2814
rect 11948 2544 12484 2788
rect 11948 2518 12484 2544
rect 185 2372 12241 2382
rect 185 2256 12241 2372
rect 185 2246 12241 2256
rect 6182 -3200 6238 -3198
rect 6182 -3252 6184 -3200
rect 6184 -3252 6236 -3200
rect 6236 -3252 6238 -3200
rect 6182 -3254 6238 -3252
rect 4464 -3536 4520 -3534
rect 4464 -3588 4466 -3536
rect 4466 -3588 4518 -3536
rect 4518 -3588 4520 -3536
rect 4464 -3590 4520 -3588
rect 7896 -3534 7952 -3532
rect 7896 -3586 7898 -3534
rect 7898 -3586 7950 -3534
rect 7950 -3586 7952 -3534
rect 7896 -3588 7952 -3586
rect 4758 -10195 7774 -10193
rect -224 -10444 312 -10418
rect -224 -10688 312 -10444
rect 4758 -10567 7774 -10195
rect 4758 -10569 7774 -10567
rect 11948 -10444 12484 -10418
rect -224 -10714 312 -10688
rect 11948 -10688 12484 -10444
rect 11948 -10714 12484 -10688
<< metal3 >>
rect -266 2814 354 2821
rect -266 2778 -224 2814
rect 312 2778 354 2814
rect -266 2554 -228 2778
rect 316 2554 354 2778
rect -266 2518 -224 2554
rect 312 2518 354 2554
rect -266 2511 354 2518
rect 11906 2814 12526 2821
rect 11906 2778 11948 2814
rect 12484 2778 12526 2814
rect 11906 2554 11944 2778
rect 12488 2554 12526 2778
rect 11906 2518 11948 2554
rect 12484 2518 12526 2554
rect 11906 2511 12526 2518
rect 110 2386 12310 2438
rect 110 2242 181 2386
rect 12245 2242 12310 2386
rect 110 2192 12310 2242
rect 6158 -3198 6258 -3176
rect 6158 -3254 6182 -3198
rect 6238 -3254 6258 -3198
rect 6158 -3512 6258 -3254
rect 4434 -3532 7988 -3512
rect 4434 -3534 7896 -3532
rect 4434 -3590 4464 -3534
rect 4520 -3588 7896 -3534
rect 7952 -3588 7988 -3532
rect 4520 -3590 7988 -3588
rect 4434 -3612 7988 -3590
rect 4664 -10189 7854 -10100
rect -266 -10418 354 -10411
rect -266 -10454 -224 -10418
rect 312 -10454 354 -10418
rect -266 -10678 -228 -10454
rect 316 -10678 354 -10454
rect 4664 -10573 4754 -10189
rect 7778 -10573 7854 -10189
rect 4664 -10646 7854 -10573
rect 11906 -10418 12526 -10411
rect 11906 -10454 11948 -10418
rect 12484 -10454 12526 -10418
rect -266 -10714 -224 -10678
rect 312 -10714 354 -10678
rect -266 -10721 354 -10714
rect 11906 -10678 11944 -10454
rect 12488 -10678 12526 -10454
rect 11906 -10714 11948 -10678
rect 12484 -10714 12526 -10678
rect 11906 -10721 12526 -10714
<< via3 >>
rect -228 2554 -224 2778
rect -224 2554 312 2778
rect 312 2554 316 2778
rect 11944 2554 11948 2778
rect 11948 2554 12484 2778
rect 12484 2554 12488 2778
rect 181 2382 12245 2386
rect 181 2246 185 2382
rect 185 2246 12241 2382
rect 12241 2246 12245 2382
rect 181 2242 12245 2246
rect -228 -10678 -224 -10454
rect -224 -10678 312 -10454
rect 312 -10678 316 -10454
rect 4754 -10193 7778 -10189
rect 4754 -10569 4758 -10193
rect 4758 -10569 7774 -10193
rect 7774 -10569 7778 -10193
rect 4754 -10573 7778 -10569
rect 11944 -10678 11948 -10454
rect 11948 -10678 12484 -10454
rect 12484 -10678 12488 -10454
<< metal4 >>
rect -440 2778 12700 3000
rect -440 2554 -228 2778
rect 316 2554 11944 2778
rect 12488 2554 12700 2778
rect -440 2386 12700 2554
rect -440 2242 181 2386
rect 12245 2242 12700 2386
rect -440 2200 12700 2242
rect -440 -10189 12700 -10100
rect -440 -10454 4754 -10189
rect -440 -10678 -228 -10454
rect 316 -10573 4754 -10454
rect 7778 -10454 12700 -10189
rect 7778 -10573 11944 -10454
rect 316 -10678 11944 -10573
rect 12488 -10678 12700 -10454
rect -440 -10900 12700 -10678
use ntap  ntap_69
timestamp 1626065694
transform 1 0 266 0 1 -5512
box 250 218 480 436
use ntap  ntap_68
timestamp 1626065694
transform 1 0 1124 0 1 -5512
box 250 218 480 436
use ntap  ntap_67
timestamp 1626065694
transform 1 0 1982 0 1 -5512
box 250 218 480 436
use ntap  ntap_66
timestamp 1626065694
transform 1 0 2840 0 1 -5512
box 250 218 480 436
use ntap  ntap_65
timestamp 1626065694
transform 1 0 3698 0 1 -5512
box 250 218 480 436
use ntap  ntap_64
timestamp 1626065694
transform 1 0 4556 0 1 -5512
box 250 218 480 436
use ntap  ntap_63
timestamp 1626065694
transform 1 0 5414 0 1 -5512
box 250 218 480 436
use ntap  ntap_62
timestamp 1626065694
transform 1 0 6272 0 1 -5512
box 250 218 480 436
use ntap  ntap_61
timestamp 1626065694
transform 1 0 7130 0 1 -5512
box 250 218 480 436
use ntap  ntap_60
timestamp 1626065694
transform 1 0 7988 0 1 -5512
box 250 218 480 436
use ntap  ntap_59
timestamp 1626065694
transform 1 0 8846 0 1 -5512
box 250 218 480 436
use ntap  ntap_58
timestamp 1626065694
transform 1 0 9704 0 1 -5512
box 250 218 480 436
use ntap  ntap_57
timestamp 1626065694
transform 1 0 10562 0 1 -5512
box 250 218 480 436
use ntap  ntap_56
timestamp 1626065694
transform 1 0 11420 0 1 -5512
box 250 218 480 436
use ntap  ntap_55
timestamp 1626065694
transform 1 0 278 0 1 -3768
box 250 218 480 436
use ntap  ntap_54
timestamp 1626065694
transform 1 0 1136 0 1 -3768
box 250 218 480 436
use ntap  ntap_53
timestamp 1626065694
transform 1 0 1994 0 1 -3768
box 250 218 480 436
use ntap  ntap_52
timestamp 1626065694
transform 1 0 2852 0 1 -3768
box 250 218 480 436
use ntap  ntap_51
timestamp 1626065694
transform 1 0 3710 0 1 -3768
box 250 218 480 436
use ntap  ntap_50
timestamp 1626065694
transform 1 0 4568 0 1 -3768
box 250 218 480 436
use ntap  ntap_49
timestamp 1626065694
transform 1 0 5426 0 1 -3768
box 250 218 480 436
use ntap  ntap_48
timestamp 1626065694
transform 1 0 6284 0 1 -3768
box 250 218 480 436
use ntap  ntap_47
timestamp 1626065694
transform 1 0 7142 0 1 -3768
box 250 218 480 436
use ntap  ntap_46
timestamp 1626065694
transform 1 0 8000 0 1 -3768
box 250 218 480 436
use ntap  ntap_45
timestamp 1626065694
transform 1 0 8858 0 1 -3768
box 250 218 480 436
use ntap  ntap_44
timestamp 1626065694
transform 1 0 9716 0 1 -3768
box 250 218 480 436
use ntap  ntap_43
timestamp 1626065694
transform 1 0 10574 0 1 -3768
box 250 218 480 436
use ntap  ntap_42
timestamp 1626065694
transform 1 0 11432 0 1 -3768
box 250 218 480 436
use ntap  ntap_41
timestamp 1626065694
transform 1 0 278 0 1 -2032
box 250 218 480 436
use ntap  ntap_40
timestamp 1626065694
transform 1 0 1136 0 1 -2032
box 250 218 480 436
use ntap  ntap_39
timestamp 1626065694
transform 1 0 1994 0 1 -2032
box 250 218 480 436
use ntap  ntap_38
timestamp 1626065694
transform 1 0 2852 0 1 -2032
box 250 218 480 436
use ntap  ntap_37
timestamp 1626065694
transform 1 0 3710 0 1 -2032
box 250 218 480 436
use ntap  ntap_36
timestamp 1626065694
transform 1 0 4568 0 1 -2032
box 250 218 480 436
use ntap  ntap_35
timestamp 1626065694
transform 1 0 5426 0 1 -2032
box 250 218 480 436
use ntap  ntap_34
timestamp 1626065694
transform 1 0 6284 0 1 -2032
box 250 218 480 436
use ntap  ntap_33
timestamp 1626065694
transform 1 0 7142 0 1 -2032
box 250 218 480 436
use ntap  ntap_32
timestamp 1626065694
transform 1 0 8000 0 1 -2032
box 250 218 480 436
use ntap  ntap_31
timestamp 1626065694
transform 1 0 8858 0 1 -2032
box 250 218 480 436
use ntap  ntap_30
timestamp 1626065694
transform 1 0 9716 0 1 -2032
box 250 218 480 436
use ntap  ntap_29
timestamp 1626065694
transform 1 0 10574 0 1 -2032
box 250 218 480 436
use ntap  ntap_28
timestamp 1626065694
transform 1 0 11432 0 1 -2032
box 250 218 480 436
use ntap  ntap_27
timestamp 1626065694
transform 1 0 282 0 1 -290
box 250 218 480 436
use ntap  ntap_26
timestamp 1626065694
transform 1 0 1140 0 1 -290
box 250 218 480 436
use ntap  ntap_25
timestamp 1626065694
transform 1 0 1998 0 1 -290
box 250 218 480 436
use ntap  ntap_24
timestamp 1626065694
transform 1 0 2856 0 1 -290
box 250 218 480 436
use ntap  ntap_23
timestamp 1626065694
transform 1 0 3714 0 1 -290
box 250 218 480 436
use ntap  ntap_22
timestamp 1626065694
transform 1 0 4572 0 1 -290
box 250 218 480 436
use ntap  ntap_21
timestamp 1626065694
transform 1 0 5430 0 1 -290
box 250 218 480 436
use ntap  ntap_20
timestamp 1626065694
transform 1 0 6288 0 1 -290
box 250 218 480 436
use ntap  ntap_19
timestamp 1626065694
transform 1 0 7146 0 1 -290
box 250 218 480 436
use ntap  ntap_18
timestamp 1626065694
transform 1 0 8004 0 1 -290
box 250 218 480 436
use ntap  ntap_17
timestamp 1626065694
transform 1 0 8862 0 1 -290
box 250 218 480 436
use ntap  ntap_16
timestamp 1626065694
transform 1 0 9720 0 1 -290
box 250 218 480 436
use ntap  ntap_15
timestamp 1626065694
transform 1 0 10578 0 1 -290
box 250 218 480 436
use ntap  ntap_14
timestamp 1626065694
transform 1 0 11436 0 1 -290
box 250 218 480 436
use ntap  ntap_13
timestamp 1626065694
transform 1 0 266 0 1 1474
box 250 218 480 436
use ntap  ntap_12
timestamp 1626065694
transform 1 0 1124 0 1 1474
box 250 218 480 436
use ntap  ntap_11
timestamp 1626065694
transform 1 0 1982 0 1 1474
box 250 218 480 436
use ntap  ntap_10
timestamp 1626065694
transform 1 0 2840 0 1 1474
box 250 218 480 436
use ntap  ntap_9
timestamp 1626065694
transform 1 0 3698 0 1 1474
box 250 218 480 436
use ntap  ntap_8
timestamp 1626065694
transform 1 0 4556 0 1 1474
box 250 218 480 436
use ntap  ntap_7
timestamp 1626065694
transform 1 0 5414 0 1 1474
box 250 218 480 436
use ntap  ntap_6
timestamp 1626065694
transform 1 0 6272 0 1 1474
box 250 218 480 436
use ntap  ntap_5
timestamp 1626065694
transform 1 0 7130 0 1 1474
box 250 218 480 436
use ntap  ntap_4
timestamp 1626065694
transform 1 0 7988 0 1 1474
box 250 218 480 436
use ntap  ntap_3
timestamp 1626065694
transform 1 0 8846 0 1 1474
box 250 218 480 436
use ntap  ntap_2
timestamp 1626065694
transform 1 0 9704 0 1 1474
box 250 218 480 436
use ntap  ntap_1
timestamp 1626065694
transform 1 0 10562 0 1 1474
box 250 218 480 436
use ntap  ntap_0
timestamp 1626065694
transform 1 0 11420 0 1 1474
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_8WETQ2  sky130_fd_pr__pfet_01v8_8WETQ2_4
timestamp 1626065694
transform 1 0 6209 0 1 -6056
box -6071 -700 6071 700
use sky130_fd_pr__pfet_01v8_8WETQ2  sky130_fd_pr__pfet_01v8_8WETQ2_3
timestamp 1626065694
transform 1 0 6209 0 1 -4316
box -6071 -700 6071 700
use sky130_fd_pr__pfet_01v8_8WETQ2  sky130_fd_pr__pfet_01v8_8WETQ2_2
timestamp 1626065694
transform 1 0 6209 0 1 -2576
box -6071 -700 6071 700
use sky130_fd_pr__pfet_01v8_8WETQ2  sky130_fd_pr__pfet_01v8_8WETQ2_1
timestamp 1626065694
transform 1 0 6209 0 1 -836
box -6071 -700 6071 700
use sky130_fd_pr__pfet_01v8_8WETQ2  sky130_fd_pr__pfet_01v8_8WETQ2_0
timestamp 1626065694
transform 1 0 6209 0 1 904
box -6071 -700 6071 700
use sky130_fd_pr__nfet_01v8_C5Q2Z6  sky130_fd_pr__nfet_01v8_C5Q2Z6_1
timestamp 1626065694
transform 1 0 6301 0 1 -8660
box -1429 -288 1429 288
use sky130_fd_pr__nfet_01v8_C5Q2Z6  sky130_fd_pr__nfet_01v8_C5Q2Z6_0
timestamp 1626065694
transform 1 0 6301 0 1 -9460
box -1429 -288 1429 288
<< labels >>
flabel metal2 s 2170 120 2190 138 1 FreeSans 600 0 0 0 low_freq_pll_ibiasn
flabel metal2 s 1436 -74 1454 -64 1 FreeSans 600 0 0 0 comparator_ibiasn
flabel metal2 s 3796 12 3814 26 1 FreeSans 600 0 0 0 biquad_gm_c_filter_ibiasn4
flabel metal1 s 5340 180 5354 186 1 FreeSans 600 0 0 0 biquad_gm_c_filter_ibiasn3
flabel metal2 s 5890 -90 5904 -74 1 FreeSans 600 0 0 0 biquad_gm_c_filter_ibiasn2
flabel metal2 s 2212 16 2228 34 1 FreeSans 600 0 0 0 biquad_gm_c_filter_ibiasn1
flabel metal2 s 1210 -3580 1234 -3554 1 FreeSans 600 0 0 0 sample_and_hold_ibiasn_A
flabel metal2 s 1524 -3460 1542 -3444 1 FreeSans 600 0 0 0 peak_detector_ibiasn2
flabel metal2 s 6342 -3576 6354 -3558 1 FreeSans 600 0 0 0 peak_detector_ibiasn1
flabel metal1 s 5342 -3304 5356 -3294 1 FreeSans 600 0 0 0 diff_to_se_converter_ibiasn
flabel metal2 s 3948 -3460 3954 -3444 1 FreeSans 600 0 0 0 input_amplifier_ibiasn2
flabel metal2 s 3240 -3356 3256 -3342 1 FreeSans 600 0 0 0 input_amplifier_ibiasn1
flabel metal2 s 6058 -6832 6082 -6816 1 FreeSans 600 0 0 0 dac_8bit_ibiasn_B
flabel metal2 s 4048 -5194 4060 -5174 1 FreeSans 600 0 0 0 sample_and_hold_ibiasn_B
flabel metal2 s 2324 -5298 2344 -5282 1 FreeSans 600 0 0 0 dac_8bit_ibiasn_A
flabel metal2 s 3562 -6966 3574 -6948 1 FreeSans 600 0 0 0 vbiasp
flabel metal4 s -414 2968 -398 2984 1 FreeSans 600 0 0 0 VDD
flabel metal2 s 6620 -9826 6626 -9814 1 FreeSans 600 0 0 0 vbiasn
flabel metal2 s 5934 -9020 5950 -9006 1 FreeSans 600 0 0 0 dac_8bit_ibiasp_A
flabel metal2 s 5264 -9132 5274 -9118 1 FreeSans 600 0 0 0 dac_8bit_ibiasp_B
flabel metal4 s -398 -10890 -382 -10872 1 FreeSans 600 0 0 0 VSS
<< properties >>
string FIXED_BBOX -312 -11172 12572 -8028
<< end >>
