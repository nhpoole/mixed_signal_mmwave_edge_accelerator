magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -8960 -1660 8960 1660
<< nwell >>
rect -7700 -400 7700 400
<< pmos >>
rect -7606 -300 -6646 300
rect -6588 -300 -5628 300
rect -5570 -300 -4610 300
rect -4552 -300 -3592 300
rect -3534 -300 -2574 300
rect -2516 -300 -1556 300
rect -1498 -300 -538 300
rect -480 -300 480 300
rect 538 -300 1498 300
rect 1556 -300 2516 300
rect 2574 -300 3534 300
rect 3592 -300 4552 300
rect 4610 -300 5570 300
rect 5628 -300 6588 300
rect 6646 -300 7606 300
<< pdiff >>
rect -7664 255 -7606 300
rect -7664 221 -7652 255
rect -7618 221 -7606 255
rect -7664 187 -7606 221
rect -7664 153 -7652 187
rect -7618 153 -7606 187
rect -7664 119 -7606 153
rect -7664 85 -7652 119
rect -7618 85 -7606 119
rect -7664 51 -7606 85
rect -7664 17 -7652 51
rect -7618 17 -7606 51
rect -7664 -17 -7606 17
rect -7664 -51 -7652 -17
rect -7618 -51 -7606 -17
rect -7664 -85 -7606 -51
rect -7664 -119 -7652 -85
rect -7618 -119 -7606 -85
rect -7664 -153 -7606 -119
rect -7664 -187 -7652 -153
rect -7618 -187 -7606 -153
rect -7664 -221 -7606 -187
rect -7664 -255 -7652 -221
rect -7618 -255 -7606 -221
rect -7664 -300 -7606 -255
rect -6646 255 -6588 300
rect -6646 221 -6634 255
rect -6600 221 -6588 255
rect -6646 187 -6588 221
rect -6646 153 -6634 187
rect -6600 153 -6588 187
rect -6646 119 -6588 153
rect -6646 85 -6634 119
rect -6600 85 -6588 119
rect -6646 51 -6588 85
rect -6646 17 -6634 51
rect -6600 17 -6588 51
rect -6646 -17 -6588 17
rect -6646 -51 -6634 -17
rect -6600 -51 -6588 -17
rect -6646 -85 -6588 -51
rect -6646 -119 -6634 -85
rect -6600 -119 -6588 -85
rect -6646 -153 -6588 -119
rect -6646 -187 -6634 -153
rect -6600 -187 -6588 -153
rect -6646 -221 -6588 -187
rect -6646 -255 -6634 -221
rect -6600 -255 -6588 -221
rect -6646 -300 -6588 -255
rect -5628 255 -5570 300
rect -5628 221 -5616 255
rect -5582 221 -5570 255
rect -5628 187 -5570 221
rect -5628 153 -5616 187
rect -5582 153 -5570 187
rect -5628 119 -5570 153
rect -5628 85 -5616 119
rect -5582 85 -5570 119
rect -5628 51 -5570 85
rect -5628 17 -5616 51
rect -5582 17 -5570 51
rect -5628 -17 -5570 17
rect -5628 -51 -5616 -17
rect -5582 -51 -5570 -17
rect -5628 -85 -5570 -51
rect -5628 -119 -5616 -85
rect -5582 -119 -5570 -85
rect -5628 -153 -5570 -119
rect -5628 -187 -5616 -153
rect -5582 -187 -5570 -153
rect -5628 -221 -5570 -187
rect -5628 -255 -5616 -221
rect -5582 -255 -5570 -221
rect -5628 -300 -5570 -255
rect -4610 255 -4552 300
rect -4610 221 -4598 255
rect -4564 221 -4552 255
rect -4610 187 -4552 221
rect -4610 153 -4598 187
rect -4564 153 -4552 187
rect -4610 119 -4552 153
rect -4610 85 -4598 119
rect -4564 85 -4552 119
rect -4610 51 -4552 85
rect -4610 17 -4598 51
rect -4564 17 -4552 51
rect -4610 -17 -4552 17
rect -4610 -51 -4598 -17
rect -4564 -51 -4552 -17
rect -4610 -85 -4552 -51
rect -4610 -119 -4598 -85
rect -4564 -119 -4552 -85
rect -4610 -153 -4552 -119
rect -4610 -187 -4598 -153
rect -4564 -187 -4552 -153
rect -4610 -221 -4552 -187
rect -4610 -255 -4598 -221
rect -4564 -255 -4552 -221
rect -4610 -300 -4552 -255
rect -3592 255 -3534 300
rect -3592 221 -3580 255
rect -3546 221 -3534 255
rect -3592 187 -3534 221
rect -3592 153 -3580 187
rect -3546 153 -3534 187
rect -3592 119 -3534 153
rect -3592 85 -3580 119
rect -3546 85 -3534 119
rect -3592 51 -3534 85
rect -3592 17 -3580 51
rect -3546 17 -3534 51
rect -3592 -17 -3534 17
rect -3592 -51 -3580 -17
rect -3546 -51 -3534 -17
rect -3592 -85 -3534 -51
rect -3592 -119 -3580 -85
rect -3546 -119 -3534 -85
rect -3592 -153 -3534 -119
rect -3592 -187 -3580 -153
rect -3546 -187 -3534 -153
rect -3592 -221 -3534 -187
rect -3592 -255 -3580 -221
rect -3546 -255 -3534 -221
rect -3592 -300 -3534 -255
rect -2574 255 -2516 300
rect -2574 221 -2562 255
rect -2528 221 -2516 255
rect -2574 187 -2516 221
rect -2574 153 -2562 187
rect -2528 153 -2516 187
rect -2574 119 -2516 153
rect -2574 85 -2562 119
rect -2528 85 -2516 119
rect -2574 51 -2516 85
rect -2574 17 -2562 51
rect -2528 17 -2516 51
rect -2574 -17 -2516 17
rect -2574 -51 -2562 -17
rect -2528 -51 -2516 -17
rect -2574 -85 -2516 -51
rect -2574 -119 -2562 -85
rect -2528 -119 -2516 -85
rect -2574 -153 -2516 -119
rect -2574 -187 -2562 -153
rect -2528 -187 -2516 -153
rect -2574 -221 -2516 -187
rect -2574 -255 -2562 -221
rect -2528 -255 -2516 -221
rect -2574 -300 -2516 -255
rect -1556 255 -1498 300
rect -1556 221 -1544 255
rect -1510 221 -1498 255
rect -1556 187 -1498 221
rect -1556 153 -1544 187
rect -1510 153 -1498 187
rect -1556 119 -1498 153
rect -1556 85 -1544 119
rect -1510 85 -1498 119
rect -1556 51 -1498 85
rect -1556 17 -1544 51
rect -1510 17 -1498 51
rect -1556 -17 -1498 17
rect -1556 -51 -1544 -17
rect -1510 -51 -1498 -17
rect -1556 -85 -1498 -51
rect -1556 -119 -1544 -85
rect -1510 -119 -1498 -85
rect -1556 -153 -1498 -119
rect -1556 -187 -1544 -153
rect -1510 -187 -1498 -153
rect -1556 -221 -1498 -187
rect -1556 -255 -1544 -221
rect -1510 -255 -1498 -221
rect -1556 -300 -1498 -255
rect -538 255 -480 300
rect -538 221 -526 255
rect -492 221 -480 255
rect -538 187 -480 221
rect -538 153 -526 187
rect -492 153 -480 187
rect -538 119 -480 153
rect -538 85 -526 119
rect -492 85 -480 119
rect -538 51 -480 85
rect -538 17 -526 51
rect -492 17 -480 51
rect -538 -17 -480 17
rect -538 -51 -526 -17
rect -492 -51 -480 -17
rect -538 -85 -480 -51
rect -538 -119 -526 -85
rect -492 -119 -480 -85
rect -538 -153 -480 -119
rect -538 -187 -526 -153
rect -492 -187 -480 -153
rect -538 -221 -480 -187
rect -538 -255 -526 -221
rect -492 -255 -480 -221
rect -538 -300 -480 -255
rect 480 255 538 300
rect 480 221 492 255
rect 526 221 538 255
rect 480 187 538 221
rect 480 153 492 187
rect 526 153 538 187
rect 480 119 538 153
rect 480 85 492 119
rect 526 85 538 119
rect 480 51 538 85
rect 480 17 492 51
rect 526 17 538 51
rect 480 -17 538 17
rect 480 -51 492 -17
rect 526 -51 538 -17
rect 480 -85 538 -51
rect 480 -119 492 -85
rect 526 -119 538 -85
rect 480 -153 538 -119
rect 480 -187 492 -153
rect 526 -187 538 -153
rect 480 -221 538 -187
rect 480 -255 492 -221
rect 526 -255 538 -221
rect 480 -300 538 -255
rect 1498 255 1556 300
rect 1498 221 1510 255
rect 1544 221 1556 255
rect 1498 187 1556 221
rect 1498 153 1510 187
rect 1544 153 1556 187
rect 1498 119 1556 153
rect 1498 85 1510 119
rect 1544 85 1556 119
rect 1498 51 1556 85
rect 1498 17 1510 51
rect 1544 17 1556 51
rect 1498 -17 1556 17
rect 1498 -51 1510 -17
rect 1544 -51 1556 -17
rect 1498 -85 1556 -51
rect 1498 -119 1510 -85
rect 1544 -119 1556 -85
rect 1498 -153 1556 -119
rect 1498 -187 1510 -153
rect 1544 -187 1556 -153
rect 1498 -221 1556 -187
rect 1498 -255 1510 -221
rect 1544 -255 1556 -221
rect 1498 -300 1556 -255
rect 2516 255 2574 300
rect 2516 221 2528 255
rect 2562 221 2574 255
rect 2516 187 2574 221
rect 2516 153 2528 187
rect 2562 153 2574 187
rect 2516 119 2574 153
rect 2516 85 2528 119
rect 2562 85 2574 119
rect 2516 51 2574 85
rect 2516 17 2528 51
rect 2562 17 2574 51
rect 2516 -17 2574 17
rect 2516 -51 2528 -17
rect 2562 -51 2574 -17
rect 2516 -85 2574 -51
rect 2516 -119 2528 -85
rect 2562 -119 2574 -85
rect 2516 -153 2574 -119
rect 2516 -187 2528 -153
rect 2562 -187 2574 -153
rect 2516 -221 2574 -187
rect 2516 -255 2528 -221
rect 2562 -255 2574 -221
rect 2516 -300 2574 -255
rect 3534 255 3592 300
rect 3534 221 3546 255
rect 3580 221 3592 255
rect 3534 187 3592 221
rect 3534 153 3546 187
rect 3580 153 3592 187
rect 3534 119 3592 153
rect 3534 85 3546 119
rect 3580 85 3592 119
rect 3534 51 3592 85
rect 3534 17 3546 51
rect 3580 17 3592 51
rect 3534 -17 3592 17
rect 3534 -51 3546 -17
rect 3580 -51 3592 -17
rect 3534 -85 3592 -51
rect 3534 -119 3546 -85
rect 3580 -119 3592 -85
rect 3534 -153 3592 -119
rect 3534 -187 3546 -153
rect 3580 -187 3592 -153
rect 3534 -221 3592 -187
rect 3534 -255 3546 -221
rect 3580 -255 3592 -221
rect 3534 -300 3592 -255
rect 4552 255 4610 300
rect 4552 221 4564 255
rect 4598 221 4610 255
rect 4552 187 4610 221
rect 4552 153 4564 187
rect 4598 153 4610 187
rect 4552 119 4610 153
rect 4552 85 4564 119
rect 4598 85 4610 119
rect 4552 51 4610 85
rect 4552 17 4564 51
rect 4598 17 4610 51
rect 4552 -17 4610 17
rect 4552 -51 4564 -17
rect 4598 -51 4610 -17
rect 4552 -85 4610 -51
rect 4552 -119 4564 -85
rect 4598 -119 4610 -85
rect 4552 -153 4610 -119
rect 4552 -187 4564 -153
rect 4598 -187 4610 -153
rect 4552 -221 4610 -187
rect 4552 -255 4564 -221
rect 4598 -255 4610 -221
rect 4552 -300 4610 -255
rect 5570 255 5628 300
rect 5570 221 5582 255
rect 5616 221 5628 255
rect 5570 187 5628 221
rect 5570 153 5582 187
rect 5616 153 5628 187
rect 5570 119 5628 153
rect 5570 85 5582 119
rect 5616 85 5628 119
rect 5570 51 5628 85
rect 5570 17 5582 51
rect 5616 17 5628 51
rect 5570 -17 5628 17
rect 5570 -51 5582 -17
rect 5616 -51 5628 -17
rect 5570 -85 5628 -51
rect 5570 -119 5582 -85
rect 5616 -119 5628 -85
rect 5570 -153 5628 -119
rect 5570 -187 5582 -153
rect 5616 -187 5628 -153
rect 5570 -221 5628 -187
rect 5570 -255 5582 -221
rect 5616 -255 5628 -221
rect 5570 -300 5628 -255
rect 6588 255 6646 300
rect 6588 221 6600 255
rect 6634 221 6646 255
rect 6588 187 6646 221
rect 6588 153 6600 187
rect 6634 153 6646 187
rect 6588 119 6646 153
rect 6588 85 6600 119
rect 6634 85 6646 119
rect 6588 51 6646 85
rect 6588 17 6600 51
rect 6634 17 6646 51
rect 6588 -17 6646 17
rect 6588 -51 6600 -17
rect 6634 -51 6646 -17
rect 6588 -85 6646 -51
rect 6588 -119 6600 -85
rect 6634 -119 6646 -85
rect 6588 -153 6646 -119
rect 6588 -187 6600 -153
rect 6634 -187 6646 -153
rect 6588 -221 6646 -187
rect 6588 -255 6600 -221
rect 6634 -255 6646 -221
rect 6588 -300 6646 -255
rect 7606 255 7664 300
rect 7606 221 7618 255
rect 7652 221 7664 255
rect 7606 187 7664 221
rect 7606 153 7618 187
rect 7652 153 7664 187
rect 7606 119 7664 153
rect 7606 85 7618 119
rect 7652 85 7664 119
rect 7606 51 7664 85
rect 7606 17 7618 51
rect 7652 17 7664 51
rect 7606 -17 7664 17
rect 7606 -51 7618 -17
rect 7652 -51 7664 -17
rect 7606 -85 7664 -51
rect 7606 -119 7618 -85
rect 7652 -119 7664 -85
rect 7606 -153 7664 -119
rect 7606 -187 7618 -153
rect 7652 -187 7664 -153
rect 7606 -221 7664 -187
rect 7606 -255 7618 -221
rect 7652 -255 7664 -221
rect 7606 -300 7664 -255
<< pdiffc >>
rect -7652 221 -7618 255
rect -7652 153 -7618 187
rect -7652 85 -7618 119
rect -7652 17 -7618 51
rect -7652 -51 -7618 -17
rect -7652 -119 -7618 -85
rect -7652 -187 -7618 -153
rect -7652 -255 -7618 -221
rect -6634 221 -6600 255
rect -6634 153 -6600 187
rect -6634 85 -6600 119
rect -6634 17 -6600 51
rect -6634 -51 -6600 -17
rect -6634 -119 -6600 -85
rect -6634 -187 -6600 -153
rect -6634 -255 -6600 -221
rect -5616 221 -5582 255
rect -5616 153 -5582 187
rect -5616 85 -5582 119
rect -5616 17 -5582 51
rect -5616 -51 -5582 -17
rect -5616 -119 -5582 -85
rect -5616 -187 -5582 -153
rect -5616 -255 -5582 -221
rect -4598 221 -4564 255
rect -4598 153 -4564 187
rect -4598 85 -4564 119
rect -4598 17 -4564 51
rect -4598 -51 -4564 -17
rect -4598 -119 -4564 -85
rect -4598 -187 -4564 -153
rect -4598 -255 -4564 -221
rect -3580 221 -3546 255
rect -3580 153 -3546 187
rect -3580 85 -3546 119
rect -3580 17 -3546 51
rect -3580 -51 -3546 -17
rect -3580 -119 -3546 -85
rect -3580 -187 -3546 -153
rect -3580 -255 -3546 -221
rect -2562 221 -2528 255
rect -2562 153 -2528 187
rect -2562 85 -2528 119
rect -2562 17 -2528 51
rect -2562 -51 -2528 -17
rect -2562 -119 -2528 -85
rect -2562 -187 -2528 -153
rect -2562 -255 -2528 -221
rect -1544 221 -1510 255
rect -1544 153 -1510 187
rect -1544 85 -1510 119
rect -1544 17 -1510 51
rect -1544 -51 -1510 -17
rect -1544 -119 -1510 -85
rect -1544 -187 -1510 -153
rect -1544 -255 -1510 -221
rect -526 221 -492 255
rect -526 153 -492 187
rect -526 85 -492 119
rect -526 17 -492 51
rect -526 -51 -492 -17
rect -526 -119 -492 -85
rect -526 -187 -492 -153
rect -526 -255 -492 -221
rect 492 221 526 255
rect 492 153 526 187
rect 492 85 526 119
rect 492 17 526 51
rect 492 -51 526 -17
rect 492 -119 526 -85
rect 492 -187 526 -153
rect 492 -255 526 -221
rect 1510 221 1544 255
rect 1510 153 1544 187
rect 1510 85 1544 119
rect 1510 17 1544 51
rect 1510 -51 1544 -17
rect 1510 -119 1544 -85
rect 1510 -187 1544 -153
rect 1510 -255 1544 -221
rect 2528 221 2562 255
rect 2528 153 2562 187
rect 2528 85 2562 119
rect 2528 17 2562 51
rect 2528 -51 2562 -17
rect 2528 -119 2562 -85
rect 2528 -187 2562 -153
rect 2528 -255 2562 -221
rect 3546 221 3580 255
rect 3546 153 3580 187
rect 3546 85 3580 119
rect 3546 17 3580 51
rect 3546 -51 3580 -17
rect 3546 -119 3580 -85
rect 3546 -187 3580 -153
rect 3546 -255 3580 -221
rect 4564 221 4598 255
rect 4564 153 4598 187
rect 4564 85 4598 119
rect 4564 17 4598 51
rect 4564 -51 4598 -17
rect 4564 -119 4598 -85
rect 4564 -187 4598 -153
rect 4564 -255 4598 -221
rect 5582 221 5616 255
rect 5582 153 5616 187
rect 5582 85 5616 119
rect 5582 17 5616 51
rect 5582 -51 5616 -17
rect 5582 -119 5616 -85
rect 5582 -187 5616 -153
rect 5582 -255 5616 -221
rect 6600 221 6634 255
rect 6600 153 6634 187
rect 6600 85 6634 119
rect 6600 17 6634 51
rect 6600 -51 6634 -17
rect 6600 -119 6634 -85
rect 6600 -187 6634 -153
rect 6600 -255 6634 -221
rect 7618 221 7652 255
rect 7618 153 7652 187
rect 7618 85 7652 119
rect 7618 17 7652 51
rect 7618 -51 7652 -17
rect 7618 -119 7652 -85
rect 7618 -187 7652 -153
rect 7618 -255 7652 -221
<< poly >>
rect -7420 381 -6832 397
rect -7420 364 -7381 381
rect -7606 347 -7381 364
rect -7347 347 -7313 381
rect -7279 347 -7245 381
rect -7211 347 -7177 381
rect -7143 347 -7109 381
rect -7075 347 -7041 381
rect -7007 347 -6973 381
rect -6939 347 -6905 381
rect -6871 364 -6832 381
rect -6402 381 -5814 397
rect -6402 364 -6363 381
rect -6871 347 -6646 364
rect -7606 300 -6646 347
rect -6588 347 -6363 364
rect -6329 347 -6295 381
rect -6261 347 -6227 381
rect -6193 347 -6159 381
rect -6125 347 -6091 381
rect -6057 347 -6023 381
rect -5989 347 -5955 381
rect -5921 347 -5887 381
rect -5853 364 -5814 381
rect -5384 381 -4796 397
rect -5384 364 -5345 381
rect -5853 347 -5628 364
rect -6588 300 -5628 347
rect -5570 347 -5345 364
rect -5311 347 -5277 381
rect -5243 347 -5209 381
rect -5175 347 -5141 381
rect -5107 347 -5073 381
rect -5039 347 -5005 381
rect -4971 347 -4937 381
rect -4903 347 -4869 381
rect -4835 364 -4796 381
rect -4366 381 -3778 397
rect -4366 364 -4327 381
rect -4835 347 -4610 364
rect -5570 300 -4610 347
rect -4552 347 -4327 364
rect -4293 347 -4259 381
rect -4225 347 -4191 381
rect -4157 347 -4123 381
rect -4089 347 -4055 381
rect -4021 347 -3987 381
rect -3953 347 -3919 381
rect -3885 347 -3851 381
rect -3817 364 -3778 381
rect -3348 381 -2760 397
rect -3348 364 -3309 381
rect -3817 347 -3592 364
rect -4552 300 -3592 347
rect -3534 347 -3309 364
rect -3275 347 -3241 381
rect -3207 347 -3173 381
rect -3139 347 -3105 381
rect -3071 347 -3037 381
rect -3003 347 -2969 381
rect -2935 347 -2901 381
rect -2867 347 -2833 381
rect -2799 364 -2760 381
rect -2330 381 -1742 397
rect -2330 364 -2291 381
rect -2799 347 -2574 364
rect -3534 300 -2574 347
rect -2516 347 -2291 364
rect -2257 347 -2223 381
rect -2189 347 -2155 381
rect -2121 347 -2087 381
rect -2053 347 -2019 381
rect -1985 347 -1951 381
rect -1917 347 -1883 381
rect -1849 347 -1815 381
rect -1781 364 -1742 381
rect -1312 381 -724 397
rect -1312 364 -1273 381
rect -1781 347 -1556 364
rect -2516 300 -1556 347
rect -1498 347 -1273 364
rect -1239 347 -1205 381
rect -1171 347 -1137 381
rect -1103 347 -1069 381
rect -1035 347 -1001 381
rect -967 347 -933 381
rect -899 347 -865 381
rect -831 347 -797 381
rect -763 364 -724 381
rect -294 381 294 397
rect -294 364 -255 381
rect -763 347 -538 364
rect -1498 300 -538 347
rect -480 347 -255 364
rect -221 347 -187 381
rect -153 347 -119 381
rect -85 347 -51 381
rect -17 347 17 381
rect 51 347 85 381
rect 119 347 153 381
rect 187 347 221 381
rect 255 364 294 381
rect 724 381 1312 397
rect 724 364 763 381
rect 255 347 480 364
rect -480 300 480 347
rect 538 347 763 364
rect 797 347 831 381
rect 865 347 899 381
rect 933 347 967 381
rect 1001 347 1035 381
rect 1069 347 1103 381
rect 1137 347 1171 381
rect 1205 347 1239 381
rect 1273 364 1312 381
rect 1742 381 2330 397
rect 1742 364 1781 381
rect 1273 347 1498 364
rect 538 300 1498 347
rect 1556 347 1781 364
rect 1815 347 1849 381
rect 1883 347 1917 381
rect 1951 347 1985 381
rect 2019 347 2053 381
rect 2087 347 2121 381
rect 2155 347 2189 381
rect 2223 347 2257 381
rect 2291 364 2330 381
rect 2760 381 3348 397
rect 2760 364 2799 381
rect 2291 347 2516 364
rect 1556 300 2516 347
rect 2574 347 2799 364
rect 2833 347 2867 381
rect 2901 347 2935 381
rect 2969 347 3003 381
rect 3037 347 3071 381
rect 3105 347 3139 381
rect 3173 347 3207 381
rect 3241 347 3275 381
rect 3309 364 3348 381
rect 3778 381 4366 397
rect 3778 364 3817 381
rect 3309 347 3534 364
rect 2574 300 3534 347
rect 3592 347 3817 364
rect 3851 347 3885 381
rect 3919 347 3953 381
rect 3987 347 4021 381
rect 4055 347 4089 381
rect 4123 347 4157 381
rect 4191 347 4225 381
rect 4259 347 4293 381
rect 4327 364 4366 381
rect 4796 381 5384 397
rect 4796 364 4835 381
rect 4327 347 4552 364
rect 3592 300 4552 347
rect 4610 347 4835 364
rect 4869 347 4903 381
rect 4937 347 4971 381
rect 5005 347 5039 381
rect 5073 347 5107 381
rect 5141 347 5175 381
rect 5209 347 5243 381
rect 5277 347 5311 381
rect 5345 364 5384 381
rect 5814 381 6402 397
rect 5814 364 5853 381
rect 5345 347 5570 364
rect 4610 300 5570 347
rect 5628 347 5853 364
rect 5887 347 5921 381
rect 5955 347 5989 381
rect 6023 347 6057 381
rect 6091 347 6125 381
rect 6159 347 6193 381
rect 6227 347 6261 381
rect 6295 347 6329 381
rect 6363 364 6402 381
rect 6832 381 7420 397
rect 6832 364 6871 381
rect 6363 347 6588 364
rect 5628 300 6588 347
rect 6646 347 6871 364
rect 6905 347 6939 381
rect 6973 347 7007 381
rect 7041 347 7075 381
rect 7109 347 7143 381
rect 7177 347 7211 381
rect 7245 347 7279 381
rect 7313 347 7347 381
rect 7381 364 7420 381
rect 7381 347 7606 364
rect 6646 300 7606 347
rect -7606 -347 -6646 -300
rect -7606 -364 -7381 -347
rect -7420 -381 -7381 -364
rect -7347 -381 -7313 -347
rect -7279 -381 -7245 -347
rect -7211 -381 -7177 -347
rect -7143 -381 -7109 -347
rect -7075 -381 -7041 -347
rect -7007 -381 -6973 -347
rect -6939 -381 -6905 -347
rect -6871 -364 -6646 -347
rect -6588 -347 -5628 -300
rect -6588 -364 -6363 -347
rect -6871 -381 -6832 -364
rect -7420 -397 -6832 -381
rect -6402 -381 -6363 -364
rect -6329 -381 -6295 -347
rect -6261 -381 -6227 -347
rect -6193 -381 -6159 -347
rect -6125 -381 -6091 -347
rect -6057 -381 -6023 -347
rect -5989 -381 -5955 -347
rect -5921 -381 -5887 -347
rect -5853 -364 -5628 -347
rect -5570 -347 -4610 -300
rect -5570 -364 -5345 -347
rect -5853 -381 -5814 -364
rect -6402 -397 -5814 -381
rect -5384 -381 -5345 -364
rect -5311 -381 -5277 -347
rect -5243 -381 -5209 -347
rect -5175 -381 -5141 -347
rect -5107 -381 -5073 -347
rect -5039 -381 -5005 -347
rect -4971 -381 -4937 -347
rect -4903 -381 -4869 -347
rect -4835 -364 -4610 -347
rect -4552 -347 -3592 -300
rect -4552 -364 -4327 -347
rect -4835 -381 -4796 -364
rect -5384 -397 -4796 -381
rect -4366 -381 -4327 -364
rect -4293 -381 -4259 -347
rect -4225 -381 -4191 -347
rect -4157 -381 -4123 -347
rect -4089 -381 -4055 -347
rect -4021 -381 -3987 -347
rect -3953 -381 -3919 -347
rect -3885 -381 -3851 -347
rect -3817 -364 -3592 -347
rect -3534 -347 -2574 -300
rect -3534 -364 -3309 -347
rect -3817 -381 -3778 -364
rect -4366 -397 -3778 -381
rect -3348 -381 -3309 -364
rect -3275 -381 -3241 -347
rect -3207 -381 -3173 -347
rect -3139 -381 -3105 -347
rect -3071 -381 -3037 -347
rect -3003 -381 -2969 -347
rect -2935 -381 -2901 -347
rect -2867 -381 -2833 -347
rect -2799 -364 -2574 -347
rect -2516 -347 -1556 -300
rect -2516 -364 -2291 -347
rect -2799 -381 -2760 -364
rect -3348 -397 -2760 -381
rect -2330 -381 -2291 -364
rect -2257 -381 -2223 -347
rect -2189 -381 -2155 -347
rect -2121 -381 -2087 -347
rect -2053 -381 -2019 -347
rect -1985 -381 -1951 -347
rect -1917 -381 -1883 -347
rect -1849 -381 -1815 -347
rect -1781 -364 -1556 -347
rect -1498 -347 -538 -300
rect -1498 -364 -1273 -347
rect -1781 -381 -1742 -364
rect -2330 -397 -1742 -381
rect -1312 -381 -1273 -364
rect -1239 -381 -1205 -347
rect -1171 -381 -1137 -347
rect -1103 -381 -1069 -347
rect -1035 -381 -1001 -347
rect -967 -381 -933 -347
rect -899 -381 -865 -347
rect -831 -381 -797 -347
rect -763 -364 -538 -347
rect -480 -347 480 -300
rect -480 -364 -255 -347
rect -763 -381 -724 -364
rect -1312 -397 -724 -381
rect -294 -381 -255 -364
rect -221 -381 -187 -347
rect -153 -381 -119 -347
rect -85 -381 -51 -347
rect -17 -381 17 -347
rect 51 -381 85 -347
rect 119 -381 153 -347
rect 187 -381 221 -347
rect 255 -364 480 -347
rect 538 -347 1498 -300
rect 538 -364 763 -347
rect 255 -381 294 -364
rect -294 -397 294 -381
rect 724 -381 763 -364
rect 797 -381 831 -347
rect 865 -381 899 -347
rect 933 -381 967 -347
rect 1001 -381 1035 -347
rect 1069 -381 1103 -347
rect 1137 -381 1171 -347
rect 1205 -381 1239 -347
rect 1273 -364 1498 -347
rect 1556 -347 2516 -300
rect 1556 -364 1781 -347
rect 1273 -381 1312 -364
rect 724 -397 1312 -381
rect 1742 -381 1781 -364
rect 1815 -381 1849 -347
rect 1883 -381 1917 -347
rect 1951 -381 1985 -347
rect 2019 -381 2053 -347
rect 2087 -381 2121 -347
rect 2155 -381 2189 -347
rect 2223 -381 2257 -347
rect 2291 -364 2516 -347
rect 2574 -347 3534 -300
rect 2574 -364 2799 -347
rect 2291 -381 2330 -364
rect 1742 -397 2330 -381
rect 2760 -381 2799 -364
rect 2833 -381 2867 -347
rect 2901 -381 2935 -347
rect 2969 -381 3003 -347
rect 3037 -381 3071 -347
rect 3105 -381 3139 -347
rect 3173 -381 3207 -347
rect 3241 -381 3275 -347
rect 3309 -364 3534 -347
rect 3592 -347 4552 -300
rect 3592 -364 3817 -347
rect 3309 -381 3348 -364
rect 2760 -397 3348 -381
rect 3778 -381 3817 -364
rect 3851 -381 3885 -347
rect 3919 -381 3953 -347
rect 3987 -381 4021 -347
rect 4055 -381 4089 -347
rect 4123 -381 4157 -347
rect 4191 -381 4225 -347
rect 4259 -381 4293 -347
rect 4327 -364 4552 -347
rect 4610 -347 5570 -300
rect 4610 -364 4835 -347
rect 4327 -381 4366 -364
rect 3778 -397 4366 -381
rect 4796 -381 4835 -364
rect 4869 -381 4903 -347
rect 4937 -381 4971 -347
rect 5005 -381 5039 -347
rect 5073 -381 5107 -347
rect 5141 -381 5175 -347
rect 5209 -381 5243 -347
rect 5277 -381 5311 -347
rect 5345 -364 5570 -347
rect 5628 -347 6588 -300
rect 5628 -364 5853 -347
rect 5345 -381 5384 -364
rect 4796 -397 5384 -381
rect 5814 -381 5853 -364
rect 5887 -381 5921 -347
rect 5955 -381 5989 -347
rect 6023 -381 6057 -347
rect 6091 -381 6125 -347
rect 6159 -381 6193 -347
rect 6227 -381 6261 -347
rect 6295 -381 6329 -347
rect 6363 -364 6588 -347
rect 6646 -347 7606 -300
rect 6646 -364 6871 -347
rect 6363 -381 6402 -364
rect 5814 -397 6402 -381
rect 6832 -381 6871 -364
rect 6905 -381 6939 -347
rect 6973 -381 7007 -347
rect 7041 -381 7075 -347
rect 7109 -381 7143 -347
rect 7177 -381 7211 -347
rect 7245 -381 7279 -347
rect 7313 -381 7347 -347
rect 7381 -364 7606 -347
rect 7381 -381 7420 -364
rect 6832 -397 7420 -381
<< polycont >>
rect -7381 347 -7347 381
rect -7313 347 -7279 381
rect -7245 347 -7211 381
rect -7177 347 -7143 381
rect -7109 347 -7075 381
rect -7041 347 -7007 381
rect -6973 347 -6939 381
rect -6905 347 -6871 381
rect -6363 347 -6329 381
rect -6295 347 -6261 381
rect -6227 347 -6193 381
rect -6159 347 -6125 381
rect -6091 347 -6057 381
rect -6023 347 -5989 381
rect -5955 347 -5921 381
rect -5887 347 -5853 381
rect -5345 347 -5311 381
rect -5277 347 -5243 381
rect -5209 347 -5175 381
rect -5141 347 -5107 381
rect -5073 347 -5039 381
rect -5005 347 -4971 381
rect -4937 347 -4903 381
rect -4869 347 -4835 381
rect -4327 347 -4293 381
rect -4259 347 -4225 381
rect -4191 347 -4157 381
rect -4123 347 -4089 381
rect -4055 347 -4021 381
rect -3987 347 -3953 381
rect -3919 347 -3885 381
rect -3851 347 -3817 381
rect -3309 347 -3275 381
rect -3241 347 -3207 381
rect -3173 347 -3139 381
rect -3105 347 -3071 381
rect -3037 347 -3003 381
rect -2969 347 -2935 381
rect -2901 347 -2867 381
rect -2833 347 -2799 381
rect -2291 347 -2257 381
rect -2223 347 -2189 381
rect -2155 347 -2121 381
rect -2087 347 -2053 381
rect -2019 347 -1985 381
rect -1951 347 -1917 381
rect -1883 347 -1849 381
rect -1815 347 -1781 381
rect -1273 347 -1239 381
rect -1205 347 -1171 381
rect -1137 347 -1103 381
rect -1069 347 -1035 381
rect -1001 347 -967 381
rect -933 347 -899 381
rect -865 347 -831 381
rect -797 347 -763 381
rect -255 347 -221 381
rect -187 347 -153 381
rect -119 347 -85 381
rect -51 347 -17 381
rect 17 347 51 381
rect 85 347 119 381
rect 153 347 187 381
rect 221 347 255 381
rect 763 347 797 381
rect 831 347 865 381
rect 899 347 933 381
rect 967 347 1001 381
rect 1035 347 1069 381
rect 1103 347 1137 381
rect 1171 347 1205 381
rect 1239 347 1273 381
rect 1781 347 1815 381
rect 1849 347 1883 381
rect 1917 347 1951 381
rect 1985 347 2019 381
rect 2053 347 2087 381
rect 2121 347 2155 381
rect 2189 347 2223 381
rect 2257 347 2291 381
rect 2799 347 2833 381
rect 2867 347 2901 381
rect 2935 347 2969 381
rect 3003 347 3037 381
rect 3071 347 3105 381
rect 3139 347 3173 381
rect 3207 347 3241 381
rect 3275 347 3309 381
rect 3817 347 3851 381
rect 3885 347 3919 381
rect 3953 347 3987 381
rect 4021 347 4055 381
rect 4089 347 4123 381
rect 4157 347 4191 381
rect 4225 347 4259 381
rect 4293 347 4327 381
rect 4835 347 4869 381
rect 4903 347 4937 381
rect 4971 347 5005 381
rect 5039 347 5073 381
rect 5107 347 5141 381
rect 5175 347 5209 381
rect 5243 347 5277 381
rect 5311 347 5345 381
rect 5853 347 5887 381
rect 5921 347 5955 381
rect 5989 347 6023 381
rect 6057 347 6091 381
rect 6125 347 6159 381
rect 6193 347 6227 381
rect 6261 347 6295 381
rect 6329 347 6363 381
rect 6871 347 6905 381
rect 6939 347 6973 381
rect 7007 347 7041 381
rect 7075 347 7109 381
rect 7143 347 7177 381
rect 7211 347 7245 381
rect 7279 347 7313 381
rect 7347 347 7381 381
rect -7381 -381 -7347 -347
rect -7313 -381 -7279 -347
rect -7245 -381 -7211 -347
rect -7177 -381 -7143 -347
rect -7109 -381 -7075 -347
rect -7041 -381 -7007 -347
rect -6973 -381 -6939 -347
rect -6905 -381 -6871 -347
rect -6363 -381 -6329 -347
rect -6295 -381 -6261 -347
rect -6227 -381 -6193 -347
rect -6159 -381 -6125 -347
rect -6091 -381 -6057 -347
rect -6023 -381 -5989 -347
rect -5955 -381 -5921 -347
rect -5887 -381 -5853 -347
rect -5345 -381 -5311 -347
rect -5277 -381 -5243 -347
rect -5209 -381 -5175 -347
rect -5141 -381 -5107 -347
rect -5073 -381 -5039 -347
rect -5005 -381 -4971 -347
rect -4937 -381 -4903 -347
rect -4869 -381 -4835 -347
rect -4327 -381 -4293 -347
rect -4259 -381 -4225 -347
rect -4191 -381 -4157 -347
rect -4123 -381 -4089 -347
rect -4055 -381 -4021 -347
rect -3987 -381 -3953 -347
rect -3919 -381 -3885 -347
rect -3851 -381 -3817 -347
rect -3309 -381 -3275 -347
rect -3241 -381 -3207 -347
rect -3173 -381 -3139 -347
rect -3105 -381 -3071 -347
rect -3037 -381 -3003 -347
rect -2969 -381 -2935 -347
rect -2901 -381 -2867 -347
rect -2833 -381 -2799 -347
rect -2291 -381 -2257 -347
rect -2223 -381 -2189 -347
rect -2155 -381 -2121 -347
rect -2087 -381 -2053 -347
rect -2019 -381 -1985 -347
rect -1951 -381 -1917 -347
rect -1883 -381 -1849 -347
rect -1815 -381 -1781 -347
rect -1273 -381 -1239 -347
rect -1205 -381 -1171 -347
rect -1137 -381 -1103 -347
rect -1069 -381 -1035 -347
rect -1001 -381 -967 -347
rect -933 -381 -899 -347
rect -865 -381 -831 -347
rect -797 -381 -763 -347
rect -255 -381 -221 -347
rect -187 -381 -153 -347
rect -119 -381 -85 -347
rect -51 -381 -17 -347
rect 17 -381 51 -347
rect 85 -381 119 -347
rect 153 -381 187 -347
rect 221 -381 255 -347
rect 763 -381 797 -347
rect 831 -381 865 -347
rect 899 -381 933 -347
rect 967 -381 1001 -347
rect 1035 -381 1069 -347
rect 1103 -381 1137 -347
rect 1171 -381 1205 -347
rect 1239 -381 1273 -347
rect 1781 -381 1815 -347
rect 1849 -381 1883 -347
rect 1917 -381 1951 -347
rect 1985 -381 2019 -347
rect 2053 -381 2087 -347
rect 2121 -381 2155 -347
rect 2189 -381 2223 -347
rect 2257 -381 2291 -347
rect 2799 -381 2833 -347
rect 2867 -381 2901 -347
rect 2935 -381 2969 -347
rect 3003 -381 3037 -347
rect 3071 -381 3105 -347
rect 3139 -381 3173 -347
rect 3207 -381 3241 -347
rect 3275 -381 3309 -347
rect 3817 -381 3851 -347
rect 3885 -381 3919 -347
rect 3953 -381 3987 -347
rect 4021 -381 4055 -347
rect 4089 -381 4123 -347
rect 4157 -381 4191 -347
rect 4225 -381 4259 -347
rect 4293 -381 4327 -347
rect 4835 -381 4869 -347
rect 4903 -381 4937 -347
rect 4971 -381 5005 -347
rect 5039 -381 5073 -347
rect 5107 -381 5141 -347
rect 5175 -381 5209 -347
rect 5243 -381 5277 -347
rect 5311 -381 5345 -347
rect 5853 -381 5887 -347
rect 5921 -381 5955 -347
rect 5989 -381 6023 -347
rect 6057 -381 6091 -347
rect 6125 -381 6159 -347
rect 6193 -381 6227 -347
rect 6261 -381 6295 -347
rect 6329 -381 6363 -347
rect 6871 -381 6905 -347
rect 6939 -381 6973 -347
rect 7007 -381 7041 -347
rect 7075 -381 7109 -347
rect 7143 -381 7177 -347
rect 7211 -381 7245 -347
rect 7279 -381 7313 -347
rect 7347 -381 7381 -347
<< locali >>
rect -7420 347 -7381 381
rect -7347 347 -7323 381
rect -7279 347 -7251 381
rect -7211 347 -7179 381
rect -7143 347 -7109 381
rect -7073 347 -7041 381
rect -7001 347 -6973 381
rect -6929 347 -6905 381
rect -6871 347 -6832 381
rect -6402 347 -6363 381
rect -6329 347 -6305 381
rect -6261 347 -6233 381
rect -6193 347 -6161 381
rect -6125 347 -6091 381
rect -6055 347 -6023 381
rect -5983 347 -5955 381
rect -5911 347 -5887 381
rect -5853 347 -5814 381
rect -5384 347 -5345 381
rect -5311 347 -5287 381
rect -5243 347 -5215 381
rect -5175 347 -5143 381
rect -5107 347 -5073 381
rect -5037 347 -5005 381
rect -4965 347 -4937 381
rect -4893 347 -4869 381
rect -4835 347 -4796 381
rect -4366 347 -4327 381
rect -4293 347 -4269 381
rect -4225 347 -4197 381
rect -4157 347 -4125 381
rect -4089 347 -4055 381
rect -4019 347 -3987 381
rect -3947 347 -3919 381
rect -3875 347 -3851 381
rect -3817 347 -3778 381
rect -3348 347 -3309 381
rect -3275 347 -3251 381
rect -3207 347 -3179 381
rect -3139 347 -3107 381
rect -3071 347 -3037 381
rect -3001 347 -2969 381
rect -2929 347 -2901 381
rect -2857 347 -2833 381
rect -2799 347 -2760 381
rect -2330 347 -2291 381
rect -2257 347 -2233 381
rect -2189 347 -2161 381
rect -2121 347 -2089 381
rect -2053 347 -2019 381
rect -1983 347 -1951 381
rect -1911 347 -1883 381
rect -1839 347 -1815 381
rect -1781 347 -1742 381
rect -1312 347 -1273 381
rect -1239 347 -1215 381
rect -1171 347 -1143 381
rect -1103 347 -1071 381
rect -1035 347 -1001 381
rect -965 347 -933 381
rect -893 347 -865 381
rect -821 347 -797 381
rect -763 347 -724 381
rect -294 347 -255 381
rect -221 347 -197 381
rect -153 347 -125 381
rect -85 347 -53 381
rect -17 347 17 381
rect 53 347 85 381
rect 125 347 153 381
rect 197 347 221 381
rect 255 347 294 381
rect 724 347 763 381
rect 797 347 821 381
rect 865 347 893 381
rect 933 347 965 381
rect 1001 347 1035 381
rect 1071 347 1103 381
rect 1143 347 1171 381
rect 1215 347 1239 381
rect 1273 347 1312 381
rect 1742 347 1781 381
rect 1815 347 1839 381
rect 1883 347 1911 381
rect 1951 347 1983 381
rect 2019 347 2053 381
rect 2089 347 2121 381
rect 2161 347 2189 381
rect 2233 347 2257 381
rect 2291 347 2330 381
rect 2760 347 2799 381
rect 2833 347 2857 381
rect 2901 347 2929 381
rect 2969 347 3001 381
rect 3037 347 3071 381
rect 3107 347 3139 381
rect 3179 347 3207 381
rect 3251 347 3275 381
rect 3309 347 3348 381
rect 3778 347 3817 381
rect 3851 347 3875 381
rect 3919 347 3947 381
rect 3987 347 4019 381
rect 4055 347 4089 381
rect 4125 347 4157 381
rect 4197 347 4225 381
rect 4269 347 4293 381
rect 4327 347 4366 381
rect 4796 347 4835 381
rect 4869 347 4893 381
rect 4937 347 4965 381
rect 5005 347 5037 381
rect 5073 347 5107 381
rect 5143 347 5175 381
rect 5215 347 5243 381
rect 5287 347 5311 381
rect 5345 347 5384 381
rect 5814 347 5853 381
rect 5887 347 5911 381
rect 5955 347 5983 381
rect 6023 347 6055 381
rect 6091 347 6125 381
rect 6161 347 6193 381
rect 6233 347 6261 381
rect 6305 347 6329 381
rect 6363 347 6402 381
rect 6832 347 6871 381
rect 6905 347 6929 381
rect 6973 347 7001 381
rect 7041 347 7073 381
rect 7109 347 7143 381
rect 7179 347 7211 381
rect 7251 347 7279 381
rect 7323 347 7347 381
rect 7381 347 7420 381
rect -7652 269 -7618 304
rect -7652 197 -7618 221
rect -7652 125 -7618 153
rect -7652 53 -7618 85
rect -7652 -17 -7618 17
rect -7652 -85 -7618 -53
rect -7652 -153 -7618 -125
rect -7652 -221 -7618 -197
rect -7652 -304 -7618 -269
rect -6634 269 -6600 304
rect -6634 197 -6600 221
rect -6634 125 -6600 153
rect -6634 53 -6600 85
rect -6634 -17 -6600 17
rect -6634 -85 -6600 -53
rect -6634 -153 -6600 -125
rect -6634 -221 -6600 -197
rect -6634 -304 -6600 -269
rect -5616 269 -5582 304
rect -5616 197 -5582 221
rect -5616 125 -5582 153
rect -5616 53 -5582 85
rect -5616 -17 -5582 17
rect -5616 -85 -5582 -53
rect -5616 -153 -5582 -125
rect -5616 -221 -5582 -197
rect -5616 -304 -5582 -269
rect -4598 269 -4564 304
rect -4598 197 -4564 221
rect -4598 125 -4564 153
rect -4598 53 -4564 85
rect -4598 -17 -4564 17
rect -4598 -85 -4564 -53
rect -4598 -153 -4564 -125
rect -4598 -221 -4564 -197
rect -4598 -304 -4564 -269
rect -3580 269 -3546 304
rect -3580 197 -3546 221
rect -3580 125 -3546 153
rect -3580 53 -3546 85
rect -3580 -17 -3546 17
rect -3580 -85 -3546 -53
rect -3580 -153 -3546 -125
rect -3580 -221 -3546 -197
rect -3580 -304 -3546 -269
rect -2562 269 -2528 304
rect -2562 197 -2528 221
rect -2562 125 -2528 153
rect -2562 53 -2528 85
rect -2562 -17 -2528 17
rect -2562 -85 -2528 -53
rect -2562 -153 -2528 -125
rect -2562 -221 -2528 -197
rect -2562 -304 -2528 -269
rect -1544 269 -1510 304
rect -1544 197 -1510 221
rect -1544 125 -1510 153
rect -1544 53 -1510 85
rect -1544 -17 -1510 17
rect -1544 -85 -1510 -53
rect -1544 -153 -1510 -125
rect -1544 -221 -1510 -197
rect -1544 -304 -1510 -269
rect -526 269 -492 304
rect -526 197 -492 221
rect -526 125 -492 153
rect -526 53 -492 85
rect -526 -17 -492 17
rect -526 -85 -492 -53
rect -526 -153 -492 -125
rect -526 -221 -492 -197
rect -526 -304 -492 -269
rect 492 269 526 304
rect 492 197 526 221
rect 492 125 526 153
rect 492 53 526 85
rect 492 -17 526 17
rect 492 -85 526 -53
rect 492 -153 526 -125
rect 492 -221 526 -197
rect 492 -304 526 -269
rect 1510 269 1544 304
rect 1510 197 1544 221
rect 1510 125 1544 153
rect 1510 53 1544 85
rect 1510 -17 1544 17
rect 1510 -85 1544 -53
rect 1510 -153 1544 -125
rect 1510 -221 1544 -197
rect 1510 -304 1544 -269
rect 2528 269 2562 304
rect 2528 197 2562 221
rect 2528 125 2562 153
rect 2528 53 2562 85
rect 2528 -17 2562 17
rect 2528 -85 2562 -53
rect 2528 -153 2562 -125
rect 2528 -221 2562 -197
rect 2528 -304 2562 -269
rect 3546 269 3580 304
rect 3546 197 3580 221
rect 3546 125 3580 153
rect 3546 53 3580 85
rect 3546 -17 3580 17
rect 3546 -85 3580 -53
rect 3546 -153 3580 -125
rect 3546 -221 3580 -197
rect 3546 -304 3580 -269
rect 4564 269 4598 304
rect 4564 197 4598 221
rect 4564 125 4598 153
rect 4564 53 4598 85
rect 4564 -17 4598 17
rect 4564 -85 4598 -53
rect 4564 -153 4598 -125
rect 4564 -221 4598 -197
rect 4564 -304 4598 -269
rect 5582 269 5616 304
rect 5582 197 5616 221
rect 5582 125 5616 153
rect 5582 53 5616 85
rect 5582 -17 5616 17
rect 5582 -85 5616 -53
rect 5582 -153 5616 -125
rect 5582 -221 5616 -197
rect 5582 -304 5616 -269
rect 6600 269 6634 304
rect 6600 197 6634 221
rect 6600 125 6634 153
rect 6600 53 6634 85
rect 6600 -17 6634 17
rect 6600 -85 6634 -53
rect 6600 -153 6634 -125
rect 6600 -221 6634 -197
rect 6600 -304 6634 -269
rect 7618 269 7652 304
rect 7618 197 7652 221
rect 7618 125 7652 153
rect 7618 53 7652 85
rect 7618 -17 7652 17
rect 7618 -85 7652 -53
rect 7618 -153 7652 -125
rect 7618 -221 7652 -197
rect 7618 -304 7652 -269
rect -7420 -381 -7381 -347
rect -7347 -381 -7323 -347
rect -7279 -381 -7251 -347
rect -7211 -381 -7179 -347
rect -7143 -381 -7109 -347
rect -7073 -381 -7041 -347
rect -7001 -381 -6973 -347
rect -6929 -381 -6905 -347
rect -6871 -381 -6832 -347
rect -6402 -381 -6363 -347
rect -6329 -381 -6305 -347
rect -6261 -381 -6233 -347
rect -6193 -381 -6161 -347
rect -6125 -381 -6091 -347
rect -6055 -381 -6023 -347
rect -5983 -381 -5955 -347
rect -5911 -381 -5887 -347
rect -5853 -381 -5814 -347
rect -5384 -381 -5345 -347
rect -5311 -381 -5287 -347
rect -5243 -381 -5215 -347
rect -5175 -381 -5143 -347
rect -5107 -381 -5073 -347
rect -5037 -381 -5005 -347
rect -4965 -381 -4937 -347
rect -4893 -381 -4869 -347
rect -4835 -381 -4796 -347
rect -4366 -381 -4327 -347
rect -4293 -381 -4269 -347
rect -4225 -381 -4197 -347
rect -4157 -381 -4125 -347
rect -4089 -381 -4055 -347
rect -4019 -381 -3987 -347
rect -3947 -381 -3919 -347
rect -3875 -381 -3851 -347
rect -3817 -381 -3778 -347
rect -3348 -381 -3309 -347
rect -3275 -381 -3251 -347
rect -3207 -381 -3179 -347
rect -3139 -381 -3107 -347
rect -3071 -381 -3037 -347
rect -3001 -381 -2969 -347
rect -2929 -381 -2901 -347
rect -2857 -381 -2833 -347
rect -2799 -381 -2760 -347
rect -2330 -381 -2291 -347
rect -2257 -381 -2233 -347
rect -2189 -381 -2161 -347
rect -2121 -381 -2089 -347
rect -2053 -381 -2019 -347
rect -1983 -381 -1951 -347
rect -1911 -381 -1883 -347
rect -1839 -381 -1815 -347
rect -1781 -381 -1742 -347
rect -1312 -381 -1273 -347
rect -1239 -381 -1215 -347
rect -1171 -381 -1143 -347
rect -1103 -381 -1071 -347
rect -1035 -381 -1001 -347
rect -965 -381 -933 -347
rect -893 -381 -865 -347
rect -821 -381 -797 -347
rect -763 -381 -724 -347
rect -294 -381 -255 -347
rect -221 -381 -197 -347
rect -153 -381 -125 -347
rect -85 -381 -53 -347
rect -17 -381 17 -347
rect 53 -381 85 -347
rect 125 -381 153 -347
rect 197 -381 221 -347
rect 255 -381 294 -347
rect 724 -381 763 -347
rect 797 -381 821 -347
rect 865 -381 893 -347
rect 933 -381 965 -347
rect 1001 -381 1035 -347
rect 1071 -381 1103 -347
rect 1143 -381 1171 -347
rect 1215 -381 1239 -347
rect 1273 -381 1312 -347
rect 1742 -381 1781 -347
rect 1815 -381 1839 -347
rect 1883 -381 1911 -347
rect 1951 -381 1983 -347
rect 2019 -381 2053 -347
rect 2089 -381 2121 -347
rect 2161 -381 2189 -347
rect 2233 -381 2257 -347
rect 2291 -381 2330 -347
rect 2760 -381 2799 -347
rect 2833 -381 2857 -347
rect 2901 -381 2929 -347
rect 2969 -381 3001 -347
rect 3037 -381 3071 -347
rect 3107 -381 3139 -347
rect 3179 -381 3207 -347
rect 3251 -381 3275 -347
rect 3309 -381 3348 -347
rect 3778 -381 3817 -347
rect 3851 -381 3875 -347
rect 3919 -381 3947 -347
rect 3987 -381 4019 -347
rect 4055 -381 4089 -347
rect 4125 -381 4157 -347
rect 4197 -381 4225 -347
rect 4269 -381 4293 -347
rect 4327 -381 4366 -347
rect 4796 -381 4835 -347
rect 4869 -381 4893 -347
rect 4937 -381 4965 -347
rect 5005 -381 5037 -347
rect 5073 -381 5107 -347
rect 5143 -381 5175 -347
rect 5215 -381 5243 -347
rect 5287 -381 5311 -347
rect 5345 -381 5384 -347
rect 5814 -381 5853 -347
rect 5887 -381 5911 -347
rect 5955 -381 5983 -347
rect 6023 -381 6055 -347
rect 6091 -381 6125 -347
rect 6161 -381 6193 -347
rect 6233 -381 6261 -347
rect 6305 -381 6329 -347
rect 6363 -381 6402 -347
rect 6832 -381 6871 -347
rect 6905 -381 6929 -347
rect 6973 -381 7001 -347
rect 7041 -381 7073 -347
rect 7109 -381 7143 -347
rect 7179 -381 7211 -347
rect 7251 -381 7279 -347
rect 7323 -381 7347 -347
rect 7381 -381 7420 -347
<< viali >>
rect -7323 347 -7313 381
rect -7313 347 -7289 381
rect -7251 347 -7245 381
rect -7245 347 -7217 381
rect -7179 347 -7177 381
rect -7177 347 -7145 381
rect -7107 347 -7075 381
rect -7075 347 -7073 381
rect -7035 347 -7007 381
rect -7007 347 -7001 381
rect -6963 347 -6939 381
rect -6939 347 -6929 381
rect -6305 347 -6295 381
rect -6295 347 -6271 381
rect -6233 347 -6227 381
rect -6227 347 -6199 381
rect -6161 347 -6159 381
rect -6159 347 -6127 381
rect -6089 347 -6057 381
rect -6057 347 -6055 381
rect -6017 347 -5989 381
rect -5989 347 -5983 381
rect -5945 347 -5921 381
rect -5921 347 -5911 381
rect -5287 347 -5277 381
rect -5277 347 -5253 381
rect -5215 347 -5209 381
rect -5209 347 -5181 381
rect -5143 347 -5141 381
rect -5141 347 -5109 381
rect -5071 347 -5039 381
rect -5039 347 -5037 381
rect -4999 347 -4971 381
rect -4971 347 -4965 381
rect -4927 347 -4903 381
rect -4903 347 -4893 381
rect -4269 347 -4259 381
rect -4259 347 -4235 381
rect -4197 347 -4191 381
rect -4191 347 -4163 381
rect -4125 347 -4123 381
rect -4123 347 -4091 381
rect -4053 347 -4021 381
rect -4021 347 -4019 381
rect -3981 347 -3953 381
rect -3953 347 -3947 381
rect -3909 347 -3885 381
rect -3885 347 -3875 381
rect -3251 347 -3241 381
rect -3241 347 -3217 381
rect -3179 347 -3173 381
rect -3173 347 -3145 381
rect -3107 347 -3105 381
rect -3105 347 -3073 381
rect -3035 347 -3003 381
rect -3003 347 -3001 381
rect -2963 347 -2935 381
rect -2935 347 -2929 381
rect -2891 347 -2867 381
rect -2867 347 -2857 381
rect -2233 347 -2223 381
rect -2223 347 -2199 381
rect -2161 347 -2155 381
rect -2155 347 -2127 381
rect -2089 347 -2087 381
rect -2087 347 -2055 381
rect -2017 347 -1985 381
rect -1985 347 -1983 381
rect -1945 347 -1917 381
rect -1917 347 -1911 381
rect -1873 347 -1849 381
rect -1849 347 -1839 381
rect -1215 347 -1205 381
rect -1205 347 -1181 381
rect -1143 347 -1137 381
rect -1137 347 -1109 381
rect -1071 347 -1069 381
rect -1069 347 -1037 381
rect -999 347 -967 381
rect -967 347 -965 381
rect -927 347 -899 381
rect -899 347 -893 381
rect -855 347 -831 381
rect -831 347 -821 381
rect -197 347 -187 381
rect -187 347 -163 381
rect -125 347 -119 381
rect -119 347 -91 381
rect -53 347 -51 381
rect -51 347 -19 381
rect 19 347 51 381
rect 51 347 53 381
rect 91 347 119 381
rect 119 347 125 381
rect 163 347 187 381
rect 187 347 197 381
rect 821 347 831 381
rect 831 347 855 381
rect 893 347 899 381
rect 899 347 927 381
rect 965 347 967 381
rect 967 347 999 381
rect 1037 347 1069 381
rect 1069 347 1071 381
rect 1109 347 1137 381
rect 1137 347 1143 381
rect 1181 347 1205 381
rect 1205 347 1215 381
rect 1839 347 1849 381
rect 1849 347 1873 381
rect 1911 347 1917 381
rect 1917 347 1945 381
rect 1983 347 1985 381
rect 1985 347 2017 381
rect 2055 347 2087 381
rect 2087 347 2089 381
rect 2127 347 2155 381
rect 2155 347 2161 381
rect 2199 347 2223 381
rect 2223 347 2233 381
rect 2857 347 2867 381
rect 2867 347 2891 381
rect 2929 347 2935 381
rect 2935 347 2963 381
rect 3001 347 3003 381
rect 3003 347 3035 381
rect 3073 347 3105 381
rect 3105 347 3107 381
rect 3145 347 3173 381
rect 3173 347 3179 381
rect 3217 347 3241 381
rect 3241 347 3251 381
rect 3875 347 3885 381
rect 3885 347 3909 381
rect 3947 347 3953 381
rect 3953 347 3981 381
rect 4019 347 4021 381
rect 4021 347 4053 381
rect 4091 347 4123 381
rect 4123 347 4125 381
rect 4163 347 4191 381
rect 4191 347 4197 381
rect 4235 347 4259 381
rect 4259 347 4269 381
rect 4893 347 4903 381
rect 4903 347 4927 381
rect 4965 347 4971 381
rect 4971 347 4999 381
rect 5037 347 5039 381
rect 5039 347 5071 381
rect 5109 347 5141 381
rect 5141 347 5143 381
rect 5181 347 5209 381
rect 5209 347 5215 381
rect 5253 347 5277 381
rect 5277 347 5287 381
rect 5911 347 5921 381
rect 5921 347 5945 381
rect 5983 347 5989 381
rect 5989 347 6017 381
rect 6055 347 6057 381
rect 6057 347 6089 381
rect 6127 347 6159 381
rect 6159 347 6161 381
rect 6199 347 6227 381
rect 6227 347 6233 381
rect 6271 347 6295 381
rect 6295 347 6305 381
rect 6929 347 6939 381
rect 6939 347 6963 381
rect 7001 347 7007 381
rect 7007 347 7035 381
rect 7073 347 7075 381
rect 7075 347 7107 381
rect 7145 347 7177 381
rect 7177 347 7179 381
rect 7217 347 7245 381
rect 7245 347 7251 381
rect 7289 347 7313 381
rect 7313 347 7323 381
rect -7652 255 -7618 269
rect -7652 235 -7618 255
rect -7652 187 -7618 197
rect -7652 163 -7618 187
rect -7652 119 -7618 125
rect -7652 91 -7618 119
rect -7652 51 -7618 53
rect -7652 19 -7618 51
rect -7652 -51 -7618 -19
rect -7652 -53 -7618 -51
rect -7652 -119 -7618 -91
rect -7652 -125 -7618 -119
rect -7652 -187 -7618 -163
rect -7652 -197 -7618 -187
rect -7652 -255 -7618 -235
rect -7652 -269 -7618 -255
rect -6634 255 -6600 269
rect -6634 235 -6600 255
rect -6634 187 -6600 197
rect -6634 163 -6600 187
rect -6634 119 -6600 125
rect -6634 91 -6600 119
rect -6634 51 -6600 53
rect -6634 19 -6600 51
rect -6634 -51 -6600 -19
rect -6634 -53 -6600 -51
rect -6634 -119 -6600 -91
rect -6634 -125 -6600 -119
rect -6634 -187 -6600 -163
rect -6634 -197 -6600 -187
rect -6634 -255 -6600 -235
rect -6634 -269 -6600 -255
rect -5616 255 -5582 269
rect -5616 235 -5582 255
rect -5616 187 -5582 197
rect -5616 163 -5582 187
rect -5616 119 -5582 125
rect -5616 91 -5582 119
rect -5616 51 -5582 53
rect -5616 19 -5582 51
rect -5616 -51 -5582 -19
rect -5616 -53 -5582 -51
rect -5616 -119 -5582 -91
rect -5616 -125 -5582 -119
rect -5616 -187 -5582 -163
rect -5616 -197 -5582 -187
rect -5616 -255 -5582 -235
rect -5616 -269 -5582 -255
rect -4598 255 -4564 269
rect -4598 235 -4564 255
rect -4598 187 -4564 197
rect -4598 163 -4564 187
rect -4598 119 -4564 125
rect -4598 91 -4564 119
rect -4598 51 -4564 53
rect -4598 19 -4564 51
rect -4598 -51 -4564 -19
rect -4598 -53 -4564 -51
rect -4598 -119 -4564 -91
rect -4598 -125 -4564 -119
rect -4598 -187 -4564 -163
rect -4598 -197 -4564 -187
rect -4598 -255 -4564 -235
rect -4598 -269 -4564 -255
rect -3580 255 -3546 269
rect -3580 235 -3546 255
rect -3580 187 -3546 197
rect -3580 163 -3546 187
rect -3580 119 -3546 125
rect -3580 91 -3546 119
rect -3580 51 -3546 53
rect -3580 19 -3546 51
rect -3580 -51 -3546 -19
rect -3580 -53 -3546 -51
rect -3580 -119 -3546 -91
rect -3580 -125 -3546 -119
rect -3580 -187 -3546 -163
rect -3580 -197 -3546 -187
rect -3580 -255 -3546 -235
rect -3580 -269 -3546 -255
rect -2562 255 -2528 269
rect -2562 235 -2528 255
rect -2562 187 -2528 197
rect -2562 163 -2528 187
rect -2562 119 -2528 125
rect -2562 91 -2528 119
rect -2562 51 -2528 53
rect -2562 19 -2528 51
rect -2562 -51 -2528 -19
rect -2562 -53 -2528 -51
rect -2562 -119 -2528 -91
rect -2562 -125 -2528 -119
rect -2562 -187 -2528 -163
rect -2562 -197 -2528 -187
rect -2562 -255 -2528 -235
rect -2562 -269 -2528 -255
rect -1544 255 -1510 269
rect -1544 235 -1510 255
rect -1544 187 -1510 197
rect -1544 163 -1510 187
rect -1544 119 -1510 125
rect -1544 91 -1510 119
rect -1544 51 -1510 53
rect -1544 19 -1510 51
rect -1544 -51 -1510 -19
rect -1544 -53 -1510 -51
rect -1544 -119 -1510 -91
rect -1544 -125 -1510 -119
rect -1544 -187 -1510 -163
rect -1544 -197 -1510 -187
rect -1544 -255 -1510 -235
rect -1544 -269 -1510 -255
rect -526 255 -492 269
rect -526 235 -492 255
rect -526 187 -492 197
rect -526 163 -492 187
rect -526 119 -492 125
rect -526 91 -492 119
rect -526 51 -492 53
rect -526 19 -492 51
rect -526 -51 -492 -19
rect -526 -53 -492 -51
rect -526 -119 -492 -91
rect -526 -125 -492 -119
rect -526 -187 -492 -163
rect -526 -197 -492 -187
rect -526 -255 -492 -235
rect -526 -269 -492 -255
rect 492 255 526 269
rect 492 235 526 255
rect 492 187 526 197
rect 492 163 526 187
rect 492 119 526 125
rect 492 91 526 119
rect 492 51 526 53
rect 492 19 526 51
rect 492 -51 526 -19
rect 492 -53 526 -51
rect 492 -119 526 -91
rect 492 -125 526 -119
rect 492 -187 526 -163
rect 492 -197 526 -187
rect 492 -255 526 -235
rect 492 -269 526 -255
rect 1510 255 1544 269
rect 1510 235 1544 255
rect 1510 187 1544 197
rect 1510 163 1544 187
rect 1510 119 1544 125
rect 1510 91 1544 119
rect 1510 51 1544 53
rect 1510 19 1544 51
rect 1510 -51 1544 -19
rect 1510 -53 1544 -51
rect 1510 -119 1544 -91
rect 1510 -125 1544 -119
rect 1510 -187 1544 -163
rect 1510 -197 1544 -187
rect 1510 -255 1544 -235
rect 1510 -269 1544 -255
rect 2528 255 2562 269
rect 2528 235 2562 255
rect 2528 187 2562 197
rect 2528 163 2562 187
rect 2528 119 2562 125
rect 2528 91 2562 119
rect 2528 51 2562 53
rect 2528 19 2562 51
rect 2528 -51 2562 -19
rect 2528 -53 2562 -51
rect 2528 -119 2562 -91
rect 2528 -125 2562 -119
rect 2528 -187 2562 -163
rect 2528 -197 2562 -187
rect 2528 -255 2562 -235
rect 2528 -269 2562 -255
rect 3546 255 3580 269
rect 3546 235 3580 255
rect 3546 187 3580 197
rect 3546 163 3580 187
rect 3546 119 3580 125
rect 3546 91 3580 119
rect 3546 51 3580 53
rect 3546 19 3580 51
rect 3546 -51 3580 -19
rect 3546 -53 3580 -51
rect 3546 -119 3580 -91
rect 3546 -125 3580 -119
rect 3546 -187 3580 -163
rect 3546 -197 3580 -187
rect 3546 -255 3580 -235
rect 3546 -269 3580 -255
rect 4564 255 4598 269
rect 4564 235 4598 255
rect 4564 187 4598 197
rect 4564 163 4598 187
rect 4564 119 4598 125
rect 4564 91 4598 119
rect 4564 51 4598 53
rect 4564 19 4598 51
rect 4564 -51 4598 -19
rect 4564 -53 4598 -51
rect 4564 -119 4598 -91
rect 4564 -125 4598 -119
rect 4564 -187 4598 -163
rect 4564 -197 4598 -187
rect 4564 -255 4598 -235
rect 4564 -269 4598 -255
rect 5582 255 5616 269
rect 5582 235 5616 255
rect 5582 187 5616 197
rect 5582 163 5616 187
rect 5582 119 5616 125
rect 5582 91 5616 119
rect 5582 51 5616 53
rect 5582 19 5616 51
rect 5582 -51 5616 -19
rect 5582 -53 5616 -51
rect 5582 -119 5616 -91
rect 5582 -125 5616 -119
rect 5582 -187 5616 -163
rect 5582 -197 5616 -187
rect 5582 -255 5616 -235
rect 5582 -269 5616 -255
rect 6600 255 6634 269
rect 6600 235 6634 255
rect 6600 187 6634 197
rect 6600 163 6634 187
rect 6600 119 6634 125
rect 6600 91 6634 119
rect 6600 51 6634 53
rect 6600 19 6634 51
rect 6600 -51 6634 -19
rect 6600 -53 6634 -51
rect 6600 -119 6634 -91
rect 6600 -125 6634 -119
rect 6600 -187 6634 -163
rect 6600 -197 6634 -187
rect 6600 -255 6634 -235
rect 6600 -269 6634 -255
rect 7618 255 7652 269
rect 7618 235 7652 255
rect 7618 187 7652 197
rect 7618 163 7652 187
rect 7618 119 7652 125
rect 7618 91 7652 119
rect 7618 51 7652 53
rect 7618 19 7652 51
rect 7618 -51 7652 -19
rect 7618 -53 7652 -51
rect 7618 -119 7652 -91
rect 7618 -125 7652 -119
rect 7618 -187 7652 -163
rect 7618 -197 7652 -187
rect 7618 -255 7652 -235
rect 7618 -269 7652 -255
rect -7323 -381 -7313 -347
rect -7313 -381 -7289 -347
rect -7251 -381 -7245 -347
rect -7245 -381 -7217 -347
rect -7179 -381 -7177 -347
rect -7177 -381 -7145 -347
rect -7107 -381 -7075 -347
rect -7075 -381 -7073 -347
rect -7035 -381 -7007 -347
rect -7007 -381 -7001 -347
rect -6963 -381 -6939 -347
rect -6939 -381 -6929 -347
rect -6305 -381 -6295 -347
rect -6295 -381 -6271 -347
rect -6233 -381 -6227 -347
rect -6227 -381 -6199 -347
rect -6161 -381 -6159 -347
rect -6159 -381 -6127 -347
rect -6089 -381 -6057 -347
rect -6057 -381 -6055 -347
rect -6017 -381 -5989 -347
rect -5989 -381 -5983 -347
rect -5945 -381 -5921 -347
rect -5921 -381 -5911 -347
rect -5287 -381 -5277 -347
rect -5277 -381 -5253 -347
rect -5215 -381 -5209 -347
rect -5209 -381 -5181 -347
rect -5143 -381 -5141 -347
rect -5141 -381 -5109 -347
rect -5071 -381 -5039 -347
rect -5039 -381 -5037 -347
rect -4999 -381 -4971 -347
rect -4971 -381 -4965 -347
rect -4927 -381 -4903 -347
rect -4903 -381 -4893 -347
rect -4269 -381 -4259 -347
rect -4259 -381 -4235 -347
rect -4197 -381 -4191 -347
rect -4191 -381 -4163 -347
rect -4125 -381 -4123 -347
rect -4123 -381 -4091 -347
rect -4053 -381 -4021 -347
rect -4021 -381 -4019 -347
rect -3981 -381 -3953 -347
rect -3953 -381 -3947 -347
rect -3909 -381 -3885 -347
rect -3885 -381 -3875 -347
rect -3251 -381 -3241 -347
rect -3241 -381 -3217 -347
rect -3179 -381 -3173 -347
rect -3173 -381 -3145 -347
rect -3107 -381 -3105 -347
rect -3105 -381 -3073 -347
rect -3035 -381 -3003 -347
rect -3003 -381 -3001 -347
rect -2963 -381 -2935 -347
rect -2935 -381 -2929 -347
rect -2891 -381 -2867 -347
rect -2867 -381 -2857 -347
rect -2233 -381 -2223 -347
rect -2223 -381 -2199 -347
rect -2161 -381 -2155 -347
rect -2155 -381 -2127 -347
rect -2089 -381 -2087 -347
rect -2087 -381 -2055 -347
rect -2017 -381 -1985 -347
rect -1985 -381 -1983 -347
rect -1945 -381 -1917 -347
rect -1917 -381 -1911 -347
rect -1873 -381 -1849 -347
rect -1849 -381 -1839 -347
rect -1215 -381 -1205 -347
rect -1205 -381 -1181 -347
rect -1143 -381 -1137 -347
rect -1137 -381 -1109 -347
rect -1071 -381 -1069 -347
rect -1069 -381 -1037 -347
rect -999 -381 -967 -347
rect -967 -381 -965 -347
rect -927 -381 -899 -347
rect -899 -381 -893 -347
rect -855 -381 -831 -347
rect -831 -381 -821 -347
rect -197 -381 -187 -347
rect -187 -381 -163 -347
rect -125 -381 -119 -347
rect -119 -381 -91 -347
rect -53 -381 -51 -347
rect -51 -381 -19 -347
rect 19 -381 51 -347
rect 51 -381 53 -347
rect 91 -381 119 -347
rect 119 -381 125 -347
rect 163 -381 187 -347
rect 187 -381 197 -347
rect 821 -381 831 -347
rect 831 -381 855 -347
rect 893 -381 899 -347
rect 899 -381 927 -347
rect 965 -381 967 -347
rect 967 -381 999 -347
rect 1037 -381 1069 -347
rect 1069 -381 1071 -347
rect 1109 -381 1137 -347
rect 1137 -381 1143 -347
rect 1181 -381 1205 -347
rect 1205 -381 1215 -347
rect 1839 -381 1849 -347
rect 1849 -381 1873 -347
rect 1911 -381 1917 -347
rect 1917 -381 1945 -347
rect 1983 -381 1985 -347
rect 1985 -381 2017 -347
rect 2055 -381 2087 -347
rect 2087 -381 2089 -347
rect 2127 -381 2155 -347
rect 2155 -381 2161 -347
rect 2199 -381 2223 -347
rect 2223 -381 2233 -347
rect 2857 -381 2867 -347
rect 2867 -381 2891 -347
rect 2929 -381 2935 -347
rect 2935 -381 2963 -347
rect 3001 -381 3003 -347
rect 3003 -381 3035 -347
rect 3073 -381 3105 -347
rect 3105 -381 3107 -347
rect 3145 -381 3173 -347
rect 3173 -381 3179 -347
rect 3217 -381 3241 -347
rect 3241 -381 3251 -347
rect 3875 -381 3885 -347
rect 3885 -381 3909 -347
rect 3947 -381 3953 -347
rect 3953 -381 3981 -347
rect 4019 -381 4021 -347
rect 4021 -381 4053 -347
rect 4091 -381 4123 -347
rect 4123 -381 4125 -347
rect 4163 -381 4191 -347
rect 4191 -381 4197 -347
rect 4235 -381 4259 -347
rect 4259 -381 4269 -347
rect 4893 -381 4903 -347
rect 4903 -381 4927 -347
rect 4965 -381 4971 -347
rect 4971 -381 4999 -347
rect 5037 -381 5039 -347
rect 5039 -381 5071 -347
rect 5109 -381 5141 -347
rect 5141 -381 5143 -347
rect 5181 -381 5209 -347
rect 5209 -381 5215 -347
rect 5253 -381 5277 -347
rect 5277 -381 5287 -347
rect 5911 -381 5921 -347
rect 5921 -381 5945 -347
rect 5983 -381 5989 -347
rect 5989 -381 6017 -347
rect 6055 -381 6057 -347
rect 6057 -381 6089 -347
rect 6127 -381 6159 -347
rect 6159 -381 6161 -347
rect 6199 -381 6227 -347
rect 6227 -381 6233 -347
rect 6271 -381 6295 -347
rect 6295 -381 6305 -347
rect 6929 -381 6939 -347
rect 6939 -381 6963 -347
rect 7001 -381 7007 -347
rect 7007 -381 7035 -347
rect 7073 -381 7075 -347
rect 7075 -381 7107 -347
rect 7145 -381 7177 -347
rect 7177 -381 7179 -347
rect 7217 -381 7245 -347
rect 7245 -381 7251 -347
rect 7289 -381 7313 -347
rect 7313 -381 7323 -347
<< metal1 >>
rect -7370 381 -6882 387
rect -7370 347 -7323 381
rect -7289 347 -7251 381
rect -7217 347 -7179 381
rect -7145 347 -7107 381
rect -7073 347 -7035 381
rect -7001 347 -6963 381
rect -6929 347 -6882 381
rect -7370 341 -6882 347
rect -6352 381 -5864 387
rect -6352 347 -6305 381
rect -6271 347 -6233 381
rect -6199 347 -6161 381
rect -6127 347 -6089 381
rect -6055 347 -6017 381
rect -5983 347 -5945 381
rect -5911 347 -5864 381
rect -6352 341 -5864 347
rect -5334 381 -4846 387
rect -5334 347 -5287 381
rect -5253 347 -5215 381
rect -5181 347 -5143 381
rect -5109 347 -5071 381
rect -5037 347 -4999 381
rect -4965 347 -4927 381
rect -4893 347 -4846 381
rect -5334 341 -4846 347
rect -4316 381 -3828 387
rect -4316 347 -4269 381
rect -4235 347 -4197 381
rect -4163 347 -4125 381
rect -4091 347 -4053 381
rect -4019 347 -3981 381
rect -3947 347 -3909 381
rect -3875 347 -3828 381
rect -4316 341 -3828 347
rect -3298 381 -2810 387
rect -3298 347 -3251 381
rect -3217 347 -3179 381
rect -3145 347 -3107 381
rect -3073 347 -3035 381
rect -3001 347 -2963 381
rect -2929 347 -2891 381
rect -2857 347 -2810 381
rect -3298 341 -2810 347
rect -2280 381 -1792 387
rect -2280 347 -2233 381
rect -2199 347 -2161 381
rect -2127 347 -2089 381
rect -2055 347 -2017 381
rect -1983 347 -1945 381
rect -1911 347 -1873 381
rect -1839 347 -1792 381
rect -2280 341 -1792 347
rect -1262 381 -774 387
rect -1262 347 -1215 381
rect -1181 347 -1143 381
rect -1109 347 -1071 381
rect -1037 347 -999 381
rect -965 347 -927 381
rect -893 347 -855 381
rect -821 347 -774 381
rect -1262 341 -774 347
rect -244 381 244 387
rect -244 347 -197 381
rect -163 347 -125 381
rect -91 347 -53 381
rect -19 347 19 381
rect 53 347 91 381
rect 125 347 163 381
rect 197 347 244 381
rect -244 341 244 347
rect 774 381 1262 387
rect 774 347 821 381
rect 855 347 893 381
rect 927 347 965 381
rect 999 347 1037 381
rect 1071 347 1109 381
rect 1143 347 1181 381
rect 1215 347 1262 381
rect 774 341 1262 347
rect 1792 381 2280 387
rect 1792 347 1839 381
rect 1873 347 1911 381
rect 1945 347 1983 381
rect 2017 347 2055 381
rect 2089 347 2127 381
rect 2161 347 2199 381
rect 2233 347 2280 381
rect 1792 341 2280 347
rect 2810 381 3298 387
rect 2810 347 2857 381
rect 2891 347 2929 381
rect 2963 347 3001 381
rect 3035 347 3073 381
rect 3107 347 3145 381
rect 3179 347 3217 381
rect 3251 347 3298 381
rect 2810 341 3298 347
rect 3828 381 4316 387
rect 3828 347 3875 381
rect 3909 347 3947 381
rect 3981 347 4019 381
rect 4053 347 4091 381
rect 4125 347 4163 381
rect 4197 347 4235 381
rect 4269 347 4316 381
rect 3828 341 4316 347
rect 4846 381 5334 387
rect 4846 347 4893 381
rect 4927 347 4965 381
rect 4999 347 5037 381
rect 5071 347 5109 381
rect 5143 347 5181 381
rect 5215 347 5253 381
rect 5287 347 5334 381
rect 4846 341 5334 347
rect 5864 381 6352 387
rect 5864 347 5911 381
rect 5945 347 5983 381
rect 6017 347 6055 381
rect 6089 347 6127 381
rect 6161 347 6199 381
rect 6233 347 6271 381
rect 6305 347 6352 381
rect 5864 341 6352 347
rect 6882 381 7370 387
rect 6882 347 6929 381
rect 6963 347 7001 381
rect 7035 347 7073 381
rect 7107 347 7145 381
rect 7179 347 7217 381
rect 7251 347 7289 381
rect 7323 347 7370 381
rect 6882 341 7370 347
rect -7658 269 -7612 300
rect -7658 235 -7652 269
rect -7618 235 -7612 269
rect -7658 197 -7612 235
rect -7658 163 -7652 197
rect -7618 163 -7612 197
rect -7658 125 -7612 163
rect -7658 91 -7652 125
rect -7618 91 -7612 125
rect -7658 53 -7612 91
rect -7658 19 -7652 53
rect -7618 19 -7612 53
rect -7658 -19 -7612 19
rect -7658 -53 -7652 -19
rect -7618 -53 -7612 -19
rect -7658 -91 -7612 -53
rect -7658 -125 -7652 -91
rect -7618 -125 -7612 -91
rect -7658 -163 -7612 -125
rect -7658 -197 -7652 -163
rect -7618 -197 -7612 -163
rect -7658 -235 -7612 -197
rect -7658 -269 -7652 -235
rect -7618 -269 -7612 -235
rect -7658 -300 -7612 -269
rect -6640 269 -6594 300
rect -6640 235 -6634 269
rect -6600 235 -6594 269
rect -6640 197 -6594 235
rect -6640 163 -6634 197
rect -6600 163 -6594 197
rect -6640 125 -6594 163
rect -6640 91 -6634 125
rect -6600 91 -6594 125
rect -6640 53 -6594 91
rect -6640 19 -6634 53
rect -6600 19 -6594 53
rect -6640 -19 -6594 19
rect -6640 -53 -6634 -19
rect -6600 -53 -6594 -19
rect -6640 -91 -6594 -53
rect -6640 -125 -6634 -91
rect -6600 -125 -6594 -91
rect -6640 -163 -6594 -125
rect -6640 -197 -6634 -163
rect -6600 -197 -6594 -163
rect -6640 -235 -6594 -197
rect -6640 -269 -6634 -235
rect -6600 -269 -6594 -235
rect -6640 -300 -6594 -269
rect -5622 269 -5576 300
rect -5622 235 -5616 269
rect -5582 235 -5576 269
rect -5622 197 -5576 235
rect -5622 163 -5616 197
rect -5582 163 -5576 197
rect -5622 125 -5576 163
rect -5622 91 -5616 125
rect -5582 91 -5576 125
rect -5622 53 -5576 91
rect -5622 19 -5616 53
rect -5582 19 -5576 53
rect -5622 -19 -5576 19
rect -5622 -53 -5616 -19
rect -5582 -53 -5576 -19
rect -5622 -91 -5576 -53
rect -5622 -125 -5616 -91
rect -5582 -125 -5576 -91
rect -5622 -163 -5576 -125
rect -5622 -197 -5616 -163
rect -5582 -197 -5576 -163
rect -5622 -235 -5576 -197
rect -5622 -269 -5616 -235
rect -5582 -269 -5576 -235
rect -5622 -300 -5576 -269
rect -4604 269 -4558 300
rect -4604 235 -4598 269
rect -4564 235 -4558 269
rect -4604 197 -4558 235
rect -4604 163 -4598 197
rect -4564 163 -4558 197
rect -4604 125 -4558 163
rect -4604 91 -4598 125
rect -4564 91 -4558 125
rect -4604 53 -4558 91
rect -4604 19 -4598 53
rect -4564 19 -4558 53
rect -4604 -19 -4558 19
rect -4604 -53 -4598 -19
rect -4564 -53 -4558 -19
rect -4604 -91 -4558 -53
rect -4604 -125 -4598 -91
rect -4564 -125 -4558 -91
rect -4604 -163 -4558 -125
rect -4604 -197 -4598 -163
rect -4564 -197 -4558 -163
rect -4604 -235 -4558 -197
rect -4604 -269 -4598 -235
rect -4564 -269 -4558 -235
rect -4604 -300 -4558 -269
rect -3586 269 -3540 300
rect -3586 235 -3580 269
rect -3546 235 -3540 269
rect -3586 197 -3540 235
rect -3586 163 -3580 197
rect -3546 163 -3540 197
rect -3586 125 -3540 163
rect -3586 91 -3580 125
rect -3546 91 -3540 125
rect -3586 53 -3540 91
rect -3586 19 -3580 53
rect -3546 19 -3540 53
rect -3586 -19 -3540 19
rect -3586 -53 -3580 -19
rect -3546 -53 -3540 -19
rect -3586 -91 -3540 -53
rect -3586 -125 -3580 -91
rect -3546 -125 -3540 -91
rect -3586 -163 -3540 -125
rect -3586 -197 -3580 -163
rect -3546 -197 -3540 -163
rect -3586 -235 -3540 -197
rect -3586 -269 -3580 -235
rect -3546 -269 -3540 -235
rect -3586 -300 -3540 -269
rect -2568 269 -2522 300
rect -2568 235 -2562 269
rect -2528 235 -2522 269
rect -2568 197 -2522 235
rect -2568 163 -2562 197
rect -2528 163 -2522 197
rect -2568 125 -2522 163
rect -2568 91 -2562 125
rect -2528 91 -2522 125
rect -2568 53 -2522 91
rect -2568 19 -2562 53
rect -2528 19 -2522 53
rect -2568 -19 -2522 19
rect -2568 -53 -2562 -19
rect -2528 -53 -2522 -19
rect -2568 -91 -2522 -53
rect -2568 -125 -2562 -91
rect -2528 -125 -2522 -91
rect -2568 -163 -2522 -125
rect -2568 -197 -2562 -163
rect -2528 -197 -2522 -163
rect -2568 -235 -2522 -197
rect -2568 -269 -2562 -235
rect -2528 -269 -2522 -235
rect -2568 -300 -2522 -269
rect -1550 269 -1504 300
rect -1550 235 -1544 269
rect -1510 235 -1504 269
rect -1550 197 -1504 235
rect -1550 163 -1544 197
rect -1510 163 -1504 197
rect -1550 125 -1504 163
rect -1550 91 -1544 125
rect -1510 91 -1504 125
rect -1550 53 -1504 91
rect -1550 19 -1544 53
rect -1510 19 -1504 53
rect -1550 -19 -1504 19
rect -1550 -53 -1544 -19
rect -1510 -53 -1504 -19
rect -1550 -91 -1504 -53
rect -1550 -125 -1544 -91
rect -1510 -125 -1504 -91
rect -1550 -163 -1504 -125
rect -1550 -197 -1544 -163
rect -1510 -197 -1504 -163
rect -1550 -235 -1504 -197
rect -1550 -269 -1544 -235
rect -1510 -269 -1504 -235
rect -1550 -300 -1504 -269
rect -532 269 -486 300
rect -532 235 -526 269
rect -492 235 -486 269
rect -532 197 -486 235
rect -532 163 -526 197
rect -492 163 -486 197
rect -532 125 -486 163
rect -532 91 -526 125
rect -492 91 -486 125
rect -532 53 -486 91
rect -532 19 -526 53
rect -492 19 -486 53
rect -532 -19 -486 19
rect -532 -53 -526 -19
rect -492 -53 -486 -19
rect -532 -91 -486 -53
rect -532 -125 -526 -91
rect -492 -125 -486 -91
rect -532 -163 -486 -125
rect -532 -197 -526 -163
rect -492 -197 -486 -163
rect -532 -235 -486 -197
rect -532 -269 -526 -235
rect -492 -269 -486 -235
rect -532 -300 -486 -269
rect 486 269 532 300
rect 486 235 492 269
rect 526 235 532 269
rect 486 197 532 235
rect 486 163 492 197
rect 526 163 532 197
rect 486 125 532 163
rect 486 91 492 125
rect 526 91 532 125
rect 486 53 532 91
rect 486 19 492 53
rect 526 19 532 53
rect 486 -19 532 19
rect 486 -53 492 -19
rect 526 -53 532 -19
rect 486 -91 532 -53
rect 486 -125 492 -91
rect 526 -125 532 -91
rect 486 -163 532 -125
rect 486 -197 492 -163
rect 526 -197 532 -163
rect 486 -235 532 -197
rect 486 -269 492 -235
rect 526 -269 532 -235
rect 486 -300 532 -269
rect 1504 269 1550 300
rect 1504 235 1510 269
rect 1544 235 1550 269
rect 1504 197 1550 235
rect 1504 163 1510 197
rect 1544 163 1550 197
rect 1504 125 1550 163
rect 1504 91 1510 125
rect 1544 91 1550 125
rect 1504 53 1550 91
rect 1504 19 1510 53
rect 1544 19 1550 53
rect 1504 -19 1550 19
rect 1504 -53 1510 -19
rect 1544 -53 1550 -19
rect 1504 -91 1550 -53
rect 1504 -125 1510 -91
rect 1544 -125 1550 -91
rect 1504 -163 1550 -125
rect 1504 -197 1510 -163
rect 1544 -197 1550 -163
rect 1504 -235 1550 -197
rect 1504 -269 1510 -235
rect 1544 -269 1550 -235
rect 1504 -300 1550 -269
rect 2522 269 2568 300
rect 2522 235 2528 269
rect 2562 235 2568 269
rect 2522 197 2568 235
rect 2522 163 2528 197
rect 2562 163 2568 197
rect 2522 125 2568 163
rect 2522 91 2528 125
rect 2562 91 2568 125
rect 2522 53 2568 91
rect 2522 19 2528 53
rect 2562 19 2568 53
rect 2522 -19 2568 19
rect 2522 -53 2528 -19
rect 2562 -53 2568 -19
rect 2522 -91 2568 -53
rect 2522 -125 2528 -91
rect 2562 -125 2568 -91
rect 2522 -163 2568 -125
rect 2522 -197 2528 -163
rect 2562 -197 2568 -163
rect 2522 -235 2568 -197
rect 2522 -269 2528 -235
rect 2562 -269 2568 -235
rect 2522 -300 2568 -269
rect 3540 269 3586 300
rect 3540 235 3546 269
rect 3580 235 3586 269
rect 3540 197 3586 235
rect 3540 163 3546 197
rect 3580 163 3586 197
rect 3540 125 3586 163
rect 3540 91 3546 125
rect 3580 91 3586 125
rect 3540 53 3586 91
rect 3540 19 3546 53
rect 3580 19 3586 53
rect 3540 -19 3586 19
rect 3540 -53 3546 -19
rect 3580 -53 3586 -19
rect 3540 -91 3586 -53
rect 3540 -125 3546 -91
rect 3580 -125 3586 -91
rect 3540 -163 3586 -125
rect 3540 -197 3546 -163
rect 3580 -197 3586 -163
rect 3540 -235 3586 -197
rect 3540 -269 3546 -235
rect 3580 -269 3586 -235
rect 3540 -300 3586 -269
rect 4558 269 4604 300
rect 4558 235 4564 269
rect 4598 235 4604 269
rect 4558 197 4604 235
rect 4558 163 4564 197
rect 4598 163 4604 197
rect 4558 125 4604 163
rect 4558 91 4564 125
rect 4598 91 4604 125
rect 4558 53 4604 91
rect 4558 19 4564 53
rect 4598 19 4604 53
rect 4558 -19 4604 19
rect 4558 -53 4564 -19
rect 4598 -53 4604 -19
rect 4558 -91 4604 -53
rect 4558 -125 4564 -91
rect 4598 -125 4604 -91
rect 4558 -163 4604 -125
rect 4558 -197 4564 -163
rect 4598 -197 4604 -163
rect 4558 -235 4604 -197
rect 4558 -269 4564 -235
rect 4598 -269 4604 -235
rect 4558 -300 4604 -269
rect 5576 269 5622 300
rect 5576 235 5582 269
rect 5616 235 5622 269
rect 5576 197 5622 235
rect 5576 163 5582 197
rect 5616 163 5622 197
rect 5576 125 5622 163
rect 5576 91 5582 125
rect 5616 91 5622 125
rect 5576 53 5622 91
rect 5576 19 5582 53
rect 5616 19 5622 53
rect 5576 -19 5622 19
rect 5576 -53 5582 -19
rect 5616 -53 5622 -19
rect 5576 -91 5622 -53
rect 5576 -125 5582 -91
rect 5616 -125 5622 -91
rect 5576 -163 5622 -125
rect 5576 -197 5582 -163
rect 5616 -197 5622 -163
rect 5576 -235 5622 -197
rect 5576 -269 5582 -235
rect 5616 -269 5622 -235
rect 5576 -300 5622 -269
rect 6594 269 6640 300
rect 6594 235 6600 269
rect 6634 235 6640 269
rect 6594 197 6640 235
rect 6594 163 6600 197
rect 6634 163 6640 197
rect 6594 125 6640 163
rect 6594 91 6600 125
rect 6634 91 6640 125
rect 6594 53 6640 91
rect 6594 19 6600 53
rect 6634 19 6640 53
rect 6594 -19 6640 19
rect 6594 -53 6600 -19
rect 6634 -53 6640 -19
rect 6594 -91 6640 -53
rect 6594 -125 6600 -91
rect 6634 -125 6640 -91
rect 6594 -163 6640 -125
rect 6594 -197 6600 -163
rect 6634 -197 6640 -163
rect 6594 -235 6640 -197
rect 6594 -269 6600 -235
rect 6634 -269 6640 -235
rect 6594 -300 6640 -269
rect 7612 269 7658 300
rect 7612 235 7618 269
rect 7652 235 7658 269
rect 7612 197 7658 235
rect 7612 163 7618 197
rect 7652 163 7658 197
rect 7612 125 7658 163
rect 7612 91 7618 125
rect 7652 91 7658 125
rect 7612 53 7658 91
rect 7612 19 7618 53
rect 7652 19 7658 53
rect 7612 -19 7658 19
rect 7612 -53 7618 -19
rect 7652 -53 7658 -19
rect 7612 -91 7658 -53
rect 7612 -125 7618 -91
rect 7652 -125 7658 -91
rect 7612 -163 7658 -125
rect 7612 -197 7618 -163
rect 7652 -197 7658 -163
rect 7612 -235 7658 -197
rect 7612 -269 7618 -235
rect 7652 -269 7658 -235
rect 7612 -300 7658 -269
rect -7370 -347 -6882 -341
rect -7370 -381 -7323 -347
rect -7289 -381 -7251 -347
rect -7217 -381 -7179 -347
rect -7145 -381 -7107 -347
rect -7073 -381 -7035 -347
rect -7001 -381 -6963 -347
rect -6929 -381 -6882 -347
rect -7370 -387 -6882 -381
rect -6352 -347 -5864 -341
rect -6352 -381 -6305 -347
rect -6271 -381 -6233 -347
rect -6199 -381 -6161 -347
rect -6127 -381 -6089 -347
rect -6055 -381 -6017 -347
rect -5983 -381 -5945 -347
rect -5911 -381 -5864 -347
rect -6352 -387 -5864 -381
rect -5334 -347 -4846 -341
rect -5334 -381 -5287 -347
rect -5253 -381 -5215 -347
rect -5181 -381 -5143 -347
rect -5109 -381 -5071 -347
rect -5037 -381 -4999 -347
rect -4965 -381 -4927 -347
rect -4893 -381 -4846 -347
rect -5334 -387 -4846 -381
rect -4316 -347 -3828 -341
rect -4316 -381 -4269 -347
rect -4235 -381 -4197 -347
rect -4163 -381 -4125 -347
rect -4091 -381 -4053 -347
rect -4019 -381 -3981 -347
rect -3947 -381 -3909 -347
rect -3875 -381 -3828 -347
rect -4316 -387 -3828 -381
rect -3298 -347 -2810 -341
rect -3298 -381 -3251 -347
rect -3217 -381 -3179 -347
rect -3145 -381 -3107 -347
rect -3073 -381 -3035 -347
rect -3001 -381 -2963 -347
rect -2929 -381 -2891 -347
rect -2857 -381 -2810 -347
rect -3298 -387 -2810 -381
rect -2280 -347 -1792 -341
rect -2280 -381 -2233 -347
rect -2199 -381 -2161 -347
rect -2127 -381 -2089 -347
rect -2055 -381 -2017 -347
rect -1983 -381 -1945 -347
rect -1911 -381 -1873 -347
rect -1839 -381 -1792 -347
rect -2280 -387 -1792 -381
rect -1262 -347 -774 -341
rect -1262 -381 -1215 -347
rect -1181 -381 -1143 -347
rect -1109 -381 -1071 -347
rect -1037 -381 -999 -347
rect -965 -381 -927 -347
rect -893 -381 -855 -347
rect -821 -381 -774 -347
rect -1262 -387 -774 -381
rect -244 -347 244 -341
rect -244 -381 -197 -347
rect -163 -381 -125 -347
rect -91 -381 -53 -347
rect -19 -381 19 -347
rect 53 -381 91 -347
rect 125 -381 163 -347
rect 197 -381 244 -347
rect -244 -387 244 -381
rect 774 -347 1262 -341
rect 774 -381 821 -347
rect 855 -381 893 -347
rect 927 -381 965 -347
rect 999 -381 1037 -347
rect 1071 -381 1109 -347
rect 1143 -381 1181 -347
rect 1215 -381 1262 -347
rect 774 -387 1262 -381
rect 1792 -347 2280 -341
rect 1792 -381 1839 -347
rect 1873 -381 1911 -347
rect 1945 -381 1983 -347
rect 2017 -381 2055 -347
rect 2089 -381 2127 -347
rect 2161 -381 2199 -347
rect 2233 -381 2280 -347
rect 1792 -387 2280 -381
rect 2810 -347 3298 -341
rect 2810 -381 2857 -347
rect 2891 -381 2929 -347
rect 2963 -381 3001 -347
rect 3035 -381 3073 -347
rect 3107 -381 3145 -347
rect 3179 -381 3217 -347
rect 3251 -381 3298 -347
rect 2810 -387 3298 -381
rect 3828 -347 4316 -341
rect 3828 -381 3875 -347
rect 3909 -381 3947 -347
rect 3981 -381 4019 -347
rect 4053 -381 4091 -347
rect 4125 -381 4163 -347
rect 4197 -381 4235 -347
rect 4269 -381 4316 -347
rect 3828 -387 4316 -381
rect 4846 -347 5334 -341
rect 4846 -381 4893 -347
rect 4927 -381 4965 -347
rect 4999 -381 5037 -347
rect 5071 -381 5109 -347
rect 5143 -381 5181 -347
rect 5215 -381 5253 -347
rect 5287 -381 5334 -347
rect 4846 -387 5334 -381
rect 5864 -347 6352 -341
rect 5864 -381 5911 -347
rect 5945 -381 5983 -347
rect 6017 -381 6055 -347
rect 6089 -381 6127 -347
rect 6161 -381 6199 -347
rect 6233 -381 6271 -347
rect 6305 -381 6352 -347
rect 5864 -387 6352 -381
rect 6882 -347 7370 -341
rect 6882 -381 6929 -347
rect 6963 -381 7001 -347
rect 7035 -381 7073 -347
rect 7107 -381 7145 -347
rect 7179 -381 7217 -347
rect 7251 -381 7289 -347
rect 7323 -381 7370 -347
rect 6882 -387 7370 -381
<< end >>
