magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -3660 -4438 3660 4438
<< nwell >>
rect -2000 400 2000 2400
rect -2400 -400 2400 -40
rect -2400 -2400 -2000 -400
rect 2000 -2400 2400 -400
rect -2400 -2800 2400 -2400
<< pwell >>
rect -2360 2524 2360 2760
rect -2360 316 -2124 2524
rect 2124 316 2360 2524
rect -2360 80 2360 316
rect -1960 -676 1960 -440
rect -1960 -2124 -1724 -676
rect 1724 -2124 1960 -676
rect -1960 -2360 1960 -2124
<< mvpsubdiff >>
rect -2334 2693 2334 2734
rect -2334 2591 -2091 2693
rect 2091 2591 2334 2693
rect -2334 2550 2334 2591
rect -2334 2491 -2150 2550
rect -2334 349 -2293 2491
rect -2191 349 -2150 2491
rect 2150 2491 2334 2550
rect -2334 290 -2150 349
rect 2150 349 2191 2491
rect 2293 349 2334 2491
rect 2150 290 2334 349
rect -2334 249 2334 290
rect -2334 147 -2091 249
rect 2091 147 2334 249
rect -2334 106 2334 147
rect -1934 -507 1934 -466
rect -1934 -609 -1683 -507
rect 1683 -609 1934 -507
rect -1934 -650 1934 -609
rect -1934 -703 -1750 -650
rect -1934 -2097 -1893 -703
rect -1791 -2097 -1750 -703
rect -1934 -2150 -1750 -2097
rect 1750 -703 1934 -650
rect 1750 -2097 1791 -703
rect 1893 -2097 1934 -703
rect 1750 -2150 1934 -2097
rect -1934 -2191 1934 -2150
rect -1934 -2293 -1683 -2191
rect 1683 -2293 1934 -2191
rect -1934 -2334 1934 -2293
<< mvnsubdiff >>
rect -1934 2293 1934 2334
rect -1934 2191 -1683 2293
rect 1683 2191 1934 2293
rect -1934 2150 1934 2191
rect -1934 2097 -1750 2150
rect -1934 703 -1893 2097
rect -1791 703 -1750 2097
rect -1934 650 -1750 703
rect 1750 2097 1934 2150
rect 1750 703 1791 2097
rect 1893 703 1934 2097
rect 1750 650 1934 703
rect -1934 609 1934 650
rect -1934 507 -1683 609
rect 1683 507 1934 609
rect -1934 466 1934 507
rect -2334 -147 2334 -106
rect -2334 -249 -2091 -147
rect 2091 -249 2334 -147
rect -2334 -290 2334 -249
rect -2334 -349 -2150 -290
rect -2334 -2491 -2293 -349
rect -2191 -2491 -2150 -349
rect 2150 -349 2334 -290
rect -2334 -2550 -2150 -2491
rect 2150 -2491 2191 -349
rect 2293 -2491 2334 -349
rect 2150 -2550 2334 -2491
rect -2334 -2591 2334 -2550
rect -2334 -2693 -2091 -2591
rect 2091 -2693 2334 -2591
rect -2334 -2734 2334 -2693
<< mvpsubdiffcont >>
rect -2091 2591 2091 2693
rect -2293 349 -2191 2491
rect 2191 349 2293 2491
rect -2091 147 2091 249
rect -1683 -609 1683 -507
rect -1893 -2097 -1791 -703
rect 1791 -2097 1893 -703
rect -1683 -2293 1683 -2191
<< mvnsubdiffcont >>
rect -1683 2191 1683 2293
rect -1893 703 -1791 2097
rect 1791 703 1893 2097
rect -1683 507 1683 609
rect -2091 -249 2091 -147
rect -2293 -2491 -2191 -349
rect 2191 -2491 2293 -349
rect -2091 -2693 2091 -2591
<< locali >>
rect -2322 2695 2322 2722
rect -2322 2589 -2141 2695
rect 2141 2589 2322 2695
rect -2322 2562 2322 2589
rect -2322 2491 -2162 2562
rect -2322 2445 -2293 2491
rect -2191 2445 -2162 2491
rect -2322 395 -2295 2445
rect -2189 395 -2162 2445
rect 2162 2491 2322 2562
rect 2162 2445 2191 2491
rect 2293 2445 2322 2491
rect -1922 2295 1922 2322
rect -1922 2189 -1745 2295
rect 1745 2189 1922 2295
rect -1922 2162 1922 2189
rect -1922 2097 -1762 2162
rect -1922 2065 -1893 2097
rect -1791 2065 -1762 2097
rect -1922 735 -1895 2065
rect -1789 735 -1762 2065
rect 1762 2097 1922 2162
rect 1762 2065 1791 2097
rect 1893 2065 1922 2097
rect -1603 1947 -1601 1981
rect -1567 1947 -1529 1981
rect -1495 1947 -1457 1981
rect -1423 1947 -1385 1981
rect -1351 1947 -1313 1981
rect -1279 1947 -1241 1981
rect -1207 1947 -1169 1981
rect -1135 1947 -1097 1981
rect -1063 1947 -1025 1981
rect -991 1947 -953 1981
rect -919 1947 -881 1981
rect -847 1947 -809 1981
rect -775 1947 -737 1981
rect -703 1947 -665 1981
rect -631 1947 -593 1981
rect -559 1947 -521 1981
rect -487 1947 -449 1981
rect -415 1947 -377 1981
rect -343 1947 -305 1981
rect -271 1947 -233 1981
rect -199 1947 -161 1981
rect -127 1947 -89 1981
rect -55 1947 -17 1981
rect 17 1947 55 1981
rect 89 1947 127 1981
rect 161 1947 199 1981
rect 233 1947 271 1981
rect 305 1947 343 1981
rect 377 1947 415 1981
rect 449 1947 487 1981
rect 521 1947 559 1981
rect 593 1947 631 1981
rect 665 1947 703 1981
rect 737 1947 775 1981
rect 809 1947 847 1981
rect 881 1947 919 1981
rect 953 1947 991 1981
rect 1025 1947 1063 1981
rect 1097 1947 1135 1981
rect 1169 1947 1207 1981
rect 1241 1947 1279 1981
rect 1313 1947 1351 1981
rect 1385 1947 1423 1981
rect 1457 1947 1495 1981
rect 1529 1947 1567 1981
rect 1601 1947 1603 1981
rect -1922 703 -1893 735
rect -1791 703 -1762 735
rect -1922 638 -1762 703
rect 1762 735 1789 2065
rect 1895 735 1922 2065
rect 1762 703 1791 735
rect 1893 703 1922 735
rect 1762 638 1922 703
rect -1922 611 1922 638
rect -1922 505 -1745 611
rect 1745 505 1922 611
rect -1922 478 1922 505
rect -2322 349 -2293 395
rect -2191 349 -2162 395
rect -2322 278 -2162 349
rect 2162 395 2189 2445
rect 2295 395 2322 2445
rect 2162 349 2191 395
rect 2293 349 2322 395
rect 2162 278 2322 349
rect -2322 251 2322 278
rect -2322 145 -2141 251
rect 2141 145 2322 251
rect -2322 118 2322 145
rect -2322 -145 2322 -118
rect -2322 -251 -2141 -145
rect 2141 -251 2322 -145
rect -2322 -278 2322 -251
rect -2322 -349 -2162 -278
rect -2322 -395 -2293 -349
rect -2191 -395 -2162 -349
rect -2322 -2445 -2295 -395
rect -2189 -2445 -2162 -395
rect 2162 -349 2322 -278
rect 2162 -395 2191 -349
rect 2293 -395 2322 -349
rect -1922 -505 1922 -478
rect -1922 -611 -1745 -505
rect 1745 -611 1922 -505
rect -1922 -638 1922 -611
rect -1922 -703 -1762 -638
rect -1922 -735 -1893 -703
rect -1791 -735 -1762 -703
rect -1922 -2065 -1895 -735
rect -1789 -2065 -1762 -735
rect 1762 -703 1922 -638
rect 1762 -735 1791 -703
rect 1893 -735 1922 -703
rect -1603 -1972 -1601 -1938
rect -1567 -1972 -1529 -1938
rect -1495 -1972 -1457 -1938
rect -1423 -1972 -1385 -1938
rect -1351 -1972 -1313 -1938
rect -1279 -1972 -1241 -1938
rect -1207 -1972 -1169 -1938
rect -1135 -1972 -1097 -1938
rect -1063 -1972 -1025 -1938
rect -991 -1972 -953 -1938
rect -919 -1972 -881 -1938
rect -847 -1972 -809 -1938
rect -775 -1972 -737 -1938
rect -703 -1972 -665 -1938
rect -631 -1972 -593 -1938
rect -559 -1972 -521 -1938
rect -487 -1972 -449 -1938
rect -415 -1972 -377 -1938
rect -343 -1972 -305 -1938
rect -271 -1972 -233 -1938
rect -199 -1972 -161 -1938
rect -127 -1972 -89 -1938
rect -55 -1972 -17 -1938
rect 17 -1972 55 -1938
rect 89 -1972 127 -1938
rect 161 -1972 199 -1938
rect 233 -1972 271 -1938
rect 305 -1972 343 -1938
rect 377 -1972 415 -1938
rect 449 -1972 487 -1938
rect 521 -1972 559 -1938
rect 593 -1972 631 -1938
rect 665 -1972 703 -1938
rect 737 -1972 775 -1938
rect 809 -1972 847 -1938
rect 881 -1972 919 -1938
rect 953 -1972 991 -1938
rect 1025 -1972 1063 -1938
rect 1097 -1972 1135 -1938
rect 1169 -1972 1207 -1938
rect 1241 -1972 1279 -1938
rect 1313 -1972 1351 -1938
rect 1385 -1972 1423 -1938
rect 1457 -1972 1495 -1938
rect 1529 -1972 1567 -1938
rect 1601 -1972 1603 -1938
rect -1922 -2097 -1893 -2065
rect -1791 -2097 -1762 -2065
rect -1922 -2162 -1762 -2097
rect 1762 -2065 1789 -735
rect 1895 -2065 1922 -735
rect 1762 -2097 1791 -2065
rect 1893 -2097 1922 -2065
rect 1762 -2162 1922 -2097
rect -1922 -2189 1922 -2162
rect -1922 -2295 -1745 -2189
rect 1745 -2295 1922 -2189
rect -1922 -2322 1922 -2295
rect -2322 -2491 -2293 -2445
rect -2191 -2491 -2162 -2445
rect -2322 -2562 -2162 -2491
rect 2162 -2445 2189 -395
rect 2295 -2445 2322 -395
rect 2162 -2491 2191 -2445
rect 2293 -2491 2322 -2445
rect 2162 -2562 2322 -2491
rect -2322 -2589 2322 -2562
rect -2322 -2695 -2141 -2589
rect 2141 -2695 2322 -2589
rect -2322 -2722 2322 -2695
<< viali >>
rect -2141 2693 2141 2695
rect -2141 2591 -2091 2693
rect -2091 2591 2091 2693
rect 2091 2591 2141 2693
rect -2141 2589 2141 2591
rect -2295 395 -2293 2445
rect -2293 395 -2191 2445
rect -2191 395 -2189 2445
rect -1745 2293 1745 2295
rect -1745 2191 -1683 2293
rect -1683 2191 1683 2293
rect 1683 2191 1745 2293
rect -1745 2189 1745 2191
rect -1895 735 -1893 2065
rect -1893 735 -1791 2065
rect -1791 735 -1789 2065
rect -1601 1947 -1567 1981
rect -1529 1947 -1495 1981
rect -1457 1947 -1423 1981
rect -1385 1947 -1351 1981
rect -1313 1947 -1279 1981
rect -1241 1947 -1207 1981
rect -1169 1947 -1135 1981
rect -1097 1947 -1063 1981
rect -1025 1947 -991 1981
rect -953 1947 -919 1981
rect -881 1947 -847 1981
rect -809 1947 -775 1981
rect -737 1947 -703 1981
rect -665 1947 -631 1981
rect -593 1947 -559 1981
rect -521 1947 -487 1981
rect -449 1947 -415 1981
rect -377 1947 -343 1981
rect -305 1947 -271 1981
rect -233 1947 -199 1981
rect -161 1947 -127 1981
rect -89 1947 -55 1981
rect -17 1947 17 1981
rect 55 1947 89 1981
rect 127 1947 161 1981
rect 199 1947 233 1981
rect 271 1947 305 1981
rect 343 1947 377 1981
rect 415 1947 449 1981
rect 487 1947 521 1981
rect 559 1947 593 1981
rect 631 1947 665 1981
rect 703 1947 737 1981
rect 775 1947 809 1981
rect 847 1947 881 1981
rect 919 1947 953 1981
rect 991 1947 1025 1981
rect 1063 1947 1097 1981
rect 1135 1947 1169 1981
rect 1207 1947 1241 1981
rect 1279 1947 1313 1981
rect 1351 1947 1385 1981
rect 1423 1947 1457 1981
rect 1495 1947 1529 1981
rect 1567 1947 1601 1981
rect 1789 735 1791 2065
rect 1791 735 1893 2065
rect 1893 735 1895 2065
rect -1745 609 1745 611
rect -1745 507 -1683 609
rect -1683 507 1683 609
rect 1683 507 1745 609
rect -1745 505 1745 507
rect 2189 395 2191 2445
rect 2191 395 2293 2445
rect 2293 395 2295 2445
rect -2141 249 2141 251
rect -2141 147 -2091 249
rect -2091 147 2091 249
rect 2091 147 2141 249
rect -2141 145 2141 147
rect -2141 -147 2141 -145
rect -2141 -249 -2091 -147
rect -2091 -249 2091 -147
rect 2091 -249 2141 -147
rect -2141 -251 2141 -249
rect -2295 -2445 -2293 -395
rect -2293 -2445 -2191 -395
rect -2191 -2445 -2189 -395
rect -1745 -507 1745 -505
rect -1745 -609 -1683 -507
rect -1683 -609 1683 -507
rect 1683 -609 1745 -507
rect -1745 -611 1745 -609
rect -1895 -2065 -1893 -735
rect -1893 -2065 -1791 -735
rect -1791 -2065 -1789 -735
rect -1601 -1972 -1567 -1938
rect -1529 -1972 -1495 -1938
rect -1457 -1972 -1423 -1938
rect -1385 -1972 -1351 -1938
rect -1313 -1972 -1279 -1938
rect -1241 -1972 -1207 -1938
rect -1169 -1972 -1135 -1938
rect -1097 -1972 -1063 -1938
rect -1025 -1972 -991 -1938
rect -953 -1972 -919 -1938
rect -881 -1972 -847 -1938
rect -809 -1972 -775 -1938
rect -737 -1972 -703 -1938
rect -665 -1972 -631 -1938
rect -593 -1972 -559 -1938
rect -521 -1972 -487 -1938
rect -449 -1972 -415 -1938
rect -377 -1972 -343 -1938
rect -305 -1972 -271 -1938
rect -233 -1972 -199 -1938
rect -161 -1972 -127 -1938
rect -89 -1972 -55 -1938
rect -17 -1972 17 -1938
rect 55 -1972 89 -1938
rect 127 -1972 161 -1938
rect 199 -1972 233 -1938
rect 271 -1972 305 -1938
rect 343 -1972 377 -1938
rect 415 -1972 449 -1938
rect 487 -1972 521 -1938
rect 559 -1972 593 -1938
rect 631 -1972 665 -1938
rect 703 -1972 737 -1938
rect 775 -1972 809 -1938
rect 847 -1972 881 -1938
rect 919 -1972 953 -1938
rect 991 -1972 1025 -1938
rect 1063 -1972 1097 -1938
rect 1135 -1972 1169 -1938
rect 1207 -1972 1241 -1938
rect 1279 -1972 1313 -1938
rect 1351 -1972 1385 -1938
rect 1423 -1972 1457 -1938
rect 1495 -1972 1529 -1938
rect 1567 -1972 1601 -1938
rect 1789 -2065 1791 -735
rect 1791 -2065 1893 -735
rect 1893 -2065 1895 -735
rect -1745 -2191 1745 -2189
rect -1745 -2293 -1683 -2191
rect -1683 -2293 1683 -2191
rect 1683 -2293 1745 -2191
rect -1745 -2295 1745 -2293
rect 2189 -2445 2191 -395
rect 2191 -2445 2293 -395
rect 2293 -2445 2295 -395
rect -2141 -2591 2141 -2589
rect -2141 -2693 -2091 -2591
rect -2091 -2693 2091 -2591
rect 2091 -2693 2141 -2591
rect -2141 -2695 2141 -2693
<< metal1 >>
rect -2400 3100 2400 3178
rect -2400 2856 -2330 3100
rect 2330 2856 2400 3100
rect -2400 2824 2400 2856
rect -2328 2695 2328 2728
rect -2328 2589 -2141 2695
rect 2141 2589 2328 2695
rect -2328 2460 2328 2589
rect -2328 2445 -2060 2460
rect -2328 395 -2295 2445
rect -2189 395 -2060 2445
rect 2061 2445 2328 2460
rect -2000 2300 2000 2400
rect -2000 2184 -1914 2300
rect 1914 2184 2000 2300
rect -2000 2156 2000 2184
rect -2000 2065 -1756 2156
rect -2000 735 -1895 2065
rect -1789 735 -1756 2065
rect -1603 1987 -1557 2156
rect -1287 1987 -1241 2156
rect -971 1987 -925 2156
rect -655 1987 -609 2156
rect -339 1987 -293 2156
rect -23 1987 23 2156
rect 293 1987 339 2156
rect 609 1987 655 2156
rect 925 1987 971 2156
rect 1241 1987 1287 2156
rect 1557 1987 1603 2156
rect 1756 2065 2000 2156
rect -1615 1981 1615 1987
rect -1615 1947 -1601 1981
rect -1567 1947 -1529 1981
rect -1495 1947 -1457 1981
rect -1423 1947 -1385 1981
rect -1351 1947 -1313 1981
rect -1279 1947 -1241 1981
rect -1207 1947 -1169 1981
rect -1135 1947 -1097 1981
rect -1063 1947 -1025 1981
rect -991 1947 -953 1981
rect -919 1947 -881 1981
rect -847 1947 -809 1981
rect -775 1947 -737 1981
rect -703 1947 -665 1981
rect -631 1947 -593 1981
rect -559 1947 -521 1981
rect -487 1947 -449 1981
rect -415 1947 -377 1981
rect -343 1947 -305 1981
rect -271 1947 -233 1981
rect -199 1947 -161 1981
rect -127 1947 -89 1981
rect -55 1947 -17 1981
rect 17 1947 55 1981
rect 89 1947 127 1981
rect 161 1947 199 1981
rect 233 1947 271 1981
rect 305 1947 343 1981
rect 377 1947 415 1981
rect 449 1947 487 1981
rect 521 1947 559 1981
rect 593 1947 631 1981
rect 665 1947 703 1981
rect 737 1947 775 1981
rect 809 1947 847 1981
rect 881 1947 919 1981
rect 953 1947 991 1981
rect 1025 1947 1063 1981
rect 1097 1947 1135 1981
rect 1169 1947 1207 1981
rect 1241 1947 1279 1981
rect 1313 1947 1351 1981
rect 1385 1947 1423 1981
rect 1457 1947 1495 1981
rect 1529 1947 1567 1981
rect 1601 1947 1615 1981
rect -1615 1941 1615 1947
rect -1603 1900 -1557 1941
rect -1287 1900 -1241 1941
rect -971 1900 -925 1941
rect -655 1900 -609 1941
rect -339 1900 -293 1941
rect -23 1900 23 1941
rect 293 1900 339 1941
rect 609 1900 655 1941
rect 925 1900 971 1941
rect 1241 1900 1287 1941
rect 1557 1900 1603 1941
rect -1445 860 -1399 900
rect -1129 860 -1083 900
rect -813 860 -767 900
rect -497 860 -451 900
rect -181 860 -135 900
rect 135 860 181 900
rect 451 860 497 900
rect 767 860 813 900
rect 1083 860 1129 900
rect 1399 860 1445 900
rect -2000 644 -1756 735
rect -1455 838 1455 860
rect -1455 722 -1431 838
rect -1059 722 1059 838
rect 1431 722 1455 838
rect -1455 700 1455 722
rect 1756 735 1789 2065
rect 1895 735 2000 2065
rect 1756 644 2000 735
rect -2000 616 2000 644
rect -2000 611 53 616
rect 937 611 2000 616
rect -2000 505 -1745 611
rect 1745 505 2000 611
rect -2000 500 53 505
rect 937 500 2000 505
rect -2000 400 2000 500
rect -2328 340 -2060 395
rect 2061 395 2189 2445
rect 2295 395 2328 2445
rect 2061 340 2328 395
rect -2328 256 2328 340
rect -2328 251 -947 256
rect -63 251 2328 256
rect -2328 145 -2141 251
rect 2141 145 2328 251
rect -2328 140 -947 145
rect -63 140 2328 145
rect -2328 40 2328 140
rect -2360 -140 2360 -40
rect -2360 -145 53 -140
rect 937 -145 2360 -140
rect -2360 -251 -2141 -145
rect 2141 -251 2360 -145
rect -2360 -256 53 -251
rect 937 -256 2360 -251
rect -2360 -340 2360 -256
rect -2360 -395 -2060 -340
rect -2360 -2445 -2295 -395
rect -2189 -2445 -2060 -395
rect 2060 -395 2360 -340
rect -2000 -500 2000 -400
rect -2000 -505 -947 -500
rect -63 -505 2000 -500
rect -2000 -611 -1745 -505
rect 1745 -611 2000 -505
rect -2000 -616 -947 -611
rect -63 -616 2000 -611
rect -2000 -644 2000 -616
rect -2000 -735 -1750 -644
rect -2000 -2065 -1895 -735
rect -1789 -2065 -1750 -735
rect -1455 -722 1455 -700
rect -1455 -838 -1431 -722
rect -1059 -838 1059 -722
rect 1431 -838 1455 -722
rect -1455 -860 1455 -838
rect 1756 -735 2000 -644
rect -1445 -900 -1399 -860
rect -1129 -900 -1083 -860
rect -813 -900 -767 -860
rect -497 -900 -451 -860
rect -181 -900 -135 -860
rect 135 -900 181 -860
rect 451 -900 497 -860
rect 767 -900 813 -860
rect 1083 -900 1129 -860
rect 1399 -900 1445 -860
rect -1603 -1932 -1557 -1900
rect -1287 -1932 -1241 -1900
rect -971 -1932 -925 -1900
rect -655 -1932 -609 -1900
rect -339 -1932 -293 -1900
rect -23 -1932 23 -1900
rect 293 -1932 339 -1900
rect 609 -1932 655 -1900
rect 925 -1932 971 -1900
rect 1241 -1932 1287 -1900
rect 1557 -1932 1603 -1900
rect -1615 -1938 1615 -1932
rect -1615 -1972 -1601 -1938
rect -1567 -1972 -1529 -1938
rect -1495 -1972 -1457 -1938
rect -1423 -1972 -1385 -1938
rect -1351 -1972 -1313 -1938
rect -1279 -1972 -1241 -1938
rect -1207 -1972 -1169 -1938
rect -1135 -1972 -1097 -1938
rect -1063 -1972 -1025 -1938
rect -991 -1972 -953 -1938
rect -919 -1972 -881 -1938
rect -847 -1972 -809 -1938
rect -775 -1972 -737 -1938
rect -703 -1972 -665 -1938
rect -631 -1972 -593 -1938
rect -559 -1972 -521 -1938
rect -487 -1972 -449 -1938
rect -415 -1972 -377 -1938
rect -343 -1972 -305 -1938
rect -271 -1972 -233 -1938
rect -199 -1972 -161 -1938
rect -127 -1972 -89 -1938
rect -55 -1972 -17 -1938
rect 17 -1972 55 -1938
rect 89 -1972 127 -1938
rect 161 -1972 199 -1938
rect 233 -1972 271 -1938
rect 305 -1972 343 -1938
rect 377 -1972 415 -1938
rect 449 -1972 487 -1938
rect 521 -1972 559 -1938
rect 593 -1972 631 -1938
rect 665 -1972 703 -1938
rect 737 -1972 775 -1938
rect 809 -1972 847 -1938
rect 881 -1972 919 -1938
rect 953 -1972 991 -1938
rect 1025 -1972 1063 -1938
rect 1097 -1972 1135 -1938
rect 1169 -1972 1207 -1938
rect 1241 -1972 1279 -1938
rect 1313 -1972 1351 -1938
rect 1385 -1972 1423 -1938
rect 1457 -1972 1495 -1938
rect 1529 -1972 1567 -1938
rect 1601 -1972 1615 -1938
rect -1615 -1978 1615 -1972
rect -2000 -2156 -1750 -2065
rect -1603 -2156 -1557 -1978
rect -1287 -2156 -1241 -1978
rect -971 -2156 -925 -1978
rect -655 -2156 -609 -1978
rect -339 -2156 -293 -1978
rect -23 -2156 23 -1978
rect 293 -2156 339 -1978
rect 609 -2156 655 -1978
rect 925 -2156 971 -1978
rect 1241 -2156 1287 -1978
rect 1557 -2156 1603 -1978
rect 1756 -2065 1789 -735
rect 1895 -2065 2000 -735
rect 1756 -2156 2000 -2065
rect -2000 -2184 2000 -2156
rect -2000 -2300 -1914 -2184
rect 1914 -2300 2000 -2184
rect -2000 -2400 2000 -2300
rect -2360 -2460 -2060 -2445
rect 2060 -2445 2189 -395
rect 2295 -2445 2360 -395
rect 2060 -2460 2360 -2445
rect -2360 -2589 2360 -2460
rect -2360 -2695 -2141 -2589
rect 2141 -2695 2360 -2589
rect -2360 -2728 2360 -2695
rect -2400 -2856 2400 -2825
rect -2400 -3100 -2330 -2856
rect 2330 -3100 2400 -2856
rect -2400 -3178 2400 -3100
<< via1 >>
rect -2330 2856 2330 3100
rect -1914 2295 1914 2300
rect -1914 2189 -1745 2295
rect -1745 2189 1745 2295
rect 1745 2189 1914 2295
rect -1914 2184 1914 2189
rect -1431 722 -1059 838
rect 1059 722 1431 838
rect 53 611 937 616
rect 53 505 937 611
rect 53 500 937 505
rect -947 251 -63 256
rect -947 145 -63 251
rect -947 140 -63 145
rect 53 -145 937 -140
rect 53 -251 937 -145
rect 53 -256 937 -251
rect -947 -505 -63 -500
rect -947 -611 -63 -505
rect -947 -616 -63 -611
rect -1431 -838 -1059 -722
rect 1059 -838 1431 -722
rect -1914 -2189 1914 -2184
rect -1914 -2295 -1745 -2189
rect -1745 -2295 1745 -2189
rect 1745 -2295 1914 -2189
rect -1914 -2300 1914 -2295
rect -2330 -3100 2330 -2856
<< metal2 >>
rect -2400 3100 2400 3178
rect -2400 2856 -2330 3100
rect 2330 2856 2400 3100
rect -2400 2300 2400 2856
rect -2400 2184 -1914 2300
rect 1914 2184 2400 2300
rect -2400 2150 2400 2184
rect -1928 2146 1928 2150
rect -1445 838 -1045 870
rect -1445 722 -1431 838
rect -1059 722 -1045 838
rect -1445 284 -1045 722
rect 1045 838 1445 870
rect 1045 722 1059 838
rect 1431 722 1445 838
rect 35 616 955 654
rect 35 500 53 616
rect 937 500 955 616
rect -2400 -284 -1045 284
rect -1445 -722 -1045 -284
rect -965 256 -45 294
rect -965 140 -947 256
rect -63 140 -45 256
rect -965 -500 -45 140
rect 35 -140 955 500
rect 35 -256 53 -140
rect 937 -256 955 -140
rect 35 -294 955 -256
rect 1045 284 1445 722
rect 1045 -284 2400 284
rect -965 -616 -947 -500
rect -63 -616 -45 -500
rect -965 -654 -45 -616
rect -1445 -838 -1431 -722
rect -1059 -838 -1045 -722
rect -1445 -870 -1045 -838
rect 1045 -722 1445 -284
rect 1045 -838 1059 -722
rect 1431 -838 1445 -722
rect 1045 -870 1445 -838
rect -1928 -2150 1928 -2146
rect -2400 -2184 2400 -2150
rect -2400 -2300 -1914 -2184
rect 1914 -2300 2400 -2184
rect -2400 -2856 2400 -2300
rect -2400 -3100 -2330 -2856
rect 2330 -3100 2400 -2856
rect -2400 -3178 2400 -3100
use sky130_fd_pr__pfet_g5v0d10v5_Q5DL9H  xm2
timestamp 1626486988
transform 1 0 0 0 1 1400
box -1645 -600 1645 600
use sky130_fd_pr__nfet_g5v0d10v5_ZGGKXL  xm1
timestamp 1626486988
transform 1 0 0 0 1 -1400
box -1635 -588 1635 588
<< labels >>
flabel metal2 s -2400 -284 -2397 284 3 FreeSans 500 0 0 0 clamp
flabel metal2 s -2392 -2814 -2386 -2808 1 FreeSans 600 0 0 0 VSS
flabel metal2 s -2376 2812 -2370 2816 1 FreeSans 600 0 0 0 VDD
<< properties >>
string FIXED_BBOX -1842 -2242 1842 -558
<< end >>
