magic
tech sky130A
magscale 1 2
timestamp 1623652296
<< nwell >>
rect -3358 -906 2840 2026
rect -3358 -2066 102 -906
<< pwell >>
rect 386 -963 1356 -962
rect 386 -972 1453 -963
rect 1474 -972 2840 -962
rect 386 -2952 2840 -972
<< nmos >>
rect 584 -1932 644 -1732
rect 1130 -1846 1190 -1646
rect 1248 -1846 1308 -1646
rect 1366 -1846 1426 -1646
rect 1484 -1846 1544 -1646
rect 1602 -1846 1662 -1646
rect 1720 -1846 1780 -1646
rect 1838 -1846 1898 -1646
rect 1956 -1846 2016 -1646
rect 2488 -1932 2548 -1732
<< scnmos >>
rect 746 -1119 776 -989
rect 1022 -1119 1052 -989
rect 1261 -1119 1291 -989
rect 1345 -1119 1375 -989
rect 1719 -1119 1749 -989
rect 1803 -1119 1833 -989
rect 2042 -1119 2072 -989
rect 2318 -1119 2348 -989
<< pmos >>
rect -2990 1090 -2590 1290
rect -2532 1090 -2132 1290
rect -2074 1090 -1674 1290
rect -1616 1090 -1216 1290
rect -1158 1090 -758 1290
rect -700 1090 -300 1290
rect 638 690 838 1090
rect 896 690 1096 1090
rect 1154 690 1354 1090
rect 1412 690 1612 1090
rect 1670 690 1870 1090
rect 1928 690 2128 1090
rect 2186 690 2386 1090
rect 638 -170 838 230
rect 896 -170 1096 230
rect 1154 -170 1354 230
rect 1412 -170 1612 230
rect 1670 -170 1870 230
rect 1928 -170 2128 230
rect 2186 -170 2386 230
<< scpmoshvt >>
rect 746 -869 776 -669
rect 1022 -869 1052 -669
rect 1261 -869 1291 -669
rect 1345 -869 1375 -669
rect 1719 -869 1749 -669
rect 1803 -869 1833 -669
rect 2042 -869 2072 -669
rect 2318 -869 2348 -669
<< pmoslvt >>
rect -2931 7 -2731 407
rect -2673 7 -2473 407
rect -2415 7 -2215 407
rect -2157 7 -1957 407
rect -1899 7 -1699 407
rect -1641 7 -1441 407
rect -1383 7 -1183 407
rect -1125 7 -925 407
rect -867 7 -667 407
rect -609 7 -409 407
rect -2931 -853 -2731 -453
rect -2673 -853 -2473 -453
rect -2415 -853 -2215 -453
rect -2157 -853 -1957 -453
rect -1899 -853 -1699 -453
rect -1641 -853 -1441 -453
rect -1383 -853 -1183 -453
rect -1125 -853 -925 -453
rect -867 -853 -667 -453
rect -609 -853 -409 -453
rect -1214 -1824 -1144 -1624
rect -1086 -1824 -1016 -1624
rect -958 -1824 -888 -1624
rect -830 -1824 -760 -1624
rect -702 -1824 -632 -1624
rect -574 -1824 -504 -1624
rect -446 -1824 -376 -1624
rect -318 -1824 -248 -1624
rect -190 -1824 -120 -1624
<< ndiff >>
rect 694 -1001 746 -989
rect 694 -1035 702 -1001
rect 736 -1035 746 -1001
rect 694 -1069 746 -1035
rect 694 -1103 702 -1069
rect 736 -1103 746 -1069
rect 694 -1119 746 -1103
rect 776 -1001 828 -989
rect 776 -1035 786 -1001
rect 820 -1035 828 -1001
rect 776 -1069 828 -1035
rect 776 -1103 786 -1069
rect 820 -1103 828 -1069
rect 776 -1119 828 -1103
rect 970 -1001 1022 -989
rect 970 -1035 978 -1001
rect 1012 -1035 1022 -1001
rect 970 -1069 1022 -1035
rect 970 -1103 978 -1069
rect 1012 -1103 1022 -1069
rect 970 -1119 1022 -1103
rect 1052 -1001 1104 -989
rect 1052 -1035 1062 -1001
rect 1096 -1035 1104 -1001
rect 1052 -1069 1104 -1035
rect 1052 -1103 1062 -1069
rect 1096 -1103 1104 -1069
rect 1052 -1119 1104 -1103
rect 1209 -1005 1261 -989
rect 1209 -1039 1217 -1005
rect 1251 -1039 1261 -1005
rect 1209 -1073 1261 -1039
rect 1209 -1107 1217 -1073
rect 1251 -1107 1261 -1073
rect 1209 -1119 1261 -1107
rect 1291 -1119 1345 -989
rect 1375 -1005 1427 -989
rect 1375 -1039 1385 -1005
rect 1419 -1039 1427 -1005
rect 1375 -1073 1427 -1039
rect 1375 -1107 1385 -1073
rect 1419 -1107 1427 -1073
rect 1375 -1119 1427 -1107
rect 1667 -1005 1719 -989
rect 1667 -1039 1675 -1005
rect 1709 -1039 1719 -1005
rect 1667 -1073 1719 -1039
rect 1667 -1107 1675 -1073
rect 1709 -1107 1719 -1073
rect 1667 -1119 1719 -1107
rect 1749 -1119 1803 -989
rect 1833 -1005 1885 -989
rect 1833 -1039 1843 -1005
rect 1877 -1039 1885 -1005
rect 1833 -1073 1885 -1039
rect 1833 -1107 1843 -1073
rect 1877 -1107 1885 -1073
rect 1833 -1119 1885 -1107
rect 1990 -1001 2042 -989
rect 1990 -1035 1998 -1001
rect 2032 -1035 2042 -1001
rect 1990 -1069 2042 -1035
rect 1990 -1103 1998 -1069
rect 2032 -1103 2042 -1069
rect 1990 -1119 2042 -1103
rect 2072 -1001 2124 -989
rect 2072 -1035 2082 -1001
rect 2116 -1035 2124 -1001
rect 2072 -1069 2124 -1035
rect 2072 -1103 2082 -1069
rect 2116 -1103 2124 -1069
rect 2072 -1119 2124 -1103
rect 2266 -1001 2318 -989
rect 2266 -1035 2274 -1001
rect 2308 -1035 2318 -1001
rect 2266 -1069 2318 -1035
rect 2266 -1103 2274 -1069
rect 2308 -1103 2318 -1069
rect 2266 -1119 2318 -1103
rect 2348 -1001 2400 -989
rect 2348 -1035 2358 -1001
rect 2392 -1035 2400 -1001
rect 2348 -1069 2400 -1035
rect 2348 -1103 2358 -1069
rect 2392 -1103 2400 -1069
rect 2348 -1119 2400 -1103
rect 526 -1744 584 -1732
rect 526 -1920 538 -1744
rect 572 -1920 584 -1744
rect 526 -1932 584 -1920
rect 644 -1744 702 -1732
rect 644 -1920 656 -1744
rect 690 -1920 702 -1744
rect 644 -1932 702 -1920
rect 1072 -1658 1130 -1646
rect 1072 -1834 1084 -1658
rect 1118 -1834 1130 -1658
rect 1072 -1846 1130 -1834
rect 1190 -1658 1248 -1646
rect 1190 -1834 1202 -1658
rect 1236 -1834 1248 -1658
rect 1190 -1846 1248 -1834
rect 1308 -1658 1366 -1646
rect 1308 -1834 1320 -1658
rect 1354 -1834 1366 -1658
rect 1308 -1846 1366 -1834
rect 1426 -1658 1484 -1646
rect 1426 -1834 1438 -1658
rect 1472 -1834 1484 -1658
rect 1426 -1846 1484 -1834
rect 1544 -1658 1602 -1646
rect 1544 -1834 1556 -1658
rect 1590 -1834 1602 -1658
rect 1544 -1846 1602 -1834
rect 1662 -1658 1720 -1646
rect 1662 -1834 1674 -1658
rect 1708 -1834 1720 -1658
rect 1662 -1846 1720 -1834
rect 1780 -1658 1838 -1646
rect 1780 -1834 1792 -1658
rect 1826 -1834 1838 -1658
rect 1780 -1846 1838 -1834
rect 1898 -1658 1956 -1646
rect 1898 -1834 1910 -1658
rect 1944 -1834 1956 -1658
rect 1898 -1846 1956 -1834
rect 2016 -1658 2074 -1646
rect 2016 -1834 2028 -1658
rect 2062 -1834 2074 -1658
rect 2016 -1846 2074 -1834
rect 2430 -1744 2488 -1732
rect 2430 -1920 2442 -1744
rect 2476 -1920 2488 -1744
rect 2430 -1932 2488 -1920
rect 2548 -1744 2606 -1732
rect 2548 -1920 2560 -1744
rect 2594 -1920 2606 -1744
rect 2548 -1932 2606 -1920
<< pdiff >>
rect -3048 1278 -2990 1290
rect -3048 1102 -3036 1278
rect -3002 1102 -2990 1278
rect -3048 1090 -2990 1102
rect -2590 1278 -2532 1290
rect -2590 1102 -2578 1278
rect -2544 1102 -2532 1278
rect -2590 1090 -2532 1102
rect -2132 1278 -2074 1290
rect -2132 1102 -2120 1278
rect -2086 1102 -2074 1278
rect -2132 1090 -2074 1102
rect -1674 1278 -1616 1290
rect -1674 1102 -1662 1278
rect -1628 1102 -1616 1278
rect -1674 1090 -1616 1102
rect -1216 1278 -1158 1290
rect -1216 1102 -1204 1278
rect -1170 1102 -1158 1278
rect -1216 1090 -1158 1102
rect -758 1278 -700 1290
rect -758 1102 -746 1278
rect -712 1102 -700 1278
rect -758 1090 -700 1102
rect -300 1278 -242 1290
rect -300 1102 -288 1278
rect -254 1102 -242 1278
rect -300 1090 -242 1102
rect -2989 395 -2931 407
rect -2989 19 -2977 395
rect -2943 19 -2931 395
rect -2989 7 -2931 19
rect -2731 395 -2673 407
rect -2731 19 -2719 395
rect -2685 19 -2673 395
rect -2731 7 -2673 19
rect -2473 395 -2415 407
rect -2473 19 -2461 395
rect -2427 19 -2415 395
rect -2473 7 -2415 19
rect -2215 395 -2157 407
rect -2215 19 -2203 395
rect -2169 19 -2157 395
rect -2215 7 -2157 19
rect -1957 395 -1899 407
rect -1957 19 -1945 395
rect -1911 19 -1899 395
rect -1957 7 -1899 19
rect -1699 395 -1641 407
rect -1699 19 -1687 395
rect -1653 19 -1641 395
rect -1699 7 -1641 19
rect -1441 395 -1383 407
rect -1441 19 -1429 395
rect -1395 19 -1383 395
rect -1441 7 -1383 19
rect -1183 395 -1125 407
rect -1183 19 -1171 395
rect -1137 19 -1125 395
rect -1183 7 -1125 19
rect -925 395 -867 407
rect -925 19 -913 395
rect -879 19 -867 395
rect -925 7 -867 19
rect -667 395 -609 407
rect -667 19 -655 395
rect -621 19 -609 395
rect -667 7 -609 19
rect -409 395 -351 407
rect -409 19 -397 395
rect -363 19 -351 395
rect -409 7 -351 19
rect -2989 -465 -2931 -453
rect -2989 -841 -2977 -465
rect -2943 -841 -2931 -465
rect -2989 -853 -2931 -841
rect -2731 -465 -2673 -453
rect -2731 -841 -2719 -465
rect -2685 -841 -2673 -465
rect -2731 -853 -2673 -841
rect -2473 -465 -2415 -453
rect -2473 -841 -2461 -465
rect -2427 -841 -2415 -465
rect -2473 -853 -2415 -841
rect -2215 -465 -2157 -453
rect -2215 -841 -2203 -465
rect -2169 -841 -2157 -465
rect -2215 -853 -2157 -841
rect -1957 -465 -1899 -453
rect -1957 -841 -1945 -465
rect -1911 -841 -1899 -465
rect -1957 -853 -1899 -841
rect -1699 -465 -1641 -453
rect -1699 -841 -1687 -465
rect -1653 -841 -1641 -465
rect -1699 -853 -1641 -841
rect -1441 -465 -1383 -453
rect -1441 -841 -1429 -465
rect -1395 -841 -1383 -465
rect -1441 -853 -1383 -841
rect -1183 -465 -1125 -453
rect -1183 -841 -1171 -465
rect -1137 -841 -1125 -465
rect -1183 -853 -1125 -841
rect -925 -465 -867 -453
rect -925 -841 -913 -465
rect -879 -841 -867 -465
rect -925 -853 -867 -841
rect -667 -465 -609 -453
rect -667 -841 -655 -465
rect -621 -841 -609 -465
rect -667 -853 -609 -841
rect -409 -465 -351 -453
rect -409 -841 -397 -465
rect -363 -841 -351 -465
rect -409 -853 -351 -841
rect 580 1078 638 1090
rect 580 702 592 1078
rect 626 702 638 1078
rect 580 690 638 702
rect 838 1078 896 1090
rect 838 702 850 1078
rect 884 702 896 1078
rect 838 690 896 702
rect 1096 1078 1154 1090
rect 1096 702 1108 1078
rect 1142 702 1154 1078
rect 1096 690 1154 702
rect 1354 1078 1412 1090
rect 1354 702 1366 1078
rect 1400 702 1412 1078
rect 1354 690 1412 702
rect 1612 1078 1670 1090
rect 1612 702 1624 1078
rect 1658 702 1670 1078
rect 1612 690 1670 702
rect 1870 1078 1928 1090
rect 1870 702 1882 1078
rect 1916 702 1928 1078
rect 1870 690 1928 702
rect 2128 1078 2186 1090
rect 2128 702 2140 1078
rect 2174 702 2186 1078
rect 2128 690 2186 702
rect 2386 1078 2444 1090
rect 2386 702 2398 1078
rect 2432 702 2444 1078
rect 2386 690 2444 702
rect 580 218 638 230
rect 580 -158 592 218
rect 626 -158 638 218
rect 580 -170 638 -158
rect 838 218 896 230
rect 838 -158 850 218
rect 884 -158 896 218
rect 838 -170 896 -158
rect 1096 218 1154 230
rect 1096 -158 1108 218
rect 1142 -158 1154 218
rect 1096 -170 1154 -158
rect 1354 218 1412 230
rect 1354 -158 1366 218
rect 1400 -158 1412 218
rect 1354 -170 1412 -158
rect 1612 218 1670 230
rect 1612 -158 1624 218
rect 1658 -158 1670 218
rect 1612 -170 1670 -158
rect 1870 218 1928 230
rect 1870 -158 1882 218
rect 1916 -158 1928 218
rect 1870 -170 1928 -158
rect 2128 218 2186 230
rect 2128 -158 2140 218
rect 2174 -158 2186 218
rect 2128 -170 2186 -158
rect 2386 218 2444 230
rect 2386 -158 2398 218
rect 2432 -158 2444 218
rect 2386 -170 2444 -158
rect 694 -681 746 -669
rect 694 -715 702 -681
rect 736 -715 746 -681
rect 694 -749 746 -715
rect 694 -783 702 -749
rect 736 -783 746 -749
rect 694 -817 746 -783
rect 694 -851 702 -817
rect 736 -851 746 -817
rect 694 -869 746 -851
rect 776 -681 828 -669
rect 776 -715 786 -681
rect 820 -715 828 -681
rect 776 -749 828 -715
rect 776 -783 786 -749
rect 820 -783 828 -749
rect 776 -817 828 -783
rect 776 -851 786 -817
rect 820 -851 828 -817
rect 776 -869 828 -851
rect 970 -681 1022 -669
rect 970 -715 978 -681
rect 1012 -715 1022 -681
rect 970 -749 1022 -715
rect 970 -783 978 -749
rect 1012 -783 1022 -749
rect 970 -817 1022 -783
rect 970 -851 978 -817
rect 1012 -851 1022 -817
rect 970 -869 1022 -851
rect 1052 -681 1104 -669
rect 1052 -715 1062 -681
rect 1096 -715 1104 -681
rect 1052 -749 1104 -715
rect 1052 -783 1062 -749
rect 1096 -783 1104 -749
rect 1052 -817 1104 -783
rect 1052 -851 1062 -817
rect 1096 -851 1104 -817
rect 1052 -869 1104 -851
rect 1209 -681 1261 -669
rect 1209 -715 1217 -681
rect 1251 -715 1261 -681
rect 1209 -749 1261 -715
rect 1209 -783 1217 -749
rect 1251 -783 1261 -749
rect 1209 -817 1261 -783
rect 1209 -851 1217 -817
rect 1251 -851 1261 -817
rect 1209 -869 1261 -851
rect 1291 -681 1345 -669
rect 1291 -715 1301 -681
rect 1335 -715 1345 -681
rect 1291 -749 1345 -715
rect 1291 -783 1301 -749
rect 1335 -783 1345 -749
rect 1291 -817 1345 -783
rect 1291 -851 1301 -817
rect 1335 -851 1345 -817
rect 1291 -869 1345 -851
rect 1375 -681 1427 -669
rect 1375 -715 1385 -681
rect 1419 -715 1427 -681
rect 1375 -749 1427 -715
rect 1375 -783 1385 -749
rect 1419 -783 1427 -749
rect 1375 -817 1427 -783
rect 1375 -851 1385 -817
rect 1419 -851 1427 -817
rect 1375 -869 1427 -851
rect 1667 -681 1719 -669
rect 1667 -715 1675 -681
rect 1709 -715 1719 -681
rect 1667 -749 1719 -715
rect 1667 -783 1675 -749
rect 1709 -783 1719 -749
rect 1667 -817 1719 -783
rect 1667 -851 1675 -817
rect 1709 -851 1719 -817
rect 1667 -869 1719 -851
rect 1749 -681 1803 -669
rect 1749 -715 1759 -681
rect 1793 -715 1803 -681
rect 1749 -749 1803 -715
rect 1749 -783 1759 -749
rect 1793 -783 1803 -749
rect 1749 -817 1803 -783
rect 1749 -851 1759 -817
rect 1793 -851 1803 -817
rect 1749 -869 1803 -851
rect 1833 -681 1885 -669
rect 1833 -715 1843 -681
rect 1877 -715 1885 -681
rect 1833 -749 1885 -715
rect 1833 -783 1843 -749
rect 1877 -783 1885 -749
rect 1833 -817 1885 -783
rect 1833 -851 1843 -817
rect 1877 -851 1885 -817
rect 1833 -869 1885 -851
rect 1990 -681 2042 -669
rect 1990 -715 1998 -681
rect 2032 -715 2042 -681
rect 1990 -749 2042 -715
rect 1990 -783 1998 -749
rect 2032 -783 2042 -749
rect 1990 -817 2042 -783
rect 1990 -851 1998 -817
rect 2032 -851 2042 -817
rect 1990 -869 2042 -851
rect 2072 -681 2124 -669
rect 2072 -715 2082 -681
rect 2116 -715 2124 -681
rect 2072 -749 2124 -715
rect 2072 -783 2082 -749
rect 2116 -783 2124 -749
rect 2072 -817 2124 -783
rect 2072 -851 2082 -817
rect 2116 -851 2124 -817
rect 2072 -869 2124 -851
rect 2266 -681 2318 -669
rect 2266 -715 2274 -681
rect 2308 -715 2318 -681
rect 2266 -749 2318 -715
rect 2266 -783 2274 -749
rect 2308 -783 2318 -749
rect 2266 -817 2318 -783
rect 2266 -851 2274 -817
rect 2308 -851 2318 -817
rect 2266 -869 2318 -851
rect 2348 -681 2400 -669
rect 2348 -715 2358 -681
rect 2392 -715 2400 -681
rect 2348 -749 2400 -715
rect 2348 -783 2358 -749
rect 2392 -783 2400 -749
rect 2348 -817 2400 -783
rect 2348 -851 2358 -817
rect 2392 -851 2400 -817
rect 2348 -869 2400 -851
rect -1272 -1636 -1214 -1624
rect -1272 -1812 -1260 -1636
rect -1226 -1812 -1214 -1636
rect -1272 -1824 -1214 -1812
rect -1144 -1636 -1086 -1624
rect -1144 -1812 -1132 -1636
rect -1098 -1812 -1086 -1636
rect -1144 -1824 -1086 -1812
rect -1016 -1636 -958 -1624
rect -1016 -1812 -1004 -1636
rect -970 -1812 -958 -1636
rect -1016 -1824 -958 -1812
rect -888 -1636 -830 -1624
rect -888 -1812 -876 -1636
rect -842 -1812 -830 -1636
rect -888 -1824 -830 -1812
rect -760 -1636 -702 -1624
rect -760 -1812 -748 -1636
rect -714 -1812 -702 -1636
rect -760 -1824 -702 -1812
rect -632 -1636 -574 -1624
rect -632 -1812 -620 -1636
rect -586 -1812 -574 -1636
rect -632 -1824 -574 -1812
rect -504 -1636 -446 -1624
rect -504 -1812 -492 -1636
rect -458 -1812 -446 -1636
rect -504 -1824 -446 -1812
rect -376 -1636 -318 -1624
rect -376 -1812 -364 -1636
rect -330 -1812 -318 -1636
rect -376 -1824 -318 -1812
rect -248 -1636 -190 -1624
rect -248 -1812 -236 -1636
rect -202 -1812 -190 -1636
rect -248 -1824 -190 -1812
rect -120 -1636 -62 -1624
rect -120 -1812 -108 -1636
rect -74 -1812 -62 -1636
rect -120 -1824 -62 -1812
<< ndiffc >>
rect 702 -1035 736 -1001
rect 702 -1103 736 -1069
rect 786 -1035 820 -1001
rect 786 -1103 820 -1069
rect 978 -1035 1012 -1001
rect 978 -1103 1012 -1069
rect 1062 -1035 1096 -1001
rect 1062 -1103 1096 -1069
rect 1217 -1039 1251 -1005
rect 1217 -1107 1251 -1073
rect 1385 -1039 1419 -1005
rect 1385 -1107 1419 -1073
rect 1675 -1039 1709 -1005
rect 1675 -1107 1709 -1073
rect 1843 -1039 1877 -1005
rect 1843 -1107 1877 -1073
rect 1998 -1035 2032 -1001
rect 1998 -1103 2032 -1069
rect 2082 -1035 2116 -1001
rect 2082 -1103 2116 -1069
rect 2274 -1035 2308 -1001
rect 2274 -1103 2308 -1069
rect 2358 -1035 2392 -1001
rect 2358 -1103 2392 -1069
rect 538 -1920 572 -1744
rect 656 -1920 690 -1744
rect 1084 -1834 1118 -1658
rect 1202 -1834 1236 -1658
rect 1320 -1834 1354 -1658
rect 1438 -1834 1472 -1658
rect 1556 -1834 1590 -1658
rect 1674 -1834 1708 -1658
rect 1792 -1834 1826 -1658
rect 1910 -1834 1944 -1658
rect 2028 -1834 2062 -1658
rect 2442 -1920 2476 -1744
rect 2560 -1920 2594 -1744
<< pdiffc >>
rect -3036 1102 -3002 1278
rect -2578 1102 -2544 1278
rect -2120 1102 -2086 1278
rect -1662 1102 -1628 1278
rect -1204 1102 -1170 1278
rect -746 1102 -712 1278
rect -288 1102 -254 1278
rect -2977 19 -2943 395
rect -2719 19 -2685 395
rect -2461 19 -2427 395
rect -2203 19 -2169 395
rect -1945 19 -1911 395
rect -1687 19 -1653 395
rect -1429 19 -1395 395
rect -1171 19 -1137 395
rect -913 19 -879 395
rect -655 19 -621 395
rect -397 19 -363 395
rect -2977 -841 -2943 -465
rect -2719 -841 -2685 -465
rect -2461 -841 -2427 -465
rect -2203 -841 -2169 -465
rect -1945 -841 -1911 -465
rect -1687 -841 -1653 -465
rect -1429 -841 -1395 -465
rect -1171 -841 -1137 -465
rect -913 -841 -879 -465
rect -655 -841 -621 -465
rect -397 -841 -363 -465
rect 592 702 626 1078
rect 850 702 884 1078
rect 1108 702 1142 1078
rect 1366 702 1400 1078
rect 1624 702 1658 1078
rect 1882 702 1916 1078
rect 2140 702 2174 1078
rect 2398 702 2432 1078
rect 592 -158 626 218
rect 850 -158 884 218
rect 1108 -158 1142 218
rect 1366 -158 1400 218
rect 1624 -158 1658 218
rect 1882 -158 1916 218
rect 2140 -158 2174 218
rect 2398 -158 2432 218
rect 702 -715 736 -681
rect 702 -783 736 -749
rect 702 -851 736 -817
rect 786 -715 820 -681
rect 786 -783 820 -749
rect 786 -851 820 -817
rect 978 -715 1012 -681
rect 978 -783 1012 -749
rect 978 -851 1012 -817
rect 1062 -715 1096 -681
rect 1062 -783 1096 -749
rect 1062 -851 1096 -817
rect 1217 -715 1251 -681
rect 1217 -783 1251 -749
rect 1217 -851 1251 -817
rect 1301 -715 1335 -681
rect 1301 -783 1335 -749
rect 1301 -851 1335 -817
rect 1385 -715 1419 -681
rect 1385 -783 1419 -749
rect 1385 -851 1419 -817
rect 1675 -715 1709 -681
rect 1675 -783 1709 -749
rect 1675 -851 1709 -817
rect 1759 -715 1793 -681
rect 1759 -783 1793 -749
rect 1759 -851 1793 -817
rect 1843 -715 1877 -681
rect 1843 -783 1877 -749
rect 1843 -851 1877 -817
rect 1998 -715 2032 -681
rect 1998 -783 2032 -749
rect 1998 -851 2032 -817
rect 2082 -715 2116 -681
rect 2082 -783 2116 -749
rect 2082 -851 2116 -817
rect 2274 -715 2308 -681
rect 2274 -783 2308 -749
rect 2274 -851 2308 -817
rect 2358 -715 2392 -681
rect 2358 -783 2392 -749
rect 2358 -851 2392 -817
rect -1260 -1812 -1226 -1636
rect -1132 -1812 -1098 -1636
rect -1004 -1812 -970 -1636
rect -876 -1812 -842 -1636
rect -748 -1812 -714 -1636
rect -620 -1812 -586 -1636
rect -492 -1812 -458 -1636
rect -364 -1812 -330 -1636
rect -236 -1812 -202 -1636
rect -108 -1812 -74 -1636
<< psubdiff >>
rect 892 -1476 1054 -1376
rect 2038 -1476 2250 -1376
rect 892 -1538 992 -1476
rect 424 -1592 520 -1558
rect 708 -1592 804 -1558
rect 424 -1654 458 -1592
rect 770 -1654 804 -1592
rect 424 -2010 458 -1948
rect 770 -2010 804 -1948
rect 424 -2044 520 -2010
rect 708 -2044 804 -2010
rect 2150 -1540 2250 -1476
rect 892 -2634 992 -2100
rect 2328 -1592 2424 -1558
rect 2612 -1592 2708 -1558
rect 2328 -1654 2362 -1592
rect 2674 -1654 2708 -1592
rect 2328 -2010 2362 -1948
rect 2674 -2010 2708 -1948
rect 2328 -2044 2424 -2010
rect 2612 -2044 2708 -2010
rect 2150 -2634 2250 -2174
rect 892 -2734 1048 -2634
rect 2032 -2734 2250 -2634
<< nsubdiff >>
rect -3322 1890 -3160 1990
rect -120 1890 42 1990
rect -3322 1828 -3222 1890
rect -58 1828 42 1890
rect -3322 -1254 -3222 -1192
rect 380 1890 542 1990
rect 2622 1890 2784 1990
rect 380 1828 480 1890
rect 2684 1828 2784 1890
rect 380 -460 480 -398
rect 2684 -460 2784 -398
rect 380 -560 542 -460
rect 2622 -560 2784 -460
rect -58 -1254 42 -1192
rect -3322 -1354 -3160 -1254
rect -120 -1354 42 -1254
rect -1374 -1448 -1278 -1414
rect -56 -1448 40 -1414
rect -1374 -1608 -1340 -1448
rect -42 -1449 40 -1448
rect 6 -1608 40 -1449
rect -1374 -1996 -1340 -1840
rect 6 -1996 40 -1840
rect -1374 -2030 -1278 -1996
rect -56 -2030 40 -1996
<< psubdiffcont >>
rect 1054 -1476 2038 -1376
rect 520 -1592 708 -1558
rect 424 -1948 458 -1654
rect 770 -1948 804 -1654
rect 520 -2044 708 -2010
rect 892 -2100 992 -1538
rect 2150 -2174 2250 -1540
rect 2424 -1592 2612 -1558
rect 2328 -1948 2362 -1654
rect 2674 -1948 2708 -1654
rect 2424 -2044 2612 -2010
rect 1048 -2734 2032 -2634
<< nsubdiffcont >>
rect -3160 1890 -120 1990
rect -3322 -1192 -3222 1828
rect -58 -1192 42 1828
rect 542 1890 2622 1990
rect 380 -398 480 1828
rect 2684 -398 2784 1828
rect 542 -560 2622 -460
rect -3160 -1354 -120 -1254
rect -1278 -1448 -56 -1414
rect -1374 -1840 -1340 -1608
rect 6 -1840 40 -1608
rect -1278 -2030 -56 -1996
<< poly >>
rect -2916 1371 -2664 1387
rect -2916 1354 -2900 1371
rect -2990 1337 -2900 1354
rect -2680 1354 -2664 1371
rect -2458 1371 -2206 1387
rect -2458 1354 -2442 1371
rect -2680 1337 -2590 1354
rect -2990 1290 -2590 1337
rect -2532 1337 -2442 1354
rect -2222 1354 -2206 1371
rect -2000 1371 -1748 1387
rect -2000 1354 -1984 1371
rect -2222 1337 -2132 1354
rect -2532 1290 -2132 1337
rect -2074 1337 -1984 1354
rect -1764 1354 -1748 1371
rect -1542 1371 -1290 1387
rect -1542 1354 -1526 1371
rect -1764 1337 -1674 1354
rect -2074 1290 -1674 1337
rect -1616 1337 -1526 1354
rect -1306 1354 -1290 1371
rect -1084 1371 -832 1387
rect -1084 1354 -1068 1371
rect -1306 1337 -1216 1354
rect -1616 1290 -1216 1337
rect -1158 1337 -1068 1354
rect -848 1354 -832 1371
rect -626 1371 -374 1387
rect -626 1354 -610 1371
rect -848 1337 -758 1354
rect -1158 1290 -758 1337
rect -700 1337 -610 1354
rect -390 1354 -374 1371
rect -390 1337 -300 1354
rect -700 1290 -300 1337
rect -2990 1043 -2590 1090
rect -2990 1026 -2900 1043
rect -2916 1009 -2900 1026
rect -2680 1026 -2590 1043
rect -2532 1043 -2132 1090
rect -2532 1026 -2442 1043
rect -2680 1009 -2664 1026
rect -2916 993 -2664 1009
rect -2458 1009 -2442 1026
rect -2222 1026 -2132 1043
rect -2074 1043 -1674 1090
rect -2074 1026 -1984 1043
rect -2222 1009 -2206 1026
rect -2458 993 -2206 1009
rect -2000 1009 -1984 1026
rect -1764 1026 -1674 1043
rect -1616 1043 -1216 1090
rect -1616 1026 -1526 1043
rect -1764 1009 -1748 1026
rect -2000 993 -1748 1009
rect -1542 1009 -1526 1026
rect -1306 1026 -1216 1043
rect -1158 1043 -758 1090
rect -1158 1026 -1068 1043
rect -1306 1009 -1290 1026
rect -1542 993 -1290 1009
rect -1084 1009 -1068 1026
rect -848 1026 -758 1043
rect -700 1043 -300 1090
rect -700 1026 -610 1043
rect -848 1009 -832 1026
rect -1084 993 -832 1009
rect -626 1009 -610 1026
rect -390 1026 -300 1043
rect -390 1009 -374 1026
rect -626 993 -374 1009
rect -2897 488 -2765 504
rect -2897 471 -2881 488
rect -2931 454 -2881 471
rect -2781 471 -2765 488
rect -2639 488 -2507 504
rect -2639 471 -2623 488
rect -2781 454 -2731 471
rect -2931 407 -2731 454
rect -2673 454 -2623 471
rect -2523 471 -2507 488
rect -2381 488 -2249 504
rect -2381 471 -2365 488
rect -2523 454 -2473 471
rect -2673 407 -2473 454
rect -2415 454 -2365 471
rect -2265 471 -2249 488
rect -2123 488 -1991 504
rect -2123 471 -2107 488
rect -2265 454 -2215 471
rect -2415 407 -2215 454
rect -2157 454 -2107 471
rect -2007 471 -1991 488
rect -1865 488 -1733 504
rect -1865 471 -1849 488
rect -2007 454 -1957 471
rect -2157 407 -1957 454
rect -1899 454 -1849 471
rect -1749 471 -1733 488
rect -1607 488 -1475 504
rect -1607 471 -1591 488
rect -1749 454 -1699 471
rect -1899 407 -1699 454
rect -1641 454 -1591 471
rect -1491 471 -1475 488
rect -1349 488 -1217 504
rect -1349 471 -1333 488
rect -1491 454 -1441 471
rect -1641 407 -1441 454
rect -1383 454 -1333 471
rect -1233 471 -1217 488
rect -1091 488 -959 504
rect -1091 471 -1075 488
rect -1233 454 -1183 471
rect -1383 407 -1183 454
rect -1125 454 -1075 471
rect -975 471 -959 488
rect -833 488 -701 504
rect -833 471 -817 488
rect -975 454 -925 471
rect -1125 407 -925 454
rect -867 454 -817 471
rect -717 471 -701 488
rect -575 488 -443 504
rect -575 471 -559 488
rect -717 454 -667 471
rect -867 407 -667 454
rect -609 454 -559 471
rect -459 471 -443 488
rect -459 454 -409 471
rect -609 407 -409 454
rect -2931 -40 -2731 7
rect -2931 -57 -2881 -40
rect -2897 -74 -2881 -57
rect -2781 -57 -2731 -40
rect -2673 -40 -2473 7
rect -2673 -57 -2623 -40
rect -2781 -74 -2765 -57
rect -2897 -90 -2765 -74
rect -2639 -74 -2623 -57
rect -2523 -57 -2473 -40
rect -2415 -40 -2215 7
rect -2415 -57 -2365 -40
rect -2523 -74 -2507 -57
rect -2639 -90 -2507 -74
rect -2381 -74 -2365 -57
rect -2265 -57 -2215 -40
rect -2157 -40 -1957 7
rect -2157 -57 -2107 -40
rect -2265 -74 -2249 -57
rect -2381 -90 -2249 -74
rect -2123 -74 -2107 -57
rect -2007 -57 -1957 -40
rect -1899 -40 -1699 7
rect -1899 -57 -1849 -40
rect -2007 -74 -1991 -57
rect -2123 -90 -1991 -74
rect -1865 -74 -1849 -57
rect -1749 -57 -1699 -40
rect -1641 -40 -1441 7
rect -1641 -57 -1591 -40
rect -1749 -74 -1733 -57
rect -1865 -90 -1733 -74
rect -1607 -74 -1591 -57
rect -1491 -57 -1441 -40
rect -1383 -40 -1183 7
rect -1383 -57 -1333 -40
rect -1491 -74 -1475 -57
rect -1607 -90 -1475 -74
rect -1349 -74 -1333 -57
rect -1233 -57 -1183 -40
rect -1125 -40 -925 7
rect -1125 -57 -1075 -40
rect -1233 -74 -1217 -57
rect -1349 -90 -1217 -74
rect -1091 -74 -1075 -57
rect -975 -57 -925 -40
rect -867 -40 -667 7
rect -867 -57 -817 -40
rect -975 -74 -959 -57
rect -1091 -90 -959 -74
rect -833 -74 -817 -57
rect -717 -57 -667 -40
rect -609 -40 -409 7
rect -609 -57 -559 -40
rect -717 -74 -701 -57
rect -833 -90 -701 -74
rect -575 -74 -559 -57
rect -459 -57 -409 -40
rect -459 -74 -443 -57
rect -575 -90 -443 -74
rect -2897 -372 -2765 -356
rect -2897 -389 -2881 -372
rect -2931 -406 -2881 -389
rect -2781 -389 -2765 -372
rect -2639 -372 -2507 -356
rect -2639 -389 -2623 -372
rect -2781 -406 -2731 -389
rect -2931 -453 -2731 -406
rect -2673 -406 -2623 -389
rect -2523 -389 -2507 -372
rect -2381 -372 -2249 -356
rect -2381 -389 -2365 -372
rect -2523 -406 -2473 -389
rect -2673 -453 -2473 -406
rect -2415 -406 -2365 -389
rect -2265 -389 -2249 -372
rect -2123 -372 -1991 -356
rect -2123 -389 -2107 -372
rect -2265 -406 -2215 -389
rect -2415 -453 -2215 -406
rect -2157 -406 -2107 -389
rect -2007 -389 -1991 -372
rect -1865 -372 -1733 -356
rect -1865 -389 -1849 -372
rect -2007 -406 -1957 -389
rect -2157 -453 -1957 -406
rect -1899 -406 -1849 -389
rect -1749 -389 -1733 -372
rect -1607 -372 -1475 -356
rect -1607 -389 -1591 -372
rect -1749 -406 -1699 -389
rect -1899 -453 -1699 -406
rect -1641 -406 -1591 -389
rect -1491 -389 -1475 -372
rect -1349 -372 -1217 -356
rect -1349 -389 -1333 -372
rect -1491 -406 -1441 -389
rect -1641 -453 -1441 -406
rect -1383 -406 -1333 -389
rect -1233 -389 -1217 -372
rect -1091 -372 -959 -356
rect -1091 -389 -1075 -372
rect -1233 -406 -1183 -389
rect -1383 -453 -1183 -406
rect -1125 -406 -1075 -389
rect -975 -389 -959 -372
rect -833 -372 -701 -356
rect -833 -389 -817 -372
rect -975 -406 -925 -389
rect -1125 -453 -925 -406
rect -867 -406 -817 -389
rect -717 -389 -701 -372
rect -575 -372 -443 -356
rect -575 -389 -559 -372
rect -717 -406 -667 -389
rect -867 -453 -667 -406
rect -609 -406 -559 -389
rect -459 -389 -443 -372
rect -459 -406 -409 -389
rect -609 -453 -409 -406
rect -2931 -900 -2731 -853
rect -2931 -917 -2881 -900
rect -2897 -934 -2881 -917
rect -2781 -917 -2731 -900
rect -2673 -900 -2473 -853
rect -2673 -917 -2623 -900
rect -2781 -934 -2765 -917
rect -2897 -950 -2765 -934
rect -2639 -934 -2623 -917
rect -2523 -917 -2473 -900
rect -2415 -900 -2215 -853
rect -2415 -917 -2365 -900
rect -2523 -934 -2507 -917
rect -2639 -950 -2507 -934
rect -2381 -934 -2365 -917
rect -2265 -917 -2215 -900
rect -2157 -900 -1957 -853
rect -2157 -917 -2107 -900
rect -2265 -934 -2249 -917
rect -2381 -950 -2249 -934
rect -2123 -934 -2107 -917
rect -2007 -917 -1957 -900
rect -1899 -900 -1699 -853
rect -1899 -917 -1849 -900
rect -2007 -934 -1991 -917
rect -2123 -950 -1991 -934
rect -1865 -934 -1849 -917
rect -1749 -917 -1699 -900
rect -1641 -900 -1441 -853
rect -1641 -917 -1591 -900
rect -1749 -934 -1733 -917
rect -1865 -950 -1733 -934
rect -1607 -934 -1591 -917
rect -1491 -917 -1441 -900
rect -1383 -900 -1183 -853
rect -1383 -917 -1333 -900
rect -1491 -934 -1475 -917
rect -1607 -950 -1475 -934
rect -1349 -934 -1333 -917
rect -1233 -917 -1183 -900
rect -1125 -900 -925 -853
rect -1125 -917 -1075 -900
rect -1233 -934 -1217 -917
rect -1349 -950 -1217 -934
rect -1091 -934 -1075 -917
rect -975 -917 -925 -900
rect -867 -900 -667 -853
rect -867 -917 -817 -900
rect -975 -934 -959 -917
rect -1091 -950 -959 -934
rect -833 -934 -817 -917
rect -717 -917 -667 -900
rect -609 -900 -409 -853
rect -609 -917 -559 -900
rect -717 -934 -701 -917
rect -833 -950 -701 -934
rect -575 -934 -559 -917
rect -459 -917 -409 -900
rect -459 -934 -443 -917
rect -575 -950 -443 -934
rect 672 1171 804 1187
rect 672 1154 688 1171
rect 638 1137 688 1154
rect 788 1154 804 1171
rect 930 1171 1062 1187
rect 930 1154 946 1171
rect 788 1137 838 1154
rect 638 1090 838 1137
rect 896 1137 946 1154
rect 1046 1154 1062 1171
rect 1188 1171 1320 1187
rect 1188 1154 1204 1171
rect 1046 1137 1096 1154
rect 896 1090 1096 1137
rect 1154 1137 1204 1154
rect 1304 1154 1320 1171
rect 1446 1171 1578 1187
rect 1446 1154 1462 1171
rect 1304 1137 1354 1154
rect 1154 1090 1354 1137
rect 1412 1137 1462 1154
rect 1562 1154 1578 1171
rect 1704 1171 1836 1187
rect 1704 1154 1720 1171
rect 1562 1137 1612 1154
rect 1412 1090 1612 1137
rect 1670 1137 1720 1154
rect 1820 1154 1836 1171
rect 1962 1171 2094 1187
rect 1962 1154 1978 1171
rect 1820 1137 1870 1154
rect 1670 1090 1870 1137
rect 1928 1137 1978 1154
rect 2078 1154 2094 1171
rect 2220 1171 2352 1187
rect 2220 1154 2236 1171
rect 2078 1137 2128 1154
rect 1928 1090 2128 1137
rect 2186 1137 2236 1154
rect 2336 1154 2352 1171
rect 2336 1137 2386 1154
rect 2186 1090 2386 1137
rect 638 643 838 690
rect 638 626 688 643
rect 672 609 688 626
rect 788 626 838 643
rect 896 643 1096 690
rect 896 626 946 643
rect 788 609 804 626
rect 672 593 804 609
rect 930 609 946 626
rect 1046 626 1096 643
rect 1154 643 1354 690
rect 1154 626 1204 643
rect 1046 609 1062 626
rect 930 593 1062 609
rect 1188 609 1204 626
rect 1304 626 1354 643
rect 1412 643 1612 690
rect 1412 626 1462 643
rect 1304 609 1320 626
rect 1188 593 1320 609
rect 1446 609 1462 626
rect 1562 626 1612 643
rect 1670 643 1870 690
rect 1670 626 1720 643
rect 1562 609 1578 626
rect 1446 593 1578 609
rect 1704 609 1720 626
rect 1820 626 1870 643
rect 1928 643 2128 690
rect 1928 626 1978 643
rect 1820 609 1836 626
rect 1704 593 1836 609
rect 1962 609 1978 626
rect 2078 626 2128 643
rect 2186 643 2386 690
rect 2186 626 2236 643
rect 2078 609 2094 626
rect 1962 593 2094 609
rect 2220 609 2236 626
rect 2336 626 2386 643
rect 2336 609 2352 626
rect 2220 593 2352 609
rect 672 311 804 327
rect 672 294 688 311
rect 638 277 688 294
rect 788 294 804 311
rect 930 311 1062 327
rect 930 294 946 311
rect 788 277 838 294
rect 638 230 838 277
rect 896 277 946 294
rect 1046 294 1062 311
rect 1188 311 1320 327
rect 1188 294 1204 311
rect 1046 277 1096 294
rect 896 230 1096 277
rect 1154 277 1204 294
rect 1304 294 1320 311
rect 1446 311 1578 327
rect 1446 294 1462 311
rect 1304 277 1354 294
rect 1154 230 1354 277
rect 1412 277 1462 294
rect 1562 294 1578 311
rect 1704 311 1836 327
rect 1704 294 1720 311
rect 1562 277 1612 294
rect 1412 230 1612 277
rect 1670 277 1720 294
rect 1820 294 1836 311
rect 1962 311 2094 327
rect 1962 294 1978 311
rect 1820 277 1870 294
rect 1670 230 1870 277
rect 1928 277 1978 294
rect 2078 294 2094 311
rect 2220 311 2352 327
rect 2220 294 2236 311
rect 2078 277 2128 294
rect 1928 230 2128 277
rect 2186 277 2236 294
rect 2336 294 2352 311
rect 2336 277 2386 294
rect 2186 230 2386 277
rect 638 -217 838 -170
rect 638 -234 688 -217
rect 672 -251 688 -234
rect 788 -234 838 -217
rect 896 -217 1096 -170
rect 896 -234 946 -217
rect 788 -251 804 -234
rect 672 -267 804 -251
rect 930 -251 946 -234
rect 1046 -234 1096 -217
rect 1154 -217 1354 -170
rect 1154 -234 1204 -217
rect 1046 -251 1062 -234
rect 930 -267 1062 -251
rect 1188 -251 1204 -234
rect 1304 -234 1354 -217
rect 1412 -217 1612 -170
rect 1412 -234 1462 -217
rect 1304 -251 1320 -234
rect 1188 -267 1320 -251
rect 1446 -251 1462 -234
rect 1562 -234 1612 -217
rect 1670 -217 1870 -170
rect 1670 -234 1720 -217
rect 1562 -251 1578 -234
rect 1446 -267 1578 -251
rect 1704 -251 1720 -234
rect 1820 -234 1870 -217
rect 1928 -217 2128 -170
rect 1928 -234 1978 -217
rect 1820 -251 1836 -234
rect 1704 -267 1836 -251
rect 1962 -251 1978 -234
rect 2078 -234 2128 -217
rect 2186 -217 2386 -170
rect 2186 -234 2236 -217
rect 2078 -251 2094 -234
rect 1962 -267 2094 -251
rect 2220 -251 2236 -234
rect 2336 -234 2386 -217
rect 2336 -251 2352 -234
rect 2220 -267 2352 -251
rect 746 -669 776 -643
rect 1022 -669 1052 -643
rect 1261 -669 1291 -643
rect 1345 -669 1375 -643
rect 1719 -669 1749 -643
rect 1803 -669 1833 -643
rect 2042 -669 2072 -643
rect 2318 -669 2348 -643
rect 746 -901 776 -869
rect 1022 -901 1052 -869
rect 1261 -901 1291 -869
rect 690 -917 776 -901
rect 690 -951 706 -917
rect 740 -951 776 -917
rect 690 -967 776 -951
rect 966 -917 1052 -901
rect 966 -951 982 -917
rect 1016 -951 1052 -917
rect 966 -967 1052 -951
rect 1199 -917 1291 -901
rect 1199 -951 1214 -917
rect 1248 -951 1291 -917
rect 1199 -967 1291 -951
rect 746 -989 776 -967
rect 1022 -989 1052 -967
rect 1261 -989 1291 -967
rect 1345 -901 1375 -869
rect 1719 -901 1749 -869
rect 1345 -917 1433 -901
rect 1345 -951 1382 -917
rect 1416 -951 1433 -917
rect 1345 -967 1433 -951
rect 1661 -917 1749 -901
rect 1661 -951 1678 -917
rect 1712 -951 1749 -917
rect 1661 -967 1749 -951
rect 1345 -989 1375 -967
rect 1719 -989 1749 -967
rect 1803 -901 1833 -869
rect 2042 -901 2072 -869
rect 2318 -901 2348 -869
rect 1803 -917 1895 -901
rect 1803 -951 1846 -917
rect 1880 -951 1895 -917
rect 1803 -967 1895 -951
rect 2042 -917 2128 -901
rect 2042 -951 2078 -917
rect 2112 -951 2128 -917
rect 2042 -967 2128 -951
rect 2318 -917 2404 -901
rect 2318 -951 2354 -917
rect 2388 -951 2404 -917
rect 2318 -967 2404 -951
rect 1803 -989 1833 -967
rect 2042 -989 2072 -967
rect 2318 -989 2348 -967
rect 746 -1145 776 -1119
rect 1022 -1145 1052 -1119
rect 1261 -1145 1291 -1119
rect 1345 -1145 1375 -1119
rect 1719 -1145 1749 -1119
rect 1803 -1145 1833 -1119
rect 2042 -1145 2072 -1119
rect 2318 -1145 2348 -1119
rect -1092 -1517 -1010 -1507
rect -1092 -1567 -1076 -1517
rect -1026 -1567 -1010 -1517
rect -1092 -1577 -1010 -1567
rect -964 -1517 -882 -1507
rect -964 -1567 -948 -1517
rect -898 -1567 -882 -1517
rect -964 -1577 -882 -1567
rect -836 -1517 -754 -1507
rect -836 -1567 -820 -1517
rect -770 -1567 -754 -1517
rect -836 -1577 -754 -1567
rect -708 -1517 -626 -1507
rect -708 -1567 -692 -1517
rect -642 -1567 -626 -1517
rect -708 -1577 -626 -1567
rect -580 -1517 -498 -1507
rect -580 -1567 -564 -1517
rect -514 -1567 -498 -1517
rect -580 -1577 -498 -1567
rect -452 -1517 -370 -1507
rect -452 -1567 -436 -1517
rect -386 -1567 -370 -1517
rect -452 -1577 -370 -1567
rect -324 -1517 -242 -1507
rect -324 -1567 -308 -1517
rect -258 -1567 -242 -1517
rect -324 -1577 -242 -1567
rect -1214 -1624 -1144 -1598
rect -1086 -1624 -1016 -1577
rect -958 -1624 -888 -1577
rect -830 -1624 -760 -1577
rect -702 -1624 -632 -1577
rect -574 -1624 -504 -1577
rect -446 -1624 -376 -1577
rect -318 -1624 -248 -1577
rect -190 -1624 -120 -1598
rect -1214 -1869 -1144 -1824
rect -1086 -1850 -1016 -1824
rect -958 -1850 -888 -1824
rect -830 -1850 -760 -1824
rect -702 -1850 -632 -1824
rect -574 -1850 -504 -1824
rect -446 -1850 -376 -1824
rect -318 -1850 -248 -1824
rect -190 -1869 -120 -1824
rect -1220 -1879 -1138 -1869
rect -1220 -1929 -1204 -1879
rect -1154 -1929 -1138 -1879
rect -1220 -1939 -1138 -1929
rect -196 -1879 -114 -1869
rect -196 -1929 -180 -1879
rect -130 -1929 -114 -1879
rect -196 -1939 -114 -1929
rect 581 -1660 647 -1644
rect 581 -1694 597 -1660
rect 631 -1694 647 -1660
rect 581 -1710 647 -1694
rect 584 -1732 644 -1710
rect 584 -1958 644 -1932
rect 1248 -1542 1308 -1526
rect 1248 -1582 1258 -1542
rect 1298 -1582 1308 -1542
rect 1130 -1646 1190 -1620
rect 1248 -1646 1308 -1582
rect 1478 -1542 1550 -1532
rect 1478 -1582 1494 -1542
rect 1534 -1582 1550 -1542
rect 1478 -1592 1550 -1582
rect 1596 -1542 1668 -1532
rect 1596 -1582 1612 -1542
rect 1652 -1582 1668 -1542
rect 1596 -1592 1668 -1582
rect 1832 -1542 1904 -1532
rect 1832 -1582 1848 -1542
rect 1888 -1582 1904 -1542
rect 1832 -1592 1904 -1582
rect 1366 -1646 1426 -1620
rect 1484 -1646 1544 -1592
rect 1602 -1646 1662 -1592
rect 1720 -1646 1780 -1620
rect 1838 -1646 1898 -1592
rect 1956 -1646 2016 -1620
rect 1130 -1896 1190 -1846
rect 1248 -1872 1308 -1846
rect 1064 -1906 1190 -1896
rect 1366 -1898 1426 -1846
rect 1484 -1872 1544 -1846
rect 1602 -1872 1662 -1846
rect 1720 -1898 1780 -1846
rect 1838 -1872 1898 -1846
rect 1956 -1896 2016 -1846
rect 1064 -1946 1080 -1906
rect 1120 -1946 1190 -1906
rect 1064 -1956 1190 -1946
rect 1360 -1908 1432 -1898
rect 1360 -1948 1376 -1908
rect 1416 -1948 1432 -1908
rect 1360 -1958 1432 -1948
rect 1714 -1908 1786 -1898
rect 1714 -1948 1730 -1908
rect 1770 -1948 1786 -1908
rect 1714 -1958 1786 -1948
rect 1956 -1906 2084 -1896
rect 1956 -1946 2028 -1906
rect 2068 -1946 2084 -1906
rect 1956 -1956 2084 -1946
rect 2485 -1660 2551 -1644
rect 2485 -1694 2501 -1660
rect 2535 -1694 2551 -1660
rect 2485 -1710 2551 -1694
rect 2488 -1732 2548 -1710
rect 2488 -1958 2548 -1932
<< polycont >>
rect -2900 1337 -2680 1371
rect -2442 1337 -2222 1371
rect -1984 1337 -1764 1371
rect -1526 1337 -1306 1371
rect -1068 1337 -848 1371
rect -610 1337 -390 1371
rect -2900 1009 -2680 1043
rect -2442 1009 -2222 1043
rect -1984 1009 -1764 1043
rect -1526 1009 -1306 1043
rect -1068 1009 -848 1043
rect -610 1009 -390 1043
rect -2881 454 -2781 488
rect -2623 454 -2523 488
rect -2365 454 -2265 488
rect -2107 454 -2007 488
rect -1849 454 -1749 488
rect -1591 454 -1491 488
rect -1333 454 -1233 488
rect -1075 454 -975 488
rect -817 454 -717 488
rect -559 454 -459 488
rect -2881 -74 -2781 -40
rect -2623 -74 -2523 -40
rect -2365 -74 -2265 -40
rect -2107 -74 -2007 -40
rect -1849 -74 -1749 -40
rect -1591 -74 -1491 -40
rect -1333 -74 -1233 -40
rect -1075 -74 -975 -40
rect -817 -74 -717 -40
rect -559 -74 -459 -40
rect -2881 -406 -2781 -372
rect -2623 -406 -2523 -372
rect -2365 -406 -2265 -372
rect -2107 -406 -2007 -372
rect -1849 -406 -1749 -372
rect -1591 -406 -1491 -372
rect -1333 -406 -1233 -372
rect -1075 -406 -975 -372
rect -817 -406 -717 -372
rect -559 -406 -459 -372
rect -2881 -934 -2781 -900
rect -2623 -934 -2523 -900
rect -2365 -934 -2265 -900
rect -2107 -934 -2007 -900
rect -1849 -934 -1749 -900
rect -1591 -934 -1491 -900
rect -1333 -934 -1233 -900
rect -1075 -934 -975 -900
rect -817 -934 -717 -900
rect -559 -934 -459 -900
rect 688 1137 788 1171
rect 946 1137 1046 1171
rect 1204 1137 1304 1171
rect 1462 1137 1562 1171
rect 1720 1137 1820 1171
rect 1978 1137 2078 1171
rect 2236 1137 2336 1171
rect 688 609 788 643
rect 946 609 1046 643
rect 1204 609 1304 643
rect 1462 609 1562 643
rect 1720 609 1820 643
rect 1978 609 2078 643
rect 2236 609 2336 643
rect 688 277 788 311
rect 946 277 1046 311
rect 1204 277 1304 311
rect 1462 277 1562 311
rect 1720 277 1820 311
rect 1978 277 2078 311
rect 2236 277 2336 311
rect 688 -251 788 -217
rect 946 -251 1046 -217
rect 1204 -251 1304 -217
rect 1462 -251 1562 -217
rect 1720 -251 1820 -217
rect 1978 -251 2078 -217
rect 2236 -251 2336 -217
rect 706 -951 740 -917
rect 982 -951 1016 -917
rect 1214 -951 1248 -917
rect 1382 -951 1416 -917
rect 1678 -951 1712 -917
rect 1846 -951 1880 -917
rect 2078 -951 2112 -917
rect 2354 -951 2388 -917
rect -1076 -1567 -1026 -1517
rect -948 -1567 -898 -1517
rect -820 -1567 -770 -1517
rect -692 -1567 -642 -1517
rect -564 -1567 -514 -1517
rect -436 -1567 -386 -1517
rect -308 -1567 -258 -1517
rect -1204 -1929 -1154 -1879
rect -180 -1929 -130 -1879
rect 597 -1694 631 -1660
rect 1258 -1582 1298 -1542
rect 1494 -1582 1534 -1542
rect 1612 -1582 1652 -1542
rect 1848 -1582 1888 -1542
rect 1080 -1946 1120 -1906
rect 1376 -1948 1416 -1908
rect 1730 -1948 1770 -1908
rect 2028 -1946 2068 -1906
rect 2501 -1694 2535 -1660
<< locali >>
rect -3322 1828 -3222 1990
rect -58 1828 42 1990
rect -2916 1337 -2900 1371
rect -2680 1337 -2664 1371
rect -2458 1337 -2442 1371
rect -2222 1337 -2206 1371
rect -2000 1337 -1984 1371
rect -1764 1337 -1748 1371
rect -1542 1337 -1526 1371
rect -1306 1337 -1290 1371
rect -1084 1337 -1068 1371
rect -848 1337 -832 1371
rect -626 1337 -610 1371
rect -390 1337 -374 1371
rect -3036 1278 -3002 1294
rect -3036 1086 -3002 1102
rect -2578 1278 -2544 1294
rect -2578 1086 -2544 1102
rect -2120 1278 -2086 1294
rect -2120 1086 -2086 1102
rect -1662 1278 -1628 1294
rect -1662 1086 -1628 1102
rect -1204 1278 -1170 1294
rect -1204 1086 -1170 1102
rect -746 1278 -712 1294
rect -746 1086 -712 1102
rect -288 1278 -254 1294
rect -288 1086 -254 1102
rect -2916 1009 -2900 1043
rect -2680 1009 -2664 1043
rect -2458 1009 -2442 1043
rect -2222 1009 -2206 1043
rect -2000 1009 -1984 1043
rect -1764 1009 -1748 1043
rect -1542 1009 -1526 1043
rect -1306 1009 -1290 1043
rect -1084 1009 -1068 1043
rect -848 1009 -832 1043
rect -626 1009 -610 1043
rect -390 1009 -374 1043
rect -2897 454 -2881 488
rect -2781 454 -2765 488
rect -2639 454 -2623 488
rect -2523 454 -2507 488
rect -2381 454 -2365 488
rect -2265 454 -2249 488
rect -2123 454 -2107 488
rect -2007 454 -1991 488
rect -1865 454 -1849 488
rect -1749 454 -1733 488
rect -1607 454 -1591 488
rect -1491 454 -1475 488
rect -1349 454 -1333 488
rect -1233 454 -1217 488
rect -1091 454 -1075 488
rect -975 454 -959 488
rect -833 454 -817 488
rect -717 454 -701 488
rect -575 454 -559 488
rect -459 454 -443 488
rect -2977 395 -2943 411
rect -2977 3 -2943 19
rect -2719 395 -2685 411
rect -2719 3 -2685 19
rect -2461 395 -2427 411
rect -2461 3 -2427 19
rect -2203 395 -2169 411
rect -2203 3 -2169 19
rect -1945 395 -1911 411
rect -1945 3 -1911 19
rect -1687 395 -1653 411
rect -1687 3 -1653 19
rect -1429 395 -1395 411
rect -1429 3 -1395 19
rect -1171 395 -1137 411
rect -1171 3 -1137 19
rect -913 395 -879 411
rect -913 3 -879 19
rect -655 395 -621 411
rect -655 3 -621 19
rect -397 395 -363 411
rect -397 3 -363 19
rect -2897 -74 -2881 -40
rect -2781 -74 -2765 -40
rect -2639 -74 -2623 -40
rect -2523 -74 -2507 -40
rect -2381 -74 -2365 -40
rect -2265 -74 -2249 -40
rect -2123 -74 -2107 -40
rect -2007 -74 -1991 -40
rect -1865 -74 -1849 -40
rect -1749 -74 -1733 -40
rect -1607 -74 -1591 -40
rect -1491 -74 -1475 -40
rect -1349 -74 -1333 -40
rect -1233 -74 -1217 -40
rect -1091 -74 -1075 -40
rect -975 -74 -959 -40
rect -833 -74 -817 -40
rect -717 -74 -701 -40
rect -575 -74 -559 -40
rect -459 -74 -443 -40
rect -2897 -406 -2881 -372
rect -2781 -406 -2765 -372
rect -2639 -406 -2623 -372
rect -2523 -406 -2507 -372
rect -2381 -406 -2365 -372
rect -2265 -406 -2249 -372
rect -2123 -406 -2107 -372
rect -2007 -406 -1991 -372
rect -1865 -406 -1849 -372
rect -1749 -406 -1733 -372
rect -1607 -406 -1591 -372
rect -1491 -406 -1475 -372
rect -1349 -406 -1333 -372
rect -1233 -406 -1217 -372
rect -1091 -406 -1075 -372
rect -975 -406 -959 -372
rect -833 -406 -817 -372
rect -717 -406 -701 -372
rect -575 -406 -559 -372
rect -459 -406 -443 -372
rect -2977 -465 -2943 -449
rect -2977 -857 -2943 -841
rect -2719 -465 -2685 -449
rect -2719 -857 -2685 -841
rect -2461 -465 -2427 -449
rect -2461 -857 -2427 -841
rect -2203 -465 -2169 -449
rect -2203 -857 -2169 -841
rect -1945 -465 -1911 -449
rect -1945 -857 -1911 -841
rect -1687 -465 -1653 -449
rect -1687 -857 -1653 -841
rect -1429 -465 -1395 -449
rect -1429 -857 -1395 -841
rect -1171 -465 -1137 -449
rect -1171 -857 -1137 -841
rect -913 -465 -879 -449
rect -913 -857 -879 -841
rect -655 -465 -621 -449
rect -655 -857 -621 -841
rect -397 -465 -363 -449
rect -397 -857 -363 -841
rect -2897 -934 -2881 -900
rect -2781 -934 -2765 -900
rect -2639 -934 -2623 -900
rect -2523 -934 -2507 -900
rect -2381 -934 -2365 -900
rect -2265 -934 -2249 -900
rect -2123 -934 -2107 -900
rect -2007 -934 -1991 -900
rect -1865 -934 -1849 -900
rect -1749 -934 -1733 -900
rect -1607 -934 -1591 -900
rect -1491 -934 -1475 -900
rect -1349 -934 -1333 -900
rect -1233 -934 -1217 -900
rect -1091 -934 -1075 -900
rect -975 -934 -959 -900
rect -833 -934 -817 -900
rect -717 -934 -701 -900
rect -575 -934 -559 -900
rect -459 -934 -443 -900
rect -3322 -1354 -3222 -1192
rect 380 1828 480 1990
rect 2684 1828 2784 1990
rect 672 1137 688 1171
rect 788 1137 804 1171
rect 930 1137 946 1171
rect 1046 1137 1062 1171
rect 1188 1137 1204 1171
rect 1304 1137 1320 1171
rect 1446 1137 1462 1171
rect 1562 1137 1578 1171
rect 1704 1137 1720 1171
rect 1820 1137 1836 1171
rect 1962 1137 1978 1171
rect 2078 1137 2094 1171
rect 2220 1137 2236 1171
rect 2336 1137 2352 1171
rect 592 1078 626 1094
rect 592 686 626 702
rect 850 1078 884 1094
rect 850 686 884 702
rect 1108 1078 1142 1094
rect 1108 686 1142 702
rect 1366 1078 1400 1094
rect 1366 686 1400 702
rect 1624 1078 1658 1094
rect 1624 686 1658 702
rect 1882 1078 1916 1094
rect 1882 686 1916 702
rect 2140 1078 2174 1094
rect 2140 686 2174 702
rect 2398 1078 2432 1094
rect 2398 686 2432 702
rect 672 609 688 643
rect 788 609 804 643
rect 930 609 946 643
rect 1046 609 1062 643
rect 1188 609 1204 643
rect 1304 609 1320 643
rect 1446 609 1462 643
rect 1562 609 1578 643
rect 1704 609 1720 643
rect 1820 609 1836 643
rect 1962 609 1978 643
rect 2078 609 2094 643
rect 2220 609 2236 643
rect 2336 609 2352 643
rect 672 277 688 311
rect 788 277 804 311
rect 930 277 946 311
rect 1046 277 1062 311
rect 1188 277 1204 311
rect 1304 277 1320 311
rect 1446 277 1462 311
rect 1562 277 1578 311
rect 1704 277 1720 311
rect 1820 277 1836 311
rect 1962 277 1978 311
rect 2078 277 2094 311
rect 2220 277 2236 311
rect 2336 277 2352 311
rect 592 218 626 234
rect 592 -174 626 -158
rect 850 218 884 234
rect 850 -174 884 -158
rect 1108 218 1142 234
rect 1108 -174 1142 -158
rect 1366 218 1400 234
rect 1366 -174 1400 -158
rect 1624 218 1658 234
rect 1624 -174 1658 -158
rect 1882 218 1916 234
rect 1882 -174 1916 -158
rect 2140 218 2174 234
rect 2140 -174 2174 -158
rect 2398 218 2432 234
rect 2398 -174 2432 -158
rect 672 -251 688 -217
rect 788 -251 804 -217
rect 930 -251 946 -217
rect 1046 -251 1062 -217
rect 1188 -251 1204 -217
rect 1304 -251 1320 -217
rect 1446 -251 1462 -217
rect 1562 -251 1578 -217
rect 1704 -251 1720 -217
rect 1820 -251 1836 -217
rect 1962 -251 1978 -217
rect 2078 -251 2094 -217
rect 2220 -251 2236 -217
rect 2336 -251 2352 -217
rect 380 -560 480 -398
rect 2684 -560 2784 -398
rect 626 -639 655 -605
rect 689 -639 747 -605
rect 781 -639 839 -605
rect 873 -639 931 -605
rect 965 -639 1023 -605
rect 1057 -639 1115 -605
rect 1149 -639 1207 -605
rect 1241 -639 1299 -605
rect 1333 -639 1391 -605
rect 1425 -638 1480 -605
rect 1514 -638 1572 -605
rect 1606 -638 1669 -605
rect 1425 -639 1669 -638
rect 1703 -639 1761 -605
rect 1795 -639 1853 -605
rect 1887 -639 1945 -605
rect 1979 -639 2037 -605
rect 2071 -639 2129 -605
rect 2163 -639 2221 -605
rect 2255 -639 2313 -605
rect 2347 -639 2405 -605
rect 2439 -639 2468 -605
rect 694 -681 736 -639
rect 694 -715 702 -681
rect 694 -749 736 -715
rect 694 -783 702 -749
rect 694 -817 736 -783
rect 694 -851 702 -817
rect 694 -867 736 -851
rect 770 -681 836 -673
rect 770 -715 786 -681
rect 820 -715 836 -681
rect 770 -749 836 -715
rect 770 -783 786 -749
rect 820 -783 836 -749
rect 770 -817 836 -783
rect 770 -851 786 -817
rect 820 -851 836 -817
rect 770 -869 836 -851
rect 970 -681 1012 -639
rect 970 -715 978 -681
rect 970 -749 1012 -715
rect 970 -783 978 -749
rect 970 -817 1012 -783
rect 970 -851 978 -817
rect 970 -867 1012 -851
rect 1046 -681 1112 -673
rect 1046 -715 1062 -681
rect 1096 -715 1112 -681
rect 1046 -749 1112 -715
rect 1046 -783 1062 -749
rect 1096 -783 1112 -749
rect 1046 -817 1112 -783
rect 1046 -851 1062 -817
rect 1096 -851 1112 -817
rect 1046 -869 1112 -851
rect 1195 -681 1251 -639
rect 1195 -715 1217 -681
rect 1195 -749 1251 -715
rect 1195 -783 1217 -749
rect 1195 -817 1251 -783
rect 1195 -851 1217 -817
rect 1195 -867 1251 -851
rect 1285 -681 1351 -673
rect 1285 -715 1301 -681
rect 1335 -715 1351 -681
rect 1285 -749 1351 -715
rect 1285 -783 1301 -749
rect 1335 -783 1351 -749
rect 1285 -817 1351 -783
rect 1285 -851 1301 -817
rect 1335 -851 1351 -817
rect 1285 -869 1351 -851
rect 1385 -681 1437 -639
rect 1419 -715 1437 -681
rect 1385 -749 1437 -715
rect 1419 -783 1437 -749
rect 1385 -817 1437 -783
rect 1419 -851 1437 -817
rect 1385 -867 1437 -851
rect 1657 -681 1709 -639
rect 1657 -715 1675 -681
rect 1657 -749 1709 -715
rect 1657 -783 1675 -749
rect 1657 -817 1709 -783
rect 1657 -851 1675 -817
rect 1657 -867 1709 -851
rect 1743 -681 1809 -673
rect 1743 -715 1759 -681
rect 1793 -715 1809 -681
rect 1743 -749 1809 -715
rect 1743 -783 1759 -749
rect 1793 -783 1809 -749
rect 1743 -817 1809 -783
rect 1743 -851 1759 -817
rect 1793 -851 1809 -817
rect 1743 -869 1809 -851
rect 1843 -681 1899 -639
rect 1877 -715 1899 -681
rect 1843 -749 1899 -715
rect 1877 -783 1899 -749
rect 1843 -817 1899 -783
rect 1877 -851 1899 -817
rect 1843 -867 1899 -851
rect 1982 -681 2048 -673
rect 1982 -715 1998 -681
rect 2032 -715 2048 -681
rect 1982 -749 2048 -715
rect 1982 -783 1998 -749
rect 2032 -783 2048 -749
rect 1982 -817 2048 -783
rect 1982 -851 1998 -817
rect 2032 -851 2048 -817
rect 1982 -869 2048 -851
rect 2082 -681 2124 -639
rect 2116 -715 2124 -681
rect 2082 -749 2124 -715
rect 2116 -783 2124 -749
rect 2082 -817 2124 -783
rect 2116 -851 2124 -817
rect 2082 -867 2124 -851
rect 2258 -681 2324 -673
rect 2258 -715 2274 -681
rect 2308 -715 2324 -681
rect 2258 -749 2324 -715
rect 2258 -783 2274 -749
rect 2308 -783 2324 -749
rect 2258 -817 2324 -783
rect 2258 -851 2274 -817
rect 2308 -851 2324 -817
rect 2258 -869 2324 -851
rect 2358 -681 2400 -639
rect 2392 -715 2400 -681
rect 2358 -749 2400 -715
rect 2392 -783 2400 -749
rect 2358 -817 2400 -783
rect 2392 -851 2400 -817
rect 2358 -867 2400 -851
rect 790 -902 836 -869
rect 1066 -902 1112 -869
rect 1197 -902 1264 -901
rect 690 -950 692 -903
rect 690 -951 706 -950
rect 740 -951 756 -903
rect 790 -950 804 -902
rect 1012 -917 1032 -903
rect 690 -1001 736 -985
rect 790 -989 836 -950
rect 966 -951 982 -950
rect 1016 -951 1032 -917
rect 1066 -950 1072 -902
rect 1197 -950 1204 -902
rect 1252 -950 1264 -902
rect 690 -1035 702 -1001
rect 690 -1069 736 -1035
rect 690 -1103 702 -1069
rect 690 -1149 736 -1103
rect 770 -1001 836 -989
rect 770 -1035 786 -1001
rect 820 -1035 836 -1001
rect 770 -1069 836 -1035
rect 770 -1103 786 -1069
rect 820 -1103 836 -1069
rect 770 -1115 836 -1103
rect 966 -1001 1012 -985
rect 1066 -989 1112 -950
rect 1197 -951 1214 -950
rect 1248 -951 1264 -950
rect 1197 -955 1264 -951
rect 1298 -989 1332 -869
rect 1366 -902 1433 -901
rect 1366 -950 1378 -902
rect 1426 -950 1433 -902
rect 1366 -951 1382 -950
rect 1416 -951 1433 -950
rect 1661 -916 1728 -901
rect 1661 -950 1674 -916
rect 1708 -917 1728 -916
rect 1661 -951 1678 -950
rect 1712 -951 1728 -917
rect 1762 -989 1796 -869
rect 1830 -904 1897 -901
rect 1982 -904 2028 -869
rect 2258 -902 2304 -869
rect 1830 -917 1852 -904
rect 1830 -951 1846 -917
rect 1830 -952 1852 -951
rect 2014 -952 2028 -904
rect 2062 -917 2082 -903
rect 2062 -951 2078 -917
rect 2290 -950 2304 -902
rect 2112 -951 2128 -950
rect 1830 -955 1897 -952
rect 1982 -989 2028 -952
rect 966 -1035 978 -1001
rect 966 -1069 1012 -1035
rect 966 -1103 978 -1069
rect 966 -1149 1012 -1103
rect 1046 -1001 1112 -989
rect 1046 -1035 1062 -1001
rect 1096 -1035 1112 -1001
rect 1046 -1069 1112 -1035
rect 1046 -1103 1062 -1069
rect 1096 -1103 1112 -1069
rect 1046 -1115 1112 -1103
rect 1195 -1005 1257 -989
rect 1195 -1039 1217 -1005
rect 1251 -1039 1257 -1005
rect 1195 -1073 1257 -1039
rect 1195 -1107 1217 -1073
rect 1251 -1107 1257 -1073
rect 1195 -1149 1257 -1107
rect 1298 -1005 1437 -989
rect 1298 -1020 1385 -1005
rect 1419 -1020 1437 -1005
rect 1298 -1068 1384 -1020
rect 1432 -1068 1437 -1020
rect 1298 -1073 1437 -1068
rect 1298 -1107 1385 -1073
rect 1419 -1107 1437 -1073
rect 1298 -1115 1437 -1107
rect 1657 -1005 1796 -989
rect 1657 -1020 1675 -1005
rect 1709 -1020 1796 -1005
rect 1657 -1068 1664 -1020
rect 1712 -1068 1796 -1020
rect 1657 -1073 1796 -1068
rect 1657 -1107 1675 -1073
rect 1709 -1107 1796 -1073
rect 1657 -1115 1796 -1107
rect 1837 -1005 1899 -989
rect 1837 -1039 1843 -1005
rect 1877 -1039 1899 -1005
rect 1837 -1073 1899 -1039
rect 1837 -1107 1843 -1073
rect 1877 -1107 1899 -1073
rect 626 -1183 655 -1149
rect 689 -1183 747 -1149
rect 781 -1183 839 -1149
rect 873 -1183 931 -1149
rect 965 -1183 1023 -1149
rect 1057 -1183 1115 -1149
rect 1149 -1183 1207 -1149
rect 1241 -1183 1299 -1149
rect 1333 -1183 1391 -1149
rect 1425 -1150 1572 -1149
rect 1425 -1183 1480 -1150
rect 1514 -1182 1572 -1150
rect 1837 -1149 1899 -1107
rect 1982 -1001 2048 -989
rect 1982 -1035 1998 -1001
rect 2032 -1035 2048 -1001
rect 1982 -1069 2048 -1035
rect 1982 -1103 1998 -1069
rect 2032 -1103 2048 -1069
rect 1982 -1115 2048 -1103
rect 2082 -1001 2128 -985
rect 2116 -1035 2128 -1001
rect 2082 -1069 2128 -1035
rect 2116 -1103 2128 -1069
rect 2082 -1149 2128 -1103
rect 2258 -989 2304 -950
rect 2338 -951 2354 -903
rect 2402 -950 2404 -903
rect 2388 -951 2404 -950
rect 2258 -1001 2324 -989
rect 2258 -1035 2274 -1001
rect 2308 -1035 2324 -1001
rect 2258 -1069 2324 -1035
rect 2258 -1103 2274 -1069
rect 2308 -1103 2324 -1069
rect 2258 -1115 2324 -1103
rect 2358 -1001 2404 -985
rect 2392 -1035 2404 -1001
rect 2358 -1069 2404 -1035
rect 2392 -1103 2404 -1069
rect 2358 -1149 2404 -1103
rect 1606 -1182 1669 -1149
rect 1514 -1183 1669 -1182
rect 1703 -1183 1761 -1149
rect 1795 -1183 1853 -1149
rect 1887 -1183 1945 -1149
rect 1979 -1183 2037 -1149
rect 2071 -1183 2129 -1149
rect 2163 -1183 2221 -1149
rect 2255 -1183 2313 -1149
rect 2347 -1183 2405 -1149
rect 2439 -1183 2468 -1149
rect -58 -1354 42 -1192
rect -1374 -1449 -1278 -1414
rect -1374 -1484 -1340 -1449
rect -54 -1449 40 -1414
rect -1076 -1512 -1026 -1501
rect -948 -1512 -898 -1501
rect -820 -1512 -770 -1501
rect -692 -1507 -642 -1501
rect -564 -1507 -514 -1501
rect -436 -1507 -386 -1501
rect -308 -1507 -258 -1501
rect 6 -1506 40 -1449
rect -702 -1512 -189 -1507
rect -1212 -1517 -189 -1512
rect -1212 -1567 -1076 -1517
rect -1026 -1567 -948 -1517
rect -898 -1567 -820 -1517
rect -770 -1567 -692 -1517
rect -642 -1567 -564 -1517
rect -514 -1567 -436 -1517
rect -386 -1567 -308 -1517
rect -258 -1567 -189 -1517
rect -1212 -1572 -189 -1567
rect -1076 -1583 -1026 -1572
rect -948 -1583 -898 -1572
rect -820 -1583 -770 -1572
rect -702 -1577 -189 -1572
rect -692 -1583 -642 -1577
rect -564 -1583 -514 -1577
rect -436 -1583 -386 -1577
rect -308 -1583 -258 -1577
rect 892 -1517 992 -1376
rect 2150 -1516 2250 -1376
rect 1494 -1532 1652 -1526
rect 1848 -1532 1888 -1526
rect -1260 -1636 -1226 -1620
rect -1277 -1812 -1260 -1785
rect -1132 -1636 -1098 -1620
rect -1226 -1812 -1207 -1785
rect -1277 -1862 -1207 -1812
rect -1132 -1828 -1098 -1812
rect -1004 -1636 -970 -1620
rect -1004 -1828 -970 -1812
rect -876 -1636 -842 -1620
rect -876 -1828 -842 -1812
rect -748 -1636 -714 -1620
rect -748 -1828 -714 -1812
rect -620 -1636 -586 -1620
rect -620 -1828 -586 -1812
rect -492 -1636 -458 -1620
rect -492 -1828 -458 -1812
rect -364 -1636 -330 -1620
rect -364 -1828 -330 -1812
rect -236 -1636 -202 -1620
rect -108 -1636 -74 -1620
rect -236 -1828 -202 -1812
rect -125 -1812 -108 -1791
rect -74 -1812 -55 -1791
rect -125 -1862 -55 -1812
rect -1277 -1863 -1188 -1862
rect -132 -1863 -130 -1862
rect -1204 -1869 -1154 -1863
rect -180 -1869 -130 -1863
rect -1204 -1879 -1144 -1869
rect -1154 -1929 -1144 -1879
rect -1204 -1936 -1144 -1929
rect -1277 -1939 -1144 -1936
rect -190 -1879 -130 -1869
rect -190 -1929 -180 -1879
rect -190 -1937 -130 -1929
rect -190 -1939 -55 -1937
rect -1204 -1945 -1154 -1939
rect -180 -1945 -130 -1939
rect -1374 -1996 -1340 -1952
rect 6 -1996 40 -1952
rect -1374 -2030 -1280 -1996
rect -56 -2030 40 -1996
rect 424 -1592 520 -1558
rect 708 -1592 804 -1558
rect 424 -1654 458 -1592
rect 770 -1654 804 -1592
rect 581 -1694 597 -1660
rect 631 -1694 647 -1660
rect 538 -1744 572 -1728
rect 538 -1936 572 -1920
rect 656 -1744 690 -1728
rect 656 -1936 690 -1920
rect 424 -2010 458 -1948
rect 770 -2010 804 -1948
rect 424 -2044 520 -2010
rect 708 -2044 804 -2010
rect 1484 -1542 1662 -1532
rect 1242 -1582 1248 -1542
rect 1308 -1582 1314 -1542
rect 1484 -1582 1494 -1542
rect 1534 -1582 1612 -1542
rect 1652 -1582 1662 -1542
rect 1484 -1592 1662 -1582
rect 1494 -1598 1652 -1592
rect 1848 -1598 1888 -1592
rect 1084 -1658 1118 -1642
rect 1084 -1850 1118 -1834
rect 1202 -1658 1236 -1642
rect 1202 -1850 1236 -1834
rect 1320 -1658 1354 -1642
rect 1320 -1850 1354 -1834
rect 1438 -1658 1472 -1642
rect 1542 -1658 1602 -1598
rect 1542 -1682 1556 -1658
rect 1438 -1850 1472 -1834
rect 1590 -1682 1602 -1658
rect 1674 -1658 1708 -1642
rect 1556 -1850 1590 -1834
rect 1674 -1850 1708 -1834
rect 1792 -1658 1826 -1642
rect 1792 -1850 1826 -1834
rect 1910 -1658 1944 -1642
rect 1910 -1850 1944 -1834
rect 2028 -1658 2062 -1642
rect 2028 -1850 2062 -1834
rect 1080 -1896 1120 -1890
rect 1376 -1898 1416 -1892
rect 1730 -1898 1770 -1892
rect 2028 -1896 2068 -1890
rect 1366 -1904 1500 -1898
rect 1366 -1908 1446 -1904
rect 1366 -1948 1376 -1908
rect 1416 -1948 1446 -1908
rect 1366 -1952 1446 -1948
rect 1494 -1952 1500 -1904
rect 1080 -1962 1120 -1956
rect 1366 -1958 1500 -1952
rect 1664 -1904 1780 -1898
rect 1664 -1952 1666 -1904
rect 1714 -1908 1780 -1904
rect 1714 -1948 1730 -1908
rect 1770 -1948 1780 -1908
rect 1714 -1952 1780 -1948
rect 1664 -1958 1780 -1952
rect 1376 -1964 1416 -1958
rect 1730 -1964 1770 -1958
rect 2028 -1962 2068 -1956
rect 892 -2734 992 -2593
rect 2328 -1592 2424 -1558
rect 2612 -1592 2708 -1558
rect 2328 -1654 2362 -1592
rect 2674 -1654 2708 -1592
rect 2485 -1694 2501 -1660
rect 2535 -1694 2551 -1660
rect 2442 -1744 2476 -1728
rect 2442 -1936 2476 -1920
rect 2560 -1744 2594 -1728
rect 2560 -1936 2594 -1920
rect 2328 -2010 2362 -1948
rect 2674 -2010 2708 -1948
rect 2328 -2044 2424 -2010
rect 2612 -2044 2708 -2010
rect 2150 -2734 2250 -2593
<< viali >>
rect -3222 1890 -3160 1990
rect -3160 1890 -120 1990
rect -120 1890 -58 1990
rect -3322 -1117 -3222 1753
rect -2882 1337 -2698 1371
rect -2424 1337 -2240 1371
rect -1966 1337 -1782 1371
rect -1508 1337 -1324 1371
rect -1050 1337 -866 1371
rect -592 1337 -408 1371
rect -3036 1102 -3002 1278
rect -2578 1102 -2544 1278
rect -2120 1102 -2086 1278
rect -1662 1102 -1628 1278
rect -1204 1102 -1170 1278
rect -746 1102 -712 1278
rect -288 1102 -254 1278
rect -2882 1009 -2698 1043
rect -2424 1009 -2240 1043
rect -1966 1009 -1782 1043
rect -1508 1009 -1324 1043
rect -1050 1009 -866 1043
rect -592 1009 -408 1043
rect -2873 454 -2789 488
rect -2615 454 -2531 488
rect -2357 454 -2273 488
rect -2099 454 -2015 488
rect -1841 454 -1757 488
rect -1583 454 -1499 488
rect -1325 454 -1241 488
rect -1067 454 -983 488
rect -809 454 -725 488
rect -551 454 -467 488
rect -2977 19 -2943 395
rect -2719 19 -2685 395
rect -2461 19 -2427 395
rect -2203 19 -2169 395
rect -1945 19 -1911 395
rect -1687 19 -1653 395
rect -1429 19 -1395 395
rect -1171 19 -1137 395
rect -913 19 -879 395
rect -655 19 -621 395
rect -397 19 -363 395
rect -2873 -74 -2789 -40
rect -2615 -74 -2531 -40
rect -2357 -74 -2273 -40
rect -2099 -74 -2015 -40
rect -1841 -74 -1757 -40
rect -1583 -74 -1499 -40
rect -1325 -74 -1241 -40
rect -1067 -74 -983 -40
rect -809 -74 -725 -40
rect -551 -74 -467 -40
rect -2873 -406 -2789 -372
rect -2615 -406 -2531 -372
rect -2357 -406 -2273 -372
rect -2099 -406 -2015 -372
rect -1841 -406 -1757 -372
rect -1583 -406 -1499 -372
rect -1325 -406 -1241 -372
rect -1067 -406 -983 -372
rect -809 -406 -725 -372
rect -551 -406 -467 -372
rect -2977 -841 -2943 -465
rect -2719 -841 -2685 -465
rect -2461 -841 -2427 -465
rect -2203 -841 -2169 -465
rect -1945 -841 -1911 -465
rect -1687 -841 -1653 -465
rect -1429 -841 -1395 -465
rect -1171 -841 -1137 -465
rect -913 -841 -879 -465
rect -655 -841 -621 -465
rect -397 -841 -363 -465
rect -2873 -934 -2789 -900
rect -2615 -934 -2531 -900
rect -2357 -934 -2273 -900
rect -2099 -934 -2015 -900
rect -1841 -934 -1757 -900
rect -1583 -934 -1499 -900
rect -1325 -934 -1241 -900
rect -1067 -934 -983 -900
rect -809 -934 -725 -900
rect -551 -934 -467 -900
rect -58 -1117 42 1753
rect 480 1890 542 1990
rect 542 1890 2622 1990
rect 2622 1890 2684 1990
rect 380 -368 480 1798
rect 2688 1564 2784 1798
rect 696 1137 780 1171
rect 954 1137 1038 1171
rect 1212 1137 1296 1171
rect 1470 1137 1554 1171
rect 1728 1137 1812 1171
rect 1986 1137 2070 1171
rect 2244 1137 2328 1171
rect 592 702 626 1078
rect 850 702 884 1078
rect 1108 702 1142 1078
rect 1366 702 1400 1078
rect 1624 702 1658 1078
rect 1882 702 1916 1078
rect 2140 702 2174 1078
rect 2398 702 2432 1078
rect 696 609 780 643
rect 954 609 1038 643
rect 1212 609 1296 643
rect 1470 609 1554 643
rect 1728 609 1812 643
rect 1986 609 2070 643
rect 2244 609 2328 643
rect 696 277 780 311
rect 954 277 1038 311
rect 1212 277 1296 311
rect 1470 277 1554 311
rect 1728 277 1812 311
rect 1986 277 2070 311
rect 2244 277 2328 311
rect 592 -158 626 218
rect 850 -158 884 218
rect 1108 -158 1142 218
rect 1366 -158 1400 218
rect 1624 -158 1658 218
rect 1882 -158 1916 218
rect 2140 -158 2174 218
rect 2398 -158 2432 218
rect 696 -251 780 -217
rect 954 -251 1038 -217
rect 1212 -251 1296 -217
rect 1470 -251 1554 -217
rect 1728 -251 1812 -217
rect 1986 -251 2070 -217
rect 2244 -251 2328 -217
rect 2684 -368 2784 1564
rect 480 -560 542 -460
rect 542 -560 2622 -460
rect 2622 -560 2684 -460
rect 655 -639 689 -605
rect 747 -639 781 -605
rect 839 -639 873 -605
rect 931 -639 965 -605
rect 1023 -639 1057 -605
rect 1115 -639 1149 -605
rect 1207 -639 1241 -605
rect 1299 -639 1333 -605
rect 1391 -639 1425 -605
rect 1480 -638 1514 -604
rect 1572 -638 1606 -604
rect 1669 -639 1703 -605
rect 1761 -639 1795 -605
rect 1853 -639 1887 -605
rect 1945 -639 1979 -605
rect 2037 -639 2071 -605
rect 2129 -639 2163 -605
rect 2221 -639 2255 -605
rect 2313 -639 2347 -605
rect 2405 -639 2439 -605
rect 692 -917 740 -902
rect 692 -950 706 -917
rect 706 -950 740 -917
rect 804 -950 852 -902
rect 964 -917 1012 -902
rect 964 -950 982 -917
rect 982 -950 1012 -917
rect 1072 -950 1120 -902
rect 1204 -917 1252 -902
rect 1204 -950 1214 -917
rect 1214 -950 1248 -917
rect 1248 -950 1252 -917
rect 1378 -917 1426 -902
rect 1378 -950 1382 -917
rect 1382 -950 1416 -917
rect 1416 -950 1426 -917
rect 1674 -917 1708 -916
rect 1674 -950 1678 -917
rect 1678 -950 1708 -917
rect 1852 -917 1900 -904
rect 1852 -951 1880 -917
rect 1880 -951 1900 -917
rect 1852 -952 1900 -951
rect 1966 -952 2014 -904
rect 2082 -917 2130 -902
rect 2082 -950 2112 -917
rect 2112 -950 2130 -917
rect 2242 -950 2290 -902
rect 1384 -1039 1385 -1020
rect 1385 -1039 1419 -1020
rect 1419 -1039 1432 -1020
rect 1384 -1068 1432 -1039
rect 1664 -1039 1675 -1020
rect 1675 -1039 1709 -1020
rect 1709 -1039 1712 -1020
rect 1664 -1068 1712 -1039
rect 655 -1183 689 -1149
rect 747 -1183 781 -1149
rect 839 -1183 873 -1149
rect 931 -1183 965 -1149
rect 1023 -1183 1057 -1149
rect 1115 -1183 1149 -1149
rect 1207 -1183 1241 -1149
rect 1299 -1183 1333 -1149
rect 1391 -1183 1425 -1149
rect 1480 -1184 1514 -1150
rect 1572 -1182 1606 -1148
rect 2354 -917 2402 -902
rect 2354 -950 2388 -917
rect 2388 -950 2402 -917
rect 1669 -1183 1703 -1149
rect 1761 -1183 1795 -1149
rect 1853 -1183 1887 -1149
rect 1945 -1183 1979 -1149
rect 2037 -1183 2071 -1149
rect 2129 -1183 2163 -1149
rect 2221 -1183 2255 -1149
rect 2313 -1183 2347 -1149
rect 2405 -1183 2439 -1149
rect -3222 -1354 -3160 -1254
rect -3160 -1354 -120 -1254
rect -120 -1354 -58 -1254
rect -1278 -1448 -56 -1414
rect -56 -1448 -54 -1414
rect -1278 -1450 -54 -1448
rect -1374 -1608 -1340 -1484
rect -1272 -1572 -1212 -1512
rect -189 -1577 -119 -1507
rect -1374 -1840 -1340 -1608
rect 6 -1608 40 -1506
rect 992 -1476 1054 -1376
rect 1054 -1476 2038 -1376
rect 2038 -1476 2150 -1376
rect 892 -1538 992 -1517
rect -1374 -1952 -1340 -1840
rect -1260 -1812 -1226 -1636
rect -1132 -1812 -1098 -1636
rect -1004 -1812 -970 -1636
rect -876 -1812 -842 -1636
rect -748 -1812 -714 -1636
rect -620 -1812 -586 -1636
rect -492 -1812 -458 -1636
rect -364 -1812 -330 -1636
rect -236 -1812 -202 -1636
rect -108 -1812 -74 -1636
rect -1277 -1936 -1204 -1863
rect -130 -1937 -55 -1862
rect 6 -1840 40 -1608
rect 6 -1952 40 -1840
rect -1280 -2030 -1278 -1996
rect -1278 -2030 -56 -1996
rect 424 -1948 458 -1654
rect 597 -1694 631 -1660
rect 538 -1920 572 -1744
rect 656 -1920 690 -1744
rect 770 -1948 804 -1654
rect 892 -2100 992 -1538
rect 1248 -1542 1308 -1532
rect 1248 -1582 1258 -1542
rect 1258 -1582 1298 -1542
rect 1298 -1582 1308 -1542
rect 1248 -1592 1308 -1582
rect 1838 -1542 1898 -1532
rect 1838 -1582 1848 -1542
rect 1848 -1582 1888 -1542
rect 1888 -1582 1898 -1542
rect 1838 -1592 1898 -1582
rect 2150 -1540 2250 -1516
rect 1084 -1834 1118 -1658
rect 1202 -1834 1236 -1658
rect 1320 -1834 1354 -1658
rect 1438 -1834 1472 -1658
rect 1556 -1834 1590 -1658
rect 1674 -1834 1708 -1658
rect 1792 -1834 1826 -1658
rect 1910 -1834 1944 -1658
rect 2028 -1834 2062 -1658
rect 1070 -1906 1130 -1896
rect 1070 -1946 1080 -1906
rect 1080 -1946 1120 -1906
rect 1120 -1946 1130 -1906
rect 1070 -1956 1130 -1946
rect 1446 -1952 1494 -1904
rect 1666 -1952 1714 -1904
rect 2018 -1906 2078 -1896
rect 2018 -1946 2028 -1906
rect 2028 -1946 2068 -1906
rect 2068 -1946 2078 -1906
rect 2018 -1956 2078 -1946
rect 892 -2593 992 -2100
rect 2150 -2174 2250 -1540
rect 2328 -1948 2362 -1654
rect 2501 -1694 2535 -1660
rect 2442 -1920 2476 -1744
rect 2560 -1920 2594 -1744
rect 2674 -1948 2708 -1654
rect 2150 -2593 2250 -2174
rect 992 -2734 1048 -2634
rect 1048 -2734 2032 -2634
rect 2032 -2734 2150 -2634
<< metal1 >>
rect -3328 1990 48 1996
rect -3328 1890 -3222 1990
rect -58 1890 48 1990
rect -3328 1884 48 1890
rect -3328 1753 -3216 1884
rect -3328 -1117 -3322 1753
rect -3222 1584 -3216 1753
rect -348 1584 -330 1884
rect -3222 1564 -330 1584
rect -64 1753 48 1884
rect -3222 -1117 -3216 1564
rect -3166 710 -3106 1564
rect -2894 1371 -2686 1377
rect -2894 1337 -2882 1371
rect -2698 1337 -2686 1371
rect -2894 1331 -2686 1337
rect -2436 1371 -2228 1377
rect -2436 1337 -2424 1371
rect -2240 1337 -2228 1371
rect -2436 1331 -2228 1337
rect -3042 1278 -2996 1290
rect -3042 1122 -3036 1278
rect -3048 1102 -3036 1122
rect -3002 1122 -2996 1278
rect -2584 1278 -2538 1290
rect -2584 1144 -2578 1278
rect -3002 1102 -2988 1122
rect -3048 836 -2988 1102
rect -2590 1102 -2578 1144
rect -2544 1144 -2538 1278
rect -2134 1278 -2074 1564
rect -1978 1371 -1770 1377
rect -1978 1337 -1966 1371
rect -1782 1337 -1770 1371
rect -1978 1331 -1770 1337
rect -1520 1371 -1312 1377
rect -1520 1337 -1508 1371
rect -1324 1337 -1312 1371
rect -1520 1331 -1312 1337
rect -2134 1242 -2120 1278
rect -2544 1102 -2530 1144
rect -2894 1043 -2686 1049
rect -2894 1009 -2882 1043
rect -2698 1009 -2686 1043
rect -2894 1003 -2686 1009
rect -2820 836 -2760 1003
rect -2590 836 -2530 1102
rect -2126 1102 -2120 1242
rect -2086 1242 -2074 1278
rect -1668 1278 -1622 1290
rect -2086 1102 -2080 1242
rect -1668 1136 -1662 1278
rect -2126 1090 -2080 1102
rect -1676 1102 -1662 1136
rect -1628 1136 -1622 1278
rect -1220 1278 -1160 1564
rect -1062 1371 -854 1377
rect -1062 1337 -1050 1371
rect -866 1337 -854 1371
rect -1062 1331 -854 1337
rect -604 1371 -396 1377
rect -604 1337 -592 1371
rect -408 1337 -396 1371
rect -604 1331 -396 1337
rect -1220 1250 -1204 1278
rect -1628 1102 -1616 1136
rect -2436 1043 -2228 1049
rect -2436 1009 -2424 1043
rect -2240 1009 -2228 1043
rect -2436 1003 -2228 1009
rect -1978 1043 -1770 1049
rect -1978 1009 -1966 1043
rect -1782 1009 -1770 1043
rect -1978 1003 -1770 1009
rect -2364 953 -2304 1003
rect -1908 953 -1848 1003
rect -1676 953 -1616 1102
rect -1210 1102 -1204 1250
rect -1170 1250 -1160 1278
rect -752 1278 -706 1290
rect -1170 1102 -1164 1250
rect -752 1137 -746 1278
rect -1210 1090 -1164 1102
rect -762 1102 -746 1137
rect -712 1137 -706 1278
rect -294 1278 -248 1290
rect -294 1140 -288 1278
rect -712 1102 -702 1137
rect -1520 1043 -1312 1049
rect -1520 1009 -1508 1043
rect -1324 1009 -1312 1043
rect -1520 1003 -1312 1009
rect -1062 1043 -854 1049
rect -1062 1009 -1050 1043
rect -866 1009 -854 1043
rect -1062 1003 -854 1009
rect -1450 953 -1390 1003
rect -986 953 -926 1003
rect -2364 893 -926 953
rect -762 836 -702 1102
rect -304 1102 -288 1140
rect -254 1140 -248 1278
rect -254 1102 -244 1140
rect -604 1043 -396 1049
rect -604 1009 -592 1043
rect -408 1009 -396 1043
rect -604 1003 -396 1009
rect -530 836 -470 1003
rect -304 836 -244 1102
rect -3048 776 -244 836
rect -3166 650 -2802 710
rect -3104 536 -3098 596
rect -3038 536 -3032 596
rect -3098 -992 -3038 536
rect -2990 395 -2930 650
rect -2862 494 -2802 650
rect -2885 488 -2777 494
rect -2885 454 -2873 488
rect -2789 454 -2777 488
rect -2885 448 -2777 454
rect -2627 488 -2519 494
rect -2627 454 -2615 488
rect -2531 454 -2519 488
rect -2627 448 -2519 454
rect -2990 378 -2977 395
rect -2983 50 -2977 378
rect -2986 19 -2977 50
rect -2943 378 -2930 395
rect -2725 395 -2679 407
rect -2943 50 -2937 378
rect -2943 19 -2926 50
rect -2725 38 -2719 395
rect -2986 -192 -2926 19
rect -2730 19 -2719 38
rect -2685 38 -2679 395
rect -2476 395 -2416 776
rect -2220 654 -2214 714
rect -2154 654 -2148 714
rect -2350 536 -2344 596
rect -2284 536 -2278 596
rect -2344 494 -2284 536
rect -2369 488 -2261 494
rect -2369 454 -2357 488
rect -2273 454 -2261 488
rect -2369 448 -2261 454
rect -2685 19 -2670 38
rect -2885 -40 -2777 -34
rect -2885 -74 -2873 -40
rect -2789 -74 -2777 -40
rect -2885 -80 -2777 -74
rect -2862 -192 -2802 -80
rect -2986 -252 -2802 -192
rect -2986 -465 -2926 -252
rect -2862 -366 -2802 -252
rect -2730 -256 -2670 19
rect -2476 19 -2461 395
rect -2427 19 -2416 395
rect -2214 395 -2154 654
rect -2092 536 -2086 596
rect -2026 536 -2020 596
rect -2086 494 -2026 536
rect -2111 488 -2003 494
rect -2111 454 -2099 488
rect -2015 454 -2003 488
rect -2111 448 -2003 454
rect -2214 336 -2203 395
rect -2627 -40 -2519 -34
rect -2627 -74 -2615 -40
rect -2531 -74 -2519 -40
rect -2627 -80 -2519 -74
rect -2600 -136 -2540 -80
rect -2606 -196 -2600 -136
rect -2540 -196 -2534 -136
rect -2736 -316 -2730 -256
rect -2670 -316 -2664 -256
rect -2885 -372 -2777 -366
rect -2885 -406 -2873 -372
rect -2789 -406 -2777 -372
rect -2885 -412 -2777 -406
rect -2627 -372 -2519 -366
rect -2627 -406 -2615 -372
rect -2531 -406 -2519 -372
rect -2627 -412 -2519 -406
rect -2986 -500 -2977 -465
rect -2983 -792 -2977 -500
rect -2990 -841 -2977 -792
rect -2943 -500 -2926 -465
rect -2725 -465 -2679 -453
rect -2943 -792 -2937 -500
rect -2943 -841 -2930 -792
rect -2725 -810 -2719 -465
rect -2990 -988 -2930 -841
rect -2730 -841 -2719 -810
rect -2685 -810 -2679 -465
rect -2476 -465 -2416 19
rect -2209 19 -2203 336
rect -2169 336 -2154 395
rect -1958 395 -1898 776
rect -1853 488 -1745 494
rect -1853 454 -1841 488
rect -1757 454 -1745 488
rect -1853 448 -1745 454
rect -1595 488 -1487 494
rect -1595 454 -1583 488
rect -1499 454 -1487 488
rect -1595 448 -1487 454
rect -2169 19 -2163 336
rect -2209 7 -2163 19
rect -1958 19 -1945 395
rect -1911 19 -1898 395
rect -1693 395 -1647 407
rect -1693 60 -1687 395
rect -2369 -40 -2261 -34
rect -2369 -74 -2357 -40
rect -2273 -74 -2261 -40
rect -2369 -80 -2261 -74
rect -2111 -40 -2003 -34
rect -2111 -74 -2099 -40
rect -2015 -74 -2003 -40
rect -2111 -80 -2003 -74
rect -2352 -196 -2346 -136
rect -2286 -196 -2280 -136
rect -2092 -196 -2086 -136
rect -2026 -196 -2020 -136
rect -2346 -366 -2286 -196
rect -2222 -316 -2216 -256
rect -2156 -316 -2150 -256
rect -2369 -372 -2261 -366
rect -2369 -406 -2357 -372
rect -2273 -406 -2261 -372
rect -2369 -412 -2261 -406
rect -2476 -528 -2461 -465
rect -2685 -841 -2670 -810
rect -2885 -900 -2777 -894
rect -2885 -934 -2873 -900
rect -2789 -934 -2777 -900
rect -2885 -940 -2777 -934
rect -2860 -988 -2800 -940
rect -3104 -1052 -3098 -992
rect -3038 -1052 -3032 -992
rect -2990 -1048 -2800 -988
rect -2730 -1026 -2670 -841
rect -2467 -841 -2461 -528
rect -2427 -528 -2416 -465
rect -2216 -465 -2156 -316
rect -2086 -366 -2026 -196
rect -2111 -372 -2003 -366
rect -2111 -406 -2099 -372
rect -2015 -406 -2003 -372
rect -2111 -412 -2003 -406
rect -2216 -502 -2203 -465
rect -2427 -841 -2421 -528
rect -2467 -853 -2421 -841
rect -2209 -841 -2203 -502
rect -2169 -502 -2156 -465
rect -1958 -465 -1898 19
rect -1700 19 -1687 60
rect -1653 60 -1647 395
rect -1442 395 -1382 776
rect -1190 654 -1184 714
rect -1124 654 -1118 714
rect -1318 536 -1312 596
rect -1252 536 -1246 596
rect -1312 494 -1252 536
rect -1337 488 -1229 494
rect -1337 454 -1325 488
rect -1241 454 -1229 488
rect -1337 448 -1229 454
rect -1653 19 -1640 60
rect -1853 -40 -1745 -34
rect -1853 -74 -1841 -40
rect -1757 -74 -1745 -40
rect -1853 -80 -1745 -74
rect -1828 -136 -1768 -80
rect -1834 -196 -1828 -136
rect -1768 -196 -1762 -136
rect -1700 -256 -1640 19
rect -1442 19 -1429 395
rect -1395 19 -1382 395
rect -1184 395 -1124 654
rect -1058 536 -1052 596
rect -992 536 -986 596
rect -1052 494 -992 536
rect -1079 488 -971 494
rect -1079 454 -1067 488
rect -983 454 -971 488
rect -1079 448 -971 454
rect -1184 364 -1171 395
rect -1595 -40 -1487 -34
rect -1595 -74 -1583 -40
rect -1499 -74 -1487 -40
rect -1595 -80 -1487 -74
rect -1570 -136 -1510 -80
rect -1576 -196 -1570 -136
rect -1510 -196 -1504 -136
rect -1706 -316 -1700 -256
rect -1640 -316 -1634 -256
rect -1853 -372 -1745 -366
rect -1853 -406 -1841 -372
rect -1757 -406 -1745 -372
rect -1853 -412 -1745 -406
rect -1595 -372 -1487 -366
rect -1595 -406 -1583 -372
rect -1499 -406 -1487 -372
rect -1595 -412 -1487 -406
rect -2169 -841 -2163 -502
rect -1958 -516 -1945 -465
rect -2209 -853 -2163 -841
rect -1951 -841 -1945 -516
rect -1911 -516 -1898 -465
rect -1693 -465 -1647 -453
rect -1911 -841 -1905 -516
rect -1693 -792 -1687 -465
rect -1951 -853 -1905 -841
rect -1700 -841 -1687 -792
rect -1653 -792 -1647 -465
rect -1442 -465 -1382 19
rect -1177 19 -1171 364
rect -1137 364 -1124 395
rect -928 395 -868 776
rect -298 654 -292 714
rect -232 654 -226 714
rect -538 536 -474 596
rect -414 536 -350 596
rect -538 494 -478 536
rect -821 488 -713 494
rect -821 454 -809 488
rect -725 454 -713 488
rect -821 448 -713 454
rect -563 488 -455 494
rect -563 454 -551 488
rect -467 454 -455 488
rect -563 448 -455 454
rect -1137 19 -1131 364
rect -1177 7 -1131 19
rect -928 19 -913 395
rect -879 19 -868 395
rect -661 395 -615 407
rect -661 84 -655 395
rect -1337 -40 -1229 -34
rect -1337 -74 -1325 -40
rect -1241 -74 -1229 -40
rect -1337 -80 -1229 -74
rect -1079 -40 -971 -34
rect -1079 -74 -1067 -40
rect -983 -74 -971 -40
rect -1079 -80 -971 -74
rect -1318 -196 -1312 -136
rect -1252 -196 -1246 -136
rect -1060 -196 -1054 -136
rect -994 -196 -988 -136
rect -1312 -366 -1252 -196
rect -1190 -316 -1184 -256
rect -1124 -316 -1118 -256
rect -1337 -372 -1229 -366
rect -1337 -406 -1325 -372
rect -1241 -406 -1229 -372
rect -1337 -412 -1229 -406
rect -1442 -526 -1429 -465
rect -1653 -841 -1640 -792
rect -2627 -900 -2519 -894
rect -2627 -934 -2615 -900
rect -2531 -934 -2519 -900
rect -2627 -940 -2519 -934
rect -2369 -900 -2261 -894
rect -2369 -934 -2357 -900
rect -2273 -934 -2261 -900
rect -2369 -940 -2261 -934
rect -2111 -900 -2003 -894
rect -2111 -934 -2099 -900
rect -2015 -934 -2003 -900
rect -2111 -940 -2003 -934
rect -1853 -900 -1745 -894
rect -1853 -934 -1841 -900
rect -1757 -934 -1745 -900
rect -1853 -940 -1745 -934
rect -2604 -992 -2544 -940
rect -1828 -992 -1768 -940
rect -2732 -1108 -2670 -1026
rect -2610 -1052 -2604 -992
rect -2544 -1052 -2538 -992
rect -1834 -1052 -1828 -992
rect -1768 -1052 -1762 -992
rect -3328 -1248 -3216 -1117
rect -2738 -1168 -2732 -1108
rect -2672 -1168 -2666 -1108
rect -1700 -1110 -1640 -841
rect -1435 -841 -1429 -526
rect -1395 -526 -1382 -465
rect -1184 -465 -1124 -316
rect -1054 -366 -994 -196
rect -1079 -372 -971 -366
rect -1079 -406 -1067 -372
rect -983 -406 -971 -372
rect -1079 -412 -971 -406
rect -1184 -516 -1171 -465
rect -1395 -841 -1389 -526
rect -1435 -853 -1389 -841
rect -1177 -841 -1171 -516
rect -1137 -516 -1124 -465
rect -928 -465 -868 19
rect -672 19 -655 84
rect -621 84 -615 395
rect -410 395 -350 536
rect -410 352 -397 395
rect -621 19 -612 84
rect -403 64 -397 352
rect -821 -40 -713 -34
rect -821 -74 -809 -40
rect -725 -74 -713 -40
rect -821 -80 -713 -74
rect -796 -136 -736 -80
rect -802 -196 -796 -136
rect -736 -196 -730 -136
rect -672 -256 -612 19
rect -410 19 -397 64
rect -363 352 -350 395
rect -363 64 -357 352
rect -363 19 -350 64
rect -563 -40 -455 -34
rect -563 -74 -551 -40
rect -467 -74 -455 -40
rect -563 -80 -455 -74
rect -538 -198 -478 -80
rect -410 -198 -350 19
rect -678 -316 -672 -256
rect -612 -316 -606 -256
rect -538 -258 -350 -198
rect -538 -366 -478 -258
rect -821 -372 -713 -366
rect -821 -406 -809 -372
rect -725 -406 -713 -372
rect -821 -412 -713 -406
rect -563 -372 -455 -366
rect -563 -406 -551 -372
rect -467 -406 -455 -372
rect -563 -412 -455 -406
rect -1137 -841 -1131 -516
rect -928 -526 -913 -465
rect -1177 -853 -1131 -841
rect -919 -841 -913 -526
rect -879 -526 -868 -465
rect -661 -465 -615 -453
rect -879 -841 -873 -526
rect -661 -798 -655 -465
rect -919 -853 -873 -841
rect -670 -841 -655 -798
rect -621 -798 -615 -465
rect -410 -465 -350 -258
rect -410 -504 -397 -465
rect -621 -841 -610 -798
rect -403 -800 -397 -504
rect -1595 -900 -1487 -894
rect -1595 -934 -1583 -900
rect -1499 -934 -1487 -900
rect -1595 -940 -1487 -934
rect -1337 -900 -1229 -894
rect -1337 -934 -1325 -900
rect -1241 -934 -1229 -900
rect -1337 -940 -1229 -934
rect -1079 -900 -971 -894
rect -1079 -934 -1067 -900
rect -983 -934 -971 -900
rect -1079 -940 -971 -934
rect -821 -900 -713 -894
rect -821 -934 -809 -900
rect -725 -934 -713 -900
rect -821 -940 -713 -934
rect -1572 -992 -1512 -940
rect -800 -992 -740 -940
rect -1578 -1052 -1572 -992
rect -1512 -1052 -1506 -992
rect -806 -1052 -800 -992
rect -740 -1052 -734 -992
rect -1700 -1176 -1640 -1170
rect -670 -1110 -610 -841
rect -412 -841 -397 -800
rect -363 -504 -350 -465
rect -363 -800 -357 -504
rect -363 -841 -352 -800
rect -563 -900 -455 -894
rect -563 -934 -551 -900
rect -467 -934 -455 -900
rect -563 -940 -455 -934
rect -538 -990 -478 -940
rect -412 -990 -352 -841
rect -538 -1050 -352 -990
rect -670 -1176 -610 -1170
rect -292 -1110 -232 654
rect -292 -1176 -232 -1170
rect -64 -1117 -58 1753
rect 42 -1117 48 1753
rect 374 1990 2790 1996
rect 374 1890 480 1990
rect 2684 1890 2790 1990
rect 374 1884 2790 1890
rect 374 1798 486 1884
rect 248 366 254 426
rect 314 366 320 426
rect 102 -316 108 -256
rect 168 -316 174 -256
rect -64 -1248 48 -1117
rect -3328 -1254 48 -1248
rect -3328 -1354 -3222 -1254
rect -58 -1354 48 -1254
rect -3328 -1360 48 -1354
rect -1570 -1458 -1564 -1398
rect -1504 -1458 -1498 -1398
rect -1388 -1414 48 -1360
rect -1388 -1450 -1278 -1414
rect -54 -1450 48 -1414
rect -1564 -2076 -1504 -1458
rect -1388 -1462 48 -1450
rect -1388 -1484 -1330 -1462
rect -1388 -1952 -1374 -1484
rect -1340 -1952 -1330 -1484
rect -1278 -1506 -1206 -1500
rect -1284 -1578 -1278 -1506
rect -1218 -1512 -1206 -1506
rect -1212 -1572 -1206 -1512
rect -1218 -1578 -1206 -1572
rect -1278 -1584 -1206 -1578
rect -195 -1501 -113 -1495
rect -195 -1507 -183 -1501
rect -195 -1577 -189 -1507
rect -195 -1583 -183 -1577
rect -113 -1583 -107 -1501
rect -10 -1506 48 -1462
rect -195 -1589 -113 -1583
rect -1266 -1636 -1220 -1624
rect -1266 -1786 -1260 -1636
rect -1276 -1812 -1260 -1786
rect -1226 -1786 -1220 -1636
rect -1138 -1636 -1092 -1624
rect -1138 -1766 -1132 -1636
rect -1098 -1766 -1092 -1636
rect -1010 -1636 -964 -1624
rect -1010 -1732 -1004 -1636
rect -1226 -1812 -1203 -1786
rect -1276 -1857 -1203 -1812
rect -1152 -1826 -1146 -1766
rect -1086 -1826 -1080 -1766
rect -1016 -1812 -1004 -1732
rect -970 -1732 -964 -1636
rect -882 -1636 -836 -1624
rect -970 -1812 -956 -1732
rect -882 -1756 -876 -1636
rect -842 -1756 -836 -1636
rect -754 -1636 -708 -1624
rect -1289 -1863 -1192 -1857
rect -1289 -1936 -1277 -1863
rect -1204 -1936 -1192 -1863
rect -1016 -1874 -956 -1812
rect -896 -1816 -890 -1756
rect -830 -1816 -824 -1756
rect -754 -1788 -748 -1636
rect -762 -1812 -748 -1788
rect -714 -1788 -708 -1636
rect -626 -1636 -580 -1624
rect -626 -1746 -620 -1636
rect -586 -1746 -580 -1636
rect -498 -1636 -452 -1624
rect -714 -1812 -702 -1788
rect -638 -1806 -632 -1746
rect -572 -1806 -566 -1746
rect -498 -1774 -492 -1636
rect -882 -1824 -836 -1816
rect -762 -1874 -702 -1812
rect -626 -1812 -620 -1806
rect -586 -1812 -580 -1806
rect -626 -1824 -580 -1812
rect -506 -1812 -492 -1774
rect -458 -1774 -452 -1636
rect -370 -1636 -324 -1624
rect -370 -1748 -364 -1636
rect -330 -1748 -324 -1636
rect -242 -1636 -196 -1624
rect -242 -1746 -236 -1636
rect -202 -1746 -196 -1636
rect -114 -1636 -68 -1624
rect -458 -1812 -446 -1774
rect -386 -1808 -380 -1748
rect -320 -1808 -314 -1748
rect -252 -1806 -246 -1746
rect -186 -1806 -180 -1746
rect -114 -1759 -108 -1636
rect -506 -1874 -446 -1812
rect -370 -1812 -364 -1808
rect -330 -1812 -324 -1808
rect -370 -1824 -324 -1812
rect -250 -1812 -236 -1806
rect -202 -1812 -190 -1806
rect -250 -1874 -190 -1812
rect -129 -1812 -108 -1759
rect -74 -1759 -68 -1636
rect -74 -1812 -54 -1759
rect -129 -1856 -54 -1812
rect -1016 -1934 -190 -1874
rect -142 -1862 -43 -1856
rect -1289 -1942 -1192 -1936
rect -142 -1937 -130 -1862
rect -55 -1937 -43 -1862
rect -1388 -1979 -1330 -1952
rect -1276 -1979 -1203 -1942
rect -142 -1943 -43 -1937
rect -129 -1979 -54 -1943
rect -10 -1952 6 -1506
rect 40 -1952 48 -1506
rect -10 -1979 48 -1952
rect -1388 -1996 48 -1979
rect -1388 -2030 -1280 -1996
rect -56 -2030 48 -1996
rect -1388 -2038 48 -2030
rect -380 -2076 -320 -2070
rect -1564 -2078 -890 -2076
rect -1564 -2136 -1146 -2078
rect -1152 -2138 -1146 -2136
rect -1086 -2136 -890 -2078
rect -830 -2136 -632 -2076
rect -572 -2136 -380 -2076
rect -1086 -2138 -1080 -2136
rect -380 -2142 -320 -2136
rect 108 -2096 168 -316
rect 254 -896 314 366
rect 374 -368 380 1798
rect 480 -368 486 1798
rect 1038 1584 1056 1884
rect 2676 1798 2790 1884
rect 2676 1584 2688 1798
rect 1038 1564 2688 1584
rect 1090 1414 1150 1564
rect 578 1354 1150 1414
rect 578 1078 638 1354
rect 708 1177 768 1354
rect 834 1244 840 1304
rect 900 1244 906 1304
rect 684 1171 792 1177
rect 684 1137 696 1171
rect 780 1137 792 1171
rect 684 1131 792 1137
rect 578 1024 592 1078
rect 586 850 592 1024
rect 374 -454 486 -368
rect 574 702 592 850
rect 626 1024 638 1078
rect 840 1078 900 1244
rect 942 1171 1050 1177
rect 942 1137 954 1171
rect 1038 1137 1050 1171
rect 942 1131 1050 1137
rect 840 1038 850 1078
rect 626 850 632 1024
rect 626 702 634 850
rect 574 492 634 702
rect 844 702 850 1038
rect 884 1038 900 1078
rect 1090 1078 1150 1354
rect 1220 1244 1226 1304
rect 1286 1244 1292 1304
rect 1478 1244 1484 1304
rect 1544 1244 1550 1304
rect 1226 1177 1286 1244
rect 1484 1177 1544 1244
rect 1200 1171 1308 1177
rect 1200 1137 1212 1171
rect 1296 1137 1308 1171
rect 1200 1131 1308 1137
rect 1458 1171 1566 1177
rect 1458 1137 1470 1171
rect 1554 1137 1566 1171
rect 1458 1131 1566 1137
rect 884 702 890 1038
rect 844 690 890 702
rect 1090 702 1108 1078
rect 1142 702 1150 1078
rect 1360 1078 1406 1090
rect 1360 746 1366 1078
rect 684 643 792 649
rect 684 609 696 643
rect 780 609 792 643
rect 684 603 792 609
rect 942 643 1050 649
rect 942 609 954 643
rect 1038 609 1050 643
rect 942 603 1050 609
rect 708 492 768 603
rect 574 432 768 492
rect 574 218 634 432
rect 708 317 768 432
rect 964 426 1024 603
rect 834 366 840 426
rect 900 366 906 426
rect 958 366 964 426
rect 1024 366 1030 426
rect 684 311 792 317
rect 684 277 696 311
rect 780 277 792 311
rect 684 271 792 277
rect 574 -158 592 218
rect 626 -158 634 218
rect 840 218 900 366
rect 942 311 1050 317
rect 942 277 954 311
rect 1038 277 1050 311
rect 942 271 1050 277
rect 840 64 850 218
rect 574 -312 634 -158
rect 844 -158 850 64
rect 884 64 900 218
rect 1090 218 1150 702
rect 1354 702 1366 746
rect 1400 746 1406 1078
rect 1606 1078 1666 1564
rect 1862 1244 1868 1304
rect 1928 1244 1934 1304
rect 1716 1171 1824 1177
rect 1716 1137 1728 1171
rect 1812 1137 1824 1171
rect 1716 1131 1824 1137
rect 1400 702 1414 746
rect 1200 643 1308 649
rect 1200 609 1212 643
rect 1296 609 1308 643
rect 1200 603 1308 609
rect 1354 426 1414 702
rect 1606 702 1624 1078
rect 1658 702 1666 1078
rect 1868 1078 1928 1244
rect 1974 1171 2082 1177
rect 1974 1137 1986 1171
rect 2070 1137 2082 1171
rect 1974 1131 2082 1137
rect 1868 1046 1882 1078
rect 1458 643 1566 649
rect 1458 609 1470 643
rect 1554 609 1566 643
rect 1458 603 1566 609
rect 1220 366 1226 426
rect 1286 366 1292 426
rect 1348 366 1354 426
rect 1414 366 1420 426
rect 1474 366 1480 426
rect 1540 366 1546 426
rect 1226 317 1286 366
rect 1480 317 1540 366
rect 1200 311 1308 317
rect 1200 277 1212 311
rect 1296 277 1308 311
rect 1200 271 1308 277
rect 1458 311 1566 317
rect 1458 277 1470 311
rect 1554 277 1566 311
rect 1458 271 1566 277
rect 1090 150 1108 218
rect 884 -158 890 64
rect 844 -170 890 -158
rect 1102 -158 1108 150
rect 1142 150 1150 218
rect 1360 218 1406 230
rect 1142 -158 1148 150
rect 1360 -112 1366 218
rect 1102 -170 1148 -158
rect 1350 -158 1366 -112
rect 1400 -112 1406 218
rect 1606 218 1666 702
rect 1876 702 1882 1046
rect 1916 1046 1928 1078
rect 2124 1078 2184 1564
rect 2232 1171 2340 1177
rect 2232 1137 2244 1171
rect 2328 1137 2340 1171
rect 2232 1131 2340 1137
rect 1916 702 1922 1046
rect 1876 690 1922 702
rect 2124 702 2140 1078
rect 2174 702 2184 1078
rect 1716 643 1824 649
rect 1716 609 1728 643
rect 1812 609 1824 643
rect 1716 603 1824 609
rect 1974 643 2082 649
rect 1974 609 1986 643
rect 2070 609 2082 643
rect 1974 603 2082 609
rect 1738 426 1798 603
rect 1996 494 2056 603
rect 2124 498 2184 702
rect 2386 1078 2446 1564
rect 2502 1244 2508 1304
rect 2568 1244 2574 1304
rect 2386 702 2398 1078
rect 2432 702 2446 1078
rect 2232 643 2340 649
rect 2232 609 2244 643
rect 2328 609 2340 643
rect 2232 603 2340 609
rect 2260 498 2320 603
rect 2386 498 2446 702
rect 1990 434 1996 494
rect 2056 434 2062 494
rect 2124 438 2446 498
rect 1732 366 1738 426
rect 1798 366 1804 426
rect 1862 366 1868 426
rect 1928 366 1934 426
rect 1716 311 1824 317
rect 1716 277 1728 311
rect 1812 277 1824 311
rect 1716 271 1824 277
rect 1606 154 1624 218
rect 1400 -158 1410 -112
rect 684 -217 792 -211
rect 684 -251 696 -217
rect 780 -251 792 -217
rect 684 -257 792 -251
rect 942 -217 1050 -211
rect 942 -251 954 -217
rect 1038 -251 1050 -217
rect 942 -257 1050 -251
rect 1200 -217 1308 -211
rect 1200 -251 1212 -217
rect 1296 -251 1308 -217
rect 1200 -257 1308 -251
rect 712 -312 772 -257
rect 574 -372 772 -312
rect 960 -328 1020 -257
rect 1350 -328 1410 -158
rect 1618 -158 1624 154
rect 1658 154 1666 218
rect 1868 218 1928 366
rect 1996 317 2056 434
rect 1974 311 2082 317
rect 1974 277 1986 311
rect 2070 277 2082 311
rect 1974 271 2082 277
rect 1868 172 1882 218
rect 1658 -158 1664 154
rect 1618 -170 1664 -158
rect 1876 -158 1882 172
rect 1916 172 1928 218
rect 2124 218 2184 438
rect 2260 317 2320 438
rect 2232 311 2340 317
rect 2232 277 2244 311
rect 2328 277 2340 311
rect 2232 271 2340 277
rect 2124 172 2140 218
rect 1916 -158 1922 172
rect 1876 -170 1922 -158
rect 2134 -158 2140 172
rect 2174 172 2184 218
rect 2386 218 2446 438
rect 2386 176 2398 218
rect 2174 -158 2180 172
rect 2134 -170 2180 -158
rect 2392 -158 2398 176
rect 2432 176 2446 218
rect 2432 -158 2438 176
rect 2392 -170 2438 -158
rect 1458 -217 1566 -211
rect 1458 -251 1470 -217
rect 1554 -251 1566 -217
rect 1458 -257 1566 -251
rect 1716 -217 1824 -211
rect 1716 -251 1728 -217
rect 1812 -251 1824 -217
rect 1716 -257 1824 -251
rect 1974 -217 2082 -211
rect 1974 -251 1986 -217
rect 2070 -251 2082 -217
rect 1974 -257 2082 -251
rect 2232 -217 2340 -211
rect 2232 -251 2244 -217
rect 2328 -251 2340 -217
rect 2232 -257 2340 -251
rect 1738 -328 1798 -257
rect 2508 -328 2568 1244
rect 954 -388 960 -328
rect 1020 -388 1026 -328
rect 1344 -388 1350 -328
rect 1410 -388 1416 -328
rect 1732 -388 1738 -328
rect 1798 -388 1804 -328
rect 2502 -388 2508 -328
rect 2568 -388 2574 -328
rect 2678 -368 2684 1564
rect 2784 -368 2790 1798
rect 2678 -454 2790 -368
rect 374 -460 2790 -454
rect 374 -560 480 -460
rect 2684 -560 2790 -460
rect 374 -566 2790 -560
rect 626 -604 2470 -566
rect 626 -605 1480 -604
rect 626 -639 655 -605
rect 689 -639 747 -605
rect 781 -639 839 -605
rect 873 -639 931 -605
rect 965 -639 1023 -605
rect 1057 -639 1115 -605
rect 1149 -639 1207 -605
rect 1241 -639 1299 -605
rect 1333 -639 1391 -605
rect 1425 -638 1480 -605
rect 1514 -638 1572 -604
rect 1606 -605 2470 -604
rect 1606 -638 1669 -605
rect 1425 -639 1669 -638
rect 1703 -639 1761 -605
rect 1795 -639 1853 -605
rect 1887 -639 1945 -605
rect 1979 -639 2037 -605
rect 2071 -639 2129 -605
rect 2163 -639 2221 -605
rect 2255 -639 2313 -605
rect 2347 -639 2405 -605
rect 2439 -639 2470 -605
rect 626 -652 2470 -639
rect 626 -670 2468 -652
rect 2772 -680 2778 -620
rect 2838 -680 2844 -620
rect 798 -896 858 -890
rect 958 -896 1018 -890
rect 254 -902 752 -896
rect 254 -950 692 -902
rect 740 -950 752 -902
rect 254 -956 752 -950
rect 798 -902 1018 -896
rect 798 -950 804 -902
rect 852 -950 964 -902
rect 1012 -950 1018 -902
rect 798 -956 1018 -950
rect 1060 -902 1264 -896
rect 1060 -950 1072 -902
rect 1120 -950 1204 -902
rect 1252 -950 1264 -902
rect 1060 -956 1264 -950
rect 1366 -902 1612 -896
rect 1366 -950 1378 -902
rect 1426 -950 1612 -902
rect 1846 -898 1906 -892
rect 1960 -898 2020 -892
rect 2076 -896 2136 -890
rect 2236 -896 2296 -890
rect 1846 -904 2028 -898
rect 1366 -956 1612 -950
rect 254 -1988 314 -956
rect 798 -962 858 -956
rect 958 -962 1018 -956
rect 1378 -1014 1438 -1008
rect 1552 -1014 1612 -956
rect 1652 -964 1658 -904
rect 1718 -964 1724 -904
rect 1846 -952 1852 -904
rect 1900 -952 1966 -904
rect 2014 -952 2028 -904
rect 1846 -958 2028 -952
rect 2076 -902 2296 -896
rect 2076 -950 2082 -902
rect 2130 -950 2242 -902
rect 2290 -950 2296 -902
rect 2076 -956 2296 -950
rect 1846 -964 1906 -958
rect 1960 -964 2020 -958
rect 2076 -962 2136 -956
rect 2236 -962 2296 -956
rect 2348 -896 2408 -890
rect 2778 -896 2838 -680
rect 2348 -902 2838 -896
rect 2348 -950 2354 -902
rect 2402 -950 2838 -902
rect 2348 -956 2838 -950
rect 2348 -962 2408 -956
rect 1658 -1014 1718 -1008
rect 1372 -1074 1378 -1014
rect 1438 -1074 1444 -1014
rect 1552 -1020 1718 -1014
rect 1552 -1068 1664 -1020
rect 1712 -1068 1718 -1020
rect 1552 -1074 1718 -1068
rect 1378 -1080 1438 -1074
rect 1658 -1080 1718 -1074
rect 626 -1148 2468 -1118
rect 626 -1149 1572 -1148
rect 626 -1183 655 -1149
rect 689 -1183 747 -1149
rect 781 -1183 839 -1149
rect 873 -1183 931 -1149
rect 965 -1183 1023 -1149
rect 1057 -1183 1115 -1149
rect 1149 -1183 1207 -1149
rect 1241 -1183 1299 -1149
rect 1333 -1183 1391 -1149
rect 1425 -1150 1572 -1149
rect 1425 -1183 1480 -1150
rect 626 -1184 1480 -1183
rect 1514 -1182 1572 -1150
rect 1606 -1149 2468 -1148
rect 1606 -1182 1669 -1149
rect 1514 -1183 1669 -1182
rect 1703 -1183 1761 -1149
rect 1795 -1183 1853 -1149
rect 1887 -1183 1945 -1149
rect 1979 -1183 2037 -1149
rect 2071 -1183 2129 -1149
rect 2163 -1183 2221 -1149
rect 2255 -1183 2313 -1149
rect 2347 -1183 2405 -1149
rect 2439 -1183 2468 -1149
rect 1514 -1184 2468 -1183
rect 626 -1214 2468 -1184
rect 886 -1376 2256 -1214
rect 886 -1476 992 -1376
rect 2150 -1476 2256 -1376
rect 886 -1482 2256 -1476
rect 886 -1517 998 -1482
rect 412 -1654 472 -1640
rect 412 -1948 424 -1654
rect 458 -1948 472 -1654
rect 558 -1702 564 -1602
rect 664 -1702 670 -1602
rect 756 -1654 820 -1642
rect 532 -1744 578 -1732
rect 650 -1734 696 -1732
rect 532 -1764 538 -1744
rect 248 -2048 254 -1988
rect 314 -2048 320 -1988
rect 108 -2162 168 -2156
rect 412 -2282 472 -1948
rect 526 -1920 538 -1764
rect 572 -1764 578 -1744
rect 642 -1744 702 -1734
rect 572 -1920 586 -1764
rect 526 -1988 586 -1920
rect 642 -1920 656 -1744
rect 690 -1794 702 -1744
rect 690 -1920 704 -1794
rect 642 -1926 704 -1920
rect 642 -1988 702 -1926
rect 756 -1948 770 -1654
rect 804 -1948 820 -1654
rect 520 -2048 526 -1988
rect 586 -2048 592 -1988
rect 636 -2048 642 -1988
rect 702 -2048 708 -1988
rect 756 -2282 820 -1948
rect 886 -2282 892 -1517
rect 322 -2308 892 -2282
rect 992 -2280 998 -1517
rect 2144 -1516 2256 -1482
rect 1130 -1532 1190 -1526
rect 1242 -1532 1314 -1520
rect 1832 -1532 1904 -1520
rect 1190 -1592 1248 -1532
rect 1308 -1592 1838 -1532
rect 1898 -1592 1904 -1532
rect 1130 -1598 1190 -1592
rect 1242 -1604 1314 -1592
rect 1078 -1658 1124 -1646
rect 1078 -1814 1084 -1658
rect 1070 -1834 1084 -1814
rect 1118 -1814 1124 -1658
rect 1196 -1658 1242 -1646
rect 1196 -1814 1202 -1658
rect 1118 -1834 1130 -1814
rect 1070 -1884 1130 -1834
rect 1188 -1834 1202 -1814
rect 1236 -1814 1242 -1658
rect 1314 -1658 1360 -1646
rect 1314 -1808 1320 -1658
rect 1236 -1834 1248 -1814
rect 1064 -1896 1136 -1884
rect 1064 -1956 1070 -1896
rect 1130 -1956 1136 -1896
rect 1064 -1968 1136 -1956
rect 1070 -2280 1130 -1968
rect 1188 -2098 1248 -1834
rect 1310 -1834 1320 -1808
rect 1354 -1808 1360 -1658
rect 1424 -1658 1484 -1592
rect 1424 -1680 1438 -1658
rect 1354 -1834 1370 -1808
rect 1182 -2158 1188 -2098
rect 1248 -2158 1254 -2098
rect 1310 -2280 1370 -1834
rect 1432 -1834 1438 -1680
rect 1472 -1680 1484 -1658
rect 1550 -1658 1596 -1646
rect 1472 -1834 1478 -1680
rect 1550 -1822 1556 -1658
rect 1432 -1846 1478 -1834
rect 1542 -1834 1556 -1822
rect 1590 -1822 1596 -1658
rect 1662 -1658 1722 -1592
rect 1832 -1604 1904 -1592
rect 1662 -1672 1674 -1658
rect 1590 -1834 1602 -1822
rect 1440 -1898 1500 -1892
rect 1434 -1958 1440 -1898
rect 1500 -1958 1506 -1898
rect 1440 -1964 1500 -1958
rect 1542 -2280 1602 -1834
rect 1668 -1834 1674 -1672
rect 1708 -1672 1722 -1658
rect 1786 -1658 1832 -1646
rect 1708 -1834 1714 -1672
rect 1786 -1810 1792 -1658
rect 1668 -1846 1714 -1834
rect 1778 -1834 1792 -1810
rect 1826 -1810 1832 -1658
rect 1904 -1658 1950 -1646
rect 1904 -1810 1910 -1658
rect 1826 -1834 1838 -1810
rect 1660 -1898 1720 -1892
rect 1654 -1958 1660 -1898
rect 1720 -1958 1726 -1898
rect 1660 -1964 1720 -1958
rect 1778 -2280 1838 -1834
rect 1896 -1834 1910 -1810
rect 1944 -1810 1950 -1658
rect 2022 -1658 2068 -1646
rect 2022 -1792 2028 -1658
rect 1944 -1834 1956 -1810
rect 1896 -2098 1956 -1834
rect 2018 -1834 2028 -1792
rect 2062 -1792 2068 -1658
rect 2062 -1834 2078 -1792
rect 2018 -1884 2078 -1834
rect 2012 -1896 2084 -1884
rect 2012 -1956 2018 -1896
rect 2078 -1956 2084 -1896
rect 2012 -1968 2084 -1956
rect 1890 -2158 1896 -2098
rect 1956 -2158 1962 -2098
rect 2018 -2280 2078 -1968
rect 2144 -2280 2150 -1516
rect 992 -2308 2150 -2280
rect 2250 -2280 2256 -1516
rect 2316 -1654 2376 -1642
rect 2316 -1948 2328 -1654
rect 2362 -1948 2376 -1654
rect 2462 -1704 2468 -1604
rect 2568 -1704 2574 -1604
rect 2662 -1654 2722 -1644
rect 2436 -1744 2482 -1732
rect 2436 -1884 2442 -1744
rect 2316 -2280 2376 -1948
rect 2426 -1920 2442 -1884
rect 2476 -1884 2482 -1744
rect 2554 -1744 2600 -1732
rect 2554 -1878 2560 -1744
rect 2476 -1920 2486 -1884
rect 2426 -2098 2486 -1920
rect 2546 -1920 2560 -1878
rect 2594 -1878 2600 -1744
rect 2594 -1920 2606 -1878
rect 2546 -1998 2606 -1920
rect 2662 -1948 2674 -1654
rect 2708 -1948 2722 -1654
rect 2540 -2058 2546 -1998
rect 2606 -2058 2612 -1998
rect 2420 -2158 2426 -2098
rect 2486 -2158 2492 -2098
rect 2662 -2280 2722 -1948
rect 2778 -1998 2838 -956
rect 2772 -2058 2778 -1998
rect 2838 -2058 2844 -1998
rect 2250 -2308 2810 -2280
rect 322 -2614 346 -2308
rect 2790 -2614 2810 -2308
rect 322 -2632 2810 -2614
rect 886 -2634 2256 -2632
rect 886 -2734 992 -2634
rect 2150 -2734 2256 -2634
rect 886 -2740 2256 -2734
<< via1 >>
rect -3216 1584 -348 1884
rect -3098 536 -3038 596
rect -2214 654 -2154 714
rect -2344 536 -2284 596
rect -2086 536 -2026 596
rect -2600 -196 -2540 -136
rect -2730 -316 -2670 -256
rect -2346 -196 -2286 -136
rect -2086 -196 -2026 -136
rect -2216 -316 -2156 -256
rect -3098 -1052 -3038 -992
rect -1184 654 -1124 714
rect -1312 536 -1252 596
rect -1828 -196 -1768 -136
rect -1052 536 -992 596
rect -1570 -196 -1510 -136
rect -1700 -316 -1640 -256
rect -292 654 -232 714
rect -474 536 -414 596
rect -1312 -196 -1252 -136
rect -1054 -196 -994 -136
rect -1184 -316 -1124 -256
rect -2604 -1052 -2544 -992
rect -1828 -1052 -1768 -992
rect -2732 -1168 -2672 -1108
rect -796 -196 -736 -136
rect -672 -316 -612 -256
rect -1572 -1052 -1512 -992
rect -800 -1052 -740 -992
rect -1700 -1170 -1640 -1110
rect -670 -1170 -610 -1110
rect -292 -1170 -232 -1110
rect 254 366 314 426
rect 108 -316 168 -256
rect -1564 -1458 -1504 -1398
rect -1278 -1512 -1218 -1506
rect -1278 -1572 -1272 -1512
rect -1272 -1572 -1218 -1512
rect -1278 -1578 -1218 -1572
rect -183 -1507 -113 -1501
rect -183 -1577 -119 -1507
rect -119 -1577 -113 -1507
rect -183 -1583 -113 -1577
rect -1146 -1812 -1132 -1766
rect -1132 -1812 -1098 -1766
rect -1098 -1812 -1086 -1766
rect -1146 -1826 -1086 -1812
rect -890 -1812 -876 -1756
rect -876 -1812 -842 -1756
rect -842 -1812 -830 -1756
rect -890 -1816 -830 -1812
rect -632 -1806 -620 -1746
rect -620 -1806 -586 -1746
rect -586 -1806 -572 -1746
rect -380 -1808 -364 -1748
rect -364 -1808 -330 -1748
rect -330 -1808 -320 -1748
rect -246 -1806 -236 -1746
rect -236 -1806 -202 -1746
rect -202 -1806 -186 -1746
rect -1146 -2138 -1086 -2078
rect -890 -2136 -830 -2076
rect -632 -2136 -572 -2076
rect -380 -2136 -320 -2076
rect 1056 1584 2676 1884
rect 840 1244 900 1304
rect 1226 1244 1286 1304
rect 1484 1244 1544 1304
rect 840 366 900 426
rect 964 366 1024 426
rect 1868 1244 1928 1304
rect 1226 366 1286 426
rect 1354 366 1414 426
rect 1480 366 1540 426
rect 2508 1244 2568 1304
rect 1996 434 2056 494
rect 1738 366 1798 426
rect 1868 366 1928 426
rect 960 -388 1020 -328
rect 1350 -388 1410 -328
rect 1738 -388 1798 -328
rect 2508 -388 2568 -328
rect 2778 -680 2838 -620
rect 1658 -916 1718 -904
rect 1658 -950 1674 -916
rect 1674 -950 1708 -916
rect 1708 -950 1718 -916
rect 1658 -964 1718 -950
rect 1378 -1020 1438 -1014
rect 1378 -1068 1384 -1020
rect 1384 -1068 1432 -1020
rect 1432 -1068 1438 -1020
rect 1378 -1074 1438 -1068
rect 564 -1660 664 -1602
rect 564 -1694 597 -1660
rect 597 -1694 631 -1660
rect 631 -1694 664 -1660
rect 564 -1702 664 -1694
rect 254 -2048 314 -1988
rect 108 -2156 168 -2096
rect 526 -2048 586 -1988
rect 642 -2048 702 -1988
rect 1130 -1592 1190 -1532
rect 1188 -2158 1248 -2098
rect 1440 -1904 1500 -1898
rect 1440 -1952 1446 -1904
rect 1446 -1952 1494 -1904
rect 1494 -1952 1500 -1904
rect 1440 -1958 1500 -1952
rect 1660 -1904 1720 -1898
rect 1660 -1952 1666 -1904
rect 1666 -1952 1714 -1904
rect 1714 -1952 1720 -1904
rect 1660 -1958 1720 -1952
rect 1896 -2158 1956 -2098
rect 2468 -1660 2568 -1604
rect 2468 -1694 2501 -1660
rect 2501 -1694 2535 -1660
rect 2535 -1694 2568 -1660
rect 2468 -1704 2568 -1694
rect 2546 -2058 2606 -1998
rect 2426 -2158 2486 -2098
rect 2778 -2058 2838 -1998
rect 346 -2593 892 -2308
rect 892 -2593 992 -2308
rect 992 -2593 2150 -2308
rect 2150 -2593 2250 -2308
rect 2250 -2593 2790 -2308
rect 346 -2614 2790 -2593
<< metal2 >>
rect -3216 1884 -348 1894
rect 1056 1884 2676 1894
rect -348 1584 -112 1650
rect -3216 1574 -112 1584
rect 1056 1574 2676 1584
rect -2214 714 -2154 720
rect -1184 714 -1124 720
rect -292 714 -232 720
rect -2154 654 -1184 714
rect -1124 654 -292 714
rect -2214 648 -2154 654
rect -1184 648 -1124 654
rect -292 648 -232 654
rect -3098 596 -3038 602
rect -2344 596 -2284 602
rect -2086 596 -2026 602
rect -1312 596 -1252 602
rect -1052 596 -992 602
rect -3038 536 -2344 596
rect -2284 536 -2086 596
rect -2026 536 -1312 596
rect -1252 536 -1052 596
rect -3098 530 -3038 536
rect -2344 530 -2284 536
rect -2086 530 -2026 536
rect -1312 530 -1252 536
rect -1052 530 -992 536
rect -474 596 -414 602
rect -172 596 -112 1574
rect 840 1304 900 1310
rect 1226 1304 1286 1310
rect 1484 1304 1544 1310
rect 1868 1304 1928 1310
rect 2508 1304 2568 1310
rect 900 1244 1226 1304
rect 1286 1244 1484 1304
rect 1544 1244 1868 1304
rect 1928 1244 2508 1304
rect 840 1238 900 1244
rect 1226 1238 1286 1244
rect 1484 1238 1544 1244
rect 1868 1238 1928 1244
rect 2508 1238 2568 1244
rect -414 536 -112 596
rect -474 530 -414 536
rect 1996 494 2056 500
rect 1987 434 1996 494
rect 2056 434 2065 494
rect 254 426 314 432
rect 840 426 900 432
rect 964 426 1024 432
rect 1226 426 1286 432
rect 1354 426 1414 432
rect 1480 426 1540 432
rect 1738 426 1798 432
rect 1868 426 1928 432
rect 1996 428 2056 434
rect 314 366 840 426
rect 900 366 964 426
rect 1024 366 1226 426
rect 1286 366 1354 426
rect 1414 366 1480 426
rect 1540 366 1738 426
rect 1798 366 1868 426
rect 254 360 314 366
rect 840 360 900 366
rect 964 360 1024 366
rect 1226 360 1286 366
rect 1354 360 1414 366
rect 1480 360 1540 366
rect 1738 360 1798 366
rect 1868 360 1928 366
rect -2600 -136 -2540 -130
rect -2346 -136 -2286 -130
rect -2086 -136 -2026 -130
rect -1828 -136 -1768 -130
rect -1570 -136 -1510 -130
rect -1312 -136 -1252 -130
rect -1054 -136 -994 -130
rect -796 -136 -736 -130
rect -2540 -196 -2346 -136
rect -2286 -196 -2086 -136
rect -2026 -196 -1828 -136
rect -1768 -196 -1570 -136
rect -1510 -196 -1312 -136
rect -1252 -196 -1054 -136
rect -994 -196 -796 -136
rect -2600 -202 -2540 -196
rect -2346 -202 -2286 -196
rect -2086 -202 -2026 -196
rect -1828 -202 -1768 -196
rect -1570 -202 -1510 -196
rect -1312 -202 -1252 -196
rect -1054 -202 -994 -196
rect -796 -202 -736 -196
rect -2730 -256 -2670 -250
rect -2216 -256 -2156 -250
rect -1700 -256 -1640 -250
rect -1184 -256 -1124 -250
rect -672 -256 -612 -250
rect 108 -256 168 -250
rect -2670 -316 -2216 -256
rect -2156 -316 -1700 -256
rect -1640 -316 -1184 -256
rect -1124 -316 -672 -256
rect -612 -316 108 -256
rect -2730 -322 -2670 -316
rect -2216 -322 -2156 -316
rect -1700 -322 -1640 -316
rect -1184 -322 -1124 -316
rect -672 -322 -612 -316
rect 108 -322 168 -316
rect 960 -328 1020 -322
rect 1350 -328 1410 -322
rect 1738 -328 1798 -322
rect 2508 -328 2568 -322
rect 1020 -388 1350 -328
rect 1410 -388 1738 -328
rect 1798 -388 2508 -328
rect 2568 -388 2838 -328
rect 960 -394 1020 -388
rect 1350 -394 1410 -388
rect 1738 -394 1798 -388
rect 2508 -394 2568 -388
rect 1484 -570 2616 -510
rect 1484 -904 1544 -570
rect 1658 -904 1718 -898
rect 1484 -964 1658 -904
rect -3098 -992 -3038 -986
rect -2604 -992 -2544 -986
rect -1828 -992 -1768 -986
rect -1572 -992 -1512 -986
rect -800 -992 -740 -986
rect -3038 -1052 -2604 -992
rect -2544 -1052 -1828 -992
rect -1768 -1052 -1572 -992
rect -1512 -1052 -800 -992
rect -3098 -1058 -3038 -1052
rect -2604 -1058 -2544 -1052
rect -1828 -1058 -1768 -1052
rect -1572 -1058 -1512 -1052
rect -800 -1058 -740 -1052
rect 1378 -1014 1438 -1008
rect 1484 -1014 1544 -964
rect 1658 -970 1718 -964
rect 2556 -962 2616 -570
rect 2778 -620 2838 -388
rect 2778 -686 2838 -680
rect 1438 -1074 1544 -1014
rect 2556 -1022 2844 -962
rect 1378 -1080 1438 -1074
rect -2732 -1108 -2672 -1102
rect -2672 -1110 586 -1108
rect -2672 -1168 -1700 -1110
rect -2732 -1174 -2672 -1168
rect -1706 -1170 -1700 -1168
rect -1640 -1168 -670 -1110
rect -1640 -1170 -1634 -1168
rect -1564 -1398 -1504 -1168
rect -676 -1170 -670 -1168
rect -610 -1168 -292 -1110
rect -610 -1170 -604 -1168
rect -298 -1170 -292 -1168
rect -232 -1168 586 -1110
rect -232 -1170 -226 -1168
rect 526 -1208 586 -1168
rect 526 -1268 1018 -1208
rect -1564 -1464 -1504 -1458
rect -1278 -1506 -1218 -1500
rect -183 -1501 -113 -1495
rect -1287 -1578 -1278 -1506
rect -1218 -1578 -1209 -1506
rect -1278 -1584 -1218 -1578
rect -192 -1583 -183 -1501
rect -113 -1583 -104 -1501
rect 958 -1532 1018 -1268
rect -183 -1589 -113 -1583
rect 958 -1592 1130 -1532
rect 1190 -1592 1196 -1532
rect 564 -1602 664 -1596
rect 560 -1697 564 -1607
rect 664 -1697 668 -1607
rect 564 -1708 664 -1702
rect -632 -1746 -572 -1740
rect -890 -1756 -830 -1750
rect -1146 -1766 -1086 -1760
rect -1146 -2078 -1086 -1826
rect -1146 -2144 -1086 -2138
rect -890 -2076 -830 -1816
rect -890 -2142 -830 -2136
rect -632 -2076 -572 -1806
rect -380 -1748 -320 -1742
rect -380 -2076 -320 -1808
rect -246 -1746 -186 -1740
rect -386 -2136 -380 -2076
rect -320 -2136 -314 -2076
rect -246 -2098 -186 -1806
rect 254 -1988 314 -1982
rect 526 -1988 586 -1982
rect 642 -1988 702 -1982
rect 958 -1988 1018 -1592
rect 2468 -1604 2568 -1598
rect 2464 -1699 2468 -1609
rect 2568 -1699 2572 -1609
rect 2468 -1710 2568 -1704
rect 1434 -1958 1440 -1898
rect 1500 -1958 1660 -1898
rect 1720 -1958 1726 -1898
rect 314 -2048 526 -1988
rect 636 -2048 642 -1988
rect 702 -2048 1018 -1988
rect 254 -2054 314 -2048
rect 526 -2054 586 -2048
rect 642 -2054 702 -2048
rect 102 -2098 108 -2096
rect -632 -2142 -572 -2136
rect -246 -2156 108 -2098
rect 168 -2098 174 -2096
rect 1188 -2098 1248 -2092
rect 1542 -2098 1602 -1958
rect 2546 -1998 2606 -1992
rect 2778 -1998 2838 -1992
rect 2606 -2058 2778 -1998
rect 2546 -2064 2606 -2058
rect 2778 -2064 2838 -2058
rect 1896 -2098 1956 -2092
rect 2426 -2098 2486 -2092
rect 168 -2156 1188 -2098
rect -246 -2158 1188 -2156
rect 1248 -2158 1896 -2098
rect 1956 -2158 2426 -2098
rect 1188 -2164 1248 -2158
rect 2426 -2164 2486 -2158
rect 346 -2308 2790 -2298
rect 346 -2624 2790 -2614
<< via2 >>
rect -3216 1584 -348 1884
rect 1056 1584 2676 1884
rect 1996 434 2056 494
rect -1278 -1578 -1218 -1506
rect -183 -1583 -113 -1501
rect 569 -1697 659 -1607
rect 2473 -1699 2563 -1609
rect 346 -2614 2790 -2308
<< metal3 >>
rect -3226 1884 -338 1889
rect -3226 1584 -3216 1884
rect -348 1584 -338 1884
rect -3226 1579 -338 1584
rect 1046 1884 2686 1889
rect 1046 1584 1056 1884
rect 2676 1584 2686 1884
rect 1046 1579 2686 1584
rect 1978 499 2078 516
rect 1978 494 1997 499
rect 1978 434 1996 494
rect 1978 429 1997 434
rect 2061 429 2078 499
rect 1978 416 2078 429
rect 2946 -1238 3046 -1232
rect -2188 -1590 -2182 -1490
rect -2082 -1590 -2076 -1490
rect -1298 -1501 -1196 -1492
rect -1298 -1583 -1283 -1501
rect -1219 -1506 -1196 -1501
rect -1218 -1578 -1196 -1506
rect -1219 -1583 -1196 -1578
rect -2182 -2858 -2082 -1590
rect -1298 -1592 -1196 -1583
rect -202 -1496 -96 -1488
rect -202 -1501 -178 -1496
rect -202 -1583 -183 -1501
rect -202 -1588 -178 -1583
rect -108 -1588 -96 -1496
rect -202 -1596 -96 -1588
rect 564 -1603 664 -1602
rect 559 -1701 565 -1603
rect 663 -1701 669 -1603
rect 2468 -1605 2568 -1604
rect 564 -1702 664 -1701
rect 2463 -1703 2469 -1605
rect 2567 -1703 2573 -1605
rect 2468 -1704 2568 -1703
rect 336 -2308 2800 -2303
rect 336 -2614 346 -2308
rect 2790 -2614 2800 -2308
rect 336 -2619 2800 -2614
rect 2946 -2858 3046 -1338
rect -2182 -2958 3046 -2858
<< via3 >>
rect -3216 1584 -348 1884
rect 1056 1584 2676 1884
rect 1997 494 2061 499
rect 1997 434 2056 494
rect 2056 434 2061 494
rect 1997 429 2061 434
rect 2946 -1338 3046 -1238
rect -2182 -1590 -2082 -1490
rect -1283 -1506 -1219 -1501
rect -1283 -1578 -1278 -1506
rect -1278 -1578 -1219 -1506
rect -1283 -1583 -1219 -1578
rect -178 -1501 -108 -1496
rect -178 -1583 -113 -1501
rect -113 -1583 -108 -1501
rect -178 -1588 -108 -1583
rect 565 -1607 663 -1603
rect 565 -1697 569 -1607
rect 569 -1697 659 -1607
rect 659 -1697 663 -1607
rect 565 -1701 663 -1697
rect 2469 -1609 2567 -1605
rect 2469 -1699 2473 -1609
rect 2473 -1699 2563 -1609
rect 2563 -1699 2567 -1609
rect 2469 -1703 2567 -1699
rect 346 -2614 2790 -2308
<< metal4 >>
rect -3400 1884 2890 2278
rect -3400 1584 -3216 1884
rect -348 1584 1056 1884
rect 2676 1584 2890 1884
rect -3400 1478 2890 1584
rect 1976 499 3044 516
rect 1976 429 1997 499
rect 2061 429 3044 499
rect 1976 416 3044 429
rect 2944 -1237 3044 416
rect 2944 -1238 3047 -1237
rect 2944 -1244 2946 -1238
rect 2468 -1338 2946 -1244
rect 3046 -1338 3047 -1238
rect 2468 -1339 3047 -1338
rect 2468 -1344 3044 -1339
rect -2183 -1490 -2081 -1489
rect -2183 -1492 -2182 -1490
rect -2190 -1590 -2182 -1492
rect -2082 -1492 -2081 -1490
rect -2082 -1496 668 -1492
rect -2082 -1501 -178 -1496
rect -2082 -1583 -1283 -1501
rect -1219 -1583 -178 -1501
rect -2082 -1588 -178 -1583
rect -108 -1588 668 -1496
rect -2082 -1590 668 -1588
rect -2190 -1592 668 -1590
rect 564 -1603 668 -1592
rect 564 -1701 565 -1603
rect 663 -1701 668 -1603
rect 564 -1702 668 -1701
rect 568 -1706 668 -1702
rect 2468 -1605 2568 -1344
rect 2468 -1703 2469 -1605
rect 2567 -1703 2568 -1605
rect 2468 -1704 2568 -1703
rect -3400 -2308 2890 -2214
rect -3400 -2614 346 -2308
rect 2790 -2614 2890 -2308
rect -3400 -3014 2890 -2614
<< labels >>
flabel metal4 324 2134 340 2140 1 FreeSans 480 0 0 0 VDD
port 7 n power bidirectional
flabel metal1 -3086 -112 -3072 -100 1 FreeSans 480 0 0 0 vip
port 1 n
flabel metal1 -2316 -232 -2306 -222 1 FreeSans 480 0 0 0 vim
port 2 n
flabel metal1 -276 278 -262 298 1 FreeSans 480 0 0 0 vlatchm
flabel metal1 -2710 -188 -2696 -178 1 FreeSans 480 0 0 0 vlatchp
flabel metal1 -1664 800 -1646 814 1 FreeSans 480 0 0 0 vtailp
flabel metal1 -1746 918 -1726 930 1 FreeSans 480 0 0 0 ibiasp
port 6 n
flabel via1 862 368 878 384 1 FreeSans 480 0 0 0 vcompm
flabel metal1 2526 590 2546 614 1 FreeSans 480 0 0 0 vcompp
flabel metal4 -186 -2534 -160 -2514 1 FreeSans 480 0 0 0 VSS
port 8 n ground bidirectional
flabel metal1 1360 -1568 1366 -1562 1 FreeSans 480 0 0 0 vlatchm
flabel metal2 1448 -2134 1456 -2126 1 FreeSans 480 0 0 0 vlatchp
flabel metal1 1156 -934 1162 -928 1 FreeSans 160 0 0 0 vcompm_buf
flabel metal1 900 -934 906 -930 1 FreeSans 160 0 0 0 vcompmb
flabel metal1 1924 -930 1928 -926 1 FreeSans 160 0 0 0 vcompp_buf
flabel metal1 2178 -932 2184 -928 1 FreeSans 160 0 0 0 vcomppb
flabel metal2 2674 -990 2680 -984 1 FreeSans 480 0 0 0 vop
port 3 n
flabel metal1 1606 -1052 1612 -1044 1 FreeSans 480 0 0 0 vom
port 4 n
flabel metal4 -1548 -1552 -1528 -1534 1 FreeSans 480 0 0 0 clk
port 5 n
flabel locali 1762 -1081 1796 -1047 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_1/Y
flabel locali 1762 -1013 1796 -979 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_1/Y
flabel locali 1762 -945 1796 -911 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_1/Y
flabel locali 1854 -945 1888 -911 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_1/B
flabel locali 1670 -945 1704 -911 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_1/A
flabel nwell 1854 -639 1888 -605 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_1/VPB
flabel pwell 1854 -1183 1888 -1149 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_1/VNB
flabel metal1 1854 -1183 1888 -1149 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_1/VGND
flabel metal1 1854 -639 1888 -605 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_1/VPWR
rlabel comment 1916 -1166 1916 -1166 6 sky130_fd_sc_hd__nand2_1_1/nand2_1
flabel locali 1298 -1081 1332 -1047 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/Y
flabel locali 1298 -1013 1332 -979 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/Y
flabel locali 1298 -945 1332 -911 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/Y
flabel locali 1206 -945 1240 -911 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/B
flabel locali 1390 -945 1424 -911 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/A
flabel nwell 1206 -639 1240 -605 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VPB
flabel pwell 1206 -1183 1240 -1149 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VNB
flabel metal1 1206 -1183 1240 -1149 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VGND
flabel metal1 1206 -639 1240 -605 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VPWR
rlabel comment 1178 -1166 1178 -1166 4 sky130_fd_sc_hd__nand2_1_0/nand2_1
flabel locali 790 -877 824 -843 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 790 -945 824 -911 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 698 -945 732 -911 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/A
flabel nwell 655 -639 689 -605 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 655 -1183 689 -1149 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 655 -1183 689 -1149 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 655 -639 689 -605 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 626 -1166 626 -1166 4 sky130_fd_sc_hd__inv_1_0/inv_1
flabel locali 1066 -877 1100 -843 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/Y
flabel locali 1066 -945 1100 -911 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/Y
flabel locali 974 -945 1008 -911 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/A
flabel nwell 931 -639 965 -605 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VPB
flabel pwell 931 -1183 965 -1149 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VNB
flabel metal1 931 -1183 965 -1149 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VGND
flabel metal1 931 -639 965 -605 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VPWR
rlabel comment 902 -1166 902 -1166 4 sky130_fd_sc_hd__inv_1_1/inv_1
flabel locali 1994 -877 2028 -843 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_2/Y
flabel locali 1994 -945 2028 -911 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_2/Y
flabel locali 2086 -945 2120 -911 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_2/A
flabel nwell 2129 -639 2163 -605 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_2/VPB
flabel pwell 2129 -1183 2163 -1149 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_2/VNB
flabel metal1 2129 -1183 2163 -1149 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_2/VGND
flabel metal1 2129 -639 2163 -605 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_2/VPWR
rlabel comment 2192 -1166 2192 -1166 6 sky130_fd_sc_hd__inv_1_2/inv_1
flabel locali 2270 -877 2304 -843 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_3/Y
flabel locali 2270 -945 2304 -911 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_3/Y
flabel locali 2362 -945 2396 -911 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_3/A
flabel nwell 2405 -639 2439 -605 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_3/VPB
flabel pwell 2405 -1183 2439 -1149 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_3/VNB
flabel metal1 2405 -1183 2439 -1149 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_3/VGND
flabel metal1 2405 -639 2439 -605 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_3/VPWR
rlabel comment 2468 -1166 2468 -1166 6 sky130_fd_sc_hd__inv_1_3/inv_1
<< end >>
