magic
tech sky130A
magscale 1 2
timestamp 1626064199
<< obsli1 >>
rect 0 0 513728 512992
<< obsm1 >>
rect 0 0 513728 512992
<< obsm2 >>
rect 0 0 513728 512992
<< obsm3 >>
rect 0 0 513728 512992
<< metal4 >>
rect 808 0 2440 512992
rect 3256 0 4888 512992
rect 5440 816 6112 512176
rect 8160 3264 8832 509728
rect 16320 816 16992 512176
rect 19040 158432 19712 509728
rect 19968 407204 20328 493392
rect 27200 493032 27872 512176
rect 20688 407924 21048 492672
rect 29920 492312 30592 509728
rect 38080 493032 38752 512176
rect 40800 492312 41472 509728
rect 48960 493032 49632 512176
rect 51680 492312 52352 509728
rect 59840 493032 60512 512176
rect 62560 492312 63232 509728
rect 70720 493032 71392 512176
rect 73440 492312 74112 509728
rect 81600 493032 82272 512176
rect 84320 492312 84992 509728
rect 92480 493032 93152 512176
rect 95200 492312 95872 509728
rect 103360 493032 104032 512176
rect 106080 492312 106752 509728
rect 107604 492312 108276 509728
rect 109404 493032 110076 512176
rect 114240 493032 114912 512176
rect 116960 492312 117632 509728
rect 125120 493032 125792 512176
rect 127840 492312 128512 509728
rect 136000 493032 136672 512176
rect 138720 492312 139392 509728
rect 146880 493032 147552 512176
rect 149600 492312 150272 509728
rect 157760 493032 158432 512176
rect 21680 491332 22028 491680
rect 22360 490652 22708 491000
rect 19968 315544 20328 401732
rect 27200 401372 27872 407564
rect 20688 316264 21048 401012
rect 29920 400652 30592 408284
rect 38080 401372 38752 407564
rect 40800 400652 41472 408284
rect 48960 401372 49632 407564
rect 51680 400652 52352 408284
rect 59840 401372 60512 407564
rect 62560 400652 63232 408284
rect 70720 401372 71392 407564
rect 73440 400652 74112 408284
rect 81600 401372 82272 407564
rect 84320 400652 84992 408284
rect 92480 401372 93152 407564
rect 95200 400652 95872 408284
rect 103360 401372 104032 407564
rect 106080 400652 106752 408284
rect 107604 400652 108276 408284
rect 109404 401372 110076 407564
rect 114240 401372 114912 407564
rect 116960 400652 117632 408284
rect 125120 401372 125792 407564
rect 127840 400652 128512 408284
rect 136000 401372 136672 407564
rect 138720 400652 139392 408284
rect 146880 401372 147552 407564
rect 149600 400652 150272 408284
rect 158388 407924 158748 492672
rect 157760 401372 158432 407564
rect 159108 407204 159468 493392
rect 21680 399672 22028 400020
rect 22360 398992 22708 399340
rect 19968 164572 20328 304072
rect 27200 303712 27872 315904
rect 20688 165292 21048 303352
rect 29920 302992 30592 316624
rect 38080 303712 38752 315904
rect 40800 302992 41472 316624
rect 48960 303712 49632 315904
rect 51680 302992 52352 316624
rect 59840 303712 60512 315904
rect 62560 302992 63232 316624
rect 70720 303712 71392 315904
rect 73440 302992 74112 316624
rect 81600 303712 82272 315904
rect 84320 302992 84992 316624
rect 92480 303712 93152 315904
rect 95200 302992 95872 316624
rect 103360 303712 104032 315904
rect 106080 310075 106752 316624
rect 21680 302012 22028 302360
rect 22360 166964 22708 167312
rect 18816 153824 19712 158432
rect 19040 3264 19712 153824
rect 19968 19600 20328 159100
rect 27200 158740 27872 164932
rect 20688 20320 21048 158380
rect 29920 158020 30592 165652
rect 38080 158740 38752 164932
rect 40800 158020 41472 165652
rect 48960 158740 49632 164932
rect 51680 158020 52352 165652
rect 59840 158740 60512 164932
rect 62560 158020 63232 165652
rect 70720 158740 71392 164932
rect 73440 158020 74112 165652
rect 81600 158740 82272 164932
rect 84320 158020 84992 165652
rect 92480 158740 93152 164932
rect 95200 158020 95872 165652
rect 105076 165292 105436 303352
rect 103360 158740 104032 164932
rect 105796 164572 106156 304072
rect 21680 157040 22028 157388
rect 22360 21992 22708 22340
rect 27200 816 27872 19960
rect 29920 3264 30592 20680
rect 38080 816 38752 19960
rect 40800 3264 41472 20680
rect 48960 816 49632 19960
rect 51680 3264 52352 20680
rect 59840 816 60512 19960
rect 62560 3264 63232 20680
rect 70720 816 71392 19960
rect 73440 3264 74112 20680
rect 81600 816 82272 19960
rect 84320 3264 84992 20680
rect 92480 816 93152 19960
rect 95200 3264 95872 20680
rect 105076 20320 105436 158380
rect 103360 816 104032 19960
rect 105796 19600 106156 159100
rect 106636 153824 107308 158432
rect 106080 3264 106752 16993
rect 107604 3264 108276 316624
rect 109404 816 110076 315904
rect 111628 164572 111988 304072
rect 114240 303712 114912 315904
rect 112348 165292 112708 303352
rect 116960 302992 117632 316624
rect 125120 303712 125792 315904
rect 127840 302992 128512 316624
rect 136000 303712 136672 315904
rect 138720 302992 139392 316624
rect 146880 303712 147552 315904
rect 149600 302992 150272 316624
rect 158388 316264 158748 401012
rect 157760 303712 158432 315904
rect 159108 315544 159468 401732
rect 160480 302992 161152 509728
rect 162704 303712 163376 512176
rect 164940 407204 165300 493392
rect 168640 493032 169312 512176
rect 165660 407924 166020 492672
rect 171360 492312 172032 509728
rect 179520 493032 180192 512176
rect 182240 492312 182912 509728
rect 190400 493032 191072 512176
rect 193120 492312 193792 509728
rect 201280 493032 201952 512176
rect 204000 492312 204672 509728
rect 212160 493032 212832 512176
rect 214880 492312 215552 509728
rect 223040 493032 223712 512176
rect 225760 492312 226432 509728
rect 233920 493032 234592 512176
rect 236640 492312 237312 509728
rect 244800 493032 245472 512176
rect 247520 492312 248192 509728
rect 255680 493032 256352 512176
rect 258400 492312 259072 509728
rect 266560 493032 267232 512176
rect 269280 492312 269952 509728
rect 277440 493032 278112 512176
rect 280160 492312 280832 509728
rect 288320 493032 288992 512176
rect 291040 492312 291712 509728
rect 299200 493032 299872 512176
rect 301920 492312 302592 509728
rect 302380 491332 302728 491680
rect 167332 490652 167680 491000
rect 164940 315544 165300 401732
rect 168640 401372 169312 407564
rect 165660 316264 166020 401012
rect 171360 400652 172032 408284
rect 179520 401372 180192 407564
rect 182240 400652 182912 408284
rect 190400 401372 191072 407564
rect 193120 400652 193792 408284
rect 201280 401372 201952 407564
rect 204000 400652 204672 408284
rect 212160 401372 212832 407564
rect 214880 400652 215552 408284
rect 223040 401372 223712 407564
rect 225760 400652 226432 408284
rect 233920 401372 234592 407564
rect 236640 400652 237312 408284
rect 244800 401372 245472 407564
rect 247520 400652 248192 408284
rect 255680 401372 256352 407564
rect 258400 400652 259072 408284
rect 266560 401372 267232 407564
rect 269280 400652 269952 408284
rect 277440 401372 278112 407564
rect 280160 400652 280832 408284
rect 288320 401372 288992 407564
rect 291040 400652 291712 408284
rect 299200 401372 299872 407564
rect 301920 400652 302592 408284
rect 303360 407924 303720 492672
rect 304080 407204 304440 493392
rect 166652 399672 167000 400020
rect 301700 398992 302048 399340
rect 168640 303712 169312 315904
rect 171360 302992 172032 316624
rect 179520 303712 180192 315904
rect 182240 302992 182912 316624
rect 190400 303712 191072 315904
rect 193120 302992 193792 316624
rect 195756 302012 196104 302360
rect 195076 166964 195424 167312
rect 110476 153824 111148 158432
rect 111628 19600 111988 159100
rect 114240 158740 114912 164932
rect 112348 20320 112708 158380
rect 116960 158020 117632 165652
rect 125120 158740 125792 164932
rect 127840 158020 128512 165652
rect 136000 158740 136672 164932
rect 138720 158020 139392 165652
rect 146880 158740 147552 164932
rect 149600 158020 150272 165652
rect 157760 158740 158432 164932
rect 160480 158020 161152 165652
rect 162704 158740 163376 164932
rect 168640 158740 169312 164932
rect 171360 158020 172032 165652
rect 179520 158740 180192 164932
rect 182240 158020 182912 165652
rect 190400 158740 191072 164932
rect 193120 158020 193792 165652
rect 196736 165292 197096 303352
rect 197456 164572 197816 304072
rect 195756 157040 196104 157388
rect 195076 156360 195424 156708
rect 114240 816 114912 19960
rect 116960 3264 117632 20680
rect 125120 816 125792 19960
rect 127840 3264 128512 20680
rect 136000 816 136672 19960
rect 138720 3264 139392 20680
rect 146880 816 147552 19960
rect 149600 3264 150272 20680
rect 157760 816 158432 19960
rect 160480 3264 161152 20680
rect 162704 816 163376 19960
rect 168640 816 169312 19960
rect 171360 3264 172032 20680
rect 179520 816 180192 19960
rect 182240 3264 182912 20680
rect 190400 816 191072 19960
rect 193120 3264 193792 20680
rect 196736 20320 197096 158380
rect 197456 19600 197816 159100
rect 198296 153824 198968 158432
rect 201280 816 201952 315904
rect 204000 3264 204672 316624
rect 209288 111260 209648 197448
rect 212160 197088 212832 315904
rect 210008 111980 210368 196728
rect 214880 196368 215552 316624
rect 223040 197088 223712 315904
rect 225760 196368 226432 316624
rect 233920 197088 234592 315904
rect 236640 196368 237312 316624
rect 244800 197088 245472 315904
rect 247520 196368 248192 316624
rect 255680 197088 256352 315904
rect 258400 196368 259072 316624
rect 266560 197088 267232 315904
rect 269280 196368 269952 316624
rect 277440 197088 278112 315904
rect 280160 196368 280832 316624
rect 288320 197088 288992 315904
rect 291040 196368 291712 316624
rect 299200 197088 299872 315904
rect 301920 196368 302592 316624
rect 303360 316264 303720 401012
rect 304080 315544 304440 401732
rect 310080 197088 310752 512176
rect 312800 196368 313472 509728
rect 315912 353892 316272 493392
rect 320960 493032 321632 512176
rect 316632 354612 316992 492672
rect 323680 492312 324352 509728
rect 331840 493032 332512 512176
rect 334560 492312 335232 509728
rect 342720 493032 343392 512176
rect 345440 492312 346112 509728
rect 350304 492312 350976 509728
rect 352104 493032 352776 512176
rect 353600 493032 354272 512176
rect 356320 492312 356992 509728
rect 364480 493032 365152 512176
rect 367200 492312 367872 509728
rect 375360 493032 376032 512176
rect 378080 492312 378752 509728
rect 386240 493032 386912 512176
rect 388960 492312 389632 509728
rect 397120 493032 397792 512176
rect 399840 492312 400512 509728
rect 400040 491332 400388 491680
rect 318304 356284 318652 356632
rect 315912 208920 316272 348420
rect 320960 348060 321632 354252
rect 316632 209640 316992 347700
rect 323680 347340 324352 354972
rect 331840 348060 332512 354252
rect 334560 347340 335232 354972
rect 342720 348060 343392 354252
rect 345440 347340 346112 354972
rect 350304 347340 350976 354972
rect 352104 348060 352776 354252
rect 353600 348060 354272 354252
rect 356320 347340 356992 354972
rect 364480 348060 365152 354252
rect 367200 347340 367872 354972
rect 375360 348060 376032 354252
rect 378080 347340 378752 354972
rect 386240 348060 386912 354252
rect 388960 347340 389632 354972
rect 397120 348060 397792 354252
rect 399840 347340 400512 354972
rect 401020 354612 401380 492672
rect 401740 353892 402100 493392
rect 318304 211312 318652 211660
rect 400040 210632 400388 210980
rect 320960 197088 321632 209280
rect 323680 196368 324352 210000
rect 331840 197088 332512 209280
rect 334560 196368 335232 210000
rect 342720 197088 343392 209280
rect 345440 196368 346112 210000
rect 346048 194708 346396 195056
rect 346728 112972 347076 113320
rect 209288 19600 209648 105788
rect 212160 105428 212832 111620
rect 210008 20320 210368 105068
rect 214880 104708 215552 112340
rect 223040 105428 223712 111620
rect 225760 104708 226432 112340
rect 233920 105428 234592 111620
rect 236640 104708 237312 112340
rect 244800 105428 245472 111620
rect 247520 104708 248192 112340
rect 255680 105428 256352 111620
rect 258400 104708 259072 112340
rect 266560 105428 267232 111620
rect 269280 104708 269952 112340
rect 277440 105428 278112 111620
rect 280160 104708 280832 112340
rect 288320 105428 288992 111620
rect 291040 104708 291712 112340
rect 299200 105428 299872 111620
rect 301920 104708 302592 112340
rect 310080 105428 310752 111620
rect 312800 104708 313472 112340
rect 320960 105428 321632 111620
rect 323680 104708 324352 112340
rect 331840 105428 332512 111620
rect 334560 104708 335232 112340
rect 342720 105428 343392 111620
rect 345440 104708 346112 112340
rect 347708 111980 348068 196728
rect 348428 111260 348788 197448
rect 346048 103048 346396 103396
rect 346728 21312 347076 21660
rect 212160 816 212832 19960
rect 214880 3264 215552 20680
rect 223040 816 223712 19960
rect 225760 3264 226432 20680
rect 233920 816 234592 19960
rect 236640 3264 237312 20680
rect 244800 816 245472 19960
rect 247520 3264 248192 20680
rect 255680 816 256352 19960
rect 258400 3264 259072 20680
rect 266560 816 267232 19960
rect 269280 3264 269952 20680
rect 277440 816 278112 19960
rect 280160 3264 280832 20680
rect 288320 816 288992 19960
rect 291040 3264 291712 20680
rect 299200 816 299872 19960
rect 301920 3264 302592 20680
rect 310080 816 310752 19960
rect 312800 3264 313472 20680
rect 320960 816 321632 19960
rect 323680 3264 324352 20680
rect 331840 816 332512 19960
rect 334560 3264 335232 20680
rect 342720 816 343392 19960
rect 345440 3264 346112 20680
rect 347708 20320 348068 105068
rect 348428 19600 348788 105788
rect 350304 3264 350976 210000
rect 352104 816 352776 209280
rect 353600 197448 354272 209280
rect 353600 197088 354620 197448
rect 354260 111620 354620 197088
rect 354980 111980 355340 196728
rect 356320 196368 356992 210000
rect 364480 197088 365152 209280
rect 367200 196368 367872 210000
rect 375360 197088 376032 209280
rect 378080 196368 378752 210000
rect 386240 197088 386912 209280
rect 388960 196368 389632 210000
rect 397120 197088 397792 209280
rect 399840 196368 400512 210000
rect 401020 209640 401380 347700
rect 401740 208920 402100 348420
rect 403704 196368 404376 509728
rect 405504 197088 406176 512176
rect 408000 493872 408672 512176
rect 407572 353892 407932 493392
rect 408292 354612 408652 492672
rect 410720 492312 411392 509728
rect 418880 493032 419552 512176
rect 421600 492312 422272 509728
rect 429760 493032 430432 512176
rect 432480 492312 433152 509728
rect 440640 493032 441312 512176
rect 443360 492312 444032 509728
rect 451520 493032 452192 512176
rect 454240 492312 454912 509728
rect 462400 493032 463072 512176
rect 465120 492312 465792 509728
rect 473280 493032 473952 512176
rect 476000 492312 476672 509728
rect 484160 493032 484832 512176
rect 486880 492312 487552 509728
rect 491020 490652 491368 491000
rect 491700 355604 492048 355952
rect 408000 350880 408672 351554
rect 407572 208920 407932 348420
rect 408292 209640 408652 347700
rect 410720 347340 411392 354972
rect 418880 348060 419552 354252
rect 421600 347340 422272 354972
rect 429760 348060 430432 354252
rect 432480 347340 433152 354972
rect 440640 348060 441312 354252
rect 443360 347340 444032 354972
rect 451520 348060 452192 354252
rect 454240 347340 454912 354972
rect 462400 348060 463072 354252
rect 465120 347340 465792 354972
rect 473280 348060 473952 354252
rect 476000 347340 476672 354972
rect 484160 348060 484832 354252
rect 486880 347340 487552 354972
rect 492680 354612 493040 492672
rect 493400 353892 493760 493392
rect 491020 211312 491368 211660
rect 491700 210632 492048 210980
rect 408000 197088 408672 208440
rect 410720 196368 411392 210000
rect 418880 197088 419552 209280
rect 421600 196368 422272 210000
rect 429760 197088 430432 209280
rect 432480 196368 433152 210000
rect 440640 197088 441312 209280
rect 443360 196368 444032 210000
rect 451520 197088 452192 209280
rect 454240 196368 454912 210000
rect 462400 197088 463072 209280
rect 465120 196368 465792 210000
rect 473280 197088 473952 209280
rect 476000 196368 476672 210000
rect 484160 197088 484832 209280
rect 486880 196368 487552 210000
rect 492680 209640 493040 347700
rect 493400 208920 493760 348420
rect 491700 195388 492048 195736
rect 356652 194708 357000 195056
rect 353600 111260 354620 111620
rect 353600 105788 354272 111260
rect 353600 105428 354620 105788
rect 354260 19960 354620 105428
rect 354980 20320 355340 105068
rect 356320 104708 356992 112340
rect 364480 105428 365152 111620
rect 367200 104708 367872 112340
rect 375360 105428 376032 111620
rect 378080 104708 378752 112340
rect 386240 105428 386912 111620
rect 388960 104708 389632 112340
rect 397120 105428 397792 111620
rect 399840 104708 400512 112340
rect 403704 104708 404376 112340
rect 405504 105428 406176 111620
rect 408000 105428 408672 111620
rect 410720 104708 411392 112340
rect 418880 105428 419552 111620
rect 421600 104708 422272 112340
rect 429760 105428 430432 111620
rect 432480 104708 433152 112340
rect 440640 105428 441312 111620
rect 443360 104708 444032 112340
rect 451520 105428 452192 111620
rect 454240 104708 454912 112340
rect 462400 105428 463072 111620
rect 465120 104708 465792 112340
rect 473280 105428 473952 111620
rect 476000 104708 476672 112340
rect 484160 105428 484832 111620
rect 486880 104708 487552 112340
rect 492680 111980 493040 196728
rect 493400 111260 493760 197448
rect 356652 103048 357000 103396
rect 491700 21312 492048 21660
rect 353600 19600 354620 19960
rect 353600 816 354272 19600
rect 356320 3264 356992 20680
rect 364480 816 365152 19960
rect 367200 3264 367872 20680
rect 375360 816 376032 19960
rect 378080 3264 378752 20680
rect 386240 816 386912 19960
rect 388960 3264 389632 20680
rect 397120 816 397792 19960
rect 399840 3264 400512 20680
rect 403704 3264 404376 20680
rect 405504 816 406176 19960
rect 408000 816 408672 19960
rect 410720 3264 411392 20680
rect 418880 816 419552 19960
rect 421600 3264 422272 20680
rect 429760 816 430432 19960
rect 432480 3264 433152 20680
rect 440640 816 441312 19960
rect 443360 3264 444032 20680
rect 451520 816 452192 19960
rect 454240 3264 454912 20680
rect 462400 816 463072 19960
rect 465120 3264 465792 20680
rect 473280 816 473952 19960
rect 476000 3264 476672 20680
rect 484160 816 484832 19960
rect 486880 3264 487552 20680
rect 492680 20320 493040 105068
rect 493400 19600 493760 105788
rect 495040 816 495712 512176
rect 497760 3264 498432 509728
rect 505920 816 506592 512176
rect 508840 0 510472 512992
rect 511288 0 512920 512992
<< obsm4 >>
rect 0 0 808 512992
rect 2440 0 3256 512992
rect 4888 512176 508840 512992
rect 4888 816 5440 512176
rect 6112 509728 16320 512176
rect 6112 3264 8160 509728
rect 8832 3264 16320 509728
rect 6112 816 16320 3264
rect 16992 509728 27200 512176
rect 16992 158432 19040 509728
rect 19712 493392 27200 509728
rect 19712 407204 19968 493392
rect 20328 493032 27200 493392
rect 27872 509728 38080 512176
rect 27872 493032 29920 509728
rect 20328 492672 29920 493032
rect 20328 407924 20688 492672
rect 21048 492312 29920 492672
rect 30592 493032 38080 509728
rect 38752 509728 48960 512176
rect 38752 493032 40800 509728
rect 30592 492312 40800 493032
rect 41472 493032 48960 509728
rect 49632 509728 59840 512176
rect 49632 493032 51680 509728
rect 41472 492312 51680 493032
rect 52352 493032 59840 509728
rect 60512 509728 70720 512176
rect 60512 493032 62560 509728
rect 52352 492312 62560 493032
rect 63232 493032 70720 509728
rect 71392 509728 81600 512176
rect 71392 493032 73440 509728
rect 63232 492312 73440 493032
rect 74112 493032 81600 509728
rect 82272 509728 92480 512176
rect 82272 493032 84320 509728
rect 74112 492312 84320 493032
rect 84992 493032 92480 509728
rect 93152 509728 103360 512176
rect 93152 493032 95200 509728
rect 84992 492312 95200 493032
rect 95872 493032 103360 509728
rect 104032 509728 109404 512176
rect 104032 493032 106080 509728
rect 95872 492312 106080 493032
rect 106752 492312 107604 509728
rect 108276 493032 109404 509728
rect 110076 493032 114240 512176
rect 114912 509728 125120 512176
rect 114912 493032 116960 509728
rect 108276 492312 116960 493032
rect 117632 493032 125120 509728
rect 125792 509728 136000 512176
rect 125792 493032 127840 509728
rect 117632 492312 127840 493032
rect 128512 493032 136000 509728
rect 136672 509728 146880 512176
rect 136672 493032 138720 509728
rect 128512 492312 138720 493032
rect 139392 493032 146880 509728
rect 147552 509728 157760 512176
rect 147552 493032 149600 509728
rect 139392 492312 149600 493032
rect 150272 493032 157760 509728
rect 158432 509728 162704 512176
rect 158432 493392 160480 509728
rect 158432 493032 159108 493392
rect 150272 492672 159108 493032
rect 150272 492312 158388 492672
rect 21048 491680 158388 492312
rect 21048 491332 21680 491680
rect 22028 491332 158388 491680
rect 21048 491000 158388 491332
rect 21048 490652 22360 491000
rect 22708 490652 158388 491000
rect 21048 408284 158388 490652
rect 21048 407924 29920 408284
rect 20328 407564 29920 407924
rect 20328 407204 27200 407564
rect 19712 401732 27200 407204
rect 19712 315544 19968 401732
rect 20328 401372 27200 401732
rect 27872 401372 29920 407564
rect 20328 401012 29920 401372
rect 20328 316264 20688 401012
rect 21048 400652 29920 401012
rect 30592 407564 40800 408284
rect 30592 401372 38080 407564
rect 38752 401372 40800 407564
rect 30592 400652 40800 401372
rect 41472 407564 51680 408284
rect 41472 401372 48960 407564
rect 49632 401372 51680 407564
rect 41472 400652 51680 401372
rect 52352 407564 62560 408284
rect 52352 401372 59840 407564
rect 60512 401372 62560 407564
rect 52352 400652 62560 401372
rect 63232 407564 73440 408284
rect 63232 401372 70720 407564
rect 71392 401372 73440 407564
rect 63232 400652 73440 401372
rect 74112 407564 84320 408284
rect 74112 401372 81600 407564
rect 82272 401372 84320 407564
rect 74112 400652 84320 401372
rect 84992 407564 95200 408284
rect 84992 401372 92480 407564
rect 93152 401372 95200 407564
rect 84992 400652 95200 401372
rect 95872 407564 106080 408284
rect 95872 401372 103360 407564
rect 104032 401372 106080 407564
rect 95872 400652 106080 401372
rect 106752 400652 107604 408284
rect 108276 407564 116960 408284
rect 108276 401372 109404 407564
rect 110076 401372 114240 407564
rect 114912 401372 116960 407564
rect 108276 400652 116960 401372
rect 117632 407564 127840 408284
rect 117632 401372 125120 407564
rect 125792 401372 127840 407564
rect 117632 400652 127840 401372
rect 128512 407564 138720 408284
rect 128512 401372 136000 407564
rect 136672 401372 138720 407564
rect 128512 400652 138720 401372
rect 139392 407564 149600 408284
rect 139392 401372 146880 407564
rect 147552 401372 149600 407564
rect 139392 400652 149600 401372
rect 150272 407924 158388 408284
rect 158748 407924 159108 492672
rect 150272 407564 159108 407924
rect 150272 401372 157760 407564
rect 158432 407204 159108 407564
rect 159468 407204 160480 493392
rect 158432 401732 160480 407204
rect 158432 401372 159108 401732
rect 150272 401012 159108 401372
rect 150272 400652 158388 401012
rect 21048 400020 158388 400652
rect 21048 399672 21680 400020
rect 22028 399672 158388 400020
rect 21048 399340 158388 399672
rect 21048 398992 22360 399340
rect 22708 398992 158388 399340
rect 21048 316624 158388 398992
rect 21048 316264 29920 316624
rect 20328 315904 29920 316264
rect 20328 315544 27200 315904
rect 19712 304072 27200 315544
rect 19712 164572 19968 304072
rect 20328 303712 27200 304072
rect 27872 303712 29920 315904
rect 20328 303352 29920 303712
rect 20328 165292 20688 303352
rect 21048 302992 29920 303352
rect 30592 315904 40800 316624
rect 30592 303712 38080 315904
rect 38752 303712 40800 315904
rect 30592 302992 40800 303712
rect 41472 315904 51680 316624
rect 41472 303712 48960 315904
rect 49632 303712 51680 315904
rect 41472 302992 51680 303712
rect 52352 315904 62560 316624
rect 52352 303712 59840 315904
rect 60512 303712 62560 315904
rect 52352 302992 62560 303712
rect 63232 315904 73440 316624
rect 63232 303712 70720 315904
rect 71392 303712 73440 315904
rect 63232 302992 73440 303712
rect 74112 315904 84320 316624
rect 74112 303712 81600 315904
rect 82272 303712 84320 315904
rect 74112 302992 84320 303712
rect 84992 315904 95200 316624
rect 84992 303712 92480 315904
rect 93152 303712 95200 315904
rect 84992 302992 95200 303712
rect 95872 315904 106080 316624
rect 95872 303712 103360 315904
rect 104032 310075 106080 315904
rect 106752 310075 107604 316624
rect 104032 304072 107604 310075
rect 104032 303712 105796 304072
rect 95872 303352 105796 303712
rect 95872 302992 105076 303352
rect 21048 302360 105076 302992
rect 21048 302012 21680 302360
rect 22028 302012 105076 302360
rect 21048 167312 105076 302012
rect 21048 166964 22360 167312
rect 22708 166964 105076 167312
rect 21048 165652 105076 166964
rect 21048 165292 29920 165652
rect 20328 164932 29920 165292
rect 20328 164572 27200 164932
rect 19712 159100 27200 164572
rect 16992 153824 18816 158432
rect 16992 3264 19040 153824
rect 19712 19600 19968 159100
rect 20328 158740 27200 159100
rect 27872 158740 29920 164932
rect 20328 158380 29920 158740
rect 20328 20320 20688 158380
rect 21048 158020 29920 158380
rect 30592 164932 40800 165652
rect 30592 158740 38080 164932
rect 38752 158740 40800 164932
rect 30592 158020 40800 158740
rect 41472 164932 51680 165652
rect 41472 158740 48960 164932
rect 49632 158740 51680 164932
rect 41472 158020 51680 158740
rect 52352 164932 62560 165652
rect 52352 158740 59840 164932
rect 60512 158740 62560 164932
rect 52352 158020 62560 158740
rect 63232 164932 73440 165652
rect 63232 158740 70720 164932
rect 71392 158740 73440 164932
rect 63232 158020 73440 158740
rect 74112 164932 84320 165652
rect 74112 158740 81600 164932
rect 82272 158740 84320 164932
rect 74112 158020 84320 158740
rect 84992 164932 95200 165652
rect 84992 158740 92480 164932
rect 93152 158740 95200 164932
rect 84992 158020 95200 158740
rect 95872 165292 105076 165652
rect 105436 165292 105796 303352
rect 95872 164932 105796 165292
rect 95872 158740 103360 164932
rect 104032 164572 105796 164932
rect 106156 164572 107604 304072
rect 104032 159100 107604 164572
rect 104032 158740 105796 159100
rect 95872 158380 105796 158740
rect 95872 158020 105076 158380
rect 21048 157388 105076 158020
rect 21048 157040 21680 157388
rect 22028 157040 105076 157388
rect 21048 22340 105076 157040
rect 21048 21992 22360 22340
rect 22708 21992 105076 22340
rect 21048 20680 105076 21992
rect 21048 20320 29920 20680
rect 20328 19960 29920 20320
rect 20328 19600 27200 19960
rect 19712 3264 27200 19600
rect 16992 816 27200 3264
rect 27872 3264 29920 19960
rect 30592 19960 40800 20680
rect 30592 3264 38080 19960
rect 27872 816 38080 3264
rect 38752 3264 40800 19960
rect 41472 19960 51680 20680
rect 41472 3264 48960 19960
rect 38752 816 48960 3264
rect 49632 3264 51680 19960
rect 52352 19960 62560 20680
rect 52352 3264 59840 19960
rect 49632 816 59840 3264
rect 60512 3264 62560 19960
rect 63232 19960 73440 20680
rect 63232 3264 70720 19960
rect 60512 816 70720 3264
rect 71392 3264 73440 19960
rect 74112 19960 84320 20680
rect 74112 3264 81600 19960
rect 71392 816 81600 3264
rect 82272 3264 84320 19960
rect 84992 19960 95200 20680
rect 84992 3264 92480 19960
rect 82272 816 92480 3264
rect 93152 3264 95200 19960
rect 95872 20320 105076 20680
rect 105436 20320 105796 158380
rect 95872 19960 105796 20320
rect 95872 3264 103360 19960
rect 93152 816 103360 3264
rect 104032 19600 105796 19960
rect 106156 158432 107604 159100
rect 106156 153824 106636 158432
rect 107308 153824 107604 158432
rect 106156 19600 107604 153824
rect 104032 16993 107604 19600
rect 104032 3264 106080 16993
rect 106752 3264 107604 16993
rect 108276 315904 116960 316624
rect 108276 3264 109404 315904
rect 104032 816 109404 3264
rect 110076 304072 114240 315904
rect 110076 164572 111628 304072
rect 111988 303712 114240 304072
rect 114912 303712 116960 315904
rect 111988 303352 116960 303712
rect 111988 165292 112348 303352
rect 112708 302992 116960 303352
rect 117632 315904 127840 316624
rect 117632 303712 125120 315904
rect 125792 303712 127840 315904
rect 117632 302992 127840 303712
rect 128512 315904 138720 316624
rect 128512 303712 136000 315904
rect 136672 303712 138720 315904
rect 128512 302992 138720 303712
rect 139392 315904 149600 316624
rect 139392 303712 146880 315904
rect 147552 303712 149600 315904
rect 139392 302992 149600 303712
rect 150272 316264 158388 316624
rect 158748 316264 159108 401012
rect 150272 315904 159108 316264
rect 150272 303712 157760 315904
rect 158432 315544 159108 315904
rect 159468 315544 160480 401732
rect 158432 303712 160480 315544
rect 150272 302992 160480 303712
rect 161152 303712 162704 509728
rect 163376 493392 168640 512176
rect 163376 407204 164940 493392
rect 165300 493032 168640 493392
rect 169312 509728 179520 512176
rect 169312 493032 171360 509728
rect 165300 492672 171360 493032
rect 165300 407924 165660 492672
rect 166020 492312 171360 492672
rect 172032 493032 179520 509728
rect 180192 509728 190400 512176
rect 180192 493032 182240 509728
rect 172032 492312 182240 493032
rect 182912 493032 190400 509728
rect 191072 509728 201280 512176
rect 191072 493032 193120 509728
rect 182912 492312 193120 493032
rect 193792 493032 201280 509728
rect 201952 509728 212160 512176
rect 201952 493032 204000 509728
rect 193792 492312 204000 493032
rect 204672 493032 212160 509728
rect 212832 509728 223040 512176
rect 212832 493032 214880 509728
rect 204672 492312 214880 493032
rect 215552 493032 223040 509728
rect 223712 509728 233920 512176
rect 223712 493032 225760 509728
rect 215552 492312 225760 493032
rect 226432 493032 233920 509728
rect 234592 509728 244800 512176
rect 234592 493032 236640 509728
rect 226432 492312 236640 493032
rect 237312 493032 244800 509728
rect 245472 509728 255680 512176
rect 245472 493032 247520 509728
rect 237312 492312 247520 493032
rect 248192 493032 255680 509728
rect 256352 509728 266560 512176
rect 256352 493032 258400 509728
rect 248192 492312 258400 493032
rect 259072 493032 266560 509728
rect 267232 509728 277440 512176
rect 267232 493032 269280 509728
rect 259072 492312 269280 493032
rect 269952 493032 277440 509728
rect 278112 509728 288320 512176
rect 278112 493032 280160 509728
rect 269952 492312 280160 493032
rect 280832 493032 288320 509728
rect 288992 509728 299200 512176
rect 288992 493032 291040 509728
rect 280832 492312 291040 493032
rect 291712 493032 299200 509728
rect 299872 509728 310080 512176
rect 299872 493032 301920 509728
rect 291712 492312 301920 493032
rect 302592 493392 310080 509728
rect 302592 492672 304080 493392
rect 302592 492312 303360 492672
rect 166020 491680 303360 492312
rect 166020 491332 302380 491680
rect 302728 491332 303360 491680
rect 166020 491000 303360 491332
rect 166020 490652 167332 491000
rect 167680 490652 303360 491000
rect 166020 408284 303360 490652
rect 166020 407924 171360 408284
rect 165300 407564 171360 407924
rect 165300 407204 168640 407564
rect 163376 401732 168640 407204
rect 163376 315544 164940 401732
rect 165300 401372 168640 401732
rect 169312 401372 171360 407564
rect 165300 401012 171360 401372
rect 165300 316264 165660 401012
rect 166020 400652 171360 401012
rect 172032 407564 182240 408284
rect 172032 401372 179520 407564
rect 180192 401372 182240 407564
rect 172032 400652 182240 401372
rect 182912 407564 193120 408284
rect 182912 401372 190400 407564
rect 191072 401372 193120 407564
rect 182912 400652 193120 401372
rect 193792 407564 204000 408284
rect 193792 401372 201280 407564
rect 201952 401372 204000 407564
rect 193792 400652 204000 401372
rect 204672 407564 214880 408284
rect 204672 401372 212160 407564
rect 212832 401372 214880 407564
rect 204672 400652 214880 401372
rect 215552 407564 225760 408284
rect 215552 401372 223040 407564
rect 223712 401372 225760 407564
rect 215552 400652 225760 401372
rect 226432 407564 236640 408284
rect 226432 401372 233920 407564
rect 234592 401372 236640 407564
rect 226432 400652 236640 401372
rect 237312 407564 247520 408284
rect 237312 401372 244800 407564
rect 245472 401372 247520 407564
rect 237312 400652 247520 401372
rect 248192 407564 258400 408284
rect 248192 401372 255680 407564
rect 256352 401372 258400 407564
rect 248192 400652 258400 401372
rect 259072 407564 269280 408284
rect 259072 401372 266560 407564
rect 267232 401372 269280 407564
rect 259072 400652 269280 401372
rect 269952 407564 280160 408284
rect 269952 401372 277440 407564
rect 278112 401372 280160 407564
rect 269952 400652 280160 401372
rect 280832 407564 291040 408284
rect 280832 401372 288320 407564
rect 288992 401372 291040 407564
rect 280832 400652 291040 401372
rect 291712 407564 301920 408284
rect 291712 401372 299200 407564
rect 299872 401372 301920 407564
rect 291712 400652 301920 401372
rect 302592 407924 303360 408284
rect 303720 407924 304080 492672
rect 302592 407204 304080 407924
rect 304440 407204 310080 493392
rect 302592 401732 310080 407204
rect 302592 401012 304080 401732
rect 302592 400652 303360 401012
rect 166020 400020 303360 400652
rect 166020 399672 166652 400020
rect 167000 399672 303360 400020
rect 166020 399340 303360 399672
rect 166020 398992 301700 399340
rect 302048 398992 303360 399340
rect 166020 316624 303360 398992
rect 166020 316264 171360 316624
rect 165300 315904 171360 316264
rect 165300 315544 168640 315904
rect 163376 303712 168640 315544
rect 169312 303712 171360 315904
rect 161152 302992 171360 303712
rect 172032 315904 182240 316624
rect 172032 303712 179520 315904
rect 180192 303712 182240 315904
rect 172032 302992 182240 303712
rect 182912 315904 193120 316624
rect 182912 303712 190400 315904
rect 191072 303712 193120 315904
rect 182912 302992 193120 303712
rect 193792 315904 204000 316624
rect 193792 304072 201280 315904
rect 193792 303352 197456 304072
rect 193792 302992 196736 303352
rect 112708 302360 196736 302992
rect 112708 302012 195756 302360
rect 196104 302012 196736 302360
rect 112708 167312 196736 302012
rect 112708 166964 195076 167312
rect 195424 166964 196736 167312
rect 112708 165652 196736 166964
rect 112708 165292 116960 165652
rect 111988 164932 116960 165292
rect 111988 164572 114240 164932
rect 110076 159100 114240 164572
rect 110076 158432 111628 159100
rect 110076 153824 110476 158432
rect 111148 153824 111628 158432
rect 110076 19600 111628 153824
rect 111988 158740 114240 159100
rect 114912 158740 116960 164932
rect 111988 158380 116960 158740
rect 111988 20320 112348 158380
rect 112708 158020 116960 158380
rect 117632 164932 127840 165652
rect 117632 158740 125120 164932
rect 125792 158740 127840 164932
rect 117632 158020 127840 158740
rect 128512 164932 138720 165652
rect 128512 158740 136000 164932
rect 136672 158740 138720 164932
rect 128512 158020 138720 158740
rect 139392 164932 149600 165652
rect 139392 158740 146880 164932
rect 147552 158740 149600 164932
rect 139392 158020 149600 158740
rect 150272 164932 160480 165652
rect 150272 158740 157760 164932
rect 158432 158740 160480 164932
rect 150272 158020 160480 158740
rect 161152 164932 171360 165652
rect 161152 158740 162704 164932
rect 163376 158740 168640 164932
rect 169312 158740 171360 164932
rect 161152 158020 171360 158740
rect 172032 164932 182240 165652
rect 172032 158740 179520 164932
rect 180192 158740 182240 164932
rect 172032 158020 182240 158740
rect 182912 164932 193120 165652
rect 182912 158740 190400 164932
rect 191072 158740 193120 164932
rect 182912 158020 193120 158740
rect 193792 165292 196736 165652
rect 197096 165292 197456 303352
rect 193792 164572 197456 165292
rect 197816 164572 201280 304072
rect 193792 159100 201280 164572
rect 193792 158380 197456 159100
rect 193792 158020 196736 158380
rect 112708 157388 196736 158020
rect 112708 157040 195756 157388
rect 196104 157040 196736 157388
rect 112708 156708 196736 157040
rect 112708 156360 195076 156708
rect 195424 156360 196736 156708
rect 112708 20680 196736 156360
rect 112708 20320 116960 20680
rect 111988 19960 116960 20320
rect 111988 19600 114240 19960
rect 110076 816 114240 19600
rect 114912 3264 116960 19960
rect 117632 19960 127840 20680
rect 117632 3264 125120 19960
rect 114912 816 125120 3264
rect 125792 3264 127840 19960
rect 128512 19960 138720 20680
rect 128512 3264 136000 19960
rect 125792 816 136000 3264
rect 136672 3264 138720 19960
rect 139392 19960 149600 20680
rect 139392 3264 146880 19960
rect 136672 816 146880 3264
rect 147552 3264 149600 19960
rect 150272 19960 160480 20680
rect 150272 3264 157760 19960
rect 147552 816 157760 3264
rect 158432 3264 160480 19960
rect 161152 19960 171360 20680
rect 161152 3264 162704 19960
rect 158432 816 162704 3264
rect 163376 816 168640 19960
rect 169312 3264 171360 19960
rect 172032 19960 182240 20680
rect 172032 3264 179520 19960
rect 169312 816 179520 3264
rect 180192 3264 182240 19960
rect 182912 19960 193120 20680
rect 182912 3264 190400 19960
rect 180192 816 190400 3264
rect 191072 3264 193120 19960
rect 193792 20320 196736 20680
rect 197096 20320 197456 158380
rect 193792 19600 197456 20320
rect 197816 158432 201280 159100
rect 197816 153824 198296 158432
rect 198968 153824 201280 158432
rect 197816 19600 201280 153824
rect 193792 3264 201280 19600
rect 191072 816 201280 3264
rect 201952 3264 204000 315904
rect 204672 315904 214880 316624
rect 204672 197448 212160 315904
rect 204672 111260 209288 197448
rect 209648 197088 212160 197448
rect 212832 197088 214880 315904
rect 209648 196728 214880 197088
rect 209648 111980 210008 196728
rect 210368 196368 214880 196728
rect 215552 315904 225760 316624
rect 215552 197088 223040 315904
rect 223712 197088 225760 315904
rect 215552 196368 225760 197088
rect 226432 315904 236640 316624
rect 226432 197088 233920 315904
rect 234592 197088 236640 315904
rect 226432 196368 236640 197088
rect 237312 315904 247520 316624
rect 237312 197088 244800 315904
rect 245472 197088 247520 315904
rect 237312 196368 247520 197088
rect 248192 315904 258400 316624
rect 248192 197088 255680 315904
rect 256352 197088 258400 315904
rect 248192 196368 258400 197088
rect 259072 315904 269280 316624
rect 259072 197088 266560 315904
rect 267232 197088 269280 315904
rect 259072 196368 269280 197088
rect 269952 315904 280160 316624
rect 269952 197088 277440 315904
rect 278112 197088 280160 315904
rect 269952 196368 280160 197088
rect 280832 315904 291040 316624
rect 280832 197088 288320 315904
rect 288992 197088 291040 315904
rect 280832 196368 291040 197088
rect 291712 315904 301920 316624
rect 291712 197088 299200 315904
rect 299872 197088 301920 315904
rect 291712 196368 301920 197088
rect 302592 316264 303360 316624
rect 303720 316264 304080 401012
rect 302592 315544 304080 316264
rect 304440 315544 310080 401732
rect 302592 197088 310080 315544
rect 310752 509728 320960 512176
rect 310752 197088 312800 509728
rect 302592 196368 312800 197088
rect 313472 493392 320960 509728
rect 313472 353892 315912 493392
rect 316272 493032 320960 493392
rect 321632 509728 331840 512176
rect 321632 493032 323680 509728
rect 316272 492672 323680 493032
rect 316272 354612 316632 492672
rect 316992 492312 323680 492672
rect 324352 493032 331840 509728
rect 332512 509728 342720 512176
rect 332512 493032 334560 509728
rect 324352 492312 334560 493032
rect 335232 493032 342720 509728
rect 343392 509728 352104 512176
rect 343392 493032 345440 509728
rect 335232 492312 345440 493032
rect 346112 492312 350304 509728
rect 350976 493032 352104 509728
rect 352776 493032 353600 512176
rect 354272 509728 364480 512176
rect 354272 493032 356320 509728
rect 350976 492312 356320 493032
rect 356992 493032 364480 509728
rect 365152 509728 375360 512176
rect 365152 493032 367200 509728
rect 356992 492312 367200 493032
rect 367872 493032 375360 509728
rect 376032 509728 386240 512176
rect 376032 493032 378080 509728
rect 367872 492312 378080 493032
rect 378752 493032 386240 509728
rect 386912 509728 397120 512176
rect 386912 493032 388960 509728
rect 378752 492312 388960 493032
rect 389632 493032 397120 509728
rect 397792 509728 405504 512176
rect 397792 493032 399840 509728
rect 389632 492312 399840 493032
rect 400512 493392 403704 509728
rect 400512 492672 401740 493392
rect 400512 492312 401020 492672
rect 316992 491680 401020 492312
rect 316992 491332 400040 491680
rect 400388 491332 401020 491680
rect 316992 356632 401020 491332
rect 316992 356284 318304 356632
rect 318652 356284 401020 356632
rect 316992 354972 401020 356284
rect 316992 354612 323680 354972
rect 316272 354252 323680 354612
rect 316272 353892 320960 354252
rect 313472 348420 320960 353892
rect 313472 208920 315912 348420
rect 316272 348060 320960 348420
rect 321632 348060 323680 354252
rect 316272 347700 323680 348060
rect 316272 209640 316632 347700
rect 316992 347340 323680 347700
rect 324352 354252 334560 354972
rect 324352 348060 331840 354252
rect 332512 348060 334560 354252
rect 324352 347340 334560 348060
rect 335232 354252 345440 354972
rect 335232 348060 342720 354252
rect 343392 348060 345440 354252
rect 335232 347340 345440 348060
rect 346112 347340 350304 354972
rect 350976 354252 356320 354972
rect 350976 348060 352104 354252
rect 352776 348060 353600 354252
rect 354272 348060 356320 354252
rect 350976 347340 356320 348060
rect 356992 354252 367200 354972
rect 356992 348060 364480 354252
rect 365152 348060 367200 354252
rect 356992 347340 367200 348060
rect 367872 354252 378080 354972
rect 367872 348060 375360 354252
rect 376032 348060 378080 354252
rect 367872 347340 378080 348060
rect 378752 354252 388960 354972
rect 378752 348060 386240 354252
rect 386912 348060 388960 354252
rect 378752 347340 388960 348060
rect 389632 354252 399840 354972
rect 389632 348060 397120 354252
rect 397792 348060 399840 354252
rect 389632 347340 399840 348060
rect 400512 354612 401020 354972
rect 401380 354612 401740 492672
rect 400512 353892 401740 354612
rect 402100 353892 403704 493392
rect 400512 348420 403704 353892
rect 400512 347700 401740 348420
rect 400512 347340 401020 347700
rect 316992 211660 401020 347340
rect 316992 211312 318304 211660
rect 318652 211312 401020 211660
rect 316992 210980 401020 211312
rect 316992 210632 400040 210980
rect 400388 210632 401020 210980
rect 316992 210000 401020 210632
rect 316992 209640 323680 210000
rect 316272 209280 323680 209640
rect 316272 208920 320960 209280
rect 313472 197088 320960 208920
rect 321632 197088 323680 209280
rect 313472 196368 323680 197088
rect 324352 209280 334560 210000
rect 324352 197088 331840 209280
rect 332512 197088 334560 209280
rect 324352 196368 334560 197088
rect 335232 209280 345440 210000
rect 335232 197088 342720 209280
rect 343392 197088 345440 209280
rect 335232 196368 345440 197088
rect 346112 197448 350304 210000
rect 346112 196728 348428 197448
rect 346112 196368 347708 196728
rect 210368 195056 347708 196368
rect 210368 194708 346048 195056
rect 346396 194708 347708 195056
rect 210368 113320 347708 194708
rect 210368 112972 346728 113320
rect 347076 112972 347708 113320
rect 210368 112340 347708 112972
rect 210368 111980 214880 112340
rect 209648 111620 214880 111980
rect 209648 111260 212160 111620
rect 204672 105788 212160 111260
rect 204672 19600 209288 105788
rect 209648 105428 212160 105788
rect 212832 105428 214880 111620
rect 209648 105068 214880 105428
rect 209648 20320 210008 105068
rect 210368 104708 214880 105068
rect 215552 111620 225760 112340
rect 215552 105428 223040 111620
rect 223712 105428 225760 111620
rect 215552 104708 225760 105428
rect 226432 111620 236640 112340
rect 226432 105428 233920 111620
rect 234592 105428 236640 111620
rect 226432 104708 236640 105428
rect 237312 111620 247520 112340
rect 237312 105428 244800 111620
rect 245472 105428 247520 111620
rect 237312 104708 247520 105428
rect 248192 111620 258400 112340
rect 248192 105428 255680 111620
rect 256352 105428 258400 111620
rect 248192 104708 258400 105428
rect 259072 111620 269280 112340
rect 259072 105428 266560 111620
rect 267232 105428 269280 111620
rect 259072 104708 269280 105428
rect 269952 111620 280160 112340
rect 269952 105428 277440 111620
rect 278112 105428 280160 111620
rect 269952 104708 280160 105428
rect 280832 111620 291040 112340
rect 280832 105428 288320 111620
rect 288992 105428 291040 111620
rect 280832 104708 291040 105428
rect 291712 111620 301920 112340
rect 291712 105428 299200 111620
rect 299872 105428 301920 111620
rect 291712 104708 301920 105428
rect 302592 111620 312800 112340
rect 302592 105428 310080 111620
rect 310752 105428 312800 111620
rect 302592 104708 312800 105428
rect 313472 111620 323680 112340
rect 313472 105428 320960 111620
rect 321632 105428 323680 111620
rect 313472 104708 323680 105428
rect 324352 111620 334560 112340
rect 324352 105428 331840 111620
rect 332512 105428 334560 111620
rect 324352 104708 334560 105428
rect 335232 111620 345440 112340
rect 335232 105428 342720 111620
rect 343392 105428 345440 111620
rect 335232 104708 345440 105428
rect 346112 111980 347708 112340
rect 348068 111980 348428 196728
rect 346112 111260 348428 111980
rect 348788 111260 350304 197448
rect 346112 105788 350304 111260
rect 346112 105068 348428 105788
rect 346112 104708 347708 105068
rect 210368 103396 347708 104708
rect 210368 103048 346048 103396
rect 346396 103048 347708 103396
rect 210368 21660 347708 103048
rect 210368 21312 346728 21660
rect 347076 21312 347708 21660
rect 210368 20680 347708 21312
rect 210368 20320 214880 20680
rect 209648 19960 214880 20320
rect 209648 19600 212160 19960
rect 204672 3264 212160 19600
rect 201952 816 212160 3264
rect 212832 3264 214880 19960
rect 215552 19960 225760 20680
rect 215552 3264 223040 19960
rect 212832 816 223040 3264
rect 223712 3264 225760 19960
rect 226432 19960 236640 20680
rect 226432 3264 233920 19960
rect 223712 816 233920 3264
rect 234592 3264 236640 19960
rect 237312 19960 247520 20680
rect 237312 3264 244800 19960
rect 234592 816 244800 3264
rect 245472 3264 247520 19960
rect 248192 19960 258400 20680
rect 248192 3264 255680 19960
rect 245472 816 255680 3264
rect 256352 3264 258400 19960
rect 259072 19960 269280 20680
rect 259072 3264 266560 19960
rect 256352 816 266560 3264
rect 267232 3264 269280 19960
rect 269952 19960 280160 20680
rect 269952 3264 277440 19960
rect 267232 816 277440 3264
rect 278112 3264 280160 19960
rect 280832 19960 291040 20680
rect 280832 3264 288320 19960
rect 278112 816 288320 3264
rect 288992 3264 291040 19960
rect 291712 19960 301920 20680
rect 291712 3264 299200 19960
rect 288992 816 299200 3264
rect 299872 3264 301920 19960
rect 302592 19960 312800 20680
rect 302592 3264 310080 19960
rect 299872 816 310080 3264
rect 310752 3264 312800 19960
rect 313472 19960 323680 20680
rect 313472 3264 320960 19960
rect 310752 816 320960 3264
rect 321632 3264 323680 19960
rect 324352 19960 334560 20680
rect 324352 3264 331840 19960
rect 321632 816 331840 3264
rect 332512 3264 334560 19960
rect 335232 19960 345440 20680
rect 335232 3264 342720 19960
rect 332512 816 342720 3264
rect 343392 3264 345440 19960
rect 346112 20320 347708 20680
rect 348068 20320 348428 105068
rect 346112 19600 348428 20320
rect 348788 19600 350304 105788
rect 346112 3264 350304 19600
rect 350976 209280 356320 210000
rect 350976 3264 352104 209280
rect 343392 816 352104 3264
rect 352776 197088 353600 209280
rect 354272 197448 356320 209280
rect 352776 111620 354260 197088
rect 354620 196728 356320 197448
rect 354620 111980 354980 196728
rect 355340 196368 356320 196728
rect 356992 209280 367200 210000
rect 356992 197088 364480 209280
rect 365152 197088 367200 209280
rect 356992 196368 367200 197088
rect 367872 209280 378080 210000
rect 367872 197088 375360 209280
rect 376032 197088 378080 209280
rect 367872 196368 378080 197088
rect 378752 209280 388960 210000
rect 378752 197088 386240 209280
rect 386912 197088 388960 209280
rect 378752 196368 388960 197088
rect 389632 209280 399840 210000
rect 389632 197088 397120 209280
rect 397792 197088 399840 209280
rect 389632 196368 399840 197088
rect 400512 209640 401020 210000
rect 401380 209640 401740 347700
rect 400512 208920 401740 209640
rect 402100 208920 403704 348420
rect 400512 196368 403704 208920
rect 404376 197088 405504 509728
rect 406176 493872 408000 512176
rect 408672 509728 418880 512176
rect 408672 493872 410720 509728
rect 406176 493392 410720 493872
rect 406176 353892 407572 493392
rect 407932 492672 410720 493392
rect 407932 354612 408292 492672
rect 408652 492312 410720 492672
rect 411392 493032 418880 509728
rect 419552 509728 429760 512176
rect 419552 493032 421600 509728
rect 411392 492312 421600 493032
rect 422272 493032 429760 509728
rect 430432 509728 440640 512176
rect 430432 493032 432480 509728
rect 422272 492312 432480 493032
rect 433152 493032 440640 509728
rect 441312 509728 451520 512176
rect 441312 493032 443360 509728
rect 433152 492312 443360 493032
rect 444032 493032 451520 509728
rect 452192 509728 462400 512176
rect 452192 493032 454240 509728
rect 444032 492312 454240 493032
rect 454912 493032 462400 509728
rect 463072 509728 473280 512176
rect 463072 493032 465120 509728
rect 454912 492312 465120 493032
rect 465792 493032 473280 509728
rect 473952 509728 484160 512176
rect 473952 493032 476000 509728
rect 465792 492312 476000 493032
rect 476672 493032 484160 509728
rect 484832 509728 495040 512176
rect 484832 493032 486880 509728
rect 476672 492312 486880 493032
rect 487552 493392 495040 509728
rect 487552 492672 493400 493392
rect 487552 492312 492680 492672
rect 408652 491000 492680 492312
rect 408652 490652 491020 491000
rect 491368 490652 492680 491000
rect 408652 355952 492680 490652
rect 408652 355604 491700 355952
rect 492048 355604 492680 355952
rect 408652 354972 492680 355604
rect 408652 354612 410720 354972
rect 407932 353892 410720 354612
rect 406176 351554 410720 353892
rect 406176 350880 408000 351554
rect 408672 350880 410720 351554
rect 406176 348420 410720 350880
rect 406176 208920 407572 348420
rect 407932 347700 410720 348420
rect 407932 209640 408292 347700
rect 408652 347340 410720 347700
rect 411392 354252 421600 354972
rect 411392 348060 418880 354252
rect 419552 348060 421600 354252
rect 411392 347340 421600 348060
rect 422272 354252 432480 354972
rect 422272 348060 429760 354252
rect 430432 348060 432480 354252
rect 422272 347340 432480 348060
rect 433152 354252 443360 354972
rect 433152 348060 440640 354252
rect 441312 348060 443360 354252
rect 433152 347340 443360 348060
rect 444032 354252 454240 354972
rect 444032 348060 451520 354252
rect 452192 348060 454240 354252
rect 444032 347340 454240 348060
rect 454912 354252 465120 354972
rect 454912 348060 462400 354252
rect 463072 348060 465120 354252
rect 454912 347340 465120 348060
rect 465792 354252 476000 354972
rect 465792 348060 473280 354252
rect 473952 348060 476000 354252
rect 465792 347340 476000 348060
rect 476672 354252 486880 354972
rect 476672 348060 484160 354252
rect 484832 348060 486880 354252
rect 476672 347340 486880 348060
rect 487552 354612 492680 354972
rect 493040 354612 493400 492672
rect 487552 353892 493400 354612
rect 493760 353892 495040 493392
rect 487552 348420 495040 353892
rect 487552 347700 493400 348420
rect 487552 347340 492680 347700
rect 408652 211660 492680 347340
rect 408652 211312 491020 211660
rect 491368 211312 492680 211660
rect 408652 210980 492680 211312
rect 408652 210632 491700 210980
rect 492048 210632 492680 210980
rect 408652 210000 492680 210632
rect 408652 209640 410720 210000
rect 407932 208920 410720 209640
rect 406176 208440 410720 208920
rect 406176 197088 408000 208440
rect 408672 197088 410720 208440
rect 404376 196368 410720 197088
rect 411392 209280 421600 210000
rect 411392 197088 418880 209280
rect 419552 197088 421600 209280
rect 411392 196368 421600 197088
rect 422272 209280 432480 210000
rect 422272 197088 429760 209280
rect 430432 197088 432480 209280
rect 422272 196368 432480 197088
rect 433152 209280 443360 210000
rect 433152 197088 440640 209280
rect 441312 197088 443360 209280
rect 433152 196368 443360 197088
rect 444032 209280 454240 210000
rect 444032 197088 451520 209280
rect 452192 197088 454240 209280
rect 444032 196368 454240 197088
rect 454912 209280 465120 210000
rect 454912 197088 462400 209280
rect 463072 197088 465120 209280
rect 454912 196368 465120 197088
rect 465792 209280 476000 210000
rect 465792 197088 473280 209280
rect 473952 197088 476000 209280
rect 465792 196368 476000 197088
rect 476672 209280 486880 210000
rect 476672 197088 484160 209280
rect 484832 197088 486880 209280
rect 476672 196368 486880 197088
rect 487552 209640 492680 210000
rect 493040 209640 493400 347700
rect 487552 208920 493400 209640
rect 493760 208920 495040 348420
rect 487552 197448 495040 208920
rect 487552 196728 493400 197448
rect 487552 196368 492680 196728
rect 355340 195736 492680 196368
rect 355340 195388 491700 195736
rect 492048 195388 492680 195736
rect 355340 195056 492680 195388
rect 355340 194708 356652 195056
rect 357000 194708 492680 195056
rect 355340 112340 492680 194708
rect 355340 111980 356320 112340
rect 352776 105428 353600 111620
rect 354620 111260 356320 111980
rect 354272 105788 356320 111260
rect 352776 19960 354260 105428
rect 354620 105068 356320 105788
rect 354620 20320 354980 105068
rect 355340 104708 356320 105068
rect 356992 111620 367200 112340
rect 356992 105428 364480 111620
rect 365152 105428 367200 111620
rect 356992 104708 367200 105428
rect 367872 111620 378080 112340
rect 367872 105428 375360 111620
rect 376032 105428 378080 111620
rect 367872 104708 378080 105428
rect 378752 111620 388960 112340
rect 378752 105428 386240 111620
rect 386912 105428 388960 111620
rect 378752 104708 388960 105428
rect 389632 111620 399840 112340
rect 389632 105428 397120 111620
rect 397792 105428 399840 111620
rect 389632 104708 399840 105428
rect 400512 104708 403704 112340
rect 404376 111620 410720 112340
rect 404376 105428 405504 111620
rect 406176 105428 408000 111620
rect 408672 105428 410720 111620
rect 404376 104708 410720 105428
rect 411392 111620 421600 112340
rect 411392 105428 418880 111620
rect 419552 105428 421600 111620
rect 411392 104708 421600 105428
rect 422272 111620 432480 112340
rect 422272 105428 429760 111620
rect 430432 105428 432480 111620
rect 422272 104708 432480 105428
rect 433152 111620 443360 112340
rect 433152 105428 440640 111620
rect 441312 105428 443360 111620
rect 433152 104708 443360 105428
rect 444032 111620 454240 112340
rect 444032 105428 451520 111620
rect 452192 105428 454240 111620
rect 444032 104708 454240 105428
rect 454912 111620 465120 112340
rect 454912 105428 462400 111620
rect 463072 105428 465120 111620
rect 454912 104708 465120 105428
rect 465792 111620 476000 112340
rect 465792 105428 473280 111620
rect 473952 105428 476000 111620
rect 465792 104708 476000 105428
rect 476672 111620 486880 112340
rect 476672 105428 484160 111620
rect 484832 105428 486880 111620
rect 476672 104708 486880 105428
rect 487552 111980 492680 112340
rect 493040 111980 493400 196728
rect 487552 111260 493400 111980
rect 493760 111260 495040 197448
rect 487552 105788 495040 111260
rect 487552 105068 493400 105788
rect 487552 104708 492680 105068
rect 355340 103396 492680 104708
rect 355340 103048 356652 103396
rect 357000 103048 492680 103396
rect 355340 21660 492680 103048
rect 355340 21312 491700 21660
rect 492048 21312 492680 21660
rect 355340 20680 492680 21312
rect 355340 20320 356320 20680
rect 352776 816 353600 19960
rect 354620 19600 356320 20320
rect 354272 3264 356320 19600
rect 356992 19960 367200 20680
rect 356992 3264 364480 19960
rect 354272 816 364480 3264
rect 365152 3264 367200 19960
rect 367872 19960 378080 20680
rect 367872 3264 375360 19960
rect 365152 816 375360 3264
rect 376032 3264 378080 19960
rect 378752 19960 388960 20680
rect 378752 3264 386240 19960
rect 376032 816 386240 3264
rect 386912 3264 388960 19960
rect 389632 19960 399840 20680
rect 389632 3264 397120 19960
rect 386912 816 397120 3264
rect 397792 3264 399840 19960
rect 400512 3264 403704 20680
rect 404376 19960 410720 20680
rect 404376 3264 405504 19960
rect 397792 816 405504 3264
rect 406176 816 408000 19960
rect 408672 3264 410720 19960
rect 411392 19960 421600 20680
rect 411392 3264 418880 19960
rect 408672 816 418880 3264
rect 419552 3264 421600 19960
rect 422272 19960 432480 20680
rect 422272 3264 429760 19960
rect 419552 816 429760 3264
rect 430432 3264 432480 19960
rect 433152 19960 443360 20680
rect 433152 3264 440640 19960
rect 430432 816 440640 3264
rect 441312 3264 443360 19960
rect 444032 19960 454240 20680
rect 444032 3264 451520 19960
rect 441312 816 451520 3264
rect 452192 3264 454240 19960
rect 454912 19960 465120 20680
rect 454912 3264 462400 19960
rect 452192 816 462400 3264
rect 463072 3264 465120 19960
rect 465792 19960 476000 20680
rect 465792 3264 473280 19960
rect 463072 816 473280 3264
rect 473952 3264 476000 19960
rect 476672 19960 486880 20680
rect 476672 3264 484160 19960
rect 473952 816 484160 3264
rect 484832 3264 486880 19960
rect 487552 20320 492680 20680
rect 493040 20320 493400 105068
rect 487552 19600 493400 20320
rect 493760 19600 495040 105788
rect 487552 3264 495040 19600
rect 484832 816 495040 3264
rect 495712 509728 505920 512176
rect 495712 3264 497760 509728
rect 498432 3264 505920 509728
rect 495712 816 505920 3264
rect 506592 816 508840 512176
rect 4888 0 508840 816
rect 510472 0 511288 512992
rect 512920 0 513728 512992
<< metal5 >>
rect 0 510544 513728 512176
rect 0 508096 513728 509728
rect 3256 505920 510472 506592
rect 808 503200 512920 503872
rect 3256 495040 510472 495712
rect 19968 493032 159468 493392
rect 164940 493032 304440 493392
rect 315912 493032 402100 493392
rect 407572 493032 493760 493392
rect 808 492320 16992 492992
rect 20688 492312 158748 492672
rect 165660 492312 303720 492672
rect 310077 492320 310752 492992
rect 316632 492312 401380 492672
rect 408292 492312 493040 492672
rect 495040 492320 512920 492992
rect 19968 491332 22028 491680
rect 20688 490652 22708 491000
rect 167332 490652 167680 492312
rect 302380 491332 304440 491680
rect 400040 491332 402100 491680
rect 491020 490652 493040 491000
rect 3256 484160 21048 484832
rect 158388 484160 166020 484832
rect 303360 484160 316992 484832
rect 401020 484160 408652 484832
rect 492680 484160 510472 484832
rect 808 481440 20328 482112
rect 159108 481440 165300 482112
rect 304080 481440 316272 482112
rect 401740 481440 407932 482112
rect 493400 481440 512920 482112
rect 3256 473280 21048 473952
rect 158388 473280 166020 473952
rect 303360 473280 316992 473952
rect 401020 473280 408652 473952
rect 492680 473280 510472 473952
rect 808 470560 20328 471232
rect 159108 470560 165300 471232
rect 304080 470560 316272 471232
rect 401740 470560 407932 471232
rect 493400 470560 512920 471232
rect 3256 462400 21048 463072
rect 158388 462400 166020 463072
rect 303360 462400 316992 463072
rect 401020 462400 408652 463072
rect 492680 462400 510472 463072
rect 808 459680 20328 460352
rect 159108 459680 165300 460352
rect 304080 459680 316272 460352
rect 401740 459680 407932 460352
rect 493400 459680 512920 460352
rect 3256 451520 21048 452192
rect 158388 451520 166020 452192
rect 303360 451520 316992 452192
rect 401020 451520 408652 452192
rect 492680 451520 510472 452192
rect 808 448800 20328 449472
rect 159108 448800 165300 449472
rect 304080 448800 316272 449472
rect 401740 448800 407932 449472
rect 493400 448800 512920 449472
rect 3256 440640 21048 441312
rect 158388 440640 166020 441312
rect 303360 440640 316992 441312
rect 401020 440640 408652 441312
rect 492680 440640 510472 441312
rect 808 437920 20328 438592
rect 159108 437920 165300 438592
rect 304080 437920 316272 438592
rect 401740 437920 407932 438592
rect 493400 437920 512920 438592
rect 3256 429760 21048 430432
rect 158388 429760 166020 430432
rect 303360 429760 316992 430432
rect 401020 429760 408652 430432
rect 492680 429760 510472 430432
rect 808 427040 20328 427712
rect 159108 427040 165300 427712
rect 304080 427040 316272 427712
rect 401740 427040 407932 427712
rect 493400 427040 512920 427712
rect 3256 418880 21048 419552
rect 158388 418880 166020 419552
rect 303360 418880 316992 419552
rect 401020 418880 408652 419552
rect 492680 418880 510472 419552
rect 808 416160 20328 416832
rect 159108 416160 165300 416832
rect 304080 416160 316272 416832
rect 401740 416160 407932 416832
rect 493400 416160 512920 416832
rect 3256 408284 21048 408672
rect 158388 408284 166020 408672
rect 303360 408284 316992 408672
rect 3256 408000 316992 408284
rect 401020 408000 408652 408672
rect 492680 408000 510472 408672
rect 20688 407924 158748 408000
rect 165660 407924 303720 408000
rect 19968 407204 159468 407564
rect 164940 407204 304440 407564
rect 808 405280 316272 405952
rect 401740 405280 407932 405952
rect 493400 405280 512920 405952
rect 19968 401372 159468 401732
rect 164940 401372 304440 401732
rect 20688 400652 158748 401012
rect 165660 400652 303720 401012
rect 19968 399672 22028 400020
rect 164940 399672 167000 400020
rect 20688 398992 22708 399340
rect 301700 398992 302048 400652
rect 3256 397120 21048 397792
rect 158388 397120 166020 397792
rect 303360 397120 316992 397792
rect 401020 397120 408652 397792
rect 492680 397120 510472 397792
rect 808 394400 20328 395072
rect 159108 394400 165300 395072
rect 304080 394400 316272 395072
rect 401740 394400 407932 395072
rect 493400 394400 512920 395072
rect 3256 386240 21048 386912
rect 158388 386240 166020 386912
rect 303360 386240 316992 386912
rect 401020 386240 408652 386912
rect 492680 386240 510472 386912
rect 808 383520 20328 384192
rect 159108 383520 165300 384192
rect 304080 383520 316272 384192
rect 401740 383520 407932 384192
rect 493400 383520 512920 384192
rect 3256 375360 21048 376032
rect 158388 375360 166020 376032
rect 303360 375360 316992 376032
rect 401020 375360 408652 376032
rect 492680 375360 510472 376032
rect 808 372640 20328 373312
rect 159108 372640 165300 373312
rect 304080 372640 316272 373312
rect 401740 372640 407932 373312
rect 493400 372640 512920 373312
rect 3256 364480 21048 365152
rect 158388 364480 166020 365152
rect 303360 364480 316992 365152
rect 401020 364480 408652 365152
rect 492680 364480 510472 365152
rect 808 361760 20328 362432
rect 159108 361760 165300 362432
rect 304080 361760 316272 362432
rect 401740 361760 407932 362432
rect 493400 361760 512920 362432
rect 316632 356284 318652 356632
rect 491700 355604 493760 355952
rect 316632 354612 401380 354972
rect 408292 354612 493040 354972
rect 3256 353600 21048 354272
rect 158388 353600 166020 354272
rect 303360 353600 313472 354272
rect 315912 353892 402100 354252
rect 407572 353892 493760 354252
rect 497760 353600 510472 354272
rect 808 350880 20328 351552
rect 159108 350880 165300 351552
rect 304080 350880 512920 351552
rect 315912 348060 402100 348420
rect 407572 348060 493760 348420
rect 316632 347340 401380 347700
rect 408292 347340 493040 347700
rect 3256 342720 21048 343392
rect 158388 342720 166020 343392
rect 303360 342720 316992 343392
rect 401020 342720 408652 343392
rect 492680 342720 510472 343392
rect 808 340000 20328 340672
rect 159108 340000 165300 340672
rect 304080 340000 316272 340672
rect 401740 340000 407932 340672
rect 493400 340000 512920 340672
rect 3256 331840 21048 332512
rect 158388 331840 166020 332512
rect 303360 331840 316992 332512
rect 401020 331840 408652 332512
rect 492680 331840 510472 332512
rect 808 329120 20328 329792
rect 159108 329120 165300 329792
rect 304080 329120 316272 329792
rect 401740 329120 407932 329792
rect 493400 329120 512920 329792
rect 3256 320960 21048 321632
rect 158388 320960 166020 321632
rect 303360 320960 316992 321632
rect 401020 320960 408652 321632
rect 492680 320960 510472 321632
rect 808 318240 20328 318912
rect 159108 318240 165300 318912
rect 304080 318240 316272 318912
rect 401740 318240 407932 318912
rect 493400 318240 512920 318912
rect 20688 316264 158748 316624
rect 165660 316264 303720 316624
rect 19968 315544 159468 315904
rect 164940 315544 304440 315904
rect 3256 310080 316992 310752
rect 401020 310080 408652 310752
rect 492680 310080 510472 310752
rect 808 307360 316272 308032
rect 401740 307360 407932 308032
rect 493400 307360 512920 308032
rect 19968 303712 106156 304072
rect 111628 303712 197816 304072
rect 20688 302992 105436 303352
rect 112348 302992 197096 303352
rect 19968 302012 22028 302360
rect 195756 302012 197816 302360
rect 3256 299200 21048 299872
rect 105076 299200 112708 299872
rect 196736 299200 316992 299872
rect 401020 299200 408652 299872
rect 492680 299200 510472 299872
rect 808 296480 20328 297152
rect 105796 296480 111988 297152
rect 197456 296480 316272 297152
rect 401740 296480 407932 297152
rect 493400 296480 512920 297152
rect 3256 288320 21048 288992
rect 105076 288320 112708 288992
rect 196736 288320 316992 288992
rect 401020 288320 408652 288992
rect 492680 288320 510472 288992
rect 808 285600 20328 286272
rect 105796 285600 111988 286272
rect 197456 285600 316272 286272
rect 401740 285600 407932 286272
rect 493400 285600 512920 286272
rect 3256 277440 21048 278112
rect 105076 277440 112708 278112
rect 196736 277440 316992 278112
rect 401020 277440 408652 278112
rect 492680 277440 510472 278112
rect 808 274720 20328 275392
rect 105796 274720 111988 275392
rect 197456 274720 316272 275392
rect 401740 274720 407932 275392
rect 493400 274720 512920 275392
rect 3256 266560 21048 267232
rect 105076 266560 112708 267232
rect 196736 266560 316992 267232
rect 401020 266560 408652 267232
rect 492680 266560 510472 267232
rect 808 263840 20328 264512
rect 105796 263840 111988 264512
rect 197456 263840 316272 264512
rect 401740 263840 407932 264512
rect 493400 263840 512920 264512
rect 3256 255680 21048 256352
rect 105076 255680 112708 256352
rect 196736 255680 316992 256352
rect 401020 255680 408652 256352
rect 492680 255680 510472 256352
rect 808 252960 20328 253632
rect 105796 252960 111988 253632
rect 197456 252960 316272 253632
rect 401740 252960 407932 253632
rect 493400 252960 512920 253632
rect 3256 244800 21048 245472
rect 105076 244800 112708 245472
rect 196736 244800 316992 245472
rect 401020 244800 408652 245472
rect 492680 244800 510472 245472
rect 808 242080 20328 242752
rect 105796 242080 111988 242752
rect 197456 242080 316272 242752
rect 401740 242080 407932 242752
rect 493400 242080 512920 242752
rect 3256 233920 21048 234592
rect 105076 233920 112708 234592
rect 196736 233920 316992 234592
rect 401020 233920 408652 234592
rect 492680 233920 510472 234592
rect 808 231200 20328 231872
rect 105796 231200 111988 231872
rect 197456 231200 316272 231872
rect 401740 231200 407932 231872
rect 493400 231200 512920 231872
rect 3256 223040 21048 223712
rect 105076 223040 112708 223712
rect 196736 223040 316992 223712
rect 401020 223040 408652 223712
rect 492680 223040 510472 223712
rect 808 220320 20328 220992
rect 105796 220320 111988 220992
rect 197456 220320 316272 220992
rect 401740 220320 407932 220992
rect 493400 220320 512920 220992
rect 3256 212160 21048 212832
rect 105076 212160 112708 212832
rect 196736 212160 316992 212832
rect 401020 212160 408652 212832
rect 492680 212160 510472 212832
rect 316632 211312 318652 211660
rect 491020 211312 493040 211660
rect 400040 210632 402100 210980
rect 491700 210632 493760 210980
rect 808 209440 20328 210112
rect 105796 209440 111988 210112
rect 197456 209440 310753 210112
rect 316632 209640 401380 210000
rect 408292 209640 493040 210000
rect 495040 209440 512920 210112
rect 315912 208920 402100 209280
rect 407572 208920 493760 209280
rect 3256 201280 21048 201952
rect 105076 201280 112708 201952
rect 196736 201280 510472 201952
rect 808 198560 20328 199232
rect 105796 198560 111988 199232
rect 197456 198560 512920 199232
rect 209288 197088 348788 197448
rect 353600 197088 493760 197448
rect 210008 196368 348068 196728
rect 354980 196368 493040 196728
rect 346048 194708 346396 196368
rect 356652 194708 357000 196368
rect 491700 195388 493760 195736
rect 3256 190400 21048 191072
rect 105076 190400 112708 191072
rect 196736 190400 210368 191072
rect 347708 190400 355340 191072
rect 492680 190400 510472 191072
rect 808 187680 20328 188352
rect 105796 187680 111988 188352
rect 197456 187680 209648 188352
rect 348428 187680 354620 188352
rect 493400 187680 512920 188352
rect 3256 179520 21048 180192
rect 105076 179520 112708 180192
rect 196736 179520 210368 180192
rect 347708 179520 355340 180192
rect 492680 179520 510472 180192
rect 808 176800 20328 177472
rect 105796 176800 111988 177472
rect 197456 176800 209648 177472
rect 348428 176800 354620 177472
rect 493400 176800 512920 177472
rect 3256 168640 21048 169312
rect 105076 168640 112708 169312
rect 196736 168640 210368 169312
rect 347708 168640 355340 169312
rect 492680 168640 510472 169312
rect 20688 166964 22708 167312
rect 195076 166964 197096 167312
rect 808 165920 20328 166592
rect 105796 165920 111988 166592
rect 197456 165920 209648 166592
rect 348428 165920 354620 166592
rect 493400 165920 512920 166592
rect 20688 165292 105436 165652
rect 112348 165292 197096 165652
rect 19968 164572 106156 164932
rect 111628 164572 197816 164932
rect 19968 158740 106156 159100
rect 111628 158740 197816 159100
rect 3256 157760 19488 158432
rect 20688 158020 105436 158380
rect 106636 157760 111148 158432
rect 112348 158020 197096 158380
rect 198296 157760 210368 158432
rect 347708 157760 355340 158432
rect 492680 157760 510472 158432
rect 19968 157040 22028 157388
rect 195756 157040 197816 157388
rect 195076 156360 197096 156708
rect 808 155040 20328 155712
rect 105796 155040 111988 155712
rect 197456 155040 209648 155712
rect 348428 155040 354620 155712
rect 493400 155040 512920 155712
rect 18816 153824 21048 154496
rect 105076 153824 107308 154496
rect 110476 153824 112708 154496
rect 196736 153824 198968 154496
rect 3256 146880 21048 147552
rect 105076 146880 112708 147552
rect 196736 146880 210368 147552
rect 347708 146880 355340 147552
rect 492680 146880 510472 147552
rect 808 144160 20328 144832
rect 105796 144160 111988 144832
rect 197456 144160 209648 144832
rect 348428 144160 354620 144832
rect 493400 144160 512920 144832
rect 3256 136000 21048 136672
rect 105076 136000 112708 136672
rect 196736 136000 210368 136672
rect 347708 136000 355340 136672
rect 492680 136000 510472 136672
rect 808 133280 20328 133952
rect 105796 133280 111988 133952
rect 197456 133280 209648 133952
rect 348428 133280 354620 133952
rect 493400 133280 512920 133952
rect 3256 125120 21048 125792
rect 105076 125120 112708 125792
rect 196736 125120 210368 125792
rect 347708 125120 355340 125792
rect 492680 125120 510472 125792
rect 808 122400 20328 123072
rect 105796 122400 111988 123072
rect 197456 122400 209648 123072
rect 348428 122400 354620 123072
rect 493400 122400 512920 123072
rect 3256 114240 21048 114912
rect 105076 114240 112708 114912
rect 196736 114240 210368 114912
rect 347708 114240 355340 114912
rect 492680 114240 510472 114912
rect 346728 112972 348788 113320
rect 808 111520 20328 112192
rect 105796 111520 111988 112192
rect 197456 111620 209648 112192
rect 210008 111980 348068 112340
rect 348428 111620 354620 112192
rect 354980 111980 493040 112340
rect 493400 111620 512920 112192
rect 197456 111520 512920 111620
rect 209288 111260 348788 111520
rect 353600 111260 493760 111520
rect 209288 105428 348788 105788
rect 353600 105428 493760 105788
rect 210008 104708 348068 105068
rect 354980 104708 493040 105068
rect 3256 103360 21048 104032
rect 105076 103360 112708 104032
rect 196736 103360 210368 104032
rect 346048 103048 346396 104708
rect 347708 103360 355340 104032
rect 356652 103048 357000 104708
rect 492680 103360 510472 104032
rect 808 100640 20328 101312
rect 105796 100640 111988 101312
rect 197456 100640 209648 101312
rect 348428 100640 354620 101312
rect 493400 100640 512920 101312
rect 3256 92480 21048 93152
rect 105076 92480 112708 93152
rect 196736 92480 210368 93152
rect 347708 92480 355340 93152
rect 492680 92480 510472 93152
rect 808 89760 20328 90432
rect 105796 89760 111988 90432
rect 197456 89760 209648 90432
rect 348428 89760 354620 90432
rect 493400 89760 512920 90432
rect 3256 81600 21048 82272
rect 105076 81600 112708 82272
rect 196736 81600 210368 82272
rect 347708 81600 355340 82272
rect 492680 81600 510472 82272
rect 808 78880 20328 79552
rect 105796 78880 111988 79552
rect 197456 78880 209648 79552
rect 348428 78880 354620 79552
rect 493400 78880 512920 79552
rect 3256 70720 21048 71392
rect 105076 70720 112708 71392
rect 196736 70720 210368 71392
rect 347708 70720 355340 71392
rect 492680 70720 510472 71392
rect 808 68000 20328 68672
rect 105796 68000 111988 68672
rect 197456 68000 209648 68672
rect 348428 68000 354620 68672
rect 493400 68000 512920 68672
rect 3256 59840 21048 60512
rect 105076 59840 112708 60512
rect 196736 59840 210368 60512
rect 347708 59840 355340 60512
rect 492680 59840 510472 60512
rect 808 57120 20328 57792
rect 105796 57120 111988 57792
rect 197456 57120 209648 57792
rect 348428 57120 354620 57792
rect 493400 57120 512920 57792
rect 3256 48960 21048 49632
rect 105076 48960 112708 49632
rect 196736 48960 210368 49632
rect 347708 48960 355340 49632
rect 492680 48960 510472 49632
rect 808 46240 20328 46912
rect 105796 46240 111988 46912
rect 197456 46240 209648 46912
rect 348428 46240 354620 46912
rect 493400 46240 512920 46912
rect 3256 38080 21048 38752
rect 105076 38080 112708 38752
rect 196736 38080 210368 38752
rect 347708 38080 355340 38752
rect 492680 38080 510472 38752
rect 808 35360 20328 36032
rect 105796 35360 111988 36032
rect 197456 35360 209648 36032
rect 348428 35360 354620 36032
rect 493400 35360 512920 36032
rect 3256 27200 21048 27872
rect 105076 27200 112708 27872
rect 196736 27200 210368 27872
rect 347708 27200 355340 27872
rect 492680 27200 510472 27872
rect 808 24480 20328 25152
rect 105796 24480 111988 25152
rect 197456 24480 209648 25152
rect 348428 24480 354620 25152
rect 493400 24480 512920 25152
rect 20688 21992 22708 22340
rect 346728 21312 348788 21660
rect 491700 21312 493760 21660
rect 20688 20320 105436 20680
rect 112348 20320 197096 20680
rect 210008 20320 348068 20680
rect 354980 20320 493040 20680
rect 19968 19600 106156 19960
rect 111628 19600 197816 19960
rect 209288 19600 348788 19960
rect 353600 19600 493760 19960
rect 3256 16320 510472 16992
rect 808 13600 512920 14272
rect 3256 5440 510472 6112
rect 0 3264 513728 4896
rect 0 816 513728 2448
<< obsm5 >>
rect 0 512176 513728 512992
rect 0 509728 513728 510544
rect 0 506592 513728 508096
rect 0 505920 3256 506592
rect 510472 505920 513728 506592
rect 0 503872 513728 505920
rect 0 503200 808 503872
rect 512920 503200 513728 503872
rect 0 495712 513728 503200
rect 0 495040 3256 495712
rect 510472 495040 513728 495712
rect 0 493392 513728 495040
rect 0 493032 19968 493392
rect 159468 493032 164940 493392
rect 304440 493032 315912 493392
rect 402100 493032 407572 493392
rect 493760 493032 513728 493392
rect 0 492992 513728 493032
rect 0 492320 808 492992
rect 16992 492672 310077 492992
rect 16992 492320 20688 492672
rect 0 492312 20688 492320
rect 158748 492312 165660 492672
rect 303720 492320 310077 492672
rect 310752 492672 495040 492992
rect 310752 492320 316632 492672
rect 303720 492312 316632 492320
rect 401380 492312 408292 492672
rect 493040 492320 495040 492672
rect 512920 492320 513728 492992
rect 493040 492312 513728 492320
rect 0 491680 167332 492312
rect 0 491332 19968 491680
rect 22028 491332 167332 491680
rect 0 491000 167332 491332
rect 0 490652 20688 491000
rect 22708 490652 167332 491000
rect 167680 491680 513728 492312
rect 167680 491332 302380 491680
rect 304440 491332 400040 491680
rect 402100 491332 513728 491680
rect 167680 491000 513728 491332
rect 167680 490652 491020 491000
rect 493040 490652 513728 491000
rect 0 484832 513728 490652
rect 0 484160 3256 484832
rect 21048 484160 158388 484832
rect 166020 484160 303360 484832
rect 316992 484160 401020 484832
rect 408652 484160 492680 484832
rect 510472 484160 513728 484832
rect 0 482112 513728 484160
rect 0 481440 808 482112
rect 20328 481440 159108 482112
rect 165300 481440 304080 482112
rect 316272 481440 401740 482112
rect 407932 481440 493400 482112
rect 512920 481440 513728 482112
rect 0 473952 513728 481440
rect 0 473280 3256 473952
rect 21048 473280 158388 473952
rect 166020 473280 303360 473952
rect 316992 473280 401020 473952
rect 408652 473280 492680 473952
rect 510472 473280 513728 473952
rect 0 471232 513728 473280
rect 0 470560 808 471232
rect 20328 470560 159108 471232
rect 165300 470560 304080 471232
rect 316272 470560 401740 471232
rect 407932 470560 493400 471232
rect 512920 470560 513728 471232
rect 0 463072 513728 470560
rect 0 462400 3256 463072
rect 21048 462400 158388 463072
rect 166020 462400 303360 463072
rect 316992 462400 401020 463072
rect 408652 462400 492680 463072
rect 510472 462400 513728 463072
rect 0 460352 513728 462400
rect 0 459680 808 460352
rect 20328 459680 159108 460352
rect 165300 459680 304080 460352
rect 316272 459680 401740 460352
rect 407932 459680 493400 460352
rect 512920 459680 513728 460352
rect 0 452192 513728 459680
rect 0 451520 3256 452192
rect 21048 451520 158388 452192
rect 166020 451520 303360 452192
rect 316992 451520 401020 452192
rect 408652 451520 492680 452192
rect 510472 451520 513728 452192
rect 0 449472 513728 451520
rect 0 448800 808 449472
rect 20328 448800 159108 449472
rect 165300 448800 304080 449472
rect 316272 448800 401740 449472
rect 407932 448800 493400 449472
rect 512920 448800 513728 449472
rect 0 441312 513728 448800
rect 0 440640 3256 441312
rect 21048 440640 158388 441312
rect 166020 440640 303360 441312
rect 316992 440640 401020 441312
rect 408652 440640 492680 441312
rect 510472 440640 513728 441312
rect 0 438592 513728 440640
rect 0 437920 808 438592
rect 20328 437920 159108 438592
rect 165300 437920 304080 438592
rect 316272 437920 401740 438592
rect 407932 437920 493400 438592
rect 512920 437920 513728 438592
rect 0 430432 513728 437920
rect 0 429760 3256 430432
rect 21048 429760 158388 430432
rect 166020 429760 303360 430432
rect 316992 429760 401020 430432
rect 408652 429760 492680 430432
rect 510472 429760 513728 430432
rect 0 427712 513728 429760
rect 0 427040 808 427712
rect 20328 427040 159108 427712
rect 165300 427040 304080 427712
rect 316272 427040 401740 427712
rect 407932 427040 493400 427712
rect 512920 427040 513728 427712
rect 0 419552 513728 427040
rect 0 418880 3256 419552
rect 21048 418880 158388 419552
rect 166020 418880 303360 419552
rect 316992 418880 401020 419552
rect 408652 418880 492680 419552
rect 510472 418880 513728 419552
rect 0 416832 513728 418880
rect 0 416160 808 416832
rect 20328 416160 159108 416832
rect 165300 416160 304080 416832
rect 316272 416160 401740 416832
rect 407932 416160 493400 416832
rect 512920 416160 513728 416832
rect 0 408672 513728 416160
rect 0 408000 3256 408672
rect 21048 408284 158388 408672
rect 166020 408284 303360 408672
rect 316992 408000 401020 408672
rect 408652 408000 492680 408672
rect 510472 408000 513728 408672
rect 0 407924 20688 408000
rect 158748 407924 165660 408000
rect 303720 407924 513728 408000
rect 0 407564 513728 407924
rect 0 407204 19968 407564
rect 159468 407204 164940 407564
rect 304440 407204 513728 407564
rect 0 405952 513728 407204
rect 0 405280 808 405952
rect 316272 405280 401740 405952
rect 407932 405280 493400 405952
rect 512920 405280 513728 405952
rect 0 401732 513728 405280
rect 0 401372 19968 401732
rect 159468 401372 164940 401732
rect 304440 401372 513728 401732
rect 0 401012 513728 401372
rect 0 400652 20688 401012
rect 158748 400652 165660 401012
rect 303720 400652 513728 401012
rect 0 400020 301700 400652
rect 0 399672 19968 400020
rect 22028 399672 164940 400020
rect 167000 399672 301700 400020
rect 0 399340 301700 399672
rect 0 398992 20688 399340
rect 22708 398992 301700 399340
rect 302048 398992 513728 400652
rect 0 397792 513728 398992
rect 0 397120 3256 397792
rect 21048 397120 158388 397792
rect 166020 397120 303360 397792
rect 316992 397120 401020 397792
rect 408652 397120 492680 397792
rect 510472 397120 513728 397792
rect 0 395072 513728 397120
rect 0 394400 808 395072
rect 20328 394400 159108 395072
rect 165300 394400 304080 395072
rect 316272 394400 401740 395072
rect 407932 394400 493400 395072
rect 512920 394400 513728 395072
rect 0 386912 513728 394400
rect 0 386240 3256 386912
rect 21048 386240 158388 386912
rect 166020 386240 303360 386912
rect 316992 386240 401020 386912
rect 408652 386240 492680 386912
rect 510472 386240 513728 386912
rect 0 384192 513728 386240
rect 0 383520 808 384192
rect 20328 383520 159108 384192
rect 165300 383520 304080 384192
rect 316272 383520 401740 384192
rect 407932 383520 493400 384192
rect 512920 383520 513728 384192
rect 0 376032 513728 383520
rect 0 375360 3256 376032
rect 21048 375360 158388 376032
rect 166020 375360 303360 376032
rect 316992 375360 401020 376032
rect 408652 375360 492680 376032
rect 510472 375360 513728 376032
rect 0 373312 513728 375360
rect 0 372640 808 373312
rect 20328 372640 159108 373312
rect 165300 372640 304080 373312
rect 316272 372640 401740 373312
rect 407932 372640 493400 373312
rect 512920 372640 513728 373312
rect 0 365152 513728 372640
rect 0 364480 3256 365152
rect 21048 364480 158388 365152
rect 166020 364480 303360 365152
rect 316992 364480 401020 365152
rect 408652 364480 492680 365152
rect 510472 364480 513728 365152
rect 0 362432 513728 364480
rect 0 361760 808 362432
rect 20328 361760 159108 362432
rect 165300 361760 304080 362432
rect 316272 361760 401740 362432
rect 407932 361760 493400 362432
rect 512920 361760 513728 362432
rect 0 356632 513728 361760
rect 0 356284 316632 356632
rect 318652 356284 513728 356632
rect 0 355952 513728 356284
rect 0 355604 491700 355952
rect 493760 355604 513728 355952
rect 0 354972 513728 355604
rect 0 354612 316632 354972
rect 401380 354612 408292 354972
rect 493040 354612 513728 354972
rect 0 354272 513728 354612
rect 0 353600 3256 354272
rect 21048 353600 158388 354272
rect 166020 353600 303360 354272
rect 313472 354252 497760 354272
rect 313472 353892 315912 354252
rect 402100 353892 407572 354252
rect 493760 353892 497760 354252
rect 313472 353600 497760 353892
rect 510472 353600 513728 354272
rect 0 351552 513728 353600
rect 0 350880 808 351552
rect 20328 350880 159108 351552
rect 165300 350880 304080 351552
rect 512920 350880 513728 351552
rect 0 348420 513728 350880
rect 0 348060 315912 348420
rect 402100 348060 407572 348420
rect 493760 348060 513728 348420
rect 0 347700 513728 348060
rect 0 347340 316632 347700
rect 401380 347340 408292 347700
rect 493040 347340 513728 347700
rect 0 343392 513728 347340
rect 0 342720 3256 343392
rect 21048 342720 158388 343392
rect 166020 342720 303360 343392
rect 316992 342720 401020 343392
rect 408652 342720 492680 343392
rect 510472 342720 513728 343392
rect 0 340672 513728 342720
rect 0 340000 808 340672
rect 20328 340000 159108 340672
rect 165300 340000 304080 340672
rect 316272 340000 401740 340672
rect 407932 340000 493400 340672
rect 512920 340000 513728 340672
rect 0 332512 513728 340000
rect 0 331840 3256 332512
rect 21048 331840 158388 332512
rect 166020 331840 303360 332512
rect 316992 331840 401020 332512
rect 408652 331840 492680 332512
rect 510472 331840 513728 332512
rect 0 329792 513728 331840
rect 0 329120 808 329792
rect 20328 329120 159108 329792
rect 165300 329120 304080 329792
rect 316272 329120 401740 329792
rect 407932 329120 493400 329792
rect 512920 329120 513728 329792
rect 0 321632 513728 329120
rect 0 320960 3256 321632
rect 21048 320960 158388 321632
rect 166020 320960 303360 321632
rect 316992 320960 401020 321632
rect 408652 320960 492680 321632
rect 510472 320960 513728 321632
rect 0 318912 513728 320960
rect 0 318240 808 318912
rect 20328 318240 159108 318912
rect 165300 318240 304080 318912
rect 316272 318240 401740 318912
rect 407932 318240 493400 318912
rect 512920 318240 513728 318912
rect 0 316624 513728 318240
rect 0 316264 20688 316624
rect 158748 316264 165660 316624
rect 303720 316264 513728 316624
rect 0 315904 513728 316264
rect 0 315544 19968 315904
rect 159468 315544 164940 315904
rect 304440 315544 513728 315904
rect 0 310752 513728 315544
rect 0 310080 3256 310752
rect 316992 310080 401020 310752
rect 408652 310080 492680 310752
rect 510472 310080 513728 310752
rect 0 308032 513728 310080
rect 0 307360 808 308032
rect 316272 307360 401740 308032
rect 407932 307360 493400 308032
rect 512920 307360 513728 308032
rect 0 304072 513728 307360
rect 0 303712 19968 304072
rect 106156 303712 111628 304072
rect 197816 303712 513728 304072
rect 0 303352 513728 303712
rect 0 302992 20688 303352
rect 105436 302992 112348 303352
rect 197096 302992 513728 303352
rect 0 302360 513728 302992
rect 0 302012 19968 302360
rect 22028 302012 195756 302360
rect 197816 302012 513728 302360
rect 0 299872 513728 302012
rect 0 299200 3256 299872
rect 21048 299200 105076 299872
rect 112708 299200 196736 299872
rect 316992 299200 401020 299872
rect 408652 299200 492680 299872
rect 510472 299200 513728 299872
rect 0 297152 513728 299200
rect 0 296480 808 297152
rect 20328 296480 105796 297152
rect 111988 296480 197456 297152
rect 316272 296480 401740 297152
rect 407932 296480 493400 297152
rect 512920 296480 513728 297152
rect 0 288992 513728 296480
rect 0 288320 3256 288992
rect 21048 288320 105076 288992
rect 112708 288320 196736 288992
rect 316992 288320 401020 288992
rect 408652 288320 492680 288992
rect 510472 288320 513728 288992
rect 0 286272 513728 288320
rect 0 285600 808 286272
rect 20328 285600 105796 286272
rect 111988 285600 197456 286272
rect 316272 285600 401740 286272
rect 407932 285600 493400 286272
rect 512920 285600 513728 286272
rect 0 278112 513728 285600
rect 0 277440 3256 278112
rect 21048 277440 105076 278112
rect 112708 277440 196736 278112
rect 316992 277440 401020 278112
rect 408652 277440 492680 278112
rect 510472 277440 513728 278112
rect 0 275392 513728 277440
rect 0 274720 808 275392
rect 20328 274720 105796 275392
rect 111988 274720 197456 275392
rect 316272 274720 401740 275392
rect 407932 274720 493400 275392
rect 512920 274720 513728 275392
rect 0 267232 513728 274720
rect 0 266560 3256 267232
rect 21048 266560 105076 267232
rect 112708 266560 196736 267232
rect 316992 266560 401020 267232
rect 408652 266560 492680 267232
rect 510472 266560 513728 267232
rect 0 264512 513728 266560
rect 0 263840 808 264512
rect 20328 263840 105796 264512
rect 111988 263840 197456 264512
rect 316272 263840 401740 264512
rect 407932 263840 493400 264512
rect 512920 263840 513728 264512
rect 0 256352 513728 263840
rect 0 255680 3256 256352
rect 21048 255680 105076 256352
rect 112708 255680 196736 256352
rect 316992 255680 401020 256352
rect 408652 255680 492680 256352
rect 510472 255680 513728 256352
rect 0 253632 513728 255680
rect 0 252960 808 253632
rect 20328 252960 105796 253632
rect 111988 252960 197456 253632
rect 316272 252960 401740 253632
rect 407932 252960 493400 253632
rect 512920 252960 513728 253632
rect 0 245472 513728 252960
rect 0 244800 3256 245472
rect 21048 244800 105076 245472
rect 112708 244800 196736 245472
rect 316992 244800 401020 245472
rect 408652 244800 492680 245472
rect 510472 244800 513728 245472
rect 0 242752 513728 244800
rect 0 242080 808 242752
rect 20328 242080 105796 242752
rect 111988 242080 197456 242752
rect 316272 242080 401740 242752
rect 407932 242080 493400 242752
rect 512920 242080 513728 242752
rect 0 234592 513728 242080
rect 0 233920 3256 234592
rect 21048 233920 105076 234592
rect 112708 233920 196736 234592
rect 316992 233920 401020 234592
rect 408652 233920 492680 234592
rect 510472 233920 513728 234592
rect 0 231872 513728 233920
rect 0 231200 808 231872
rect 20328 231200 105796 231872
rect 111988 231200 197456 231872
rect 316272 231200 401740 231872
rect 407932 231200 493400 231872
rect 512920 231200 513728 231872
rect 0 223712 513728 231200
rect 0 223040 3256 223712
rect 21048 223040 105076 223712
rect 112708 223040 196736 223712
rect 316992 223040 401020 223712
rect 408652 223040 492680 223712
rect 510472 223040 513728 223712
rect 0 220992 513728 223040
rect 0 220320 808 220992
rect 20328 220320 105796 220992
rect 111988 220320 197456 220992
rect 316272 220320 401740 220992
rect 407932 220320 493400 220992
rect 512920 220320 513728 220992
rect 0 212832 513728 220320
rect 0 212160 3256 212832
rect 21048 212160 105076 212832
rect 112708 212160 196736 212832
rect 316992 212160 401020 212832
rect 408652 212160 492680 212832
rect 510472 212160 513728 212832
rect 0 211660 513728 212160
rect 0 211312 316632 211660
rect 318652 211312 491020 211660
rect 493040 211312 513728 211660
rect 0 210980 513728 211312
rect 0 210632 400040 210980
rect 402100 210632 491700 210980
rect 493760 210632 513728 210980
rect 0 210112 513728 210632
rect 0 209440 808 210112
rect 20328 209440 105796 210112
rect 111988 209440 197456 210112
rect 310753 210000 495040 210112
rect 310753 209640 316632 210000
rect 401380 209640 408292 210000
rect 493040 209640 495040 210000
rect 310753 209440 495040 209640
rect 512920 209440 513728 210112
rect 0 209280 513728 209440
rect 0 208920 315912 209280
rect 402100 208920 407572 209280
rect 493760 208920 513728 209280
rect 0 201952 513728 208920
rect 0 201280 3256 201952
rect 21048 201280 105076 201952
rect 112708 201280 196736 201952
rect 510472 201280 513728 201952
rect 0 199232 513728 201280
rect 0 198560 808 199232
rect 20328 198560 105796 199232
rect 111988 198560 197456 199232
rect 512920 198560 513728 199232
rect 0 197448 513728 198560
rect 0 197088 209288 197448
rect 348788 197088 353600 197448
rect 493760 197088 513728 197448
rect 0 196728 513728 197088
rect 0 196368 210008 196728
rect 348068 196368 354980 196728
rect 493040 196368 513728 196728
rect 0 194708 346048 196368
rect 346396 194708 356652 196368
rect 357000 195736 513728 196368
rect 357000 195388 491700 195736
rect 493760 195388 513728 195736
rect 357000 194708 513728 195388
rect 0 191072 513728 194708
rect 0 190400 3256 191072
rect 21048 190400 105076 191072
rect 112708 190400 196736 191072
rect 210368 190400 347708 191072
rect 355340 190400 492680 191072
rect 510472 190400 513728 191072
rect 0 188352 513728 190400
rect 0 187680 808 188352
rect 20328 187680 105796 188352
rect 111988 187680 197456 188352
rect 209648 187680 348428 188352
rect 354620 187680 493400 188352
rect 512920 187680 513728 188352
rect 0 180192 513728 187680
rect 0 179520 3256 180192
rect 21048 179520 105076 180192
rect 112708 179520 196736 180192
rect 210368 179520 347708 180192
rect 355340 179520 492680 180192
rect 510472 179520 513728 180192
rect 0 177472 513728 179520
rect 0 176800 808 177472
rect 20328 176800 105796 177472
rect 111988 176800 197456 177472
rect 209648 176800 348428 177472
rect 354620 176800 493400 177472
rect 512920 176800 513728 177472
rect 0 169312 513728 176800
rect 0 168640 3256 169312
rect 21048 168640 105076 169312
rect 112708 168640 196736 169312
rect 210368 168640 347708 169312
rect 355340 168640 492680 169312
rect 510472 168640 513728 169312
rect 0 167312 513728 168640
rect 0 166964 20688 167312
rect 22708 166964 195076 167312
rect 197096 166964 513728 167312
rect 0 166592 513728 166964
rect 0 165920 808 166592
rect 20328 165920 105796 166592
rect 111988 165920 197456 166592
rect 209648 165920 348428 166592
rect 354620 165920 493400 166592
rect 512920 165920 513728 166592
rect 0 165652 513728 165920
rect 0 165292 20688 165652
rect 105436 165292 112348 165652
rect 197096 165292 513728 165652
rect 0 164932 513728 165292
rect 0 164572 19968 164932
rect 106156 164572 111628 164932
rect 197816 164572 513728 164932
rect 0 159100 513728 164572
rect 0 158740 19968 159100
rect 106156 158740 111628 159100
rect 197816 158740 513728 159100
rect 0 158432 513728 158740
rect 0 157760 3256 158432
rect 19488 158380 106636 158432
rect 19488 158020 20688 158380
rect 105436 158020 106636 158380
rect 19488 157760 106636 158020
rect 111148 158380 198296 158432
rect 111148 158020 112348 158380
rect 197096 158020 198296 158380
rect 111148 157760 198296 158020
rect 210368 157760 347708 158432
rect 355340 157760 492680 158432
rect 510472 157760 513728 158432
rect 0 157388 513728 157760
rect 0 157040 19968 157388
rect 22028 157040 195756 157388
rect 197816 157040 513728 157388
rect 0 156708 513728 157040
rect 0 156360 195076 156708
rect 197096 156360 513728 156708
rect 0 155712 513728 156360
rect 0 155040 808 155712
rect 20328 155040 105796 155712
rect 111988 155040 197456 155712
rect 209648 155040 348428 155712
rect 354620 155040 493400 155712
rect 512920 155040 513728 155712
rect 0 154496 513728 155040
rect 0 153824 18816 154496
rect 21048 153824 105076 154496
rect 107308 153824 110476 154496
rect 112708 153824 196736 154496
rect 198968 153824 513728 154496
rect 0 147552 513728 153824
rect 0 146880 3256 147552
rect 21048 146880 105076 147552
rect 112708 146880 196736 147552
rect 210368 146880 347708 147552
rect 355340 146880 492680 147552
rect 510472 146880 513728 147552
rect 0 144832 513728 146880
rect 0 144160 808 144832
rect 20328 144160 105796 144832
rect 111988 144160 197456 144832
rect 209648 144160 348428 144832
rect 354620 144160 493400 144832
rect 512920 144160 513728 144832
rect 0 136672 513728 144160
rect 0 136000 3256 136672
rect 21048 136000 105076 136672
rect 112708 136000 196736 136672
rect 210368 136000 347708 136672
rect 355340 136000 492680 136672
rect 510472 136000 513728 136672
rect 0 133952 513728 136000
rect 0 133280 808 133952
rect 20328 133280 105796 133952
rect 111988 133280 197456 133952
rect 209648 133280 348428 133952
rect 354620 133280 493400 133952
rect 512920 133280 513728 133952
rect 0 125792 513728 133280
rect 0 125120 3256 125792
rect 21048 125120 105076 125792
rect 112708 125120 196736 125792
rect 210368 125120 347708 125792
rect 355340 125120 492680 125792
rect 510472 125120 513728 125792
rect 0 123072 513728 125120
rect 0 122400 808 123072
rect 20328 122400 105796 123072
rect 111988 122400 197456 123072
rect 209648 122400 348428 123072
rect 354620 122400 493400 123072
rect 512920 122400 513728 123072
rect 0 114912 513728 122400
rect 0 114240 3256 114912
rect 21048 114240 105076 114912
rect 112708 114240 196736 114912
rect 210368 114240 347708 114912
rect 355340 114240 492680 114912
rect 510472 114240 513728 114912
rect 0 113320 513728 114240
rect 0 112972 346728 113320
rect 348788 112972 513728 113320
rect 0 112340 513728 112972
rect 0 112192 210008 112340
rect 0 111520 808 112192
rect 20328 111520 105796 112192
rect 111988 111520 197456 112192
rect 209648 111980 210008 112192
rect 348068 112192 354980 112340
rect 348068 111980 348428 112192
rect 209648 111620 348428 111980
rect 354620 111980 354980 112192
rect 493040 112192 513728 112340
rect 493040 111980 493400 112192
rect 354620 111620 493400 111980
rect 512920 111520 513728 112192
rect 0 111260 209288 111520
rect 348788 111260 353600 111520
rect 493760 111260 513728 111520
rect 0 105788 513728 111260
rect 0 105428 209288 105788
rect 348788 105428 353600 105788
rect 493760 105428 513728 105788
rect 0 105068 513728 105428
rect 0 104708 210008 105068
rect 348068 104708 354980 105068
rect 493040 104708 513728 105068
rect 0 104032 346048 104708
rect 0 103360 3256 104032
rect 21048 103360 105076 104032
rect 112708 103360 196736 104032
rect 210368 103360 346048 104032
rect 0 103048 346048 103360
rect 346396 104032 356652 104708
rect 346396 103360 347708 104032
rect 355340 103360 356652 104032
rect 346396 103048 356652 103360
rect 357000 104032 513728 104708
rect 357000 103360 492680 104032
rect 510472 103360 513728 104032
rect 357000 103048 513728 103360
rect 0 101312 513728 103048
rect 0 100640 808 101312
rect 20328 100640 105796 101312
rect 111988 100640 197456 101312
rect 209648 100640 348428 101312
rect 354620 100640 493400 101312
rect 512920 100640 513728 101312
rect 0 93152 513728 100640
rect 0 92480 3256 93152
rect 21048 92480 105076 93152
rect 112708 92480 196736 93152
rect 210368 92480 347708 93152
rect 355340 92480 492680 93152
rect 510472 92480 513728 93152
rect 0 90432 513728 92480
rect 0 89760 808 90432
rect 20328 89760 105796 90432
rect 111988 89760 197456 90432
rect 209648 89760 348428 90432
rect 354620 89760 493400 90432
rect 512920 89760 513728 90432
rect 0 82272 513728 89760
rect 0 81600 3256 82272
rect 21048 81600 105076 82272
rect 112708 81600 196736 82272
rect 210368 81600 347708 82272
rect 355340 81600 492680 82272
rect 510472 81600 513728 82272
rect 0 79552 513728 81600
rect 0 78880 808 79552
rect 20328 78880 105796 79552
rect 111988 78880 197456 79552
rect 209648 78880 348428 79552
rect 354620 78880 493400 79552
rect 512920 78880 513728 79552
rect 0 71392 513728 78880
rect 0 70720 3256 71392
rect 21048 70720 105076 71392
rect 112708 70720 196736 71392
rect 210368 70720 347708 71392
rect 355340 70720 492680 71392
rect 510472 70720 513728 71392
rect 0 68672 513728 70720
rect 0 68000 808 68672
rect 20328 68000 105796 68672
rect 111988 68000 197456 68672
rect 209648 68000 348428 68672
rect 354620 68000 493400 68672
rect 512920 68000 513728 68672
rect 0 60512 513728 68000
rect 0 59840 3256 60512
rect 21048 59840 105076 60512
rect 112708 59840 196736 60512
rect 210368 59840 347708 60512
rect 355340 59840 492680 60512
rect 510472 59840 513728 60512
rect 0 57792 513728 59840
rect 0 57120 808 57792
rect 20328 57120 105796 57792
rect 111988 57120 197456 57792
rect 209648 57120 348428 57792
rect 354620 57120 493400 57792
rect 512920 57120 513728 57792
rect 0 49632 513728 57120
rect 0 48960 3256 49632
rect 21048 48960 105076 49632
rect 112708 48960 196736 49632
rect 210368 48960 347708 49632
rect 355340 48960 492680 49632
rect 510472 48960 513728 49632
rect 0 46912 513728 48960
rect 0 46240 808 46912
rect 20328 46240 105796 46912
rect 111988 46240 197456 46912
rect 209648 46240 348428 46912
rect 354620 46240 493400 46912
rect 512920 46240 513728 46912
rect 0 38752 513728 46240
rect 0 38080 3256 38752
rect 21048 38080 105076 38752
rect 112708 38080 196736 38752
rect 210368 38080 347708 38752
rect 355340 38080 492680 38752
rect 510472 38080 513728 38752
rect 0 36032 513728 38080
rect 0 35360 808 36032
rect 20328 35360 105796 36032
rect 111988 35360 197456 36032
rect 209648 35360 348428 36032
rect 354620 35360 493400 36032
rect 512920 35360 513728 36032
rect 0 27872 513728 35360
rect 0 27200 3256 27872
rect 21048 27200 105076 27872
rect 112708 27200 196736 27872
rect 210368 27200 347708 27872
rect 355340 27200 492680 27872
rect 510472 27200 513728 27872
rect 0 25152 513728 27200
rect 0 24480 808 25152
rect 20328 24480 105796 25152
rect 111988 24480 197456 25152
rect 209648 24480 348428 25152
rect 354620 24480 493400 25152
rect 512920 24480 513728 25152
rect 0 22340 513728 24480
rect 0 21992 20688 22340
rect 22708 21992 513728 22340
rect 0 21660 513728 21992
rect 0 21312 346728 21660
rect 348788 21312 491700 21660
rect 493760 21312 513728 21660
rect 0 20680 513728 21312
rect 0 20320 20688 20680
rect 105436 20320 112348 20680
rect 197096 20320 210008 20680
rect 348068 20320 354980 20680
rect 493040 20320 513728 20680
rect 0 19960 513728 20320
rect 0 19600 19968 19960
rect 106156 19600 111628 19960
rect 197816 19600 209288 19960
rect 348788 19600 353600 19960
rect 493760 19600 513728 19960
rect 0 16992 513728 19600
rect 0 16320 3256 16992
rect 510472 16320 513728 16992
rect 0 14272 513728 16320
rect 0 13600 808 14272
rect 512920 13600 513728 14272
rect 0 6112 513728 13600
rect 0 5440 3256 6112
rect 510472 5440 513728 6112
rect 0 4896 513728 5440
rect 0 2448 513728 3264
rect 0 0 513728 816
<< labels >>
rlabel metal2 s 216 512895 244 512992 6 clk
port 1 nsew signal input
rlabel metal2 s 73356 512895 73384 512992 6 rst_n
port 2 nsew signal input
rlabel metal2 s 146772 512895 146800 512992 6 load_en
port 3 nsew signal input
rlabel metal2 s 220096 512895 220124 512992 6 debug_en
port 4 nsew signal input
rlabel metal2 s 366836 512895 366864 512992 6 serial_in
port 5 nsew signal input
rlabel metal2 s 513484 512895 513512 512992 6 sram_select[1]
port 6 nsew signal input
rlabel metal2 s 440252 512895 440280 512992 6 sram_select[0]
port 7 nsew signal input
rlabel metal2 s 0 512944 97 512972 6 frequency_adc_done
port 8 nsew signal input
rlabel metal2 s 0 241352 97 241380 6 amplitude_adc_done
port 9 nsew signal input
rlabel metal2 s 0 271544 97 271572 6 sig_frequency[7]
port 10 nsew signal input
rlabel metal2 s 0 301736 97 301764 6 sig_frequency[6]
port 11 nsew signal input
rlabel metal2 s 0 331860 97 331888 6 sig_frequency[5]
port 12 nsew signal input
rlabel metal2 s 0 362052 97 362080 6 sig_frequency[4]
port 13 nsew signal input
rlabel metal2 s 0 392244 97 392272 6 sig_frequency[3]
port 14 nsew signal input
rlabel metal2 s 0 422368 97 422396 6 sig_frequency[2]
port 15 nsew signal input
rlabel metal2 s 0 452560 97 452588 6 sig_frequency[1]
port 16 nsew signal input
rlabel metal2 s 0 482752 97 482780 6 sig_frequency[0]
port 17 nsew signal input
rlabel metal2 s 0 20 97 48 6 sig_amplitude[7]
port 18 nsew signal input
rlabel metal2 s 0 30144 97 30172 6 sig_amplitude[6]
port 19 nsew signal input
rlabel metal2 s 0 60336 97 60364 6 sig_amplitude[5]
port 20 nsew signal input
rlabel metal2 s 0 90528 97 90556 6 sig_amplitude[4]
port 21 nsew signal input
rlabel metal2 s 0 120652 97 120680 6 sig_amplitude[3]
port 22 nsew signal input
rlabel metal2 s 0 150844 97 150872 6 sig_amplitude[2]
port 23 nsew signal input
rlabel metal2 s 0 181036 97 181064 6 sig_amplitude[1]
port 24 nsew signal input
rlabel metal2 s 0 211160 97 211188 6 sig_amplitude[0]
port 25 nsew signal input
rlabel metal2 s 293512 512895 293540 512992 6 adc_bypass_en
port 26 nsew signal input
rlabel metal2 s 513631 512944 513728 512972 6 serial_out
port 27 nsew signal output
rlabel metal2 s 513631 256516 513728 256544 6 serial_out_valid
port 28 nsew signal output
rlabel metal2 s 513631 20 513728 48 6 freq_eval_done
port 29 nsew signal output
rlabel metal5 s 512096 510544 513728 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 0 510544 1632 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 512096 816 513728 2448 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 0 816 1632 2448 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 511288 511360 512920 512992 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 511288 0 512920 1632 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 808 511360 2440 512992 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 808 0 2440 1632 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 495040 492320 495712 492992 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 400040 491332 400388 491680 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 310080 492320 310752 492992 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 302380 491332 302728 491680 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 491700 355604 492048 355952 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 166652 399672 167000 400020 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 21680 491332 22028 491680 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 16320 492320 16992 492992 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 21680 399672 22028 400020 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 195756 302012 196104 302360 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 21680 302012 22028 302360 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 491700 210632 492048 210980 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 491700 195388 492048 195736 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 400040 210632 400388 210980 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 353600 197088 354620 197448 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 111260 493760 112192 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 491700 21312 492048 21660 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 353600 105428 354620 105788 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 353600 111260 354620 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 346728 112972 347076 113320 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 348428 111260 348788 112192 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 353600 19600 354620 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 346728 21312 347076 21660 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 195756 157040 196104 157388 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 21680 157040 22028 157388 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 209288 111260 209648 112192 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 495041 492320 512920 492992 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 481440 512920 482112 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 470560 512920 471232 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 459680 512920 460352 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 481440 407932 482112 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 400214 491332 402100 491680 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 470560 407932 471232 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 459680 407932 460352 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 407572 493032 493760 493392 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 437920 512920 438592 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 427040 512920 427712 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 416160 512920 416832 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 405280 512920 405952 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 394400 512920 395072 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 437920 407932 438592 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 427040 407932 427712 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 416160 407932 416832 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 405280 407932 405952 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 394400 407932 395072 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 448800 512920 449472 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 448800 407932 449472 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 310077 492320 310749 492992 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 302514 491332 304440 491680 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 304080 481440 316272 482112 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 304080 470560 316272 471232 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 304080 459680 316272 460352 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 304080 437920 316272 438592 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 304080 427040 316272 427712 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 304080 416160 316272 416832 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 304080 394400 316272 395072 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 304080 448800 316272 449472 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 315912 493032 402100 493392 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 383520 512920 384192 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 372640 512920 373312 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 491874 355604 493760 355952 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 361760 512920 362432 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 340000 512920 340672 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 329120 512920 329792 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 383520 407932 384192 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 372640 407932 373312 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 361760 407932 362432 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 340000 407932 340672 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 329120 407932 329792 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 407572 348060 493760 348420 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 407572 353892 493760 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 318240 512920 318912 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 307360 512920 308032 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 296480 512920 297152 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 285600 512920 286272 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 274720 512920 275392 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 263840 512920 264512 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 318240 407932 318912 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 307360 407932 308032 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 296480 407932 297152 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 285600 407932 286272 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 274720 407932 275392 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 263840 407932 264512 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 304080 383520 316272 384192 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 304080 372640 316272 373312 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 304080 361760 316272 362432 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 304080 340000 316272 340672 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 304080 329120 316272 329792 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 304080 318240 316272 318912 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 304080 350880 512920 351552 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 315912 348060 402100 348420 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 315912 353892 402100 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 159108 481440 165300 482112 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 159108 470560 165300 471232 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 159108 459680 165300 460352 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 159108 437920 165300 438592 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 159108 427040 165300 427712 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 164940 399672 166866 400020 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 159108 416160 165300 416832 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 159108 394400 165300 395072 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 159108 448800 165300 449472 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 19968 491332 21894 491680 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 492320 16991 492992 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 481440 20328 482112 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 470560 20328 471232 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 459680 20328 460352 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 437920 20328 438592 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 427040 20328 427712 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 416160 20328 416832 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 19968 399672 21894 400020 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 394400 20328 395072 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 448800 20328 449472 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 19968 493032 159468 493392 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 19968 407204 159468 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 19968 401372 159468 401732 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 159108 383520 165300 384192 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 159108 372640 165300 373312 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 159108 361760 165300 362432 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 159108 350880 165300 351552 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 159108 340000 165300 340672 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 159108 329120 165300 329792 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 195930 302012 197816 302360 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 159108 318240 165300 318912 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 383520 20328 384192 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 372640 20328 373312 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 361760 20328 362432 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 350880 20328 351552 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 340000 20328 340672 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 329120 20328 329792 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 296480 111988 297152 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 285600 111988 286272 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 274720 111988 275392 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 263840 111988 264512 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 318240 20328 318912 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 19968 302012 21854 302360 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 296480 20328 297152 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 285600 20328 286272 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 274720 20328 275392 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 263840 20328 264512 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 19968 303712 106156 304072 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 19968 315544 159468 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 111628 303712 197816 304072 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 0 510544 513728 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 503200 512920 503872 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 164940 493032 304440 493392 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 164940 407204 304440 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 164940 401372 304440 401732 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 405280 316272 405952 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 164940 315544 304440 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 307360 316272 308032 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 296480 316272 297152 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 285600 316272 286272 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 274720 316272 275392 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 263840 316272 264512 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 252960 512920 253632 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 242080 512920 242752 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 231200 512920 231872 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 491874 210632 493760 210980 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 220320 512920 220992 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 495040 209440 512920 210112 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 491834 195388 493760 195736 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 252960 407932 253632 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 242080 407932 242752 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 231200 407932 231872 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 401740 220320 407932 220992 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 400214 210632 402100 210980 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 407572 208920 493760 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 187680 512920 188352 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 176800 512920 177472 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 165920 512920 166592 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 155040 512920 155712 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 144160 512920 144832 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 133280 512920 133952 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 348428 187680 354620 188352 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 348428 176800 354620 177472 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 348428 165920 354620 166592 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 348428 155040 354620 155712 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 348428 144160 354620 144832 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 348428 133280 354620 133952 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 315912 208920 402100 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 354260 197088 493760 197448 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 122400 512920 123072 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 100640 512920 101312 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 111520 512920 112192 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 89760 512920 90432 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 78880 512920 79552 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 68000 512920 68672 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 57120 512920 57792 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 46240 512920 46912 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 35360 512920 36032 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 491834 21312 493760 21660 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 493400 24480 512920 25152 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 346862 112972 348788 113320 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 348428 122400 354620 123072 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 348428 100640 354620 101312 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 348428 111520 354620 112192 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 348428 89760 354620 90432 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 348428 78880 354620 79552 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 348428 68000 354620 68672 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 348428 57120 354620 57792 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 348428 46240 354620 46912 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 348428 35360 354620 36032 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 346862 21312 348788 21660 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 348428 24480 354620 25152 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 354260 19600 493760 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 354260 105428 493760 105788 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 354260 111260 493760 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 176800 209648 177472 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 187680 209648 188352 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 165920 209648 166592 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 195930 157040 197816 157388 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 144160 209648 144832 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 155040 209648 155712 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 133280 209648 133952 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 252960 111988 253632 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 242080 111988 242752 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 231200 111988 231872 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 220320 111988 220992 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 209440 111988 210112 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 198560 111988 199232 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 252960 20328 253632 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 242080 20328 242752 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 231200 20328 231872 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 220320 20328 220992 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 209440 20328 210112 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 198560 20328 199232 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 187680 111988 188352 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 176800 111988 177472 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 165920 111988 166592 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 155040 111988 155712 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 144160 111988 144832 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 133280 111988 133952 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 187680 20328 188352 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 176800 20328 177472 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 165920 20328 166592 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 19968 157040 21854 157388 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 155040 20328 155712 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 144160 20328 144832 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 133280 20328 133952 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 19968 158740 106156 159100 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 19968 164572 106156 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 111628 158740 197816 159100 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 111628 164572 197816 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 122400 209648 123072 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 100640 209648 101312 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 111520 209648 112192 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 89760 209648 90432 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 78880 209648 79552 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 68000 209648 68672 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 57120 209648 57792 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 46240 209648 46912 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 35360 209648 36032 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 24480 209648 25152 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 122400 111988 123072 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 100640 111988 101312 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 111520 111988 112192 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 89760 111988 90432 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 78880 111988 79552 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 68000 111988 68672 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 122400 20328 123072 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 100640 20328 101312 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 111520 20328 112192 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 89760 20328 90432 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 78880 20328 79552 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 68000 20328 68672 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 57120 111988 57792 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 46240 111988 46912 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 35360 111988 36032 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 105796 24480 111988 25152 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 57120 20328 57792 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 46240 20328 46912 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 35360 20328 36032 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 24480 20328 25152 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 19968 19600 106156 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 111628 19600 197816 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 252960 316272 253632 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 242080 316272 242752 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 231200 316272 231872 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 220320 316272 220992 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 209440 310753 210112 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 209288 197088 348788 197448 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 197456 198560 512920 199232 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 209288 111260 348788 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 209288 105428 348788 105788 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 209288 19600 348788 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 0 816 513728 2448 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 808 13600 512920 14272 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 400040 491332 400388 491680 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 302380 491332 302728 491680 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 491700 355604 492048 355952 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 166652 399672 167000 400020 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 21680 491332 22028 491680 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 21680 399672 22028 400020 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 195756 302012 196104 302360 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 21680 302012 22028 302360 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 491700 210632 492048 210980 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 491700 195388 492048 195736 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 400040 210632 400388 210980 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 353600 197088 354620 197448 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 491700 21312 492048 21660 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 353600 105428 354620 105788 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 353600 111260 354620 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 346728 112972 347076 113320 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 353600 19600 354620 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 346728 21312 347076 21660 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 195756 157040 196104 157388 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 21680 157040 22028 157388 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 484160 493032 484832 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 451520 493032 452192 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 462400 493032 463072 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 473280 493032 473952 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 418880 493032 419552 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 429760 493032 430432 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 440640 493032 441312 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 408000 493872 408672 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 386240 493032 386912 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 397120 493032 397792 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 353600 493032 354272 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 364480 493032 365152 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 375360 493032 376032 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 331840 493032 332512 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 342720 493032 343392 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 352104 493032 352776 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 299200 493032 299872 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 266560 493032 267232 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 277440 493032 278112 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 288320 493032 288992 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 320960 493032 321632 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 299200 401372 299872 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 277440 401372 278112 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 266560 401372 267232 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 288320 401372 288992 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 304080 407204 304440 493392 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 484160 348060 484832 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 473280 348060 473952 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 451520 348060 452192 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 462400 348060 463072 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 408000 350880 408672 351554 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 386240 348060 386912 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 397120 348060 397792 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 418880 348060 419552 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 429760 348060 430432 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 440640 348060 441312 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 375360 348060 376032 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 364480 348060 365152 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 353600 348060 354272 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 352104 348060 352776 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 342720 348060 343392 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 331840 348060 332512 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 320960 348060 321632 354252 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 304080 315544 304440 401732 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 315912 353892 316272 493392 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 401740 353892 402100 493392 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 407572 353892 407932 493392 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 493400 353892 493760 493392 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 255680 493032 256352 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 244800 493032 245472 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 233920 493032 234592 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 201280 493032 201952 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 212160 493032 212832 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 223040 493032 223712 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 168640 493032 169312 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 179520 493032 180192 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 190400 493032 191072 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 136000 493032 136672 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 146880 493032 147552 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 157760 493032 158432 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 255680 401372 256352 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 244800 401372 245472 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 233920 401372 234592 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 223040 401372 223712 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 212160 401372 212832 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 201280 401372 201952 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 190400 401372 191072 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 179520 401372 180192 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 168640 401372 169312 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 157760 401372 158432 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 146880 401372 147552 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 136000 401372 136672 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 159108 407204 159468 493392 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 164940 407204 165300 493392 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 125120 493032 125792 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 103360 493032 104032 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 109404 493032 110076 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 114240 493032 114912 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 70720 493032 71392 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 81600 493032 82272 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 92480 493032 93152 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 38080 493032 38752 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 48960 493032 49632 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 59840 493032 60512 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 27200 493032 27872 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 125120 401372 125792 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 114240 401372 114912 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 109404 401372 110076 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 103360 401372 104032 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 92480 401372 93152 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 81600 401372 82272 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 70720 401372 71392 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 59840 401372 60512 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 48960 401372 49632 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 38080 401372 38752 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 27200 401372 27872 407564 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 19968 407204 20328 493392 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 168640 303712 169312 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 179520 303712 180192 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 190400 303712 191072 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 136000 303712 136672 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 146880 303712 147552 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 157760 303712 158432 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 103360 303712 104032 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 114240 303712 114912 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 125120 303712 125792 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 92480 303712 93152 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 81600 303712 82272 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 70720 303712 71392 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 59840 303712 60512 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 48960 303712 49632 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 38080 303712 38752 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 27200 303712 27872 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 162704 303712 163376 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 19968 315544 20328 401732 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 159108 315544 159468 401732 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 164940 315544 165300 401732 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 484160 197088 484832 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 451520 197088 452192 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 462400 197088 463072 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 473280 197088 473952 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 418880 197088 419552 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 429760 197088 430432 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 440640 197088 441312 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 397120 197088 397792 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 386240 197088 386912 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 408000 197088 408672 208440 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 375360 197088 376032 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 364480 197088 365152 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 353600 197088 354272 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 342720 197088 343392 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 331840 197088 332512 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 320960 197088 321632 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 484160 105428 484832 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 473280 105428 473952 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 462400 105428 463072 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 451520 105428 452192 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 440640 105428 441312 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 429760 105428 430432 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 418880 105428 419552 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 405504 105428 406176 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 408000 105428 408672 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 397120 105428 397792 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 386240 105428 386912 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 484160 816 484832 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 473280 816 473952 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 451520 816 452192 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 462400 816 463072 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 418880 816 419552 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 429760 816 430432 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 440640 816 441312 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 386240 816 386912 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 397120 816 397792 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 405504 816 406176 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 408000 816 408672 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 493400 19600 493760 105788 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 375360 105428 376032 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 364480 105428 365152 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 353600 105428 354272 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 342720 105428 343392 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 331840 105428 332512 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 310080 105428 310752 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 299200 105428 299872 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 277440 105428 278112 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 266560 105428 267232 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 288320 105428 288992 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 320960 105428 321632 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 375360 816 376032 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 364480 816 365152 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 353600 816 354272 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 331840 816 332512 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 342720 816 343392 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 299200 816 299872 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 310080 816 310752 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 266560 816 267232 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 277440 816 278112 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 288320 816 288992 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 320960 816 321632 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 348428 19600 348788 105788 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 354260 19600 354620 105788 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 352104 816 352776 209280 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 348428 111260 348788 197448 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 354260 111260 354620 197448 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 493400 111260 493760 197448 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 190400 158740 191072 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 179520 158740 180192 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 168640 158740 169312 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 162704 158740 163376 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 157760 158740 158432 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 146880 158740 147552 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 136000 158740 136672 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 103360 158740 104032 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 114240 158740 114912 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 125120 158740 125792 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 81600 158740 82272 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 70720 158740 71392 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 92480 158740 93152 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 27200 158740 27872 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 38080 158740 38752 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 48960 158740 49632 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 59840 158740 60512 164932 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 255680 105428 256352 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 244800 105428 245472 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 233920 105428 234592 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 223040 105428 223712 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 212160 105428 212832 111620 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 233920 816 234592 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 244800 816 245472 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 255680 816 256352 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 212160 816 212832 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 223040 816 223712 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 162704 816 163376 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 168640 816 169312 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 179520 816 180192 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 190400 816 191072 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 136000 816 136672 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 146880 816 147552 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 157760 816 158432 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 209288 19600 209648 105788 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 103360 816 104032 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 114240 816 114912 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 125120 816 125792 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 70720 816 71392 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 81600 816 82272 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 92480 816 93152 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 38080 816 38752 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 48960 816 49632 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 59840 816 60512 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 27200 816 27872 19960 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 209288 111260 209648 197448 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 19968 19600 20328 159100 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 105796 19600 106156 159100 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 111628 19600 111988 159100 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 197456 19600 197816 159100 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 511288 0 512920 512992 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 405504 197088 406176 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 495040 816 495712 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 505920 816 506592 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 401740 208920 402100 348420 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 407572 208920 407932 348420 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 493400 208920 493760 348420 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 299200 197088 299872 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 310080 197088 310752 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 315912 208920 316272 348420 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 266560 197088 267232 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 277440 197088 278112 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 288320 197088 288992 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 212160 197088 212832 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 223040 197088 223712 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 233920 197088 234592 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 244800 197088 245472 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 255680 197088 256352 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 201280 816 201952 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 197456 164572 197816 304072 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 808 0 2440 512992 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 109404 816 110076 315904 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 5440 816 6112 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 16320 816 16992 512176 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 19968 164572 20328 304072 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 105796 164572 106156 304072 6 VSS
port 30 nsew ground bidirectional
rlabel metal4 s 111628 164572 111988 304072 6 VSS
port 30 nsew ground bidirectional
rlabel metal5 s 512096 508096 513728 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 0 508096 1632 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 512096 3264 513728 4896 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 0 3264 1632 4896 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 508840 511360 510472 512992 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 508840 0 510472 1632 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 3256 511360 4888 512992 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 3256 0 4888 1632 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 491020 490652 491368 491000 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 303360 407924 303720 408672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 301700 398992 302048 399340 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 497760 353600 498432 354272 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 318304 356284 318652 356632 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 312800 353600 313472 354272 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 167332 490652 167680 491000 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 165660 407924 166020 408672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 158388 407924 158748 408672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 22360 490652 22708 491000 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 20688 407924 21048 408672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 22360 398992 22708 399340 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 491020 211312 491368 211660 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 356652 194708 357000 195056 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 346048 194708 346396 195056 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 318304 211312 318652 211660 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 356652 103048 357000 103396 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 346048 103048 346396 103396 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 195076 166964 195424 167312 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 195076 156360 195424 156708 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 22360 166964 22708 167312 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 22360 21992 22708 22340 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 491194 490652 493040 491000 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 484160 510472 484832 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 473280 510472 473952 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 462400 510472 463072 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 451520 510472 452192 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 484160 408652 484832 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 473280 408652 473952 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 451520 408652 452192 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 462400 408652 463072 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 408292 492312 493040 492672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 440640 510472 441312 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 429760 510472 430432 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 418880 510472 419552 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 408000 510472 408672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 397120 510472 397792 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 386240 510472 386912 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 440640 408652 441312 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 418880 408652 419552 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 429760 408652 430432 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 408000 408652 408672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 386240 408652 386912 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 397120 408652 397792 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 303360 484160 316992 484832 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 303360 473280 316992 473952 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 303360 451520 316992 452192 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 303360 462400 316992 463072 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 303360 440640 316992 441312 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 303360 418880 316992 419552 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 303360 429760 316992 430432 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 303360 408000 316992 408672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 303360 386240 316992 386912 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 303360 397120 316992 397792 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 301700 399166 302048 401012 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 316632 492312 401380 492672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 375360 510472 376032 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 497762 353600 510472 354272 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 364480 510472 365152 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 342720 510472 343392 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 331840 510472 332512 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 320960 510472 321632 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 375360 408652 376032 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 364480 408652 365152 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 342720 408652 343392 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 320960 408652 321632 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 331840 408652 332512 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 408292 347340 493040 347700 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 408292 354612 493040 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 310080 510472 310752 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 299200 510472 299872 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 277440 510472 278112 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 266560 510472 267232 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 288320 510472 288992 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 310080 408652 310752 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 299200 408652 299872 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 277440 408652 278112 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 266560 408652 267232 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 288320 408652 288992 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 303360 375360 316992 376032 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 316632 356284 318478 356632 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 303360 353600 313471 354272 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 303360 364480 316992 365152 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 303360 342720 316992 343392 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 303360 320960 316992 321632 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 303360 331840 316992 332512 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 316632 347340 401380 347700 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 316632 354612 401380 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 167332 490826 167680 492672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 158388 484160 166020 484832 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 158388 473280 166020 473952 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 158388 462400 166020 463072 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 158388 451520 166020 452192 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 158388 440640 166020 441312 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 158388 429760 166020 430432 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 158388 418880 166020 419552 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 158388 408000 166020 408672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 158388 397120 166020 397792 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 158388 386240 166020 386912 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 20688 490652 22574 491000 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 484160 21048 484832 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 473280 21048 473952 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 462400 21048 463072 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 451520 21048 452192 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 440640 21048 441312 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 429760 21048 430432 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 418880 21048 419552 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 408000 21048 408672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 20688 398992 22574 399340 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 397120 21048 397792 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 386240 21048 386912 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 20688 492312 158748 492672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 20688 407924 158748 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 20688 400652 158748 401012 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 158388 375360 166020 376032 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 158388 364480 166020 365152 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 158388 353600 166020 354272 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 158388 342720 166020 343392 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 158388 331840 166020 332512 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 158388 320960 166020 321632 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 375360 21048 376032 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 364480 21048 365152 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 353600 21048 354272 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 342720 21048 343392 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 331840 21048 332512 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 320960 21048 321632 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 299200 112708 299872 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 277440 112708 278112 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 266560 112708 267232 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 288320 112708 288992 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 299200 21048 299872 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 277440 21048 278112 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 266560 21048 267232 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 288320 21048 288992 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 20688 302992 105436 303352 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 20688 316264 158748 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 112348 302992 197096 303352 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 505920 510472 506592 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 0 508096 513728 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 495040 510472 495712 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 165660 492312 303720 492672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 165660 400652 303720 401012 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 165660 407924 303720 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 310080 316992 310752 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 165660 316264 303720 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 299200 316992 299872 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 277440 316992 278112 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 266560 316992 267232 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 288320 316992 288992 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 255680 510472 256352 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 244800 510472 245472 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 233920 510472 234592 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 491194 211312 493040 211660 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 223040 510472 223712 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 212160 510472 212832 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 244800 408652 245472 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 255680 408652 256352 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 233920 408652 234592 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 212160 408652 212832 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 401020 223040 408652 223712 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 408292 209640 493040 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 190400 510472 191072 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 179520 510472 180192 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 168640 510472 169312 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 157760 510472 158432 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 146880 510472 147552 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 136000 510472 136672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 356652 194882 357000 196728 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 346048 194882 346396 196728 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 316632 211312 318478 211660 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 347708 190400 355340 191072 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 347708 179520 355340 180192 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 347708 168640 355340 169312 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 347708 157760 355340 158432 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 347708 146880 355340 147552 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 347708 136000 355340 136672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 316632 209640 401380 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 354980 196368 493040 196728 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 125120 510472 125792 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 114240 510472 114912 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 103360 510472 104032 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 92480 510472 93152 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 81600 510472 82272 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 70720 510472 71392 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 59840 510472 60512 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 48960 510472 49632 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 38080 510472 38752 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 492680 27200 510472 27872 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 356652 103222 357000 105068 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 346048 103222 346396 105068 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 347708 125120 355340 125792 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 347708 114240 355340 114912 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 347708 103360 355340 104032 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 347708 92480 355340 93152 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 347708 81600 355340 82272 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 347708 70720 355340 71392 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 347708 59840 355340 60512 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 347708 48960 355340 49632 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 347708 38080 355340 38752 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 347708 27200 355340 27872 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 354980 20320 493040 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 354980 104708 493040 105068 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 354980 111980 493040 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 179520 210368 180192 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 190400 210368 191072 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 195250 166964 197096 167312 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 168640 210368 169312 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 153824 198968 154496 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 195250 156360 197096 156708 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 198296 157760 210368 158432 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 146880 210368 147552 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 136000 210368 136672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 244800 112708 245472 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 255680 112708 256352 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 233920 112708 234592 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 212160 112708 212832 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 223040 112708 223712 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 201280 112708 201952 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 255680 21048 256352 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 244800 21048 245472 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 233920 21048 234592 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 223040 21048 223712 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 212160 21048 212832 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 201280 21048 201952 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 179520 112708 180192 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 190400 112708 191072 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 168640 112708 169312 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 106636 157760 111148 158432 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 153824 107308 154496 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 110476 153824 112708 154496 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 146880 112708 147552 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 136000 112708 136672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 190400 21048 191072 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 179520 21048 180192 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 20688 166964 22534 167312 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 168640 21048 169312 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 18816 153824 21048 154496 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 157760 19488 158432 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 146880 21048 147552 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 136000 21048 136672 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 20688 158020 105436 158380 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 20688 165292 105436 165652 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 112348 158020 197096 158380 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 112348 165292 197096 165652 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 114240 210368 114912 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 125120 210368 125792 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 103360 210368 104032 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 81600 210368 82272 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 92480 210368 93152 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 70720 210368 71392 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 48960 210368 49632 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 59840 210368 60512 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 38080 210368 38752 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 27200 210368 27872 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 114240 112708 114912 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 125120 112708 125792 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 103360 112708 104032 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 81600 112708 82272 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 92480 112708 93152 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 70720 112708 71392 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 125120 21048 125792 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 114240 21048 114912 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 103360 21048 104032 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 92480 21048 93152 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 81600 21048 82272 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 70720 21048 71392 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 48960 112708 49632 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 59840 112708 60512 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 38080 112708 38752 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 105076 27200 112708 27872 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 59840 21048 60512 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 48960 21048 49632 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 38080 21048 38752 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 20688 21992 22534 22340 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 27200 21048 27872 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 20688 20320 105436 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 112348 20320 197096 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 255680 316992 256352 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 244800 316992 245472 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 233920 316992 234592 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 223040 316992 223712 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 212160 316992 212832 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 196736 201280 510472 201952 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 210008 196368 348068 196728 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 210008 104708 348068 105068 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 210008 111980 348068 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 16320 510472 16992 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 210008 20320 348068 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 3256 5440 510472 6112 6 VDD
port 31 nsew power bidirectional
rlabel metal5 s 0 3264 513728 4896 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 491020 490652 491368 491000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 301700 398992 302048 399340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 318304 356284 318652 356632 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 167332 490652 167680 491000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 22360 490652 22708 491000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 22360 398992 22708 399340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 491020 211312 491368 211660 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 356652 194708 357000 195056 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 346048 194708 346396 195056 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 318304 211312 318652 211660 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 356652 103048 357000 103396 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 346048 103048 346396 103396 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 195076 166964 195424 167312 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 195076 156360 195424 156708 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 22360 166964 22708 167312 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 18816 153824 19712 154496 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 22360 21992 22708 22340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 486880 492312 487552 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 454240 492312 454912 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 465120 492312 465792 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 476000 492312 476672 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 421600 492312 422272 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 432480 492312 433152 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 443360 492312 444032 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 388960 492312 389632 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 399840 492312 400512 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 410720 492312 411392 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 356320 492312 356992 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 367200 492312 367872 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 378080 492312 378752 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 323680 492312 324352 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 334560 492312 335232 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 345440 492312 346112 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 350304 492312 350976 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 291040 492312 291712 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 301920 492312 302592 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 258400 492312 259072 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 269280 492312 269952 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 280160 492312 280832 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 291040 400652 291712 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 301920 400652 302592 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 258400 400652 259072 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 269280 400652 269952 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 280160 400652 280832 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 303360 407924 303720 492672 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 454240 347340 454912 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 465120 347340 465792 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 476000 347340 476672 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 486880 347340 487552 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 388960 347340 389632 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 399840 347340 400512 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 410720 347340 411392 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 421600 347340 422272 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 432480 347340 433152 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 443360 347340 444032 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 367200 347340 367872 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 356320 347340 356992 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 378080 347340 378752 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 350304 347340 350976 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 345440 347340 346112 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 334560 347340 335232 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 323680 347340 324352 354972 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 303360 316264 303720 401012 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 316632 354612 316992 492672 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 401020 354612 401380 492672 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 408292 354612 408652 492672 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 492680 354612 493040 492672 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 225760 492312 226432 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 236640 492312 237312 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 247520 492312 248192 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 193120 492312 193792 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 204000 492312 204672 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 214880 492312 215552 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 171360 492312 172032 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 182240 492312 182912 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 138720 492312 139392 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 149600 492312 150272 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 225760 400652 226432 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 236640 400652 237312 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 247520 400652 248192 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 193120 400652 193792 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 204000 400652 204672 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 214880 400652 215552 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 171360 400652 172032 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 182240 400652 182912 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 138720 400652 139392 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 149600 400652 150272 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 158388 407924 158748 492672 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 165660 407924 166020 492672 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 106080 492312 106752 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 107604 492312 108276 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 116960 492312 117632 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 73440 492312 74112 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 84320 492312 84992 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 95200 492312 95872 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 40800 492312 41472 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 51680 492312 52352 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 62560 492312 63232 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 29920 492312 30592 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 106080 400652 106752 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 107604 400652 108276 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 116960 400652 117632 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 73440 400652 74112 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 84320 400652 84992 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 95200 400652 95872 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 40800 400652 41472 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 51680 400652 52352 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 62560 400652 63232 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 29920 400652 30592 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 20688 407924 21048 492672 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 127840 492312 128512 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 127840 400652 128512 408284 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 193120 302992 193792 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 171360 302992 172032 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 182240 302992 182912 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 138720 302992 139392 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 149600 302992 150272 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 106080 310075 106752 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 116960 302992 117632 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 73440 302992 74112 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 84320 302992 84992 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 95200 302992 95872 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 40800 302992 41472 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 51680 302992 52352 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 62560 302992 63232 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 29920 302992 30592 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 127840 302992 128512 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 160480 302992 161152 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 20688 316264 21048 401012 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 158388 316264 158748 401012 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 165660 316264 166020 401012 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 486880 196368 487552 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 454240 196368 454912 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 465120 196368 465792 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 476000 196368 476672 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 421600 196368 422272 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 432480 196368 433152 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 443360 196368 444032 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 388960 196368 389632 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 399840 196368 400512 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 410720 196368 411392 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 356320 196368 356992 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 367200 196368 367872 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 378080 196368 378752 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 323680 196368 324352 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 334560 196368 335232 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 345440 196368 346112 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 486880 104708 487552 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 454240 104708 454912 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 465120 104708 465792 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 476000 104708 476672 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 421600 104708 422272 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 432480 104708 433152 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 443360 104708 444032 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 388960 104708 389632 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 399840 104708 400512 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 403704 104708 404376 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 410720 104708 411392 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 486880 3264 487552 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 454240 3264 454912 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 465120 3264 465792 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 476000 3264 476672 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 421600 3264 422272 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 432480 3264 433152 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 443360 3264 444032 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 388960 3264 389632 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 399840 3264 400512 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 403704 3264 404376 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 410720 3264 411392 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 492680 20320 493040 105068 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 356320 104708 356992 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 367200 104708 367872 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 378080 104708 378752 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 323680 104708 324352 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 334560 104708 335232 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 345440 104708 346112 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 291040 104708 291712 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 301920 104708 302592 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 312800 104708 313472 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 258400 104708 259072 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 269280 104708 269952 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 280160 104708 280832 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 356320 3264 356992 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 367200 3264 367872 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 378080 3264 378752 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 323680 3264 324352 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 334560 3264 335232 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 345440 3264 346112 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 291040 3264 291712 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 301920 3264 302592 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 312800 3264 313472 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 258400 3264 259072 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 269280 3264 269952 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 280160 3264 280832 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 347708 20320 348068 105068 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 354980 20320 355340 105068 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 350304 3264 350976 210000 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 347708 111980 348068 196728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 354980 111980 355340 196728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 492680 111980 493040 196728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 198296 153824 198968 158432 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 193120 158020 193792 165652 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 171360 158020 172032 165652 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 182240 158020 182912 165652 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 149600 158020 150272 165652 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 138720 158020 139392 165652 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 160480 158020 161152 165652 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 106636 153824 107308 158432 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 110476 153824 111148 158432 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 116960 158020 117632 165652 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 95200 158020 95872 165652 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 84320 158020 84992 165652 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 73440 158020 74112 165652 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 18816 153824 19488 158432 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 29920 158020 30592 165652 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 40800 158020 41472 165652 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 51680 158020 52352 165652 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 62560 158020 63232 165652 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 127840 158020 128512 165652 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 225760 104708 226432 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 236640 104708 237312 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 247520 104708 248192 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 214880 104708 215552 112340 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 225760 3264 226432 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 236640 3264 237312 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 247520 3264 248192 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 193120 3264 193792 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 214880 3264 215552 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 171360 3264 172032 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 182240 3264 182912 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 138720 3264 139392 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 149600 3264 150272 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 160480 3264 161152 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 210008 20320 210368 105068 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 106080 3264 106752 16993 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 116960 3264 117632 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 73440 3264 74112 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 84320 3264 84992 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 95200 3264 95872 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 40800 3264 41472 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 51680 3264 52352 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 62560 3264 63232 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 29920 3264 30592 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 127840 3264 128512 20680 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 210008 111980 210368 196728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 20688 20320 21048 158380 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 105076 20320 105436 158380 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 112348 20320 112708 158380 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 196736 20320 197096 158380 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 492680 209640 493040 347700 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 408292 209640 408652 347700 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 401020 209640 401380 347700 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 497760 3264 498432 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 403704 196368 404376 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 508840 0 510472 512992 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 316632 209640 316992 347700 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 312800 196368 313472 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 301920 196368 302592 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 291040 196368 291712 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 280160 196368 280832 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 269280 196368 269952 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 258400 196368 259072 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 196736 165292 197096 303352 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 204000 3264 204672 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 247520 196368 248192 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 236640 196368 237312 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 225760 196368 226432 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 214880 196368 215552 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 112348 165292 112708 303352 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 105076 165292 105436 303352 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 20688 165292 21048 303352 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 19040 3264 19712 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 8160 3264 8832 509728 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 107604 3264 108276 316624 6 VDD
port 31 nsew power bidirectional
rlabel metal4 s 3256 0 4888 512992 6 VDD
port 31 nsew power bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 513728 512992
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
