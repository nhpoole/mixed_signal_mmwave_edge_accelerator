magic
tech sky130A
timestamp 1626486988
<< checkpaint >>
rect -720 -798 720 798
<< metal4 >>
rect -90 139 90 168
rect -90 21 -59 139
rect 59 21 90 139
rect -90 -168 90 21
<< via4 >>
rect -59 21 59 139
<< metal5 >>
rect -90 139 90 168
rect -90 21 -59 139
rect 59 21 90 139
rect -90 -168 90 21
<< end >>
