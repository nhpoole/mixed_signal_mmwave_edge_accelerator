magic
tech sky130A
magscale 1 2
timestamp 1624237933
<< nwell >>
rect -12316 15828 -7807 16346
rect 11254 16156 35770 30898
rect -12316 15507 -7032 15828
rect -12316 15506 -7807 15507
<< pwell >>
rect -10458 15448 -10428 15450
rect -10458 15412 -10407 15448
rect -12316 14792 -10407 15412
rect -10348 15267 -10162 15449
rect -7858 15448 -7828 15450
rect -7858 15412 -7807 15448
rect -10183 15263 -10162 15267
rect -10183 15229 -10149 15263
rect -9716 14792 -7807 15412
rect -7748 15267 -7562 15449
rect -7298 15267 -7112 15449
rect -7583 15263 -7562 15267
rect -7133 15263 -7112 15267
rect -7583 15229 -7549 15263
rect -7133 15229 -7099 15263
rect -1446 -718 35870 15398
<< nmos >>
rect -12120 15002 -11920 15202
rect -11862 15002 -11662 15202
rect -11604 15002 -11404 15202
rect -11346 15002 -11146 15202
rect -11088 15002 -10888 15202
rect -10830 15002 -10630 15202
rect -9520 15002 -9320 15202
rect -9262 15002 -9062 15202
rect -9004 15002 -8804 15202
rect -8746 15002 -8546 15202
rect -8488 15002 -8288 15202
rect -8230 15002 -8030 15202
rect 13540 13904 14500 14504
rect 14558 13904 15518 14504
rect 15576 13904 16536 14504
rect 16594 13904 17554 14504
rect 17612 13904 18572 14504
rect 18630 13904 19590 14504
rect 19648 13904 20608 14504
rect 20666 13904 21626 14504
rect 21684 13904 22644 14504
rect 22702 13904 23662 14504
rect 23720 13904 24680 14504
rect 24738 13904 25698 14504
rect 25756 13904 26716 14504
rect 26774 13904 27734 14504
rect 27792 13904 28752 14504
rect 28810 13904 29770 14504
rect 29828 13904 30788 14504
rect 30846 13904 31806 14504
rect 31864 13904 32824 14504
rect 32882 13904 33842 14504
rect 13540 13086 14500 13686
rect 14558 13086 15518 13686
rect 15576 13086 16536 13686
rect 16594 13086 17554 13686
rect 17612 13086 18572 13686
rect 18630 13086 19590 13686
rect 19648 13086 20608 13686
rect 20666 13086 21626 13686
rect 21684 13086 22644 13686
rect 22702 13086 23662 13686
rect 23720 13086 24680 13686
rect 24738 13086 25698 13686
rect 25756 13086 26716 13686
rect 26774 13086 27734 13686
rect 27792 13086 28752 13686
rect 28810 13086 29770 13686
rect 29828 13086 30788 13686
rect 30846 13086 31806 13686
rect 31864 13086 32824 13686
rect 32882 13086 33842 13686
rect 13540 11708 14500 12308
rect 14558 11708 15518 12308
rect 15576 11708 16536 12308
rect 16594 11708 17554 12308
rect 17612 11708 18572 12308
rect 18630 11708 19590 12308
rect 19648 11708 20608 12308
rect 20666 11708 21626 12308
rect 21684 11708 22644 12308
rect 22702 11708 23662 12308
rect 23720 11708 24680 12308
rect 24738 11708 25698 12308
rect 25756 11708 26716 12308
rect 26774 11708 27734 12308
rect 27792 11708 28752 12308
rect 28810 11708 29770 12308
rect 29828 11708 30788 12308
rect 30846 11708 31806 12308
rect 31864 11708 32824 12308
rect 32882 11708 33842 12308
rect 13540 10476 14500 11076
rect 14558 10476 15518 11076
rect 15576 10476 16536 11076
rect 16594 10476 17554 11076
rect 17612 10476 18572 11076
rect 18630 10476 19590 11076
rect 19648 10476 20608 11076
rect 20666 10476 21626 11076
rect 21684 10476 22644 11076
rect 22702 10476 23662 11076
rect 23720 10476 24680 11076
rect 24738 10476 25698 11076
rect 25756 10476 26716 11076
rect 26774 10476 27734 11076
rect 27792 10476 28752 11076
rect 28810 10476 29770 11076
rect 29828 10476 30788 11076
rect 30846 10476 31806 11076
rect 31864 10476 32824 11076
rect 32882 10476 33842 11076
rect 13538 9242 14498 9842
rect 14556 9242 15516 9842
rect 15574 9242 16534 9842
rect 16592 9242 17552 9842
rect 17610 9242 18570 9842
rect 18628 9242 19588 9842
rect 19646 9242 20606 9842
rect 20664 9242 21624 9842
rect 21682 9242 22642 9842
rect 22700 9242 23660 9842
rect 23718 9242 24678 9842
rect 24736 9242 25696 9842
rect 25754 9242 26714 9842
rect 26772 9242 27732 9842
rect 27790 9242 28750 9842
rect 28808 9242 29768 9842
rect 29826 9242 30786 9842
rect 30844 9242 31804 9842
rect 31862 9242 32822 9842
rect 32880 9242 33840 9842
rect 13538 8008 14498 8608
rect 14556 8008 15516 8608
rect 15574 8008 16534 8608
rect 16592 8008 17552 8608
rect 17610 8008 18570 8608
rect 18628 8008 19588 8608
rect 19646 8008 20606 8608
rect 20664 8008 21624 8608
rect 21682 8008 22642 8608
rect 22700 8008 23660 8608
rect 23718 8008 24678 8608
rect 24736 8008 25696 8608
rect 25754 8008 26714 8608
rect 26772 8008 27732 8608
rect 27790 8008 28750 8608
rect 28808 8008 29768 8608
rect 29826 8008 30786 8608
rect 30844 8008 31804 8608
rect 31862 8008 32822 8608
rect 32880 8008 33840 8608
rect 13538 6776 14498 7376
rect 14556 6776 15516 7376
rect 15574 6776 16534 7376
rect 16592 6776 17552 7376
rect 17610 6776 18570 7376
rect 18628 6776 19588 7376
rect 19646 6776 20606 7376
rect 20664 6776 21624 7376
rect 21682 6776 22642 7376
rect 22700 6776 23660 7376
rect 23718 6776 24678 7376
rect 24736 6776 25696 7376
rect 25754 6776 26714 7376
rect 26772 6776 27732 7376
rect 27790 6776 28750 7376
rect 28808 6776 29768 7376
rect 29826 6776 30786 7376
rect 30844 6776 31804 7376
rect 31862 6776 32822 7376
rect 32880 6776 33840 7376
rect 13538 5542 14498 6142
rect 14556 5542 15516 6142
rect 15574 5542 16534 6142
rect 16592 5542 17552 6142
rect 17610 5542 18570 6142
rect 18628 5542 19588 6142
rect 19646 5542 20606 6142
rect 20664 5542 21624 6142
rect 21682 5542 22642 6142
rect 22700 5542 23660 6142
rect 23718 5542 24678 6142
rect 24736 5542 25696 6142
rect 25754 5542 26714 6142
rect 26772 5542 27732 6142
rect 27790 5542 28750 6142
rect 28808 5542 29768 6142
rect 29826 5542 30786 6142
rect 30844 5542 31804 6142
rect 31862 5542 32822 6142
rect 32880 5542 33840 6142
rect 13538 4308 14498 4908
rect 14556 4308 15516 4908
rect 15574 4308 16534 4908
rect 16592 4308 17552 4908
rect 17610 4308 18570 4908
rect 18628 4308 19588 4908
rect 19646 4308 20606 4908
rect 20664 4308 21624 4908
rect 21682 4308 22642 4908
rect 22700 4308 23660 4908
rect 23718 4308 24678 4908
rect 24736 4308 25696 4908
rect 25754 4308 26714 4908
rect 26772 4308 27732 4908
rect 27790 4308 28750 4908
rect 28808 4308 29768 4908
rect 29826 4308 30786 4908
rect 30844 4308 31804 4908
rect 31862 4308 32822 4908
rect 32880 4308 33840 4908
rect 13538 3076 14498 3676
rect 14556 3076 15516 3676
rect 15574 3076 16534 3676
rect 16592 3076 17552 3676
rect 17610 3076 18570 3676
rect 18628 3076 19588 3676
rect 19646 3076 20606 3676
rect 20664 3076 21624 3676
rect 21682 3076 22642 3676
rect 22700 3076 23660 3676
rect 23718 3076 24678 3676
rect 24736 3076 25696 3676
rect 25754 3076 26714 3676
rect 26772 3076 27732 3676
rect 27790 3076 28750 3676
rect 28808 3076 29768 3676
rect 29826 3076 30786 3676
rect 30844 3076 31804 3676
rect 31862 3076 32822 3676
rect 32880 3076 33840 3676
rect 13538 1842 14498 2442
rect 14556 1842 15516 2442
rect 15574 1842 16534 2442
rect 16592 1842 17552 2442
rect 17610 1842 18570 2442
rect 18628 1842 19588 2442
rect 19646 1842 20606 2442
rect 20664 1842 21624 2442
rect 21682 1842 22642 2442
rect 22700 1842 23660 2442
rect 23718 1842 24678 2442
rect 24736 1842 25696 2442
rect 25754 1842 26714 2442
rect 26772 1842 27732 2442
rect 27790 1842 28750 2442
rect 28808 1842 29768 2442
rect 29826 1842 30786 2442
rect 30844 1842 31804 2442
rect 31862 1842 32822 2442
rect 32880 1842 33840 2442
rect 908 800 1868 1400
rect 1926 800 2886 1400
rect 2944 800 3904 1400
rect 3962 800 4922 1400
rect 4980 800 5940 1400
rect 5998 800 6958 1400
rect 7016 800 7976 1400
rect 8034 800 8994 1400
rect 9052 800 10012 1400
rect 10070 800 11030 1400
rect 13538 610 14498 1210
rect 14556 610 15516 1210
rect 15574 610 16534 1210
rect 16592 610 17552 1210
rect 17610 610 18570 1210
rect 18628 610 19588 1210
rect 19646 610 20606 1210
rect 20664 610 21624 1210
rect 21682 610 22642 1210
rect 22700 610 23660 1210
rect 23718 610 24678 1210
rect 24736 610 25696 1210
rect 25754 610 26714 1210
rect 26772 610 27732 1210
rect 27790 610 28750 1210
rect 28808 610 29768 1210
rect 29826 610 30786 1210
rect 30844 610 31804 1210
rect 31862 610 32822 1210
rect 32880 610 33840 1210
<< scnmos >>
rect -10270 15293 -10240 15423
rect -7670 15293 -7640 15423
rect -7220 15293 -7190 15423
<< pmos >>
rect 18432 20868 19392 21468
rect 19450 20868 20410 21468
rect 20468 20868 21428 21468
rect 21486 20868 22446 21468
rect 22504 20868 23464 21468
rect 23522 20868 24482 21468
rect 24540 20868 25500 21468
rect 25558 20868 26518 21468
rect 26576 20868 27536 21468
rect 27594 20868 28554 21468
rect 28612 20868 29572 21468
rect 29630 20868 30590 21468
rect 30648 20868 31608 21468
rect 31666 20868 32626 21468
rect 32684 20868 33644 21468
rect 18432 19612 19392 20212
rect 19450 19612 20410 20212
rect 20468 19612 21428 20212
rect 21486 19612 22446 20212
rect 22504 19612 23464 20212
rect 23522 19612 24482 20212
rect 24540 19612 25500 20212
rect 25558 19612 26518 20212
rect 26576 19612 27536 20212
rect 27594 19612 28554 20212
rect 28612 19612 29572 20212
rect 29630 19612 30590 20212
rect 30648 19612 31608 20212
rect 31666 19612 32626 20212
rect 32684 19612 33644 20212
rect 18432 18356 19392 18956
rect 19450 18356 20410 18956
rect 20468 18356 21428 18956
rect 21486 18356 22446 18956
rect 22504 18356 23464 18956
rect 23522 18356 24482 18956
rect 24540 18356 25500 18956
rect 25558 18356 26518 18956
rect 26576 18356 27536 18956
rect 27594 18356 28554 18956
rect 28612 18356 29572 18956
rect 29630 18356 30590 18956
rect 30648 18356 31608 18956
rect 31666 18356 32626 18956
rect 32684 18356 33644 18956
rect 18432 17100 19392 17700
rect 19450 17100 20410 17700
rect 20468 17100 21428 17700
rect 21486 17100 22446 17700
rect 22504 17100 23464 17700
rect 23522 17100 24482 17700
rect 24540 17100 25500 17700
rect 25558 17100 26518 17700
rect 26576 17100 27536 17700
rect 27594 17100 28554 17700
rect 28612 17100 29572 17700
rect 29630 17100 30590 17700
rect 30648 17100 31608 17700
rect 31666 17100 32626 17700
rect 32684 17100 33644 17700
<< scpmoshvt >>
rect -10270 15543 -10240 15743
rect -7670 15543 -7640 15743
rect -7220 15543 -7190 15743
<< pmoslvt >>
rect 17446 27414 18406 28014
rect 18464 27414 19424 28014
rect 19482 27414 20442 28014
rect 20500 27414 21460 28014
rect 21518 27414 22478 28014
rect 22536 27414 23496 28014
rect 23554 27414 24514 28014
rect 24572 27414 25532 28014
rect 25590 27414 26550 28014
rect 26608 27414 27568 28014
rect 27626 27414 28586 28014
rect 28644 27414 29604 28014
rect 29662 27414 30622 28014
rect 30680 27414 31640 28014
rect 31698 27414 32658 28014
rect 32716 27414 33676 28014
rect 17446 26278 18406 26878
rect 18464 26278 19424 26878
rect 19482 26278 20442 26878
rect 20500 26278 21460 26878
rect 21518 26278 22478 26878
rect 22536 26278 23496 26878
rect 23554 26278 24514 26878
rect 24572 26278 25532 26878
rect 25590 26278 26550 26878
rect 26608 26278 27568 26878
rect 27626 26278 28586 26878
rect 28644 26278 29604 26878
rect 29662 26278 30622 26878
rect 30680 26278 31640 26878
rect 31698 26278 32658 26878
rect 32716 26278 33676 26878
rect 17446 25142 18406 25742
rect 18464 25142 19424 25742
rect 19482 25142 20442 25742
rect 20500 25142 21460 25742
rect 21518 25142 22478 25742
rect 22536 25142 23496 25742
rect 23554 25142 24514 25742
rect 24572 25142 25532 25742
rect 25590 25142 26550 25742
rect 26608 25142 27568 25742
rect 27626 25142 28586 25742
rect 28644 25142 29604 25742
rect 29662 25142 30622 25742
rect 30680 25142 31640 25742
rect 31698 25142 32658 25742
rect 32716 25142 33676 25742
rect 18640 23504 19600 24104
rect 19658 23504 20618 24104
rect 20676 23504 21636 24104
rect 21694 23504 22654 24104
rect 22712 23504 23672 24104
rect 23730 23504 24690 24104
rect 24748 23504 25708 24104
rect 25766 23504 26726 24104
rect 26784 23504 27744 24104
rect 27802 23504 28762 24104
rect 28820 23504 29780 24104
rect 29838 23504 30798 24104
rect 30856 23504 31816 24104
rect 31874 23504 32834 24104
rect 18640 22472 19600 23072
rect 19658 22472 20618 23072
rect 20676 22472 21636 23072
rect 21694 22472 22654 23072
rect 22712 22472 23672 23072
rect 23730 22472 24690 23072
rect 24748 22472 25708 23072
rect 25766 22472 26726 23072
rect 26784 22472 27744 23072
rect 27802 22472 28762 23072
rect 28820 22472 29780 23072
rect 29838 22472 30798 23072
rect 30856 22472 31816 23072
rect 31874 22472 32834 23072
rect 13128 20764 14088 21364
rect 14146 20764 15106 21364
rect 15164 20764 16124 21364
rect 16182 20764 17142 21364
rect 13128 19732 14088 20332
rect 14146 19732 15106 20332
rect 15164 19732 16124 20332
rect 16182 19732 17142 20332
rect 13128 18700 14088 19300
rect 14146 18700 15106 19300
rect 15164 18700 16124 19300
rect 16182 18700 17142 19300
rect 13128 17668 14088 18268
rect 14146 17668 15106 18268
rect 15164 17668 16124 18268
rect 16182 17668 17142 18268
<< pmoshvt >>
rect -12120 15726 -11920 16126
rect -11862 15726 -11662 16126
rect -11604 15726 -11404 16126
rect -11346 15726 -11146 16126
rect -11088 15726 -10888 16126
rect -10830 15726 -10630 16126
rect -9520 15726 -9320 16126
rect -9262 15726 -9062 16126
rect -9004 15726 -8804 16126
rect -8746 15726 -8546 16126
rect -8488 15726 -8288 16126
rect -8230 15726 -8030 16126
<< nmoslvt >>
rect 1774 13428 2734 14028
rect 2792 13428 3752 14028
rect 3810 13428 4770 14028
rect 4828 13428 5788 14028
rect 5846 13428 6806 14028
rect 6864 13428 7824 14028
rect 7882 13428 8842 14028
rect 8900 13428 9860 14028
rect 9918 13428 10878 14028
rect 1774 12610 2734 13210
rect 2792 12610 3752 13210
rect 3810 12610 4770 13210
rect 4828 12610 5788 13210
rect 5846 12610 6806 13210
rect 6864 12610 7824 13210
rect 7882 12610 8842 13210
rect 8900 12610 9860 13210
rect 9918 12610 10878 13210
rect 1774 11792 2734 12392
rect 2792 11792 3752 12392
rect 3810 11792 4770 12392
rect 4828 11792 5788 12392
rect 5846 11792 6806 12392
rect 6864 11792 7824 12392
rect 7882 11792 8842 12392
rect 8900 11792 9860 12392
rect 9918 11792 10878 12392
rect 1774 10974 2734 11574
rect 2792 10974 3752 11574
rect 3810 10974 4770 11574
rect 4828 10974 5788 11574
rect 5846 10974 6806 11574
rect 6864 10974 7824 11574
rect 7882 10974 8842 11574
rect 8900 10974 9860 11574
rect 9918 10974 10878 11574
rect 1774 10156 2734 10756
rect 2792 10156 3752 10756
rect 3810 10156 4770 10756
rect 4828 10156 5788 10756
rect 5846 10156 6806 10756
rect 6864 10156 7824 10756
rect 7882 10156 8842 10756
rect 8900 10156 9860 10756
rect 9918 10156 10878 10756
rect 1774 9338 2734 9938
rect 2792 9338 3752 9938
rect 3810 9338 4770 9938
rect 4828 9338 5788 9938
rect 5846 9338 6806 9938
rect 6864 9338 7824 9938
rect 7882 9338 8842 9938
rect 8900 9338 9860 9938
rect 9918 9338 10878 9938
rect 1774 8520 2734 9120
rect 2792 8520 3752 9120
rect 3810 8520 4770 9120
rect 4828 8520 5788 9120
rect 5846 8520 6806 9120
rect 6864 8520 7824 9120
rect 7882 8520 8842 9120
rect 8900 8520 9860 9120
rect 9918 8520 10878 9120
rect 1774 7702 2734 8302
rect 2792 7702 3752 8302
rect 3810 7702 4770 8302
rect 4828 7702 5788 8302
rect 5846 7702 6806 8302
rect 6864 7702 7824 8302
rect 7882 7702 8842 8302
rect 8900 7702 9860 8302
rect 9918 7702 10878 8302
rect 450 5678 1410 6278
rect 1468 5678 2428 6278
rect 2486 5678 3446 6278
rect 3504 5678 4464 6278
rect 4522 5678 5482 6278
rect 5540 5678 6500 6278
rect 6558 5678 7518 6278
rect 7576 5678 8536 6278
rect 8594 5678 9554 6278
rect 9612 5678 10572 6278
rect 10630 5678 11590 6278
rect 450 4566 1410 5166
rect 1468 4566 2428 5166
rect 2486 4566 3446 5166
rect 3504 4566 4464 5166
rect 4522 4566 5482 5166
rect 5540 4566 6500 5166
rect 6558 4566 7518 5166
rect 7576 4566 8536 5166
rect 8594 4566 9554 5166
rect 9612 4566 10572 5166
rect 10630 4566 11590 5166
rect 450 3454 1410 4054
rect 1468 3454 2428 4054
rect 2486 3454 3446 4054
rect 3504 3454 4464 4054
rect 4522 3454 5482 4054
rect 5540 3454 6500 4054
rect 6558 3454 7518 4054
rect 7576 3454 8536 4054
rect 8594 3454 9554 4054
rect 9612 3454 10572 4054
rect 10630 3454 11590 4054
rect 450 2342 1410 2942
rect 1468 2342 2428 2942
rect 2486 2342 3446 2942
rect 3504 2342 4464 2942
rect 4522 2342 5482 2942
rect 5540 2342 6500 2942
rect 6558 2342 7518 2942
rect 7576 2342 8536 2942
rect 8594 2342 9554 2942
rect 9612 2342 10572 2942
rect 10630 2342 11590 2942
<< ndiff >>
rect -10322 15411 -10270 15423
rect -10322 15377 -10314 15411
rect -10280 15377 -10270 15411
rect -10322 15343 -10270 15377
rect -10322 15309 -10314 15343
rect -10280 15309 -10270 15343
rect -10322 15293 -10270 15309
rect -10240 15411 -10188 15423
rect -10240 15377 -10230 15411
rect -10196 15377 -10188 15411
rect -10240 15343 -10188 15377
rect -7722 15411 -7670 15423
rect -7722 15377 -7714 15411
rect -7680 15377 -7670 15411
rect -10240 15309 -10230 15343
rect -10196 15309 -10188 15343
rect -10240 15293 -10188 15309
rect -12178 15190 -12120 15202
rect -12178 15014 -12166 15190
rect -12132 15014 -12120 15190
rect -12178 15002 -12120 15014
rect -11920 15190 -11862 15202
rect -11920 15014 -11908 15190
rect -11874 15014 -11862 15190
rect -11920 15002 -11862 15014
rect -11662 15190 -11604 15202
rect -11662 15014 -11650 15190
rect -11616 15014 -11604 15190
rect -11662 15002 -11604 15014
rect -11404 15190 -11346 15202
rect -11404 15014 -11392 15190
rect -11358 15014 -11346 15190
rect -11404 15002 -11346 15014
rect -11146 15190 -11088 15202
rect -11146 15014 -11134 15190
rect -11100 15014 -11088 15190
rect -11146 15002 -11088 15014
rect -10888 15190 -10830 15202
rect -10888 15014 -10876 15190
rect -10842 15014 -10830 15190
rect -10888 15002 -10830 15014
rect -10630 15190 -10572 15202
rect -10630 15014 -10618 15190
rect -10584 15014 -10572 15190
rect -10630 15002 -10572 15014
rect -7722 15343 -7670 15377
rect -7722 15309 -7714 15343
rect -7680 15309 -7670 15343
rect -7722 15293 -7670 15309
rect -7640 15411 -7588 15423
rect -7640 15377 -7630 15411
rect -7596 15377 -7588 15411
rect -7640 15343 -7588 15377
rect -7640 15309 -7630 15343
rect -7596 15309 -7588 15343
rect -7640 15293 -7588 15309
rect -7272 15411 -7220 15423
rect -7272 15377 -7264 15411
rect -7230 15377 -7220 15411
rect -7272 15343 -7220 15377
rect -7272 15309 -7264 15343
rect -7230 15309 -7220 15343
rect -7272 15293 -7220 15309
rect -7190 15411 -7138 15423
rect -7190 15377 -7180 15411
rect -7146 15377 -7138 15411
rect -7190 15343 -7138 15377
rect -7190 15309 -7180 15343
rect -7146 15309 -7138 15343
rect -7190 15293 -7138 15309
rect -9578 15190 -9520 15202
rect -9578 15014 -9566 15190
rect -9532 15014 -9520 15190
rect -9578 15002 -9520 15014
rect -9320 15190 -9262 15202
rect -9320 15014 -9308 15190
rect -9274 15014 -9262 15190
rect -9320 15002 -9262 15014
rect -9062 15190 -9004 15202
rect -9062 15014 -9050 15190
rect -9016 15014 -9004 15190
rect -9062 15002 -9004 15014
rect -8804 15190 -8746 15202
rect -8804 15014 -8792 15190
rect -8758 15014 -8746 15190
rect -8804 15002 -8746 15014
rect -8546 15190 -8488 15202
rect -8546 15014 -8534 15190
rect -8500 15014 -8488 15190
rect -8546 15002 -8488 15014
rect -8288 15190 -8230 15202
rect -8288 15014 -8276 15190
rect -8242 15014 -8230 15190
rect -8288 15002 -8230 15014
rect -8030 15190 -7972 15202
rect -8030 15014 -8018 15190
rect -7984 15014 -7972 15190
rect -8030 15002 -7972 15014
rect 13482 14492 13540 14504
rect 1716 14016 1774 14028
rect 1716 13440 1728 14016
rect 1762 13440 1774 14016
rect 1716 13428 1774 13440
rect 2734 14016 2792 14028
rect 2734 13440 2746 14016
rect 2780 13440 2792 14016
rect 2734 13428 2792 13440
rect 3752 14016 3810 14028
rect 3752 13440 3764 14016
rect 3798 13440 3810 14016
rect 3752 13428 3810 13440
rect 4770 14016 4828 14028
rect 4770 13440 4782 14016
rect 4816 13440 4828 14016
rect 4770 13428 4828 13440
rect 5788 14016 5846 14028
rect 5788 13440 5800 14016
rect 5834 13440 5846 14016
rect 5788 13428 5846 13440
rect 6806 14016 6864 14028
rect 6806 13440 6818 14016
rect 6852 13440 6864 14016
rect 6806 13428 6864 13440
rect 7824 14016 7882 14028
rect 7824 13440 7836 14016
rect 7870 13440 7882 14016
rect 7824 13428 7882 13440
rect 8842 14016 8900 14028
rect 8842 13440 8854 14016
rect 8888 13440 8900 14016
rect 8842 13428 8900 13440
rect 9860 14016 9918 14028
rect 9860 13440 9872 14016
rect 9906 13440 9918 14016
rect 9860 13428 9918 13440
rect 10878 14016 10936 14028
rect 10878 13440 10890 14016
rect 10924 13440 10936 14016
rect 13482 13916 13494 14492
rect 13528 13916 13540 14492
rect 13482 13904 13540 13916
rect 14500 14492 14558 14504
rect 14500 13916 14512 14492
rect 14546 13916 14558 14492
rect 14500 13904 14558 13916
rect 15518 14492 15576 14504
rect 15518 13916 15530 14492
rect 15564 13916 15576 14492
rect 15518 13904 15576 13916
rect 16536 14492 16594 14504
rect 16536 13916 16548 14492
rect 16582 13916 16594 14492
rect 16536 13904 16594 13916
rect 17554 14492 17612 14504
rect 17554 13916 17566 14492
rect 17600 13916 17612 14492
rect 17554 13904 17612 13916
rect 18572 14492 18630 14504
rect 18572 13916 18584 14492
rect 18618 13916 18630 14492
rect 18572 13904 18630 13916
rect 19590 14492 19648 14504
rect 19590 13916 19602 14492
rect 19636 13916 19648 14492
rect 19590 13904 19648 13916
rect 20608 14492 20666 14504
rect 20608 13916 20620 14492
rect 20654 13916 20666 14492
rect 20608 13904 20666 13916
rect 21626 14492 21684 14504
rect 21626 13916 21638 14492
rect 21672 13916 21684 14492
rect 21626 13904 21684 13916
rect 22644 14492 22702 14504
rect 22644 13916 22656 14492
rect 22690 13916 22702 14492
rect 22644 13904 22702 13916
rect 23662 14492 23720 14504
rect 23662 13916 23674 14492
rect 23708 13916 23720 14492
rect 23662 13904 23720 13916
rect 24680 14492 24738 14504
rect 24680 13916 24692 14492
rect 24726 13916 24738 14492
rect 24680 13904 24738 13916
rect 25698 14492 25756 14504
rect 25698 13916 25710 14492
rect 25744 13916 25756 14492
rect 25698 13904 25756 13916
rect 26716 14492 26774 14504
rect 26716 13916 26728 14492
rect 26762 13916 26774 14492
rect 26716 13904 26774 13916
rect 27734 14492 27792 14504
rect 27734 13916 27746 14492
rect 27780 13916 27792 14492
rect 27734 13904 27792 13916
rect 28752 14492 28810 14504
rect 28752 13916 28764 14492
rect 28798 13916 28810 14492
rect 28752 13904 28810 13916
rect 29770 14492 29828 14504
rect 29770 13916 29782 14492
rect 29816 13916 29828 14492
rect 29770 13904 29828 13916
rect 30788 14492 30846 14504
rect 30788 13916 30800 14492
rect 30834 13916 30846 14492
rect 30788 13904 30846 13916
rect 31806 14492 31864 14504
rect 31806 13916 31818 14492
rect 31852 13916 31864 14492
rect 31806 13904 31864 13916
rect 32824 14492 32882 14504
rect 32824 13916 32836 14492
rect 32870 13916 32882 14492
rect 32824 13904 32882 13916
rect 33842 14492 33900 14504
rect 33842 13916 33854 14492
rect 33888 13916 33900 14492
rect 33842 13904 33900 13916
rect 10878 13428 10936 13440
rect 13482 13674 13540 13686
rect 1716 13198 1774 13210
rect 1716 12622 1728 13198
rect 1762 12622 1774 13198
rect 1716 12610 1774 12622
rect 2734 13198 2792 13210
rect 2734 12622 2746 13198
rect 2780 12622 2792 13198
rect 2734 12610 2792 12622
rect 3752 13198 3810 13210
rect 3752 12622 3764 13198
rect 3798 12622 3810 13198
rect 3752 12610 3810 12622
rect 4770 13198 4828 13210
rect 4770 12622 4782 13198
rect 4816 12622 4828 13198
rect 4770 12610 4828 12622
rect 5788 13198 5846 13210
rect 5788 12622 5800 13198
rect 5834 12622 5846 13198
rect 5788 12610 5846 12622
rect 6806 13198 6864 13210
rect 6806 12622 6818 13198
rect 6852 12622 6864 13198
rect 6806 12610 6864 12622
rect 7824 13198 7882 13210
rect 7824 12622 7836 13198
rect 7870 12622 7882 13198
rect 7824 12610 7882 12622
rect 8842 13198 8900 13210
rect 8842 12622 8854 13198
rect 8888 12622 8900 13198
rect 8842 12610 8900 12622
rect 9860 13198 9918 13210
rect 9860 12622 9872 13198
rect 9906 12622 9918 13198
rect 9860 12610 9918 12622
rect 10878 13198 10936 13210
rect 10878 12622 10890 13198
rect 10924 12622 10936 13198
rect 13482 13098 13494 13674
rect 13528 13098 13540 13674
rect 13482 13086 13540 13098
rect 14500 13674 14558 13686
rect 14500 13098 14512 13674
rect 14546 13098 14558 13674
rect 14500 13086 14558 13098
rect 15518 13674 15576 13686
rect 15518 13098 15530 13674
rect 15564 13098 15576 13674
rect 15518 13086 15576 13098
rect 16536 13674 16594 13686
rect 16536 13098 16548 13674
rect 16582 13098 16594 13674
rect 16536 13086 16594 13098
rect 17554 13674 17612 13686
rect 17554 13098 17566 13674
rect 17600 13098 17612 13674
rect 17554 13086 17612 13098
rect 18572 13674 18630 13686
rect 18572 13098 18584 13674
rect 18618 13098 18630 13674
rect 18572 13086 18630 13098
rect 19590 13674 19648 13686
rect 19590 13098 19602 13674
rect 19636 13098 19648 13674
rect 19590 13086 19648 13098
rect 20608 13674 20666 13686
rect 20608 13098 20620 13674
rect 20654 13098 20666 13674
rect 20608 13086 20666 13098
rect 21626 13674 21684 13686
rect 21626 13098 21638 13674
rect 21672 13098 21684 13674
rect 21626 13086 21684 13098
rect 22644 13674 22702 13686
rect 22644 13098 22656 13674
rect 22690 13098 22702 13674
rect 22644 13086 22702 13098
rect 23662 13674 23720 13686
rect 23662 13098 23674 13674
rect 23708 13098 23720 13674
rect 23662 13086 23720 13098
rect 24680 13674 24738 13686
rect 24680 13098 24692 13674
rect 24726 13098 24738 13674
rect 24680 13086 24738 13098
rect 25698 13674 25756 13686
rect 25698 13098 25710 13674
rect 25744 13098 25756 13674
rect 25698 13086 25756 13098
rect 26716 13674 26774 13686
rect 26716 13098 26728 13674
rect 26762 13098 26774 13674
rect 26716 13086 26774 13098
rect 27734 13674 27792 13686
rect 27734 13098 27746 13674
rect 27780 13098 27792 13674
rect 27734 13086 27792 13098
rect 28752 13674 28810 13686
rect 28752 13098 28764 13674
rect 28798 13098 28810 13674
rect 28752 13086 28810 13098
rect 29770 13674 29828 13686
rect 29770 13098 29782 13674
rect 29816 13098 29828 13674
rect 29770 13086 29828 13098
rect 30788 13674 30846 13686
rect 30788 13098 30800 13674
rect 30834 13098 30846 13674
rect 30788 13086 30846 13098
rect 31806 13674 31864 13686
rect 31806 13098 31818 13674
rect 31852 13098 31864 13674
rect 31806 13086 31864 13098
rect 32824 13674 32882 13686
rect 32824 13098 32836 13674
rect 32870 13098 32882 13674
rect 32824 13086 32882 13098
rect 33842 13674 33900 13686
rect 33842 13098 33854 13674
rect 33888 13098 33900 13674
rect 33842 13086 33900 13098
rect 10878 12610 10936 12622
rect 1716 12380 1774 12392
rect 1716 11804 1728 12380
rect 1762 11804 1774 12380
rect 1716 11792 1774 11804
rect 2734 12380 2792 12392
rect 2734 11804 2746 12380
rect 2780 11804 2792 12380
rect 2734 11792 2792 11804
rect 3752 12380 3810 12392
rect 3752 11804 3764 12380
rect 3798 11804 3810 12380
rect 3752 11792 3810 11804
rect 4770 12380 4828 12392
rect 4770 11804 4782 12380
rect 4816 11804 4828 12380
rect 4770 11792 4828 11804
rect 5788 12380 5846 12392
rect 5788 11804 5800 12380
rect 5834 11804 5846 12380
rect 5788 11792 5846 11804
rect 6806 12380 6864 12392
rect 6806 11804 6818 12380
rect 6852 11804 6864 12380
rect 6806 11792 6864 11804
rect 7824 12380 7882 12392
rect 7824 11804 7836 12380
rect 7870 11804 7882 12380
rect 7824 11792 7882 11804
rect 8842 12380 8900 12392
rect 8842 11804 8854 12380
rect 8888 11804 8900 12380
rect 8842 11792 8900 11804
rect 9860 12380 9918 12392
rect 9860 11804 9872 12380
rect 9906 11804 9918 12380
rect 9860 11792 9918 11804
rect 10878 12380 10936 12392
rect 10878 11804 10890 12380
rect 10924 11804 10936 12380
rect 10878 11792 10936 11804
rect 13482 12296 13540 12308
rect 13482 11720 13494 12296
rect 13528 11720 13540 12296
rect 13482 11708 13540 11720
rect 14500 12296 14558 12308
rect 14500 11720 14512 12296
rect 14546 11720 14558 12296
rect 14500 11708 14558 11720
rect 15518 12296 15576 12308
rect 15518 11720 15530 12296
rect 15564 11720 15576 12296
rect 15518 11708 15576 11720
rect 16536 12296 16594 12308
rect 16536 11720 16548 12296
rect 16582 11720 16594 12296
rect 16536 11708 16594 11720
rect 17554 12296 17612 12308
rect 17554 11720 17566 12296
rect 17600 11720 17612 12296
rect 17554 11708 17612 11720
rect 18572 12296 18630 12308
rect 18572 11720 18584 12296
rect 18618 11720 18630 12296
rect 18572 11708 18630 11720
rect 19590 12296 19648 12308
rect 19590 11720 19602 12296
rect 19636 11720 19648 12296
rect 19590 11708 19648 11720
rect 20608 12296 20666 12308
rect 20608 11720 20620 12296
rect 20654 11720 20666 12296
rect 20608 11708 20666 11720
rect 21626 12296 21684 12308
rect 21626 11720 21638 12296
rect 21672 11720 21684 12296
rect 21626 11708 21684 11720
rect 22644 12296 22702 12308
rect 22644 11720 22656 12296
rect 22690 11720 22702 12296
rect 22644 11708 22702 11720
rect 23662 12296 23720 12308
rect 23662 11720 23674 12296
rect 23708 11720 23720 12296
rect 23662 11708 23720 11720
rect 24680 12296 24738 12308
rect 24680 11720 24692 12296
rect 24726 11720 24738 12296
rect 24680 11708 24738 11720
rect 25698 12296 25756 12308
rect 25698 11720 25710 12296
rect 25744 11720 25756 12296
rect 25698 11708 25756 11720
rect 26716 12296 26774 12308
rect 26716 11720 26728 12296
rect 26762 11720 26774 12296
rect 26716 11708 26774 11720
rect 27734 12296 27792 12308
rect 27734 11720 27746 12296
rect 27780 11720 27792 12296
rect 27734 11708 27792 11720
rect 28752 12296 28810 12308
rect 28752 11720 28764 12296
rect 28798 11720 28810 12296
rect 28752 11708 28810 11720
rect 29770 12296 29828 12308
rect 29770 11720 29782 12296
rect 29816 11720 29828 12296
rect 29770 11708 29828 11720
rect 30788 12296 30846 12308
rect 30788 11720 30800 12296
rect 30834 11720 30846 12296
rect 30788 11708 30846 11720
rect 31806 12296 31864 12308
rect 31806 11720 31818 12296
rect 31852 11720 31864 12296
rect 31806 11708 31864 11720
rect 32824 12296 32882 12308
rect 32824 11720 32836 12296
rect 32870 11720 32882 12296
rect 32824 11708 32882 11720
rect 33842 12296 33900 12308
rect 33842 11720 33854 12296
rect 33888 11720 33900 12296
rect 33842 11708 33900 11720
rect 1716 11562 1774 11574
rect 1716 10986 1728 11562
rect 1762 10986 1774 11562
rect 1716 10974 1774 10986
rect 2734 11562 2792 11574
rect 2734 10986 2746 11562
rect 2780 10986 2792 11562
rect 2734 10974 2792 10986
rect 3752 11562 3810 11574
rect 3752 10986 3764 11562
rect 3798 10986 3810 11562
rect 3752 10974 3810 10986
rect 4770 11562 4828 11574
rect 4770 10986 4782 11562
rect 4816 10986 4828 11562
rect 4770 10974 4828 10986
rect 5788 11562 5846 11574
rect 5788 10986 5800 11562
rect 5834 10986 5846 11562
rect 5788 10974 5846 10986
rect 6806 11562 6864 11574
rect 6806 10986 6818 11562
rect 6852 10986 6864 11562
rect 6806 10974 6864 10986
rect 7824 11562 7882 11574
rect 7824 10986 7836 11562
rect 7870 10986 7882 11562
rect 7824 10974 7882 10986
rect 8842 11562 8900 11574
rect 8842 10986 8854 11562
rect 8888 10986 8900 11562
rect 8842 10974 8900 10986
rect 9860 11562 9918 11574
rect 9860 10986 9872 11562
rect 9906 10986 9918 11562
rect 9860 10974 9918 10986
rect 10878 11562 10936 11574
rect 10878 10986 10890 11562
rect 10924 10986 10936 11562
rect 10878 10974 10936 10986
rect 13482 11064 13540 11076
rect 1716 10744 1774 10756
rect 1716 10168 1728 10744
rect 1762 10168 1774 10744
rect 1716 10156 1774 10168
rect 2734 10744 2792 10756
rect 2734 10168 2746 10744
rect 2780 10168 2792 10744
rect 2734 10156 2792 10168
rect 3752 10744 3810 10756
rect 3752 10168 3764 10744
rect 3798 10168 3810 10744
rect 3752 10156 3810 10168
rect 4770 10744 4828 10756
rect 4770 10168 4782 10744
rect 4816 10168 4828 10744
rect 4770 10156 4828 10168
rect 5788 10744 5846 10756
rect 5788 10168 5800 10744
rect 5834 10168 5846 10744
rect 5788 10156 5846 10168
rect 6806 10744 6864 10756
rect 6806 10168 6818 10744
rect 6852 10168 6864 10744
rect 6806 10156 6864 10168
rect 7824 10744 7882 10756
rect 7824 10168 7836 10744
rect 7870 10168 7882 10744
rect 7824 10156 7882 10168
rect 8842 10744 8900 10756
rect 8842 10168 8854 10744
rect 8888 10168 8900 10744
rect 8842 10156 8900 10168
rect 9860 10744 9918 10756
rect 9860 10168 9872 10744
rect 9906 10168 9918 10744
rect 9860 10156 9918 10168
rect 10878 10744 10936 10756
rect 10878 10168 10890 10744
rect 10924 10168 10936 10744
rect 13482 10488 13494 11064
rect 13528 10488 13540 11064
rect 13482 10476 13540 10488
rect 14500 11064 14558 11076
rect 14500 10488 14512 11064
rect 14546 10488 14558 11064
rect 14500 10476 14558 10488
rect 15518 11064 15576 11076
rect 15518 10488 15530 11064
rect 15564 10488 15576 11064
rect 15518 10476 15576 10488
rect 16536 11064 16594 11076
rect 16536 10488 16548 11064
rect 16582 10488 16594 11064
rect 16536 10476 16594 10488
rect 17554 11064 17612 11076
rect 17554 10488 17566 11064
rect 17600 10488 17612 11064
rect 17554 10476 17612 10488
rect 18572 11064 18630 11076
rect 18572 10488 18584 11064
rect 18618 10488 18630 11064
rect 18572 10476 18630 10488
rect 19590 11064 19648 11076
rect 19590 10488 19602 11064
rect 19636 10488 19648 11064
rect 19590 10476 19648 10488
rect 20608 11064 20666 11076
rect 20608 10488 20620 11064
rect 20654 10488 20666 11064
rect 20608 10476 20666 10488
rect 21626 11064 21684 11076
rect 21626 10488 21638 11064
rect 21672 10488 21684 11064
rect 21626 10476 21684 10488
rect 22644 11064 22702 11076
rect 22644 10488 22656 11064
rect 22690 10488 22702 11064
rect 22644 10476 22702 10488
rect 23662 11064 23720 11076
rect 23662 10488 23674 11064
rect 23708 10488 23720 11064
rect 23662 10476 23720 10488
rect 24680 11064 24738 11076
rect 24680 10488 24692 11064
rect 24726 10488 24738 11064
rect 24680 10476 24738 10488
rect 25698 11064 25756 11076
rect 25698 10488 25710 11064
rect 25744 10488 25756 11064
rect 25698 10476 25756 10488
rect 26716 11064 26774 11076
rect 26716 10488 26728 11064
rect 26762 10488 26774 11064
rect 26716 10476 26774 10488
rect 27734 11064 27792 11076
rect 27734 10488 27746 11064
rect 27780 10488 27792 11064
rect 27734 10476 27792 10488
rect 28752 11064 28810 11076
rect 28752 10488 28764 11064
rect 28798 10488 28810 11064
rect 28752 10476 28810 10488
rect 29770 11064 29828 11076
rect 29770 10488 29782 11064
rect 29816 10488 29828 11064
rect 29770 10476 29828 10488
rect 30788 11064 30846 11076
rect 30788 10488 30800 11064
rect 30834 10488 30846 11064
rect 30788 10476 30846 10488
rect 31806 11064 31864 11076
rect 31806 10488 31818 11064
rect 31852 10488 31864 11064
rect 31806 10476 31864 10488
rect 32824 11064 32882 11076
rect 32824 10488 32836 11064
rect 32870 10488 32882 11064
rect 32824 10476 32882 10488
rect 33842 11064 33900 11076
rect 33842 10488 33854 11064
rect 33888 10488 33900 11064
rect 33842 10476 33900 10488
rect 10878 10156 10936 10168
rect 1716 9926 1774 9938
rect 1716 9350 1728 9926
rect 1762 9350 1774 9926
rect 1716 9338 1774 9350
rect 2734 9926 2792 9938
rect 2734 9350 2746 9926
rect 2780 9350 2792 9926
rect 2734 9338 2792 9350
rect 3752 9926 3810 9938
rect 3752 9350 3764 9926
rect 3798 9350 3810 9926
rect 3752 9338 3810 9350
rect 4770 9926 4828 9938
rect 4770 9350 4782 9926
rect 4816 9350 4828 9926
rect 4770 9338 4828 9350
rect 5788 9926 5846 9938
rect 5788 9350 5800 9926
rect 5834 9350 5846 9926
rect 5788 9338 5846 9350
rect 6806 9926 6864 9938
rect 6806 9350 6818 9926
rect 6852 9350 6864 9926
rect 6806 9338 6864 9350
rect 7824 9926 7882 9938
rect 7824 9350 7836 9926
rect 7870 9350 7882 9926
rect 7824 9338 7882 9350
rect 8842 9926 8900 9938
rect 8842 9350 8854 9926
rect 8888 9350 8900 9926
rect 8842 9338 8900 9350
rect 9860 9926 9918 9938
rect 9860 9350 9872 9926
rect 9906 9350 9918 9926
rect 9860 9338 9918 9350
rect 10878 9926 10936 9938
rect 10878 9350 10890 9926
rect 10924 9350 10936 9926
rect 10878 9338 10936 9350
rect 13480 9830 13538 9842
rect 13480 9254 13492 9830
rect 13526 9254 13538 9830
rect 13480 9242 13538 9254
rect 14498 9830 14556 9842
rect 14498 9254 14510 9830
rect 14544 9254 14556 9830
rect 14498 9242 14556 9254
rect 15516 9830 15574 9842
rect 15516 9254 15528 9830
rect 15562 9254 15574 9830
rect 15516 9242 15574 9254
rect 16534 9830 16592 9842
rect 16534 9254 16546 9830
rect 16580 9254 16592 9830
rect 16534 9242 16592 9254
rect 17552 9830 17610 9842
rect 17552 9254 17564 9830
rect 17598 9254 17610 9830
rect 17552 9242 17610 9254
rect 18570 9830 18628 9842
rect 18570 9254 18582 9830
rect 18616 9254 18628 9830
rect 18570 9242 18628 9254
rect 19588 9830 19646 9842
rect 19588 9254 19600 9830
rect 19634 9254 19646 9830
rect 19588 9242 19646 9254
rect 20606 9830 20664 9842
rect 20606 9254 20618 9830
rect 20652 9254 20664 9830
rect 20606 9242 20664 9254
rect 21624 9830 21682 9842
rect 21624 9254 21636 9830
rect 21670 9254 21682 9830
rect 21624 9242 21682 9254
rect 22642 9830 22700 9842
rect 22642 9254 22654 9830
rect 22688 9254 22700 9830
rect 22642 9242 22700 9254
rect 23660 9830 23718 9842
rect 23660 9254 23672 9830
rect 23706 9254 23718 9830
rect 23660 9242 23718 9254
rect 24678 9830 24736 9842
rect 24678 9254 24690 9830
rect 24724 9254 24736 9830
rect 24678 9242 24736 9254
rect 25696 9830 25754 9842
rect 25696 9254 25708 9830
rect 25742 9254 25754 9830
rect 25696 9242 25754 9254
rect 26714 9830 26772 9842
rect 26714 9254 26726 9830
rect 26760 9254 26772 9830
rect 26714 9242 26772 9254
rect 27732 9830 27790 9842
rect 27732 9254 27744 9830
rect 27778 9254 27790 9830
rect 27732 9242 27790 9254
rect 28750 9830 28808 9842
rect 28750 9254 28762 9830
rect 28796 9254 28808 9830
rect 28750 9242 28808 9254
rect 29768 9830 29826 9842
rect 29768 9254 29780 9830
rect 29814 9254 29826 9830
rect 29768 9242 29826 9254
rect 30786 9830 30844 9842
rect 30786 9254 30798 9830
rect 30832 9254 30844 9830
rect 30786 9242 30844 9254
rect 31804 9830 31862 9842
rect 31804 9254 31816 9830
rect 31850 9254 31862 9830
rect 31804 9242 31862 9254
rect 32822 9830 32880 9842
rect 32822 9254 32834 9830
rect 32868 9254 32880 9830
rect 32822 9242 32880 9254
rect 33840 9830 33898 9842
rect 33840 9254 33852 9830
rect 33886 9254 33898 9830
rect 33840 9242 33898 9254
rect 1716 9108 1774 9120
rect 1716 8532 1728 9108
rect 1762 8532 1774 9108
rect 1716 8520 1774 8532
rect 2734 9108 2792 9120
rect 2734 8532 2746 9108
rect 2780 8532 2792 9108
rect 2734 8520 2792 8532
rect 3752 9108 3810 9120
rect 3752 8532 3764 9108
rect 3798 8532 3810 9108
rect 3752 8520 3810 8532
rect 4770 9108 4828 9120
rect 4770 8532 4782 9108
rect 4816 8532 4828 9108
rect 4770 8520 4828 8532
rect 5788 9108 5846 9120
rect 5788 8532 5800 9108
rect 5834 8532 5846 9108
rect 5788 8520 5846 8532
rect 6806 9108 6864 9120
rect 6806 8532 6818 9108
rect 6852 8532 6864 9108
rect 6806 8520 6864 8532
rect 7824 9108 7882 9120
rect 7824 8532 7836 9108
rect 7870 8532 7882 9108
rect 7824 8520 7882 8532
rect 8842 9108 8900 9120
rect 8842 8532 8854 9108
rect 8888 8532 8900 9108
rect 8842 8520 8900 8532
rect 9860 9108 9918 9120
rect 9860 8532 9872 9108
rect 9906 8532 9918 9108
rect 9860 8520 9918 8532
rect 10878 9108 10936 9120
rect 10878 8532 10890 9108
rect 10924 8532 10936 9108
rect 10878 8520 10936 8532
rect 13480 8596 13538 8608
rect 1716 8290 1774 8302
rect 1716 7714 1728 8290
rect 1762 7714 1774 8290
rect 1716 7702 1774 7714
rect 2734 8290 2792 8302
rect 2734 7714 2746 8290
rect 2780 7714 2792 8290
rect 2734 7702 2792 7714
rect 3752 8290 3810 8302
rect 3752 7714 3764 8290
rect 3798 7714 3810 8290
rect 3752 7702 3810 7714
rect 4770 8290 4828 8302
rect 4770 7714 4782 8290
rect 4816 7714 4828 8290
rect 4770 7702 4828 7714
rect 5788 8290 5846 8302
rect 5788 7714 5800 8290
rect 5834 7714 5846 8290
rect 5788 7702 5846 7714
rect 6806 8290 6864 8302
rect 6806 7714 6818 8290
rect 6852 7714 6864 8290
rect 6806 7702 6864 7714
rect 7824 8290 7882 8302
rect 7824 7714 7836 8290
rect 7870 7714 7882 8290
rect 7824 7702 7882 7714
rect 8842 8290 8900 8302
rect 8842 7714 8854 8290
rect 8888 7714 8900 8290
rect 8842 7702 8900 7714
rect 9860 8290 9918 8302
rect 9860 7714 9872 8290
rect 9906 7714 9918 8290
rect 9860 7702 9918 7714
rect 10878 8290 10936 8302
rect 10878 7714 10890 8290
rect 10924 7714 10936 8290
rect 13480 8020 13492 8596
rect 13526 8020 13538 8596
rect 13480 8008 13538 8020
rect 14498 8596 14556 8608
rect 14498 8020 14510 8596
rect 14544 8020 14556 8596
rect 14498 8008 14556 8020
rect 15516 8596 15574 8608
rect 15516 8020 15528 8596
rect 15562 8020 15574 8596
rect 15516 8008 15574 8020
rect 16534 8596 16592 8608
rect 16534 8020 16546 8596
rect 16580 8020 16592 8596
rect 16534 8008 16592 8020
rect 17552 8596 17610 8608
rect 17552 8020 17564 8596
rect 17598 8020 17610 8596
rect 17552 8008 17610 8020
rect 18570 8596 18628 8608
rect 18570 8020 18582 8596
rect 18616 8020 18628 8596
rect 18570 8008 18628 8020
rect 19588 8596 19646 8608
rect 19588 8020 19600 8596
rect 19634 8020 19646 8596
rect 19588 8008 19646 8020
rect 20606 8596 20664 8608
rect 20606 8020 20618 8596
rect 20652 8020 20664 8596
rect 20606 8008 20664 8020
rect 21624 8596 21682 8608
rect 21624 8020 21636 8596
rect 21670 8020 21682 8596
rect 21624 8008 21682 8020
rect 22642 8596 22700 8608
rect 22642 8020 22654 8596
rect 22688 8020 22700 8596
rect 22642 8008 22700 8020
rect 23660 8596 23718 8608
rect 23660 8020 23672 8596
rect 23706 8020 23718 8596
rect 23660 8008 23718 8020
rect 24678 8596 24736 8608
rect 24678 8020 24690 8596
rect 24724 8020 24736 8596
rect 24678 8008 24736 8020
rect 25696 8596 25754 8608
rect 25696 8020 25708 8596
rect 25742 8020 25754 8596
rect 25696 8008 25754 8020
rect 26714 8596 26772 8608
rect 26714 8020 26726 8596
rect 26760 8020 26772 8596
rect 26714 8008 26772 8020
rect 27732 8596 27790 8608
rect 27732 8020 27744 8596
rect 27778 8020 27790 8596
rect 27732 8008 27790 8020
rect 28750 8596 28808 8608
rect 28750 8020 28762 8596
rect 28796 8020 28808 8596
rect 28750 8008 28808 8020
rect 29768 8596 29826 8608
rect 29768 8020 29780 8596
rect 29814 8020 29826 8596
rect 29768 8008 29826 8020
rect 30786 8596 30844 8608
rect 30786 8020 30798 8596
rect 30832 8020 30844 8596
rect 30786 8008 30844 8020
rect 31804 8596 31862 8608
rect 31804 8020 31816 8596
rect 31850 8020 31862 8596
rect 31804 8008 31862 8020
rect 32822 8596 32880 8608
rect 32822 8020 32834 8596
rect 32868 8020 32880 8596
rect 32822 8008 32880 8020
rect 33840 8596 33898 8608
rect 33840 8020 33852 8596
rect 33886 8020 33898 8596
rect 33840 8008 33898 8020
rect 10878 7702 10936 7714
rect 13480 7364 13538 7376
rect 13480 6788 13492 7364
rect 13526 6788 13538 7364
rect 13480 6776 13538 6788
rect 14498 7364 14556 7376
rect 14498 6788 14510 7364
rect 14544 6788 14556 7364
rect 14498 6776 14556 6788
rect 15516 7364 15574 7376
rect 15516 6788 15528 7364
rect 15562 6788 15574 7364
rect 15516 6776 15574 6788
rect 16534 7364 16592 7376
rect 16534 6788 16546 7364
rect 16580 6788 16592 7364
rect 16534 6776 16592 6788
rect 17552 7364 17610 7376
rect 17552 6788 17564 7364
rect 17598 6788 17610 7364
rect 17552 6776 17610 6788
rect 18570 7364 18628 7376
rect 18570 6788 18582 7364
rect 18616 6788 18628 7364
rect 18570 6776 18628 6788
rect 19588 7364 19646 7376
rect 19588 6788 19600 7364
rect 19634 6788 19646 7364
rect 19588 6776 19646 6788
rect 20606 7364 20664 7376
rect 20606 6788 20618 7364
rect 20652 6788 20664 7364
rect 20606 6776 20664 6788
rect 21624 7364 21682 7376
rect 21624 6788 21636 7364
rect 21670 6788 21682 7364
rect 21624 6776 21682 6788
rect 22642 7364 22700 7376
rect 22642 6788 22654 7364
rect 22688 6788 22700 7364
rect 22642 6776 22700 6788
rect 23660 7364 23718 7376
rect 23660 6788 23672 7364
rect 23706 6788 23718 7364
rect 23660 6776 23718 6788
rect 24678 7364 24736 7376
rect 24678 6788 24690 7364
rect 24724 6788 24736 7364
rect 24678 6776 24736 6788
rect 25696 7364 25754 7376
rect 25696 6788 25708 7364
rect 25742 6788 25754 7364
rect 25696 6776 25754 6788
rect 26714 7364 26772 7376
rect 26714 6788 26726 7364
rect 26760 6788 26772 7364
rect 26714 6776 26772 6788
rect 27732 7364 27790 7376
rect 27732 6788 27744 7364
rect 27778 6788 27790 7364
rect 27732 6776 27790 6788
rect 28750 7364 28808 7376
rect 28750 6788 28762 7364
rect 28796 6788 28808 7364
rect 28750 6776 28808 6788
rect 29768 7364 29826 7376
rect 29768 6788 29780 7364
rect 29814 6788 29826 7364
rect 29768 6776 29826 6788
rect 30786 7364 30844 7376
rect 30786 6788 30798 7364
rect 30832 6788 30844 7364
rect 30786 6776 30844 6788
rect 31804 7364 31862 7376
rect 31804 6788 31816 7364
rect 31850 6788 31862 7364
rect 31804 6776 31862 6788
rect 32822 7364 32880 7376
rect 32822 6788 32834 7364
rect 32868 6788 32880 7364
rect 32822 6776 32880 6788
rect 33840 7364 33898 7376
rect 33840 6788 33852 7364
rect 33886 6788 33898 7364
rect 33840 6776 33898 6788
rect 392 6266 450 6278
rect 392 5690 404 6266
rect 438 5690 450 6266
rect 392 5678 450 5690
rect 1410 6266 1468 6278
rect 1410 5690 1422 6266
rect 1456 5690 1468 6266
rect 1410 5678 1468 5690
rect 2428 6266 2486 6278
rect 2428 5690 2440 6266
rect 2474 5690 2486 6266
rect 2428 5678 2486 5690
rect 3446 6266 3504 6278
rect 3446 5690 3458 6266
rect 3492 5690 3504 6266
rect 3446 5678 3504 5690
rect 4464 6266 4522 6278
rect 4464 5690 4476 6266
rect 4510 5690 4522 6266
rect 4464 5678 4522 5690
rect 5482 6266 5540 6278
rect 5482 5690 5494 6266
rect 5528 5690 5540 6266
rect 5482 5678 5540 5690
rect 6500 6266 6558 6278
rect 6500 5690 6512 6266
rect 6546 5690 6558 6266
rect 6500 5678 6558 5690
rect 7518 6266 7576 6278
rect 7518 5690 7530 6266
rect 7564 5690 7576 6266
rect 7518 5678 7576 5690
rect 8536 6266 8594 6278
rect 8536 5690 8548 6266
rect 8582 5690 8594 6266
rect 8536 5678 8594 5690
rect 9554 6266 9612 6278
rect 9554 5690 9566 6266
rect 9600 5690 9612 6266
rect 9554 5678 9612 5690
rect 10572 6266 10630 6278
rect 10572 5690 10584 6266
rect 10618 5690 10630 6266
rect 10572 5678 10630 5690
rect 11590 6266 11648 6278
rect 11590 5690 11602 6266
rect 11636 5690 11648 6266
rect 11590 5678 11648 5690
rect 13480 6130 13538 6142
rect 13480 5554 13492 6130
rect 13526 5554 13538 6130
rect 13480 5542 13538 5554
rect 14498 6130 14556 6142
rect 14498 5554 14510 6130
rect 14544 5554 14556 6130
rect 14498 5542 14556 5554
rect 15516 6130 15574 6142
rect 15516 5554 15528 6130
rect 15562 5554 15574 6130
rect 15516 5542 15574 5554
rect 16534 6130 16592 6142
rect 16534 5554 16546 6130
rect 16580 5554 16592 6130
rect 16534 5542 16592 5554
rect 17552 6130 17610 6142
rect 17552 5554 17564 6130
rect 17598 5554 17610 6130
rect 17552 5542 17610 5554
rect 18570 6130 18628 6142
rect 18570 5554 18582 6130
rect 18616 5554 18628 6130
rect 18570 5542 18628 5554
rect 19588 6130 19646 6142
rect 19588 5554 19600 6130
rect 19634 5554 19646 6130
rect 19588 5542 19646 5554
rect 20606 6130 20664 6142
rect 20606 5554 20618 6130
rect 20652 5554 20664 6130
rect 20606 5542 20664 5554
rect 21624 6130 21682 6142
rect 21624 5554 21636 6130
rect 21670 5554 21682 6130
rect 21624 5542 21682 5554
rect 22642 6130 22700 6142
rect 22642 5554 22654 6130
rect 22688 5554 22700 6130
rect 22642 5542 22700 5554
rect 23660 6130 23718 6142
rect 23660 5554 23672 6130
rect 23706 5554 23718 6130
rect 23660 5542 23718 5554
rect 24678 6130 24736 6142
rect 24678 5554 24690 6130
rect 24724 5554 24736 6130
rect 24678 5542 24736 5554
rect 25696 6130 25754 6142
rect 25696 5554 25708 6130
rect 25742 5554 25754 6130
rect 25696 5542 25754 5554
rect 26714 6130 26772 6142
rect 26714 5554 26726 6130
rect 26760 5554 26772 6130
rect 26714 5542 26772 5554
rect 27732 6130 27790 6142
rect 27732 5554 27744 6130
rect 27778 5554 27790 6130
rect 27732 5542 27790 5554
rect 28750 6130 28808 6142
rect 28750 5554 28762 6130
rect 28796 5554 28808 6130
rect 28750 5542 28808 5554
rect 29768 6130 29826 6142
rect 29768 5554 29780 6130
rect 29814 5554 29826 6130
rect 29768 5542 29826 5554
rect 30786 6130 30844 6142
rect 30786 5554 30798 6130
rect 30832 5554 30844 6130
rect 30786 5542 30844 5554
rect 31804 6130 31862 6142
rect 31804 5554 31816 6130
rect 31850 5554 31862 6130
rect 31804 5542 31862 5554
rect 32822 6130 32880 6142
rect 32822 5554 32834 6130
rect 32868 5554 32880 6130
rect 32822 5542 32880 5554
rect 33840 6130 33898 6142
rect 33840 5554 33852 6130
rect 33886 5554 33898 6130
rect 33840 5542 33898 5554
rect 392 5154 450 5166
rect 392 4578 404 5154
rect 438 4578 450 5154
rect 392 4566 450 4578
rect 1410 5154 1468 5166
rect 1410 4578 1422 5154
rect 1456 4578 1468 5154
rect 1410 4566 1468 4578
rect 2428 5154 2486 5166
rect 2428 4578 2440 5154
rect 2474 4578 2486 5154
rect 2428 4566 2486 4578
rect 3446 5154 3504 5166
rect 3446 4578 3458 5154
rect 3492 4578 3504 5154
rect 3446 4566 3504 4578
rect 4464 5154 4522 5166
rect 4464 4578 4476 5154
rect 4510 4578 4522 5154
rect 4464 4566 4522 4578
rect 5482 5154 5540 5166
rect 5482 4578 5494 5154
rect 5528 4578 5540 5154
rect 5482 4566 5540 4578
rect 6500 5154 6558 5166
rect 6500 4578 6512 5154
rect 6546 4578 6558 5154
rect 6500 4566 6558 4578
rect 7518 5154 7576 5166
rect 7518 4578 7530 5154
rect 7564 4578 7576 5154
rect 7518 4566 7576 4578
rect 8536 5154 8594 5166
rect 8536 4578 8548 5154
rect 8582 4578 8594 5154
rect 8536 4566 8594 4578
rect 9554 5154 9612 5166
rect 9554 4578 9566 5154
rect 9600 4578 9612 5154
rect 9554 4566 9612 4578
rect 10572 5154 10630 5166
rect 10572 4578 10584 5154
rect 10618 4578 10630 5154
rect 10572 4566 10630 4578
rect 11590 5154 11648 5166
rect 11590 4578 11602 5154
rect 11636 4578 11648 5154
rect 11590 4566 11648 4578
rect 13480 4896 13538 4908
rect 13480 4320 13492 4896
rect 13526 4320 13538 4896
rect 13480 4308 13538 4320
rect 14498 4896 14556 4908
rect 14498 4320 14510 4896
rect 14544 4320 14556 4896
rect 14498 4308 14556 4320
rect 15516 4896 15574 4908
rect 15516 4320 15528 4896
rect 15562 4320 15574 4896
rect 15516 4308 15574 4320
rect 16534 4896 16592 4908
rect 16534 4320 16546 4896
rect 16580 4320 16592 4896
rect 16534 4308 16592 4320
rect 17552 4896 17610 4908
rect 17552 4320 17564 4896
rect 17598 4320 17610 4896
rect 17552 4308 17610 4320
rect 18570 4896 18628 4908
rect 18570 4320 18582 4896
rect 18616 4320 18628 4896
rect 18570 4308 18628 4320
rect 19588 4896 19646 4908
rect 19588 4320 19600 4896
rect 19634 4320 19646 4896
rect 19588 4308 19646 4320
rect 20606 4896 20664 4908
rect 20606 4320 20618 4896
rect 20652 4320 20664 4896
rect 20606 4308 20664 4320
rect 21624 4896 21682 4908
rect 21624 4320 21636 4896
rect 21670 4320 21682 4896
rect 21624 4308 21682 4320
rect 22642 4896 22700 4908
rect 22642 4320 22654 4896
rect 22688 4320 22700 4896
rect 22642 4308 22700 4320
rect 23660 4896 23718 4908
rect 23660 4320 23672 4896
rect 23706 4320 23718 4896
rect 23660 4308 23718 4320
rect 24678 4896 24736 4908
rect 24678 4320 24690 4896
rect 24724 4320 24736 4896
rect 24678 4308 24736 4320
rect 25696 4896 25754 4908
rect 25696 4320 25708 4896
rect 25742 4320 25754 4896
rect 25696 4308 25754 4320
rect 26714 4896 26772 4908
rect 26714 4320 26726 4896
rect 26760 4320 26772 4896
rect 26714 4308 26772 4320
rect 27732 4896 27790 4908
rect 27732 4320 27744 4896
rect 27778 4320 27790 4896
rect 27732 4308 27790 4320
rect 28750 4896 28808 4908
rect 28750 4320 28762 4896
rect 28796 4320 28808 4896
rect 28750 4308 28808 4320
rect 29768 4896 29826 4908
rect 29768 4320 29780 4896
rect 29814 4320 29826 4896
rect 29768 4308 29826 4320
rect 30786 4896 30844 4908
rect 30786 4320 30798 4896
rect 30832 4320 30844 4896
rect 30786 4308 30844 4320
rect 31804 4896 31862 4908
rect 31804 4320 31816 4896
rect 31850 4320 31862 4896
rect 31804 4308 31862 4320
rect 32822 4896 32880 4908
rect 32822 4320 32834 4896
rect 32868 4320 32880 4896
rect 32822 4308 32880 4320
rect 33840 4896 33898 4908
rect 33840 4320 33852 4896
rect 33886 4320 33898 4896
rect 33840 4308 33898 4320
rect 392 4042 450 4054
rect 392 3466 404 4042
rect 438 3466 450 4042
rect 392 3454 450 3466
rect 1410 4042 1468 4054
rect 1410 3466 1422 4042
rect 1456 3466 1468 4042
rect 1410 3454 1468 3466
rect 2428 4042 2486 4054
rect 2428 3466 2440 4042
rect 2474 3466 2486 4042
rect 2428 3454 2486 3466
rect 3446 4042 3504 4054
rect 3446 3466 3458 4042
rect 3492 3466 3504 4042
rect 3446 3454 3504 3466
rect 4464 4042 4522 4054
rect 4464 3466 4476 4042
rect 4510 3466 4522 4042
rect 4464 3454 4522 3466
rect 5482 4042 5540 4054
rect 5482 3466 5494 4042
rect 5528 3466 5540 4042
rect 5482 3454 5540 3466
rect 6500 4042 6558 4054
rect 6500 3466 6512 4042
rect 6546 3466 6558 4042
rect 6500 3454 6558 3466
rect 7518 4042 7576 4054
rect 7518 3466 7530 4042
rect 7564 3466 7576 4042
rect 7518 3454 7576 3466
rect 8536 4042 8594 4054
rect 8536 3466 8548 4042
rect 8582 3466 8594 4042
rect 8536 3454 8594 3466
rect 9554 4042 9612 4054
rect 9554 3466 9566 4042
rect 9600 3466 9612 4042
rect 9554 3454 9612 3466
rect 10572 4042 10630 4054
rect 10572 3466 10584 4042
rect 10618 3466 10630 4042
rect 10572 3454 10630 3466
rect 11590 4042 11648 4054
rect 11590 3466 11602 4042
rect 11636 3466 11648 4042
rect 11590 3454 11648 3466
rect 13480 3664 13538 3676
rect 13480 3088 13492 3664
rect 13526 3088 13538 3664
rect 13480 3076 13538 3088
rect 14498 3664 14556 3676
rect 14498 3088 14510 3664
rect 14544 3088 14556 3664
rect 14498 3076 14556 3088
rect 15516 3664 15574 3676
rect 15516 3088 15528 3664
rect 15562 3088 15574 3664
rect 15516 3076 15574 3088
rect 16534 3664 16592 3676
rect 16534 3088 16546 3664
rect 16580 3088 16592 3664
rect 16534 3076 16592 3088
rect 17552 3664 17610 3676
rect 17552 3088 17564 3664
rect 17598 3088 17610 3664
rect 17552 3076 17610 3088
rect 18570 3664 18628 3676
rect 18570 3088 18582 3664
rect 18616 3088 18628 3664
rect 18570 3076 18628 3088
rect 19588 3664 19646 3676
rect 19588 3088 19600 3664
rect 19634 3088 19646 3664
rect 19588 3076 19646 3088
rect 20606 3664 20664 3676
rect 20606 3088 20618 3664
rect 20652 3088 20664 3664
rect 20606 3076 20664 3088
rect 21624 3664 21682 3676
rect 21624 3088 21636 3664
rect 21670 3088 21682 3664
rect 21624 3076 21682 3088
rect 22642 3664 22700 3676
rect 22642 3088 22654 3664
rect 22688 3088 22700 3664
rect 22642 3076 22700 3088
rect 23660 3664 23718 3676
rect 23660 3088 23672 3664
rect 23706 3088 23718 3664
rect 23660 3076 23718 3088
rect 24678 3664 24736 3676
rect 24678 3088 24690 3664
rect 24724 3088 24736 3664
rect 24678 3076 24736 3088
rect 25696 3664 25754 3676
rect 25696 3088 25708 3664
rect 25742 3088 25754 3664
rect 25696 3076 25754 3088
rect 26714 3664 26772 3676
rect 26714 3088 26726 3664
rect 26760 3088 26772 3664
rect 26714 3076 26772 3088
rect 27732 3664 27790 3676
rect 27732 3088 27744 3664
rect 27778 3088 27790 3664
rect 27732 3076 27790 3088
rect 28750 3664 28808 3676
rect 28750 3088 28762 3664
rect 28796 3088 28808 3664
rect 28750 3076 28808 3088
rect 29768 3664 29826 3676
rect 29768 3088 29780 3664
rect 29814 3088 29826 3664
rect 29768 3076 29826 3088
rect 30786 3664 30844 3676
rect 30786 3088 30798 3664
rect 30832 3088 30844 3664
rect 30786 3076 30844 3088
rect 31804 3664 31862 3676
rect 31804 3088 31816 3664
rect 31850 3088 31862 3664
rect 31804 3076 31862 3088
rect 32822 3664 32880 3676
rect 32822 3088 32834 3664
rect 32868 3088 32880 3664
rect 32822 3076 32880 3088
rect 33840 3664 33898 3676
rect 33840 3088 33852 3664
rect 33886 3088 33898 3664
rect 33840 3076 33898 3088
rect 392 2930 450 2942
rect 392 2354 404 2930
rect 438 2354 450 2930
rect 392 2342 450 2354
rect 1410 2930 1468 2942
rect 1410 2354 1422 2930
rect 1456 2354 1468 2930
rect 1410 2342 1468 2354
rect 2428 2930 2486 2942
rect 2428 2354 2440 2930
rect 2474 2354 2486 2930
rect 2428 2342 2486 2354
rect 3446 2930 3504 2942
rect 3446 2354 3458 2930
rect 3492 2354 3504 2930
rect 3446 2342 3504 2354
rect 4464 2930 4522 2942
rect 4464 2354 4476 2930
rect 4510 2354 4522 2930
rect 4464 2342 4522 2354
rect 5482 2930 5540 2942
rect 5482 2354 5494 2930
rect 5528 2354 5540 2930
rect 5482 2342 5540 2354
rect 6500 2930 6558 2942
rect 6500 2354 6512 2930
rect 6546 2354 6558 2930
rect 6500 2342 6558 2354
rect 7518 2930 7576 2942
rect 7518 2354 7530 2930
rect 7564 2354 7576 2930
rect 7518 2342 7576 2354
rect 8536 2930 8594 2942
rect 8536 2354 8548 2930
rect 8582 2354 8594 2930
rect 8536 2342 8594 2354
rect 9554 2930 9612 2942
rect 9554 2354 9566 2930
rect 9600 2354 9612 2930
rect 9554 2342 9612 2354
rect 10572 2930 10630 2942
rect 10572 2354 10584 2930
rect 10618 2354 10630 2930
rect 10572 2342 10630 2354
rect 11590 2930 11648 2942
rect 11590 2354 11602 2930
rect 11636 2354 11648 2930
rect 11590 2342 11648 2354
rect 13480 2430 13538 2442
rect 13480 1854 13492 2430
rect 13526 1854 13538 2430
rect 13480 1842 13538 1854
rect 14498 2430 14556 2442
rect 14498 1854 14510 2430
rect 14544 1854 14556 2430
rect 14498 1842 14556 1854
rect 15516 2430 15574 2442
rect 15516 1854 15528 2430
rect 15562 1854 15574 2430
rect 15516 1842 15574 1854
rect 16534 2430 16592 2442
rect 16534 1854 16546 2430
rect 16580 1854 16592 2430
rect 16534 1842 16592 1854
rect 17552 2430 17610 2442
rect 17552 1854 17564 2430
rect 17598 1854 17610 2430
rect 17552 1842 17610 1854
rect 18570 2430 18628 2442
rect 18570 1854 18582 2430
rect 18616 1854 18628 2430
rect 18570 1842 18628 1854
rect 19588 2430 19646 2442
rect 19588 1854 19600 2430
rect 19634 1854 19646 2430
rect 19588 1842 19646 1854
rect 20606 2430 20664 2442
rect 20606 1854 20618 2430
rect 20652 1854 20664 2430
rect 20606 1842 20664 1854
rect 21624 2430 21682 2442
rect 21624 1854 21636 2430
rect 21670 1854 21682 2430
rect 21624 1842 21682 1854
rect 22642 2430 22700 2442
rect 22642 1854 22654 2430
rect 22688 1854 22700 2430
rect 22642 1842 22700 1854
rect 23660 2430 23718 2442
rect 23660 1854 23672 2430
rect 23706 1854 23718 2430
rect 23660 1842 23718 1854
rect 24678 2430 24736 2442
rect 24678 1854 24690 2430
rect 24724 1854 24736 2430
rect 24678 1842 24736 1854
rect 25696 2430 25754 2442
rect 25696 1854 25708 2430
rect 25742 1854 25754 2430
rect 25696 1842 25754 1854
rect 26714 2430 26772 2442
rect 26714 1854 26726 2430
rect 26760 1854 26772 2430
rect 26714 1842 26772 1854
rect 27732 2430 27790 2442
rect 27732 1854 27744 2430
rect 27778 1854 27790 2430
rect 27732 1842 27790 1854
rect 28750 2430 28808 2442
rect 28750 1854 28762 2430
rect 28796 1854 28808 2430
rect 28750 1842 28808 1854
rect 29768 2430 29826 2442
rect 29768 1854 29780 2430
rect 29814 1854 29826 2430
rect 29768 1842 29826 1854
rect 30786 2430 30844 2442
rect 30786 1854 30798 2430
rect 30832 1854 30844 2430
rect 30786 1842 30844 1854
rect 31804 2430 31862 2442
rect 31804 1854 31816 2430
rect 31850 1854 31862 2430
rect 31804 1842 31862 1854
rect 32822 2430 32880 2442
rect 32822 1854 32834 2430
rect 32868 1854 32880 2430
rect 32822 1842 32880 1854
rect 33840 2430 33898 2442
rect 33840 1854 33852 2430
rect 33886 1854 33898 2430
rect 33840 1842 33898 1854
rect 850 1388 908 1400
rect 850 812 862 1388
rect 896 812 908 1388
rect 850 800 908 812
rect 1868 1388 1926 1400
rect 1868 812 1880 1388
rect 1914 812 1926 1388
rect 1868 800 1926 812
rect 2886 1388 2944 1400
rect 2886 812 2898 1388
rect 2932 812 2944 1388
rect 2886 800 2944 812
rect 3904 1388 3962 1400
rect 3904 812 3916 1388
rect 3950 812 3962 1388
rect 3904 800 3962 812
rect 4922 1388 4980 1400
rect 4922 812 4934 1388
rect 4968 812 4980 1388
rect 4922 800 4980 812
rect 5940 1388 5998 1400
rect 5940 812 5952 1388
rect 5986 812 5998 1388
rect 5940 800 5998 812
rect 6958 1388 7016 1400
rect 6958 812 6970 1388
rect 7004 812 7016 1388
rect 6958 800 7016 812
rect 7976 1388 8034 1400
rect 7976 812 7988 1388
rect 8022 812 8034 1388
rect 7976 800 8034 812
rect 8994 1388 9052 1400
rect 8994 812 9006 1388
rect 9040 812 9052 1388
rect 8994 800 9052 812
rect 10012 1388 10070 1400
rect 10012 812 10024 1388
rect 10058 812 10070 1388
rect 10012 800 10070 812
rect 11030 1388 11088 1400
rect 11030 812 11042 1388
rect 11076 812 11088 1388
rect 11030 800 11088 812
rect 13480 1198 13538 1210
rect 13480 622 13492 1198
rect 13526 622 13538 1198
rect 13480 610 13538 622
rect 14498 1198 14556 1210
rect 14498 622 14510 1198
rect 14544 622 14556 1198
rect 14498 610 14556 622
rect 15516 1198 15574 1210
rect 15516 622 15528 1198
rect 15562 622 15574 1198
rect 15516 610 15574 622
rect 16534 1198 16592 1210
rect 16534 622 16546 1198
rect 16580 622 16592 1198
rect 16534 610 16592 622
rect 17552 1198 17610 1210
rect 17552 622 17564 1198
rect 17598 622 17610 1198
rect 17552 610 17610 622
rect 18570 1198 18628 1210
rect 18570 622 18582 1198
rect 18616 622 18628 1198
rect 18570 610 18628 622
rect 19588 1198 19646 1210
rect 19588 622 19600 1198
rect 19634 622 19646 1198
rect 19588 610 19646 622
rect 20606 1198 20664 1210
rect 20606 622 20618 1198
rect 20652 622 20664 1198
rect 20606 610 20664 622
rect 21624 1198 21682 1210
rect 21624 622 21636 1198
rect 21670 622 21682 1198
rect 21624 610 21682 622
rect 22642 1198 22700 1210
rect 22642 622 22654 1198
rect 22688 622 22700 1198
rect 22642 610 22700 622
rect 23660 1198 23718 1210
rect 23660 622 23672 1198
rect 23706 622 23718 1198
rect 23660 610 23718 622
rect 24678 1198 24736 1210
rect 24678 622 24690 1198
rect 24724 622 24736 1198
rect 24678 610 24736 622
rect 25696 1198 25754 1210
rect 25696 622 25708 1198
rect 25742 622 25754 1198
rect 25696 610 25754 622
rect 26714 1198 26772 1210
rect 26714 622 26726 1198
rect 26760 622 26772 1198
rect 26714 610 26772 622
rect 27732 1198 27790 1210
rect 27732 622 27744 1198
rect 27778 622 27790 1198
rect 27732 610 27790 622
rect 28750 1198 28808 1210
rect 28750 622 28762 1198
rect 28796 622 28808 1198
rect 28750 610 28808 622
rect 29768 1198 29826 1210
rect 29768 622 29780 1198
rect 29814 622 29826 1198
rect 29768 610 29826 622
rect 30786 1198 30844 1210
rect 30786 622 30798 1198
rect 30832 622 30844 1198
rect 30786 610 30844 622
rect 31804 1198 31862 1210
rect 31804 622 31816 1198
rect 31850 622 31862 1198
rect 31804 610 31862 622
rect 32822 1198 32880 1210
rect 32822 622 32834 1198
rect 32868 622 32880 1198
rect 32822 610 32880 622
rect 33840 1198 33898 1210
rect 33840 622 33852 1198
rect 33886 622 33898 1198
rect 33840 610 33898 622
<< pdiff >>
rect 17388 28002 17446 28014
rect 17388 27426 17400 28002
rect 17434 27426 17446 28002
rect 17388 27414 17446 27426
rect 18406 28002 18464 28014
rect 18406 27426 18418 28002
rect 18452 27426 18464 28002
rect 18406 27414 18464 27426
rect 19424 28002 19482 28014
rect 19424 27426 19436 28002
rect 19470 27426 19482 28002
rect 19424 27414 19482 27426
rect 20442 28002 20500 28014
rect 20442 27426 20454 28002
rect 20488 27426 20500 28002
rect 20442 27414 20500 27426
rect 21460 28002 21518 28014
rect 21460 27426 21472 28002
rect 21506 27426 21518 28002
rect 21460 27414 21518 27426
rect 22478 28002 22536 28014
rect 22478 27426 22490 28002
rect 22524 27426 22536 28002
rect 22478 27414 22536 27426
rect 23496 28002 23554 28014
rect 23496 27426 23508 28002
rect 23542 27426 23554 28002
rect 23496 27414 23554 27426
rect 24514 28002 24572 28014
rect 24514 27426 24526 28002
rect 24560 27426 24572 28002
rect 24514 27414 24572 27426
rect 25532 28002 25590 28014
rect 25532 27426 25544 28002
rect 25578 27426 25590 28002
rect 25532 27414 25590 27426
rect 26550 28002 26608 28014
rect 26550 27426 26562 28002
rect 26596 27426 26608 28002
rect 26550 27414 26608 27426
rect 27568 28002 27626 28014
rect 27568 27426 27580 28002
rect 27614 27426 27626 28002
rect 27568 27414 27626 27426
rect 28586 28002 28644 28014
rect 28586 27426 28598 28002
rect 28632 27426 28644 28002
rect 28586 27414 28644 27426
rect 29604 28002 29662 28014
rect 29604 27426 29616 28002
rect 29650 27426 29662 28002
rect 29604 27414 29662 27426
rect 30622 28002 30680 28014
rect 30622 27426 30634 28002
rect 30668 27426 30680 28002
rect 30622 27414 30680 27426
rect 31640 28002 31698 28014
rect 31640 27426 31652 28002
rect 31686 27426 31698 28002
rect 31640 27414 31698 27426
rect 32658 28002 32716 28014
rect 32658 27426 32670 28002
rect 32704 27426 32716 28002
rect 32658 27414 32716 27426
rect 33676 28002 33734 28014
rect 33676 27426 33688 28002
rect 33722 27426 33734 28002
rect 33676 27414 33734 27426
rect 17388 26866 17446 26878
rect 17388 26290 17400 26866
rect 17434 26290 17446 26866
rect 17388 26278 17446 26290
rect 18406 26866 18464 26878
rect 18406 26290 18418 26866
rect 18452 26290 18464 26866
rect 18406 26278 18464 26290
rect 19424 26866 19482 26878
rect 19424 26290 19436 26866
rect 19470 26290 19482 26866
rect 19424 26278 19482 26290
rect 20442 26866 20500 26878
rect 20442 26290 20454 26866
rect 20488 26290 20500 26866
rect 20442 26278 20500 26290
rect 21460 26866 21518 26878
rect 21460 26290 21472 26866
rect 21506 26290 21518 26866
rect 21460 26278 21518 26290
rect 22478 26866 22536 26878
rect 22478 26290 22490 26866
rect 22524 26290 22536 26866
rect 22478 26278 22536 26290
rect 23496 26866 23554 26878
rect 23496 26290 23508 26866
rect 23542 26290 23554 26866
rect 23496 26278 23554 26290
rect 24514 26866 24572 26878
rect 24514 26290 24526 26866
rect 24560 26290 24572 26866
rect 24514 26278 24572 26290
rect 25532 26866 25590 26878
rect 25532 26290 25544 26866
rect 25578 26290 25590 26866
rect 25532 26278 25590 26290
rect 26550 26866 26608 26878
rect 26550 26290 26562 26866
rect 26596 26290 26608 26866
rect 26550 26278 26608 26290
rect 27568 26866 27626 26878
rect 27568 26290 27580 26866
rect 27614 26290 27626 26866
rect 27568 26278 27626 26290
rect 28586 26866 28644 26878
rect 28586 26290 28598 26866
rect 28632 26290 28644 26866
rect 28586 26278 28644 26290
rect 29604 26866 29662 26878
rect 29604 26290 29616 26866
rect 29650 26290 29662 26866
rect 29604 26278 29662 26290
rect 30622 26866 30680 26878
rect 30622 26290 30634 26866
rect 30668 26290 30680 26866
rect 30622 26278 30680 26290
rect 31640 26866 31698 26878
rect 31640 26290 31652 26866
rect 31686 26290 31698 26866
rect 31640 26278 31698 26290
rect 32658 26866 32716 26878
rect 32658 26290 32670 26866
rect 32704 26290 32716 26866
rect 32658 26278 32716 26290
rect 33676 26866 33734 26878
rect 33676 26290 33688 26866
rect 33722 26290 33734 26866
rect 33676 26278 33734 26290
rect 17388 25730 17446 25742
rect 17388 25154 17400 25730
rect 17434 25154 17446 25730
rect 17388 25142 17446 25154
rect 18406 25730 18464 25742
rect 18406 25154 18418 25730
rect 18452 25154 18464 25730
rect 18406 25142 18464 25154
rect 19424 25730 19482 25742
rect 19424 25154 19436 25730
rect 19470 25154 19482 25730
rect 19424 25142 19482 25154
rect 20442 25730 20500 25742
rect 20442 25154 20454 25730
rect 20488 25154 20500 25730
rect 20442 25142 20500 25154
rect 21460 25730 21518 25742
rect 21460 25154 21472 25730
rect 21506 25154 21518 25730
rect 21460 25142 21518 25154
rect 22478 25730 22536 25742
rect 22478 25154 22490 25730
rect 22524 25154 22536 25730
rect 22478 25142 22536 25154
rect 23496 25730 23554 25742
rect 23496 25154 23508 25730
rect 23542 25154 23554 25730
rect 23496 25142 23554 25154
rect 24514 25730 24572 25742
rect 24514 25154 24526 25730
rect 24560 25154 24572 25730
rect 24514 25142 24572 25154
rect 25532 25730 25590 25742
rect 25532 25154 25544 25730
rect 25578 25154 25590 25730
rect 25532 25142 25590 25154
rect 26550 25730 26608 25742
rect 26550 25154 26562 25730
rect 26596 25154 26608 25730
rect 26550 25142 26608 25154
rect 27568 25730 27626 25742
rect 27568 25154 27580 25730
rect 27614 25154 27626 25730
rect 27568 25142 27626 25154
rect 28586 25730 28644 25742
rect 28586 25154 28598 25730
rect 28632 25154 28644 25730
rect 28586 25142 28644 25154
rect 29604 25730 29662 25742
rect 29604 25154 29616 25730
rect 29650 25154 29662 25730
rect 29604 25142 29662 25154
rect 30622 25730 30680 25742
rect 30622 25154 30634 25730
rect 30668 25154 30680 25730
rect 30622 25142 30680 25154
rect 31640 25730 31698 25742
rect 31640 25154 31652 25730
rect 31686 25154 31698 25730
rect 31640 25142 31698 25154
rect 32658 25730 32716 25742
rect 32658 25154 32670 25730
rect 32704 25154 32716 25730
rect 32658 25142 32716 25154
rect 33676 25730 33734 25742
rect 33676 25154 33688 25730
rect 33722 25154 33734 25730
rect 33676 25142 33734 25154
rect 18582 24092 18640 24104
rect 18582 23516 18594 24092
rect 18628 23516 18640 24092
rect 18582 23504 18640 23516
rect 19600 24092 19658 24104
rect 19600 23516 19612 24092
rect 19646 23516 19658 24092
rect 19600 23504 19658 23516
rect 20618 24092 20676 24104
rect 20618 23516 20630 24092
rect 20664 23516 20676 24092
rect 20618 23504 20676 23516
rect 21636 24092 21694 24104
rect 21636 23516 21648 24092
rect 21682 23516 21694 24092
rect 21636 23504 21694 23516
rect 22654 24092 22712 24104
rect 22654 23516 22666 24092
rect 22700 23516 22712 24092
rect 22654 23504 22712 23516
rect 23672 24092 23730 24104
rect 23672 23516 23684 24092
rect 23718 23516 23730 24092
rect 23672 23504 23730 23516
rect 24690 24092 24748 24104
rect 24690 23516 24702 24092
rect 24736 23516 24748 24092
rect 24690 23504 24748 23516
rect 25708 24092 25766 24104
rect 25708 23516 25720 24092
rect 25754 23516 25766 24092
rect 25708 23504 25766 23516
rect 26726 24092 26784 24104
rect 26726 23516 26738 24092
rect 26772 23516 26784 24092
rect 26726 23504 26784 23516
rect 27744 24092 27802 24104
rect 27744 23516 27756 24092
rect 27790 23516 27802 24092
rect 27744 23504 27802 23516
rect 28762 24092 28820 24104
rect 28762 23516 28774 24092
rect 28808 23516 28820 24092
rect 28762 23504 28820 23516
rect 29780 24092 29838 24104
rect 29780 23516 29792 24092
rect 29826 23516 29838 24092
rect 29780 23504 29838 23516
rect 30798 24092 30856 24104
rect 30798 23516 30810 24092
rect 30844 23516 30856 24092
rect 30798 23504 30856 23516
rect 31816 24092 31874 24104
rect 31816 23516 31828 24092
rect 31862 23516 31874 24092
rect 31816 23504 31874 23516
rect 32834 24092 32892 24104
rect 32834 23516 32846 24092
rect 32880 23516 32892 24092
rect 32834 23504 32892 23516
rect 18582 23060 18640 23072
rect 18582 22484 18594 23060
rect 18628 22484 18640 23060
rect 18582 22472 18640 22484
rect 19600 23060 19658 23072
rect 19600 22484 19612 23060
rect 19646 22484 19658 23060
rect 19600 22472 19658 22484
rect 20618 23060 20676 23072
rect 20618 22484 20630 23060
rect 20664 22484 20676 23060
rect 20618 22472 20676 22484
rect 21636 23060 21694 23072
rect 21636 22484 21648 23060
rect 21682 22484 21694 23060
rect 21636 22472 21694 22484
rect 22654 23060 22712 23072
rect 22654 22484 22666 23060
rect 22700 22484 22712 23060
rect 22654 22472 22712 22484
rect 23672 23060 23730 23072
rect 23672 22484 23684 23060
rect 23718 22484 23730 23060
rect 23672 22472 23730 22484
rect 24690 23060 24748 23072
rect 24690 22484 24702 23060
rect 24736 22484 24748 23060
rect 24690 22472 24748 22484
rect 25708 23060 25766 23072
rect 25708 22484 25720 23060
rect 25754 22484 25766 23060
rect 25708 22472 25766 22484
rect 26726 23060 26784 23072
rect 26726 22484 26738 23060
rect 26772 22484 26784 23060
rect 26726 22472 26784 22484
rect 27744 23060 27802 23072
rect 27744 22484 27756 23060
rect 27790 22484 27802 23060
rect 27744 22472 27802 22484
rect 28762 23060 28820 23072
rect 28762 22484 28774 23060
rect 28808 22484 28820 23060
rect 28762 22472 28820 22484
rect 29780 23060 29838 23072
rect 29780 22484 29792 23060
rect 29826 22484 29838 23060
rect 29780 22472 29838 22484
rect 30798 23060 30856 23072
rect 30798 22484 30810 23060
rect 30844 22484 30856 23060
rect 30798 22472 30856 22484
rect 31816 23060 31874 23072
rect 31816 22484 31828 23060
rect 31862 22484 31874 23060
rect 31816 22472 31874 22484
rect 32834 23060 32892 23072
rect 32834 22484 32846 23060
rect 32880 22484 32892 23060
rect 32834 22472 32892 22484
rect 18374 21456 18432 21468
rect 13070 21352 13128 21364
rect 13070 20776 13082 21352
rect 13116 20776 13128 21352
rect 13070 20764 13128 20776
rect 14088 21352 14146 21364
rect 14088 20776 14100 21352
rect 14134 20776 14146 21352
rect 14088 20764 14146 20776
rect 15106 21352 15164 21364
rect 15106 20776 15118 21352
rect 15152 20776 15164 21352
rect 15106 20764 15164 20776
rect 16124 21352 16182 21364
rect 16124 20776 16136 21352
rect 16170 20776 16182 21352
rect 16124 20764 16182 20776
rect 17142 21352 17200 21364
rect 17142 20776 17154 21352
rect 17188 20776 17200 21352
rect 18374 20880 18386 21456
rect 18420 20880 18432 21456
rect 18374 20868 18432 20880
rect 19392 21456 19450 21468
rect 19392 20880 19404 21456
rect 19438 20880 19450 21456
rect 19392 20868 19450 20880
rect 20410 21456 20468 21468
rect 20410 20880 20422 21456
rect 20456 20880 20468 21456
rect 20410 20868 20468 20880
rect 21428 21456 21486 21468
rect 21428 20880 21440 21456
rect 21474 20880 21486 21456
rect 21428 20868 21486 20880
rect 22446 21456 22504 21468
rect 22446 20880 22458 21456
rect 22492 20880 22504 21456
rect 22446 20868 22504 20880
rect 23464 21456 23522 21468
rect 23464 20880 23476 21456
rect 23510 20880 23522 21456
rect 23464 20868 23522 20880
rect 24482 21456 24540 21468
rect 24482 20880 24494 21456
rect 24528 20880 24540 21456
rect 24482 20868 24540 20880
rect 25500 21456 25558 21468
rect 25500 20880 25512 21456
rect 25546 20880 25558 21456
rect 25500 20868 25558 20880
rect 26518 21456 26576 21468
rect 26518 20880 26530 21456
rect 26564 20880 26576 21456
rect 26518 20868 26576 20880
rect 27536 21456 27594 21468
rect 27536 20880 27548 21456
rect 27582 20880 27594 21456
rect 27536 20868 27594 20880
rect 28554 21456 28612 21468
rect 28554 20880 28566 21456
rect 28600 20880 28612 21456
rect 28554 20868 28612 20880
rect 29572 21456 29630 21468
rect 29572 20880 29584 21456
rect 29618 20880 29630 21456
rect 29572 20868 29630 20880
rect 30590 21456 30648 21468
rect 30590 20880 30602 21456
rect 30636 20880 30648 21456
rect 30590 20868 30648 20880
rect 31608 21456 31666 21468
rect 31608 20880 31620 21456
rect 31654 20880 31666 21456
rect 31608 20868 31666 20880
rect 32626 21456 32684 21468
rect 32626 20880 32638 21456
rect 32672 20880 32684 21456
rect 32626 20868 32684 20880
rect 33644 21456 33702 21468
rect 33644 20880 33656 21456
rect 33690 20880 33702 21456
rect 33644 20868 33702 20880
rect 17142 20764 17200 20776
rect 13070 20320 13128 20332
rect 13070 19744 13082 20320
rect 13116 19744 13128 20320
rect 13070 19732 13128 19744
rect 14088 20320 14146 20332
rect 14088 19744 14100 20320
rect 14134 19744 14146 20320
rect 14088 19732 14146 19744
rect 15106 20320 15164 20332
rect 15106 19744 15118 20320
rect 15152 19744 15164 20320
rect 15106 19732 15164 19744
rect 16124 20320 16182 20332
rect 16124 19744 16136 20320
rect 16170 19744 16182 20320
rect 16124 19732 16182 19744
rect 17142 20320 17200 20332
rect 17142 19744 17154 20320
rect 17188 19744 17200 20320
rect 17142 19732 17200 19744
rect 18374 20200 18432 20212
rect 18374 19624 18386 20200
rect 18420 19624 18432 20200
rect 18374 19612 18432 19624
rect 19392 20200 19450 20212
rect 19392 19624 19404 20200
rect 19438 19624 19450 20200
rect 19392 19612 19450 19624
rect 20410 20200 20468 20212
rect 20410 19624 20422 20200
rect 20456 19624 20468 20200
rect 20410 19612 20468 19624
rect 21428 20200 21486 20212
rect 21428 19624 21440 20200
rect 21474 19624 21486 20200
rect 21428 19612 21486 19624
rect 22446 20200 22504 20212
rect 22446 19624 22458 20200
rect 22492 19624 22504 20200
rect 22446 19612 22504 19624
rect 23464 20200 23522 20212
rect 23464 19624 23476 20200
rect 23510 19624 23522 20200
rect 23464 19612 23522 19624
rect 24482 20200 24540 20212
rect 24482 19624 24494 20200
rect 24528 19624 24540 20200
rect 24482 19612 24540 19624
rect 25500 20200 25558 20212
rect 25500 19624 25512 20200
rect 25546 19624 25558 20200
rect 25500 19612 25558 19624
rect 26518 20200 26576 20212
rect 26518 19624 26530 20200
rect 26564 19624 26576 20200
rect 26518 19612 26576 19624
rect 27536 20200 27594 20212
rect 27536 19624 27548 20200
rect 27582 19624 27594 20200
rect 27536 19612 27594 19624
rect 28554 20200 28612 20212
rect 28554 19624 28566 20200
rect 28600 19624 28612 20200
rect 28554 19612 28612 19624
rect 29572 20200 29630 20212
rect 29572 19624 29584 20200
rect 29618 19624 29630 20200
rect 29572 19612 29630 19624
rect 30590 20200 30648 20212
rect 30590 19624 30602 20200
rect 30636 19624 30648 20200
rect 30590 19612 30648 19624
rect 31608 20200 31666 20212
rect 31608 19624 31620 20200
rect 31654 19624 31666 20200
rect 31608 19612 31666 19624
rect 32626 20200 32684 20212
rect 32626 19624 32638 20200
rect 32672 19624 32684 20200
rect 32626 19612 32684 19624
rect 33644 20200 33702 20212
rect 33644 19624 33656 20200
rect 33690 19624 33702 20200
rect 33644 19612 33702 19624
rect 13070 19288 13128 19300
rect 13070 18712 13082 19288
rect 13116 18712 13128 19288
rect 13070 18700 13128 18712
rect 14088 19288 14146 19300
rect 14088 18712 14100 19288
rect 14134 18712 14146 19288
rect 14088 18700 14146 18712
rect 15106 19288 15164 19300
rect 15106 18712 15118 19288
rect 15152 18712 15164 19288
rect 15106 18700 15164 18712
rect 16124 19288 16182 19300
rect 16124 18712 16136 19288
rect 16170 18712 16182 19288
rect 16124 18700 16182 18712
rect 17142 19288 17200 19300
rect 17142 18712 17154 19288
rect 17188 18712 17200 19288
rect 17142 18700 17200 18712
rect 18374 18944 18432 18956
rect 18374 18368 18386 18944
rect 18420 18368 18432 18944
rect 18374 18356 18432 18368
rect 19392 18944 19450 18956
rect 19392 18368 19404 18944
rect 19438 18368 19450 18944
rect 19392 18356 19450 18368
rect 20410 18944 20468 18956
rect 20410 18368 20422 18944
rect 20456 18368 20468 18944
rect 20410 18356 20468 18368
rect 21428 18944 21486 18956
rect 21428 18368 21440 18944
rect 21474 18368 21486 18944
rect 21428 18356 21486 18368
rect 22446 18944 22504 18956
rect 22446 18368 22458 18944
rect 22492 18368 22504 18944
rect 22446 18356 22504 18368
rect 23464 18944 23522 18956
rect 23464 18368 23476 18944
rect 23510 18368 23522 18944
rect 23464 18356 23522 18368
rect 24482 18944 24540 18956
rect 24482 18368 24494 18944
rect 24528 18368 24540 18944
rect 24482 18356 24540 18368
rect 25500 18944 25558 18956
rect 25500 18368 25512 18944
rect 25546 18368 25558 18944
rect 25500 18356 25558 18368
rect 26518 18944 26576 18956
rect 26518 18368 26530 18944
rect 26564 18368 26576 18944
rect 26518 18356 26576 18368
rect 27536 18944 27594 18956
rect 27536 18368 27548 18944
rect 27582 18368 27594 18944
rect 27536 18356 27594 18368
rect 28554 18944 28612 18956
rect 28554 18368 28566 18944
rect 28600 18368 28612 18944
rect 28554 18356 28612 18368
rect 29572 18944 29630 18956
rect 29572 18368 29584 18944
rect 29618 18368 29630 18944
rect 29572 18356 29630 18368
rect 30590 18944 30648 18956
rect 30590 18368 30602 18944
rect 30636 18368 30648 18944
rect 30590 18356 30648 18368
rect 31608 18944 31666 18956
rect 31608 18368 31620 18944
rect 31654 18368 31666 18944
rect 31608 18356 31666 18368
rect 32626 18944 32684 18956
rect 32626 18368 32638 18944
rect 32672 18368 32684 18944
rect 32626 18356 32684 18368
rect 33644 18944 33702 18956
rect 33644 18368 33656 18944
rect 33690 18368 33702 18944
rect 33644 18356 33702 18368
rect 13070 18256 13128 18268
rect 13070 17680 13082 18256
rect 13116 17680 13128 18256
rect 13070 17668 13128 17680
rect 14088 18256 14146 18268
rect 14088 17680 14100 18256
rect 14134 17680 14146 18256
rect 14088 17668 14146 17680
rect 15106 18256 15164 18268
rect 15106 17680 15118 18256
rect 15152 17680 15164 18256
rect 15106 17668 15164 17680
rect 16124 18256 16182 18268
rect 16124 17680 16136 18256
rect 16170 17680 16182 18256
rect 16124 17668 16182 17680
rect 17142 18256 17200 18268
rect 17142 17680 17154 18256
rect 17188 17680 17200 18256
rect 17142 17668 17200 17680
rect 18374 17688 18432 17700
rect 18374 17112 18386 17688
rect 18420 17112 18432 17688
rect 18374 17100 18432 17112
rect 19392 17688 19450 17700
rect 19392 17112 19404 17688
rect 19438 17112 19450 17688
rect 19392 17100 19450 17112
rect 20410 17688 20468 17700
rect 20410 17112 20422 17688
rect 20456 17112 20468 17688
rect 20410 17100 20468 17112
rect 21428 17688 21486 17700
rect 21428 17112 21440 17688
rect 21474 17112 21486 17688
rect 21428 17100 21486 17112
rect 22446 17688 22504 17700
rect 22446 17112 22458 17688
rect 22492 17112 22504 17688
rect 22446 17100 22504 17112
rect 23464 17688 23522 17700
rect 23464 17112 23476 17688
rect 23510 17112 23522 17688
rect 23464 17100 23522 17112
rect 24482 17688 24540 17700
rect 24482 17112 24494 17688
rect 24528 17112 24540 17688
rect 24482 17100 24540 17112
rect 25500 17688 25558 17700
rect 25500 17112 25512 17688
rect 25546 17112 25558 17688
rect 25500 17100 25558 17112
rect 26518 17688 26576 17700
rect 26518 17112 26530 17688
rect 26564 17112 26576 17688
rect 26518 17100 26576 17112
rect 27536 17688 27594 17700
rect 27536 17112 27548 17688
rect 27582 17112 27594 17688
rect 27536 17100 27594 17112
rect 28554 17688 28612 17700
rect 28554 17112 28566 17688
rect 28600 17112 28612 17688
rect 28554 17100 28612 17112
rect 29572 17688 29630 17700
rect 29572 17112 29584 17688
rect 29618 17112 29630 17688
rect 29572 17100 29630 17112
rect 30590 17688 30648 17700
rect 30590 17112 30602 17688
rect 30636 17112 30648 17688
rect 30590 17100 30648 17112
rect 31608 17688 31666 17700
rect 31608 17112 31620 17688
rect 31654 17112 31666 17688
rect 31608 17100 31666 17112
rect 32626 17688 32684 17700
rect 32626 17112 32638 17688
rect 32672 17112 32684 17688
rect 32626 17100 32684 17112
rect 33644 17688 33702 17700
rect 33644 17112 33656 17688
rect 33690 17112 33702 17688
rect 33644 17100 33702 17112
rect -12178 16114 -12120 16126
rect -12178 15738 -12166 16114
rect -12132 15738 -12120 16114
rect -12178 15726 -12120 15738
rect -11920 16114 -11862 16126
rect -11920 15738 -11908 16114
rect -11874 15738 -11862 16114
rect -11920 15726 -11862 15738
rect -11662 16114 -11604 16126
rect -11662 15738 -11650 16114
rect -11616 15738 -11604 16114
rect -11662 15726 -11604 15738
rect -11404 16114 -11346 16126
rect -11404 15738 -11392 16114
rect -11358 15738 -11346 16114
rect -11404 15726 -11346 15738
rect -11146 16114 -11088 16126
rect -11146 15738 -11134 16114
rect -11100 15738 -11088 16114
rect -11146 15726 -11088 15738
rect -10888 16114 -10830 16126
rect -10888 15738 -10876 16114
rect -10842 15738 -10830 16114
rect -10888 15726 -10830 15738
rect -10630 16114 -10572 16126
rect -10630 15738 -10618 16114
rect -10584 15738 -10572 16114
rect -10630 15726 -10572 15738
rect -10322 15731 -10270 15743
rect -10322 15697 -10314 15731
rect -10280 15697 -10270 15731
rect -10322 15663 -10270 15697
rect -10322 15629 -10314 15663
rect -10280 15629 -10270 15663
rect -10322 15595 -10270 15629
rect -10322 15561 -10314 15595
rect -10280 15561 -10270 15595
rect -10322 15543 -10270 15561
rect -10240 15731 -10188 15743
rect -10240 15697 -10230 15731
rect -10196 15697 -10188 15731
rect -10240 15663 -10188 15697
rect -10240 15629 -10230 15663
rect -10196 15629 -10188 15663
rect -10240 15595 -10188 15629
rect -10240 15561 -10230 15595
rect -10196 15561 -10188 15595
rect -10240 15543 -10188 15561
rect -9578 16114 -9520 16126
rect -9578 15738 -9566 16114
rect -9532 15738 -9520 16114
rect -9578 15726 -9520 15738
rect -9320 16114 -9262 16126
rect -9320 15738 -9308 16114
rect -9274 15738 -9262 16114
rect -9320 15726 -9262 15738
rect -9062 16114 -9004 16126
rect -9062 15738 -9050 16114
rect -9016 15738 -9004 16114
rect -9062 15726 -9004 15738
rect -8804 16114 -8746 16126
rect -8804 15738 -8792 16114
rect -8758 15738 -8746 16114
rect -8804 15726 -8746 15738
rect -8546 16114 -8488 16126
rect -8546 15738 -8534 16114
rect -8500 15738 -8488 16114
rect -8546 15726 -8488 15738
rect -8288 16114 -8230 16126
rect -8288 15738 -8276 16114
rect -8242 15738 -8230 16114
rect -8288 15726 -8230 15738
rect -8030 16114 -7972 16126
rect -8030 15738 -8018 16114
rect -7984 15738 -7972 16114
rect -8030 15726 -7972 15738
rect -7722 15731 -7670 15743
rect -7722 15697 -7714 15731
rect -7680 15697 -7670 15731
rect -7722 15663 -7670 15697
rect -7722 15629 -7714 15663
rect -7680 15629 -7670 15663
rect -7722 15595 -7670 15629
rect -7722 15561 -7714 15595
rect -7680 15561 -7670 15595
rect -7722 15543 -7670 15561
rect -7640 15731 -7588 15743
rect -7640 15697 -7630 15731
rect -7596 15697 -7588 15731
rect -7640 15663 -7588 15697
rect -7640 15629 -7630 15663
rect -7596 15629 -7588 15663
rect -7640 15595 -7588 15629
rect -7640 15561 -7630 15595
rect -7596 15561 -7588 15595
rect -7640 15543 -7588 15561
rect -7272 15731 -7220 15743
rect -7272 15697 -7264 15731
rect -7230 15697 -7220 15731
rect -7272 15663 -7220 15697
rect -7272 15629 -7264 15663
rect -7230 15629 -7220 15663
rect -7272 15595 -7220 15629
rect -7272 15561 -7264 15595
rect -7230 15561 -7220 15595
rect -7272 15543 -7220 15561
rect -7190 15731 -7138 15743
rect -7190 15697 -7180 15731
rect -7146 15697 -7138 15731
rect -7190 15663 -7138 15697
rect -7190 15629 -7180 15663
rect -7146 15629 -7138 15663
rect -7190 15595 -7138 15629
rect -7190 15561 -7180 15595
rect -7146 15561 -7138 15595
rect -7190 15543 -7138 15561
<< ndiffc >>
rect -10314 15377 -10280 15411
rect -10314 15309 -10280 15343
rect -10230 15377 -10196 15411
rect -7714 15377 -7680 15411
rect -10230 15309 -10196 15343
rect -12166 15014 -12132 15190
rect -11908 15014 -11874 15190
rect -11650 15014 -11616 15190
rect -11392 15014 -11358 15190
rect -11134 15014 -11100 15190
rect -10876 15014 -10842 15190
rect -10618 15014 -10584 15190
rect -7714 15309 -7680 15343
rect -7630 15377 -7596 15411
rect -7630 15309 -7596 15343
rect -7264 15377 -7230 15411
rect -7264 15309 -7230 15343
rect -7180 15377 -7146 15411
rect -7180 15309 -7146 15343
rect -9566 15014 -9532 15190
rect -9308 15014 -9274 15190
rect -9050 15014 -9016 15190
rect -8792 15014 -8758 15190
rect -8534 15014 -8500 15190
rect -8276 15014 -8242 15190
rect -8018 15014 -7984 15190
rect 1728 13440 1762 14016
rect 2746 13440 2780 14016
rect 3764 13440 3798 14016
rect 4782 13440 4816 14016
rect 5800 13440 5834 14016
rect 6818 13440 6852 14016
rect 7836 13440 7870 14016
rect 8854 13440 8888 14016
rect 9872 13440 9906 14016
rect 10890 13440 10924 14016
rect 13494 13916 13528 14492
rect 14512 13916 14546 14492
rect 15530 13916 15564 14492
rect 16548 13916 16582 14492
rect 17566 13916 17600 14492
rect 18584 13916 18618 14492
rect 19602 13916 19636 14492
rect 20620 13916 20654 14492
rect 21638 13916 21672 14492
rect 22656 13916 22690 14492
rect 23674 13916 23708 14492
rect 24692 13916 24726 14492
rect 25710 13916 25744 14492
rect 26728 13916 26762 14492
rect 27746 13916 27780 14492
rect 28764 13916 28798 14492
rect 29782 13916 29816 14492
rect 30800 13916 30834 14492
rect 31818 13916 31852 14492
rect 32836 13916 32870 14492
rect 33854 13916 33888 14492
rect 1728 12622 1762 13198
rect 2746 12622 2780 13198
rect 3764 12622 3798 13198
rect 4782 12622 4816 13198
rect 5800 12622 5834 13198
rect 6818 12622 6852 13198
rect 7836 12622 7870 13198
rect 8854 12622 8888 13198
rect 9872 12622 9906 13198
rect 10890 12622 10924 13198
rect 13494 13098 13528 13674
rect 14512 13098 14546 13674
rect 15530 13098 15564 13674
rect 16548 13098 16582 13674
rect 17566 13098 17600 13674
rect 18584 13098 18618 13674
rect 19602 13098 19636 13674
rect 20620 13098 20654 13674
rect 21638 13098 21672 13674
rect 22656 13098 22690 13674
rect 23674 13098 23708 13674
rect 24692 13098 24726 13674
rect 25710 13098 25744 13674
rect 26728 13098 26762 13674
rect 27746 13098 27780 13674
rect 28764 13098 28798 13674
rect 29782 13098 29816 13674
rect 30800 13098 30834 13674
rect 31818 13098 31852 13674
rect 32836 13098 32870 13674
rect 33854 13098 33888 13674
rect 1728 11804 1762 12380
rect 2746 11804 2780 12380
rect 3764 11804 3798 12380
rect 4782 11804 4816 12380
rect 5800 11804 5834 12380
rect 6818 11804 6852 12380
rect 7836 11804 7870 12380
rect 8854 11804 8888 12380
rect 9872 11804 9906 12380
rect 10890 11804 10924 12380
rect 13494 11720 13528 12296
rect 14512 11720 14546 12296
rect 15530 11720 15564 12296
rect 16548 11720 16582 12296
rect 17566 11720 17600 12296
rect 18584 11720 18618 12296
rect 19602 11720 19636 12296
rect 20620 11720 20654 12296
rect 21638 11720 21672 12296
rect 22656 11720 22690 12296
rect 23674 11720 23708 12296
rect 24692 11720 24726 12296
rect 25710 11720 25744 12296
rect 26728 11720 26762 12296
rect 27746 11720 27780 12296
rect 28764 11720 28798 12296
rect 29782 11720 29816 12296
rect 30800 11720 30834 12296
rect 31818 11720 31852 12296
rect 32836 11720 32870 12296
rect 33854 11720 33888 12296
rect 1728 10986 1762 11562
rect 2746 10986 2780 11562
rect 3764 10986 3798 11562
rect 4782 10986 4816 11562
rect 5800 10986 5834 11562
rect 6818 10986 6852 11562
rect 7836 10986 7870 11562
rect 8854 10986 8888 11562
rect 9872 10986 9906 11562
rect 10890 10986 10924 11562
rect 1728 10168 1762 10744
rect 2746 10168 2780 10744
rect 3764 10168 3798 10744
rect 4782 10168 4816 10744
rect 5800 10168 5834 10744
rect 6818 10168 6852 10744
rect 7836 10168 7870 10744
rect 8854 10168 8888 10744
rect 9872 10168 9906 10744
rect 10890 10168 10924 10744
rect 13494 10488 13528 11064
rect 14512 10488 14546 11064
rect 15530 10488 15564 11064
rect 16548 10488 16582 11064
rect 17566 10488 17600 11064
rect 18584 10488 18618 11064
rect 19602 10488 19636 11064
rect 20620 10488 20654 11064
rect 21638 10488 21672 11064
rect 22656 10488 22690 11064
rect 23674 10488 23708 11064
rect 24692 10488 24726 11064
rect 25710 10488 25744 11064
rect 26728 10488 26762 11064
rect 27746 10488 27780 11064
rect 28764 10488 28798 11064
rect 29782 10488 29816 11064
rect 30800 10488 30834 11064
rect 31818 10488 31852 11064
rect 32836 10488 32870 11064
rect 33854 10488 33888 11064
rect 1728 9350 1762 9926
rect 2746 9350 2780 9926
rect 3764 9350 3798 9926
rect 4782 9350 4816 9926
rect 5800 9350 5834 9926
rect 6818 9350 6852 9926
rect 7836 9350 7870 9926
rect 8854 9350 8888 9926
rect 9872 9350 9906 9926
rect 10890 9350 10924 9926
rect 13492 9254 13526 9830
rect 14510 9254 14544 9830
rect 15528 9254 15562 9830
rect 16546 9254 16580 9830
rect 17564 9254 17598 9830
rect 18582 9254 18616 9830
rect 19600 9254 19634 9830
rect 20618 9254 20652 9830
rect 21636 9254 21670 9830
rect 22654 9254 22688 9830
rect 23672 9254 23706 9830
rect 24690 9254 24724 9830
rect 25708 9254 25742 9830
rect 26726 9254 26760 9830
rect 27744 9254 27778 9830
rect 28762 9254 28796 9830
rect 29780 9254 29814 9830
rect 30798 9254 30832 9830
rect 31816 9254 31850 9830
rect 32834 9254 32868 9830
rect 33852 9254 33886 9830
rect 1728 8532 1762 9108
rect 2746 8532 2780 9108
rect 3764 8532 3798 9108
rect 4782 8532 4816 9108
rect 5800 8532 5834 9108
rect 6818 8532 6852 9108
rect 7836 8532 7870 9108
rect 8854 8532 8888 9108
rect 9872 8532 9906 9108
rect 10890 8532 10924 9108
rect 1728 7714 1762 8290
rect 2746 7714 2780 8290
rect 3764 7714 3798 8290
rect 4782 7714 4816 8290
rect 5800 7714 5834 8290
rect 6818 7714 6852 8290
rect 7836 7714 7870 8290
rect 8854 7714 8888 8290
rect 9872 7714 9906 8290
rect 10890 7714 10924 8290
rect 13492 8020 13526 8596
rect 14510 8020 14544 8596
rect 15528 8020 15562 8596
rect 16546 8020 16580 8596
rect 17564 8020 17598 8596
rect 18582 8020 18616 8596
rect 19600 8020 19634 8596
rect 20618 8020 20652 8596
rect 21636 8020 21670 8596
rect 22654 8020 22688 8596
rect 23672 8020 23706 8596
rect 24690 8020 24724 8596
rect 25708 8020 25742 8596
rect 26726 8020 26760 8596
rect 27744 8020 27778 8596
rect 28762 8020 28796 8596
rect 29780 8020 29814 8596
rect 30798 8020 30832 8596
rect 31816 8020 31850 8596
rect 32834 8020 32868 8596
rect 33852 8020 33886 8596
rect 13492 6788 13526 7364
rect 14510 6788 14544 7364
rect 15528 6788 15562 7364
rect 16546 6788 16580 7364
rect 17564 6788 17598 7364
rect 18582 6788 18616 7364
rect 19600 6788 19634 7364
rect 20618 6788 20652 7364
rect 21636 6788 21670 7364
rect 22654 6788 22688 7364
rect 23672 6788 23706 7364
rect 24690 6788 24724 7364
rect 25708 6788 25742 7364
rect 26726 6788 26760 7364
rect 27744 6788 27778 7364
rect 28762 6788 28796 7364
rect 29780 6788 29814 7364
rect 30798 6788 30832 7364
rect 31816 6788 31850 7364
rect 32834 6788 32868 7364
rect 33852 6788 33886 7364
rect 404 5690 438 6266
rect 1422 5690 1456 6266
rect 2440 5690 2474 6266
rect 3458 5690 3492 6266
rect 4476 5690 4510 6266
rect 5494 5690 5528 6266
rect 6512 5690 6546 6266
rect 7530 5690 7564 6266
rect 8548 5690 8582 6266
rect 9566 5690 9600 6266
rect 10584 5690 10618 6266
rect 11602 5690 11636 6266
rect 13492 5554 13526 6130
rect 14510 5554 14544 6130
rect 15528 5554 15562 6130
rect 16546 5554 16580 6130
rect 17564 5554 17598 6130
rect 18582 5554 18616 6130
rect 19600 5554 19634 6130
rect 20618 5554 20652 6130
rect 21636 5554 21670 6130
rect 22654 5554 22688 6130
rect 23672 5554 23706 6130
rect 24690 5554 24724 6130
rect 25708 5554 25742 6130
rect 26726 5554 26760 6130
rect 27744 5554 27778 6130
rect 28762 5554 28796 6130
rect 29780 5554 29814 6130
rect 30798 5554 30832 6130
rect 31816 5554 31850 6130
rect 32834 5554 32868 6130
rect 33852 5554 33886 6130
rect 404 4578 438 5154
rect 1422 4578 1456 5154
rect 2440 4578 2474 5154
rect 3458 4578 3492 5154
rect 4476 4578 4510 5154
rect 5494 4578 5528 5154
rect 6512 4578 6546 5154
rect 7530 4578 7564 5154
rect 8548 4578 8582 5154
rect 9566 4578 9600 5154
rect 10584 4578 10618 5154
rect 11602 4578 11636 5154
rect 13492 4320 13526 4896
rect 14510 4320 14544 4896
rect 15528 4320 15562 4896
rect 16546 4320 16580 4896
rect 17564 4320 17598 4896
rect 18582 4320 18616 4896
rect 19600 4320 19634 4896
rect 20618 4320 20652 4896
rect 21636 4320 21670 4896
rect 22654 4320 22688 4896
rect 23672 4320 23706 4896
rect 24690 4320 24724 4896
rect 25708 4320 25742 4896
rect 26726 4320 26760 4896
rect 27744 4320 27778 4896
rect 28762 4320 28796 4896
rect 29780 4320 29814 4896
rect 30798 4320 30832 4896
rect 31816 4320 31850 4896
rect 32834 4320 32868 4896
rect 33852 4320 33886 4896
rect 404 3466 438 4042
rect 1422 3466 1456 4042
rect 2440 3466 2474 4042
rect 3458 3466 3492 4042
rect 4476 3466 4510 4042
rect 5494 3466 5528 4042
rect 6512 3466 6546 4042
rect 7530 3466 7564 4042
rect 8548 3466 8582 4042
rect 9566 3466 9600 4042
rect 10584 3466 10618 4042
rect 11602 3466 11636 4042
rect 13492 3088 13526 3664
rect 14510 3088 14544 3664
rect 15528 3088 15562 3664
rect 16546 3088 16580 3664
rect 17564 3088 17598 3664
rect 18582 3088 18616 3664
rect 19600 3088 19634 3664
rect 20618 3088 20652 3664
rect 21636 3088 21670 3664
rect 22654 3088 22688 3664
rect 23672 3088 23706 3664
rect 24690 3088 24724 3664
rect 25708 3088 25742 3664
rect 26726 3088 26760 3664
rect 27744 3088 27778 3664
rect 28762 3088 28796 3664
rect 29780 3088 29814 3664
rect 30798 3088 30832 3664
rect 31816 3088 31850 3664
rect 32834 3088 32868 3664
rect 33852 3088 33886 3664
rect 404 2354 438 2930
rect 1422 2354 1456 2930
rect 2440 2354 2474 2930
rect 3458 2354 3492 2930
rect 4476 2354 4510 2930
rect 5494 2354 5528 2930
rect 6512 2354 6546 2930
rect 7530 2354 7564 2930
rect 8548 2354 8582 2930
rect 9566 2354 9600 2930
rect 10584 2354 10618 2930
rect 11602 2354 11636 2930
rect 13492 1854 13526 2430
rect 14510 1854 14544 2430
rect 15528 1854 15562 2430
rect 16546 1854 16580 2430
rect 17564 1854 17598 2430
rect 18582 1854 18616 2430
rect 19600 1854 19634 2430
rect 20618 1854 20652 2430
rect 21636 1854 21670 2430
rect 22654 1854 22688 2430
rect 23672 1854 23706 2430
rect 24690 1854 24724 2430
rect 25708 1854 25742 2430
rect 26726 1854 26760 2430
rect 27744 1854 27778 2430
rect 28762 1854 28796 2430
rect 29780 1854 29814 2430
rect 30798 1854 30832 2430
rect 31816 1854 31850 2430
rect 32834 1854 32868 2430
rect 33852 1854 33886 2430
rect 862 812 896 1388
rect 1880 812 1914 1388
rect 2898 812 2932 1388
rect 3916 812 3950 1388
rect 4934 812 4968 1388
rect 5952 812 5986 1388
rect 6970 812 7004 1388
rect 7988 812 8022 1388
rect 9006 812 9040 1388
rect 10024 812 10058 1388
rect 11042 812 11076 1388
rect 13492 622 13526 1198
rect 14510 622 14544 1198
rect 15528 622 15562 1198
rect 16546 622 16580 1198
rect 17564 622 17598 1198
rect 18582 622 18616 1198
rect 19600 622 19634 1198
rect 20618 622 20652 1198
rect 21636 622 21670 1198
rect 22654 622 22688 1198
rect 23672 622 23706 1198
rect 24690 622 24724 1198
rect 25708 622 25742 1198
rect 26726 622 26760 1198
rect 27744 622 27778 1198
rect 28762 622 28796 1198
rect 29780 622 29814 1198
rect 30798 622 30832 1198
rect 31816 622 31850 1198
rect 32834 622 32868 1198
rect 33852 622 33886 1198
<< pdiffc >>
rect 17400 27426 17434 28002
rect 18418 27426 18452 28002
rect 19436 27426 19470 28002
rect 20454 27426 20488 28002
rect 21472 27426 21506 28002
rect 22490 27426 22524 28002
rect 23508 27426 23542 28002
rect 24526 27426 24560 28002
rect 25544 27426 25578 28002
rect 26562 27426 26596 28002
rect 27580 27426 27614 28002
rect 28598 27426 28632 28002
rect 29616 27426 29650 28002
rect 30634 27426 30668 28002
rect 31652 27426 31686 28002
rect 32670 27426 32704 28002
rect 33688 27426 33722 28002
rect 17400 26290 17434 26866
rect 18418 26290 18452 26866
rect 19436 26290 19470 26866
rect 20454 26290 20488 26866
rect 21472 26290 21506 26866
rect 22490 26290 22524 26866
rect 23508 26290 23542 26866
rect 24526 26290 24560 26866
rect 25544 26290 25578 26866
rect 26562 26290 26596 26866
rect 27580 26290 27614 26866
rect 28598 26290 28632 26866
rect 29616 26290 29650 26866
rect 30634 26290 30668 26866
rect 31652 26290 31686 26866
rect 32670 26290 32704 26866
rect 33688 26290 33722 26866
rect 17400 25154 17434 25730
rect 18418 25154 18452 25730
rect 19436 25154 19470 25730
rect 20454 25154 20488 25730
rect 21472 25154 21506 25730
rect 22490 25154 22524 25730
rect 23508 25154 23542 25730
rect 24526 25154 24560 25730
rect 25544 25154 25578 25730
rect 26562 25154 26596 25730
rect 27580 25154 27614 25730
rect 28598 25154 28632 25730
rect 29616 25154 29650 25730
rect 30634 25154 30668 25730
rect 31652 25154 31686 25730
rect 32670 25154 32704 25730
rect 33688 25154 33722 25730
rect 18594 23516 18628 24092
rect 19612 23516 19646 24092
rect 20630 23516 20664 24092
rect 21648 23516 21682 24092
rect 22666 23516 22700 24092
rect 23684 23516 23718 24092
rect 24702 23516 24736 24092
rect 25720 23516 25754 24092
rect 26738 23516 26772 24092
rect 27756 23516 27790 24092
rect 28774 23516 28808 24092
rect 29792 23516 29826 24092
rect 30810 23516 30844 24092
rect 31828 23516 31862 24092
rect 32846 23516 32880 24092
rect 18594 22484 18628 23060
rect 19612 22484 19646 23060
rect 20630 22484 20664 23060
rect 21648 22484 21682 23060
rect 22666 22484 22700 23060
rect 23684 22484 23718 23060
rect 24702 22484 24736 23060
rect 25720 22484 25754 23060
rect 26738 22484 26772 23060
rect 27756 22484 27790 23060
rect 28774 22484 28808 23060
rect 29792 22484 29826 23060
rect 30810 22484 30844 23060
rect 31828 22484 31862 23060
rect 32846 22484 32880 23060
rect 13082 20776 13116 21352
rect 14100 20776 14134 21352
rect 15118 20776 15152 21352
rect 16136 20776 16170 21352
rect 17154 20776 17188 21352
rect 18386 20880 18420 21456
rect 19404 20880 19438 21456
rect 20422 20880 20456 21456
rect 21440 20880 21474 21456
rect 22458 20880 22492 21456
rect 23476 20880 23510 21456
rect 24494 20880 24528 21456
rect 25512 20880 25546 21456
rect 26530 20880 26564 21456
rect 27548 20880 27582 21456
rect 28566 20880 28600 21456
rect 29584 20880 29618 21456
rect 30602 20880 30636 21456
rect 31620 20880 31654 21456
rect 32638 20880 32672 21456
rect 33656 20880 33690 21456
rect 13082 19744 13116 20320
rect 14100 19744 14134 20320
rect 15118 19744 15152 20320
rect 16136 19744 16170 20320
rect 17154 19744 17188 20320
rect 18386 19624 18420 20200
rect 19404 19624 19438 20200
rect 20422 19624 20456 20200
rect 21440 19624 21474 20200
rect 22458 19624 22492 20200
rect 23476 19624 23510 20200
rect 24494 19624 24528 20200
rect 25512 19624 25546 20200
rect 26530 19624 26564 20200
rect 27548 19624 27582 20200
rect 28566 19624 28600 20200
rect 29584 19624 29618 20200
rect 30602 19624 30636 20200
rect 31620 19624 31654 20200
rect 32638 19624 32672 20200
rect 33656 19624 33690 20200
rect 13082 18712 13116 19288
rect 14100 18712 14134 19288
rect 15118 18712 15152 19288
rect 16136 18712 16170 19288
rect 17154 18712 17188 19288
rect 18386 18368 18420 18944
rect 19404 18368 19438 18944
rect 20422 18368 20456 18944
rect 21440 18368 21474 18944
rect 22458 18368 22492 18944
rect 23476 18368 23510 18944
rect 24494 18368 24528 18944
rect 25512 18368 25546 18944
rect 26530 18368 26564 18944
rect 27548 18368 27582 18944
rect 28566 18368 28600 18944
rect 29584 18368 29618 18944
rect 30602 18368 30636 18944
rect 31620 18368 31654 18944
rect 32638 18368 32672 18944
rect 33656 18368 33690 18944
rect 13082 17680 13116 18256
rect 14100 17680 14134 18256
rect 15118 17680 15152 18256
rect 16136 17680 16170 18256
rect 17154 17680 17188 18256
rect 18386 17112 18420 17688
rect 19404 17112 19438 17688
rect 20422 17112 20456 17688
rect 21440 17112 21474 17688
rect 22458 17112 22492 17688
rect 23476 17112 23510 17688
rect 24494 17112 24528 17688
rect 25512 17112 25546 17688
rect 26530 17112 26564 17688
rect 27548 17112 27582 17688
rect 28566 17112 28600 17688
rect 29584 17112 29618 17688
rect 30602 17112 30636 17688
rect 31620 17112 31654 17688
rect 32638 17112 32672 17688
rect 33656 17112 33690 17688
rect -12166 15738 -12132 16114
rect -11908 15738 -11874 16114
rect -11650 15738 -11616 16114
rect -11392 15738 -11358 16114
rect -11134 15738 -11100 16114
rect -10876 15738 -10842 16114
rect -10618 15738 -10584 16114
rect -10314 15697 -10280 15731
rect -10314 15629 -10280 15663
rect -10314 15561 -10280 15595
rect -10230 15697 -10196 15731
rect -10230 15629 -10196 15663
rect -10230 15561 -10196 15595
rect -9566 15738 -9532 16114
rect -9308 15738 -9274 16114
rect -9050 15738 -9016 16114
rect -8792 15738 -8758 16114
rect -8534 15738 -8500 16114
rect -8276 15738 -8242 16114
rect -8018 15738 -7984 16114
rect -7714 15697 -7680 15731
rect -7714 15629 -7680 15663
rect -7714 15561 -7680 15595
rect -7630 15697 -7596 15731
rect -7630 15629 -7596 15663
rect -7630 15561 -7596 15595
rect -7264 15697 -7230 15731
rect -7264 15629 -7230 15663
rect -7264 15561 -7230 15595
rect -7180 15697 -7146 15731
rect -7180 15629 -7146 15663
rect -7180 15561 -7146 15595
<< psubdiff >>
rect -12280 15342 -12184 15376
rect -10566 15342 -10470 15376
rect -12280 15280 -12246 15342
rect -10504 15280 -10470 15342
rect -9680 15342 -9584 15376
rect -7966 15342 -7870 15376
rect -12280 14862 -12246 14924
rect -9680 15280 -9646 15342
rect -10504 14862 -10470 14924
rect -12280 14828 -12184 14862
rect -10566 14828 -10470 14862
rect -7904 15280 -7870 15342
rect -9680 14862 -9646 14924
rect -7904 14862 -7870 14924
rect -9680 14828 -9584 14862
rect -7966 14828 -7870 14862
rect -1410 15262 -1248 15362
rect 35672 15262 35834 15362
rect -1410 15200 -1310 15262
rect 35734 15200 35834 15262
rect 13998 14756 14080 14780
rect 13998 14722 14022 14756
rect 14056 14722 14080 14756
rect 13998 14698 14080 14722
rect 15016 14756 15098 14780
rect 15016 14722 15040 14756
rect 15074 14722 15098 14756
rect 15016 14698 15098 14722
rect 16034 14756 16116 14780
rect 16034 14722 16058 14756
rect 16092 14722 16116 14756
rect 16034 14698 16116 14722
rect 17052 14756 17134 14780
rect 17052 14722 17076 14756
rect 17110 14722 17134 14756
rect 17052 14698 17134 14722
rect 18070 14756 18152 14780
rect 18070 14722 18094 14756
rect 18128 14722 18152 14756
rect 18070 14698 18152 14722
rect 19088 14756 19170 14780
rect 19088 14722 19112 14756
rect 19146 14722 19170 14756
rect 19088 14698 19170 14722
rect 20106 14756 20188 14780
rect 20106 14722 20130 14756
rect 20164 14722 20188 14756
rect 20106 14698 20188 14722
rect 21124 14756 21206 14780
rect 21124 14722 21148 14756
rect 21182 14722 21206 14756
rect 21124 14698 21206 14722
rect 22142 14756 22224 14780
rect 22142 14722 22166 14756
rect 22200 14722 22224 14756
rect 22142 14698 22224 14722
rect 23160 14756 23242 14780
rect 23160 14722 23184 14756
rect 23218 14722 23242 14756
rect 23160 14698 23242 14722
rect 24178 14756 24260 14780
rect 24178 14722 24202 14756
rect 24236 14722 24260 14756
rect 24178 14698 24260 14722
rect 25196 14756 25278 14780
rect 25196 14722 25220 14756
rect 25254 14722 25278 14756
rect 25196 14698 25278 14722
rect 26214 14756 26296 14780
rect 26214 14722 26238 14756
rect 26272 14722 26296 14756
rect 26214 14698 26296 14722
rect 27232 14756 27314 14780
rect 27232 14722 27256 14756
rect 27290 14722 27314 14756
rect 27232 14698 27314 14722
rect 28250 14756 28332 14780
rect 28250 14722 28274 14756
rect 28308 14722 28332 14756
rect 28250 14698 28332 14722
rect 29268 14756 29350 14780
rect 29268 14722 29292 14756
rect 29326 14722 29350 14756
rect 29268 14698 29350 14722
rect 30286 14756 30368 14780
rect 30286 14722 30310 14756
rect 30344 14722 30368 14756
rect 30286 14698 30368 14722
rect 31304 14756 31386 14780
rect 31304 14722 31328 14756
rect 31362 14722 31386 14756
rect 31304 14698 31386 14722
rect 32322 14756 32404 14780
rect 32322 14722 32346 14756
rect 32380 14722 32404 14756
rect 32322 14698 32404 14722
rect 33340 14756 33422 14780
rect 33340 14722 33364 14756
rect 33398 14722 33422 14756
rect 33340 14698 33422 14722
rect 1704 14154 1786 14178
rect 1704 14120 1728 14154
rect 1762 14120 1786 14154
rect 1704 14096 1786 14120
rect 2722 14154 2804 14178
rect 2722 14120 2746 14154
rect 2780 14120 2804 14154
rect 2722 14096 2804 14120
rect 3740 14154 3822 14178
rect 3740 14120 3764 14154
rect 3798 14120 3822 14154
rect 3740 14096 3822 14120
rect 4758 14154 4840 14178
rect 4758 14120 4782 14154
rect 4816 14120 4840 14154
rect 4758 14096 4840 14120
rect 5776 14154 5858 14178
rect 5776 14120 5800 14154
rect 5834 14120 5858 14154
rect 5776 14096 5858 14120
rect 6794 14154 6876 14178
rect 6794 14120 6818 14154
rect 6852 14120 6876 14154
rect 6794 14096 6876 14120
rect 7812 14154 7894 14178
rect 7812 14120 7836 14154
rect 7870 14120 7894 14154
rect 7812 14096 7894 14120
rect 8830 14154 8912 14178
rect 8830 14120 8854 14154
rect 8888 14120 8912 14154
rect 8830 14096 8912 14120
rect 9848 14154 9930 14178
rect 9848 14120 9872 14154
rect 9906 14120 9930 14154
rect 9848 14096 9930 14120
rect 10876 14154 10958 14178
rect 10876 14120 10900 14154
rect 10934 14120 10958 14154
rect 10876 14096 10958 14120
rect 1704 13336 1786 13360
rect 1704 13302 1728 13336
rect 1762 13302 1786 13336
rect 1704 13278 1786 13302
rect 2722 13336 2804 13360
rect 2722 13302 2746 13336
rect 2780 13302 2804 13336
rect 2722 13278 2804 13302
rect 3740 13336 3822 13360
rect 3740 13302 3764 13336
rect 3798 13302 3822 13336
rect 3740 13278 3822 13302
rect 4758 13336 4840 13360
rect 4758 13302 4782 13336
rect 4816 13302 4840 13336
rect 4758 13278 4840 13302
rect 5776 13336 5858 13360
rect 5776 13302 5800 13336
rect 5834 13302 5858 13336
rect 5776 13278 5858 13302
rect 6794 13336 6876 13360
rect 6794 13302 6818 13336
rect 6852 13302 6876 13336
rect 6794 13278 6876 13302
rect 7812 13336 7894 13360
rect 7812 13302 7836 13336
rect 7870 13302 7894 13336
rect 7812 13278 7894 13302
rect 8830 13336 8912 13360
rect 8830 13302 8854 13336
rect 8888 13302 8912 13336
rect 8830 13278 8912 13302
rect 9848 13336 9930 13360
rect 9848 13302 9872 13336
rect 9906 13302 9930 13336
rect 9848 13278 9930 13302
rect 10876 13336 10958 13360
rect 10876 13302 10900 13336
rect 10934 13302 10958 13336
rect 10876 13278 10958 13302
rect 14010 12730 14092 12754
rect 14010 12696 14034 12730
rect 14068 12696 14092 12730
rect 14010 12672 14092 12696
rect 15028 12730 15110 12754
rect 15028 12696 15052 12730
rect 15086 12696 15110 12730
rect 15028 12672 15110 12696
rect 16046 12730 16128 12754
rect 16046 12696 16070 12730
rect 16104 12696 16128 12730
rect 16046 12672 16128 12696
rect 17064 12730 17146 12754
rect 17064 12696 17088 12730
rect 17122 12696 17146 12730
rect 17064 12672 17146 12696
rect 18082 12730 18164 12754
rect 18082 12696 18106 12730
rect 18140 12696 18164 12730
rect 18082 12672 18164 12696
rect 19100 12730 19182 12754
rect 19100 12696 19124 12730
rect 19158 12696 19182 12730
rect 19100 12672 19182 12696
rect 20118 12730 20200 12754
rect 20118 12696 20142 12730
rect 20176 12696 20200 12730
rect 20118 12672 20200 12696
rect 21136 12730 21218 12754
rect 21136 12696 21160 12730
rect 21194 12696 21218 12730
rect 21136 12672 21218 12696
rect 22154 12730 22236 12754
rect 22154 12696 22178 12730
rect 22212 12696 22236 12730
rect 22154 12672 22236 12696
rect 23172 12730 23254 12754
rect 23172 12696 23196 12730
rect 23230 12696 23254 12730
rect 23172 12672 23254 12696
rect 24190 12730 24272 12754
rect 24190 12696 24214 12730
rect 24248 12696 24272 12730
rect 24190 12672 24272 12696
rect 25208 12730 25290 12754
rect 25208 12696 25232 12730
rect 25266 12696 25290 12730
rect 25208 12672 25290 12696
rect 26226 12730 26308 12754
rect 26226 12696 26250 12730
rect 26284 12696 26308 12730
rect 26226 12672 26308 12696
rect 27244 12730 27326 12754
rect 27244 12696 27268 12730
rect 27302 12696 27326 12730
rect 27244 12672 27326 12696
rect 28262 12730 28344 12754
rect 28262 12696 28286 12730
rect 28320 12696 28344 12730
rect 28262 12672 28344 12696
rect 29280 12730 29362 12754
rect 29280 12696 29304 12730
rect 29338 12696 29362 12730
rect 29280 12672 29362 12696
rect 30298 12730 30380 12754
rect 30298 12696 30322 12730
rect 30356 12696 30380 12730
rect 30298 12672 30380 12696
rect 31316 12730 31398 12754
rect 31316 12696 31340 12730
rect 31374 12696 31398 12730
rect 31316 12672 31398 12696
rect 32334 12730 32416 12754
rect 32334 12696 32358 12730
rect 32392 12696 32416 12730
rect 32334 12672 32416 12696
rect 33352 12730 33434 12754
rect 33352 12696 33376 12730
rect 33410 12696 33434 12730
rect 33352 12672 33434 12696
rect 1704 12518 1786 12542
rect 1704 12484 1728 12518
rect 1762 12484 1786 12518
rect 1704 12460 1786 12484
rect 2722 12518 2804 12542
rect 2722 12484 2746 12518
rect 2780 12484 2804 12518
rect 2722 12460 2804 12484
rect 3740 12518 3822 12542
rect 3740 12484 3764 12518
rect 3798 12484 3822 12518
rect 3740 12460 3822 12484
rect 4758 12518 4840 12542
rect 4758 12484 4782 12518
rect 4816 12484 4840 12518
rect 4758 12460 4840 12484
rect 5776 12518 5858 12542
rect 5776 12484 5800 12518
rect 5834 12484 5858 12518
rect 5776 12460 5858 12484
rect 6794 12518 6876 12542
rect 6794 12484 6818 12518
rect 6852 12484 6876 12518
rect 6794 12460 6876 12484
rect 7812 12518 7894 12542
rect 7812 12484 7836 12518
rect 7870 12484 7894 12518
rect 7812 12460 7894 12484
rect 8830 12518 8912 12542
rect 8830 12484 8854 12518
rect 8888 12484 8912 12518
rect 8830 12460 8912 12484
rect 9848 12518 9930 12542
rect 9848 12484 9872 12518
rect 9906 12484 9930 12518
rect 9848 12460 9930 12484
rect 10876 12518 10958 12542
rect 10876 12484 10900 12518
rect 10934 12484 10958 12518
rect 10876 12460 10958 12484
rect 1704 11700 1786 11724
rect 1704 11666 1728 11700
rect 1762 11666 1786 11700
rect 1704 11642 1786 11666
rect 2722 11700 2804 11724
rect 2722 11666 2746 11700
rect 2780 11666 2804 11700
rect 2722 11642 2804 11666
rect 3740 11700 3822 11724
rect 3740 11666 3764 11700
rect 3798 11666 3822 11700
rect 3740 11642 3822 11666
rect 4758 11700 4840 11724
rect 4758 11666 4782 11700
rect 4816 11666 4840 11700
rect 4758 11642 4840 11666
rect 5776 11700 5858 11724
rect 5776 11666 5800 11700
rect 5834 11666 5858 11700
rect 5776 11642 5858 11666
rect 6794 11700 6876 11724
rect 6794 11666 6818 11700
rect 6852 11666 6876 11700
rect 6794 11642 6876 11666
rect 7812 11700 7894 11724
rect 7812 11666 7836 11700
rect 7870 11666 7894 11700
rect 7812 11642 7894 11666
rect 8830 11700 8912 11724
rect 8830 11666 8854 11700
rect 8888 11666 8912 11700
rect 8830 11642 8912 11666
rect 9848 11700 9930 11724
rect 9848 11666 9872 11700
rect 9906 11666 9930 11700
rect 9848 11642 9930 11666
rect 10876 11700 10958 11724
rect 10876 11666 10900 11700
rect 10934 11666 10958 11700
rect 10876 11642 10958 11666
rect 13998 11424 14080 11448
rect 13998 11390 14022 11424
rect 14056 11390 14080 11424
rect 13998 11366 14080 11390
rect 15016 11424 15098 11448
rect 15016 11390 15040 11424
rect 15074 11390 15098 11424
rect 15016 11366 15098 11390
rect 16034 11424 16116 11448
rect 16034 11390 16058 11424
rect 16092 11390 16116 11424
rect 16034 11366 16116 11390
rect 17052 11424 17134 11448
rect 17052 11390 17076 11424
rect 17110 11390 17134 11424
rect 17052 11366 17134 11390
rect 18070 11424 18152 11448
rect 18070 11390 18094 11424
rect 18128 11390 18152 11424
rect 18070 11366 18152 11390
rect 19088 11424 19170 11448
rect 19088 11390 19112 11424
rect 19146 11390 19170 11424
rect 19088 11366 19170 11390
rect 20106 11424 20188 11448
rect 20106 11390 20130 11424
rect 20164 11390 20188 11424
rect 20106 11366 20188 11390
rect 21124 11424 21206 11448
rect 21124 11390 21148 11424
rect 21182 11390 21206 11424
rect 21124 11366 21206 11390
rect 22142 11424 22224 11448
rect 22142 11390 22166 11424
rect 22200 11390 22224 11424
rect 22142 11366 22224 11390
rect 23160 11424 23242 11448
rect 23160 11390 23184 11424
rect 23218 11390 23242 11424
rect 23160 11366 23242 11390
rect 24178 11424 24260 11448
rect 24178 11390 24202 11424
rect 24236 11390 24260 11424
rect 24178 11366 24260 11390
rect 25196 11424 25278 11448
rect 25196 11390 25220 11424
rect 25254 11390 25278 11424
rect 25196 11366 25278 11390
rect 26214 11424 26296 11448
rect 26214 11390 26238 11424
rect 26272 11390 26296 11424
rect 26214 11366 26296 11390
rect 27232 11424 27314 11448
rect 27232 11390 27256 11424
rect 27290 11390 27314 11424
rect 27232 11366 27314 11390
rect 28250 11424 28332 11448
rect 28250 11390 28274 11424
rect 28308 11390 28332 11424
rect 28250 11366 28332 11390
rect 29268 11424 29350 11448
rect 29268 11390 29292 11424
rect 29326 11390 29350 11424
rect 29268 11366 29350 11390
rect 30286 11424 30368 11448
rect 30286 11390 30310 11424
rect 30344 11390 30368 11424
rect 30286 11366 30368 11390
rect 31304 11424 31386 11448
rect 31304 11390 31328 11424
rect 31362 11390 31386 11424
rect 31304 11366 31386 11390
rect 32322 11424 32404 11448
rect 32322 11390 32346 11424
rect 32380 11390 32404 11424
rect 32322 11366 32404 11390
rect 33340 11424 33422 11448
rect 33340 11390 33364 11424
rect 33398 11390 33422 11424
rect 33340 11366 33422 11390
rect 1704 10882 1786 10906
rect 1704 10848 1728 10882
rect 1762 10848 1786 10882
rect 1704 10824 1786 10848
rect 2722 10882 2804 10906
rect 2722 10848 2746 10882
rect 2780 10848 2804 10882
rect 2722 10824 2804 10848
rect 3740 10882 3822 10906
rect 3740 10848 3764 10882
rect 3798 10848 3822 10882
rect 3740 10824 3822 10848
rect 4758 10882 4840 10906
rect 4758 10848 4782 10882
rect 4816 10848 4840 10882
rect 4758 10824 4840 10848
rect 5776 10882 5858 10906
rect 5776 10848 5800 10882
rect 5834 10848 5858 10882
rect 5776 10824 5858 10848
rect 6794 10882 6876 10906
rect 6794 10848 6818 10882
rect 6852 10848 6876 10882
rect 6794 10824 6876 10848
rect 7812 10882 7894 10906
rect 7812 10848 7836 10882
rect 7870 10848 7894 10882
rect 7812 10824 7894 10848
rect 8830 10882 8912 10906
rect 8830 10848 8854 10882
rect 8888 10848 8912 10882
rect 8830 10824 8912 10848
rect 9848 10882 9930 10906
rect 9848 10848 9872 10882
rect 9906 10848 9930 10882
rect 9848 10824 9930 10848
rect 10876 10882 10958 10906
rect 10876 10848 10900 10882
rect 10934 10848 10958 10882
rect 10876 10824 10958 10848
rect 13986 10188 14068 10212
rect 1704 10064 1786 10088
rect 1704 10030 1728 10064
rect 1762 10030 1786 10064
rect 1704 10006 1786 10030
rect 2722 10064 2804 10088
rect 2722 10030 2746 10064
rect 2780 10030 2804 10064
rect 2722 10006 2804 10030
rect 3740 10064 3822 10088
rect 3740 10030 3764 10064
rect 3798 10030 3822 10064
rect 3740 10006 3822 10030
rect 4758 10064 4840 10088
rect 4758 10030 4782 10064
rect 4816 10030 4840 10064
rect 4758 10006 4840 10030
rect 5776 10064 5858 10088
rect 5776 10030 5800 10064
rect 5834 10030 5858 10064
rect 5776 10006 5858 10030
rect 6794 10064 6876 10088
rect 6794 10030 6818 10064
rect 6852 10030 6876 10064
rect 6794 10006 6876 10030
rect 7812 10064 7894 10088
rect 7812 10030 7836 10064
rect 7870 10030 7894 10064
rect 7812 10006 7894 10030
rect 8830 10064 8912 10088
rect 13986 10154 14010 10188
rect 14044 10154 14068 10188
rect 13986 10130 14068 10154
rect 15004 10188 15086 10212
rect 15004 10154 15028 10188
rect 15062 10154 15086 10188
rect 15004 10130 15086 10154
rect 16022 10188 16104 10212
rect 16022 10154 16046 10188
rect 16080 10154 16104 10188
rect 16022 10130 16104 10154
rect 17040 10188 17122 10212
rect 17040 10154 17064 10188
rect 17098 10154 17122 10188
rect 17040 10130 17122 10154
rect 18058 10188 18140 10212
rect 18058 10154 18082 10188
rect 18116 10154 18140 10188
rect 18058 10130 18140 10154
rect 19076 10188 19158 10212
rect 19076 10154 19100 10188
rect 19134 10154 19158 10188
rect 19076 10130 19158 10154
rect 20094 10188 20176 10212
rect 20094 10154 20118 10188
rect 20152 10154 20176 10188
rect 20094 10130 20176 10154
rect 21112 10188 21194 10212
rect 21112 10154 21136 10188
rect 21170 10154 21194 10188
rect 21112 10130 21194 10154
rect 22130 10188 22212 10212
rect 22130 10154 22154 10188
rect 22188 10154 22212 10188
rect 22130 10130 22212 10154
rect 23148 10188 23230 10212
rect 23148 10154 23172 10188
rect 23206 10154 23230 10188
rect 23148 10130 23230 10154
rect 24166 10188 24248 10212
rect 24166 10154 24190 10188
rect 24224 10154 24248 10188
rect 24166 10130 24248 10154
rect 25184 10188 25266 10212
rect 25184 10154 25208 10188
rect 25242 10154 25266 10188
rect 25184 10130 25266 10154
rect 26202 10188 26284 10212
rect 26202 10154 26226 10188
rect 26260 10154 26284 10188
rect 26202 10130 26284 10154
rect 27220 10188 27302 10212
rect 27220 10154 27244 10188
rect 27278 10154 27302 10188
rect 27220 10130 27302 10154
rect 28238 10188 28320 10212
rect 28238 10154 28262 10188
rect 28296 10154 28320 10188
rect 28238 10130 28320 10154
rect 29256 10188 29338 10212
rect 29256 10154 29280 10188
rect 29314 10154 29338 10188
rect 29256 10130 29338 10154
rect 30274 10188 30356 10212
rect 30274 10154 30298 10188
rect 30332 10154 30356 10188
rect 30274 10130 30356 10154
rect 31292 10188 31374 10212
rect 31292 10154 31316 10188
rect 31350 10154 31374 10188
rect 31292 10130 31374 10154
rect 32310 10188 32392 10212
rect 32310 10154 32334 10188
rect 32368 10154 32392 10188
rect 32310 10130 32392 10154
rect 33328 10188 33410 10212
rect 33328 10154 33352 10188
rect 33386 10154 33410 10188
rect 33328 10130 33410 10154
rect 8830 10030 8854 10064
rect 8888 10030 8912 10064
rect 8830 10006 8912 10030
rect 9848 10064 9930 10088
rect 9848 10030 9872 10064
rect 9906 10030 9930 10064
rect 9848 10006 9930 10030
rect 10876 10064 10958 10088
rect 10876 10030 10900 10064
rect 10934 10030 10958 10064
rect 10876 10006 10958 10030
rect 1704 9246 1786 9270
rect 1704 9212 1728 9246
rect 1762 9212 1786 9246
rect 1704 9188 1786 9212
rect 2722 9246 2804 9270
rect 2722 9212 2746 9246
rect 2780 9212 2804 9246
rect 2722 9188 2804 9212
rect 3740 9246 3822 9270
rect 3740 9212 3764 9246
rect 3798 9212 3822 9246
rect 3740 9188 3822 9212
rect 4758 9246 4840 9270
rect 4758 9212 4782 9246
rect 4816 9212 4840 9246
rect 4758 9188 4840 9212
rect 5776 9246 5858 9270
rect 5776 9212 5800 9246
rect 5834 9212 5858 9246
rect 5776 9188 5858 9212
rect 6794 9246 6876 9270
rect 6794 9212 6818 9246
rect 6852 9212 6876 9246
rect 6794 9188 6876 9212
rect 7812 9246 7894 9270
rect 7812 9212 7836 9246
rect 7870 9212 7894 9246
rect 7812 9188 7894 9212
rect 8830 9246 8912 9270
rect 8830 9212 8854 9246
rect 8888 9212 8912 9246
rect 8830 9188 8912 9212
rect 9848 9246 9930 9270
rect 9848 9212 9872 9246
rect 9906 9212 9930 9246
rect 9848 9188 9930 9212
rect 10876 9246 10958 9270
rect 10876 9212 10900 9246
rect 10934 9212 10958 9246
rect 10876 9188 10958 9212
rect 13986 8964 14068 8988
rect 13986 8930 14010 8964
rect 14044 8930 14068 8964
rect 13986 8906 14068 8930
rect 15004 8964 15086 8988
rect 15004 8930 15028 8964
rect 15062 8930 15086 8964
rect 15004 8906 15086 8930
rect 16022 8964 16104 8988
rect 16022 8930 16046 8964
rect 16080 8930 16104 8964
rect 16022 8906 16104 8930
rect 17040 8964 17122 8988
rect 17040 8930 17064 8964
rect 17098 8930 17122 8964
rect 17040 8906 17122 8930
rect 18058 8964 18140 8988
rect 18058 8930 18082 8964
rect 18116 8930 18140 8964
rect 18058 8906 18140 8930
rect 19076 8964 19158 8988
rect 19076 8930 19100 8964
rect 19134 8930 19158 8964
rect 19076 8906 19158 8930
rect 20094 8964 20176 8988
rect 20094 8930 20118 8964
rect 20152 8930 20176 8964
rect 20094 8906 20176 8930
rect 21112 8964 21194 8988
rect 21112 8930 21136 8964
rect 21170 8930 21194 8964
rect 21112 8906 21194 8930
rect 22130 8964 22212 8988
rect 22130 8930 22154 8964
rect 22188 8930 22212 8964
rect 22130 8906 22212 8930
rect 23148 8964 23230 8988
rect 23148 8930 23172 8964
rect 23206 8930 23230 8964
rect 23148 8906 23230 8930
rect 24166 8964 24248 8988
rect 24166 8930 24190 8964
rect 24224 8930 24248 8964
rect 24166 8906 24248 8930
rect 25184 8964 25266 8988
rect 25184 8930 25208 8964
rect 25242 8930 25266 8964
rect 25184 8906 25266 8930
rect 26202 8964 26284 8988
rect 26202 8930 26226 8964
rect 26260 8930 26284 8964
rect 26202 8906 26284 8930
rect 27220 8964 27302 8988
rect 27220 8930 27244 8964
rect 27278 8930 27302 8964
rect 27220 8906 27302 8930
rect 28238 8964 28320 8988
rect 28238 8930 28262 8964
rect 28296 8930 28320 8964
rect 28238 8906 28320 8930
rect 29256 8964 29338 8988
rect 29256 8930 29280 8964
rect 29314 8930 29338 8964
rect 29256 8906 29338 8930
rect 30274 8964 30356 8988
rect 30274 8930 30298 8964
rect 30332 8930 30356 8964
rect 30274 8906 30356 8930
rect 31292 8964 31374 8988
rect 31292 8930 31316 8964
rect 31350 8930 31374 8964
rect 31292 8906 31374 8930
rect 32310 8964 32392 8988
rect 32310 8930 32334 8964
rect 32368 8930 32392 8964
rect 32310 8906 32392 8930
rect 33328 8964 33410 8988
rect 33328 8930 33352 8964
rect 33386 8930 33410 8964
rect 33328 8906 33410 8930
rect 1704 8428 1786 8452
rect 1704 8394 1728 8428
rect 1762 8394 1786 8428
rect 1704 8370 1786 8394
rect 2722 8428 2804 8452
rect 2722 8394 2746 8428
rect 2780 8394 2804 8428
rect 2722 8370 2804 8394
rect 3740 8428 3822 8452
rect 3740 8394 3764 8428
rect 3798 8394 3822 8428
rect 3740 8370 3822 8394
rect 4758 8428 4840 8452
rect 4758 8394 4782 8428
rect 4816 8394 4840 8428
rect 4758 8370 4840 8394
rect 5776 8428 5858 8452
rect 5776 8394 5800 8428
rect 5834 8394 5858 8428
rect 5776 8370 5858 8394
rect 6794 8428 6876 8452
rect 6794 8394 6818 8428
rect 6852 8394 6876 8428
rect 6794 8370 6876 8394
rect 7812 8428 7894 8452
rect 7812 8394 7836 8428
rect 7870 8394 7894 8428
rect 7812 8370 7894 8394
rect 8830 8428 8912 8452
rect 8830 8394 8854 8428
rect 8888 8394 8912 8428
rect 8830 8370 8912 8394
rect 9848 8428 9930 8452
rect 9848 8394 9872 8428
rect 9906 8394 9930 8428
rect 9848 8370 9930 8394
rect 10876 8428 10958 8452
rect 10876 8394 10900 8428
rect 10934 8394 10958 8428
rect 10876 8370 10958 8394
rect 13998 7728 14080 7752
rect 13998 7694 14022 7728
rect 14056 7694 14080 7728
rect 13998 7670 14080 7694
rect 15016 7728 15098 7752
rect 15016 7694 15040 7728
rect 15074 7694 15098 7728
rect 15016 7670 15098 7694
rect 16034 7728 16116 7752
rect 16034 7694 16058 7728
rect 16092 7694 16116 7728
rect 16034 7670 16116 7694
rect 17052 7728 17134 7752
rect 17052 7694 17076 7728
rect 17110 7694 17134 7728
rect 17052 7670 17134 7694
rect 18070 7728 18152 7752
rect 18070 7694 18094 7728
rect 18128 7694 18152 7728
rect 18070 7670 18152 7694
rect 19088 7728 19170 7752
rect 19088 7694 19112 7728
rect 19146 7694 19170 7728
rect 19088 7670 19170 7694
rect 20106 7728 20188 7752
rect 20106 7694 20130 7728
rect 20164 7694 20188 7728
rect 20106 7670 20188 7694
rect 21124 7728 21206 7752
rect 21124 7694 21148 7728
rect 21182 7694 21206 7728
rect 21124 7670 21206 7694
rect 22142 7728 22224 7752
rect 22142 7694 22166 7728
rect 22200 7694 22224 7728
rect 22142 7670 22224 7694
rect 23160 7728 23242 7752
rect 23160 7694 23184 7728
rect 23218 7694 23242 7728
rect 23160 7670 23242 7694
rect 24178 7728 24260 7752
rect 24178 7694 24202 7728
rect 24236 7694 24260 7728
rect 24178 7670 24260 7694
rect 25196 7728 25278 7752
rect 25196 7694 25220 7728
rect 25254 7694 25278 7728
rect 25196 7670 25278 7694
rect 26214 7728 26296 7752
rect 26214 7694 26238 7728
rect 26272 7694 26296 7728
rect 26214 7670 26296 7694
rect 27232 7728 27314 7752
rect 27232 7694 27256 7728
rect 27290 7694 27314 7728
rect 27232 7670 27314 7694
rect 28250 7728 28332 7752
rect 28250 7694 28274 7728
rect 28308 7694 28332 7728
rect 28250 7670 28332 7694
rect 29268 7728 29350 7752
rect 29268 7694 29292 7728
rect 29326 7694 29350 7728
rect 29268 7670 29350 7694
rect 30286 7728 30368 7752
rect 30286 7694 30310 7728
rect 30344 7694 30368 7728
rect 30286 7670 30368 7694
rect 31304 7728 31386 7752
rect 31304 7694 31328 7728
rect 31362 7694 31386 7728
rect 31304 7670 31386 7694
rect 32322 7728 32404 7752
rect 32322 7694 32346 7728
rect 32380 7694 32404 7728
rect 32322 7670 32404 7694
rect 33340 7728 33422 7752
rect 33340 7694 33364 7728
rect 33398 7694 33422 7728
rect 33340 7670 33422 7694
rect 1692 7534 1774 7558
rect 1692 7500 1716 7534
rect 1750 7500 1774 7534
rect 1692 7476 1774 7500
rect 2710 7534 2792 7558
rect 2710 7500 2734 7534
rect 2768 7500 2792 7534
rect 2710 7476 2792 7500
rect 3728 7534 3810 7558
rect 3728 7500 3752 7534
rect 3786 7500 3810 7534
rect 3728 7476 3810 7500
rect 4746 7534 4828 7558
rect 4746 7500 4770 7534
rect 4804 7500 4828 7534
rect 4746 7476 4828 7500
rect 5764 7534 5846 7558
rect 5764 7500 5788 7534
rect 5822 7500 5846 7534
rect 5764 7476 5846 7500
rect 6782 7534 6864 7558
rect 6782 7500 6806 7534
rect 6840 7500 6864 7534
rect 6782 7476 6864 7500
rect 7800 7534 7882 7558
rect 7800 7500 7824 7534
rect 7858 7500 7882 7534
rect 7800 7476 7882 7500
rect 8818 7534 8900 7558
rect 8818 7500 8842 7534
rect 8876 7500 8900 7534
rect 8818 7476 8900 7500
rect 9836 7534 9918 7558
rect 9836 7500 9860 7534
rect 9894 7500 9918 7534
rect 9836 7476 9918 7500
rect 10864 7534 10946 7558
rect 10864 7500 10888 7534
rect 10922 7500 10946 7534
rect 10864 7476 10946 7500
rect 896 6586 978 6610
rect 896 6552 920 6586
rect 954 6552 978 6586
rect 896 6528 978 6552
rect 1914 6586 1996 6610
rect 1914 6552 1938 6586
rect 1972 6552 1996 6586
rect 1914 6528 1996 6552
rect 2932 6586 3014 6610
rect 2932 6552 2956 6586
rect 2990 6552 3014 6586
rect 2932 6528 3014 6552
rect 3950 6586 4032 6610
rect 3950 6552 3974 6586
rect 4008 6552 4032 6586
rect 3950 6528 4032 6552
rect 4968 6586 5050 6610
rect 4968 6552 4992 6586
rect 5026 6552 5050 6586
rect 4968 6528 5050 6552
rect 5986 6586 6068 6610
rect 5986 6552 6010 6586
rect 6044 6552 6068 6586
rect 5986 6528 6068 6552
rect 7004 6586 7086 6610
rect 7004 6552 7028 6586
rect 7062 6552 7086 6586
rect 7004 6528 7086 6552
rect 8022 6586 8104 6610
rect 8022 6552 8046 6586
rect 8080 6552 8104 6586
rect 8022 6528 8104 6552
rect 9040 6586 9122 6610
rect 9040 6552 9064 6586
rect 9098 6552 9122 6586
rect 9040 6528 9122 6552
rect 10058 6586 10140 6610
rect 10058 6552 10082 6586
rect 10116 6552 10140 6586
rect 10058 6528 10140 6552
rect 11076 6586 11158 6610
rect 11076 6552 11100 6586
rect 11134 6552 11158 6586
rect 11076 6528 11158 6552
rect 13998 6480 14080 6504
rect 13998 6446 14022 6480
rect 14056 6446 14080 6480
rect 13998 6422 14080 6446
rect 15016 6480 15098 6504
rect 15016 6446 15040 6480
rect 15074 6446 15098 6480
rect 15016 6422 15098 6446
rect 16034 6480 16116 6504
rect 16034 6446 16058 6480
rect 16092 6446 16116 6480
rect 16034 6422 16116 6446
rect 17052 6480 17134 6504
rect 17052 6446 17076 6480
rect 17110 6446 17134 6480
rect 17052 6422 17134 6446
rect 18070 6480 18152 6504
rect 18070 6446 18094 6480
rect 18128 6446 18152 6480
rect 18070 6422 18152 6446
rect 19088 6480 19170 6504
rect 19088 6446 19112 6480
rect 19146 6446 19170 6480
rect 19088 6422 19170 6446
rect 20106 6480 20188 6504
rect 20106 6446 20130 6480
rect 20164 6446 20188 6480
rect 20106 6422 20188 6446
rect 21124 6480 21206 6504
rect 21124 6446 21148 6480
rect 21182 6446 21206 6480
rect 21124 6422 21206 6446
rect 22142 6480 22224 6504
rect 22142 6446 22166 6480
rect 22200 6446 22224 6480
rect 22142 6422 22224 6446
rect 23160 6480 23242 6504
rect 23160 6446 23184 6480
rect 23218 6446 23242 6480
rect 23160 6422 23242 6446
rect 24178 6480 24260 6504
rect 24178 6446 24202 6480
rect 24236 6446 24260 6480
rect 24178 6422 24260 6446
rect 25196 6480 25278 6504
rect 25196 6446 25220 6480
rect 25254 6446 25278 6480
rect 25196 6422 25278 6446
rect 26214 6480 26296 6504
rect 26214 6446 26238 6480
rect 26272 6446 26296 6480
rect 26214 6422 26296 6446
rect 27232 6480 27314 6504
rect 27232 6446 27256 6480
rect 27290 6446 27314 6480
rect 27232 6422 27314 6446
rect 28250 6480 28332 6504
rect 28250 6446 28274 6480
rect 28308 6446 28332 6480
rect 28250 6422 28332 6446
rect 29268 6480 29350 6504
rect 29268 6446 29292 6480
rect 29326 6446 29350 6480
rect 29268 6422 29350 6446
rect 30286 6480 30368 6504
rect 30286 6446 30310 6480
rect 30344 6446 30368 6480
rect 30286 6422 30368 6446
rect 31304 6480 31386 6504
rect 31304 6446 31328 6480
rect 31362 6446 31386 6480
rect 31304 6422 31386 6446
rect 32322 6480 32404 6504
rect 32322 6446 32346 6480
rect 32380 6446 32404 6480
rect 32322 6422 32404 6446
rect 33340 6480 33422 6504
rect 33340 6446 33364 6480
rect 33398 6446 33422 6480
rect 33340 6422 33422 6446
rect 908 5444 990 5468
rect 908 5410 932 5444
rect 966 5410 990 5444
rect 908 5386 990 5410
rect 1926 5444 2008 5468
rect 1926 5410 1950 5444
rect 1984 5410 2008 5444
rect 1926 5386 2008 5410
rect 2944 5444 3026 5468
rect 2944 5410 2968 5444
rect 3002 5410 3026 5444
rect 2944 5386 3026 5410
rect 3962 5444 4044 5468
rect 3962 5410 3986 5444
rect 4020 5410 4044 5444
rect 3962 5386 4044 5410
rect 4980 5444 5062 5468
rect 4980 5410 5004 5444
rect 5038 5410 5062 5444
rect 4980 5386 5062 5410
rect 5998 5444 6080 5468
rect 5998 5410 6022 5444
rect 6056 5410 6080 5444
rect 5998 5386 6080 5410
rect 7016 5444 7098 5468
rect 7016 5410 7040 5444
rect 7074 5410 7098 5444
rect 7016 5386 7098 5410
rect 8034 5444 8116 5468
rect 8034 5410 8058 5444
rect 8092 5410 8116 5444
rect 8034 5386 8116 5410
rect 9052 5444 9134 5468
rect 9052 5410 9076 5444
rect 9110 5410 9134 5444
rect 9052 5386 9134 5410
rect 10070 5444 10152 5468
rect 10070 5410 10094 5444
rect 10128 5410 10152 5444
rect 10070 5386 10152 5410
rect 11088 5444 11170 5468
rect 11088 5410 11112 5444
rect 11146 5410 11170 5444
rect 11088 5386 11170 5410
rect 13974 5244 14056 5268
rect 13974 5210 13998 5244
rect 14032 5210 14056 5244
rect 13974 5186 14056 5210
rect 14992 5244 15074 5268
rect 14992 5210 15016 5244
rect 15050 5210 15074 5244
rect 14992 5186 15074 5210
rect 16010 5244 16092 5268
rect 16010 5210 16034 5244
rect 16068 5210 16092 5244
rect 16010 5186 16092 5210
rect 17028 5244 17110 5268
rect 17028 5210 17052 5244
rect 17086 5210 17110 5244
rect 17028 5186 17110 5210
rect 18046 5244 18128 5268
rect 18046 5210 18070 5244
rect 18104 5210 18128 5244
rect 18046 5186 18128 5210
rect 19064 5244 19146 5268
rect 19064 5210 19088 5244
rect 19122 5210 19146 5244
rect 19064 5186 19146 5210
rect 20082 5244 20164 5268
rect 20082 5210 20106 5244
rect 20140 5210 20164 5244
rect 20082 5186 20164 5210
rect 21100 5244 21182 5268
rect 21100 5210 21124 5244
rect 21158 5210 21182 5244
rect 21100 5186 21182 5210
rect 22118 5244 22200 5268
rect 22118 5210 22142 5244
rect 22176 5210 22200 5244
rect 22118 5186 22200 5210
rect 23136 5244 23218 5268
rect 23136 5210 23160 5244
rect 23194 5210 23218 5244
rect 23136 5186 23218 5210
rect 24154 5244 24236 5268
rect 24154 5210 24178 5244
rect 24212 5210 24236 5244
rect 24154 5186 24236 5210
rect 25172 5244 25254 5268
rect 25172 5210 25196 5244
rect 25230 5210 25254 5244
rect 25172 5186 25254 5210
rect 26190 5244 26272 5268
rect 26190 5210 26214 5244
rect 26248 5210 26272 5244
rect 26190 5186 26272 5210
rect 27208 5244 27290 5268
rect 27208 5210 27232 5244
rect 27266 5210 27290 5244
rect 27208 5186 27290 5210
rect 28226 5244 28308 5268
rect 28226 5210 28250 5244
rect 28284 5210 28308 5244
rect 28226 5186 28308 5210
rect 29244 5244 29326 5268
rect 29244 5210 29268 5244
rect 29302 5210 29326 5244
rect 29244 5186 29326 5210
rect 30262 5244 30344 5268
rect 30262 5210 30286 5244
rect 30320 5210 30344 5244
rect 30262 5186 30344 5210
rect 31280 5244 31362 5268
rect 31280 5210 31304 5244
rect 31338 5210 31362 5244
rect 31280 5186 31362 5210
rect 32298 5244 32380 5268
rect 32298 5210 32322 5244
rect 32356 5210 32380 5244
rect 32298 5186 32380 5210
rect 33316 5244 33398 5268
rect 33316 5210 33340 5244
rect 33374 5210 33398 5244
rect 33316 5186 33398 5210
rect 886 4336 968 4360
rect 886 4302 910 4336
rect 944 4302 968 4336
rect 886 4278 968 4302
rect 1904 4336 1986 4360
rect 1904 4302 1928 4336
rect 1962 4302 1986 4336
rect 1904 4278 1986 4302
rect 2922 4336 3004 4360
rect 2922 4302 2946 4336
rect 2980 4302 3004 4336
rect 2922 4278 3004 4302
rect 3940 4336 4022 4360
rect 3940 4302 3964 4336
rect 3998 4302 4022 4336
rect 3940 4278 4022 4302
rect 4958 4336 5040 4360
rect 4958 4302 4982 4336
rect 5016 4302 5040 4336
rect 4958 4278 5040 4302
rect 5976 4336 6058 4360
rect 5976 4302 6000 4336
rect 6034 4302 6058 4336
rect 5976 4278 6058 4302
rect 6994 4336 7076 4360
rect 6994 4302 7018 4336
rect 7052 4302 7076 4336
rect 6994 4278 7076 4302
rect 8012 4336 8094 4360
rect 8012 4302 8036 4336
rect 8070 4302 8094 4336
rect 8012 4278 8094 4302
rect 9030 4336 9112 4360
rect 9030 4302 9054 4336
rect 9088 4302 9112 4336
rect 9030 4278 9112 4302
rect 10048 4336 10130 4360
rect 10048 4302 10072 4336
rect 10106 4302 10130 4336
rect 10048 4278 10130 4302
rect 11066 4336 11148 4360
rect 11066 4302 11090 4336
rect 11124 4302 11148 4336
rect 11066 4278 11148 4302
rect 13986 4020 14068 4044
rect 13986 3986 14010 4020
rect 14044 3986 14068 4020
rect 13986 3962 14068 3986
rect 15004 4020 15086 4044
rect 15004 3986 15028 4020
rect 15062 3986 15086 4020
rect 15004 3962 15086 3986
rect 16022 4020 16104 4044
rect 16022 3986 16046 4020
rect 16080 3986 16104 4020
rect 16022 3962 16104 3986
rect 17040 4020 17122 4044
rect 17040 3986 17064 4020
rect 17098 3986 17122 4020
rect 17040 3962 17122 3986
rect 18058 4020 18140 4044
rect 18058 3986 18082 4020
rect 18116 3986 18140 4020
rect 18058 3962 18140 3986
rect 19076 4020 19158 4044
rect 19076 3986 19100 4020
rect 19134 3986 19158 4020
rect 19076 3962 19158 3986
rect 20094 4020 20176 4044
rect 20094 3986 20118 4020
rect 20152 3986 20176 4020
rect 20094 3962 20176 3986
rect 21112 4020 21194 4044
rect 21112 3986 21136 4020
rect 21170 3986 21194 4020
rect 21112 3962 21194 3986
rect 22130 4020 22212 4044
rect 22130 3986 22154 4020
rect 22188 3986 22212 4020
rect 22130 3962 22212 3986
rect 23148 4020 23230 4044
rect 23148 3986 23172 4020
rect 23206 3986 23230 4020
rect 23148 3962 23230 3986
rect 24166 4020 24248 4044
rect 24166 3986 24190 4020
rect 24224 3986 24248 4020
rect 24166 3962 24248 3986
rect 25184 4020 25266 4044
rect 25184 3986 25208 4020
rect 25242 3986 25266 4020
rect 25184 3962 25266 3986
rect 26202 4020 26284 4044
rect 26202 3986 26226 4020
rect 26260 3986 26284 4020
rect 26202 3962 26284 3986
rect 27220 4020 27302 4044
rect 27220 3986 27244 4020
rect 27278 3986 27302 4020
rect 27220 3962 27302 3986
rect 28238 4020 28320 4044
rect 28238 3986 28262 4020
rect 28296 3986 28320 4020
rect 28238 3962 28320 3986
rect 29256 4020 29338 4044
rect 29256 3986 29280 4020
rect 29314 3986 29338 4020
rect 29256 3962 29338 3986
rect 30274 4020 30356 4044
rect 30274 3986 30298 4020
rect 30332 3986 30356 4020
rect 30274 3962 30356 3986
rect 31292 4020 31374 4044
rect 31292 3986 31316 4020
rect 31350 3986 31374 4020
rect 31292 3962 31374 3986
rect 32310 4020 32392 4044
rect 32310 3986 32334 4020
rect 32368 3986 32392 4020
rect 32310 3962 32392 3986
rect 33328 4020 33410 4044
rect 33328 3986 33352 4020
rect 33386 3986 33410 4020
rect 33328 3962 33410 3986
rect 886 3230 968 3254
rect 886 3196 910 3230
rect 944 3196 968 3230
rect 886 3172 968 3196
rect 1904 3230 1986 3254
rect 1904 3196 1928 3230
rect 1962 3196 1986 3230
rect 1904 3172 1986 3196
rect 2922 3230 3004 3254
rect 2922 3196 2946 3230
rect 2980 3196 3004 3230
rect 2922 3172 3004 3196
rect 3940 3230 4022 3254
rect 3940 3196 3964 3230
rect 3998 3196 4022 3230
rect 3940 3172 4022 3196
rect 4958 3230 5040 3254
rect 4958 3196 4982 3230
rect 5016 3196 5040 3230
rect 4958 3172 5040 3196
rect 5976 3230 6058 3254
rect 5976 3196 6000 3230
rect 6034 3196 6058 3230
rect 5976 3172 6058 3196
rect 6994 3230 7076 3254
rect 6994 3196 7018 3230
rect 7052 3196 7076 3230
rect 6994 3172 7076 3196
rect 8012 3230 8094 3254
rect 8012 3196 8036 3230
rect 8070 3196 8094 3230
rect 8012 3172 8094 3196
rect 9030 3230 9112 3254
rect 9030 3196 9054 3230
rect 9088 3196 9112 3230
rect 9030 3172 9112 3196
rect 10048 3230 10130 3254
rect 10048 3196 10072 3230
rect 10106 3196 10130 3230
rect 10048 3172 10130 3196
rect 11066 3230 11148 3254
rect 11066 3196 11090 3230
rect 11124 3196 11148 3230
rect 11066 3172 11148 3196
rect 13986 2784 14068 2808
rect 13986 2750 14010 2784
rect 14044 2750 14068 2784
rect 13986 2726 14068 2750
rect 15004 2784 15086 2808
rect 15004 2750 15028 2784
rect 15062 2750 15086 2784
rect 15004 2726 15086 2750
rect 16022 2784 16104 2808
rect 16022 2750 16046 2784
rect 16080 2750 16104 2784
rect 16022 2726 16104 2750
rect 17040 2784 17122 2808
rect 17040 2750 17064 2784
rect 17098 2750 17122 2784
rect 17040 2726 17122 2750
rect 18058 2784 18140 2808
rect 18058 2750 18082 2784
rect 18116 2750 18140 2784
rect 18058 2726 18140 2750
rect 19076 2784 19158 2808
rect 19076 2750 19100 2784
rect 19134 2750 19158 2784
rect 19076 2726 19158 2750
rect 20094 2784 20176 2808
rect 20094 2750 20118 2784
rect 20152 2750 20176 2784
rect 20094 2726 20176 2750
rect 21112 2784 21194 2808
rect 21112 2750 21136 2784
rect 21170 2750 21194 2784
rect 21112 2726 21194 2750
rect 22130 2784 22212 2808
rect 22130 2750 22154 2784
rect 22188 2750 22212 2784
rect 22130 2726 22212 2750
rect 23148 2784 23230 2808
rect 23148 2750 23172 2784
rect 23206 2750 23230 2784
rect 23148 2726 23230 2750
rect 24166 2784 24248 2808
rect 24166 2750 24190 2784
rect 24224 2750 24248 2784
rect 24166 2726 24248 2750
rect 25184 2784 25266 2808
rect 25184 2750 25208 2784
rect 25242 2750 25266 2784
rect 25184 2726 25266 2750
rect 26202 2784 26284 2808
rect 26202 2750 26226 2784
rect 26260 2750 26284 2784
rect 26202 2726 26284 2750
rect 27220 2784 27302 2808
rect 27220 2750 27244 2784
rect 27278 2750 27302 2784
rect 27220 2726 27302 2750
rect 28238 2784 28320 2808
rect 28238 2750 28262 2784
rect 28296 2750 28320 2784
rect 28238 2726 28320 2750
rect 29256 2784 29338 2808
rect 29256 2750 29280 2784
rect 29314 2750 29338 2784
rect 29256 2726 29338 2750
rect 30274 2784 30356 2808
rect 30274 2750 30298 2784
rect 30332 2750 30356 2784
rect 30274 2726 30356 2750
rect 31292 2784 31374 2808
rect 31292 2750 31316 2784
rect 31350 2750 31374 2784
rect 31292 2726 31374 2750
rect 32310 2784 32392 2808
rect 32310 2750 32334 2784
rect 32368 2750 32392 2784
rect 32310 2726 32392 2750
rect 33328 2784 33410 2808
rect 33328 2750 33352 2784
rect 33386 2750 33410 2784
rect 33328 2726 33410 2750
rect 886 1888 968 1912
rect 886 1854 910 1888
rect 944 1854 968 1888
rect 886 1830 968 1854
rect 1904 1888 1986 1912
rect 1904 1854 1928 1888
rect 1962 1854 1986 1888
rect 1904 1830 1986 1854
rect 2922 1888 3004 1912
rect 2922 1854 2946 1888
rect 2980 1854 3004 1888
rect 2922 1830 3004 1854
rect 3940 1888 4022 1912
rect 3940 1854 3964 1888
rect 3998 1854 4022 1888
rect 3940 1830 4022 1854
rect 4958 1888 5040 1912
rect 4958 1854 4982 1888
rect 5016 1854 5040 1888
rect 4958 1830 5040 1854
rect 5976 1888 6058 1912
rect 5976 1854 6000 1888
rect 6034 1854 6058 1888
rect 5976 1830 6058 1854
rect 6994 1888 7076 1912
rect 6994 1854 7018 1888
rect 7052 1854 7076 1888
rect 6994 1830 7076 1854
rect 8012 1888 8094 1912
rect 8012 1854 8036 1888
rect 8070 1854 8094 1888
rect 8012 1830 8094 1854
rect 9030 1888 9112 1912
rect 9030 1854 9054 1888
rect 9088 1854 9112 1888
rect 9030 1830 9112 1854
rect 10048 1888 10130 1912
rect 10048 1854 10072 1888
rect 10106 1854 10130 1888
rect 10048 1830 10130 1854
rect 11066 1888 11148 1912
rect 11066 1854 11090 1888
rect 11124 1854 11148 1888
rect 11066 1830 11148 1854
rect 13998 1538 14080 1562
rect 13998 1504 14022 1538
rect 14056 1504 14080 1538
rect 13998 1480 14080 1504
rect 15016 1538 15098 1562
rect 15016 1504 15040 1538
rect 15074 1504 15098 1538
rect 15016 1480 15098 1504
rect 16034 1538 16116 1562
rect 16034 1504 16058 1538
rect 16092 1504 16116 1538
rect 16034 1480 16116 1504
rect 17052 1538 17134 1562
rect 17052 1504 17076 1538
rect 17110 1504 17134 1538
rect 17052 1480 17134 1504
rect 18070 1538 18152 1562
rect 18070 1504 18094 1538
rect 18128 1504 18152 1538
rect 18070 1480 18152 1504
rect 19088 1538 19170 1562
rect 19088 1504 19112 1538
rect 19146 1504 19170 1538
rect 19088 1480 19170 1504
rect 20106 1538 20188 1562
rect 20106 1504 20130 1538
rect 20164 1504 20188 1538
rect 20106 1480 20188 1504
rect 21124 1538 21206 1562
rect 21124 1504 21148 1538
rect 21182 1504 21206 1538
rect 21124 1480 21206 1504
rect 22142 1538 22224 1562
rect 22142 1504 22166 1538
rect 22200 1504 22224 1538
rect 22142 1480 22224 1504
rect 23160 1538 23242 1562
rect 23160 1504 23184 1538
rect 23218 1504 23242 1538
rect 23160 1480 23242 1504
rect 24178 1538 24260 1562
rect 24178 1504 24202 1538
rect 24236 1504 24260 1538
rect 24178 1480 24260 1504
rect 25196 1538 25278 1562
rect 25196 1504 25220 1538
rect 25254 1504 25278 1538
rect 25196 1480 25278 1504
rect 26214 1538 26296 1562
rect 26214 1504 26238 1538
rect 26272 1504 26296 1538
rect 26214 1480 26296 1504
rect 27232 1538 27314 1562
rect 27232 1504 27256 1538
rect 27290 1504 27314 1538
rect 27232 1480 27314 1504
rect 28250 1538 28332 1562
rect 28250 1504 28274 1538
rect 28308 1504 28332 1538
rect 28250 1480 28332 1504
rect 29268 1538 29350 1562
rect 29268 1504 29292 1538
rect 29326 1504 29350 1538
rect 29268 1480 29350 1504
rect 30286 1538 30368 1562
rect 30286 1504 30310 1538
rect 30344 1504 30368 1538
rect 30286 1480 30368 1504
rect 31304 1538 31386 1562
rect 31304 1504 31328 1538
rect 31362 1504 31386 1538
rect 31304 1480 31386 1504
rect 32322 1538 32404 1562
rect 32322 1504 32346 1538
rect 32380 1504 32404 1538
rect 32322 1480 32404 1504
rect 33340 1538 33422 1562
rect 33340 1504 33364 1538
rect 33398 1504 33422 1538
rect 33340 1480 33422 1504
rect 696 442 778 466
rect 696 408 720 442
rect 754 408 778 442
rect 696 384 778 408
rect 1714 442 1796 466
rect 1714 408 1738 442
rect 1772 408 1796 442
rect 1714 384 1796 408
rect 2732 442 2814 466
rect 2732 408 2756 442
rect 2790 408 2814 442
rect 2732 384 2814 408
rect 3750 442 3832 466
rect 3750 408 3774 442
rect 3808 408 3832 442
rect 3750 384 3832 408
rect 4768 442 4850 466
rect 4768 408 4792 442
rect 4826 408 4850 442
rect 4768 384 4850 408
rect 5786 442 5868 466
rect 5786 408 5810 442
rect 5844 408 5868 442
rect 5786 384 5868 408
rect 6804 442 6886 466
rect 6804 408 6828 442
rect 6862 408 6886 442
rect 6804 384 6886 408
rect 7822 442 7904 466
rect 7822 408 7846 442
rect 7880 408 7904 442
rect 7822 384 7904 408
rect 8840 442 8922 466
rect 8840 408 8864 442
rect 8898 408 8922 442
rect 8840 384 8922 408
rect 9858 442 9940 466
rect 9858 408 9882 442
rect 9916 408 9940 442
rect 9858 384 9940 408
rect 10876 442 10958 466
rect 10876 408 10900 442
rect 10934 408 10958 442
rect 10876 384 10958 408
rect 13986 360 14068 384
rect 13986 326 14010 360
rect 14044 326 14068 360
rect 13986 302 14068 326
rect 15004 360 15086 384
rect 15004 326 15028 360
rect 15062 326 15086 360
rect 15004 302 15086 326
rect 16022 360 16104 384
rect 16022 326 16046 360
rect 16080 326 16104 360
rect 16022 302 16104 326
rect 17040 360 17122 384
rect 17040 326 17064 360
rect 17098 326 17122 360
rect 17040 302 17122 326
rect 18058 360 18140 384
rect 18058 326 18082 360
rect 18116 326 18140 360
rect 18058 302 18140 326
rect 19076 360 19158 384
rect 19076 326 19100 360
rect 19134 326 19158 360
rect 19076 302 19158 326
rect 20094 360 20176 384
rect 20094 326 20118 360
rect 20152 326 20176 360
rect 20094 302 20176 326
rect 21112 360 21194 384
rect 21112 326 21136 360
rect 21170 326 21194 360
rect 21112 302 21194 326
rect 22130 360 22212 384
rect 22130 326 22154 360
rect 22188 326 22212 360
rect 22130 302 22212 326
rect 23148 360 23230 384
rect 23148 326 23172 360
rect 23206 326 23230 360
rect 23148 302 23230 326
rect 24166 360 24248 384
rect 24166 326 24190 360
rect 24224 326 24248 360
rect 24166 302 24248 326
rect 25184 360 25266 384
rect 25184 326 25208 360
rect 25242 326 25266 360
rect 25184 302 25266 326
rect 26202 360 26284 384
rect 26202 326 26226 360
rect 26260 326 26284 360
rect 26202 302 26284 326
rect 27220 360 27302 384
rect 27220 326 27244 360
rect 27278 326 27302 360
rect 27220 302 27302 326
rect 28238 360 28320 384
rect 28238 326 28262 360
rect 28296 326 28320 360
rect 28238 302 28320 326
rect 29256 360 29338 384
rect 29256 326 29280 360
rect 29314 326 29338 360
rect 29256 302 29338 326
rect 30274 360 30356 384
rect 30274 326 30298 360
rect 30332 326 30356 360
rect 30274 302 30356 326
rect 31292 360 31374 384
rect 31292 326 31316 360
rect 31350 326 31374 360
rect 31292 302 31374 326
rect 32310 360 32392 384
rect 32310 326 32334 360
rect 32368 326 32392 360
rect 32310 302 32392 326
rect 33328 360 33410 384
rect 33328 326 33352 360
rect 33386 326 33410 360
rect 33328 302 33410 326
rect -1410 -582 -1310 -520
rect 35734 -582 35834 -520
rect -1410 -682 -1248 -582
rect 35672 -682 35834 -582
<< nsubdiff >>
rect 11290 30762 11452 30862
rect 35572 30762 35734 30862
rect 11290 30700 11390 30762
rect 35634 30700 35734 30762
rect 17884 28318 17966 28344
rect 17884 28284 17908 28318
rect 17942 28284 17966 28318
rect 17884 28260 17966 28284
rect 18902 28318 18984 28344
rect 18902 28284 18926 28318
rect 18960 28284 18984 28318
rect 18902 28260 18984 28284
rect 19920 28318 20002 28344
rect 19920 28284 19944 28318
rect 19978 28284 20002 28318
rect 19920 28260 20002 28284
rect 20938 28318 21020 28344
rect 20938 28284 20962 28318
rect 20996 28284 21020 28318
rect 20938 28260 21020 28284
rect 21956 28318 22038 28344
rect 21956 28284 21980 28318
rect 22014 28284 22038 28318
rect 21956 28260 22038 28284
rect 22974 28318 23056 28344
rect 22974 28284 22998 28318
rect 23032 28284 23056 28318
rect 22974 28260 23056 28284
rect 23992 28318 24074 28344
rect 23992 28284 24016 28318
rect 24050 28284 24074 28318
rect 23992 28260 24074 28284
rect 25010 28318 25092 28344
rect 25010 28284 25034 28318
rect 25068 28284 25092 28318
rect 25010 28260 25092 28284
rect 26028 28318 26110 28344
rect 26028 28284 26052 28318
rect 26086 28284 26110 28318
rect 26028 28260 26110 28284
rect 27046 28318 27128 28344
rect 27046 28284 27070 28318
rect 27104 28284 27128 28318
rect 27046 28260 27128 28284
rect 28064 28318 28146 28344
rect 28064 28284 28088 28318
rect 28122 28284 28146 28318
rect 28064 28260 28146 28284
rect 29082 28318 29164 28344
rect 29082 28284 29106 28318
rect 29140 28284 29164 28318
rect 29082 28260 29164 28284
rect 30100 28318 30182 28344
rect 30100 28284 30124 28318
rect 30158 28284 30182 28318
rect 30100 28260 30182 28284
rect 31118 28318 31200 28344
rect 31118 28284 31142 28318
rect 31176 28284 31200 28318
rect 31118 28260 31200 28284
rect 32136 28318 32218 28344
rect 32136 28284 32160 28318
rect 32194 28284 32218 28318
rect 32136 28260 32218 28284
rect 33154 28318 33236 28344
rect 33154 28284 33178 28318
rect 33212 28284 33236 28318
rect 33154 28260 33236 28284
rect 17906 27164 17988 27190
rect 17906 27130 17930 27164
rect 17964 27130 17988 27164
rect 17906 27106 17988 27130
rect 18924 27164 19006 27190
rect 18924 27130 18948 27164
rect 18982 27130 19006 27164
rect 18924 27106 19006 27130
rect 19942 27164 20024 27190
rect 19942 27130 19966 27164
rect 20000 27130 20024 27164
rect 19942 27106 20024 27130
rect 20960 27164 21042 27190
rect 20960 27130 20984 27164
rect 21018 27130 21042 27164
rect 20960 27106 21042 27130
rect 21978 27164 22060 27190
rect 21978 27130 22002 27164
rect 22036 27130 22060 27164
rect 21978 27106 22060 27130
rect 22996 27164 23078 27190
rect 22996 27130 23020 27164
rect 23054 27130 23078 27164
rect 22996 27106 23078 27130
rect 24014 27164 24096 27190
rect 24014 27130 24038 27164
rect 24072 27130 24096 27164
rect 24014 27106 24096 27130
rect 25032 27164 25114 27190
rect 25032 27130 25056 27164
rect 25090 27130 25114 27164
rect 25032 27106 25114 27130
rect 26050 27164 26132 27190
rect 26050 27130 26074 27164
rect 26108 27130 26132 27164
rect 26050 27106 26132 27130
rect 27068 27164 27150 27190
rect 27068 27130 27092 27164
rect 27126 27130 27150 27164
rect 27068 27106 27150 27130
rect 28086 27164 28168 27190
rect 28086 27130 28110 27164
rect 28144 27130 28168 27164
rect 28086 27106 28168 27130
rect 29104 27164 29186 27190
rect 29104 27130 29128 27164
rect 29162 27130 29186 27164
rect 29104 27106 29186 27130
rect 30122 27164 30204 27190
rect 30122 27130 30146 27164
rect 30180 27130 30204 27164
rect 30122 27106 30204 27130
rect 31140 27164 31222 27190
rect 31140 27130 31164 27164
rect 31198 27130 31222 27164
rect 31140 27106 31222 27130
rect 32158 27164 32240 27190
rect 32158 27130 32182 27164
rect 32216 27130 32240 27164
rect 32158 27106 32240 27130
rect 33176 27164 33258 27190
rect 33176 27130 33200 27164
rect 33234 27130 33258 27164
rect 33176 27106 33258 27130
rect 17884 26032 17966 26058
rect 17884 25998 17908 26032
rect 17942 25998 17966 26032
rect 17884 25974 17966 25998
rect 18902 26032 18984 26058
rect 18902 25998 18926 26032
rect 18960 25998 18984 26032
rect 18902 25974 18984 25998
rect 19920 26032 20002 26058
rect 19920 25998 19944 26032
rect 19978 25998 20002 26032
rect 19920 25974 20002 25998
rect 20938 26032 21020 26058
rect 20938 25998 20962 26032
rect 20996 25998 21020 26032
rect 20938 25974 21020 25998
rect 21956 26032 22038 26058
rect 21956 25998 21980 26032
rect 22014 25998 22038 26032
rect 21956 25974 22038 25998
rect 22974 26032 23056 26058
rect 22974 25998 22998 26032
rect 23032 25998 23056 26032
rect 22974 25974 23056 25998
rect 23992 26032 24074 26058
rect 23992 25998 24016 26032
rect 24050 25998 24074 26032
rect 23992 25974 24074 25998
rect 25010 26032 25092 26058
rect 25010 25998 25034 26032
rect 25068 25998 25092 26032
rect 25010 25974 25092 25998
rect 26028 26032 26110 26058
rect 26028 25998 26052 26032
rect 26086 25998 26110 26032
rect 26028 25974 26110 25998
rect 27046 26032 27128 26058
rect 27046 25998 27070 26032
rect 27104 25998 27128 26032
rect 27046 25974 27128 25998
rect 28064 26032 28146 26058
rect 28064 25998 28088 26032
rect 28122 25998 28146 26032
rect 28064 25974 28146 25998
rect 29082 26032 29164 26058
rect 29082 25998 29106 26032
rect 29140 25998 29164 26032
rect 29082 25974 29164 25998
rect 30100 26032 30182 26058
rect 30100 25998 30124 26032
rect 30158 25998 30182 26032
rect 30100 25974 30182 25998
rect 31118 26032 31200 26058
rect 31118 25998 31142 26032
rect 31176 25998 31200 26032
rect 31118 25974 31200 25998
rect 32136 26032 32218 26058
rect 32136 25998 32160 26032
rect 32194 25998 32218 26032
rect 32136 25974 32218 25998
rect 33154 26032 33236 26058
rect 33154 25998 33178 26032
rect 33212 25998 33236 26032
rect 33154 25974 33236 25998
rect 17884 24650 17966 24676
rect 17884 24616 17908 24650
rect 17942 24616 17966 24650
rect 17884 24592 17966 24616
rect 18902 24650 18984 24676
rect 18902 24616 18926 24650
rect 18960 24616 18984 24650
rect 18902 24592 18984 24616
rect 19920 24650 20002 24676
rect 19920 24616 19944 24650
rect 19978 24616 20002 24650
rect 19920 24592 20002 24616
rect 20938 24650 21020 24676
rect 20938 24616 20962 24650
rect 20996 24616 21020 24650
rect 20938 24592 21020 24616
rect 21956 24650 22038 24676
rect 21956 24616 21980 24650
rect 22014 24616 22038 24650
rect 21956 24592 22038 24616
rect 22974 24650 23056 24676
rect 22974 24616 22998 24650
rect 23032 24616 23056 24650
rect 22974 24592 23056 24616
rect 23992 24650 24074 24676
rect 23992 24616 24016 24650
rect 24050 24616 24074 24650
rect 23992 24592 24074 24616
rect 25010 24650 25092 24676
rect 25010 24616 25034 24650
rect 25068 24616 25092 24650
rect 25010 24592 25092 24616
rect 26028 24650 26110 24676
rect 26028 24616 26052 24650
rect 26086 24616 26110 24650
rect 26028 24592 26110 24616
rect 27046 24650 27128 24676
rect 27046 24616 27070 24650
rect 27104 24616 27128 24650
rect 27046 24592 27128 24616
rect 28064 24650 28146 24676
rect 28064 24616 28088 24650
rect 28122 24616 28146 24650
rect 28064 24592 28146 24616
rect 29082 24650 29164 24676
rect 29082 24616 29106 24650
rect 29140 24616 29164 24650
rect 29082 24592 29164 24616
rect 30100 24650 30182 24676
rect 30100 24616 30124 24650
rect 30158 24616 30182 24650
rect 30100 24592 30182 24616
rect 31118 24650 31200 24676
rect 31118 24616 31142 24650
rect 31176 24616 31200 24650
rect 31118 24592 31200 24616
rect 32136 24650 32218 24676
rect 32136 24616 32160 24650
rect 32194 24616 32218 24650
rect 32136 24592 32218 24616
rect 33154 24650 33236 24676
rect 33154 24616 33178 24650
rect 33212 24616 33236 24650
rect 33154 24592 33236 24616
rect 18572 23302 18654 23328
rect 18572 23268 18596 23302
rect 18630 23268 18654 23302
rect 18572 23244 18654 23268
rect 19590 23302 19672 23328
rect 19590 23268 19614 23302
rect 19648 23268 19672 23302
rect 19590 23244 19672 23268
rect 20608 23302 20690 23328
rect 20608 23268 20632 23302
rect 20666 23268 20690 23302
rect 20608 23244 20690 23268
rect 21626 23302 21708 23328
rect 21626 23268 21650 23302
rect 21684 23268 21708 23302
rect 21626 23244 21708 23268
rect 22644 23302 22726 23328
rect 22644 23268 22668 23302
rect 22702 23268 22726 23302
rect 22644 23244 22726 23268
rect 23662 23302 23744 23328
rect 23662 23268 23686 23302
rect 23720 23268 23744 23302
rect 23662 23244 23744 23268
rect 24680 23302 24762 23328
rect 24680 23268 24704 23302
rect 24738 23268 24762 23302
rect 24680 23244 24762 23268
rect 25698 23302 25780 23328
rect 25698 23268 25722 23302
rect 25756 23268 25780 23302
rect 25698 23244 25780 23268
rect 26716 23302 26798 23328
rect 26716 23268 26740 23302
rect 26774 23268 26798 23302
rect 26716 23244 26798 23268
rect 27734 23302 27816 23328
rect 27734 23268 27758 23302
rect 27792 23268 27816 23302
rect 27734 23244 27816 23268
rect 28752 23302 28834 23328
rect 28752 23268 28776 23302
rect 28810 23268 28834 23302
rect 28752 23244 28834 23268
rect 29770 23302 29852 23328
rect 29770 23268 29794 23302
rect 29828 23268 29852 23302
rect 29770 23244 29852 23268
rect 30788 23302 30870 23328
rect 30788 23268 30812 23302
rect 30846 23268 30870 23302
rect 30788 23244 30870 23268
rect 31806 23302 31888 23328
rect 31806 23268 31830 23302
rect 31864 23268 31888 23302
rect 31806 23244 31888 23268
rect 32824 23302 32906 23328
rect 32824 23268 32848 23302
rect 32882 23268 32906 23302
rect 32824 23244 32906 23268
rect 18178 22024 18260 22050
rect 18178 21990 18202 22024
rect 18236 21990 18260 22024
rect 18178 21966 18260 21990
rect 19196 22024 19278 22050
rect 19196 21990 19220 22024
rect 19254 21990 19278 22024
rect 19196 21966 19278 21990
rect 20214 22024 20296 22050
rect 20214 21990 20238 22024
rect 20272 21990 20296 22024
rect 20214 21966 20296 21990
rect 21232 22024 21314 22050
rect 21232 21990 21256 22024
rect 21290 21990 21314 22024
rect 21232 21966 21314 21990
rect 22250 22024 22332 22050
rect 22250 21990 22274 22024
rect 22308 21990 22332 22024
rect 22250 21966 22332 21990
rect 23268 22024 23350 22050
rect 23268 21990 23292 22024
rect 23326 21990 23350 22024
rect 23268 21966 23350 21990
rect 24286 22024 24368 22050
rect 24286 21990 24310 22024
rect 24344 21990 24368 22024
rect 24286 21966 24368 21990
rect 25304 22024 25386 22050
rect 25304 21990 25328 22024
rect 25362 21990 25386 22024
rect 25304 21966 25386 21990
rect 26322 22024 26404 22050
rect 26322 21990 26346 22024
rect 26380 21990 26404 22024
rect 26322 21966 26404 21990
rect 27340 22024 27422 22050
rect 27340 21990 27364 22024
rect 27398 21990 27422 22024
rect 27340 21966 27422 21990
rect 28358 22024 28440 22050
rect 28358 21990 28382 22024
rect 28416 21990 28440 22024
rect 28358 21966 28440 21990
rect 29376 22024 29458 22050
rect 29376 21990 29400 22024
rect 29434 21990 29458 22024
rect 29376 21966 29458 21990
rect 30394 22024 30476 22050
rect 30394 21990 30418 22024
rect 30452 21990 30476 22024
rect 30394 21966 30476 21990
rect 31412 22024 31494 22050
rect 31412 21990 31436 22024
rect 31470 21990 31494 22024
rect 31412 21966 31494 21990
rect 32430 22024 32512 22050
rect 32430 21990 32454 22024
rect 32488 21990 32512 22024
rect 32430 21966 32512 21990
rect 33448 22024 33530 22050
rect 33448 21990 33472 22024
rect 33506 21990 33530 22024
rect 33448 21966 33530 21990
rect 13580 21714 13662 21740
rect 13580 21680 13604 21714
rect 13638 21680 13662 21714
rect 13580 21656 13662 21680
rect 14598 21714 14680 21740
rect 14598 21680 14622 21714
rect 14656 21680 14680 21714
rect 14598 21656 14680 21680
rect 15616 21714 15698 21740
rect 15616 21680 15640 21714
rect 15674 21680 15698 21714
rect 15616 21656 15698 21680
rect 16634 21714 16716 21740
rect 16634 21680 16658 21714
rect 16692 21680 16716 21714
rect 16634 21656 16716 21680
rect 13056 20560 13138 20586
rect 13056 20526 13080 20560
rect 13114 20526 13138 20560
rect 13056 20502 13138 20526
rect 14074 20560 14156 20586
rect 14074 20526 14098 20560
rect 14132 20526 14156 20560
rect 14074 20502 14156 20526
rect 15092 20560 15174 20586
rect 15092 20526 15116 20560
rect 15150 20526 15174 20560
rect 15092 20502 15174 20526
rect 16110 20560 16192 20586
rect 16110 20526 16134 20560
rect 16168 20526 16192 20560
rect 16110 20502 16192 20526
rect 18268 20576 18350 20602
rect 18268 20542 18292 20576
rect 18326 20542 18350 20576
rect 18268 20518 18350 20542
rect 19286 20576 19368 20602
rect 19286 20542 19310 20576
rect 19344 20542 19368 20576
rect 19286 20518 19368 20542
rect 20304 20576 20386 20602
rect 20304 20542 20328 20576
rect 20362 20542 20386 20576
rect 20304 20518 20386 20542
rect 21322 20576 21404 20602
rect 21322 20542 21346 20576
rect 21380 20542 21404 20576
rect 21322 20518 21404 20542
rect 22340 20576 22422 20602
rect 22340 20542 22364 20576
rect 22398 20542 22422 20576
rect 22340 20518 22422 20542
rect 23358 20576 23440 20602
rect 23358 20542 23382 20576
rect 23416 20542 23440 20576
rect 23358 20518 23440 20542
rect 24376 20576 24458 20602
rect 24376 20542 24400 20576
rect 24434 20542 24458 20576
rect 24376 20518 24458 20542
rect 25394 20576 25476 20602
rect 25394 20542 25418 20576
rect 25452 20542 25476 20576
rect 25394 20518 25476 20542
rect 26412 20576 26494 20602
rect 26412 20542 26436 20576
rect 26470 20542 26494 20576
rect 26412 20518 26494 20542
rect 27430 20576 27512 20602
rect 27430 20542 27454 20576
rect 27488 20542 27512 20576
rect 27430 20518 27512 20542
rect 28448 20576 28530 20602
rect 28448 20542 28472 20576
rect 28506 20542 28530 20576
rect 28448 20518 28530 20542
rect 29466 20576 29548 20602
rect 29466 20542 29490 20576
rect 29524 20542 29548 20576
rect 29466 20518 29548 20542
rect 30484 20576 30566 20602
rect 30484 20542 30508 20576
rect 30542 20542 30566 20576
rect 30484 20518 30566 20542
rect 31502 20576 31584 20602
rect 31502 20542 31526 20576
rect 31560 20542 31584 20576
rect 31502 20518 31584 20542
rect 32520 20576 32602 20602
rect 32520 20542 32544 20576
rect 32578 20542 32602 20576
rect 32520 20518 32602 20542
rect 33538 20576 33620 20602
rect 33538 20542 33562 20576
rect 33596 20542 33620 20576
rect 33538 20518 33620 20542
rect 13066 19532 13148 19558
rect 13066 19498 13090 19532
rect 13124 19498 13148 19532
rect 13066 19474 13148 19498
rect 14084 19532 14166 19558
rect 14084 19498 14108 19532
rect 14142 19498 14166 19532
rect 14084 19474 14166 19498
rect 15102 19532 15184 19558
rect 15102 19498 15126 19532
rect 15160 19498 15184 19532
rect 15102 19474 15184 19498
rect 16120 19532 16202 19558
rect 16120 19498 16144 19532
rect 16178 19498 16202 19532
rect 16120 19474 16202 19498
rect 18292 19308 18374 19334
rect 18292 19274 18316 19308
rect 18350 19274 18374 19308
rect 18292 19250 18374 19274
rect 19310 19308 19392 19334
rect 19310 19274 19334 19308
rect 19368 19274 19392 19308
rect 19310 19250 19392 19274
rect 20328 19308 20410 19334
rect 20328 19274 20352 19308
rect 20386 19274 20410 19308
rect 20328 19250 20410 19274
rect 21346 19308 21428 19334
rect 21346 19274 21370 19308
rect 21404 19274 21428 19308
rect 21346 19250 21428 19274
rect 22364 19308 22446 19334
rect 22364 19274 22388 19308
rect 22422 19274 22446 19308
rect 22364 19250 22446 19274
rect 23382 19308 23464 19334
rect 23382 19274 23406 19308
rect 23440 19274 23464 19308
rect 23382 19250 23464 19274
rect 24400 19308 24482 19334
rect 24400 19274 24424 19308
rect 24458 19274 24482 19308
rect 24400 19250 24482 19274
rect 25418 19308 25500 19334
rect 25418 19274 25442 19308
rect 25476 19274 25500 19308
rect 25418 19250 25500 19274
rect 26436 19308 26518 19334
rect 26436 19274 26460 19308
rect 26494 19274 26518 19308
rect 26436 19250 26518 19274
rect 27454 19308 27536 19334
rect 27454 19274 27478 19308
rect 27512 19274 27536 19308
rect 27454 19250 27536 19274
rect 28472 19308 28554 19334
rect 28472 19274 28496 19308
rect 28530 19274 28554 19308
rect 28472 19250 28554 19274
rect 29490 19308 29572 19334
rect 29490 19274 29514 19308
rect 29548 19274 29572 19308
rect 29490 19250 29572 19274
rect 30508 19308 30590 19334
rect 30508 19274 30532 19308
rect 30566 19274 30590 19308
rect 30508 19250 30590 19274
rect 31526 19308 31608 19334
rect 31526 19274 31550 19308
rect 31584 19274 31608 19308
rect 31526 19250 31608 19274
rect 32544 19308 32626 19334
rect 32544 19274 32568 19308
rect 32602 19274 32626 19308
rect 32544 19250 32626 19274
rect 33562 19308 33644 19334
rect 33562 19274 33586 19308
rect 33620 19274 33644 19308
rect 33562 19250 33644 19274
rect 13056 18504 13138 18530
rect 13056 18470 13080 18504
rect 13114 18470 13138 18504
rect 13056 18446 13138 18470
rect 14074 18504 14156 18530
rect 14074 18470 14098 18504
rect 14132 18470 14156 18504
rect 14074 18446 14156 18470
rect 15092 18504 15174 18530
rect 15092 18470 15116 18504
rect 15150 18470 15174 18504
rect 15092 18446 15174 18470
rect 16110 18504 16192 18530
rect 16110 18470 16134 18504
rect 16168 18470 16192 18504
rect 16110 18446 16192 18470
rect 18156 18064 18238 18090
rect 18156 18030 18180 18064
rect 18214 18030 18238 18064
rect 18156 18006 18238 18030
rect 19174 18064 19256 18090
rect 19174 18030 19198 18064
rect 19232 18030 19256 18064
rect 19174 18006 19256 18030
rect 20192 18064 20274 18090
rect 20192 18030 20216 18064
rect 20250 18030 20274 18064
rect 20192 18006 20274 18030
rect 21210 18064 21292 18090
rect 21210 18030 21234 18064
rect 21268 18030 21292 18064
rect 21210 18006 21292 18030
rect 22228 18064 22310 18090
rect 22228 18030 22252 18064
rect 22286 18030 22310 18064
rect 22228 18006 22310 18030
rect 23246 18064 23328 18090
rect 23246 18030 23270 18064
rect 23304 18030 23328 18064
rect 23246 18006 23328 18030
rect 24264 18064 24346 18090
rect 24264 18030 24288 18064
rect 24322 18030 24346 18064
rect 24264 18006 24346 18030
rect 25282 18064 25364 18090
rect 25282 18030 25306 18064
rect 25340 18030 25364 18064
rect 25282 18006 25364 18030
rect 26300 18064 26382 18090
rect 26300 18030 26324 18064
rect 26358 18030 26382 18064
rect 26300 18006 26382 18030
rect 27318 18064 27400 18090
rect 27318 18030 27342 18064
rect 27376 18030 27400 18064
rect 27318 18006 27400 18030
rect 28336 18064 28418 18090
rect 28336 18030 28360 18064
rect 28394 18030 28418 18064
rect 28336 18006 28418 18030
rect 29354 18064 29436 18090
rect 29354 18030 29378 18064
rect 29412 18030 29436 18064
rect 29354 18006 29436 18030
rect 30372 18064 30454 18090
rect 30372 18030 30396 18064
rect 30430 18030 30454 18064
rect 30372 18006 30454 18030
rect 31390 18064 31472 18090
rect 31390 18030 31414 18064
rect 31448 18030 31472 18064
rect 31390 18006 31472 18030
rect 32408 18064 32490 18090
rect 32408 18030 32432 18064
rect 32466 18030 32490 18064
rect 32408 18006 32490 18030
rect 33426 18064 33508 18090
rect 33426 18030 33450 18064
rect 33484 18030 33508 18064
rect 33426 18006 33508 18030
rect 13580 17352 13662 17378
rect 13580 17318 13604 17352
rect 13638 17318 13662 17352
rect 13580 17294 13662 17318
rect 14598 17352 14680 17378
rect 14598 17318 14622 17352
rect 14656 17318 14680 17352
rect 14598 17294 14680 17318
rect 15616 17352 15698 17378
rect 15616 17318 15640 17352
rect 15674 17318 15698 17352
rect 15616 17294 15698 17318
rect 16634 17352 16716 17378
rect 16634 17318 16658 17352
rect 16692 17318 16716 17352
rect 16634 17294 16716 17318
rect -12280 16275 -12184 16309
rect -10566 16275 -10470 16309
rect -12280 16213 -12246 16275
rect -10504 16213 -10470 16275
rect -12280 15577 -12246 15639
rect -9680 16275 -9584 16309
rect -7966 16275 -7870 16309
rect -9680 16213 -9646 16275
rect -10504 15577 -10470 15639
rect -12280 15543 -12184 15577
rect -10566 15543 -10470 15577
rect -7904 16213 -7870 16275
rect -9680 15577 -9646 15639
rect 11290 16292 11390 16354
rect 35634 16292 35734 16354
rect 11290 16192 11452 16292
rect 35572 16192 35734 16292
rect -7904 15577 -7870 15639
rect -9680 15543 -9584 15577
rect -7966 15543 -7870 15577
<< psubdiffcont >>
rect -12184 15342 -10566 15376
rect -12280 14924 -12246 15280
rect -9584 15342 -7966 15376
rect -10504 14924 -10470 15280
rect -12184 14828 -10566 14862
rect -9680 14924 -9646 15280
rect -7904 14924 -7870 15280
rect -9584 14828 -7966 14862
rect -1248 15262 35672 15362
rect -1410 -520 -1310 15200
rect 14022 14722 14056 14756
rect 15040 14722 15074 14756
rect 16058 14722 16092 14756
rect 17076 14722 17110 14756
rect 18094 14722 18128 14756
rect 19112 14722 19146 14756
rect 20130 14722 20164 14756
rect 21148 14722 21182 14756
rect 22166 14722 22200 14756
rect 23184 14722 23218 14756
rect 24202 14722 24236 14756
rect 25220 14722 25254 14756
rect 26238 14722 26272 14756
rect 27256 14722 27290 14756
rect 28274 14722 28308 14756
rect 29292 14722 29326 14756
rect 30310 14722 30344 14756
rect 31328 14722 31362 14756
rect 32346 14722 32380 14756
rect 33364 14722 33398 14756
rect 1728 14120 1762 14154
rect 2746 14120 2780 14154
rect 3764 14120 3798 14154
rect 4782 14120 4816 14154
rect 5800 14120 5834 14154
rect 6818 14120 6852 14154
rect 7836 14120 7870 14154
rect 8854 14120 8888 14154
rect 9872 14120 9906 14154
rect 10900 14120 10934 14154
rect 1728 13302 1762 13336
rect 2746 13302 2780 13336
rect 3764 13302 3798 13336
rect 4782 13302 4816 13336
rect 5800 13302 5834 13336
rect 6818 13302 6852 13336
rect 7836 13302 7870 13336
rect 8854 13302 8888 13336
rect 9872 13302 9906 13336
rect 10900 13302 10934 13336
rect 14034 12696 14068 12730
rect 15052 12696 15086 12730
rect 16070 12696 16104 12730
rect 17088 12696 17122 12730
rect 18106 12696 18140 12730
rect 19124 12696 19158 12730
rect 20142 12696 20176 12730
rect 21160 12696 21194 12730
rect 22178 12696 22212 12730
rect 23196 12696 23230 12730
rect 24214 12696 24248 12730
rect 25232 12696 25266 12730
rect 26250 12696 26284 12730
rect 27268 12696 27302 12730
rect 28286 12696 28320 12730
rect 29304 12696 29338 12730
rect 30322 12696 30356 12730
rect 31340 12696 31374 12730
rect 32358 12696 32392 12730
rect 33376 12696 33410 12730
rect 1728 12484 1762 12518
rect 2746 12484 2780 12518
rect 3764 12484 3798 12518
rect 4782 12484 4816 12518
rect 5800 12484 5834 12518
rect 6818 12484 6852 12518
rect 7836 12484 7870 12518
rect 8854 12484 8888 12518
rect 9872 12484 9906 12518
rect 10900 12484 10934 12518
rect 1728 11666 1762 11700
rect 2746 11666 2780 11700
rect 3764 11666 3798 11700
rect 4782 11666 4816 11700
rect 5800 11666 5834 11700
rect 6818 11666 6852 11700
rect 7836 11666 7870 11700
rect 8854 11666 8888 11700
rect 9872 11666 9906 11700
rect 10900 11666 10934 11700
rect 14022 11390 14056 11424
rect 15040 11390 15074 11424
rect 16058 11390 16092 11424
rect 17076 11390 17110 11424
rect 18094 11390 18128 11424
rect 19112 11390 19146 11424
rect 20130 11390 20164 11424
rect 21148 11390 21182 11424
rect 22166 11390 22200 11424
rect 23184 11390 23218 11424
rect 24202 11390 24236 11424
rect 25220 11390 25254 11424
rect 26238 11390 26272 11424
rect 27256 11390 27290 11424
rect 28274 11390 28308 11424
rect 29292 11390 29326 11424
rect 30310 11390 30344 11424
rect 31328 11390 31362 11424
rect 32346 11390 32380 11424
rect 33364 11390 33398 11424
rect 1728 10848 1762 10882
rect 2746 10848 2780 10882
rect 3764 10848 3798 10882
rect 4782 10848 4816 10882
rect 5800 10848 5834 10882
rect 6818 10848 6852 10882
rect 7836 10848 7870 10882
rect 8854 10848 8888 10882
rect 9872 10848 9906 10882
rect 10900 10848 10934 10882
rect 1728 10030 1762 10064
rect 2746 10030 2780 10064
rect 3764 10030 3798 10064
rect 4782 10030 4816 10064
rect 5800 10030 5834 10064
rect 6818 10030 6852 10064
rect 7836 10030 7870 10064
rect 14010 10154 14044 10188
rect 15028 10154 15062 10188
rect 16046 10154 16080 10188
rect 17064 10154 17098 10188
rect 18082 10154 18116 10188
rect 19100 10154 19134 10188
rect 20118 10154 20152 10188
rect 21136 10154 21170 10188
rect 22154 10154 22188 10188
rect 23172 10154 23206 10188
rect 24190 10154 24224 10188
rect 25208 10154 25242 10188
rect 26226 10154 26260 10188
rect 27244 10154 27278 10188
rect 28262 10154 28296 10188
rect 29280 10154 29314 10188
rect 30298 10154 30332 10188
rect 31316 10154 31350 10188
rect 32334 10154 32368 10188
rect 33352 10154 33386 10188
rect 8854 10030 8888 10064
rect 9872 10030 9906 10064
rect 10900 10030 10934 10064
rect 1728 9212 1762 9246
rect 2746 9212 2780 9246
rect 3764 9212 3798 9246
rect 4782 9212 4816 9246
rect 5800 9212 5834 9246
rect 6818 9212 6852 9246
rect 7836 9212 7870 9246
rect 8854 9212 8888 9246
rect 9872 9212 9906 9246
rect 10900 9212 10934 9246
rect 14010 8930 14044 8964
rect 15028 8930 15062 8964
rect 16046 8930 16080 8964
rect 17064 8930 17098 8964
rect 18082 8930 18116 8964
rect 19100 8930 19134 8964
rect 20118 8930 20152 8964
rect 21136 8930 21170 8964
rect 22154 8930 22188 8964
rect 23172 8930 23206 8964
rect 24190 8930 24224 8964
rect 25208 8930 25242 8964
rect 26226 8930 26260 8964
rect 27244 8930 27278 8964
rect 28262 8930 28296 8964
rect 29280 8930 29314 8964
rect 30298 8930 30332 8964
rect 31316 8930 31350 8964
rect 32334 8930 32368 8964
rect 33352 8930 33386 8964
rect 1728 8394 1762 8428
rect 2746 8394 2780 8428
rect 3764 8394 3798 8428
rect 4782 8394 4816 8428
rect 5800 8394 5834 8428
rect 6818 8394 6852 8428
rect 7836 8394 7870 8428
rect 8854 8394 8888 8428
rect 9872 8394 9906 8428
rect 10900 8394 10934 8428
rect 14022 7694 14056 7728
rect 15040 7694 15074 7728
rect 16058 7694 16092 7728
rect 17076 7694 17110 7728
rect 18094 7694 18128 7728
rect 19112 7694 19146 7728
rect 20130 7694 20164 7728
rect 21148 7694 21182 7728
rect 22166 7694 22200 7728
rect 23184 7694 23218 7728
rect 24202 7694 24236 7728
rect 25220 7694 25254 7728
rect 26238 7694 26272 7728
rect 27256 7694 27290 7728
rect 28274 7694 28308 7728
rect 29292 7694 29326 7728
rect 30310 7694 30344 7728
rect 31328 7694 31362 7728
rect 32346 7694 32380 7728
rect 33364 7694 33398 7728
rect 1716 7500 1750 7534
rect 2734 7500 2768 7534
rect 3752 7500 3786 7534
rect 4770 7500 4804 7534
rect 5788 7500 5822 7534
rect 6806 7500 6840 7534
rect 7824 7500 7858 7534
rect 8842 7500 8876 7534
rect 9860 7500 9894 7534
rect 10888 7500 10922 7534
rect 920 6552 954 6586
rect 1938 6552 1972 6586
rect 2956 6552 2990 6586
rect 3974 6552 4008 6586
rect 4992 6552 5026 6586
rect 6010 6552 6044 6586
rect 7028 6552 7062 6586
rect 8046 6552 8080 6586
rect 9064 6552 9098 6586
rect 10082 6552 10116 6586
rect 11100 6552 11134 6586
rect 14022 6446 14056 6480
rect 15040 6446 15074 6480
rect 16058 6446 16092 6480
rect 17076 6446 17110 6480
rect 18094 6446 18128 6480
rect 19112 6446 19146 6480
rect 20130 6446 20164 6480
rect 21148 6446 21182 6480
rect 22166 6446 22200 6480
rect 23184 6446 23218 6480
rect 24202 6446 24236 6480
rect 25220 6446 25254 6480
rect 26238 6446 26272 6480
rect 27256 6446 27290 6480
rect 28274 6446 28308 6480
rect 29292 6446 29326 6480
rect 30310 6446 30344 6480
rect 31328 6446 31362 6480
rect 32346 6446 32380 6480
rect 33364 6446 33398 6480
rect 932 5410 966 5444
rect 1950 5410 1984 5444
rect 2968 5410 3002 5444
rect 3986 5410 4020 5444
rect 5004 5410 5038 5444
rect 6022 5410 6056 5444
rect 7040 5410 7074 5444
rect 8058 5410 8092 5444
rect 9076 5410 9110 5444
rect 10094 5410 10128 5444
rect 11112 5410 11146 5444
rect 13998 5210 14032 5244
rect 15016 5210 15050 5244
rect 16034 5210 16068 5244
rect 17052 5210 17086 5244
rect 18070 5210 18104 5244
rect 19088 5210 19122 5244
rect 20106 5210 20140 5244
rect 21124 5210 21158 5244
rect 22142 5210 22176 5244
rect 23160 5210 23194 5244
rect 24178 5210 24212 5244
rect 25196 5210 25230 5244
rect 26214 5210 26248 5244
rect 27232 5210 27266 5244
rect 28250 5210 28284 5244
rect 29268 5210 29302 5244
rect 30286 5210 30320 5244
rect 31304 5210 31338 5244
rect 32322 5210 32356 5244
rect 33340 5210 33374 5244
rect 910 4302 944 4336
rect 1928 4302 1962 4336
rect 2946 4302 2980 4336
rect 3964 4302 3998 4336
rect 4982 4302 5016 4336
rect 6000 4302 6034 4336
rect 7018 4302 7052 4336
rect 8036 4302 8070 4336
rect 9054 4302 9088 4336
rect 10072 4302 10106 4336
rect 11090 4302 11124 4336
rect 14010 3986 14044 4020
rect 15028 3986 15062 4020
rect 16046 3986 16080 4020
rect 17064 3986 17098 4020
rect 18082 3986 18116 4020
rect 19100 3986 19134 4020
rect 20118 3986 20152 4020
rect 21136 3986 21170 4020
rect 22154 3986 22188 4020
rect 23172 3986 23206 4020
rect 24190 3986 24224 4020
rect 25208 3986 25242 4020
rect 26226 3986 26260 4020
rect 27244 3986 27278 4020
rect 28262 3986 28296 4020
rect 29280 3986 29314 4020
rect 30298 3986 30332 4020
rect 31316 3986 31350 4020
rect 32334 3986 32368 4020
rect 33352 3986 33386 4020
rect 910 3196 944 3230
rect 1928 3196 1962 3230
rect 2946 3196 2980 3230
rect 3964 3196 3998 3230
rect 4982 3196 5016 3230
rect 6000 3196 6034 3230
rect 7018 3196 7052 3230
rect 8036 3196 8070 3230
rect 9054 3196 9088 3230
rect 10072 3196 10106 3230
rect 11090 3196 11124 3230
rect 14010 2750 14044 2784
rect 15028 2750 15062 2784
rect 16046 2750 16080 2784
rect 17064 2750 17098 2784
rect 18082 2750 18116 2784
rect 19100 2750 19134 2784
rect 20118 2750 20152 2784
rect 21136 2750 21170 2784
rect 22154 2750 22188 2784
rect 23172 2750 23206 2784
rect 24190 2750 24224 2784
rect 25208 2750 25242 2784
rect 26226 2750 26260 2784
rect 27244 2750 27278 2784
rect 28262 2750 28296 2784
rect 29280 2750 29314 2784
rect 30298 2750 30332 2784
rect 31316 2750 31350 2784
rect 32334 2750 32368 2784
rect 33352 2750 33386 2784
rect 910 1854 944 1888
rect 1928 1854 1962 1888
rect 2946 1854 2980 1888
rect 3964 1854 3998 1888
rect 4982 1854 5016 1888
rect 6000 1854 6034 1888
rect 7018 1854 7052 1888
rect 8036 1854 8070 1888
rect 9054 1854 9088 1888
rect 10072 1854 10106 1888
rect 11090 1854 11124 1888
rect 14022 1504 14056 1538
rect 15040 1504 15074 1538
rect 16058 1504 16092 1538
rect 17076 1504 17110 1538
rect 18094 1504 18128 1538
rect 19112 1504 19146 1538
rect 20130 1504 20164 1538
rect 21148 1504 21182 1538
rect 22166 1504 22200 1538
rect 23184 1504 23218 1538
rect 24202 1504 24236 1538
rect 25220 1504 25254 1538
rect 26238 1504 26272 1538
rect 27256 1504 27290 1538
rect 28274 1504 28308 1538
rect 29292 1504 29326 1538
rect 30310 1504 30344 1538
rect 31328 1504 31362 1538
rect 32346 1504 32380 1538
rect 33364 1504 33398 1538
rect 720 408 754 442
rect 1738 408 1772 442
rect 2756 408 2790 442
rect 3774 408 3808 442
rect 4792 408 4826 442
rect 5810 408 5844 442
rect 6828 408 6862 442
rect 7846 408 7880 442
rect 8864 408 8898 442
rect 9882 408 9916 442
rect 10900 408 10934 442
rect 14010 326 14044 360
rect 15028 326 15062 360
rect 16046 326 16080 360
rect 17064 326 17098 360
rect 18082 326 18116 360
rect 19100 326 19134 360
rect 20118 326 20152 360
rect 21136 326 21170 360
rect 22154 326 22188 360
rect 23172 326 23206 360
rect 24190 326 24224 360
rect 25208 326 25242 360
rect 26226 326 26260 360
rect 27244 326 27278 360
rect 28262 326 28296 360
rect 29280 326 29314 360
rect 30298 326 30332 360
rect 31316 326 31350 360
rect 32334 326 32368 360
rect 33352 326 33386 360
rect 35734 -520 35834 15200
rect -1248 -682 35672 -582
<< nsubdiffcont >>
rect 11452 30762 35572 30862
rect 11290 16354 11390 30700
rect 17908 28284 17942 28318
rect 18926 28284 18960 28318
rect 19944 28284 19978 28318
rect 20962 28284 20996 28318
rect 21980 28284 22014 28318
rect 22998 28284 23032 28318
rect 24016 28284 24050 28318
rect 25034 28284 25068 28318
rect 26052 28284 26086 28318
rect 27070 28284 27104 28318
rect 28088 28284 28122 28318
rect 29106 28284 29140 28318
rect 30124 28284 30158 28318
rect 31142 28284 31176 28318
rect 32160 28284 32194 28318
rect 33178 28284 33212 28318
rect 17930 27130 17964 27164
rect 18948 27130 18982 27164
rect 19966 27130 20000 27164
rect 20984 27130 21018 27164
rect 22002 27130 22036 27164
rect 23020 27130 23054 27164
rect 24038 27130 24072 27164
rect 25056 27130 25090 27164
rect 26074 27130 26108 27164
rect 27092 27130 27126 27164
rect 28110 27130 28144 27164
rect 29128 27130 29162 27164
rect 30146 27130 30180 27164
rect 31164 27130 31198 27164
rect 32182 27130 32216 27164
rect 33200 27130 33234 27164
rect 17908 25998 17942 26032
rect 18926 25998 18960 26032
rect 19944 25998 19978 26032
rect 20962 25998 20996 26032
rect 21980 25998 22014 26032
rect 22998 25998 23032 26032
rect 24016 25998 24050 26032
rect 25034 25998 25068 26032
rect 26052 25998 26086 26032
rect 27070 25998 27104 26032
rect 28088 25998 28122 26032
rect 29106 25998 29140 26032
rect 30124 25998 30158 26032
rect 31142 25998 31176 26032
rect 32160 25998 32194 26032
rect 33178 25998 33212 26032
rect 17908 24616 17942 24650
rect 18926 24616 18960 24650
rect 19944 24616 19978 24650
rect 20962 24616 20996 24650
rect 21980 24616 22014 24650
rect 22998 24616 23032 24650
rect 24016 24616 24050 24650
rect 25034 24616 25068 24650
rect 26052 24616 26086 24650
rect 27070 24616 27104 24650
rect 28088 24616 28122 24650
rect 29106 24616 29140 24650
rect 30124 24616 30158 24650
rect 31142 24616 31176 24650
rect 32160 24616 32194 24650
rect 33178 24616 33212 24650
rect 18596 23268 18630 23302
rect 19614 23268 19648 23302
rect 20632 23268 20666 23302
rect 21650 23268 21684 23302
rect 22668 23268 22702 23302
rect 23686 23268 23720 23302
rect 24704 23268 24738 23302
rect 25722 23268 25756 23302
rect 26740 23268 26774 23302
rect 27758 23268 27792 23302
rect 28776 23268 28810 23302
rect 29794 23268 29828 23302
rect 30812 23268 30846 23302
rect 31830 23268 31864 23302
rect 32848 23268 32882 23302
rect 18202 21990 18236 22024
rect 19220 21990 19254 22024
rect 20238 21990 20272 22024
rect 21256 21990 21290 22024
rect 22274 21990 22308 22024
rect 23292 21990 23326 22024
rect 24310 21990 24344 22024
rect 25328 21990 25362 22024
rect 26346 21990 26380 22024
rect 27364 21990 27398 22024
rect 28382 21990 28416 22024
rect 29400 21990 29434 22024
rect 30418 21990 30452 22024
rect 31436 21990 31470 22024
rect 32454 21990 32488 22024
rect 33472 21990 33506 22024
rect 13604 21680 13638 21714
rect 14622 21680 14656 21714
rect 15640 21680 15674 21714
rect 16658 21680 16692 21714
rect 13080 20526 13114 20560
rect 14098 20526 14132 20560
rect 15116 20526 15150 20560
rect 16134 20526 16168 20560
rect 18292 20542 18326 20576
rect 19310 20542 19344 20576
rect 20328 20542 20362 20576
rect 21346 20542 21380 20576
rect 22364 20542 22398 20576
rect 23382 20542 23416 20576
rect 24400 20542 24434 20576
rect 25418 20542 25452 20576
rect 26436 20542 26470 20576
rect 27454 20542 27488 20576
rect 28472 20542 28506 20576
rect 29490 20542 29524 20576
rect 30508 20542 30542 20576
rect 31526 20542 31560 20576
rect 32544 20542 32578 20576
rect 33562 20542 33596 20576
rect 13090 19498 13124 19532
rect 14108 19498 14142 19532
rect 15126 19498 15160 19532
rect 16144 19498 16178 19532
rect 18316 19274 18350 19308
rect 19334 19274 19368 19308
rect 20352 19274 20386 19308
rect 21370 19274 21404 19308
rect 22388 19274 22422 19308
rect 23406 19274 23440 19308
rect 24424 19274 24458 19308
rect 25442 19274 25476 19308
rect 26460 19274 26494 19308
rect 27478 19274 27512 19308
rect 28496 19274 28530 19308
rect 29514 19274 29548 19308
rect 30532 19274 30566 19308
rect 31550 19274 31584 19308
rect 32568 19274 32602 19308
rect 33586 19274 33620 19308
rect 13080 18470 13114 18504
rect 14098 18470 14132 18504
rect 15116 18470 15150 18504
rect 16134 18470 16168 18504
rect 18180 18030 18214 18064
rect 19198 18030 19232 18064
rect 20216 18030 20250 18064
rect 21234 18030 21268 18064
rect 22252 18030 22286 18064
rect 23270 18030 23304 18064
rect 24288 18030 24322 18064
rect 25306 18030 25340 18064
rect 26324 18030 26358 18064
rect 27342 18030 27376 18064
rect 28360 18030 28394 18064
rect 29378 18030 29412 18064
rect 30396 18030 30430 18064
rect 31414 18030 31448 18064
rect 32432 18030 32466 18064
rect 33450 18030 33484 18064
rect 13604 17318 13638 17352
rect 14622 17318 14656 17352
rect 15640 17318 15674 17352
rect 16658 17318 16692 17352
rect -12184 16275 -10566 16309
rect -12280 15639 -12246 16213
rect -10504 15639 -10470 16213
rect -9584 16275 -7966 16309
rect -12184 15543 -10566 15577
rect -9680 15639 -9646 16213
rect -7904 15639 -7870 16213
rect 35634 16354 35734 30700
rect 11452 16192 35572 16292
rect -9584 15543 -7966 15577
<< poly >>
rect 17632 28095 18220 28111
rect 17632 28078 17648 28095
rect 17446 28061 17648 28078
rect 18204 28078 18220 28095
rect 18650 28095 19238 28111
rect 18650 28078 18666 28095
rect 18204 28061 18406 28078
rect 17446 28014 18406 28061
rect 18464 28061 18666 28078
rect 19222 28078 19238 28095
rect 19668 28095 20256 28111
rect 19668 28078 19684 28095
rect 19222 28061 19424 28078
rect 18464 28014 19424 28061
rect 19482 28061 19684 28078
rect 20240 28078 20256 28095
rect 20686 28095 21274 28111
rect 20686 28078 20702 28095
rect 20240 28061 20442 28078
rect 19482 28014 20442 28061
rect 20500 28061 20702 28078
rect 21258 28078 21274 28095
rect 21704 28095 22292 28111
rect 21704 28078 21720 28095
rect 21258 28061 21460 28078
rect 20500 28014 21460 28061
rect 21518 28061 21720 28078
rect 22276 28078 22292 28095
rect 22722 28095 23310 28111
rect 22722 28078 22738 28095
rect 22276 28061 22478 28078
rect 21518 28014 22478 28061
rect 22536 28061 22738 28078
rect 23294 28078 23310 28095
rect 23740 28095 24328 28111
rect 23740 28078 23756 28095
rect 23294 28061 23496 28078
rect 22536 28014 23496 28061
rect 23554 28061 23756 28078
rect 24312 28078 24328 28095
rect 24758 28095 25346 28111
rect 24758 28078 24774 28095
rect 24312 28061 24514 28078
rect 23554 28014 24514 28061
rect 24572 28061 24774 28078
rect 25330 28078 25346 28095
rect 25776 28095 26364 28111
rect 25776 28078 25792 28095
rect 25330 28061 25532 28078
rect 24572 28014 25532 28061
rect 25590 28061 25792 28078
rect 26348 28078 26364 28095
rect 26794 28095 27382 28111
rect 26794 28078 26810 28095
rect 26348 28061 26550 28078
rect 25590 28014 26550 28061
rect 26608 28061 26810 28078
rect 27366 28078 27382 28095
rect 27812 28095 28400 28111
rect 27812 28078 27828 28095
rect 27366 28061 27568 28078
rect 26608 28014 27568 28061
rect 27626 28061 27828 28078
rect 28384 28078 28400 28095
rect 28830 28095 29418 28111
rect 28830 28078 28846 28095
rect 28384 28061 28586 28078
rect 27626 28014 28586 28061
rect 28644 28061 28846 28078
rect 29402 28078 29418 28095
rect 29848 28095 30436 28111
rect 29848 28078 29864 28095
rect 29402 28061 29604 28078
rect 28644 28014 29604 28061
rect 29662 28061 29864 28078
rect 30420 28078 30436 28095
rect 30866 28095 31454 28111
rect 30866 28078 30882 28095
rect 30420 28061 30622 28078
rect 29662 28014 30622 28061
rect 30680 28061 30882 28078
rect 31438 28078 31454 28095
rect 31884 28095 32472 28111
rect 31884 28078 31900 28095
rect 31438 28061 31640 28078
rect 30680 28014 31640 28061
rect 31698 28061 31900 28078
rect 32456 28078 32472 28095
rect 32902 28095 33490 28111
rect 32902 28078 32918 28095
rect 32456 28061 32658 28078
rect 31698 28014 32658 28061
rect 32716 28061 32918 28078
rect 33474 28078 33490 28095
rect 33474 28061 33676 28078
rect 32716 28014 33676 28061
rect 17446 27367 18406 27414
rect 17446 27350 17648 27367
rect 17632 27333 17648 27350
rect 18204 27350 18406 27367
rect 18464 27367 19424 27414
rect 18464 27350 18666 27367
rect 18204 27333 18220 27350
rect 17632 27317 18220 27333
rect 18650 27333 18666 27350
rect 19222 27350 19424 27367
rect 19482 27367 20442 27414
rect 19482 27350 19684 27367
rect 19222 27333 19238 27350
rect 18650 27317 19238 27333
rect 19668 27333 19684 27350
rect 20240 27350 20442 27367
rect 20500 27367 21460 27414
rect 20500 27350 20702 27367
rect 20240 27333 20256 27350
rect 19668 27317 20256 27333
rect 20686 27333 20702 27350
rect 21258 27350 21460 27367
rect 21518 27367 22478 27414
rect 21518 27350 21720 27367
rect 21258 27333 21274 27350
rect 20686 27317 21274 27333
rect 21704 27333 21720 27350
rect 22276 27350 22478 27367
rect 22536 27367 23496 27414
rect 22536 27350 22738 27367
rect 22276 27333 22292 27350
rect 21704 27317 22292 27333
rect 22722 27333 22738 27350
rect 23294 27350 23496 27367
rect 23554 27367 24514 27414
rect 23554 27350 23756 27367
rect 23294 27333 23310 27350
rect 22722 27317 23310 27333
rect 23740 27333 23756 27350
rect 24312 27350 24514 27367
rect 24572 27367 25532 27414
rect 24572 27350 24774 27367
rect 24312 27333 24328 27350
rect 23740 27317 24328 27333
rect 24758 27333 24774 27350
rect 25330 27350 25532 27367
rect 25590 27367 26550 27414
rect 25590 27350 25792 27367
rect 25330 27333 25346 27350
rect 24758 27317 25346 27333
rect 25776 27333 25792 27350
rect 26348 27350 26550 27367
rect 26608 27367 27568 27414
rect 26608 27350 26810 27367
rect 26348 27333 26364 27350
rect 25776 27317 26364 27333
rect 26794 27333 26810 27350
rect 27366 27350 27568 27367
rect 27626 27367 28586 27414
rect 27626 27350 27828 27367
rect 27366 27333 27382 27350
rect 26794 27317 27382 27333
rect 27812 27333 27828 27350
rect 28384 27350 28586 27367
rect 28644 27367 29604 27414
rect 28644 27350 28846 27367
rect 28384 27333 28400 27350
rect 27812 27317 28400 27333
rect 28830 27333 28846 27350
rect 29402 27350 29604 27367
rect 29662 27367 30622 27414
rect 29662 27350 29864 27367
rect 29402 27333 29418 27350
rect 28830 27317 29418 27333
rect 29848 27333 29864 27350
rect 30420 27350 30622 27367
rect 30680 27367 31640 27414
rect 30680 27350 30882 27367
rect 30420 27333 30436 27350
rect 29848 27317 30436 27333
rect 30866 27333 30882 27350
rect 31438 27350 31640 27367
rect 31698 27367 32658 27414
rect 31698 27350 31900 27367
rect 31438 27333 31454 27350
rect 30866 27317 31454 27333
rect 31884 27333 31900 27350
rect 32456 27350 32658 27367
rect 32716 27367 33676 27414
rect 32716 27350 32918 27367
rect 32456 27333 32472 27350
rect 31884 27317 32472 27333
rect 32902 27333 32918 27350
rect 33474 27350 33676 27367
rect 33474 27333 33490 27350
rect 32902 27317 33490 27333
rect 17632 26959 18220 26975
rect 17632 26942 17648 26959
rect 17446 26925 17648 26942
rect 18204 26942 18220 26959
rect 18650 26959 19238 26975
rect 18650 26942 18666 26959
rect 18204 26925 18406 26942
rect 17446 26878 18406 26925
rect 18464 26925 18666 26942
rect 19222 26942 19238 26959
rect 19668 26959 20256 26975
rect 19668 26942 19684 26959
rect 19222 26925 19424 26942
rect 18464 26878 19424 26925
rect 19482 26925 19684 26942
rect 20240 26942 20256 26959
rect 20686 26959 21274 26975
rect 20686 26942 20702 26959
rect 20240 26925 20442 26942
rect 19482 26878 20442 26925
rect 20500 26925 20702 26942
rect 21258 26942 21274 26959
rect 21704 26959 22292 26975
rect 21704 26942 21720 26959
rect 21258 26925 21460 26942
rect 20500 26878 21460 26925
rect 21518 26925 21720 26942
rect 22276 26942 22292 26959
rect 22722 26959 23310 26975
rect 22722 26942 22738 26959
rect 22276 26925 22478 26942
rect 21518 26878 22478 26925
rect 22536 26925 22738 26942
rect 23294 26942 23310 26959
rect 23740 26959 24328 26975
rect 23740 26942 23756 26959
rect 23294 26925 23496 26942
rect 22536 26878 23496 26925
rect 23554 26925 23756 26942
rect 24312 26942 24328 26959
rect 24758 26959 25346 26975
rect 24758 26942 24774 26959
rect 24312 26925 24514 26942
rect 23554 26878 24514 26925
rect 24572 26925 24774 26942
rect 25330 26942 25346 26959
rect 25776 26959 26364 26975
rect 25776 26942 25792 26959
rect 25330 26925 25532 26942
rect 24572 26878 25532 26925
rect 25590 26925 25792 26942
rect 26348 26942 26364 26959
rect 26794 26959 27382 26975
rect 26794 26942 26810 26959
rect 26348 26925 26550 26942
rect 25590 26878 26550 26925
rect 26608 26925 26810 26942
rect 27366 26942 27382 26959
rect 27812 26959 28400 26975
rect 27812 26942 27828 26959
rect 27366 26925 27568 26942
rect 26608 26878 27568 26925
rect 27626 26925 27828 26942
rect 28384 26942 28400 26959
rect 28830 26959 29418 26975
rect 28830 26942 28846 26959
rect 28384 26925 28586 26942
rect 27626 26878 28586 26925
rect 28644 26925 28846 26942
rect 29402 26942 29418 26959
rect 29848 26959 30436 26975
rect 29848 26942 29864 26959
rect 29402 26925 29604 26942
rect 28644 26878 29604 26925
rect 29662 26925 29864 26942
rect 30420 26942 30436 26959
rect 30866 26959 31454 26975
rect 30866 26942 30882 26959
rect 30420 26925 30622 26942
rect 29662 26878 30622 26925
rect 30680 26925 30882 26942
rect 31438 26942 31454 26959
rect 31884 26959 32472 26975
rect 31884 26942 31900 26959
rect 31438 26925 31640 26942
rect 30680 26878 31640 26925
rect 31698 26925 31900 26942
rect 32456 26942 32472 26959
rect 32902 26959 33490 26975
rect 32902 26942 32918 26959
rect 32456 26925 32658 26942
rect 31698 26878 32658 26925
rect 32716 26925 32918 26942
rect 33474 26942 33490 26959
rect 33474 26925 33676 26942
rect 32716 26878 33676 26925
rect 17446 26231 18406 26278
rect 17446 26214 17648 26231
rect 17632 26197 17648 26214
rect 18204 26214 18406 26231
rect 18464 26231 19424 26278
rect 18464 26214 18666 26231
rect 18204 26197 18220 26214
rect 17632 26181 18220 26197
rect 18650 26197 18666 26214
rect 19222 26214 19424 26231
rect 19482 26231 20442 26278
rect 19482 26214 19684 26231
rect 19222 26197 19238 26214
rect 18650 26181 19238 26197
rect 19668 26197 19684 26214
rect 20240 26214 20442 26231
rect 20500 26231 21460 26278
rect 20500 26214 20702 26231
rect 20240 26197 20256 26214
rect 19668 26181 20256 26197
rect 20686 26197 20702 26214
rect 21258 26214 21460 26231
rect 21518 26231 22478 26278
rect 21518 26214 21720 26231
rect 21258 26197 21274 26214
rect 20686 26181 21274 26197
rect 21704 26197 21720 26214
rect 22276 26214 22478 26231
rect 22536 26231 23496 26278
rect 22536 26214 22738 26231
rect 22276 26197 22292 26214
rect 21704 26181 22292 26197
rect 22722 26197 22738 26214
rect 23294 26214 23496 26231
rect 23554 26231 24514 26278
rect 23554 26214 23756 26231
rect 23294 26197 23310 26214
rect 22722 26181 23310 26197
rect 23740 26197 23756 26214
rect 24312 26214 24514 26231
rect 24572 26231 25532 26278
rect 24572 26214 24774 26231
rect 24312 26197 24328 26214
rect 23740 26181 24328 26197
rect 24758 26197 24774 26214
rect 25330 26214 25532 26231
rect 25590 26231 26550 26278
rect 25590 26214 25792 26231
rect 25330 26197 25346 26214
rect 24758 26181 25346 26197
rect 25776 26197 25792 26214
rect 26348 26214 26550 26231
rect 26608 26231 27568 26278
rect 26608 26214 26810 26231
rect 26348 26197 26364 26214
rect 25776 26181 26364 26197
rect 26794 26197 26810 26214
rect 27366 26214 27568 26231
rect 27626 26231 28586 26278
rect 27626 26214 27828 26231
rect 27366 26197 27382 26214
rect 26794 26181 27382 26197
rect 27812 26197 27828 26214
rect 28384 26214 28586 26231
rect 28644 26231 29604 26278
rect 28644 26214 28846 26231
rect 28384 26197 28400 26214
rect 27812 26181 28400 26197
rect 28830 26197 28846 26214
rect 29402 26214 29604 26231
rect 29662 26231 30622 26278
rect 29662 26214 29864 26231
rect 29402 26197 29418 26214
rect 28830 26181 29418 26197
rect 29848 26197 29864 26214
rect 30420 26214 30622 26231
rect 30680 26231 31640 26278
rect 30680 26214 30882 26231
rect 30420 26197 30436 26214
rect 29848 26181 30436 26197
rect 30866 26197 30882 26214
rect 31438 26214 31640 26231
rect 31698 26231 32658 26278
rect 31698 26214 31900 26231
rect 31438 26197 31454 26214
rect 30866 26181 31454 26197
rect 31884 26197 31900 26214
rect 32456 26214 32658 26231
rect 32716 26231 33676 26278
rect 32716 26214 32918 26231
rect 32456 26197 32472 26214
rect 31884 26181 32472 26197
rect 32902 26197 32918 26214
rect 33474 26214 33676 26231
rect 33474 26197 33490 26214
rect 32902 26181 33490 26197
rect 17632 25823 18220 25839
rect 17632 25806 17648 25823
rect 17446 25789 17648 25806
rect 18204 25806 18220 25823
rect 18650 25823 19238 25839
rect 18650 25806 18666 25823
rect 18204 25789 18406 25806
rect 17446 25742 18406 25789
rect 18464 25789 18666 25806
rect 19222 25806 19238 25823
rect 19668 25823 20256 25839
rect 19668 25806 19684 25823
rect 19222 25789 19424 25806
rect 18464 25742 19424 25789
rect 19482 25789 19684 25806
rect 20240 25806 20256 25823
rect 20686 25823 21274 25839
rect 20686 25806 20702 25823
rect 20240 25789 20442 25806
rect 19482 25742 20442 25789
rect 20500 25789 20702 25806
rect 21258 25806 21274 25823
rect 21704 25823 22292 25839
rect 21704 25806 21720 25823
rect 21258 25789 21460 25806
rect 20500 25742 21460 25789
rect 21518 25789 21720 25806
rect 22276 25806 22292 25823
rect 22722 25823 23310 25839
rect 22722 25806 22738 25823
rect 22276 25789 22478 25806
rect 21518 25742 22478 25789
rect 22536 25789 22738 25806
rect 23294 25806 23310 25823
rect 23740 25823 24328 25839
rect 23740 25806 23756 25823
rect 23294 25789 23496 25806
rect 22536 25742 23496 25789
rect 23554 25789 23756 25806
rect 24312 25806 24328 25823
rect 24758 25823 25346 25839
rect 24758 25806 24774 25823
rect 24312 25789 24514 25806
rect 23554 25742 24514 25789
rect 24572 25789 24774 25806
rect 25330 25806 25346 25823
rect 25776 25823 26364 25839
rect 25776 25806 25792 25823
rect 25330 25789 25532 25806
rect 24572 25742 25532 25789
rect 25590 25789 25792 25806
rect 26348 25806 26364 25823
rect 26794 25823 27382 25839
rect 26794 25806 26810 25823
rect 26348 25789 26550 25806
rect 25590 25742 26550 25789
rect 26608 25789 26810 25806
rect 27366 25806 27382 25823
rect 27812 25823 28400 25839
rect 27812 25806 27828 25823
rect 27366 25789 27568 25806
rect 26608 25742 27568 25789
rect 27626 25789 27828 25806
rect 28384 25806 28400 25823
rect 28830 25823 29418 25839
rect 28830 25806 28846 25823
rect 28384 25789 28586 25806
rect 27626 25742 28586 25789
rect 28644 25789 28846 25806
rect 29402 25806 29418 25823
rect 29848 25823 30436 25839
rect 29848 25806 29864 25823
rect 29402 25789 29604 25806
rect 28644 25742 29604 25789
rect 29662 25789 29864 25806
rect 30420 25806 30436 25823
rect 30866 25823 31454 25839
rect 30866 25806 30882 25823
rect 30420 25789 30622 25806
rect 29662 25742 30622 25789
rect 30680 25789 30882 25806
rect 31438 25806 31454 25823
rect 31884 25823 32472 25839
rect 31884 25806 31900 25823
rect 31438 25789 31640 25806
rect 30680 25742 31640 25789
rect 31698 25789 31900 25806
rect 32456 25806 32472 25823
rect 32902 25823 33490 25839
rect 32902 25806 32918 25823
rect 32456 25789 32658 25806
rect 31698 25742 32658 25789
rect 32716 25789 32918 25806
rect 33474 25806 33490 25823
rect 33474 25789 33676 25806
rect 32716 25742 33676 25789
rect 17446 25095 18406 25142
rect 17446 25078 17648 25095
rect 17632 25061 17648 25078
rect 18204 25078 18406 25095
rect 18464 25095 19424 25142
rect 18464 25078 18666 25095
rect 18204 25061 18220 25078
rect 17632 25045 18220 25061
rect 18650 25061 18666 25078
rect 19222 25078 19424 25095
rect 19482 25095 20442 25142
rect 19482 25078 19684 25095
rect 19222 25061 19238 25078
rect 18650 25045 19238 25061
rect 19668 25061 19684 25078
rect 20240 25078 20442 25095
rect 20500 25095 21460 25142
rect 20500 25078 20702 25095
rect 20240 25061 20256 25078
rect 19668 25045 20256 25061
rect 20686 25061 20702 25078
rect 21258 25078 21460 25095
rect 21518 25095 22478 25142
rect 21518 25078 21720 25095
rect 21258 25061 21274 25078
rect 20686 25045 21274 25061
rect 21704 25061 21720 25078
rect 22276 25078 22478 25095
rect 22536 25095 23496 25142
rect 22536 25078 22738 25095
rect 22276 25061 22292 25078
rect 21704 25045 22292 25061
rect 22722 25061 22738 25078
rect 23294 25078 23496 25095
rect 23554 25095 24514 25142
rect 23554 25078 23756 25095
rect 23294 25061 23310 25078
rect 22722 25045 23310 25061
rect 23740 25061 23756 25078
rect 24312 25078 24514 25095
rect 24572 25095 25532 25142
rect 24572 25078 24774 25095
rect 24312 25061 24328 25078
rect 23740 25045 24328 25061
rect 24758 25061 24774 25078
rect 25330 25078 25532 25095
rect 25590 25095 26550 25142
rect 25590 25078 25792 25095
rect 25330 25061 25346 25078
rect 24758 25045 25346 25061
rect 25776 25061 25792 25078
rect 26348 25078 26550 25095
rect 26608 25095 27568 25142
rect 26608 25078 26810 25095
rect 26348 25061 26364 25078
rect 25776 25045 26364 25061
rect 26794 25061 26810 25078
rect 27366 25078 27568 25095
rect 27626 25095 28586 25142
rect 27626 25078 27828 25095
rect 27366 25061 27382 25078
rect 26794 25045 27382 25061
rect 27812 25061 27828 25078
rect 28384 25078 28586 25095
rect 28644 25095 29604 25142
rect 28644 25078 28846 25095
rect 28384 25061 28400 25078
rect 27812 25045 28400 25061
rect 28830 25061 28846 25078
rect 29402 25078 29604 25095
rect 29662 25095 30622 25142
rect 29662 25078 29864 25095
rect 29402 25061 29418 25078
rect 28830 25045 29418 25061
rect 29848 25061 29864 25078
rect 30420 25078 30622 25095
rect 30680 25095 31640 25142
rect 30680 25078 30882 25095
rect 30420 25061 30436 25078
rect 29848 25045 30436 25061
rect 30866 25061 30882 25078
rect 31438 25078 31640 25095
rect 31698 25095 32658 25142
rect 31698 25078 31900 25095
rect 31438 25061 31454 25078
rect 30866 25045 31454 25061
rect 31884 25061 31900 25078
rect 32456 25078 32658 25095
rect 32716 25095 33676 25142
rect 32716 25078 32918 25095
rect 32456 25061 32472 25078
rect 31884 25045 32472 25061
rect 32902 25061 32918 25078
rect 33474 25078 33676 25095
rect 33474 25061 33490 25078
rect 32902 25045 33490 25061
rect 18826 24185 19414 24201
rect 18826 24168 18842 24185
rect 18640 24151 18842 24168
rect 19398 24168 19414 24185
rect 19844 24185 20432 24201
rect 19844 24168 19860 24185
rect 19398 24151 19600 24168
rect 18640 24104 19600 24151
rect 19658 24151 19860 24168
rect 20416 24168 20432 24185
rect 20862 24185 21450 24201
rect 20862 24168 20878 24185
rect 20416 24151 20618 24168
rect 19658 24104 20618 24151
rect 20676 24151 20878 24168
rect 21434 24168 21450 24185
rect 21880 24185 22468 24201
rect 21880 24168 21896 24185
rect 21434 24151 21636 24168
rect 20676 24104 21636 24151
rect 21694 24151 21896 24168
rect 22452 24168 22468 24185
rect 22898 24185 23486 24201
rect 22898 24168 22914 24185
rect 22452 24151 22654 24168
rect 21694 24104 22654 24151
rect 22712 24151 22914 24168
rect 23470 24168 23486 24185
rect 23916 24185 24504 24201
rect 23916 24168 23932 24185
rect 23470 24151 23672 24168
rect 22712 24104 23672 24151
rect 23730 24151 23932 24168
rect 24488 24168 24504 24185
rect 24934 24185 25522 24201
rect 24934 24168 24950 24185
rect 24488 24151 24690 24168
rect 23730 24104 24690 24151
rect 24748 24151 24950 24168
rect 25506 24168 25522 24185
rect 25952 24185 26540 24201
rect 25952 24168 25968 24185
rect 25506 24151 25708 24168
rect 24748 24104 25708 24151
rect 25766 24151 25968 24168
rect 26524 24168 26540 24185
rect 26970 24185 27558 24201
rect 26970 24168 26986 24185
rect 26524 24151 26726 24168
rect 25766 24104 26726 24151
rect 26784 24151 26986 24168
rect 27542 24168 27558 24185
rect 27988 24185 28576 24201
rect 27988 24168 28004 24185
rect 27542 24151 27744 24168
rect 26784 24104 27744 24151
rect 27802 24151 28004 24168
rect 28560 24168 28576 24185
rect 29006 24185 29594 24201
rect 29006 24168 29022 24185
rect 28560 24151 28762 24168
rect 27802 24104 28762 24151
rect 28820 24151 29022 24168
rect 29578 24168 29594 24185
rect 30024 24185 30612 24201
rect 30024 24168 30040 24185
rect 29578 24151 29780 24168
rect 28820 24104 29780 24151
rect 29838 24151 30040 24168
rect 30596 24168 30612 24185
rect 31042 24185 31630 24201
rect 31042 24168 31058 24185
rect 30596 24151 30798 24168
rect 29838 24104 30798 24151
rect 30856 24151 31058 24168
rect 31614 24168 31630 24185
rect 32060 24185 32648 24201
rect 32060 24168 32076 24185
rect 31614 24151 31816 24168
rect 30856 24104 31816 24151
rect 31874 24151 32076 24168
rect 32632 24168 32648 24185
rect 32632 24151 32834 24168
rect 31874 24104 32834 24151
rect 18640 23457 19600 23504
rect 18640 23440 18842 23457
rect 18826 23423 18842 23440
rect 19398 23440 19600 23457
rect 19658 23457 20618 23504
rect 19658 23440 19860 23457
rect 19398 23423 19414 23440
rect 18826 23407 19414 23423
rect 19844 23423 19860 23440
rect 20416 23440 20618 23457
rect 20676 23457 21636 23504
rect 20676 23440 20878 23457
rect 20416 23423 20432 23440
rect 19844 23407 20432 23423
rect 20862 23423 20878 23440
rect 21434 23440 21636 23457
rect 21694 23457 22654 23504
rect 21694 23440 21896 23457
rect 21434 23423 21450 23440
rect 20862 23407 21450 23423
rect 21880 23423 21896 23440
rect 22452 23440 22654 23457
rect 22712 23457 23672 23504
rect 22712 23440 22914 23457
rect 22452 23423 22468 23440
rect 21880 23407 22468 23423
rect 22898 23423 22914 23440
rect 23470 23440 23672 23457
rect 23730 23457 24690 23504
rect 23730 23440 23932 23457
rect 23470 23423 23486 23440
rect 22898 23407 23486 23423
rect 23916 23423 23932 23440
rect 24488 23440 24690 23457
rect 24748 23457 25708 23504
rect 24748 23440 24950 23457
rect 24488 23423 24504 23440
rect 23916 23407 24504 23423
rect 24934 23423 24950 23440
rect 25506 23440 25708 23457
rect 25766 23457 26726 23504
rect 25766 23440 25968 23457
rect 25506 23423 25522 23440
rect 24934 23407 25522 23423
rect 25952 23423 25968 23440
rect 26524 23440 26726 23457
rect 26784 23457 27744 23504
rect 26784 23440 26986 23457
rect 26524 23423 26540 23440
rect 25952 23407 26540 23423
rect 26970 23423 26986 23440
rect 27542 23440 27744 23457
rect 27802 23457 28762 23504
rect 27802 23440 28004 23457
rect 27542 23423 27558 23440
rect 26970 23407 27558 23423
rect 27988 23423 28004 23440
rect 28560 23440 28762 23457
rect 28820 23457 29780 23504
rect 28820 23440 29022 23457
rect 28560 23423 28576 23440
rect 27988 23407 28576 23423
rect 29006 23423 29022 23440
rect 29578 23440 29780 23457
rect 29838 23457 30798 23504
rect 29838 23440 30040 23457
rect 29578 23423 29594 23440
rect 29006 23407 29594 23423
rect 30024 23423 30040 23440
rect 30596 23440 30798 23457
rect 30856 23457 31816 23504
rect 30856 23440 31058 23457
rect 30596 23423 30612 23440
rect 30024 23407 30612 23423
rect 31042 23423 31058 23440
rect 31614 23440 31816 23457
rect 31874 23457 32834 23504
rect 31874 23440 32076 23457
rect 31614 23423 31630 23440
rect 31042 23407 31630 23423
rect 32060 23423 32076 23440
rect 32632 23440 32834 23457
rect 32632 23423 32648 23440
rect 32060 23407 32648 23423
rect 18826 23153 19414 23169
rect 18826 23136 18842 23153
rect 18640 23119 18842 23136
rect 19398 23136 19414 23153
rect 19844 23153 20432 23169
rect 19844 23136 19860 23153
rect 19398 23119 19600 23136
rect 18640 23072 19600 23119
rect 19658 23119 19860 23136
rect 20416 23136 20432 23153
rect 20862 23153 21450 23169
rect 20862 23136 20878 23153
rect 20416 23119 20618 23136
rect 19658 23072 20618 23119
rect 20676 23119 20878 23136
rect 21434 23136 21450 23153
rect 21880 23153 22468 23169
rect 21880 23136 21896 23153
rect 21434 23119 21636 23136
rect 20676 23072 21636 23119
rect 21694 23119 21896 23136
rect 22452 23136 22468 23153
rect 22898 23153 23486 23169
rect 22898 23136 22914 23153
rect 22452 23119 22654 23136
rect 21694 23072 22654 23119
rect 22712 23119 22914 23136
rect 23470 23136 23486 23153
rect 23916 23153 24504 23169
rect 23916 23136 23932 23153
rect 23470 23119 23672 23136
rect 22712 23072 23672 23119
rect 23730 23119 23932 23136
rect 24488 23136 24504 23153
rect 24934 23153 25522 23169
rect 24934 23136 24950 23153
rect 24488 23119 24690 23136
rect 23730 23072 24690 23119
rect 24748 23119 24950 23136
rect 25506 23136 25522 23153
rect 25952 23153 26540 23169
rect 25952 23136 25968 23153
rect 25506 23119 25708 23136
rect 24748 23072 25708 23119
rect 25766 23119 25968 23136
rect 26524 23136 26540 23153
rect 26970 23153 27558 23169
rect 26970 23136 26986 23153
rect 26524 23119 26726 23136
rect 25766 23072 26726 23119
rect 26784 23119 26986 23136
rect 27542 23136 27558 23153
rect 27988 23153 28576 23169
rect 27988 23136 28004 23153
rect 27542 23119 27744 23136
rect 26784 23072 27744 23119
rect 27802 23119 28004 23136
rect 28560 23136 28576 23153
rect 29006 23153 29594 23169
rect 29006 23136 29022 23153
rect 28560 23119 28762 23136
rect 27802 23072 28762 23119
rect 28820 23119 29022 23136
rect 29578 23136 29594 23153
rect 30024 23153 30612 23169
rect 30024 23136 30040 23153
rect 29578 23119 29780 23136
rect 28820 23072 29780 23119
rect 29838 23119 30040 23136
rect 30596 23136 30612 23153
rect 31042 23153 31630 23169
rect 31042 23136 31058 23153
rect 30596 23119 30798 23136
rect 29838 23072 30798 23119
rect 30856 23119 31058 23136
rect 31614 23136 31630 23153
rect 32060 23153 32648 23169
rect 32060 23136 32076 23153
rect 31614 23119 31816 23136
rect 30856 23072 31816 23119
rect 31874 23119 32076 23136
rect 32632 23136 32648 23153
rect 32632 23119 32834 23136
rect 31874 23072 32834 23119
rect 18640 22425 19600 22472
rect 18640 22408 18842 22425
rect 18826 22391 18842 22408
rect 19398 22408 19600 22425
rect 19658 22425 20618 22472
rect 19658 22408 19860 22425
rect 19398 22391 19414 22408
rect 18826 22375 19414 22391
rect 19844 22391 19860 22408
rect 20416 22408 20618 22425
rect 20676 22425 21636 22472
rect 20676 22408 20878 22425
rect 20416 22391 20432 22408
rect 19844 22375 20432 22391
rect 20862 22391 20878 22408
rect 21434 22408 21636 22425
rect 21694 22425 22654 22472
rect 21694 22408 21896 22425
rect 21434 22391 21450 22408
rect 20862 22375 21450 22391
rect 21880 22391 21896 22408
rect 22452 22408 22654 22425
rect 22712 22425 23672 22472
rect 22712 22408 22914 22425
rect 22452 22391 22468 22408
rect 21880 22375 22468 22391
rect 22898 22391 22914 22408
rect 23470 22408 23672 22425
rect 23730 22425 24690 22472
rect 23730 22408 23932 22425
rect 23470 22391 23486 22408
rect 22898 22375 23486 22391
rect 23916 22391 23932 22408
rect 24488 22408 24690 22425
rect 24748 22425 25708 22472
rect 24748 22408 24950 22425
rect 24488 22391 24504 22408
rect 23916 22375 24504 22391
rect 24934 22391 24950 22408
rect 25506 22408 25708 22425
rect 25766 22425 26726 22472
rect 25766 22408 25968 22425
rect 25506 22391 25522 22408
rect 24934 22375 25522 22391
rect 25952 22391 25968 22408
rect 26524 22408 26726 22425
rect 26784 22425 27744 22472
rect 26784 22408 26986 22425
rect 26524 22391 26540 22408
rect 25952 22375 26540 22391
rect 26970 22391 26986 22408
rect 27542 22408 27744 22425
rect 27802 22425 28762 22472
rect 27802 22408 28004 22425
rect 27542 22391 27558 22408
rect 26970 22375 27558 22391
rect 27988 22391 28004 22408
rect 28560 22408 28762 22425
rect 28820 22425 29780 22472
rect 28820 22408 29022 22425
rect 28560 22391 28576 22408
rect 27988 22375 28576 22391
rect 29006 22391 29022 22408
rect 29578 22408 29780 22425
rect 29838 22425 30798 22472
rect 29838 22408 30040 22425
rect 29578 22391 29594 22408
rect 29006 22375 29594 22391
rect 30024 22391 30040 22408
rect 30596 22408 30798 22425
rect 30856 22425 31816 22472
rect 30856 22408 31058 22425
rect 30596 22391 30612 22408
rect 30024 22375 30612 22391
rect 31042 22391 31058 22408
rect 31614 22408 31816 22425
rect 31874 22425 32834 22472
rect 31874 22408 32076 22425
rect 31614 22391 31630 22408
rect 31042 22375 31630 22391
rect 32060 22391 32076 22408
rect 32632 22408 32834 22425
rect 32632 22391 32648 22408
rect 32060 22375 32648 22391
rect 18618 21549 19206 21565
rect 18618 21532 18634 21549
rect 18432 21515 18634 21532
rect 19190 21532 19206 21549
rect 19636 21549 20224 21565
rect 19636 21532 19652 21549
rect 19190 21515 19392 21532
rect 18432 21468 19392 21515
rect 19450 21515 19652 21532
rect 20208 21532 20224 21549
rect 20654 21549 21242 21565
rect 20654 21532 20670 21549
rect 20208 21515 20410 21532
rect 19450 21468 20410 21515
rect 20468 21515 20670 21532
rect 21226 21532 21242 21549
rect 21672 21549 22260 21565
rect 21672 21532 21688 21549
rect 21226 21515 21428 21532
rect 20468 21468 21428 21515
rect 21486 21515 21688 21532
rect 22244 21532 22260 21549
rect 22690 21549 23278 21565
rect 22690 21532 22706 21549
rect 22244 21515 22446 21532
rect 21486 21468 22446 21515
rect 22504 21515 22706 21532
rect 23262 21532 23278 21549
rect 23708 21549 24296 21565
rect 23708 21532 23724 21549
rect 23262 21515 23464 21532
rect 22504 21468 23464 21515
rect 23522 21515 23724 21532
rect 24280 21532 24296 21549
rect 24726 21549 25314 21565
rect 24726 21532 24742 21549
rect 24280 21515 24482 21532
rect 23522 21468 24482 21515
rect 24540 21515 24742 21532
rect 25298 21532 25314 21549
rect 25744 21549 26332 21565
rect 25744 21532 25760 21549
rect 25298 21515 25500 21532
rect 24540 21468 25500 21515
rect 25558 21515 25760 21532
rect 26316 21532 26332 21549
rect 26762 21549 27350 21565
rect 26762 21532 26778 21549
rect 26316 21515 26518 21532
rect 25558 21468 26518 21515
rect 26576 21515 26778 21532
rect 27334 21532 27350 21549
rect 27780 21549 28368 21565
rect 27780 21532 27796 21549
rect 27334 21515 27536 21532
rect 26576 21468 27536 21515
rect 27594 21515 27796 21532
rect 28352 21532 28368 21549
rect 28798 21549 29386 21565
rect 28798 21532 28814 21549
rect 28352 21515 28554 21532
rect 27594 21468 28554 21515
rect 28612 21515 28814 21532
rect 29370 21532 29386 21549
rect 29816 21549 30404 21565
rect 29816 21532 29832 21549
rect 29370 21515 29572 21532
rect 28612 21468 29572 21515
rect 29630 21515 29832 21532
rect 30388 21532 30404 21549
rect 30834 21549 31422 21565
rect 30834 21532 30850 21549
rect 30388 21515 30590 21532
rect 29630 21468 30590 21515
rect 30648 21515 30850 21532
rect 31406 21532 31422 21549
rect 31852 21549 32440 21565
rect 31852 21532 31868 21549
rect 31406 21515 31608 21532
rect 30648 21468 31608 21515
rect 31666 21515 31868 21532
rect 32424 21532 32440 21549
rect 32870 21549 33458 21565
rect 32870 21532 32886 21549
rect 32424 21515 32626 21532
rect 31666 21468 32626 21515
rect 32684 21515 32886 21532
rect 33442 21532 33458 21549
rect 33442 21515 33644 21532
rect 32684 21468 33644 21515
rect 13314 21445 13902 21461
rect 13314 21428 13330 21445
rect 13128 21411 13330 21428
rect 13886 21428 13902 21445
rect 14332 21445 14920 21461
rect 14332 21428 14348 21445
rect 13886 21411 14088 21428
rect 13128 21364 14088 21411
rect 14146 21411 14348 21428
rect 14904 21428 14920 21445
rect 15350 21445 15938 21461
rect 15350 21428 15366 21445
rect 14904 21411 15106 21428
rect 14146 21364 15106 21411
rect 15164 21411 15366 21428
rect 15922 21428 15938 21445
rect 16368 21445 16956 21461
rect 16368 21428 16384 21445
rect 15922 21411 16124 21428
rect 15164 21364 16124 21411
rect 16182 21411 16384 21428
rect 16940 21428 16956 21445
rect 16940 21411 17142 21428
rect 16182 21364 17142 21411
rect 18432 20821 19392 20868
rect 18432 20804 18634 20821
rect 18618 20787 18634 20804
rect 19190 20804 19392 20821
rect 19450 20821 20410 20868
rect 19450 20804 19652 20821
rect 19190 20787 19206 20804
rect 18618 20771 19206 20787
rect 19636 20787 19652 20804
rect 20208 20804 20410 20821
rect 20468 20821 21428 20868
rect 20468 20804 20670 20821
rect 20208 20787 20224 20804
rect 19636 20771 20224 20787
rect 20654 20787 20670 20804
rect 21226 20804 21428 20821
rect 21486 20821 22446 20868
rect 21486 20804 21688 20821
rect 21226 20787 21242 20804
rect 20654 20771 21242 20787
rect 21672 20787 21688 20804
rect 22244 20804 22446 20821
rect 22504 20821 23464 20868
rect 22504 20804 22706 20821
rect 22244 20787 22260 20804
rect 21672 20771 22260 20787
rect 22690 20787 22706 20804
rect 23262 20804 23464 20821
rect 23522 20821 24482 20868
rect 23522 20804 23724 20821
rect 23262 20787 23278 20804
rect 22690 20771 23278 20787
rect 23708 20787 23724 20804
rect 24280 20804 24482 20821
rect 24540 20821 25500 20868
rect 24540 20804 24742 20821
rect 24280 20787 24296 20804
rect 23708 20771 24296 20787
rect 24726 20787 24742 20804
rect 25298 20804 25500 20821
rect 25558 20821 26518 20868
rect 25558 20804 25760 20821
rect 25298 20787 25314 20804
rect 24726 20771 25314 20787
rect 25744 20787 25760 20804
rect 26316 20804 26518 20821
rect 26576 20821 27536 20868
rect 26576 20804 26778 20821
rect 26316 20787 26332 20804
rect 25744 20771 26332 20787
rect 26762 20787 26778 20804
rect 27334 20804 27536 20821
rect 27594 20821 28554 20868
rect 27594 20804 27796 20821
rect 27334 20787 27350 20804
rect 26762 20771 27350 20787
rect 27780 20787 27796 20804
rect 28352 20804 28554 20821
rect 28612 20821 29572 20868
rect 28612 20804 28814 20821
rect 28352 20787 28368 20804
rect 27780 20771 28368 20787
rect 28798 20787 28814 20804
rect 29370 20804 29572 20821
rect 29630 20821 30590 20868
rect 29630 20804 29832 20821
rect 29370 20787 29386 20804
rect 28798 20771 29386 20787
rect 29816 20787 29832 20804
rect 30388 20804 30590 20821
rect 30648 20821 31608 20868
rect 30648 20804 30850 20821
rect 30388 20787 30404 20804
rect 29816 20771 30404 20787
rect 30834 20787 30850 20804
rect 31406 20804 31608 20821
rect 31666 20821 32626 20868
rect 31666 20804 31868 20821
rect 31406 20787 31422 20804
rect 30834 20771 31422 20787
rect 31852 20787 31868 20804
rect 32424 20804 32626 20821
rect 32684 20821 33644 20868
rect 32684 20804 32886 20821
rect 32424 20787 32440 20804
rect 31852 20771 32440 20787
rect 32870 20787 32886 20804
rect 33442 20804 33644 20821
rect 33442 20787 33458 20804
rect 32870 20771 33458 20787
rect 13128 20717 14088 20764
rect 13128 20700 13330 20717
rect 13314 20683 13330 20700
rect 13886 20700 14088 20717
rect 14146 20717 15106 20764
rect 14146 20700 14348 20717
rect 13886 20683 13902 20700
rect 13314 20667 13902 20683
rect 14332 20683 14348 20700
rect 14904 20700 15106 20717
rect 15164 20717 16124 20764
rect 15164 20700 15366 20717
rect 14904 20683 14920 20700
rect 14332 20667 14920 20683
rect 15350 20683 15366 20700
rect 15922 20700 16124 20717
rect 16182 20717 17142 20764
rect 16182 20700 16384 20717
rect 15922 20683 15938 20700
rect 15350 20667 15938 20683
rect 16368 20683 16384 20700
rect 16940 20700 17142 20717
rect 16940 20683 16956 20700
rect 16368 20667 16956 20683
rect 13314 20413 13902 20429
rect 13314 20396 13330 20413
rect 13128 20379 13330 20396
rect 13886 20396 13902 20413
rect 14332 20413 14920 20429
rect 14332 20396 14348 20413
rect 13886 20379 14088 20396
rect 13128 20332 14088 20379
rect 14146 20379 14348 20396
rect 14904 20396 14920 20413
rect 15350 20413 15938 20429
rect 15350 20396 15366 20413
rect 14904 20379 15106 20396
rect 14146 20332 15106 20379
rect 15164 20379 15366 20396
rect 15922 20396 15938 20413
rect 16368 20413 16956 20429
rect 16368 20396 16384 20413
rect 15922 20379 16124 20396
rect 15164 20332 16124 20379
rect 16182 20379 16384 20396
rect 16940 20396 16956 20413
rect 16940 20379 17142 20396
rect 16182 20332 17142 20379
rect 18618 20293 19206 20309
rect 18618 20276 18634 20293
rect 18432 20259 18634 20276
rect 19190 20276 19206 20293
rect 19636 20293 20224 20309
rect 19636 20276 19652 20293
rect 19190 20259 19392 20276
rect 18432 20212 19392 20259
rect 19450 20259 19652 20276
rect 20208 20276 20224 20293
rect 20654 20293 21242 20309
rect 20654 20276 20670 20293
rect 20208 20259 20410 20276
rect 19450 20212 20410 20259
rect 20468 20259 20670 20276
rect 21226 20276 21242 20293
rect 21672 20293 22260 20309
rect 21672 20276 21688 20293
rect 21226 20259 21428 20276
rect 20468 20212 21428 20259
rect 21486 20259 21688 20276
rect 22244 20276 22260 20293
rect 22690 20293 23278 20309
rect 22690 20276 22706 20293
rect 22244 20259 22446 20276
rect 21486 20212 22446 20259
rect 22504 20259 22706 20276
rect 23262 20276 23278 20293
rect 23708 20293 24296 20309
rect 23708 20276 23724 20293
rect 23262 20259 23464 20276
rect 22504 20212 23464 20259
rect 23522 20259 23724 20276
rect 24280 20276 24296 20293
rect 24726 20293 25314 20309
rect 24726 20276 24742 20293
rect 24280 20259 24482 20276
rect 23522 20212 24482 20259
rect 24540 20259 24742 20276
rect 25298 20276 25314 20293
rect 25744 20293 26332 20309
rect 25744 20276 25760 20293
rect 25298 20259 25500 20276
rect 24540 20212 25500 20259
rect 25558 20259 25760 20276
rect 26316 20276 26332 20293
rect 26762 20293 27350 20309
rect 26762 20276 26778 20293
rect 26316 20259 26518 20276
rect 25558 20212 26518 20259
rect 26576 20259 26778 20276
rect 27334 20276 27350 20293
rect 27780 20293 28368 20309
rect 27780 20276 27796 20293
rect 27334 20259 27536 20276
rect 26576 20212 27536 20259
rect 27594 20259 27796 20276
rect 28352 20276 28368 20293
rect 28798 20293 29386 20309
rect 28798 20276 28814 20293
rect 28352 20259 28554 20276
rect 27594 20212 28554 20259
rect 28612 20259 28814 20276
rect 29370 20276 29386 20293
rect 29816 20293 30404 20309
rect 29816 20276 29832 20293
rect 29370 20259 29572 20276
rect 28612 20212 29572 20259
rect 29630 20259 29832 20276
rect 30388 20276 30404 20293
rect 30834 20293 31422 20309
rect 30834 20276 30850 20293
rect 30388 20259 30590 20276
rect 29630 20212 30590 20259
rect 30648 20259 30850 20276
rect 31406 20276 31422 20293
rect 31852 20293 32440 20309
rect 31852 20276 31868 20293
rect 31406 20259 31608 20276
rect 30648 20212 31608 20259
rect 31666 20259 31868 20276
rect 32424 20276 32440 20293
rect 32870 20293 33458 20309
rect 32870 20276 32886 20293
rect 32424 20259 32626 20276
rect 31666 20212 32626 20259
rect 32684 20259 32886 20276
rect 33442 20276 33458 20293
rect 33442 20259 33644 20276
rect 32684 20212 33644 20259
rect 13128 19685 14088 19732
rect 13128 19668 13330 19685
rect 13314 19651 13330 19668
rect 13886 19668 14088 19685
rect 14146 19685 15106 19732
rect 14146 19668 14348 19685
rect 13886 19651 13902 19668
rect 13314 19635 13902 19651
rect 14332 19651 14348 19668
rect 14904 19668 15106 19685
rect 15164 19685 16124 19732
rect 15164 19668 15366 19685
rect 14904 19651 14920 19668
rect 14332 19635 14920 19651
rect 15350 19651 15366 19668
rect 15922 19668 16124 19685
rect 16182 19685 17142 19732
rect 16182 19668 16384 19685
rect 15922 19651 15938 19668
rect 15350 19635 15938 19651
rect 16368 19651 16384 19668
rect 16940 19668 17142 19685
rect 16940 19651 16956 19668
rect 16368 19635 16956 19651
rect 18432 19565 19392 19612
rect 18432 19548 18634 19565
rect 18618 19531 18634 19548
rect 19190 19548 19392 19565
rect 19450 19565 20410 19612
rect 19450 19548 19652 19565
rect 19190 19531 19206 19548
rect 18618 19515 19206 19531
rect 19636 19531 19652 19548
rect 20208 19548 20410 19565
rect 20468 19565 21428 19612
rect 20468 19548 20670 19565
rect 20208 19531 20224 19548
rect 19636 19515 20224 19531
rect 20654 19531 20670 19548
rect 21226 19548 21428 19565
rect 21486 19565 22446 19612
rect 21486 19548 21688 19565
rect 21226 19531 21242 19548
rect 20654 19515 21242 19531
rect 21672 19531 21688 19548
rect 22244 19548 22446 19565
rect 22504 19565 23464 19612
rect 22504 19548 22706 19565
rect 22244 19531 22260 19548
rect 21672 19515 22260 19531
rect 22690 19531 22706 19548
rect 23262 19548 23464 19565
rect 23522 19565 24482 19612
rect 23522 19548 23724 19565
rect 23262 19531 23278 19548
rect 22690 19515 23278 19531
rect 23708 19531 23724 19548
rect 24280 19548 24482 19565
rect 24540 19565 25500 19612
rect 24540 19548 24742 19565
rect 24280 19531 24296 19548
rect 23708 19515 24296 19531
rect 24726 19531 24742 19548
rect 25298 19548 25500 19565
rect 25558 19565 26518 19612
rect 25558 19548 25760 19565
rect 25298 19531 25314 19548
rect 24726 19515 25314 19531
rect 25744 19531 25760 19548
rect 26316 19548 26518 19565
rect 26576 19565 27536 19612
rect 26576 19548 26778 19565
rect 26316 19531 26332 19548
rect 25744 19515 26332 19531
rect 26762 19531 26778 19548
rect 27334 19548 27536 19565
rect 27594 19565 28554 19612
rect 27594 19548 27796 19565
rect 27334 19531 27350 19548
rect 26762 19515 27350 19531
rect 27780 19531 27796 19548
rect 28352 19548 28554 19565
rect 28612 19565 29572 19612
rect 28612 19548 28814 19565
rect 28352 19531 28368 19548
rect 27780 19515 28368 19531
rect 28798 19531 28814 19548
rect 29370 19548 29572 19565
rect 29630 19565 30590 19612
rect 29630 19548 29832 19565
rect 29370 19531 29386 19548
rect 28798 19515 29386 19531
rect 29816 19531 29832 19548
rect 30388 19548 30590 19565
rect 30648 19565 31608 19612
rect 30648 19548 30850 19565
rect 30388 19531 30404 19548
rect 29816 19515 30404 19531
rect 30834 19531 30850 19548
rect 31406 19548 31608 19565
rect 31666 19565 32626 19612
rect 31666 19548 31868 19565
rect 31406 19531 31422 19548
rect 30834 19515 31422 19531
rect 31852 19531 31868 19548
rect 32424 19548 32626 19565
rect 32684 19565 33644 19612
rect 32684 19548 32886 19565
rect 32424 19531 32440 19548
rect 31852 19515 32440 19531
rect 32870 19531 32886 19548
rect 33442 19548 33644 19565
rect 33442 19531 33458 19548
rect 32870 19515 33458 19531
rect 13314 19381 13902 19397
rect 13314 19364 13330 19381
rect 13128 19347 13330 19364
rect 13886 19364 13902 19381
rect 14332 19381 14920 19397
rect 14332 19364 14348 19381
rect 13886 19347 14088 19364
rect 13128 19300 14088 19347
rect 14146 19347 14348 19364
rect 14904 19364 14920 19381
rect 15350 19381 15938 19397
rect 15350 19364 15366 19381
rect 14904 19347 15106 19364
rect 14146 19300 15106 19347
rect 15164 19347 15366 19364
rect 15922 19364 15938 19381
rect 16368 19381 16956 19397
rect 16368 19364 16384 19381
rect 15922 19347 16124 19364
rect 15164 19300 16124 19347
rect 16182 19347 16384 19364
rect 16940 19364 16956 19381
rect 16940 19347 17142 19364
rect 16182 19300 17142 19347
rect 18618 19037 19206 19053
rect 18618 19020 18634 19037
rect 18432 19003 18634 19020
rect 19190 19020 19206 19037
rect 19636 19037 20224 19053
rect 19636 19020 19652 19037
rect 19190 19003 19392 19020
rect 18432 18956 19392 19003
rect 19450 19003 19652 19020
rect 20208 19020 20224 19037
rect 20654 19037 21242 19053
rect 20654 19020 20670 19037
rect 20208 19003 20410 19020
rect 19450 18956 20410 19003
rect 20468 19003 20670 19020
rect 21226 19020 21242 19037
rect 21672 19037 22260 19053
rect 21672 19020 21688 19037
rect 21226 19003 21428 19020
rect 20468 18956 21428 19003
rect 21486 19003 21688 19020
rect 22244 19020 22260 19037
rect 22690 19037 23278 19053
rect 22690 19020 22706 19037
rect 22244 19003 22446 19020
rect 21486 18956 22446 19003
rect 22504 19003 22706 19020
rect 23262 19020 23278 19037
rect 23708 19037 24296 19053
rect 23708 19020 23724 19037
rect 23262 19003 23464 19020
rect 22504 18956 23464 19003
rect 23522 19003 23724 19020
rect 24280 19020 24296 19037
rect 24726 19037 25314 19053
rect 24726 19020 24742 19037
rect 24280 19003 24482 19020
rect 23522 18956 24482 19003
rect 24540 19003 24742 19020
rect 25298 19020 25314 19037
rect 25744 19037 26332 19053
rect 25744 19020 25760 19037
rect 25298 19003 25500 19020
rect 24540 18956 25500 19003
rect 25558 19003 25760 19020
rect 26316 19020 26332 19037
rect 26762 19037 27350 19053
rect 26762 19020 26778 19037
rect 26316 19003 26518 19020
rect 25558 18956 26518 19003
rect 26576 19003 26778 19020
rect 27334 19020 27350 19037
rect 27780 19037 28368 19053
rect 27780 19020 27796 19037
rect 27334 19003 27536 19020
rect 26576 18956 27536 19003
rect 27594 19003 27796 19020
rect 28352 19020 28368 19037
rect 28798 19037 29386 19053
rect 28798 19020 28814 19037
rect 28352 19003 28554 19020
rect 27594 18956 28554 19003
rect 28612 19003 28814 19020
rect 29370 19020 29386 19037
rect 29816 19037 30404 19053
rect 29816 19020 29832 19037
rect 29370 19003 29572 19020
rect 28612 18956 29572 19003
rect 29630 19003 29832 19020
rect 30388 19020 30404 19037
rect 30834 19037 31422 19053
rect 30834 19020 30850 19037
rect 30388 19003 30590 19020
rect 29630 18956 30590 19003
rect 30648 19003 30850 19020
rect 31406 19020 31422 19037
rect 31852 19037 32440 19053
rect 31852 19020 31868 19037
rect 31406 19003 31608 19020
rect 30648 18956 31608 19003
rect 31666 19003 31868 19020
rect 32424 19020 32440 19037
rect 32870 19037 33458 19053
rect 32870 19020 32886 19037
rect 32424 19003 32626 19020
rect 31666 18956 32626 19003
rect 32684 19003 32886 19020
rect 33442 19020 33458 19037
rect 33442 19003 33644 19020
rect 32684 18956 33644 19003
rect 13128 18653 14088 18700
rect 13128 18636 13330 18653
rect 13314 18619 13330 18636
rect 13886 18636 14088 18653
rect 14146 18653 15106 18700
rect 14146 18636 14348 18653
rect 13886 18619 13902 18636
rect 13314 18603 13902 18619
rect 14332 18619 14348 18636
rect 14904 18636 15106 18653
rect 15164 18653 16124 18700
rect 15164 18636 15366 18653
rect 14904 18619 14920 18636
rect 14332 18603 14920 18619
rect 15350 18619 15366 18636
rect 15922 18636 16124 18653
rect 16182 18653 17142 18700
rect 16182 18636 16384 18653
rect 15922 18619 15938 18636
rect 15350 18603 15938 18619
rect 16368 18619 16384 18636
rect 16940 18636 17142 18653
rect 16940 18619 16956 18636
rect 16368 18603 16956 18619
rect 13314 18349 13902 18365
rect 13314 18332 13330 18349
rect 13128 18315 13330 18332
rect 13886 18332 13902 18349
rect 14332 18349 14920 18365
rect 14332 18332 14348 18349
rect 13886 18315 14088 18332
rect 13128 18268 14088 18315
rect 14146 18315 14348 18332
rect 14904 18332 14920 18349
rect 15350 18349 15938 18365
rect 15350 18332 15366 18349
rect 14904 18315 15106 18332
rect 14146 18268 15106 18315
rect 15164 18315 15366 18332
rect 15922 18332 15938 18349
rect 16368 18349 16956 18365
rect 16368 18332 16384 18349
rect 15922 18315 16124 18332
rect 15164 18268 16124 18315
rect 16182 18315 16384 18332
rect 16940 18332 16956 18349
rect 16940 18315 17142 18332
rect 16182 18268 17142 18315
rect 18432 18309 19392 18356
rect 18432 18292 18634 18309
rect 18618 18275 18634 18292
rect 19190 18292 19392 18309
rect 19450 18309 20410 18356
rect 19450 18292 19652 18309
rect 19190 18275 19206 18292
rect 18618 18259 19206 18275
rect 19636 18275 19652 18292
rect 20208 18292 20410 18309
rect 20468 18309 21428 18356
rect 20468 18292 20670 18309
rect 20208 18275 20224 18292
rect 19636 18259 20224 18275
rect 20654 18275 20670 18292
rect 21226 18292 21428 18309
rect 21486 18309 22446 18356
rect 21486 18292 21688 18309
rect 21226 18275 21242 18292
rect 20654 18259 21242 18275
rect 21672 18275 21688 18292
rect 22244 18292 22446 18309
rect 22504 18309 23464 18356
rect 22504 18292 22706 18309
rect 22244 18275 22260 18292
rect 21672 18259 22260 18275
rect 22690 18275 22706 18292
rect 23262 18292 23464 18309
rect 23522 18309 24482 18356
rect 23522 18292 23724 18309
rect 23262 18275 23278 18292
rect 22690 18259 23278 18275
rect 23708 18275 23724 18292
rect 24280 18292 24482 18309
rect 24540 18309 25500 18356
rect 24540 18292 24742 18309
rect 24280 18275 24296 18292
rect 23708 18259 24296 18275
rect 24726 18275 24742 18292
rect 25298 18292 25500 18309
rect 25558 18309 26518 18356
rect 25558 18292 25760 18309
rect 25298 18275 25314 18292
rect 24726 18259 25314 18275
rect 25744 18275 25760 18292
rect 26316 18292 26518 18309
rect 26576 18309 27536 18356
rect 26576 18292 26778 18309
rect 26316 18275 26332 18292
rect 25744 18259 26332 18275
rect 26762 18275 26778 18292
rect 27334 18292 27536 18309
rect 27594 18309 28554 18356
rect 27594 18292 27796 18309
rect 27334 18275 27350 18292
rect 26762 18259 27350 18275
rect 27780 18275 27796 18292
rect 28352 18292 28554 18309
rect 28612 18309 29572 18356
rect 28612 18292 28814 18309
rect 28352 18275 28368 18292
rect 27780 18259 28368 18275
rect 28798 18275 28814 18292
rect 29370 18292 29572 18309
rect 29630 18309 30590 18356
rect 29630 18292 29832 18309
rect 29370 18275 29386 18292
rect 28798 18259 29386 18275
rect 29816 18275 29832 18292
rect 30388 18292 30590 18309
rect 30648 18309 31608 18356
rect 30648 18292 30850 18309
rect 30388 18275 30404 18292
rect 29816 18259 30404 18275
rect 30834 18275 30850 18292
rect 31406 18292 31608 18309
rect 31666 18309 32626 18356
rect 31666 18292 31868 18309
rect 31406 18275 31422 18292
rect 30834 18259 31422 18275
rect 31852 18275 31868 18292
rect 32424 18292 32626 18309
rect 32684 18309 33644 18356
rect 32684 18292 32886 18309
rect 32424 18275 32440 18292
rect 31852 18259 32440 18275
rect 32870 18275 32886 18292
rect 33442 18292 33644 18309
rect 33442 18275 33458 18292
rect 32870 18259 33458 18275
rect 18618 17781 19206 17797
rect 18618 17764 18634 17781
rect 18432 17747 18634 17764
rect 19190 17764 19206 17781
rect 19636 17781 20224 17797
rect 19636 17764 19652 17781
rect 19190 17747 19392 17764
rect 18432 17700 19392 17747
rect 19450 17747 19652 17764
rect 20208 17764 20224 17781
rect 20654 17781 21242 17797
rect 20654 17764 20670 17781
rect 20208 17747 20410 17764
rect 19450 17700 20410 17747
rect 20468 17747 20670 17764
rect 21226 17764 21242 17781
rect 21672 17781 22260 17797
rect 21672 17764 21688 17781
rect 21226 17747 21428 17764
rect 20468 17700 21428 17747
rect 21486 17747 21688 17764
rect 22244 17764 22260 17781
rect 22690 17781 23278 17797
rect 22690 17764 22706 17781
rect 22244 17747 22446 17764
rect 21486 17700 22446 17747
rect 22504 17747 22706 17764
rect 23262 17764 23278 17781
rect 23708 17781 24296 17797
rect 23708 17764 23724 17781
rect 23262 17747 23464 17764
rect 22504 17700 23464 17747
rect 23522 17747 23724 17764
rect 24280 17764 24296 17781
rect 24726 17781 25314 17797
rect 24726 17764 24742 17781
rect 24280 17747 24482 17764
rect 23522 17700 24482 17747
rect 24540 17747 24742 17764
rect 25298 17764 25314 17781
rect 25744 17781 26332 17797
rect 25744 17764 25760 17781
rect 25298 17747 25500 17764
rect 24540 17700 25500 17747
rect 25558 17747 25760 17764
rect 26316 17764 26332 17781
rect 26762 17781 27350 17797
rect 26762 17764 26778 17781
rect 26316 17747 26518 17764
rect 25558 17700 26518 17747
rect 26576 17747 26778 17764
rect 27334 17764 27350 17781
rect 27780 17781 28368 17797
rect 27780 17764 27796 17781
rect 27334 17747 27536 17764
rect 26576 17700 27536 17747
rect 27594 17747 27796 17764
rect 28352 17764 28368 17781
rect 28798 17781 29386 17797
rect 28798 17764 28814 17781
rect 28352 17747 28554 17764
rect 27594 17700 28554 17747
rect 28612 17747 28814 17764
rect 29370 17764 29386 17781
rect 29816 17781 30404 17797
rect 29816 17764 29832 17781
rect 29370 17747 29572 17764
rect 28612 17700 29572 17747
rect 29630 17747 29832 17764
rect 30388 17764 30404 17781
rect 30834 17781 31422 17797
rect 30834 17764 30850 17781
rect 30388 17747 30590 17764
rect 29630 17700 30590 17747
rect 30648 17747 30850 17764
rect 31406 17764 31422 17781
rect 31852 17781 32440 17797
rect 31852 17764 31868 17781
rect 31406 17747 31608 17764
rect 30648 17700 31608 17747
rect 31666 17747 31868 17764
rect 32424 17764 32440 17781
rect 32870 17781 33458 17797
rect 32870 17764 32886 17781
rect 32424 17747 32626 17764
rect 31666 17700 32626 17747
rect 32684 17747 32886 17764
rect 33442 17764 33458 17781
rect 33442 17747 33644 17764
rect 32684 17700 33644 17747
rect 13128 17621 14088 17668
rect 13128 17604 13330 17621
rect 13314 17587 13330 17604
rect 13886 17604 14088 17621
rect 14146 17621 15106 17668
rect 14146 17604 14348 17621
rect 13886 17587 13902 17604
rect 13314 17571 13902 17587
rect 14332 17587 14348 17604
rect 14904 17604 15106 17621
rect 15164 17621 16124 17668
rect 15164 17604 15366 17621
rect 14904 17587 14920 17604
rect 14332 17571 14920 17587
rect 15350 17587 15366 17604
rect 15922 17604 16124 17621
rect 16182 17621 17142 17668
rect 16182 17604 16384 17621
rect 15922 17587 15938 17604
rect 15350 17571 15938 17587
rect 16368 17587 16384 17604
rect 16940 17604 17142 17621
rect 16940 17587 16956 17604
rect 16368 17571 16956 17587
rect 18432 17053 19392 17100
rect 18432 17036 18634 17053
rect 18618 17019 18634 17036
rect 19190 17036 19392 17053
rect 19450 17053 20410 17100
rect 19450 17036 19652 17053
rect 19190 17019 19206 17036
rect 18618 17003 19206 17019
rect 19636 17019 19652 17036
rect 20208 17036 20410 17053
rect 20468 17053 21428 17100
rect 20468 17036 20670 17053
rect 20208 17019 20224 17036
rect 19636 17003 20224 17019
rect 20654 17019 20670 17036
rect 21226 17036 21428 17053
rect 21486 17053 22446 17100
rect 21486 17036 21688 17053
rect 21226 17019 21242 17036
rect 20654 17003 21242 17019
rect 21672 17019 21688 17036
rect 22244 17036 22446 17053
rect 22504 17053 23464 17100
rect 22504 17036 22706 17053
rect 22244 17019 22260 17036
rect 21672 17003 22260 17019
rect 22690 17019 22706 17036
rect 23262 17036 23464 17053
rect 23522 17053 24482 17100
rect 23522 17036 23724 17053
rect 23262 17019 23278 17036
rect 22690 17003 23278 17019
rect 23708 17019 23724 17036
rect 24280 17036 24482 17053
rect 24540 17053 25500 17100
rect 24540 17036 24742 17053
rect 24280 17019 24296 17036
rect 23708 17003 24296 17019
rect 24726 17019 24742 17036
rect 25298 17036 25500 17053
rect 25558 17053 26518 17100
rect 25558 17036 25760 17053
rect 25298 17019 25314 17036
rect 24726 17003 25314 17019
rect 25744 17019 25760 17036
rect 26316 17036 26518 17053
rect 26576 17053 27536 17100
rect 26576 17036 26778 17053
rect 26316 17019 26332 17036
rect 25744 17003 26332 17019
rect 26762 17019 26778 17036
rect 27334 17036 27536 17053
rect 27594 17053 28554 17100
rect 27594 17036 27796 17053
rect 27334 17019 27350 17036
rect 26762 17003 27350 17019
rect 27780 17019 27796 17036
rect 28352 17036 28554 17053
rect 28612 17053 29572 17100
rect 28612 17036 28814 17053
rect 28352 17019 28368 17036
rect 27780 17003 28368 17019
rect 28798 17019 28814 17036
rect 29370 17036 29572 17053
rect 29630 17053 30590 17100
rect 29630 17036 29832 17053
rect 29370 17019 29386 17036
rect 28798 17003 29386 17019
rect 29816 17019 29832 17036
rect 30388 17036 30590 17053
rect 30648 17053 31608 17100
rect 30648 17036 30850 17053
rect 30388 17019 30404 17036
rect 29816 17003 30404 17019
rect 30834 17019 30850 17036
rect 31406 17036 31608 17053
rect 31666 17053 32626 17100
rect 31666 17036 31868 17053
rect 31406 17019 31422 17036
rect 30834 17003 31422 17019
rect 31852 17019 31868 17036
rect 32424 17036 32626 17053
rect 32684 17053 33644 17100
rect 32684 17036 32886 17053
rect 32424 17019 32440 17036
rect 31852 17003 32440 17019
rect 32870 17019 32886 17036
rect 33442 17036 33644 17053
rect 33442 17019 33458 17036
rect 32870 17003 33458 17019
rect -12086 16207 -11954 16223
rect -12086 16190 -12070 16207
rect -12120 16173 -12070 16190
rect -11970 16190 -11954 16207
rect -11828 16207 -11696 16223
rect -11828 16190 -11812 16207
rect -11970 16173 -11920 16190
rect -12120 16126 -11920 16173
rect -11862 16173 -11812 16190
rect -11712 16190 -11696 16207
rect -11570 16207 -11438 16223
rect -11570 16190 -11554 16207
rect -11712 16173 -11662 16190
rect -11862 16126 -11662 16173
rect -11604 16173 -11554 16190
rect -11454 16190 -11438 16207
rect -11312 16207 -11180 16223
rect -11312 16190 -11296 16207
rect -11454 16173 -11404 16190
rect -11604 16126 -11404 16173
rect -11346 16173 -11296 16190
rect -11196 16190 -11180 16207
rect -11054 16207 -10922 16223
rect -11054 16190 -11038 16207
rect -11196 16173 -11146 16190
rect -11346 16126 -11146 16173
rect -11088 16173 -11038 16190
rect -10938 16190 -10922 16207
rect -10796 16207 -10664 16223
rect -10796 16190 -10780 16207
rect -10938 16173 -10888 16190
rect -11088 16126 -10888 16173
rect -10830 16173 -10780 16190
rect -10680 16190 -10664 16207
rect -10680 16173 -10630 16190
rect -10830 16126 -10630 16173
rect -12120 15679 -11920 15726
rect -12120 15662 -12070 15679
rect -12086 15645 -12070 15662
rect -11970 15662 -11920 15679
rect -11862 15679 -11662 15726
rect -11862 15662 -11812 15679
rect -11970 15645 -11954 15662
rect -12086 15629 -11954 15645
rect -11828 15645 -11812 15662
rect -11712 15662 -11662 15679
rect -11604 15679 -11404 15726
rect -11604 15662 -11554 15679
rect -11712 15645 -11696 15662
rect -11828 15629 -11696 15645
rect -11570 15645 -11554 15662
rect -11454 15662 -11404 15679
rect -11346 15679 -11146 15726
rect -11346 15662 -11296 15679
rect -11454 15645 -11438 15662
rect -11570 15629 -11438 15645
rect -11312 15645 -11296 15662
rect -11196 15662 -11146 15679
rect -11088 15679 -10888 15726
rect -11088 15662 -11038 15679
rect -11196 15645 -11180 15662
rect -11312 15629 -11180 15645
rect -11054 15645 -11038 15662
rect -10938 15662 -10888 15679
rect -10830 15679 -10630 15726
rect -10830 15662 -10780 15679
rect -10938 15645 -10922 15662
rect -11054 15629 -10922 15645
rect -10796 15645 -10780 15662
rect -10680 15662 -10630 15679
rect -10680 15645 -10664 15662
rect -10796 15629 -10664 15645
rect -10270 15743 -10240 15769
rect -9486 16207 -9354 16223
rect -9486 16190 -9470 16207
rect -9520 16173 -9470 16190
rect -9370 16190 -9354 16207
rect -9228 16207 -9096 16223
rect -9228 16190 -9212 16207
rect -9370 16173 -9320 16190
rect -9520 16126 -9320 16173
rect -9262 16173 -9212 16190
rect -9112 16190 -9096 16207
rect -8970 16207 -8838 16223
rect -8970 16190 -8954 16207
rect -9112 16173 -9062 16190
rect -9262 16126 -9062 16173
rect -9004 16173 -8954 16190
rect -8854 16190 -8838 16207
rect -8712 16207 -8580 16223
rect -8712 16190 -8696 16207
rect -8854 16173 -8804 16190
rect -9004 16126 -8804 16173
rect -8746 16173 -8696 16190
rect -8596 16190 -8580 16207
rect -8454 16207 -8322 16223
rect -8454 16190 -8438 16207
rect -8596 16173 -8546 16190
rect -8746 16126 -8546 16173
rect -8488 16173 -8438 16190
rect -8338 16190 -8322 16207
rect -8196 16207 -8064 16223
rect -8196 16190 -8180 16207
rect -8338 16173 -8288 16190
rect -8488 16126 -8288 16173
rect -8230 16173 -8180 16190
rect -8080 16190 -8064 16207
rect -8080 16173 -8030 16190
rect -8230 16126 -8030 16173
rect -9520 15679 -9320 15726
rect -9520 15662 -9470 15679
rect -9486 15645 -9470 15662
rect -9370 15662 -9320 15679
rect -9262 15679 -9062 15726
rect -9262 15662 -9212 15679
rect -9370 15645 -9354 15662
rect -9486 15629 -9354 15645
rect -9228 15645 -9212 15662
rect -9112 15662 -9062 15679
rect -9004 15679 -8804 15726
rect -9004 15662 -8954 15679
rect -9112 15645 -9096 15662
rect -9228 15629 -9096 15645
rect -8970 15645 -8954 15662
rect -8854 15662 -8804 15679
rect -8746 15679 -8546 15726
rect -8746 15662 -8696 15679
rect -8854 15645 -8838 15662
rect -8970 15629 -8838 15645
rect -8712 15645 -8696 15662
rect -8596 15662 -8546 15679
rect -8488 15679 -8288 15726
rect -8488 15662 -8438 15679
rect -8596 15645 -8580 15662
rect -8712 15629 -8580 15645
rect -8454 15645 -8438 15662
rect -8338 15662 -8288 15679
rect -8230 15679 -8030 15726
rect -8230 15662 -8180 15679
rect -8338 15645 -8322 15662
rect -8454 15629 -8322 15645
rect -8196 15645 -8180 15662
rect -8080 15662 -8030 15679
rect -8080 15645 -8064 15662
rect -8196 15629 -8064 15645
rect -7670 15743 -7640 15769
rect -7220 15743 -7190 15769
rect -10270 15511 -10240 15543
rect -7670 15511 -7640 15543
rect -7220 15511 -7190 15543
rect -10270 15495 -10184 15511
rect -10270 15461 -10234 15495
rect -10200 15461 -10184 15495
rect -10270 15445 -10184 15461
rect -7670 15495 -7584 15511
rect -7670 15461 -7634 15495
rect -7600 15461 -7584 15495
rect -7670 15445 -7584 15461
rect -7220 15495 -7134 15511
rect -7220 15461 -7184 15495
rect -7150 15461 -7134 15495
rect -7220 15445 -7134 15461
rect -10270 15423 -10240 15445
rect -7670 15423 -7640 15445
rect -7220 15423 -7190 15445
rect -12086 15274 -11954 15290
rect -12086 15257 -12070 15274
rect -12120 15240 -12070 15257
rect -11970 15257 -11954 15274
rect -11828 15274 -11696 15290
rect -11828 15257 -11812 15274
rect -11970 15240 -11920 15257
rect -12120 15202 -11920 15240
rect -11862 15240 -11812 15257
rect -11712 15257 -11696 15274
rect -11570 15274 -11438 15290
rect -11570 15257 -11554 15274
rect -11712 15240 -11662 15257
rect -11862 15202 -11662 15240
rect -11604 15240 -11554 15257
rect -11454 15257 -11438 15274
rect -11312 15274 -11180 15290
rect -11312 15257 -11296 15274
rect -11454 15240 -11404 15257
rect -11604 15202 -11404 15240
rect -11346 15240 -11296 15257
rect -11196 15257 -11180 15274
rect -11054 15274 -10922 15290
rect -11054 15257 -11038 15274
rect -11196 15240 -11146 15257
rect -11346 15202 -11146 15240
rect -11088 15240 -11038 15257
rect -10938 15257 -10922 15274
rect -10796 15274 -10664 15290
rect -10796 15257 -10780 15274
rect -10938 15240 -10888 15257
rect -11088 15202 -10888 15240
rect -10830 15240 -10780 15257
rect -10680 15257 -10664 15274
rect -10680 15240 -10630 15257
rect -10830 15202 -10630 15240
rect -12120 14964 -11920 15002
rect -12120 14947 -12070 14964
rect -12086 14930 -12070 14947
rect -11970 14947 -11920 14964
rect -11862 14964 -11662 15002
rect -11862 14947 -11812 14964
rect -11970 14930 -11954 14947
rect -12086 14914 -11954 14930
rect -11828 14930 -11812 14947
rect -11712 14947 -11662 14964
rect -11604 14964 -11404 15002
rect -11604 14947 -11554 14964
rect -11712 14930 -11696 14947
rect -11828 14914 -11696 14930
rect -11570 14930 -11554 14947
rect -11454 14947 -11404 14964
rect -11346 14964 -11146 15002
rect -11346 14947 -11296 14964
rect -11454 14930 -11438 14947
rect -11570 14914 -11438 14930
rect -11312 14930 -11296 14947
rect -11196 14947 -11146 14964
rect -11088 14964 -10888 15002
rect -11088 14947 -11038 14964
rect -11196 14930 -11180 14947
rect -11312 14914 -11180 14930
rect -11054 14930 -11038 14947
rect -10938 14947 -10888 14964
rect -10830 14964 -10630 15002
rect -10830 14947 -10780 14964
rect -10938 14930 -10922 14947
rect -11054 14914 -10922 14930
rect -10796 14930 -10780 14947
rect -10680 14947 -10630 14964
rect -10680 14930 -10664 14947
rect -10796 14914 -10664 14930
rect -10270 15267 -10240 15293
rect -9486 15274 -9354 15290
rect -9486 15257 -9470 15274
rect -9520 15240 -9470 15257
rect -9370 15257 -9354 15274
rect -9228 15274 -9096 15290
rect -9228 15257 -9212 15274
rect -9370 15240 -9320 15257
rect -9520 15202 -9320 15240
rect -9262 15240 -9212 15257
rect -9112 15257 -9096 15274
rect -8970 15274 -8838 15290
rect -8970 15257 -8954 15274
rect -9112 15240 -9062 15257
rect -9262 15202 -9062 15240
rect -9004 15240 -8954 15257
rect -8854 15257 -8838 15274
rect -8712 15274 -8580 15290
rect -8712 15257 -8696 15274
rect -8854 15240 -8804 15257
rect -9004 15202 -8804 15240
rect -8746 15240 -8696 15257
rect -8596 15257 -8580 15274
rect -8454 15274 -8322 15290
rect -8454 15257 -8438 15274
rect -8596 15240 -8546 15257
rect -8746 15202 -8546 15240
rect -8488 15240 -8438 15257
rect -8338 15257 -8322 15274
rect -8196 15274 -8064 15290
rect -8196 15257 -8180 15274
rect -8338 15240 -8288 15257
rect -8488 15202 -8288 15240
rect -8230 15240 -8180 15257
rect -8080 15257 -8064 15274
rect -8080 15240 -8030 15257
rect -8230 15202 -8030 15240
rect -9520 14964 -9320 15002
rect -9520 14947 -9470 14964
rect -9486 14930 -9470 14947
rect -9370 14947 -9320 14964
rect -9262 14964 -9062 15002
rect -9262 14947 -9212 14964
rect -9370 14930 -9354 14947
rect -9486 14914 -9354 14930
rect -9228 14930 -9212 14947
rect -9112 14947 -9062 14964
rect -9004 14964 -8804 15002
rect -9004 14947 -8954 14964
rect -9112 14930 -9096 14947
rect -9228 14914 -9096 14930
rect -8970 14930 -8954 14947
rect -8854 14947 -8804 14964
rect -8746 14964 -8546 15002
rect -8746 14947 -8696 14964
rect -8854 14930 -8838 14947
rect -8970 14914 -8838 14930
rect -8712 14930 -8696 14947
rect -8596 14947 -8546 14964
rect -8488 14964 -8288 15002
rect -8488 14947 -8438 14964
rect -8596 14930 -8580 14947
rect -8712 14914 -8580 14930
rect -8454 14930 -8438 14947
rect -8338 14947 -8288 14964
rect -8230 14964 -8030 15002
rect -8230 14947 -8180 14964
rect -8338 14930 -8322 14947
rect -8454 14914 -8322 14930
rect -8196 14930 -8180 14947
rect -8080 14947 -8030 14964
rect -8080 14930 -8064 14947
rect -8196 14914 -8064 14930
rect -7670 15267 -7640 15293
rect -7220 15267 -7190 15293
rect 13726 14576 14314 14592
rect 13726 14559 13742 14576
rect 13540 14542 13742 14559
rect 14298 14559 14314 14576
rect 14744 14576 15332 14592
rect 14744 14559 14760 14576
rect 14298 14542 14500 14559
rect 13540 14504 14500 14542
rect 14558 14542 14760 14559
rect 15316 14559 15332 14576
rect 15762 14576 16350 14592
rect 15762 14559 15778 14576
rect 15316 14542 15518 14559
rect 14558 14504 15518 14542
rect 15576 14542 15778 14559
rect 16334 14559 16350 14576
rect 16780 14576 17368 14592
rect 16780 14559 16796 14576
rect 16334 14542 16536 14559
rect 15576 14504 16536 14542
rect 16594 14542 16796 14559
rect 17352 14559 17368 14576
rect 17798 14576 18386 14592
rect 17798 14559 17814 14576
rect 17352 14542 17554 14559
rect 16594 14504 17554 14542
rect 17612 14542 17814 14559
rect 18370 14559 18386 14576
rect 18816 14576 19404 14592
rect 18816 14559 18832 14576
rect 18370 14542 18572 14559
rect 17612 14504 18572 14542
rect 18630 14542 18832 14559
rect 19388 14559 19404 14576
rect 19834 14576 20422 14592
rect 19834 14559 19850 14576
rect 19388 14542 19590 14559
rect 18630 14504 19590 14542
rect 19648 14542 19850 14559
rect 20406 14559 20422 14576
rect 20852 14576 21440 14592
rect 20852 14559 20868 14576
rect 20406 14542 20608 14559
rect 19648 14504 20608 14542
rect 20666 14542 20868 14559
rect 21424 14559 21440 14576
rect 21870 14576 22458 14592
rect 21870 14559 21886 14576
rect 21424 14542 21626 14559
rect 20666 14504 21626 14542
rect 21684 14542 21886 14559
rect 22442 14559 22458 14576
rect 22888 14576 23476 14592
rect 22888 14559 22904 14576
rect 22442 14542 22644 14559
rect 21684 14504 22644 14542
rect 22702 14542 22904 14559
rect 23460 14559 23476 14576
rect 23906 14576 24494 14592
rect 23906 14559 23922 14576
rect 23460 14542 23662 14559
rect 22702 14504 23662 14542
rect 23720 14542 23922 14559
rect 24478 14559 24494 14576
rect 24924 14576 25512 14592
rect 24924 14559 24940 14576
rect 24478 14542 24680 14559
rect 23720 14504 24680 14542
rect 24738 14542 24940 14559
rect 25496 14559 25512 14576
rect 25942 14576 26530 14592
rect 25942 14559 25958 14576
rect 25496 14542 25698 14559
rect 24738 14504 25698 14542
rect 25756 14542 25958 14559
rect 26514 14559 26530 14576
rect 26960 14576 27548 14592
rect 26960 14559 26976 14576
rect 26514 14542 26716 14559
rect 25756 14504 26716 14542
rect 26774 14542 26976 14559
rect 27532 14559 27548 14576
rect 27978 14576 28566 14592
rect 27978 14559 27994 14576
rect 27532 14542 27734 14559
rect 26774 14504 27734 14542
rect 27792 14542 27994 14559
rect 28550 14559 28566 14576
rect 28996 14576 29584 14592
rect 28996 14559 29012 14576
rect 28550 14542 28752 14559
rect 27792 14504 28752 14542
rect 28810 14542 29012 14559
rect 29568 14559 29584 14576
rect 30014 14576 30602 14592
rect 30014 14559 30030 14576
rect 29568 14542 29770 14559
rect 28810 14504 29770 14542
rect 29828 14542 30030 14559
rect 30586 14559 30602 14576
rect 31032 14576 31620 14592
rect 31032 14559 31048 14576
rect 30586 14542 30788 14559
rect 29828 14504 30788 14542
rect 30846 14542 31048 14559
rect 31604 14559 31620 14576
rect 32050 14576 32638 14592
rect 32050 14559 32066 14576
rect 31604 14542 31806 14559
rect 30846 14504 31806 14542
rect 31864 14542 32066 14559
rect 32622 14559 32638 14576
rect 33068 14576 33656 14592
rect 33068 14559 33084 14576
rect 32622 14542 32824 14559
rect 31864 14504 32824 14542
rect 32882 14542 33084 14559
rect 33640 14559 33656 14576
rect 33640 14542 33842 14559
rect 32882 14504 33842 14542
rect 1960 14100 2548 14116
rect 1960 14083 1976 14100
rect 1774 14066 1976 14083
rect 2532 14083 2548 14100
rect 2978 14100 3566 14116
rect 2978 14083 2994 14100
rect 2532 14066 2734 14083
rect 1774 14028 2734 14066
rect 2792 14066 2994 14083
rect 3550 14083 3566 14100
rect 3996 14100 4584 14116
rect 3996 14083 4012 14100
rect 3550 14066 3752 14083
rect 2792 14028 3752 14066
rect 3810 14066 4012 14083
rect 4568 14083 4584 14100
rect 5014 14100 5602 14116
rect 5014 14083 5030 14100
rect 4568 14066 4770 14083
rect 3810 14028 4770 14066
rect 4828 14066 5030 14083
rect 5586 14083 5602 14100
rect 6032 14100 6620 14116
rect 6032 14083 6048 14100
rect 5586 14066 5788 14083
rect 4828 14028 5788 14066
rect 5846 14066 6048 14083
rect 6604 14083 6620 14100
rect 7050 14100 7638 14116
rect 7050 14083 7066 14100
rect 6604 14066 6806 14083
rect 5846 14028 6806 14066
rect 6864 14066 7066 14083
rect 7622 14083 7638 14100
rect 8068 14100 8656 14116
rect 8068 14083 8084 14100
rect 7622 14066 7824 14083
rect 6864 14028 7824 14066
rect 7882 14066 8084 14083
rect 8640 14083 8656 14100
rect 9086 14100 9674 14116
rect 9086 14083 9102 14100
rect 8640 14066 8842 14083
rect 7882 14028 8842 14066
rect 8900 14066 9102 14083
rect 9658 14083 9674 14100
rect 10104 14100 10692 14116
rect 10104 14083 10120 14100
rect 9658 14066 9860 14083
rect 8900 14028 9860 14066
rect 9918 14066 10120 14083
rect 10676 14083 10692 14100
rect 10676 14066 10878 14083
rect 9918 14028 10878 14066
rect 13540 13866 14500 13904
rect 13540 13849 13742 13866
rect 13726 13832 13742 13849
rect 14298 13849 14500 13866
rect 14558 13866 15518 13904
rect 14558 13849 14760 13866
rect 14298 13832 14314 13849
rect 13726 13816 14314 13832
rect 14744 13832 14760 13849
rect 15316 13849 15518 13866
rect 15576 13866 16536 13904
rect 15576 13849 15778 13866
rect 15316 13832 15332 13849
rect 14744 13816 15332 13832
rect 15762 13832 15778 13849
rect 16334 13849 16536 13866
rect 16594 13866 17554 13904
rect 16594 13849 16796 13866
rect 16334 13832 16350 13849
rect 15762 13816 16350 13832
rect 16780 13832 16796 13849
rect 17352 13849 17554 13866
rect 17612 13866 18572 13904
rect 17612 13849 17814 13866
rect 17352 13832 17368 13849
rect 16780 13816 17368 13832
rect 17798 13832 17814 13849
rect 18370 13849 18572 13866
rect 18630 13866 19590 13904
rect 18630 13849 18832 13866
rect 18370 13832 18386 13849
rect 17798 13816 18386 13832
rect 18816 13832 18832 13849
rect 19388 13849 19590 13866
rect 19648 13866 20608 13904
rect 19648 13849 19850 13866
rect 19388 13832 19404 13849
rect 18816 13816 19404 13832
rect 19834 13832 19850 13849
rect 20406 13849 20608 13866
rect 20666 13866 21626 13904
rect 20666 13849 20868 13866
rect 20406 13832 20422 13849
rect 19834 13816 20422 13832
rect 20852 13832 20868 13849
rect 21424 13849 21626 13866
rect 21684 13866 22644 13904
rect 21684 13849 21886 13866
rect 21424 13832 21440 13849
rect 20852 13816 21440 13832
rect 21870 13832 21886 13849
rect 22442 13849 22644 13866
rect 22702 13866 23662 13904
rect 22702 13849 22904 13866
rect 22442 13832 22458 13849
rect 21870 13816 22458 13832
rect 22888 13832 22904 13849
rect 23460 13849 23662 13866
rect 23720 13866 24680 13904
rect 23720 13849 23922 13866
rect 23460 13832 23476 13849
rect 22888 13816 23476 13832
rect 23906 13832 23922 13849
rect 24478 13849 24680 13866
rect 24738 13866 25698 13904
rect 24738 13849 24940 13866
rect 24478 13832 24494 13849
rect 23906 13816 24494 13832
rect 24924 13832 24940 13849
rect 25496 13849 25698 13866
rect 25756 13866 26716 13904
rect 25756 13849 25958 13866
rect 25496 13832 25512 13849
rect 24924 13816 25512 13832
rect 25942 13832 25958 13849
rect 26514 13849 26716 13866
rect 26774 13866 27734 13904
rect 26774 13849 26976 13866
rect 26514 13832 26530 13849
rect 25942 13816 26530 13832
rect 26960 13832 26976 13849
rect 27532 13849 27734 13866
rect 27792 13866 28752 13904
rect 27792 13849 27994 13866
rect 27532 13832 27548 13849
rect 26960 13816 27548 13832
rect 27978 13832 27994 13849
rect 28550 13849 28752 13866
rect 28810 13866 29770 13904
rect 28810 13849 29012 13866
rect 28550 13832 28566 13849
rect 27978 13816 28566 13832
rect 28996 13832 29012 13849
rect 29568 13849 29770 13866
rect 29828 13866 30788 13904
rect 29828 13849 30030 13866
rect 29568 13832 29584 13849
rect 28996 13816 29584 13832
rect 30014 13832 30030 13849
rect 30586 13849 30788 13866
rect 30846 13866 31806 13904
rect 30846 13849 31048 13866
rect 30586 13832 30602 13849
rect 30014 13816 30602 13832
rect 31032 13832 31048 13849
rect 31604 13849 31806 13866
rect 31864 13866 32824 13904
rect 31864 13849 32066 13866
rect 31604 13832 31620 13849
rect 31032 13816 31620 13832
rect 32050 13832 32066 13849
rect 32622 13849 32824 13866
rect 32882 13866 33842 13904
rect 32882 13849 33084 13866
rect 32622 13832 32638 13849
rect 32050 13816 32638 13832
rect 33068 13832 33084 13849
rect 33640 13849 33842 13866
rect 33640 13832 33656 13849
rect 33068 13816 33656 13832
rect 13726 13758 14314 13774
rect 13726 13741 13742 13758
rect 13540 13724 13742 13741
rect 14298 13741 14314 13758
rect 14744 13758 15332 13774
rect 14744 13741 14760 13758
rect 14298 13724 14500 13741
rect 13540 13686 14500 13724
rect 14558 13724 14760 13741
rect 15316 13741 15332 13758
rect 15762 13758 16350 13774
rect 15762 13741 15778 13758
rect 15316 13724 15518 13741
rect 14558 13686 15518 13724
rect 15576 13724 15778 13741
rect 16334 13741 16350 13758
rect 16780 13758 17368 13774
rect 16780 13741 16796 13758
rect 16334 13724 16536 13741
rect 15576 13686 16536 13724
rect 16594 13724 16796 13741
rect 17352 13741 17368 13758
rect 17798 13758 18386 13774
rect 17798 13741 17814 13758
rect 17352 13724 17554 13741
rect 16594 13686 17554 13724
rect 17612 13724 17814 13741
rect 18370 13741 18386 13758
rect 18816 13758 19404 13774
rect 18816 13741 18832 13758
rect 18370 13724 18572 13741
rect 17612 13686 18572 13724
rect 18630 13724 18832 13741
rect 19388 13741 19404 13758
rect 19834 13758 20422 13774
rect 19834 13741 19850 13758
rect 19388 13724 19590 13741
rect 18630 13686 19590 13724
rect 19648 13724 19850 13741
rect 20406 13741 20422 13758
rect 20852 13758 21440 13774
rect 20852 13741 20868 13758
rect 20406 13724 20608 13741
rect 19648 13686 20608 13724
rect 20666 13724 20868 13741
rect 21424 13741 21440 13758
rect 21870 13758 22458 13774
rect 21870 13741 21886 13758
rect 21424 13724 21626 13741
rect 20666 13686 21626 13724
rect 21684 13724 21886 13741
rect 22442 13741 22458 13758
rect 22888 13758 23476 13774
rect 22888 13741 22904 13758
rect 22442 13724 22644 13741
rect 21684 13686 22644 13724
rect 22702 13724 22904 13741
rect 23460 13741 23476 13758
rect 23906 13758 24494 13774
rect 23906 13741 23922 13758
rect 23460 13724 23662 13741
rect 22702 13686 23662 13724
rect 23720 13724 23922 13741
rect 24478 13741 24494 13758
rect 24924 13758 25512 13774
rect 24924 13741 24940 13758
rect 24478 13724 24680 13741
rect 23720 13686 24680 13724
rect 24738 13724 24940 13741
rect 25496 13741 25512 13758
rect 25942 13758 26530 13774
rect 25942 13741 25958 13758
rect 25496 13724 25698 13741
rect 24738 13686 25698 13724
rect 25756 13724 25958 13741
rect 26514 13741 26530 13758
rect 26960 13758 27548 13774
rect 26960 13741 26976 13758
rect 26514 13724 26716 13741
rect 25756 13686 26716 13724
rect 26774 13724 26976 13741
rect 27532 13741 27548 13758
rect 27978 13758 28566 13774
rect 27978 13741 27994 13758
rect 27532 13724 27734 13741
rect 26774 13686 27734 13724
rect 27792 13724 27994 13741
rect 28550 13741 28566 13758
rect 28996 13758 29584 13774
rect 28996 13741 29012 13758
rect 28550 13724 28752 13741
rect 27792 13686 28752 13724
rect 28810 13724 29012 13741
rect 29568 13741 29584 13758
rect 30014 13758 30602 13774
rect 30014 13741 30030 13758
rect 29568 13724 29770 13741
rect 28810 13686 29770 13724
rect 29828 13724 30030 13741
rect 30586 13741 30602 13758
rect 31032 13758 31620 13774
rect 31032 13741 31048 13758
rect 30586 13724 30788 13741
rect 29828 13686 30788 13724
rect 30846 13724 31048 13741
rect 31604 13741 31620 13758
rect 32050 13758 32638 13774
rect 32050 13741 32066 13758
rect 31604 13724 31806 13741
rect 30846 13686 31806 13724
rect 31864 13724 32066 13741
rect 32622 13741 32638 13758
rect 33068 13758 33656 13774
rect 33068 13741 33084 13758
rect 32622 13724 32824 13741
rect 31864 13686 32824 13724
rect 32882 13724 33084 13741
rect 33640 13741 33656 13758
rect 33640 13724 33842 13741
rect 32882 13686 33842 13724
rect 1774 13390 2734 13428
rect 1774 13373 1976 13390
rect 1960 13356 1976 13373
rect 2532 13373 2734 13390
rect 2792 13390 3752 13428
rect 2792 13373 2994 13390
rect 2532 13356 2548 13373
rect 1960 13340 2548 13356
rect 2978 13356 2994 13373
rect 3550 13373 3752 13390
rect 3810 13390 4770 13428
rect 3810 13373 4012 13390
rect 3550 13356 3566 13373
rect 2978 13340 3566 13356
rect 1960 13282 2548 13298
rect 1960 13265 1976 13282
rect 1774 13248 1976 13265
rect 2532 13265 2548 13282
rect 3996 13356 4012 13373
rect 4568 13373 4770 13390
rect 4828 13390 5788 13428
rect 4828 13373 5030 13390
rect 4568 13356 4584 13373
rect 3996 13340 4584 13356
rect 2978 13282 3566 13298
rect 2978 13265 2994 13282
rect 2532 13248 2734 13265
rect 1774 13210 2734 13248
rect 2792 13248 2994 13265
rect 3550 13265 3566 13282
rect 5014 13356 5030 13373
rect 5586 13373 5788 13390
rect 5846 13390 6806 13428
rect 5846 13373 6048 13390
rect 5586 13356 5602 13373
rect 5014 13340 5602 13356
rect 3996 13282 4584 13298
rect 3996 13265 4012 13282
rect 3550 13248 3752 13265
rect 2792 13210 3752 13248
rect 3810 13248 4012 13265
rect 4568 13265 4584 13282
rect 6032 13356 6048 13373
rect 6604 13373 6806 13390
rect 6864 13390 7824 13428
rect 6864 13373 7066 13390
rect 6604 13356 6620 13373
rect 6032 13340 6620 13356
rect 5014 13282 5602 13298
rect 5014 13265 5030 13282
rect 4568 13248 4770 13265
rect 3810 13210 4770 13248
rect 4828 13248 5030 13265
rect 5586 13265 5602 13282
rect 7050 13356 7066 13373
rect 7622 13373 7824 13390
rect 7882 13390 8842 13428
rect 7882 13373 8084 13390
rect 7622 13356 7638 13373
rect 7050 13340 7638 13356
rect 6032 13282 6620 13298
rect 6032 13265 6048 13282
rect 5586 13248 5788 13265
rect 4828 13210 5788 13248
rect 5846 13248 6048 13265
rect 6604 13265 6620 13282
rect 8068 13356 8084 13373
rect 8640 13373 8842 13390
rect 8900 13390 9860 13428
rect 8900 13373 9102 13390
rect 8640 13356 8656 13373
rect 8068 13340 8656 13356
rect 7050 13282 7638 13298
rect 7050 13265 7066 13282
rect 6604 13248 6806 13265
rect 5846 13210 6806 13248
rect 6864 13248 7066 13265
rect 7622 13265 7638 13282
rect 9086 13356 9102 13373
rect 9658 13373 9860 13390
rect 9918 13390 10878 13428
rect 9918 13373 10120 13390
rect 9658 13356 9674 13373
rect 9086 13340 9674 13356
rect 8068 13282 8656 13298
rect 8068 13265 8084 13282
rect 7622 13248 7824 13265
rect 6864 13210 7824 13248
rect 7882 13248 8084 13265
rect 8640 13265 8656 13282
rect 10104 13356 10120 13373
rect 10676 13373 10878 13390
rect 10676 13356 10692 13373
rect 10104 13340 10692 13356
rect 9086 13282 9674 13298
rect 9086 13265 9102 13282
rect 8640 13248 8842 13265
rect 7882 13210 8842 13248
rect 8900 13248 9102 13265
rect 9658 13265 9674 13282
rect 10104 13282 10692 13298
rect 10104 13265 10120 13282
rect 9658 13248 9860 13265
rect 8900 13210 9860 13248
rect 9918 13248 10120 13265
rect 10676 13265 10692 13282
rect 10676 13248 10878 13265
rect 9918 13210 10878 13248
rect 13540 13048 14500 13086
rect 13540 13031 13742 13048
rect 13726 13014 13742 13031
rect 14298 13031 14500 13048
rect 14558 13048 15518 13086
rect 14558 13031 14760 13048
rect 14298 13014 14314 13031
rect 13726 12998 14314 13014
rect 14744 13014 14760 13031
rect 15316 13031 15518 13048
rect 15576 13048 16536 13086
rect 15576 13031 15778 13048
rect 15316 13014 15332 13031
rect 14744 12998 15332 13014
rect 15762 13014 15778 13031
rect 16334 13031 16536 13048
rect 16594 13048 17554 13086
rect 16594 13031 16796 13048
rect 16334 13014 16350 13031
rect 15762 12998 16350 13014
rect 16780 13014 16796 13031
rect 17352 13031 17554 13048
rect 17612 13048 18572 13086
rect 17612 13031 17814 13048
rect 17352 13014 17368 13031
rect 16780 12998 17368 13014
rect 17798 13014 17814 13031
rect 18370 13031 18572 13048
rect 18630 13048 19590 13086
rect 18630 13031 18832 13048
rect 18370 13014 18386 13031
rect 17798 12998 18386 13014
rect 18816 13014 18832 13031
rect 19388 13031 19590 13048
rect 19648 13048 20608 13086
rect 19648 13031 19850 13048
rect 19388 13014 19404 13031
rect 18816 12998 19404 13014
rect 19834 13014 19850 13031
rect 20406 13031 20608 13048
rect 20666 13048 21626 13086
rect 20666 13031 20868 13048
rect 20406 13014 20422 13031
rect 19834 12998 20422 13014
rect 20852 13014 20868 13031
rect 21424 13031 21626 13048
rect 21684 13048 22644 13086
rect 21684 13031 21886 13048
rect 21424 13014 21440 13031
rect 20852 12998 21440 13014
rect 21870 13014 21886 13031
rect 22442 13031 22644 13048
rect 22702 13048 23662 13086
rect 22702 13031 22904 13048
rect 22442 13014 22458 13031
rect 21870 12998 22458 13014
rect 22888 13014 22904 13031
rect 23460 13031 23662 13048
rect 23720 13048 24680 13086
rect 23720 13031 23922 13048
rect 23460 13014 23476 13031
rect 22888 12998 23476 13014
rect 23906 13014 23922 13031
rect 24478 13031 24680 13048
rect 24738 13048 25698 13086
rect 24738 13031 24940 13048
rect 24478 13014 24494 13031
rect 23906 12998 24494 13014
rect 24924 13014 24940 13031
rect 25496 13031 25698 13048
rect 25756 13048 26716 13086
rect 25756 13031 25958 13048
rect 25496 13014 25512 13031
rect 24924 12998 25512 13014
rect 25942 13014 25958 13031
rect 26514 13031 26716 13048
rect 26774 13048 27734 13086
rect 26774 13031 26976 13048
rect 26514 13014 26530 13031
rect 25942 12998 26530 13014
rect 26960 13014 26976 13031
rect 27532 13031 27734 13048
rect 27792 13048 28752 13086
rect 27792 13031 27994 13048
rect 27532 13014 27548 13031
rect 26960 12998 27548 13014
rect 27978 13014 27994 13031
rect 28550 13031 28752 13048
rect 28810 13048 29770 13086
rect 28810 13031 29012 13048
rect 28550 13014 28566 13031
rect 27978 12998 28566 13014
rect 28996 13014 29012 13031
rect 29568 13031 29770 13048
rect 29828 13048 30788 13086
rect 29828 13031 30030 13048
rect 29568 13014 29584 13031
rect 28996 12998 29584 13014
rect 30014 13014 30030 13031
rect 30586 13031 30788 13048
rect 30846 13048 31806 13086
rect 30846 13031 31048 13048
rect 30586 13014 30602 13031
rect 30014 12998 30602 13014
rect 31032 13014 31048 13031
rect 31604 13031 31806 13048
rect 31864 13048 32824 13086
rect 31864 13031 32066 13048
rect 31604 13014 31620 13031
rect 31032 12998 31620 13014
rect 32050 13014 32066 13031
rect 32622 13031 32824 13048
rect 32882 13048 33842 13086
rect 32882 13031 33084 13048
rect 32622 13014 32638 13031
rect 32050 12998 32638 13014
rect 33068 13014 33084 13031
rect 33640 13031 33842 13048
rect 33640 13014 33656 13031
rect 33068 12998 33656 13014
rect 1774 12572 2734 12610
rect 1774 12555 1976 12572
rect 1960 12538 1976 12555
rect 2532 12555 2734 12572
rect 2792 12572 3752 12610
rect 2792 12555 2994 12572
rect 2532 12538 2548 12555
rect 1960 12522 2548 12538
rect 2978 12538 2994 12555
rect 3550 12555 3752 12572
rect 3810 12572 4770 12610
rect 3810 12555 4012 12572
rect 3550 12538 3566 12555
rect 2978 12522 3566 12538
rect 1960 12464 2548 12480
rect 1960 12447 1976 12464
rect 1774 12430 1976 12447
rect 2532 12447 2548 12464
rect 3996 12538 4012 12555
rect 4568 12555 4770 12572
rect 4828 12572 5788 12610
rect 4828 12555 5030 12572
rect 4568 12538 4584 12555
rect 3996 12522 4584 12538
rect 2978 12464 3566 12480
rect 2978 12447 2994 12464
rect 2532 12430 2734 12447
rect 1774 12392 2734 12430
rect 2792 12430 2994 12447
rect 3550 12447 3566 12464
rect 5014 12538 5030 12555
rect 5586 12555 5788 12572
rect 5846 12572 6806 12610
rect 5846 12555 6048 12572
rect 5586 12538 5602 12555
rect 5014 12522 5602 12538
rect 3996 12464 4584 12480
rect 3996 12447 4012 12464
rect 3550 12430 3752 12447
rect 2792 12392 3752 12430
rect 3810 12430 4012 12447
rect 4568 12447 4584 12464
rect 6032 12538 6048 12555
rect 6604 12555 6806 12572
rect 6864 12572 7824 12610
rect 6864 12555 7066 12572
rect 6604 12538 6620 12555
rect 6032 12522 6620 12538
rect 5014 12464 5602 12480
rect 5014 12447 5030 12464
rect 4568 12430 4770 12447
rect 3810 12392 4770 12430
rect 4828 12430 5030 12447
rect 5586 12447 5602 12464
rect 7050 12538 7066 12555
rect 7622 12555 7824 12572
rect 7882 12572 8842 12610
rect 7882 12555 8084 12572
rect 7622 12538 7638 12555
rect 7050 12522 7638 12538
rect 6032 12464 6620 12480
rect 6032 12447 6048 12464
rect 5586 12430 5788 12447
rect 4828 12392 5788 12430
rect 5846 12430 6048 12447
rect 6604 12447 6620 12464
rect 8068 12538 8084 12555
rect 8640 12555 8842 12572
rect 8900 12572 9860 12610
rect 8900 12555 9102 12572
rect 8640 12538 8656 12555
rect 8068 12522 8656 12538
rect 7050 12464 7638 12480
rect 7050 12447 7066 12464
rect 6604 12430 6806 12447
rect 5846 12392 6806 12430
rect 6864 12430 7066 12447
rect 7622 12447 7638 12464
rect 9086 12538 9102 12555
rect 9658 12555 9860 12572
rect 9918 12572 10878 12610
rect 9918 12555 10120 12572
rect 9658 12538 9674 12555
rect 9086 12522 9674 12538
rect 8068 12464 8656 12480
rect 8068 12447 8084 12464
rect 7622 12430 7824 12447
rect 6864 12392 7824 12430
rect 7882 12430 8084 12447
rect 8640 12447 8656 12464
rect 10104 12538 10120 12555
rect 10676 12555 10878 12572
rect 10676 12538 10692 12555
rect 10104 12522 10692 12538
rect 9086 12464 9674 12480
rect 9086 12447 9102 12464
rect 8640 12430 8842 12447
rect 7882 12392 8842 12430
rect 8900 12430 9102 12447
rect 9658 12447 9674 12464
rect 10104 12464 10692 12480
rect 10104 12447 10120 12464
rect 9658 12430 9860 12447
rect 8900 12392 9860 12430
rect 9918 12430 10120 12447
rect 10676 12447 10692 12464
rect 10676 12430 10878 12447
rect 9918 12392 10878 12430
rect 13726 12380 14314 12396
rect 13726 12363 13742 12380
rect 13540 12346 13742 12363
rect 14298 12363 14314 12380
rect 14744 12380 15332 12396
rect 14744 12363 14760 12380
rect 14298 12346 14500 12363
rect 13540 12308 14500 12346
rect 14558 12346 14760 12363
rect 15316 12363 15332 12380
rect 15762 12380 16350 12396
rect 15762 12363 15778 12380
rect 15316 12346 15518 12363
rect 14558 12308 15518 12346
rect 15576 12346 15778 12363
rect 16334 12363 16350 12380
rect 16780 12380 17368 12396
rect 16780 12363 16796 12380
rect 16334 12346 16536 12363
rect 15576 12308 16536 12346
rect 16594 12346 16796 12363
rect 17352 12363 17368 12380
rect 17798 12380 18386 12396
rect 17798 12363 17814 12380
rect 17352 12346 17554 12363
rect 16594 12308 17554 12346
rect 17612 12346 17814 12363
rect 18370 12363 18386 12380
rect 18816 12380 19404 12396
rect 18816 12363 18832 12380
rect 18370 12346 18572 12363
rect 17612 12308 18572 12346
rect 18630 12346 18832 12363
rect 19388 12363 19404 12380
rect 19834 12380 20422 12396
rect 19834 12363 19850 12380
rect 19388 12346 19590 12363
rect 18630 12308 19590 12346
rect 19648 12346 19850 12363
rect 20406 12363 20422 12380
rect 20852 12380 21440 12396
rect 20852 12363 20868 12380
rect 20406 12346 20608 12363
rect 19648 12308 20608 12346
rect 20666 12346 20868 12363
rect 21424 12363 21440 12380
rect 21870 12380 22458 12396
rect 21870 12363 21886 12380
rect 21424 12346 21626 12363
rect 20666 12308 21626 12346
rect 21684 12346 21886 12363
rect 22442 12363 22458 12380
rect 22888 12380 23476 12396
rect 22888 12363 22904 12380
rect 22442 12346 22644 12363
rect 21684 12308 22644 12346
rect 22702 12346 22904 12363
rect 23460 12363 23476 12380
rect 23906 12380 24494 12396
rect 23906 12363 23922 12380
rect 23460 12346 23662 12363
rect 22702 12308 23662 12346
rect 23720 12346 23922 12363
rect 24478 12363 24494 12380
rect 24924 12380 25512 12396
rect 24924 12363 24940 12380
rect 24478 12346 24680 12363
rect 23720 12308 24680 12346
rect 24738 12346 24940 12363
rect 25496 12363 25512 12380
rect 25942 12380 26530 12396
rect 25942 12363 25958 12380
rect 25496 12346 25698 12363
rect 24738 12308 25698 12346
rect 25756 12346 25958 12363
rect 26514 12363 26530 12380
rect 26960 12380 27548 12396
rect 26960 12363 26976 12380
rect 26514 12346 26716 12363
rect 25756 12308 26716 12346
rect 26774 12346 26976 12363
rect 27532 12363 27548 12380
rect 27978 12380 28566 12396
rect 27978 12363 27994 12380
rect 27532 12346 27734 12363
rect 26774 12308 27734 12346
rect 27792 12346 27994 12363
rect 28550 12363 28566 12380
rect 28996 12380 29584 12396
rect 28996 12363 29012 12380
rect 28550 12346 28752 12363
rect 27792 12308 28752 12346
rect 28810 12346 29012 12363
rect 29568 12363 29584 12380
rect 30014 12380 30602 12396
rect 30014 12363 30030 12380
rect 29568 12346 29770 12363
rect 28810 12308 29770 12346
rect 29828 12346 30030 12363
rect 30586 12363 30602 12380
rect 31032 12380 31620 12396
rect 31032 12363 31048 12380
rect 30586 12346 30788 12363
rect 29828 12308 30788 12346
rect 30846 12346 31048 12363
rect 31604 12363 31620 12380
rect 32050 12380 32638 12396
rect 32050 12363 32066 12380
rect 31604 12346 31806 12363
rect 30846 12308 31806 12346
rect 31864 12346 32066 12363
rect 32622 12363 32638 12380
rect 33068 12380 33656 12396
rect 33068 12363 33084 12380
rect 32622 12346 32824 12363
rect 31864 12308 32824 12346
rect 32882 12346 33084 12363
rect 33640 12363 33656 12380
rect 33640 12346 33842 12363
rect 32882 12308 33842 12346
rect 1774 11754 2734 11792
rect 1774 11737 1976 11754
rect 1960 11720 1976 11737
rect 2532 11737 2734 11754
rect 2792 11754 3752 11792
rect 2792 11737 2994 11754
rect 2532 11720 2548 11737
rect 1960 11704 2548 11720
rect 2978 11720 2994 11737
rect 3550 11737 3752 11754
rect 3810 11754 4770 11792
rect 3810 11737 4012 11754
rect 3550 11720 3566 11737
rect 2978 11704 3566 11720
rect 1960 11646 2548 11662
rect 1960 11629 1976 11646
rect 1774 11612 1976 11629
rect 2532 11629 2548 11646
rect 3996 11720 4012 11737
rect 4568 11737 4770 11754
rect 4828 11754 5788 11792
rect 4828 11737 5030 11754
rect 4568 11720 4584 11737
rect 3996 11704 4584 11720
rect 2978 11646 3566 11662
rect 2978 11629 2994 11646
rect 2532 11612 2734 11629
rect 1774 11574 2734 11612
rect 2792 11612 2994 11629
rect 3550 11629 3566 11646
rect 5014 11720 5030 11737
rect 5586 11737 5788 11754
rect 5846 11754 6806 11792
rect 5846 11737 6048 11754
rect 5586 11720 5602 11737
rect 5014 11704 5602 11720
rect 3996 11646 4584 11662
rect 3996 11629 4012 11646
rect 3550 11612 3752 11629
rect 2792 11574 3752 11612
rect 3810 11612 4012 11629
rect 4568 11629 4584 11646
rect 6032 11720 6048 11737
rect 6604 11737 6806 11754
rect 6864 11754 7824 11792
rect 6864 11737 7066 11754
rect 6604 11720 6620 11737
rect 6032 11704 6620 11720
rect 5014 11646 5602 11662
rect 5014 11629 5030 11646
rect 4568 11612 4770 11629
rect 3810 11574 4770 11612
rect 4828 11612 5030 11629
rect 5586 11629 5602 11646
rect 7050 11720 7066 11737
rect 7622 11737 7824 11754
rect 7882 11754 8842 11792
rect 7882 11737 8084 11754
rect 7622 11720 7638 11737
rect 7050 11704 7638 11720
rect 6032 11646 6620 11662
rect 6032 11629 6048 11646
rect 5586 11612 5788 11629
rect 4828 11574 5788 11612
rect 5846 11612 6048 11629
rect 6604 11629 6620 11646
rect 8068 11720 8084 11737
rect 8640 11737 8842 11754
rect 8900 11754 9860 11792
rect 8900 11737 9102 11754
rect 8640 11720 8656 11737
rect 8068 11704 8656 11720
rect 7050 11646 7638 11662
rect 7050 11629 7066 11646
rect 6604 11612 6806 11629
rect 5846 11574 6806 11612
rect 6864 11612 7066 11629
rect 7622 11629 7638 11646
rect 9086 11720 9102 11737
rect 9658 11737 9860 11754
rect 9918 11754 10878 11792
rect 9918 11737 10120 11754
rect 9658 11720 9674 11737
rect 9086 11704 9674 11720
rect 8068 11646 8656 11662
rect 8068 11629 8084 11646
rect 7622 11612 7824 11629
rect 6864 11574 7824 11612
rect 7882 11612 8084 11629
rect 8640 11629 8656 11646
rect 10104 11720 10120 11737
rect 10676 11737 10878 11754
rect 10676 11720 10692 11737
rect 10104 11704 10692 11720
rect 9086 11646 9674 11662
rect 9086 11629 9102 11646
rect 8640 11612 8842 11629
rect 7882 11574 8842 11612
rect 8900 11612 9102 11629
rect 9658 11629 9674 11646
rect 10104 11646 10692 11662
rect 10104 11629 10120 11646
rect 9658 11612 9860 11629
rect 8900 11574 9860 11612
rect 9918 11612 10120 11629
rect 10676 11629 10692 11646
rect 13540 11670 14500 11708
rect 13540 11653 13742 11670
rect 13726 11636 13742 11653
rect 14298 11653 14500 11670
rect 14558 11670 15518 11708
rect 14558 11653 14760 11670
rect 14298 11636 14314 11653
rect 10676 11612 10878 11629
rect 13726 11620 14314 11636
rect 14744 11636 14760 11653
rect 15316 11653 15518 11670
rect 15576 11670 16536 11708
rect 15576 11653 15778 11670
rect 15316 11636 15332 11653
rect 14744 11620 15332 11636
rect 15762 11636 15778 11653
rect 16334 11653 16536 11670
rect 16594 11670 17554 11708
rect 16594 11653 16796 11670
rect 16334 11636 16350 11653
rect 15762 11620 16350 11636
rect 16780 11636 16796 11653
rect 17352 11653 17554 11670
rect 17612 11670 18572 11708
rect 17612 11653 17814 11670
rect 17352 11636 17368 11653
rect 16780 11620 17368 11636
rect 17798 11636 17814 11653
rect 18370 11653 18572 11670
rect 18630 11670 19590 11708
rect 18630 11653 18832 11670
rect 18370 11636 18386 11653
rect 17798 11620 18386 11636
rect 18816 11636 18832 11653
rect 19388 11653 19590 11670
rect 19648 11670 20608 11708
rect 19648 11653 19850 11670
rect 19388 11636 19404 11653
rect 18816 11620 19404 11636
rect 19834 11636 19850 11653
rect 20406 11653 20608 11670
rect 20666 11670 21626 11708
rect 20666 11653 20868 11670
rect 20406 11636 20422 11653
rect 19834 11620 20422 11636
rect 20852 11636 20868 11653
rect 21424 11653 21626 11670
rect 21684 11670 22644 11708
rect 21684 11653 21886 11670
rect 21424 11636 21440 11653
rect 20852 11620 21440 11636
rect 21870 11636 21886 11653
rect 22442 11653 22644 11670
rect 22702 11670 23662 11708
rect 22702 11653 22904 11670
rect 22442 11636 22458 11653
rect 21870 11620 22458 11636
rect 22888 11636 22904 11653
rect 23460 11653 23662 11670
rect 23720 11670 24680 11708
rect 23720 11653 23922 11670
rect 23460 11636 23476 11653
rect 22888 11620 23476 11636
rect 23906 11636 23922 11653
rect 24478 11653 24680 11670
rect 24738 11670 25698 11708
rect 24738 11653 24940 11670
rect 24478 11636 24494 11653
rect 23906 11620 24494 11636
rect 24924 11636 24940 11653
rect 25496 11653 25698 11670
rect 25756 11670 26716 11708
rect 25756 11653 25958 11670
rect 25496 11636 25512 11653
rect 24924 11620 25512 11636
rect 25942 11636 25958 11653
rect 26514 11653 26716 11670
rect 26774 11670 27734 11708
rect 26774 11653 26976 11670
rect 26514 11636 26530 11653
rect 25942 11620 26530 11636
rect 26960 11636 26976 11653
rect 27532 11653 27734 11670
rect 27792 11670 28752 11708
rect 27792 11653 27994 11670
rect 27532 11636 27548 11653
rect 26960 11620 27548 11636
rect 27978 11636 27994 11653
rect 28550 11653 28752 11670
rect 28810 11670 29770 11708
rect 28810 11653 29012 11670
rect 28550 11636 28566 11653
rect 27978 11620 28566 11636
rect 28996 11636 29012 11653
rect 29568 11653 29770 11670
rect 29828 11670 30788 11708
rect 29828 11653 30030 11670
rect 29568 11636 29584 11653
rect 28996 11620 29584 11636
rect 30014 11636 30030 11653
rect 30586 11653 30788 11670
rect 30846 11670 31806 11708
rect 30846 11653 31048 11670
rect 30586 11636 30602 11653
rect 30014 11620 30602 11636
rect 31032 11636 31048 11653
rect 31604 11653 31806 11670
rect 31864 11670 32824 11708
rect 31864 11653 32066 11670
rect 31604 11636 31620 11653
rect 31032 11620 31620 11636
rect 32050 11636 32066 11653
rect 32622 11653 32824 11670
rect 32882 11670 33842 11708
rect 32882 11653 33084 11670
rect 32622 11636 32638 11653
rect 32050 11620 32638 11636
rect 33068 11636 33084 11653
rect 33640 11653 33842 11670
rect 33640 11636 33656 11653
rect 33068 11620 33656 11636
rect 9918 11574 10878 11612
rect 13726 11148 14314 11164
rect 13726 11131 13742 11148
rect 13540 11114 13742 11131
rect 14298 11131 14314 11148
rect 14744 11148 15332 11164
rect 14744 11131 14760 11148
rect 14298 11114 14500 11131
rect 13540 11076 14500 11114
rect 14558 11114 14760 11131
rect 15316 11131 15332 11148
rect 15762 11148 16350 11164
rect 15762 11131 15778 11148
rect 15316 11114 15518 11131
rect 14558 11076 15518 11114
rect 15576 11114 15778 11131
rect 16334 11131 16350 11148
rect 16780 11148 17368 11164
rect 16780 11131 16796 11148
rect 16334 11114 16536 11131
rect 15576 11076 16536 11114
rect 16594 11114 16796 11131
rect 17352 11131 17368 11148
rect 17798 11148 18386 11164
rect 17798 11131 17814 11148
rect 17352 11114 17554 11131
rect 16594 11076 17554 11114
rect 17612 11114 17814 11131
rect 18370 11131 18386 11148
rect 18816 11148 19404 11164
rect 18816 11131 18832 11148
rect 18370 11114 18572 11131
rect 17612 11076 18572 11114
rect 18630 11114 18832 11131
rect 19388 11131 19404 11148
rect 19834 11148 20422 11164
rect 19834 11131 19850 11148
rect 19388 11114 19590 11131
rect 18630 11076 19590 11114
rect 19648 11114 19850 11131
rect 20406 11131 20422 11148
rect 20852 11148 21440 11164
rect 20852 11131 20868 11148
rect 20406 11114 20608 11131
rect 19648 11076 20608 11114
rect 20666 11114 20868 11131
rect 21424 11131 21440 11148
rect 21870 11148 22458 11164
rect 21870 11131 21886 11148
rect 21424 11114 21626 11131
rect 20666 11076 21626 11114
rect 21684 11114 21886 11131
rect 22442 11131 22458 11148
rect 22888 11148 23476 11164
rect 22888 11131 22904 11148
rect 22442 11114 22644 11131
rect 21684 11076 22644 11114
rect 22702 11114 22904 11131
rect 23460 11131 23476 11148
rect 23906 11148 24494 11164
rect 23906 11131 23922 11148
rect 23460 11114 23662 11131
rect 22702 11076 23662 11114
rect 23720 11114 23922 11131
rect 24478 11131 24494 11148
rect 24924 11148 25512 11164
rect 24924 11131 24940 11148
rect 24478 11114 24680 11131
rect 23720 11076 24680 11114
rect 24738 11114 24940 11131
rect 25496 11131 25512 11148
rect 25942 11148 26530 11164
rect 25942 11131 25958 11148
rect 25496 11114 25698 11131
rect 24738 11076 25698 11114
rect 25756 11114 25958 11131
rect 26514 11131 26530 11148
rect 26960 11148 27548 11164
rect 26960 11131 26976 11148
rect 26514 11114 26716 11131
rect 25756 11076 26716 11114
rect 26774 11114 26976 11131
rect 27532 11131 27548 11148
rect 27978 11148 28566 11164
rect 27978 11131 27994 11148
rect 27532 11114 27734 11131
rect 26774 11076 27734 11114
rect 27792 11114 27994 11131
rect 28550 11131 28566 11148
rect 28996 11148 29584 11164
rect 28996 11131 29012 11148
rect 28550 11114 28752 11131
rect 27792 11076 28752 11114
rect 28810 11114 29012 11131
rect 29568 11131 29584 11148
rect 30014 11148 30602 11164
rect 30014 11131 30030 11148
rect 29568 11114 29770 11131
rect 28810 11076 29770 11114
rect 29828 11114 30030 11131
rect 30586 11131 30602 11148
rect 31032 11148 31620 11164
rect 31032 11131 31048 11148
rect 30586 11114 30788 11131
rect 29828 11076 30788 11114
rect 30846 11114 31048 11131
rect 31604 11131 31620 11148
rect 32050 11148 32638 11164
rect 32050 11131 32066 11148
rect 31604 11114 31806 11131
rect 30846 11076 31806 11114
rect 31864 11114 32066 11131
rect 32622 11131 32638 11148
rect 33068 11148 33656 11164
rect 33068 11131 33084 11148
rect 32622 11114 32824 11131
rect 31864 11076 32824 11114
rect 32882 11114 33084 11131
rect 33640 11131 33656 11148
rect 33640 11114 33842 11131
rect 32882 11076 33842 11114
rect 1774 10936 2734 10974
rect 1774 10919 1976 10936
rect 1960 10902 1976 10919
rect 2532 10919 2734 10936
rect 2792 10936 3752 10974
rect 2792 10919 2994 10936
rect 2532 10902 2548 10919
rect 1960 10886 2548 10902
rect 2978 10902 2994 10919
rect 3550 10919 3752 10936
rect 3810 10936 4770 10974
rect 3810 10919 4012 10936
rect 3550 10902 3566 10919
rect 2978 10886 3566 10902
rect 1960 10828 2548 10844
rect 1960 10811 1976 10828
rect 1774 10794 1976 10811
rect 2532 10811 2548 10828
rect 3996 10902 4012 10919
rect 4568 10919 4770 10936
rect 4828 10936 5788 10974
rect 4828 10919 5030 10936
rect 4568 10902 4584 10919
rect 3996 10886 4584 10902
rect 2978 10828 3566 10844
rect 2978 10811 2994 10828
rect 2532 10794 2734 10811
rect 1774 10756 2734 10794
rect 2792 10794 2994 10811
rect 3550 10811 3566 10828
rect 5014 10902 5030 10919
rect 5586 10919 5788 10936
rect 5846 10936 6806 10974
rect 5846 10919 6048 10936
rect 5586 10902 5602 10919
rect 5014 10886 5602 10902
rect 3996 10828 4584 10844
rect 3996 10811 4012 10828
rect 3550 10794 3752 10811
rect 2792 10756 3752 10794
rect 3810 10794 4012 10811
rect 4568 10811 4584 10828
rect 6032 10902 6048 10919
rect 6604 10919 6806 10936
rect 6864 10936 7824 10974
rect 6864 10919 7066 10936
rect 6604 10902 6620 10919
rect 6032 10886 6620 10902
rect 5014 10828 5602 10844
rect 5014 10811 5030 10828
rect 4568 10794 4770 10811
rect 3810 10756 4770 10794
rect 4828 10794 5030 10811
rect 5586 10811 5602 10828
rect 7050 10902 7066 10919
rect 7622 10919 7824 10936
rect 7882 10936 8842 10974
rect 7882 10919 8084 10936
rect 7622 10902 7638 10919
rect 7050 10886 7638 10902
rect 6032 10828 6620 10844
rect 6032 10811 6048 10828
rect 5586 10794 5788 10811
rect 4828 10756 5788 10794
rect 5846 10794 6048 10811
rect 6604 10811 6620 10828
rect 8068 10902 8084 10919
rect 8640 10919 8842 10936
rect 8900 10936 9860 10974
rect 8900 10919 9102 10936
rect 8640 10902 8656 10919
rect 8068 10886 8656 10902
rect 7050 10828 7638 10844
rect 7050 10811 7066 10828
rect 6604 10794 6806 10811
rect 5846 10756 6806 10794
rect 6864 10794 7066 10811
rect 7622 10811 7638 10828
rect 9086 10902 9102 10919
rect 9658 10919 9860 10936
rect 9918 10936 10878 10974
rect 9918 10919 10120 10936
rect 9658 10902 9674 10919
rect 9086 10886 9674 10902
rect 8068 10828 8656 10844
rect 8068 10811 8084 10828
rect 7622 10794 7824 10811
rect 6864 10756 7824 10794
rect 7882 10794 8084 10811
rect 8640 10811 8656 10828
rect 10104 10902 10120 10919
rect 10676 10919 10878 10936
rect 10676 10902 10692 10919
rect 10104 10886 10692 10902
rect 9086 10828 9674 10844
rect 9086 10811 9102 10828
rect 8640 10794 8842 10811
rect 7882 10756 8842 10794
rect 8900 10794 9102 10811
rect 9658 10811 9674 10828
rect 10104 10828 10692 10844
rect 10104 10811 10120 10828
rect 9658 10794 9860 10811
rect 8900 10756 9860 10794
rect 9918 10794 10120 10811
rect 10676 10811 10692 10828
rect 10676 10794 10878 10811
rect 9918 10756 10878 10794
rect 13540 10438 14500 10476
rect 13540 10421 13742 10438
rect 13726 10404 13742 10421
rect 14298 10421 14500 10438
rect 14558 10438 15518 10476
rect 14558 10421 14760 10438
rect 14298 10404 14314 10421
rect 13726 10388 14314 10404
rect 14744 10404 14760 10421
rect 15316 10421 15518 10438
rect 15576 10438 16536 10476
rect 15576 10421 15778 10438
rect 15316 10404 15332 10421
rect 14744 10388 15332 10404
rect 15762 10404 15778 10421
rect 16334 10421 16536 10438
rect 16594 10438 17554 10476
rect 16594 10421 16796 10438
rect 16334 10404 16350 10421
rect 15762 10388 16350 10404
rect 16780 10404 16796 10421
rect 17352 10421 17554 10438
rect 17612 10438 18572 10476
rect 17612 10421 17814 10438
rect 17352 10404 17368 10421
rect 16780 10388 17368 10404
rect 17798 10404 17814 10421
rect 18370 10421 18572 10438
rect 18630 10438 19590 10476
rect 18630 10421 18832 10438
rect 18370 10404 18386 10421
rect 17798 10388 18386 10404
rect 18816 10404 18832 10421
rect 19388 10421 19590 10438
rect 19648 10438 20608 10476
rect 19648 10421 19850 10438
rect 19388 10404 19404 10421
rect 18816 10388 19404 10404
rect 19834 10404 19850 10421
rect 20406 10421 20608 10438
rect 20666 10438 21626 10476
rect 20666 10421 20868 10438
rect 20406 10404 20422 10421
rect 19834 10388 20422 10404
rect 20852 10404 20868 10421
rect 21424 10421 21626 10438
rect 21684 10438 22644 10476
rect 21684 10421 21886 10438
rect 21424 10404 21440 10421
rect 20852 10388 21440 10404
rect 21870 10404 21886 10421
rect 22442 10421 22644 10438
rect 22702 10438 23662 10476
rect 22702 10421 22904 10438
rect 22442 10404 22458 10421
rect 21870 10388 22458 10404
rect 22888 10404 22904 10421
rect 23460 10421 23662 10438
rect 23720 10438 24680 10476
rect 23720 10421 23922 10438
rect 23460 10404 23476 10421
rect 22888 10388 23476 10404
rect 23906 10404 23922 10421
rect 24478 10421 24680 10438
rect 24738 10438 25698 10476
rect 24738 10421 24940 10438
rect 24478 10404 24494 10421
rect 23906 10388 24494 10404
rect 24924 10404 24940 10421
rect 25496 10421 25698 10438
rect 25756 10438 26716 10476
rect 25756 10421 25958 10438
rect 25496 10404 25512 10421
rect 24924 10388 25512 10404
rect 25942 10404 25958 10421
rect 26514 10421 26716 10438
rect 26774 10438 27734 10476
rect 26774 10421 26976 10438
rect 26514 10404 26530 10421
rect 25942 10388 26530 10404
rect 26960 10404 26976 10421
rect 27532 10421 27734 10438
rect 27792 10438 28752 10476
rect 27792 10421 27994 10438
rect 27532 10404 27548 10421
rect 26960 10388 27548 10404
rect 27978 10404 27994 10421
rect 28550 10421 28752 10438
rect 28810 10438 29770 10476
rect 28810 10421 29012 10438
rect 28550 10404 28566 10421
rect 27978 10388 28566 10404
rect 28996 10404 29012 10421
rect 29568 10421 29770 10438
rect 29828 10438 30788 10476
rect 29828 10421 30030 10438
rect 29568 10404 29584 10421
rect 28996 10388 29584 10404
rect 30014 10404 30030 10421
rect 30586 10421 30788 10438
rect 30846 10438 31806 10476
rect 30846 10421 31048 10438
rect 30586 10404 30602 10421
rect 30014 10388 30602 10404
rect 31032 10404 31048 10421
rect 31604 10421 31806 10438
rect 31864 10438 32824 10476
rect 31864 10421 32066 10438
rect 31604 10404 31620 10421
rect 31032 10388 31620 10404
rect 32050 10404 32066 10421
rect 32622 10421 32824 10438
rect 32882 10438 33842 10476
rect 32882 10421 33084 10438
rect 32622 10404 32638 10421
rect 32050 10388 32638 10404
rect 33068 10404 33084 10421
rect 33640 10421 33842 10438
rect 33640 10404 33656 10421
rect 33068 10388 33656 10404
rect 1774 10118 2734 10156
rect 1774 10101 1976 10118
rect 1960 10084 1976 10101
rect 2532 10101 2734 10118
rect 2792 10118 3752 10156
rect 2792 10101 2994 10118
rect 2532 10084 2548 10101
rect 1960 10068 2548 10084
rect 2978 10084 2994 10101
rect 3550 10101 3752 10118
rect 3810 10118 4770 10156
rect 3810 10101 4012 10118
rect 3550 10084 3566 10101
rect 2978 10068 3566 10084
rect 1960 10010 2548 10026
rect 1960 9993 1976 10010
rect 1774 9976 1976 9993
rect 2532 9993 2548 10010
rect 3996 10084 4012 10101
rect 4568 10101 4770 10118
rect 4828 10118 5788 10156
rect 4828 10101 5030 10118
rect 4568 10084 4584 10101
rect 3996 10068 4584 10084
rect 2978 10010 3566 10026
rect 2978 9993 2994 10010
rect 2532 9976 2734 9993
rect 1774 9938 2734 9976
rect 2792 9976 2994 9993
rect 3550 9993 3566 10010
rect 5014 10084 5030 10101
rect 5586 10101 5788 10118
rect 5846 10118 6806 10156
rect 5846 10101 6048 10118
rect 5586 10084 5602 10101
rect 5014 10068 5602 10084
rect 3996 10010 4584 10026
rect 3996 9993 4012 10010
rect 3550 9976 3752 9993
rect 2792 9938 3752 9976
rect 3810 9976 4012 9993
rect 4568 9993 4584 10010
rect 6032 10084 6048 10101
rect 6604 10101 6806 10118
rect 6864 10118 7824 10156
rect 6864 10101 7066 10118
rect 6604 10084 6620 10101
rect 6032 10068 6620 10084
rect 5014 10010 5602 10026
rect 5014 9993 5030 10010
rect 4568 9976 4770 9993
rect 3810 9938 4770 9976
rect 4828 9976 5030 9993
rect 5586 9993 5602 10010
rect 7050 10084 7066 10101
rect 7622 10101 7824 10118
rect 7882 10118 8842 10156
rect 7882 10101 8084 10118
rect 7622 10084 7638 10101
rect 7050 10068 7638 10084
rect 6032 10010 6620 10026
rect 6032 9993 6048 10010
rect 5586 9976 5788 9993
rect 4828 9938 5788 9976
rect 5846 9976 6048 9993
rect 6604 9993 6620 10010
rect 8068 10084 8084 10101
rect 8640 10101 8842 10118
rect 8900 10118 9860 10156
rect 8900 10101 9102 10118
rect 8640 10084 8656 10101
rect 8068 10068 8656 10084
rect 7050 10010 7638 10026
rect 7050 9993 7066 10010
rect 6604 9976 6806 9993
rect 5846 9938 6806 9976
rect 6864 9976 7066 9993
rect 7622 9993 7638 10010
rect 9086 10084 9102 10101
rect 9658 10101 9860 10118
rect 9918 10118 10878 10156
rect 9918 10101 10120 10118
rect 9658 10084 9674 10101
rect 9086 10068 9674 10084
rect 8068 10010 8656 10026
rect 8068 9993 8084 10010
rect 7622 9976 7824 9993
rect 6864 9938 7824 9976
rect 7882 9976 8084 9993
rect 8640 9993 8656 10010
rect 10104 10084 10120 10101
rect 10676 10101 10878 10118
rect 10676 10084 10692 10101
rect 10104 10068 10692 10084
rect 9086 10010 9674 10026
rect 9086 9993 9102 10010
rect 8640 9976 8842 9993
rect 7882 9938 8842 9976
rect 8900 9976 9102 9993
rect 9658 9993 9674 10010
rect 10104 10010 10692 10026
rect 10104 9993 10120 10010
rect 9658 9976 9860 9993
rect 8900 9938 9860 9976
rect 9918 9976 10120 9993
rect 10676 9993 10692 10010
rect 10676 9976 10878 9993
rect 9918 9938 10878 9976
rect 13724 9914 14312 9930
rect 13724 9897 13740 9914
rect 13538 9880 13740 9897
rect 14296 9897 14312 9914
rect 14742 9914 15330 9930
rect 14742 9897 14758 9914
rect 14296 9880 14498 9897
rect 13538 9842 14498 9880
rect 14556 9880 14758 9897
rect 15314 9897 15330 9914
rect 15760 9914 16348 9930
rect 15760 9897 15776 9914
rect 15314 9880 15516 9897
rect 14556 9842 15516 9880
rect 15574 9880 15776 9897
rect 16332 9897 16348 9914
rect 16778 9914 17366 9930
rect 16778 9897 16794 9914
rect 16332 9880 16534 9897
rect 15574 9842 16534 9880
rect 16592 9880 16794 9897
rect 17350 9897 17366 9914
rect 17796 9914 18384 9930
rect 17796 9897 17812 9914
rect 17350 9880 17552 9897
rect 16592 9842 17552 9880
rect 17610 9880 17812 9897
rect 18368 9897 18384 9914
rect 18814 9914 19402 9930
rect 18814 9897 18830 9914
rect 18368 9880 18570 9897
rect 17610 9842 18570 9880
rect 18628 9880 18830 9897
rect 19386 9897 19402 9914
rect 19832 9914 20420 9930
rect 19832 9897 19848 9914
rect 19386 9880 19588 9897
rect 18628 9842 19588 9880
rect 19646 9880 19848 9897
rect 20404 9897 20420 9914
rect 20850 9914 21438 9930
rect 20850 9897 20866 9914
rect 20404 9880 20606 9897
rect 19646 9842 20606 9880
rect 20664 9880 20866 9897
rect 21422 9897 21438 9914
rect 21868 9914 22456 9930
rect 21868 9897 21884 9914
rect 21422 9880 21624 9897
rect 20664 9842 21624 9880
rect 21682 9880 21884 9897
rect 22440 9897 22456 9914
rect 22886 9914 23474 9930
rect 22886 9897 22902 9914
rect 22440 9880 22642 9897
rect 21682 9842 22642 9880
rect 22700 9880 22902 9897
rect 23458 9897 23474 9914
rect 23904 9914 24492 9930
rect 23904 9897 23920 9914
rect 23458 9880 23660 9897
rect 22700 9842 23660 9880
rect 23718 9880 23920 9897
rect 24476 9897 24492 9914
rect 24922 9914 25510 9930
rect 24922 9897 24938 9914
rect 24476 9880 24678 9897
rect 23718 9842 24678 9880
rect 24736 9880 24938 9897
rect 25494 9897 25510 9914
rect 25940 9914 26528 9930
rect 25940 9897 25956 9914
rect 25494 9880 25696 9897
rect 24736 9842 25696 9880
rect 25754 9880 25956 9897
rect 26512 9897 26528 9914
rect 26958 9914 27546 9930
rect 26958 9897 26974 9914
rect 26512 9880 26714 9897
rect 25754 9842 26714 9880
rect 26772 9880 26974 9897
rect 27530 9897 27546 9914
rect 27976 9914 28564 9930
rect 27976 9897 27992 9914
rect 27530 9880 27732 9897
rect 26772 9842 27732 9880
rect 27790 9880 27992 9897
rect 28548 9897 28564 9914
rect 28994 9914 29582 9930
rect 28994 9897 29010 9914
rect 28548 9880 28750 9897
rect 27790 9842 28750 9880
rect 28808 9880 29010 9897
rect 29566 9897 29582 9914
rect 30012 9914 30600 9930
rect 30012 9897 30028 9914
rect 29566 9880 29768 9897
rect 28808 9842 29768 9880
rect 29826 9880 30028 9897
rect 30584 9897 30600 9914
rect 31030 9914 31618 9930
rect 31030 9897 31046 9914
rect 30584 9880 30786 9897
rect 29826 9842 30786 9880
rect 30844 9880 31046 9897
rect 31602 9897 31618 9914
rect 32048 9914 32636 9930
rect 32048 9897 32064 9914
rect 31602 9880 31804 9897
rect 30844 9842 31804 9880
rect 31862 9880 32064 9897
rect 32620 9897 32636 9914
rect 33066 9914 33654 9930
rect 33066 9897 33082 9914
rect 32620 9880 32822 9897
rect 31862 9842 32822 9880
rect 32880 9880 33082 9897
rect 33638 9897 33654 9914
rect 33638 9880 33840 9897
rect 32880 9842 33840 9880
rect 1774 9300 2734 9338
rect 1774 9283 1976 9300
rect 1960 9266 1976 9283
rect 2532 9283 2734 9300
rect 2792 9300 3752 9338
rect 2792 9283 2994 9300
rect 2532 9266 2548 9283
rect 1960 9250 2548 9266
rect 2978 9266 2994 9283
rect 3550 9283 3752 9300
rect 3810 9300 4770 9338
rect 3810 9283 4012 9300
rect 3550 9266 3566 9283
rect 2978 9250 3566 9266
rect 1960 9192 2548 9208
rect 1960 9175 1976 9192
rect 1774 9158 1976 9175
rect 2532 9175 2548 9192
rect 3996 9266 4012 9283
rect 4568 9283 4770 9300
rect 4828 9300 5788 9338
rect 4828 9283 5030 9300
rect 4568 9266 4584 9283
rect 3996 9250 4584 9266
rect 2978 9192 3566 9208
rect 2978 9175 2994 9192
rect 2532 9158 2734 9175
rect 1774 9120 2734 9158
rect 2792 9158 2994 9175
rect 3550 9175 3566 9192
rect 5014 9266 5030 9283
rect 5586 9283 5788 9300
rect 5846 9300 6806 9338
rect 5846 9283 6048 9300
rect 5586 9266 5602 9283
rect 5014 9250 5602 9266
rect 3996 9192 4584 9208
rect 3996 9175 4012 9192
rect 3550 9158 3752 9175
rect 2792 9120 3752 9158
rect 3810 9158 4012 9175
rect 4568 9175 4584 9192
rect 6032 9266 6048 9283
rect 6604 9283 6806 9300
rect 6864 9300 7824 9338
rect 6864 9283 7066 9300
rect 6604 9266 6620 9283
rect 6032 9250 6620 9266
rect 5014 9192 5602 9208
rect 5014 9175 5030 9192
rect 4568 9158 4770 9175
rect 3810 9120 4770 9158
rect 4828 9158 5030 9175
rect 5586 9175 5602 9192
rect 7050 9266 7066 9283
rect 7622 9283 7824 9300
rect 7882 9300 8842 9338
rect 7882 9283 8084 9300
rect 7622 9266 7638 9283
rect 7050 9250 7638 9266
rect 6032 9192 6620 9208
rect 6032 9175 6048 9192
rect 5586 9158 5788 9175
rect 4828 9120 5788 9158
rect 5846 9158 6048 9175
rect 6604 9175 6620 9192
rect 8068 9266 8084 9283
rect 8640 9283 8842 9300
rect 8900 9300 9860 9338
rect 8900 9283 9102 9300
rect 8640 9266 8656 9283
rect 8068 9250 8656 9266
rect 7050 9192 7638 9208
rect 7050 9175 7066 9192
rect 6604 9158 6806 9175
rect 5846 9120 6806 9158
rect 6864 9158 7066 9175
rect 7622 9175 7638 9192
rect 9086 9266 9102 9283
rect 9658 9283 9860 9300
rect 9918 9300 10878 9338
rect 9918 9283 10120 9300
rect 9658 9266 9674 9283
rect 9086 9250 9674 9266
rect 8068 9192 8656 9208
rect 8068 9175 8084 9192
rect 7622 9158 7824 9175
rect 6864 9120 7824 9158
rect 7882 9158 8084 9175
rect 8640 9175 8656 9192
rect 10104 9266 10120 9283
rect 10676 9283 10878 9300
rect 10676 9266 10692 9283
rect 10104 9250 10692 9266
rect 9086 9192 9674 9208
rect 9086 9175 9102 9192
rect 8640 9158 8842 9175
rect 7882 9120 8842 9158
rect 8900 9158 9102 9175
rect 9658 9175 9674 9192
rect 10104 9192 10692 9208
rect 10104 9175 10120 9192
rect 9658 9158 9860 9175
rect 8900 9120 9860 9158
rect 9918 9158 10120 9175
rect 10676 9175 10692 9192
rect 13538 9204 14498 9242
rect 13538 9187 13740 9204
rect 10676 9158 10878 9175
rect 9918 9120 10878 9158
rect 13724 9170 13740 9187
rect 14296 9187 14498 9204
rect 14556 9204 15516 9242
rect 14556 9187 14758 9204
rect 14296 9170 14312 9187
rect 13724 9154 14312 9170
rect 14742 9170 14758 9187
rect 15314 9187 15516 9204
rect 15574 9204 16534 9242
rect 15574 9187 15776 9204
rect 15314 9170 15330 9187
rect 14742 9154 15330 9170
rect 15760 9170 15776 9187
rect 16332 9187 16534 9204
rect 16592 9204 17552 9242
rect 16592 9187 16794 9204
rect 16332 9170 16348 9187
rect 15760 9154 16348 9170
rect 16778 9170 16794 9187
rect 17350 9187 17552 9204
rect 17610 9204 18570 9242
rect 17610 9187 17812 9204
rect 17350 9170 17366 9187
rect 16778 9154 17366 9170
rect 17796 9170 17812 9187
rect 18368 9187 18570 9204
rect 18628 9204 19588 9242
rect 18628 9187 18830 9204
rect 18368 9170 18384 9187
rect 17796 9154 18384 9170
rect 18814 9170 18830 9187
rect 19386 9187 19588 9204
rect 19646 9204 20606 9242
rect 19646 9187 19848 9204
rect 19386 9170 19402 9187
rect 18814 9154 19402 9170
rect 19832 9170 19848 9187
rect 20404 9187 20606 9204
rect 20664 9204 21624 9242
rect 20664 9187 20866 9204
rect 20404 9170 20420 9187
rect 19832 9154 20420 9170
rect 20850 9170 20866 9187
rect 21422 9187 21624 9204
rect 21682 9204 22642 9242
rect 21682 9187 21884 9204
rect 21422 9170 21438 9187
rect 20850 9154 21438 9170
rect 21868 9170 21884 9187
rect 22440 9187 22642 9204
rect 22700 9204 23660 9242
rect 22700 9187 22902 9204
rect 22440 9170 22456 9187
rect 21868 9154 22456 9170
rect 22886 9170 22902 9187
rect 23458 9187 23660 9204
rect 23718 9204 24678 9242
rect 23718 9187 23920 9204
rect 23458 9170 23474 9187
rect 22886 9154 23474 9170
rect 23904 9170 23920 9187
rect 24476 9187 24678 9204
rect 24736 9204 25696 9242
rect 24736 9187 24938 9204
rect 24476 9170 24492 9187
rect 23904 9154 24492 9170
rect 24922 9170 24938 9187
rect 25494 9187 25696 9204
rect 25754 9204 26714 9242
rect 25754 9187 25956 9204
rect 25494 9170 25510 9187
rect 24922 9154 25510 9170
rect 25940 9170 25956 9187
rect 26512 9187 26714 9204
rect 26772 9204 27732 9242
rect 26772 9187 26974 9204
rect 26512 9170 26528 9187
rect 25940 9154 26528 9170
rect 26958 9170 26974 9187
rect 27530 9187 27732 9204
rect 27790 9204 28750 9242
rect 27790 9187 27992 9204
rect 27530 9170 27546 9187
rect 26958 9154 27546 9170
rect 27976 9170 27992 9187
rect 28548 9187 28750 9204
rect 28808 9204 29768 9242
rect 28808 9187 29010 9204
rect 28548 9170 28564 9187
rect 27976 9154 28564 9170
rect 28994 9170 29010 9187
rect 29566 9187 29768 9204
rect 29826 9204 30786 9242
rect 29826 9187 30028 9204
rect 29566 9170 29582 9187
rect 28994 9154 29582 9170
rect 30012 9170 30028 9187
rect 30584 9187 30786 9204
rect 30844 9204 31804 9242
rect 30844 9187 31046 9204
rect 30584 9170 30600 9187
rect 30012 9154 30600 9170
rect 31030 9170 31046 9187
rect 31602 9187 31804 9204
rect 31862 9204 32822 9242
rect 31862 9187 32064 9204
rect 31602 9170 31618 9187
rect 31030 9154 31618 9170
rect 32048 9170 32064 9187
rect 32620 9187 32822 9204
rect 32880 9204 33840 9242
rect 32880 9187 33082 9204
rect 32620 9170 32636 9187
rect 32048 9154 32636 9170
rect 33066 9170 33082 9187
rect 33638 9187 33840 9204
rect 33638 9170 33654 9187
rect 33066 9154 33654 9170
rect 13724 8680 14312 8696
rect 13724 8663 13740 8680
rect 13538 8646 13740 8663
rect 14296 8663 14312 8680
rect 14742 8680 15330 8696
rect 14742 8663 14758 8680
rect 14296 8646 14498 8663
rect 13538 8608 14498 8646
rect 14556 8646 14758 8663
rect 15314 8663 15330 8680
rect 15760 8680 16348 8696
rect 15760 8663 15776 8680
rect 15314 8646 15516 8663
rect 14556 8608 15516 8646
rect 15574 8646 15776 8663
rect 16332 8663 16348 8680
rect 16778 8680 17366 8696
rect 16778 8663 16794 8680
rect 16332 8646 16534 8663
rect 15574 8608 16534 8646
rect 16592 8646 16794 8663
rect 17350 8663 17366 8680
rect 17796 8680 18384 8696
rect 17796 8663 17812 8680
rect 17350 8646 17552 8663
rect 16592 8608 17552 8646
rect 17610 8646 17812 8663
rect 18368 8663 18384 8680
rect 18814 8680 19402 8696
rect 18814 8663 18830 8680
rect 18368 8646 18570 8663
rect 17610 8608 18570 8646
rect 18628 8646 18830 8663
rect 19386 8663 19402 8680
rect 19832 8680 20420 8696
rect 19832 8663 19848 8680
rect 19386 8646 19588 8663
rect 18628 8608 19588 8646
rect 19646 8646 19848 8663
rect 20404 8663 20420 8680
rect 20850 8680 21438 8696
rect 20850 8663 20866 8680
rect 20404 8646 20606 8663
rect 19646 8608 20606 8646
rect 20664 8646 20866 8663
rect 21422 8663 21438 8680
rect 21868 8680 22456 8696
rect 21868 8663 21884 8680
rect 21422 8646 21624 8663
rect 20664 8608 21624 8646
rect 21682 8646 21884 8663
rect 22440 8663 22456 8680
rect 22886 8680 23474 8696
rect 22886 8663 22902 8680
rect 22440 8646 22642 8663
rect 21682 8608 22642 8646
rect 22700 8646 22902 8663
rect 23458 8663 23474 8680
rect 23904 8680 24492 8696
rect 23904 8663 23920 8680
rect 23458 8646 23660 8663
rect 22700 8608 23660 8646
rect 23718 8646 23920 8663
rect 24476 8663 24492 8680
rect 24922 8680 25510 8696
rect 24922 8663 24938 8680
rect 24476 8646 24678 8663
rect 23718 8608 24678 8646
rect 24736 8646 24938 8663
rect 25494 8663 25510 8680
rect 25940 8680 26528 8696
rect 25940 8663 25956 8680
rect 25494 8646 25696 8663
rect 24736 8608 25696 8646
rect 25754 8646 25956 8663
rect 26512 8663 26528 8680
rect 26958 8680 27546 8696
rect 26958 8663 26974 8680
rect 26512 8646 26714 8663
rect 25754 8608 26714 8646
rect 26772 8646 26974 8663
rect 27530 8663 27546 8680
rect 27976 8680 28564 8696
rect 27976 8663 27992 8680
rect 27530 8646 27732 8663
rect 26772 8608 27732 8646
rect 27790 8646 27992 8663
rect 28548 8663 28564 8680
rect 28994 8680 29582 8696
rect 28994 8663 29010 8680
rect 28548 8646 28750 8663
rect 27790 8608 28750 8646
rect 28808 8646 29010 8663
rect 29566 8663 29582 8680
rect 30012 8680 30600 8696
rect 30012 8663 30028 8680
rect 29566 8646 29768 8663
rect 28808 8608 29768 8646
rect 29826 8646 30028 8663
rect 30584 8663 30600 8680
rect 31030 8680 31618 8696
rect 31030 8663 31046 8680
rect 30584 8646 30786 8663
rect 29826 8608 30786 8646
rect 30844 8646 31046 8663
rect 31602 8663 31618 8680
rect 32048 8680 32636 8696
rect 32048 8663 32064 8680
rect 31602 8646 31804 8663
rect 30844 8608 31804 8646
rect 31862 8646 32064 8663
rect 32620 8663 32636 8680
rect 33066 8680 33654 8696
rect 33066 8663 33082 8680
rect 32620 8646 32822 8663
rect 31862 8608 32822 8646
rect 32880 8646 33082 8663
rect 33638 8663 33654 8680
rect 33638 8646 33840 8663
rect 32880 8608 33840 8646
rect 1774 8482 2734 8520
rect 1774 8465 1976 8482
rect 1960 8448 1976 8465
rect 2532 8465 2734 8482
rect 2792 8482 3752 8520
rect 2792 8465 2994 8482
rect 2532 8448 2548 8465
rect 1960 8432 2548 8448
rect 2978 8448 2994 8465
rect 3550 8465 3752 8482
rect 3810 8482 4770 8520
rect 3810 8465 4012 8482
rect 3550 8448 3566 8465
rect 2978 8432 3566 8448
rect 1960 8374 2548 8390
rect 1960 8357 1976 8374
rect 1774 8340 1976 8357
rect 2532 8357 2548 8374
rect 3996 8448 4012 8465
rect 4568 8465 4770 8482
rect 4828 8482 5788 8520
rect 4828 8465 5030 8482
rect 4568 8448 4584 8465
rect 3996 8432 4584 8448
rect 2978 8374 3566 8390
rect 2978 8357 2994 8374
rect 2532 8340 2734 8357
rect 1774 8302 2734 8340
rect 2792 8340 2994 8357
rect 3550 8357 3566 8374
rect 5014 8448 5030 8465
rect 5586 8465 5788 8482
rect 5846 8482 6806 8520
rect 5846 8465 6048 8482
rect 5586 8448 5602 8465
rect 5014 8432 5602 8448
rect 3996 8374 4584 8390
rect 3996 8357 4012 8374
rect 3550 8340 3752 8357
rect 2792 8302 3752 8340
rect 3810 8340 4012 8357
rect 4568 8357 4584 8374
rect 6032 8448 6048 8465
rect 6604 8465 6806 8482
rect 6864 8482 7824 8520
rect 6864 8465 7066 8482
rect 6604 8448 6620 8465
rect 6032 8432 6620 8448
rect 5014 8374 5602 8390
rect 5014 8357 5030 8374
rect 4568 8340 4770 8357
rect 3810 8302 4770 8340
rect 4828 8340 5030 8357
rect 5586 8357 5602 8374
rect 7050 8448 7066 8465
rect 7622 8465 7824 8482
rect 7882 8482 8842 8520
rect 7882 8465 8084 8482
rect 7622 8448 7638 8465
rect 7050 8432 7638 8448
rect 6032 8374 6620 8390
rect 6032 8357 6048 8374
rect 5586 8340 5788 8357
rect 4828 8302 5788 8340
rect 5846 8340 6048 8357
rect 6604 8357 6620 8374
rect 8068 8448 8084 8465
rect 8640 8465 8842 8482
rect 8900 8482 9860 8520
rect 8900 8465 9102 8482
rect 8640 8448 8656 8465
rect 8068 8432 8656 8448
rect 7050 8374 7638 8390
rect 7050 8357 7066 8374
rect 6604 8340 6806 8357
rect 5846 8302 6806 8340
rect 6864 8340 7066 8357
rect 7622 8357 7638 8374
rect 9086 8448 9102 8465
rect 9658 8465 9860 8482
rect 9918 8482 10878 8520
rect 9918 8465 10120 8482
rect 9658 8448 9674 8465
rect 9086 8432 9674 8448
rect 8068 8374 8656 8390
rect 8068 8357 8084 8374
rect 7622 8340 7824 8357
rect 6864 8302 7824 8340
rect 7882 8340 8084 8357
rect 8640 8357 8656 8374
rect 10104 8448 10120 8465
rect 10676 8465 10878 8482
rect 10676 8448 10692 8465
rect 10104 8432 10692 8448
rect 9086 8374 9674 8390
rect 9086 8357 9102 8374
rect 8640 8340 8842 8357
rect 7882 8302 8842 8340
rect 8900 8340 9102 8357
rect 9658 8357 9674 8374
rect 10104 8374 10692 8390
rect 10104 8357 10120 8374
rect 9658 8340 9860 8357
rect 8900 8302 9860 8340
rect 9918 8340 10120 8357
rect 10676 8357 10692 8374
rect 10676 8340 10878 8357
rect 9918 8302 10878 8340
rect 13538 7970 14498 8008
rect 13538 7953 13740 7970
rect 13724 7936 13740 7953
rect 14296 7953 14498 7970
rect 14556 7970 15516 8008
rect 14556 7953 14758 7970
rect 14296 7936 14312 7953
rect 13724 7920 14312 7936
rect 14742 7936 14758 7953
rect 15314 7953 15516 7970
rect 15574 7970 16534 8008
rect 15574 7953 15776 7970
rect 15314 7936 15330 7953
rect 14742 7920 15330 7936
rect 15760 7936 15776 7953
rect 16332 7953 16534 7970
rect 16592 7970 17552 8008
rect 16592 7953 16794 7970
rect 16332 7936 16348 7953
rect 15760 7920 16348 7936
rect 16778 7936 16794 7953
rect 17350 7953 17552 7970
rect 17610 7970 18570 8008
rect 17610 7953 17812 7970
rect 17350 7936 17366 7953
rect 16778 7920 17366 7936
rect 17796 7936 17812 7953
rect 18368 7953 18570 7970
rect 18628 7970 19588 8008
rect 18628 7953 18830 7970
rect 18368 7936 18384 7953
rect 17796 7920 18384 7936
rect 18814 7936 18830 7953
rect 19386 7953 19588 7970
rect 19646 7970 20606 8008
rect 19646 7953 19848 7970
rect 19386 7936 19402 7953
rect 18814 7920 19402 7936
rect 19832 7936 19848 7953
rect 20404 7953 20606 7970
rect 20664 7970 21624 8008
rect 20664 7953 20866 7970
rect 20404 7936 20420 7953
rect 19832 7920 20420 7936
rect 20850 7936 20866 7953
rect 21422 7953 21624 7970
rect 21682 7970 22642 8008
rect 21682 7953 21884 7970
rect 21422 7936 21438 7953
rect 20850 7920 21438 7936
rect 21868 7936 21884 7953
rect 22440 7953 22642 7970
rect 22700 7970 23660 8008
rect 22700 7953 22902 7970
rect 22440 7936 22456 7953
rect 21868 7920 22456 7936
rect 22886 7936 22902 7953
rect 23458 7953 23660 7970
rect 23718 7970 24678 8008
rect 23718 7953 23920 7970
rect 23458 7936 23474 7953
rect 22886 7920 23474 7936
rect 23904 7936 23920 7953
rect 24476 7953 24678 7970
rect 24736 7970 25696 8008
rect 24736 7953 24938 7970
rect 24476 7936 24492 7953
rect 23904 7920 24492 7936
rect 24922 7936 24938 7953
rect 25494 7953 25696 7970
rect 25754 7970 26714 8008
rect 25754 7953 25956 7970
rect 25494 7936 25510 7953
rect 24922 7920 25510 7936
rect 25940 7936 25956 7953
rect 26512 7953 26714 7970
rect 26772 7970 27732 8008
rect 26772 7953 26974 7970
rect 26512 7936 26528 7953
rect 25940 7920 26528 7936
rect 26958 7936 26974 7953
rect 27530 7953 27732 7970
rect 27790 7970 28750 8008
rect 27790 7953 27992 7970
rect 27530 7936 27546 7953
rect 26958 7920 27546 7936
rect 27976 7936 27992 7953
rect 28548 7953 28750 7970
rect 28808 7970 29768 8008
rect 28808 7953 29010 7970
rect 28548 7936 28564 7953
rect 27976 7920 28564 7936
rect 28994 7936 29010 7953
rect 29566 7953 29768 7970
rect 29826 7970 30786 8008
rect 29826 7953 30028 7970
rect 29566 7936 29582 7953
rect 28994 7920 29582 7936
rect 30012 7936 30028 7953
rect 30584 7953 30786 7970
rect 30844 7970 31804 8008
rect 30844 7953 31046 7970
rect 30584 7936 30600 7953
rect 30012 7920 30600 7936
rect 31030 7936 31046 7953
rect 31602 7953 31804 7970
rect 31862 7970 32822 8008
rect 31862 7953 32064 7970
rect 31602 7936 31618 7953
rect 31030 7920 31618 7936
rect 32048 7936 32064 7953
rect 32620 7953 32822 7970
rect 32880 7970 33840 8008
rect 32880 7953 33082 7970
rect 32620 7936 32636 7953
rect 32048 7920 32636 7936
rect 33066 7936 33082 7953
rect 33638 7953 33840 7970
rect 33638 7936 33654 7953
rect 33066 7920 33654 7936
rect 1774 7664 2734 7702
rect 1774 7647 1976 7664
rect 1960 7630 1976 7647
rect 2532 7647 2734 7664
rect 2792 7664 3752 7702
rect 2792 7647 2994 7664
rect 2532 7630 2548 7647
rect 1960 7614 2548 7630
rect 2978 7630 2994 7647
rect 3550 7647 3752 7664
rect 3810 7664 4770 7702
rect 3810 7647 4012 7664
rect 3550 7630 3566 7647
rect 2978 7614 3566 7630
rect 3996 7630 4012 7647
rect 4568 7647 4770 7664
rect 4828 7664 5788 7702
rect 4828 7647 5030 7664
rect 4568 7630 4584 7647
rect 3996 7614 4584 7630
rect 5014 7630 5030 7647
rect 5586 7647 5788 7664
rect 5846 7664 6806 7702
rect 5846 7647 6048 7664
rect 5586 7630 5602 7647
rect 5014 7614 5602 7630
rect 6032 7630 6048 7647
rect 6604 7647 6806 7664
rect 6864 7664 7824 7702
rect 6864 7647 7066 7664
rect 6604 7630 6620 7647
rect 6032 7614 6620 7630
rect 7050 7630 7066 7647
rect 7622 7647 7824 7664
rect 7882 7664 8842 7702
rect 7882 7647 8084 7664
rect 7622 7630 7638 7647
rect 7050 7614 7638 7630
rect 8068 7630 8084 7647
rect 8640 7647 8842 7664
rect 8900 7664 9860 7702
rect 8900 7647 9102 7664
rect 8640 7630 8656 7647
rect 8068 7614 8656 7630
rect 9086 7630 9102 7647
rect 9658 7647 9860 7664
rect 9918 7664 10878 7702
rect 9918 7647 10120 7664
rect 9658 7630 9674 7647
rect 9086 7614 9674 7630
rect 10104 7630 10120 7647
rect 10676 7647 10878 7664
rect 10676 7630 10692 7647
rect 10104 7614 10692 7630
rect 13724 7448 14312 7464
rect 13724 7431 13740 7448
rect 13538 7414 13740 7431
rect 14296 7431 14312 7448
rect 14742 7448 15330 7464
rect 14742 7431 14758 7448
rect 14296 7414 14498 7431
rect 13538 7376 14498 7414
rect 14556 7414 14758 7431
rect 15314 7431 15330 7448
rect 15760 7448 16348 7464
rect 15760 7431 15776 7448
rect 15314 7414 15516 7431
rect 14556 7376 15516 7414
rect 15574 7414 15776 7431
rect 16332 7431 16348 7448
rect 16778 7448 17366 7464
rect 16778 7431 16794 7448
rect 16332 7414 16534 7431
rect 15574 7376 16534 7414
rect 16592 7414 16794 7431
rect 17350 7431 17366 7448
rect 17796 7448 18384 7464
rect 17796 7431 17812 7448
rect 17350 7414 17552 7431
rect 16592 7376 17552 7414
rect 17610 7414 17812 7431
rect 18368 7431 18384 7448
rect 18814 7448 19402 7464
rect 18814 7431 18830 7448
rect 18368 7414 18570 7431
rect 17610 7376 18570 7414
rect 18628 7414 18830 7431
rect 19386 7431 19402 7448
rect 19832 7448 20420 7464
rect 19832 7431 19848 7448
rect 19386 7414 19588 7431
rect 18628 7376 19588 7414
rect 19646 7414 19848 7431
rect 20404 7431 20420 7448
rect 20850 7448 21438 7464
rect 20850 7431 20866 7448
rect 20404 7414 20606 7431
rect 19646 7376 20606 7414
rect 20664 7414 20866 7431
rect 21422 7431 21438 7448
rect 21868 7448 22456 7464
rect 21868 7431 21884 7448
rect 21422 7414 21624 7431
rect 20664 7376 21624 7414
rect 21682 7414 21884 7431
rect 22440 7431 22456 7448
rect 22886 7448 23474 7464
rect 22886 7431 22902 7448
rect 22440 7414 22642 7431
rect 21682 7376 22642 7414
rect 22700 7414 22902 7431
rect 23458 7431 23474 7448
rect 23904 7448 24492 7464
rect 23904 7431 23920 7448
rect 23458 7414 23660 7431
rect 22700 7376 23660 7414
rect 23718 7414 23920 7431
rect 24476 7431 24492 7448
rect 24922 7448 25510 7464
rect 24922 7431 24938 7448
rect 24476 7414 24678 7431
rect 23718 7376 24678 7414
rect 24736 7414 24938 7431
rect 25494 7431 25510 7448
rect 25940 7448 26528 7464
rect 25940 7431 25956 7448
rect 25494 7414 25696 7431
rect 24736 7376 25696 7414
rect 25754 7414 25956 7431
rect 26512 7431 26528 7448
rect 26958 7448 27546 7464
rect 26958 7431 26974 7448
rect 26512 7414 26714 7431
rect 25754 7376 26714 7414
rect 26772 7414 26974 7431
rect 27530 7431 27546 7448
rect 27976 7448 28564 7464
rect 27976 7431 27992 7448
rect 27530 7414 27732 7431
rect 26772 7376 27732 7414
rect 27790 7414 27992 7431
rect 28548 7431 28564 7448
rect 28994 7448 29582 7464
rect 28994 7431 29010 7448
rect 28548 7414 28750 7431
rect 27790 7376 28750 7414
rect 28808 7414 29010 7431
rect 29566 7431 29582 7448
rect 30012 7448 30600 7464
rect 30012 7431 30028 7448
rect 29566 7414 29768 7431
rect 28808 7376 29768 7414
rect 29826 7414 30028 7431
rect 30584 7431 30600 7448
rect 31030 7448 31618 7464
rect 31030 7431 31046 7448
rect 30584 7414 30786 7431
rect 29826 7376 30786 7414
rect 30844 7414 31046 7431
rect 31602 7431 31618 7448
rect 32048 7448 32636 7464
rect 32048 7431 32064 7448
rect 31602 7414 31804 7431
rect 30844 7376 31804 7414
rect 31862 7414 32064 7431
rect 32620 7431 32636 7448
rect 33066 7448 33654 7464
rect 33066 7431 33082 7448
rect 32620 7414 32822 7431
rect 31862 7376 32822 7414
rect 32880 7414 33082 7431
rect 33638 7431 33654 7448
rect 33638 7414 33840 7431
rect 32880 7376 33840 7414
rect 13538 6738 14498 6776
rect 13538 6721 13740 6738
rect 13724 6704 13740 6721
rect 14296 6721 14498 6738
rect 14556 6738 15516 6776
rect 14556 6721 14758 6738
rect 14296 6704 14312 6721
rect 13724 6688 14312 6704
rect 14742 6704 14758 6721
rect 15314 6721 15516 6738
rect 15574 6738 16534 6776
rect 15574 6721 15776 6738
rect 15314 6704 15330 6721
rect 14742 6688 15330 6704
rect 15760 6704 15776 6721
rect 16332 6721 16534 6738
rect 16592 6738 17552 6776
rect 16592 6721 16794 6738
rect 16332 6704 16348 6721
rect 15760 6688 16348 6704
rect 16778 6704 16794 6721
rect 17350 6721 17552 6738
rect 17610 6738 18570 6776
rect 17610 6721 17812 6738
rect 17350 6704 17366 6721
rect 16778 6688 17366 6704
rect 17796 6704 17812 6721
rect 18368 6721 18570 6738
rect 18628 6738 19588 6776
rect 18628 6721 18830 6738
rect 18368 6704 18384 6721
rect 17796 6688 18384 6704
rect 18814 6704 18830 6721
rect 19386 6721 19588 6738
rect 19646 6738 20606 6776
rect 19646 6721 19848 6738
rect 19386 6704 19402 6721
rect 18814 6688 19402 6704
rect 19832 6704 19848 6721
rect 20404 6721 20606 6738
rect 20664 6738 21624 6776
rect 20664 6721 20866 6738
rect 20404 6704 20420 6721
rect 19832 6688 20420 6704
rect 20850 6704 20866 6721
rect 21422 6721 21624 6738
rect 21682 6738 22642 6776
rect 21682 6721 21884 6738
rect 21422 6704 21438 6721
rect 20850 6688 21438 6704
rect 21868 6704 21884 6721
rect 22440 6721 22642 6738
rect 22700 6738 23660 6776
rect 22700 6721 22902 6738
rect 22440 6704 22456 6721
rect 21868 6688 22456 6704
rect 22886 6704 22902 6721
rect 23458 6721 23660 6738
rect 23718 6738 24678 6776
rect 23718 6721 23920 6738
rect 23458 6704 23474 6721
rect 22886 6688 23474 6704
rect 23904 6704 23920 6721
rect 24476 6721 24678 6738
rect 24736 6738 25696 6776
rect 24736 6721 24938 6738
rect 24476 6704 24492 6721
rect 23904 6688 24492 6704
rect 24922 6704 24938 6721
rect 25494 6721 25696 6738
rect 25754 6738 26714 6776
rect 25754 6721 25956 6738
rect 25494 6704 25510 6721
rect 24922 6688 25510 6704
rect 25940 6704 25956 6721
rect 26512 6721 26714 6738
rect 26772 6738 27732 6776
rect 26772 6721 26974 6738
rect 26512 6704 26528 6721
rect 25940 6688 26528 6704
rect 26958 6704 26974 6721
rect 27530 6721 27732 6738
rect 27790 6738 28750 6776
rect 27790 6721 27992 6738
rect 27530 6704 27546 6721
rect 26958 6688 27546 6704
rect 27976 6704 27992 6721
rect 28548 6721 28750 6738
rect 28808 6738 29768 6776
rect 28808 6721 29010 6738
rect 28548 6704 28564 6721
rect 27976 6688 28564 6704
rect 28994 6704 29010 6721
rect 29566 6721 29768 6738
rect 29826 6738 30786 6776
rect 29826 6721 30028 6738
rect 29566 6704 29582 6721
rect 28994 6688 29582 6704
rect 30012 6704 30028 6721
rect 30584 6721 30786 6738
rect 30844 6738 31804 6776
rect 30844 6721 31046 6738
rect 30584 6704 30600 6721
rect 30012 6688 30600 6704
rect 31030 6704 31046 6721
rect 31602 6721 31804 6738
rect 31862 6738 32822 6776
rect 31862 6721 32064 6738
rect 31602 6704 31618 6721
rect 31030 6688 31618 6704
rect 32048 6704 32064 6721
rect 32620 6721 32822 6738
rect 32880 6738 33840 6776
rect 32880 6721 33082 6738
rect 32620 6704 32636 6721
rect 32048 6688 32636 6704
rect 33066 6704 33082 6721
rect 33638 6721 33840 6738
rect 33638 6704 33654 6721
rect 33066 6688 33654 6704
rect 636 6350 1224 6366
rect 636 6333 652 6350
rect 450 6316 652 6333
rect 1208 6333 1224 6350
rect 1654 6350 2242 6366
rect 1654 6333 1670 6350
rect 1208 6316 1410 6333
rect 450 6278 1410 6316
rect 1468 6316 1670 6333
rect 2226 6333 2242 6350
rect 2672 6350 3260 6366
rect 2672 6333 2688 6350
rect 2226 6316 2428 6333
rect 1468 6278 2428 6316
rect 2486 6316 2688 6333
rect 3244 6333 3260 6350
rect 3690 6350 4278 6366
rect 3690 6333 3706 6350
rect 3244 6316 3446 6333
rect 2486 6278 3446 6316
rect 3504 6316 3706 6333
rect 4262 6333 4278 6350
rect 4708 6350 5296 6366
rect 4708 6333 4724 6350
rect 4262 6316 4464 6333
rect 3504 6278 4464 6316
rect 4522 6316 4724 6333
rect 5280 6333 5296 6350
rect 5726 6350 6314 6366
rect 5726 6333 5742 6350
rect 5280 6316 5482 6333
rect 4522 6278 5482 6316
rect 5540 6316 5742 6333
rect 6298 6333 6314 6350
rect 6744 6350 7332 6366
rect 6744 6333 6760 6350
rect 6298 6316 6500 6333
rect 5540 6278 6500 6316
rect 6558 6316 6760 6333
rect 7316 6333 7332 6350
rect 7762 6350 8350 6366
rect 7762 6333 7778 6350
rect 7316 6316 7518 6333
rect 6558 6278 7518 6316
rect 7576 6316 7778 6333
rect 8334 6333 8350 6350
rect 8780 6350 9368 6366
rect 8780 6333 8796 6350
rect 8334 6316 8536 6333
rect 7576 6278 8536 6316
rect 8594 6316 8796 6333
rect 9352 6333 9368 6350
rect 9798 6350 10386 6366
rect 9798 6333 9814 6350
rect 9352 6316 9554 6333
rect 8594 6278 9554 6316
rect 9612 6316 9814 6333
rect 10370 6333 10386 6350
rect 10816 6350 11404 6366
rect 10816 6333 10832 6350
rect 10370 6316 10572 6333
rect 9612 6278 10572 6316
rect 10630 6316 10832 6333
rect 11388 6333 11404 6350
rect 11388 6316 11590 6333
rect 10630 6278 11590 6316
rect 13724 6214 14312 6230
rect 13724 6197 13740 6214
rect 13538 6180 13740 6197
rect 14296 6197 14312 6214
rect 14742 6214 15330 6230
rect 14742 6197 14758 6214
rect 14296 6180 14498 6197
rect 13538 6142 14498 6180
rect 14556 6180 14758 6197
rect 15314 6197 15330 6214
rect 15760 6214 16348 6230
rect 15760 6197 15776 6214
rect 15314 6180 15516 6197
rect 14556 6142 15516 6180
rect 15574 6180 15776 6197
rect 16332 6197 16348 6214
rect 16778 6214 17366 6230
rect 16778 6197 16794 6214
rect 16332 6180 16534 6197
rect 15574 6142 16534 6180
rect 16592 6180 16794 6197
rect 17350 6197 17366 6214
rect 17796 6214 18384 6230
rect 17796 6197 17812 6214
rect 17350 6180 17552 6197
rect 16592 6142 17552 6180
rect 17610 6180 17812 6197
rect 18368 6197 18384 6214
rect 18814 6214 19402 6230
rect 18814 6197 18830 6214
rect 18368 6180 18570 6197
rect 17610 6142 18570 6180
rect 18628 6180 18830 6197
rect 19386 6197 19402 6214
rect 19832 6214 20420 6230
rect 19832 6197 19848 6214
rect 19386 6180 19588 6197
rect 18628 6142 19588 6180
rect 19646 6180 19848 6197
rect 20404 6197 20420 6214
rect 20850 6214 21438 6230
rect 20850 6197 20866 6214
rect 20404 6180 20606 6197
rect 19646 6142 20606 6180
rect 20664 6180 20866 6197
rect 21422 6197 21438 6214
rect 21868 6214 22456 6230
rect 21868 6197 21884 6214
rect 21422 6180 21624 6197
rect 20664 6142 21624 6180
rect 21682 6180 21884 6197
rect 22440 6197 22456 6214
rect 22886 6214 23474 6230
rect 22886 6197 22902 6214
rect 22440 6180 22642 6197
rect 21682 6142 22642 6180
rect 22700 6180 22902 6197
rect 23458 6197 23474 6214
rect 23904 6214 24492 6230
rect 23904 6197 23920 6214
rect 23458 6180 23660 6197
rect 22700 6142 23660 6180
rect 23718 6180 23920 6197
rect 24476 6197 24492 6214
rect 24922 6214 25510 6230
rect 24922 6197 24938 6214
rect 24476 6180 24678 6197
rect 23718 6142 24678 6180
rect 24736 6180 24938 6197
rect 25494 6197 25510 6214
rect 25940 6214 26528 6230
rect 25940 6197 25956 6214
rect 25494 6180 25696 6197
rect 24736 6142 25696 6180
rect 25754 6180 25956 6197
rect 26512 6197 26528 6214
rect 26958 6214 27546 6230
rect 26958 6197 26974 6214
rect 26512 6180 26714 6197
rect 25754 6142 26714 6180
rect 26772 6180 26974 6197
rect 27530 6197 27546 6214
rect 27976 6214 28564 6230
rect 27976 6197 27992 6214
rect 27530 6180 27732 6197
rect 26772 6142 27732 6180
rect 27790 6180 27992 6197
rect 28548 6197 28564 6214
rect 28994 6214 29582 6230
rect 28994 6197 29010 6214
rect 28548 6180 28750 6197
rect 27790 6142 28750 6180
rect 28808 6180 29010 6197
rect 29566 6197 29582 6214
rect 30012 6214 30600 6230
rect 30012 6197 30028 6214
rect 29566 6180 29768 6197
rect 28808 6142 29768 6180
rect 29826 6180 30028 6197
rect 30584 6197 30600 6214
rect 31030 6214 31618 6230
rect 31030 6197 31046 6214
rect 30584 6180 30786 6197
rect 29826 6142 30786 6180
rect 30844 6180 31046 6197
rect 31602 6197 31618 6214
rect 32048 6214 32636 6230
rect 32048 6197 32064 6214
rect 31602 6180 31804 6197
rect 30844 6142 31804 6180
rect 31862 6180 32064 6197
rect 32620 6197 32636 6214
rect 33066 6214 33654 6230
rect 33066 6197 33082 6214
rect 32620 6180 32822 6197
rect 31862 6142 32822 6180
rect 32880 6180 33082 6197
rect 33638 6197 33654 6214
rect 33638 6180 33840 6197
rect 32880 6142 33840 6180
rect 450 5640 1410 5678
rect 450 5623 652 5640
rect 636 5606 652 5623
rect 1208 5623 1410 5640
rect 1468 5640 2428 5678
rect 1468 5623 1670 5640
rect 1208 5606 1224 5623
rect 636 5590 1224 5606
rect 1654 5606 1670 5623
rect 2226 5623 2428 5640
rect 2486 5640 3446 5678
rect 2486 5623 2688 5640
rect 2226 5606 2242 5623
rect 1654 5590 2242 5606
rect 2672 5606 2688 5623
rect 3244 5623 3446 5640
rect 3504 5640 4464 5678
rect 3504 5623 3706 5640
rect 3244 5606 3260 5623
rect 2672 5590 3260 5606
rect 3690 5606 3706 5623
rect 4262 5623 4464 5640
rect 4522 5640 5482 5678
rect 4522 5623 4724 5640
rect 4262 5606 4278 5623
rect 3690 5590 4278 5606
rect 4708 5606 4724 5623
rect 5280 5623 5482 5640
rect 5540 5640 6500 5678
rect 5540 5623 5742 5640
rect 5280 5606 5296 5623
rect 4708 5590 5296 5606
rect 5726 5606 5742 5623
rect 6298 5623 6500 5640
rect 6558 5640 7518 5678
rect 6558 5623 6760 5640
rect 6298 5606 6314 5623
rect 5726 5590 6314 5606
rect 6744 5606 6760 5623
rect 7316 5623 7518 5640
rect 7576 5640 8536 5678
rect 7576 5623 7778 5640
rect 7316 5606 7332 5623
rect 6744 5590 7332 5606
rect 7762 5606 7778 5623
rect 8334 5623 8536 5640
rect 8594 5640 9554 5678
rect 8594 5623 8796 5640
rect 8334 5606 8350 5623
rect 7762 5590 8350 5606
rect 8780 5606 8796 5623
rect 9352 5623 9554 5640
rect 9612 5640 10572 5678
rect 9612 5623 9814 5640
rect 9352 5606 9368 5623
rect 8780 5590 9368 5606
rect 9798 5606 9814 5623
rect 10370 5623 10572 5640
rect 10630 5640 11590 5678
rect 10630 5623 10832 5640
rect 10370 5606 10386 5623
rect 9798 5590 10386 5606
rect 10816 5606 10832 5623
rect 11388 5623 11590 5640
rect 11388 5606 11404 5623
rect 10816 5590 11404 5606
rect 13538 5504 14498 5542
rect 13538 5487 13740 5504
rect 13724 5470 13740 5487
rect 14296 5487 14498 5504
rect 14556 5504 15516 5542
rect 14556 5487 14758 5504
rect 14296 5470 14312 5487
rect 13724 5454 14312 5470
rect 14742 5470 14758 5487
rect 15314 5487 15516 5504
rect 15574 5504 16534 5542
rect 15574 5487 15776 5504
rect 15314 5470 15330 5487
rect 14742 5454 15330 5470
rect 15760 5470 15776 5487
rect 16332 5487 16534 5504
rect 16592 5504 17552 5542
rect 16592 5487 16794 5504
rect 16332 5470 16348 5487
rect 15760 5454 16348 5470
rect 16778 5470 16794 5487
rect 17350 5487 17552 5504
rect 17610 5504 18570 5542
rect 17610 5487 17812 5504
rect 17350 5470 17366 5487
rect 16778 5454 17366 5470
rect 17796 5470 17812 5487
rect 18368 5487 18570 5504
rect 18628 5504 19588 5542
rect 18628 5487 18830 5504
rect 18368 5470 18384 5487
rect 17796 5454 18384 5470
rect 18814 5470 18830 5487
rect 19386 5487 19588 5504
rect 19646 5504 20606 5542
rect 19646 5487 19848 5504
rect 19386 5470 19402 5487
rect 18814 5454 19402 5470
rect 19832 5470 19848 5487
rect 20404 5487 20606 5504
rect 20664 5504 21624 5542
rect 20664 5487 20866 5504
rect 20404 5470 20420 5487
rect 19832 5454 20420 5470
rect 20850 5470 20866 5487
rect 21422 5487 21624 5504
rect 21682 5504 22642 5542
rect 21682 5487 21884 5504
rect 21422 5470 21438 5487
rect 20850 5454 21438 5470
rect 21868 5470 21884 5487
rect 22440 5487 22642 5504
rect 22700 5504 23660 5542
rect 22700 5487 22902 5504
rect 22440 5470 22456 5487
rect 21868 5454 22456 5470
rect 22886 5470 22902 5487
rect 23458 5487 23660 5504
rect 23718 5504 24678 5542
rect 23718 5487 23920 5504
rect 23458 5470 23474 5487
rect 22886 5454 23474 5470
rect 23904 5470 23920 5487
rect 24476 5487 24678 5504
rect 24736 5504 25696 5542
rect 24736 5487 24938 5504
rect 24476 5470 24492 5487
rect 23904 5454 24492 5470
rect 24922 5470 24938 5487
rect 25494 5487 25696 5504
rect 25754 5504 26714 5542
rect 25754 5487 25956 5504
rect 25494 5470 25510 5487
rect 24922 5454 25510 5470
rect 25940 5470 25956 5487
rect 26512 5487 26714 5504
rect 26772 5504 27732 5542
rect 26772 5487 26974 5504
rect 26512 5470 26528 5487
rect 25940 5454 26528 5470
rect 26958 5470 26974 5487
rect 27530 5487 27732 5504
rect 27790 5504 28750 5542
rect 27790 5487 27992 5504
rect 27530 5470 27546 5487
rect 26958 5454 27546 5470
rect 27976 5470 27992 5487
rect 28548 5487 28750 5504
rect 28808 5504 29768 5542
rect 28808 5487 29010 5504
rect 28548 5470 28564 5487
rect 27976 5454 28564 5470
rect 28994 5470 29010 5487
rect 29566 5487 29768 5504
rect 29826 5504 30786 5542
rect 29826 5487 30028 5504
rect 29566 5470 29582 5487
rect 28994 5454 29582 5470
rect 30012 5470 30028 5487
rect 30584 5487 30786 5504
rect 30844 5504 31804 5542
rect 30844 5487 31046 5504
rect 30584 5470 30600 5487
rect 30012 5454 30600 5470
rect 31030 5470 31046 5487
rect 31602 5487 31804 5504
rect 31862 5504 32822 5542
rect 31862 5487 32064 5504
rect 31602 5470 31618 5487
rect 31030 5454 31618 5470
rect 32048 5470 32064 5487
rect 32620 5487 32822 5504
rect 32880 5504 33840 5542
rect 32880 5487 33082 5504
rect 32620 5470 32636 5487
rect 32048 5454 32636 5470
rect 33066 5470 33082 5487
rect 33638 5487 33840 5504
rect 33638 5470 33654 5487
rect 33066 5454 33654 5470
rect 636 5238 1224 5254
rect 636 5221 652 5238
rect 450 5204 652 5221
rect 1208 5221 1224 5238
rect 1654 5238 2242 5254
rect 1654 5221 1670 5238
rect 1208 5204 1410 5221
rect 450 5166 1410 5204
rect 1468 5204 1670 5221
rect 2226 5221 2242 5238
rect 2672 5238 3260 5254
rect 2672 5221 2688 5238
rect 2226 5204 2428 5221
rect 1468 5166 2428 5204
rect 2486 5204 2688 5221
rect 3244 5221 3260 5238
rect 3690 5238 4278 5254
rect 3690 5221 3706 5238
rect 3244 5204 3446 5221
rect 2486 5166 3446 5204
rect 3504 5204 3706 5221
rect 4262 5221 4278 5238
rect 4708 5238 5296 5254
rect 4708 5221 4724 5238
rect 4262 5204 4464 5221
rect 3504 5166 4464 5204
rect 4522 5204 4724 5221
rect 5280 5221 5296 5238
rect 5726 5238 6314 5254
rect 5726 5221 5742 5238
rect 5280 5204 5482 5221
rect 4522 5166 5482 5204
rect 5540 5204 5742 5221
rect 6298 5221 6314 5238
rect 6744 5238 7332 5254
rect 6744 5221 6760 5238
rect 6298 5204 6500 5221
rect 5540 5166 6500 5204
rect 6558 5204 6760 5221
rect 7316 5221 7332 5238
rect 7762 5238 8350 5254
rect 7762 5221 7778 5238
rect 7316 5204 7518 5221
rect 6558 5166 7518 5204
rect 7576 5204 7778 5221
rect 8334 5221 8350 5238
rect 8780 5238 9368 5254
rect 8780 5221 8796 5238
rect 8334 5204 8536 5221
rect 7576 5166 8536 5204
rect 8594 5204 8796 5221
rect 9352 5221 9368 5238
rect 9798 5238 10386 5254
rect 9798 5221 9814 5238
rect 9352 5204 9554 5221
rect 8594 5166 9554 5204
rect 9612 5204 9814 5221
rect 10370 5221 10386 5238
rect 10816 5238 11404 5254
rect 10816 5221 10832 5238
rect 10370 5204 10572 5221
rect 9612 5166 10572 5204
rect 10630 5204 10832 5221
rect 11388 5221 11404 5238
rect 11388 5204 11590 5221
rect 10630 5166 11590 5204
rect 13724 4980 14312 4996
rect 13724 4963 13740 4980
rect 13538 4946 13740 4963
rect 14296 4963 14312 4980
rect 14742 4980 15330 4996
rect 14742 4963 14758 4980
rect 14296 4946 14498 4963
rect 13538 4908 14498 4946
rect 14556 4946 14758 4963
rect 15314 4963 15330 4980
rect 15760 4980 16348 4996
rect 15760 4963 15776 4980
rect 15314 4946 15516 4963
rect 14556 4908 15516 4946
rect 15574 4946 15776 4963
rect 16332 4963 16348 4980
rect 16778 4980 17366 4996
rect 16778 4963 16794 4980
rect 16332 4946 16534 4963
rect 15574 4908 16534 4946
rect 16592 4946 16794 4963
rect 17350 4963 17366 4980
rect 17796 4980 18384 4996
rect 17796 4963 17812 4980
rect 17350 4946 17552 4963
rect 16592 4908 17552 4946
rect 17610 4946 17812 4963
rect 18368 4963 18384 4980
rect 18814 4980 19402 4996
rect 18814 4963 18830 4980
rect 18368 4946 18570 4963
rect 17610 4908 18570 4946
rect 18628 4946 18830 4963
rect 19386 4963 19402 4980
rect 19832 4980 20420 4996
rect 19832 4963 19848 4980
rect 19386 4946 19588 4963
rect 18628 4908 19588 4946
rect 19646 4946 19848 4963
rect 20404 4963 20420 4980
rect 20850 4980 21438 4996
rect 20850 4963 20866 4980
rect 20404 4946 20606 4963
rect 19646 4908 20606 4946
rect 20664 4946 20866 4963
rect 21422 4963 21438 4980
rect 21868 4980 22456 4996
rect 21868 4963 21884 4980
rect 21422 4946 21624 4963
rect 20664 4908 21624 4946
rect 21682 4946 21884 4963
rect 22440 4963 22456 4980
rect 22886 4980 23474 4996
rect 22886 4963 22902 4980
rect 22440 4946 22642 4963
rect 21682 4908 22642 4946
rect 22700 4946 22902 4963
rect 23458 4963 23474 4980
rect 23904 4980 24492 4996
rect 23904 4963 23920 4980
rect 23458 4946 23660 4963
rect 22700 4908 23660 4946
rect 23718 4946 23920 4963
rect 24476 4963 24492 4980
rect 24922 4980 25510 4996
rect 24922 4963 24938 4980
rect 24476 4946 24678 4963
rect 23718 4908 24678 4946
rect 24736 4946 24938 4963
rect 25494 4963 25510 4980
rect 25940 4980 26528 4996
rect 25940 4963 25956 4980
rect 25494 4946 25696 4963
rect 24736 4908 25696 4946
rect 25754 4946 25956 4963
rect 26512 4963 26528 4980
rect 26958 4980 27546 4996
rect 26958 4963 26974 4980
rect 26512 4946 26714 4963
rect 25754 4908 26714 4946
rect 26772 4946 26974 4963
rect 27530 4963 27546 4980
rect 27976 4980 28564 4996
rect 27976 4963 27992 4980
rect 27530 4946 27732 4963
rect 26772 4908 27732 4946
rect 27790 4946 27992 4963
rect 28548 4963 28564 4980
rect 28994 4980 29582 4996
rect 28994 4963 29010 4980
rect 28548 4946 28750 4963
rect 27790 4908 28750 4946
rect 28808 4946 29010 4963
rect 29566 4963 29582 4980
rect 30012 4980 30600 4996
rect 30012 4963 30028 4980
rect 29566 4946 29768 4963
rect 28808 4908 29768 4946
rect 29826 4946 30028 4963
rect 30584 4963 30600 4980
rect 31030 4980 31618 4996
rect 31030 4963 31046 4980
rect 30584 4946 30786 4963
rect 29826 4908 30786 4946
rect 30844 4946 31046 4963
rect 31602 4963 31618 4980
rect 32048 4980 32636 4996
rect 32048 4963 32064 4980
rect 31602 4946 31804 4963
rect 30844 4908 31804 4946
rect 31862 4946 32064 4963
rect 32620 4963 32636 4980
rect 33066 4980 33654 4996
rect 33066 4963 33082 4980
rect 32620 4946 32822 4963
rect 31862 4908 32822 4946
rect 32880 4946 33082 4963
rect 33638 4963 33654 4980
rect 33638 4946 33840 4963
rect 32880 4908 33840 4946
rect 450 4528 1410 4566
rect 450 4511 652 4528
rect 636 4494 652 4511
rect 1208 4511 1410 4528
rect 1468 4528 2428 4566
rect 1468 4511 1670 4528
rect 1208 4494 1224 4511
rect 636 4478 1224 4494
rect 1654 4494 1670 4511
rect 2226 4511 2428 4528
rect 2486 4528 3446 4566
rect 2486 4511 2688 4528
rect 2226 4494 2242 4511
rect 1654 4478 2242 4494
rect 2672 4494 2688 4511
rect 3244 4511 3446 4528
rect 3504 4528 4464 4566
rect 3504 4511 3706 4528
rect 3244 4494 3260 4511
rect 2672 4478 3260 4494
rect 3690 4494 3706 4511
rect 4262 4511 4464 4528
rect 4522 4528 5482 4566
rect 4522 4511 4724 4528
rect 4262 4494 4278 4511
rect 3690 4478 4278 4494
rect 4708 4494 4724 4511
rect 5280 4511 5482 4528
rect 5540 4528 6500 4566
rect 5540 4511 5742 4528
rect 5280 4494 5296 4511
rect 4708 4478 5296 4494
rect 5726 4494 5742 4511
rect 6298 4511 6500 4528
rect 6558 4528 7518 4566
rect 6558 4511 6760 4528
rect 6298 4494 6314 4511
rect 5726 4478 6314 4494
rect 6744 4494 6760 4511
rect 7316 4511 7518 4528
rect 7576 4528 8536 4566
rect 7576 4511 7778 4528
rect 7316 4494 7332 4511
rect 6744 4478 7332 4494
rect 7762 4494 7778 4511
rect 8334 4511 8536 4528
rect 8594 4528 9554 4566
rect 8594 4511 8796 4528
rect 8334 4494 8350 4511
rect 7762 4478 8350 4494
rect 8780 4494 8796 4511
rect 9352 4511 9554 4528
rect 9612 4528 10572 4566
rect 9612 4511 9814 4528
rect 9352 4494 9368 4511
rect 8780 4478 9368 4494
rect 9798 4494 9814 4511
rect 10370 4511 10572 4528
rect 10630 4528 11590 4566
rect 10630 4511 10832 4528
rect 10370 4494 10386 4511
rect 9798 4478 10386 4494
rect 10816 4494 10832 4511
rect 11388 4511 11590 4528
rect 11388 4494 11404 4511
rect 10816 4478 11404 4494
rect 13538 4270 14498 4308
rect 13538 4253 13740 4270
rect 13724 4236 13740 4253
rect 14296 4253 14498 4270
rect 14556 4270 15516 4308
rect 14556 4253 14758 4270
rect 14296 4236 14312 4253
rect 13724 4220 14312 4236
rect 14742 4236 14758 4253
rect 15314 4253 15516 4270
rect 15574 4270 16534 4308
rect 15574 4253 15776 4270
rect 15314 4236 15330 4253
rect 14742 4220 15330 4236
rect 15760 4236 15776 4253
rect 16332 4253 16534 4270
rect 16592 4270 17552 4308
rect 16592 4253 16794 4270
rect 16332 4236 16348 4253
rect 15760 4220 16348 4236
rect 16778 4236 16794 4253
rect 17350 4253 17552 4270
rect 17610 4270 18570 4308
rect 17610 4253 17812 4270
rect 17350 4236 17366 4253
rect 16778 4220 17366 4236
rect 17796 4236 17812 4253
rect 18368 4253 18570 4270
rect 18628 4270 19588 4308
rect 18628 4253 18830 4270
rect 18368 4236 18384 4253
rect 17796 4220 18384 4236
rect 18814 4236 18830 4253
rect 19386 4253 19588 4270
rect 19646 4270 20606 4308
rect 19646 4253 19848 4270
rect 19386 4236 19402 4253
rect 18814 4220 19402 4236
rect 19832 4236 19848 4253
rect 20404 4253 20606 4270
rect 20664 4270 21624 4308
rect 20664 4253 20866 4270
rect 20404 4236 20420 4253
rect 19832 4220 20420 4236
rect 20850 4236 20866 4253
rect 21422 4253 21624 4270
rect 21682 4270 22642 4308
rect 21682 4253 21884 4270
rect 21422 4236 21438 4253
rect 20850 4220 21438 4236
rect 21868 4236 21884 4253
rect 22440 4253 22642 4270
rect 22700 4270 23660 4308
rect 22700 4253 22902 4270
rect 22440 4236 22456 4253
rect 21868 4220 22456 4236
rect 22886 4236 22902 4253
rect 23458 4253 23660 4270
rect 23718 4270 24678 4308
rect 23718 4253 23920 4270
rect 23458 4236 23474 4253
rect 22886 4220 23474 4236
rect 23904 4236 23920 4253
rect 24476 4253 24678 4270
rect 24736 4270 25696 4308
rect 24736 4253 24938 4270
rect 24476 4236 24492 4253
rect 23904 4220 24492 4236
rect 24922 4236 24938 4253
rect 25494 4253 25696 4270
rect 25754 4270 26714 4308
rect 25754 4253 25956 4270
rect 25494 4236 25510 4253
rect 24922 4220 25510 4236
rect 25940 4236 25956 4253
rect 26512 4253 26714 4270
rect 26772 4270 27732 4308
rect 26772 4253 26974 4270
rect 26512 4236 26528 4253
rect 25940 4220 26528 4236
rect 26958 4236 26974 4253
rect 27530 4253 27732 4270
rect 27790 4270 28750 4308
rect 27790 4253 27992 4270
rect 27530 4236 27546 4253
rect 26958 4220 27546 4236
rect 27976 4236 27992 4253
rect 28548 4253 28750 4270
rect 28808 4270 29768 4308
rect 28808 4253 29010 4270
rect 28548 4236 28564 4253
rect 27976 4220 28564 4236
rect 28994 4236 29010 4253
rect 29566 4253 29768 4270
rect 29826 4270 30786 4308
rect 29826 4253 30028 4270
rect 29566 4236 29582 4253
rect 28994 4220 29582 4236
rect 30012 4236 30028 4253
rect 30584 4253 30786 4270
rect 30844 4270 31804 4308
rect 30844 4253 31046 4270
rect 30584 4236 30600 4253
rect 30012 4220 30600 4236
rect 31030 4236 31046 4253
rect 31602 4253 31804 4270
rect 31862 4270 32822 4308
rect 31862 4253 32064 4270
rect 31602 4236 31618 4253
rect 31030 4220 31618 4236
rect 32048 4236 32064 4253
rect 32620 4253 32822 4270
rect 32880 4270 33840 4308
rect 32880 4253 33082 4270
rect 32620 4236 32636 4253
rect 32048 4220 32636 4236
rect 33066 4236 33082 4253
rect 33638 4253 33840 4270
rect 33638 4236 33654 4253
rect 33066 4220 33654 4236
rect 636 4126 1224 4142
rect 636 4109 652 4126
rect 450 4092 652 4109
rect 1208 4109 1224 4126
rect 1654 4126 2242 4142
rect 1654 4109 1670 4126
rect 1208 4092 1410 4109
rect 450 4054 1410 4092
rect 1468 4092 1670 4109
rect 2226 4109 2242 4126
rect 2672 4126 3260 4142
rect 2672 4109 2688 4126
rect 2226 4092 2428 4109
rect 1468 4054 2428 4092
rect 2486 4092 2688 4109
rect 3244 4109 3260 4126
rect 3690 4126 4278 4142
rect 3690 4109 3706 4126
rect 3244 4092 3446 4109
rect 2486 4054 3446 4092
rect 3504 4092 3706 4109
rect 4262 4109 4278 4126
rect 4708 4126 5296 4142
rect 4708 4109 4724 4126
rect 4262 4092 4464 4109
rect 3504 4054 4464 4092
rect 4522 4092 4724 4109
rect 5280 4109 5296 4126
rect 5726 4126 6314 4142
rect 5726 4109 5742 4126
rect 5280 4092 5482 4109
rect 4522 4054 5482 4092
rect 5540 4092 5742 4109
rect 6298 4109 6314 4126
rect 6744 4126 7332 4142
rect 6744 4109 6760 4126
rect 6298 4092 6500 4109
rect 5540 4054 6500 4092
rect 6558 4092 6760 4109
rect 7316 4109 7332 4126
rect 7762 4126 8350 4142
rect 7762 4109 7778 4126
rect 7316 4092 7518 4109
rect 6558 4054 7518 4092
rect 7576 4092 7778 4109
rect 8334 4109 8350 4126
rect 8780 4126 9368 4142
rect 8780 4109 8796 4126
rect 8334 4092 8536 4109
rect 7576 4054 8536 4092
rect 8594 4092 8796 4109
rect 9352 4109 9368 4126
rect 9798 4126 10386 4142
rect 9798 4109 9814 4126
rect 9352 4092 9554 4109
rect 8594 4054 9554 4092
rect 9612 4092 9814 4109
rect 10370 4109 10386 4126
rect 10816 4126 11404 4142
rect 10816 4109 10832 4126
rect 10370 4092 10572 4109
rect 9612 4054 10572 4092
rect 10630 4092 10832 4109
rect 11388 4109 11404 4126
rect 11388 4092 11590 4109
rect 10630 4054 11590 4092
rect 13724 3748 14312 3764
rect 13724 3731 13740 3748
rect 13538 3714 13740 3731
rect 14296 3731 14312 3748
rect 14742 3748 15330 3764
rect 14742 3731 14758 3748
rect 14296 3714 14498 3731
rect 13538 3676 14498 3714
rect 14556 3714 14758 3731
rect 15314 3731 15330 3748
rect 15760 3748 16348 3764
rect 15760 3731 15776 3748
rect 15314 3714 15516 3731
rect 14556 3676 15516 3714
rect 15574 3714 15776 3731
rect 16332 3731 16348 3748
rect 16778 3748 17366 3764
rect 16778 3731 16794 3748
rect 16332 3714 16534 3731
rect 15574 3676 16534 3714
rect 16592 3714 16794 3731
rect 17350 3731 17366 3748
rect 17796 3748 18384 3764
rect 17796 3731 17812 3748
rect 17350 3714 17552 3731
rect 16592 3676 17552 3714
rect 17610 3714 17812 3731
rect 18368 3731 18384 3748
rect 18814 3748 19402 3764
rect 18814 3731 18830 3748
rect 18368 3714 18570 3731
rect 17610 3676 18570 3714
rect 18628 3714 18830 3731
rect 19386 3731 19402 3748
rect 19832 3748 20420 3764
rect 19832 3731 19848 3748
rect 19386 3714 19588 3731
rect 18628 3676 19588 3714
rect 19646 3714 19848 3731
rect 20404 3731 20420 3748
rect 20850 3748 21438 3764
rect 20850 3731 20866 3748
rect 20404 3714 20606 3731
rect 19646 3676 20606 3714
rect 20664 3714 20866 3731
rect 21422 3731 21438 3748
rect 21868 3748 22456 3764
rect 21868 3731 21884 3748
rect 21422 3714 21624 3731
rect 20664 3676 21624 3714
rect 21682 3714 21884 3731
rect 22440 3731 22456 3748
rect 22886 3748 23474 3764
rect 22886 3731 22902 3748
rect 22440 3714 22642 3731
rect 21682 3676 22642 3714
rect 22700 3714 22902 3731
rect 23458 3731 23474 3748
rect 23904 3748 24492 3764
rect 23904 3731 23920 3748
rect 23458 3714 23660 3731
rect 22700 3676 23660 3714
rect 23718 3714 23920 3731
rect 24476 3731 24492 3748
rect 24922 3748 25510 3764
rect 24922 3731 24938 3748
rect 24476 3714 24678 3731
rect 23718 3676 24678 3714
rect 24736 3714 24938 3731
rect 25494 3731 25510 3748
rect 25940 3748 26528 3764
rect 25940 3731 25956 3748
rect 25494 3714 25696 3731
rect 24736 3676 25696 3714
rect 25754 3714 25956 3731
rect 26512 3731 26528 3748
rect 26958 3748 27546 3764
rect 26958 3731 26974 3748
rect 26512 3714 26714 3731
rect 25754 3676 26714 3714
rect 26772 3714 26974 3731
rect 27530 3731 27546 3748
rect 27976 3748 28564 3764
rect 27976 3731 27992 3748
rect 27530 3714 27732 3731
rect 26772 3676 27732 3714
rect 27790 3714 27992 3731
rect 28548 3731 28564 3748
rect 28994 3748 29582 3764
rect 28994 3731 29010 3748
rect 28548 3714 28750 3731
rect 27790 3676 28750 3714
rect 28808 3714 29010 3731
rect 29566 3731 29582 3748
rect 30012 3748 30600 3764
rect 30012 3731 30028 3748
rect 29566 3714 29768 3731
rect 28808 3676 29768 3714
rect 29826 3714 30028 3731
rect 30584 3731 30600 3748
rect 31030 3748 31618 3764
rect 31030 3731 31046 3748
rect 30584 3714 30786 3731
rect 29826 3676 30786 3714
rect 30844 3714 31046 3731
rect 31602 3731 31618 3748
rect 32048 3748 32636 3764
rect 32048 3731 32064 3748
rect 31602 3714 31804 3731
rect 30844 3676 31804 3714
rect 31862 3714 32064 3731
rect 32620 3731 32636 3748
rect 33066 3748 33654 3764
rect 33066 3731 33082 3748
rect 32620 3714 32822 3731
rect 31862 3676 32822 3714
rect 32880 3714 33082 3731
rect 33638 3731 33654 3748
rect 33638 3714 33840 3731
rect 32880 3676 33840 3714
rect 450 3416 1410 3454
rect 450 3399 652 3416
rect 636 3382 652 3399
rect 1208 3399 1410 3416
rect 1468 3416 2428 3454
rect 1468 3399 1670 3416
rect 1208 3382 1224 3399
rect 636 3366 1224 3382
rect 1654 3382 1670 3399
rect 2226 3399 2428 3416
rect 2486 3416 3446 3454
rect 2486 3399 2688 3416
rect 2226 3382 2242 3399
rect 1654 3366 2242 3382
rect 2672 3382 2688 3399
rect 3244 3399 3446 3416
rect 3504 3416 4464 3454
rect 3504 3399 3706 3416
rect 3244 3382 3260 3399
rect 2672 3366 3260 3382
rect 3690 3382 3706 3399
rect 4262 3399 4464 3416
rect 4522 3416 5482 3454
rect 4522 3399 4724 3416
rect 4262 3382 4278 3399
rect 3690 3366 4278 3382
rect 4708 3382 4724 3399
rect 5280 3399 5482 3416
rect 5540 3416 6500 3454
rect 5540 3399 5742 3416
rect 5280 3382 5296 3399
rect 4708 3366 5296 3382
rect 5726 3382 5742 3399
rect 6298 3399 6500 3416
rect 6558 3416 7518 3454
rect 6558 3399 6760 3416
rect 6298 3382 6314 3399
rect 5726 3366 6314 3382
rect 6744 3382 6760 3399
rect 7316 3399 7518 3416
rect 7576 3416 8536 3454
rect 7576 3399 7778 3416
rect 7316 3382 7332 3399
rect 6744 3366 7332 3382
rect 7762 3382 7778 3399
rect 8334 3399 8536 3416
rect 8594 3416 9554 3454
rect 8594 3399 8796 3416
rect 8334 3382 8350 3399
rect 7762 3366 8350 3382
rect 8780 3382 8796 3399
rect 9352 3399 9554 3416
rect 9612 3416 10572 3454
rect 9612 3399 9814 3416
rect 9352 3382 9368 3399
rect 8780 3366 9368 3382
rect 9798 3382 9814 3399
rect 10370 3399 10572 3416
rect 10630 3416 11590 3454
rect 10630 3399 10832 3416
rect 10370 3382 10386 3399
rect 9798 3366 10386 3382
rect 10816 3382 10832 3399
rect 11388 3399 11590 3416
rect 11388 3382 11404 3399
rect 10816 3366 11404 3382
rect 13538 3038 14498 3076
rect 636 3014 1224 3030
rect 636 2997 652 3014
rect 450 2980 652 2997
rect 1208 2997 1224 3014
rect 1654 3014 2242 3030
rect 1654 2997 1670 3014
rect 1208 2980 1410 2997
rect 450 2942 1410 2980
rect 1468 2980 1670 2997
rect 2226 2997 2242 3014
rect 2672 3014 3260 3030
rect 2672 2997 2688 3014
rect 2226 2980 2428 2997
rect 1468 2942 2428 2980
rect 2486 2980 2688 2997
rect 3244 2997 3260 3014
rect 3690 3014 4278 3030
rect 3690 2997 3706 3014
rect 3244 2980 3446 2997
rect 2486 2942 3446 2980
rect 3504 2980 3706 2997
rect 4262 2997 4278 3014
rect 4708 3014 5296 3030
rect 4708 2997 4724 3014
rect 4262 2980 4464 2997
rect 3504 2942 4464 2980
rect 4522 2980 4724 2997
rect 5280 2997 5296 3014
rect 5726 3014 6314 3030
rect 5726 2997 5742 3014
rect 5280 2980 5482 2997
rect 4522 2942 5482 2980
rect 5540 2980 5742 2997
rect 6298 2997 6314 3014
rect 6744 3014 7332 3030
rect 6744 2997 6760 3014
rect 6298 2980 6500 2997
rect 5540 2942 6500 2980
rect 6558 2980 6760 2997
rect 7316 2997 7332 3014
rect 7762 3014 8350 3030
rect 7762 2997 7778 3014
rect 7316 2980 7518 2997
rect 6558 2942 7518 2980
rect 7576 2980 7778 2997
rect 8334 2997 8350 3014
rect 8780 3014 9368 3030
rect 8780 2997 8796 3014
rect 8334 2980 8536 2997
rect 7576 2942 8536 2980
rect 8594 2980 8796 2997
rect 9352 2997 9368 3014
rect 9798 3014 10386 3030
rect 9798 2997 9814 3014
rect 9352 2980 9554 2997
rect 8594 2942 9554 2980
rect 9612 2980 9814 2997
rect 10370 2997 10386 3014
rect 10816 3014 11404 3030
rect 13538 3021 13740 3038
rect 10816 2997 10832 3014
rect 10370 2980 10572 2997
rect 9612 2942 10572 2980
rect 10630 2980 10832 2997
rect 11388 2997 11404 3014
rect 13724 3004 13740 3021
rect 14296 3021 14498 3038
rect 14556 3038 15516 3076
rect 14556 3021 14758 3038
rect 14296 3004 14312 3021
rect 11388 2980 11590 2997
rect 13724 2988 14312 3004
rect 14742 3004 14758 3021
rect 15314 3021 15516 3038
rect 15574 3038 16534 3076
rect 15574 3021 15776 3038
rect 15314 3004 15330 3021
rect 14742 2988 15330 3004
rect 15760 3004 15776 3021
rect 16332 3021 16534 3038
rect 16592 3038 17552 3076
rect 16592 3021 16794 3038
rect 16332 3004 16348 3021
rect 15760 2988 16348 3004
rect 16778 3004 16794 3021
rect 17350 3021 17552 3038
rect 17610 3038 18570 3076
rect 17610 3021 17812 3038
rect 17350 3004 17366 3021
rect 16778 2988 17366 3004
rect 17796 3004 17812 3021
rect 18368 3021 18570 3038
rect 18628 3038 19588 3076
rect 18628 3021 18830 3038
rect 18368 3004 18384 3021
rect 17796 2988 18384 3004
rect 18814 3004 18830 3021
rect 19386 3021 19588 3038
rect 19646 3038 20606 3076
rect 19646 3021 19848 3038
rect 19386 3004 19402 3021
rect 18814 2988 19402 3004
rect 19832 3004 19848 3021
rect 20404 3021 20606 3038
rect 20664 3038 21624 3076
rect 20664 3021 20866 3038
rect 20404 3004 20420 3021
rect 19832 2988 20420 3004
rect 20850 3004 20866 3021
rect 21422 3021 21624 3038
rect 21682 3038 22642 3076
rect 21682 3021 21884 3038
rect 21422 3004 21438 3021
rect 20850 2988 21438 3004
rect 21868 3004 21884 3021
rect 22440 3021 22642 3038
rect 22700 3038 23660 3076
rect 22700 3021 22902 3038
rect 22440 3004 22456 3021
rect 21868 2988 22456 3004
rect 22886 3004 22902 3021
rect 23458 3021 23660 3038
rect 23718 3038 24678 3076
rect 23718 3021 23920 3038
rect 23458 3004 23474 3021
rect 22886 2988 23474 3004
rect 23904 3004 23920 3021
rect 24476 3021 24678 3038
rect 24736 3038 25696 3076
rect 24736 3021 24938 3038
rect 24476 3004 24492 3021
rect 23904 2988 24492 3004
rect 24922 3004 24938 3021
rect 25494 3021 25696 3038
rect 25754 3038 26714 3076
rect 25754 3021 25956 3038
rect 25494 3004 25510 3021
rect 24922 2988 25510 3004
rect 25940 3004 25956 3021
rect 26512 3021 26714 3038
rect 26772 3038 27732 3076
rect 26772 3021 26974 3038
rect 26512 3004 26528 3021
rect 25940 2988 26528 3004
rect 26958 3004 26974 3021
rect 27530 3021 27732 3038
rect 27790 3038 28750 3076
rect 27790 3021 27992 3038
rect 27530 3004 27546 3021
rect 26958 2988 27546 3004
rect 27976 3004 27992 3021
rect 28548 3021 28750 3038
rect 28808 3038 29768 3076
rect 28808 3021 29010 3038
rect 28548 3004 28564 3021
rect 27976 2988 28564 3004
rect 28994 3004 29010 3021
rect 29566 3021 29768 3038
rect 29826 3038 30786 3076
rect 29826 3021 30028 3038
rect 29566 3004 29582 3021
rect 28994 2988 29582 3004
rect 30012 3004 30028 3021
rect 30584 3021 30786 3038
rect 30844 3038 31804 3076
rect 30844 3021 31046 3038
rect 30584 3004 30600 3021
rect 30012 2988 30600 3004
rect 31030 3004 31046 3021
rect 31602 3021 31804 3038
rect 31862 3038 32822 3076
rect 31862 3021 32064 3038
rect 31602 3004 31618 3021
rect 31030 2988 31618 3004
rect 32048 3004 32064 3021
rect 32620 3021 32822 3038
rect 32880 3038 33840 3076
rect 32880 3021 33082 3038
rect 32620 3004 32636 3021
rect 32048 2988 32636 3004
rect 33066 3004 33082 3021
rect 33638 3021 33840 3038
rect 33638 3004 33654 3021
rect 33066 2988 33654 3004
rect 10630 2942 11590 2980
rect 13724 2514 14312 2530
rect 13724 2497 13740 2514
rect 13538 2480 13740 2497
rect 14296 2497 14312 2514
rect 14742 2514 15330 2530
rect 14742 2497 14758 2514
rect 14296 2480 14498 2497
rect 13538 2442 14498 2480
rect 14556 2480 14758 2497
rect 15314 2497 15330 2514
rect 15760 2514 16348 2530
rect 15760 2497 15776 2514
rect 15314 2480 15516 2497
rect 14556 2442 15516 2480
rect 15574 2480 15776 2497
rect 16332 2497 16348 2514
rect 16778 2514 17366 2530
rect 16778 2497 16794 2514
rect 16332 2480 16534 2497
rect 15574 2442 16534 2480
rect 16592 2480 16794 2497
rect 17350 2497 17366 2514
rect 17796 2514 18384 2530
rect 17796 2497 17812 2514
rect 17350 2480 17552 2497
rect 16592 2442 17552 2480
rect 17610 2480 17812 2497
rect 18368 2497 18384 2514
rect 18814 2514 19402 2530
rect 18814 2497 18830 2514
rect 18368 2480 18570 2497
rect 17610 2442 18570 2480
rect 18628 2480 18830 2497
rect 19386 2497 19402 2514
rect 19832 2514 20420 2530
rect 19832 2497 19848 2514
rect 19386 2480 19588 2497
rect 18628 2442 19588 2480
rect 19646 2480 19848 2497
rect 20404 2497 20420 2514
rect 20850 2514 21438 2530
rect 20850 2497 20866 2514
rect 20404 2480 20606 2497
rect 19646 2442 20606 2480
rect 20664 2480 20866 2497
rect 21422 2497 21438 2514
rect 21868 2514 22456 2530
rect 21868 2497 21884 2514
rect 21422 2480 21624 2497
rect 20664 2442 21624 2480
rect 21682 2480 21884 2497
rect 22440 2497 22456 2514
rect 22886 2514 23474 2530
rect 22886 2497 22902 2514
rect 22440 2480 22642 2497
rect 21682 2442 22642 2480
rect 22700 2480 22902 2497
rect 23458 2497 23474 2514
rect 23904 2514 24492 2530
rect 23904 2497 23920 2514
rect 23458 2480 23660 2497
rect 22700 2442 23660 2480
rect 23718 2480 23920 2497
rect 24476 2497 24492 2514
rect 24922 2514 25510 2530
rect 24922 2497 24938 2514
rect 24476 2480 24678 2497
rect 23718 2442 24678 2480
rect 24736 2480 24938 2497
rect 25494 2497 25510 2514
rect 25940 2514 26528 2530
rect 25940 2497 25956 2514
rect 25494 2480 25696 2497
rect 24736 2442 25696 2480
rect 25754 2480 25956 2497
rect 26512 2497 26528 2514
rect 26958 2514 27546 2530
rect 26958 2497 26974 2514
rect 26512 2480 26714 2497
rect 25754 2442 26714 2480
rect 26772 2480 26974 2497
rect 27530 2497 27546 2514
rect 27976 2514 28564 2530
rect 27976 2497 27992 2514
rect 27530 2480 27732 2497
rect 26772 2442 27732 2480
rect 27790 2480 27992 2497
rect 28548 2497 28564 2514
rect 28994 2514 29582 2530
rect 28994 2497 29010 2514
rect 28548 2480 28750 2497
rect 27790 2442 28750 2480
rect 28808 2480 29010 2497
rect 29566 2497 29582 2514
rect 30012 2514 30600 2530
rect 30012 2497 30028 2514
rect 29566 2480 29768 2497
rect 28808 2442 29768 2480
rect 29826 2480 30028 2497
rect 30584 2497 30600 2514
rect 31030 2514 31618 2530
rect 31030 2497 31046 2514
rect 30584 2480 30786 2497
rect 29826 2442 30786 2480
rect 30844 2480 31046 2497
rect 31602 2497 31618 2514
rect 32048 2514 32636 2530
rect 32048 2497 32064 2514
rect 31602 2480 31804 2497
rect 30844 2442 31804 2480
rect 31862 2480 32064 2497
rect 32620 2497 32636 2514
rect 33066 2514 33654 2530
rect 33066 2497 33082 2514
rect 32620 2480 32822 2497
rect 31862 2442 32822 2480
rect 32880 2480 33082 2497
rect 33638 2497 33654 2514
rect 33638 2480 33840 2497
rect 32880 2442 33840 2480
rect 450 2304 1410 2342
rect 450 2287 652 2304
rect 636 2270 652 2287
rect 1208 2287 1410 2304
rect 1468 2304 2428 2342
rect 1468 2287 1670 2304
rect 1208 2270 1224 2287
rect 636 2254 1224 2270
rect 1654 2270 1670 2287
rect 2226 2287 2428 2304
rect 2486 2304 3446 2342
rect 2486 2287 2688 2304
rect 2226 2270 2242 2287
rect 1654 2254 2242 2270
rect 2672 2270 2688 2287
rect 3244 2287 3446 2304
rect 3504 2304 4464 2342
rect 3504 2287 3706 2304
rect 3244 2270 3260 2287
rect 2672 2254 3260 2270
rect 3690 2270 3706 2287
rect 4262 2287 4464 2304
rect 4522 2304 5482 2342
rect 4522 2287 4724 2304
rect 4262 2270 4278 2287
rect 3690 2254 4278 2270
rect 4708 2270 4724 2287
rect 5280 2287 5482 2304
rect 5540 2304 6500 2342
rect 5540 2287 5742 2304
rect 5280 2270 5296 2287
rect 4708 2254 5296 2270
rect 5726 2270 5742 2287
rect 6298 2287 6500 2304
rect 6558 2304 7518 2342
rect 6558 2287 6760 2304
rect 6298 2270 6314 2287
rect 5726 2254 6314 2270
rect 6744 2270 6760 2287
rect 7316 2287 7518 2304
rect 7576 2304 8536 2342
rect 7576 2287 7778 2304
rect 7316 2270 7332 2287
rect 6744 2254 7332 2270
rect 7762 2270 7778 2287
rect 8334 2287 8536 2304
rect 8594 2304 9554 2342
rect 8594 2287 8796 2304
rect 8334 2270 8350 2287
rect 7762 2254 8350 2270
rect 8780 2270 8796 2287
rect 9352 2287 9554 2304
rect 9612 2304 10572 2342
rect 9612 2287 9814 2304
rect 9352 2270 9368 2287
rect 8780 2254 9368 2270
rect 9798 2270 9814 2287
rect 10370 2287 10572 2304
rect 10630 2304 11590 2342
rect 10630 2287 10832 2304
rect 10370 2270 10386 2287
rect 9798 2254 10386 2270
rect 10816 2270 10832 2287
rect 11388 2287 11590 2304
rect 11388 2270 11404 2287
rect 10816 2254 11404 2270
rect 13538 1804 14498 1842
rect 13538 1787 13740 1804
rect 13724 1770 13740 1787
rect 14296 1787 14498 1804
rect 14556 1804 15516 1842
rect 14556 1787 14758 1804
rect 14296 1770 14312 1787
rect 13724 1754 14312 1770
rect 14742 1770 14758 1787
rect 15314 1787 15516 1804
rect 15574 1804 16534 1842
rect 15574 1787 15776 1804
rect 15314 1770 15330 1787
rect 14742 1754 15330 1770
rect 15760 1770 15776 1787
rect 16332 1787 16534 1804
rect 16592 1804 17552 1842
rect 16592 1787 16794 1804
rect 16332 1770 16348 1787
rect 15760 1754 16348 1770
rect 16778 1770 16794 1787
rect 17350 1787 17552 1804
rect 17610 1804 18570 1842
rect 17610 1787 17812 1804
rect 17350 1770 17366 1787
rect 16778 1754 17366 1770
rect 17796 1770 17812 1787
rect 18368 1787 18570 1804
rect 18628 1804 19588 1842
rect 18628 1787 18830 1804
rect 18368 1770 18384 1787
rect 17796 1754 18384 1770
rect 18814 1770 18830 1787
rect 19386 1787 19588 1804
rect 19646 1804 20606 1842
rect 19646 1787 19848 1804
rect 19386 1770 19402 1787
rect 18814 1754 19402 1770
rect 19832 1770 19848 1787
rect 20404 1787 20606 1804
rect 20664 1804 21624 1842
rect 20664 1787 20866 1804
rect 20404 1770 20420 1787
rect 19832 1754 20420 1770
rect 20850 1770 20866 1787
rect 21422 1787 21624 1804
rect 21682 1804 22642 1842
rect 21682 1787 21884 1804
rect 21422 1770 21438 1787
rect 20850 1754 21438 1770
rect 21868 1770 21884 1787
rect 22440 1787 22642 1804
rect 22700 1804 23660 1842
rect 22700 1787 22902 1804
rect 22440 1770 22456 1787
rect 21868 1754 22456 1770
rect 22886 1770 22902 1787
rect 23458 1787 23660 1804
rect 23718 1804 24678 1842
rect 23718 1787 23920 1804
rect 23458 1770 23474 1787
rect 22886 1754 23474 1770
rect 23904 1770 23920 1787
rect 24476 1787 24678 1804
rect 24736 1804 25696 1842
rect 24736 1787 24938 1804
rect 24476 1770 24492 1787
rect 23904 1754 24492 1770
rect 24922 1770 24938 1787
rect 25494 1787 25696 1804
rect 25754 1804 26714 1842
rect 25754 1787 25956 1804
rect 25494 1770 25510 1787
rect 24922 1754 25510 1770
rect 25940 1770 25956 1787
rect 26512 1787 26714 1804
rect 26772 1804 27732 1842
rect 26772 1787 26974 1804
rect 26512 1770 26528 1787
rect 25940 1754 26528 1770
rect 26958 1770 26974 1787
rect 27530 1787 27732 1804
rect 27790 1804 28750 1842
rect 27790 1787 27992 1804
rect 27530 1770 27546 1787
rect 26958 1754 27546 1770
rect 27976 1770 27992 1787
rect 28548 1787 28750 1804
rect 28808 1804 29768 1842
rect 28808 1787 29010 1804
rect 28548 1770 28564 1787
rect 27976 1754 28564 1770
rect 28994 1770 29010 1787
rect 29566 1787 29768 1804
rect 29826 1804 30786 1842
rect 29826 1787 30028 1804
rect 29566 1770 29582 1787
rect 28994 1754 29582 1770
rect 30012 1770 30028 1787
rect 30584 1787 30786 1804
rect 30844 1804 31804 1842
rect 30844 1787 31046 1804
rect 30584 1770 30600 1787
rect 30012 1754 30600 1770
rect 31030 1770 31046 1787
rect 31602 1787 31804 1804
rect 31862 1804 32822 1842
rect 31862 1787 32064 1804
rect 31602 1770 31618 1787
rect 31030 1754 31618 1770
rect 32048 1770 32064 1787
rect 32620 1787 32822 1804
rect 32880 1804 33840 1842
rect 32880 1787 33082 1804
rect 32620 1770 32636 1787
rect 32048 1754 32636 1770
rect 33066 1770 33082 1787
rect 33638 1787 33840 1804
rect 33638 1770 33654 1787
rect 33066 1754 33654 1770
rect 1094 1472 1682 1488
rect 1094 1455 1110 1472
rect 908 1438 1110 1455
rect 1666 1455 1682 1472
rect 2112 1472 2700 1488
rect 2112 1455 2128 1472
rect 1666 1438 1868 1455
rect 908 1400 1868 1438
rect 1926 1438 2128 1455
rect 2684 1455 2700 1472
rect 3130 1472 3718 1488
rect 3130 1455 3146 1472
rect 2684 1438 2886 1455
rect 1926 1400 2886 1438
rect 2944 1438 3146 1455
rect 3702 1455 3718 1472
rect 4148 1472 4736 1488
rect 4148 1455 4164 1472
rect 3702 1438 3904 1455
rect 2944 1400 3904 1438
rect 3962 1438 4164 1455
rect 4720 1455 4736 1472
rect 5166 1472 5754 1488
rect 5166 1455 5182 1472
rect 4720 1438 4922 1455
rect 3962 1400 4922 1438
rect 4980 1438 5182 1455
rect 5738 1455 5754 1472
rect 6184 1472 6772 1488
rect 6184 1455 6200 1472
rect 5738 1438 5940 1455
rect 4980 1400 5940 1438
rect 5998 1438 6200 1455
rect 6756 1455 6772 1472
rect 7202 1472 7790 1488
rect 7202 1455 7218 1472
rect 6756 1438 6958 1455
rect 5998 1400 6958 1438
rect 7016 1438 7218 1455
rect 7774 1455 7790 1472
rect 8220 1472 8808 1488
rect 8220 1455 8236 1472
rect 7774 1438 7976 1455
rect 7016 1400 7976 1438
rect 8034 1438 8236 1455
rect 8792 1455 8808 1472
rect 9238 1472 9826 1488
rect 9238 1455 9254 1472
rect 8792 1438 8994 1455
rect 8034 1400 8994 1438
rect 9052 1438 9254 1455
rect 9810 1455 9826 1472
rect 10256 1472 10844 1488
rect 10256 1455 10272 1472
rect 9810 1438 10012 1455
rect 9052 1400 10012 1438
rect 10070 1438 10272 1455
rect 10828 1455 10844 1472
rect 10828 1438 11030 1455
rect 10070 1400 11030 1438
rect 13724 1282 14312 1298
rect 13724 1265 13740 1282
rect 13538 1248 13740 1265
rect 14296 1265 14312 1282
rect 14742 1282 15330 1298
rect 14742 1265 14758 1282
rect 14296 1248 14498 1265
rect 13538 1210 14498 1248
rect 14556 1248 14758 1265
rect 15314 1265 15330 1282
rect 15760 1282 16348 1298
rect 15760 1265 15776 1282
rect 15314 1248 15516 1265
rect 14556 1210 15516 1248
rect 15574 1248 15776 1265
rect 16332 1265 16348 1282
rect 16778 1282 17366 1298
rect 16778 1265 16794 1282
rect 16332 1248 16534 1265
rect 15574 1210 16534 1248
rect 16592 1248 16794 1265
rect 17350 1265 17366 1282
rect 17796 1282 18384 1298
rect 17796 1265 17812 1282
rect 17350 1248 17552 1265
rect 16592 1210 17552 1248
rect 17610 1248 17812 1265
rect 18368 1265 18384 1282
rect 18814 1282 19402 1298
rect 18814 1265 18830 1282
rect 18368 1248 18570 1265
rect 17610 1210 18570 1248
rect 18628 1248 18830 1265
rect 19386 1265 19402 1282
rect 19832 1282 20420 1298
rect 19832 1265 19848 1282
rect 19386 1248 19588 1265
rect 18628 1210 19588 1248
rect 19646 1248 19848 1265
rect 20404 1265 20420 1282
rect 20850 1282 21438 1298
rect 20850 1265 20866 1282
rect 20404 1248 20606 1265
rect 19646 1210 20606 1248
rect 20664 1248 20866 1265
rect 21422 1265 21438 1282
rect 21868 1282 22456 1298
rect 21868 1265 21884 1282
rect 21422 1248 21624 1265
rect 20664 1210 21624 1248
rect 21682 1248 21884 1265
rect 22440 1265 22456 1282
rect 22886 1282 23474 1298
rect 22886 1265 22902 1282
rect 22440 1248 22642 1265
rect 21682 1210 22642 1248
rect 22700 1248 22902 1265
rect 23458 1265 23474 1282
rect 23904 1282 24492 1298
rect 23904 1265 23920 1282
rect 23458 1248 23660 1265
rect 22700 1210 23660 1248
rect 23718 1248 23920 1265
rect 24476 1265 24492 1282
rect 24922 1282 25510 1298
rect 24922 1265 24938 1282
rect 24476 1248 24678 1265
rect 23718 1210 24678 1248
rect 24736 1248 24938 1265
rect 25494 1265 25510 1282
rect 25940 1282 26528 1298
rect 25940 1265 25956 1282
rect 25494 1248 25696 1265
rect 24736 1210 25696 1248
rect 25754 1248 25956 1265
rect 26512 1265 26528 1282
rect 26958 1282 27546 1298
rect 26958 1265 26974 1282
rect 26512 1248 26714 1265
rect 25754 1210 26714 1248
rect 26772 1248 26974 1265
rect 27530 1265 27546 1282
rect 27976 1282 28564 1298
rect 27976 1265 27992 1282
rect 27530 1248 27732 1265
rect 26772 1210 27732 1248
rect 27790 1248 27992 1265
rect 28548 1265 28564 1282
rect 28994 1282 29582 1298
rect 28994 1265 29010 1282
rect 28548 1248 28750 1265
rect 27790 1210 28750 1248
rect 28808 1248 29010 1265
rect 29566 1265 29582 1282
rect 30012 1282 30600 1298
rect 30012 1265 30028 1282
rect 29566 1248 29768 1265
rect 28808 1210 29768 1248
rect 29826 1248 30028 1265
rect 30584 1265 30600 1282
rect 31030 1282 31618 1298
rect 31030 1265 31046 1282
rect 30584 1248 30786 1265
rect 29826 1210 30786 1248
rect 30844 1248 31046 1265
rect 31602 1265 31618 1282
rect 32048 1282 32636 1298
rect 32048 1265 32064 1282
rect 31602 1248 31804 1265
rect 30844 1210 31804 1248
rect 31862 1248 32064 1265
rect 32620 1265 32636 1282
rect 33066 1282 33654 1298
rect 33066 1265 33082 1282
rect 32620 1248 32822 1265
rect 31862 1210 32822 1248
rect 32880 1248 33082 1265
rect 33638 1265 33654 1282
rect 33638 1248 33840 1265
rect 32880 1210 33840 1248
rect 908 762 1868 800
rect 908 745 1110 762
rect 1094 728 1110 745
rect 1666 745 1868 762
rect 1926 762 2886 800
rect 1926 745 2128 762
rect 1666 728 1682 745
rect 1094 712 1682 728
rect 2112 728 2128 745
rect 2684 745 2886 762
rect 2944 762 3904 800
rect 2944 745 3146 762
rect 2684 728 2700 745
rect 2112 712 2700 728
rect 3130 728 3146 745
rect 3702 745 3904 762
rect 3962 762 4922 800
rect 3962 745 4164 762
rect 3702 728 3718 745
rect 3130 712 3718 728
rect 4148 728 4164 745
rect 4720 745 4922 762
rect 4980 762 5940 800
rect 4980 745 5182 762
rect 4720 728 4736 745
rect 4148 712 4736 728
rect 5166 728 5182 745
rect 5738 745 5940 762
rect 5998 762 6958 800
rect 5998 745 6200 762
rect 5738 728 5754 745
rect 5166 712 5754 728
rect 6184 728 6200 745
rect 6756 745 6958 762
rect 7016 762 7976 800
rect 7016 745 7218 762
rect 6756 728 6772 745
rect 6184 712 6772 728
rect 7202 728 7218 745
rect 7774 745 7976 762
rect 8034 762 8994 800
rect 8034 745 8236 762
rect 7774 728 7790 745
rect 7202 712 7790 728
rect 8220 728 8236 745
rect 8792 745 8994 762
rect 9052 762 10012 800
rect 9052 745 9254 762
rect 8792 728 8808 745
rect 8220 712 8808 728
rect 9238 728 9254 745
rect 9810 745 10012 762
rect 10070 762 11030 800
rect 10070 745 10272 762
rect 9810 728 9826 745
rect 9238 712 9826 728
rect 10256 728 10272 745
rect 10828 745 11030 762
rect 10828 728 10844 745
rect 10256 712 10844 728
rect 13538 572 14498 610
rect 13538 555 13740 572
rect 13724 538 13740 555
rect 14296 555 14498 572
rect 14556 572 15516 610
rect 14556 555 14758 572
rect 14296 538 14312 555
rect 13724 522 14312 538
rect 14742 538 14758 555
rect 15314 555 15516 572
rect 15574 572 16534 610
rect 15574 555 15776 572
rect 15314 538 15330 555
rect 14742 522 15330 538
rect 15760 538 15776 555
rect 16332 555 16534 572
rect 16592 572 17552 610
rect 16592 555 16794 572
rect 16332 538 16348 555
rect 15760 522 16348 538
rect 16778 538 16794 555
rect 17350 555 17552 572
rect 17610 572 18570 610
rect 17610 555 17812 572
rect 17350 538 17366 555
rect 16778 522 17366 538
rect 17796 538 17812 555
rect 18368 555 18570 572
rect 18628 572 19588 610
rect 18628 555 18830 572
rect 18368 538 18384 555
rect 17796 522 18384 538
rect 18814 538 18830 555
rect 19386 555 19588 572
rect 19646 572 20606 610
rect 19646 555 19848 572
rect 19386 538 19402 555
rect 18814 522 19402 538
rect 19832 538 19848 555
rect 20404 555 20606 572
rect 20664 572 21624 610
rect 20664 555 20866 572
rect 20404 538 20420 555
rect 19832 522 20420 538
rect 20850 538 20866 555
rect 21422 555 21624 572
rect 21682 572 22642 610
rect 21682 555 21884 572
rect 21422 538 21438 555
rect 20850 522 21438 538
rect 21868 538 21884 555
rect 22440 555 22642 572
rect 22700 572 23660 610
rect 22700 555 22902 572
rect 22440 538 22456 555
rect 21868 522 22456 538
rect 22886 538 22902 555
rect 23458 555 23660 572
rect 23718 572 24678 610
rect 23718 555 23920 572
rect 23458 538 23474 555
rect 22886 522 23474 538
rect 23904 538 23920 555
rect 24476 555 24678 572
rect 24736 572 25696 610
rect 24736 555 24938 572
rect 24476 538 24492 555
rect 23904 522 24492 538
rect 24922 538 24938 555
rect 25494 555 25696 572
rect 25754 572 26714 610
rect 25754 555 25956 572
rect 25494 538 25510 555
rect 24922 522 25510 538
rect 25940 538 25956 555
rect 26512 555 26714 572
rect 26772 572 27732 610
rect 26772 555 26974 572
rect 26512 538 26528 555
rect 25940 522 26528 538
rect 26958 538 26974 555
rect 27530 555 27732 572
rect 27790 572 28750 610
rect 27790 555 27992 572
rect 27530 538 27546 555
rect 26958 522 27546 538
rect 27976 538 27992 555
rect 28548 555 28750 572
rect 28808 572 29768 610
rect 28808 555 29010 572
rect 28548 538 28564 555
rect 27976 522 28564 538
rect 28994 538 29010 555
rect 29566 555 29768 572
rect 29826 572 30786 610
rect 29826 555 30028 572
rect 29566 538 29582 555
rect 28994 522 29582 538
rect 30012 538 30028 555
rect 30584 555 30786 572
rect 30844 572 31804 610
rect 30844 555 31046 572
rect 30584 538 30600 555
rect 30012 522 30600 538
rect 31030 538 31046 555
rect 31602 555 31804 572
rect 31862 572 32822 610
rect 31862 555 32064 572
rect 31602 538 31618 555
rect 31030 522 31618 538
rect 32048 538 32064 555
rect 32620 555 32822 572
rect 32880 572 33840 610
rect 32880 555 33082 572
rect 32620 538 32636 555
rect 32048 522 32636 538
rect 33066 538 33082 555
rect 33638 555 33840 572
rect 33638 538 33654 555
rect 33066 522 33654 538
<< polycont >>
rect 17648 28061 18204 28095
rect 18666 28061 19222 28095
rect 19684 28061 20240 28095
rect 20702 28061 21258 28095
rect 21720 28061 22276 28095
rect 22738 28061 23294 28095
rect 23756 28061 24312 28095
rect 24774 28061 25330 28095
rect 25792 28061 26348 28095
rect 26810 28061 27366 28095
rect 27828 28061 28384 28095
rect 28846 28061 29402 28095
rect 29864 28061 30420 28095
rect 30882 28061 31438 28095
rect 31900 28061 32456 28095
rect 32918 28061 33474 28095
rect 17648 27333 18204 27367
rect 18666 27333 19222 27367
rect 19684 27333 20240 27367
rect 20702 27333 21258 27367
rect 21720 27333 22276 27367
rect 22738 27333 23294 27367
rect 23756 27333 24312 27367
rect 24774 27333 25330 27367
rect 25792 27333 26348 27367
rect 26810 27333 27366 27367
rect 27828 27333 28384 27367
rect 28846 27333 29402 27367
rect 29864 27333 30420 27367
rect 30882 27333 31438 27367
rect 31900 27333 32456 27367
rect 32918 27333 33474 27367
rect 17648 26925 18204 26959
rect 18666 26925 19222 26959
rect 19684 26925 20240 26959
rect 20702 26925 21258 26959
rect 21720 26925 22276 26959
rect 22738 26925 23294 26959
rect 23756 26925 24312 26959
rect 24774 26925 25330 26959
rect 25792 26925 26348 26959
rect 26810 26925 27366 26959
rect 27828 26925 28384 26959
rect 28846 26925 29402 26959
rect 29864 26925 30420 26959
rect 30882 26925 31438 26959
rect 31900 26925 32456 26959
rect 32918 26925 33474 26959
rect 17648 26197 18204 26231
rect 18666 26197 19222 26231
rect 19684 26197 20240 26231
rect 20702 26197 21258 26231
rect 21720 26197 22276 26231
rect 22738 26197 23294 26231
rect 23756 26197 24312 26231
rect 24774 26197 25330 26231
rect 25792 26197 26348 26231
rect 26810 26197 27366 26231
rect 27828 26197 28384 26231
rect 28846 26197 29402 26231
rect 29864 26197 30420 26231
rect 30882 26197 31438 26231
rect 31900 26197 32456 26231
rect 32918 26197 33474 26231
rect 17648 25789 18204 25823
rect 18666 25789 19222 25823
rect 19684 25789 20240 25823
rect 20702 25789 21258 25823
rect 21720 25789 22276 25823
rect 22738 25789 23294 25823
rect 23756 25789 24312 25823
rect 24774 25789 25330 25823
rect 25792 25789 26348 25823
rect 26810 25789 27366 25823
rect 27828 25789 28384 25823
rect 28846 25789 29402 25823
rect 29864 25789 30420 25823
rect 30882 25789 31438 25823
rect 31900 25789 32456 25823
rect 32918 25789 33474 25823
rect 17648 25061 18204 25095
rect 18666 25061 19222 25095
rect 19684 25061 20240 25095
rect 20702 25061 21258 25095
rect 21720 25061 22276 25095
rect 22738 25061 23294 25095
rect 23756 25061 24312 25095
rect 24774 25061 25330 25095
rect 25792 25061 26348 25095
rect 26810 25061 27366 25095
rect 27828 25061 28384 25095
rect 28846 25061 29402 25095
rect 29864 25061 30420 25095
rect 30882 25061 31438 25095
rect 31900 25061 32456 25095
rect 32918 25061 33474 25095
rect 18842 24151 19398 24185
rect 19860 24151 20416 24185
rect 20878 24151 21434 24185
rect 21896 24151 22452 24185
rect 22914 24151 23470 24185
rect 23932 24151 24488 24185
rect 24950 24151 25506 24185
rect 25968 24151 26524 24185
rect 26986 24151 27542 24185
rect 28004 24151 28560 24185
rect 29022 24151 29578 24185
rect 30040 24151 30596 24185
rect 31058 24151 31614 24185
rect 32076 24151 32632 24185
rect 18842 23423 19398 23457
rect 19860 23423 20416 23457
rect 20878 23423 21434 23457
rect 21896 23423 22452 23457
rect 22914 23423 23470 23457
rect 23932 23423 24488 23457
rect 24950 23423 25506 23457
rect 25968 23423 26524 23457
rect 26986 23423 27542 23457
rect 28004 23423 28560 23457
rect 29022 23423 29578 23457
rect 30040 23423 30596 23457
rect 31058 23423 31614 23457
rect 32076 23423 32632 23457
rect 18842 23119 19398 23153
rect 19860 23119 20416 23153
rect 20878 23119 21434 23153
rect 21896 23119 22452 23153
rect 22914 23119 23470 23153
rect 23932 23119 24488 23153
rect 24950 23119 25506 23153
rect 25968 23119 26524 23153
rect 26986 23119 27542 23153
rect 28004 23119 28560 23153
rect 29022 23119 29578 23153
rect 30040 23119 30596 23153
rect 31058 23119 31614 23153
rect 32076 23119 32632 23153
rect 18842 22391 19398 22425
rect 19860 22391 20416 22425
rect 20878 22391 21434 22425
rect 21896 22391 22452 22425
rect 22914 22391 23470 22425
rect 23932 22391 24488 22425
rect 24950 22391 25506 22425
rect 25968 22391 26524 22425
rect 26986 22391 27542 22425
rect 28004 22391 28560 22425
rect 29022 22391 29578 22425
rect 30040 22391 30596 22425
rect 31058 22391 31614 22425
rect 32076 22391 32632 22425
rect 18634 21515 19190 21549
rect 19652 21515 20208 21549
rect 20670 21515 21226 21549
rect 21688 21515 22244 21549
rect 22706 21515 23262 21549
rect 23724 21515 24280 21549
rect 24742 21515 25298 21549
rect 25760 21515 26316 21549
rect 26778 21515 27334 21549
rect 27796 21515 28352 21549
rect 28814 21515 29370 21549
rect 29832 21515 30388 21549
rect 30850 21515 31406 21549
rect 31868 21515 32424 21549
rect 32886 21515 33442 21549
rect 13330 21411 13886 21445
rect 14348 21411 14904 21445
rect 15366 21411 15922 21445
rect 16384 21411 16940 21445
rect 18634 20787 19190 20821
rect 19652 20787 20208 20821
rect 20670 20787 21226 20821
rect 21688 20787 22244 20821
rect 22706 20787 23262 20821
rect 23724 20787 24280 20821
rect 24742 20787 25298 20821
rect 25760 20787 26316 20821
rect 26778 20787 27334 20821
rect 27796 20787 28352 20821
rect 28814 20787 29370 20821
rect 29832 20787 30388 20821
rect 30850 20787 31406 20821
rect 31868 20787 32424 20821
rect 32886 20787 33442 20821
rect 13330 20683 13886 20717
rect 14348 20683 14904 20717
rect 15366 20683 15922 20717
rect 16384 20683 16940 20717
rect 13330 20379 13886 20413
rect 14348 20379 14904 20413
rect 15366 20379 15922 20413
rect 16384 20379 16940 20413
rect 18634 20259 19190 20293
rect 19652 20259 20208 20293
rect 20670 20259 21226 20293
rect 21688 20259 22244 20293
rect 22706 20259 23262 20293
rect 23724 20259 24280 20293
rect 24742 20259 25298 20293
rect 25760 20259 26316 20293
rect 26778 20259 27334 20293
rect 27796 20259 28352 20293
rect 28814 20259 29370 20293
rect 29832 20259 30388 20293
rect 30850 20259 31406 20293
rect 31868 20259 32424 20293
rect 32886 20259 33442 20293
rect 13330 19651 13886 19685
rect 14348 19651 14904 19685
rect 15366 19651 15922 19685
rect 16384 19651 16940 19685
rect 18634 19531 19190 19565
rect 19652 19531 20208 19565
rect 20670 19531 21226 19565
rect 21688 19531 22244 19565
rect 22706 19531 23262 19565
rect 23724 19531 24280 19565
rect 24742 19531 25298 19565
rect 25760 19531 26316 19565
rect 26778 19531 27334 19565
rect 27796 19531 28352 19565
rect 28814 19531 29370 19565
rect 29832 19531 30388 19565
rect 30850 19531 31406 19565
rect 31868 19531 32424 19565
rect 32886 19531 33442 19565
rect 13330 19347 13886 19381
rect 14348 19347 14904 19381
rect 15366 19347 15922 19381
rect 16384 19347 16940 19381
rect 18634 19003 19190 19037
rect 19652 19003 20208 19037
rect 20670 19003 21226 19037
rect 21688 19003 22244 19037
rect 22706 19003 23262 19037
rect 23724 19003 24280 19037
rect 24742 19003 25298 19037
rect 25760 19003 26316 19037
rect 26778 19003 27334 19037
rect 27796 19003 28352 19037
rect 28814 19003 29370 19037
rect 29832 19003 30388 19037
rect 30850 19003 31406 19037
rect 31868 19003 32424 19037
rect 32886 19003 33442 19037
rect 13330 18619 13886 18653
rect 14348 18619 14904 18653
rect 15366 18619 15922 18653
rect 16384 18619 16940 18653
rect 13330 18315 13886 18349
rect 14348 18315 14904 18349
rect 15366 18315 15922 18349
rect 16384 18315 16940 18349
rect 18634 18275 19190 18309
rect 19652 18275 20208 18309
rect 20670 18275 21226 18309
rect 21688 18275 22244 18309
rect 22706 18275 23262 18309
rect 23724 18275 24280 18309
rect 24742 18275 25298 18309
rect 25760 18275 26316 18309
rect 26778 18275 27334 18309
rect 27796 18275 28352 18309
rect 28814 18275 29370 18309
rect 29832 18275 30388 18309
rect 30850 18275 31406 18309
rect 31868 18275 32424 18309
rect 32886 18275 33442 18309
rect 18634 17747 19190 17781
rect 19652 17747 20208 17781
rect 20670 17747 21226 17781
rect 21688 17747 22244 17781
rect 22706 17747 23262 17781
rect 23724 17747 24280 17781
rect 24742 17747 25298 17781
rect 25760 17747 26316 17781
rect 26778 17747 27334 17781
rect 27796 17747 28352 17781
rect 28814 17747 29370 17781
rect 29832 17747 30388 17781
rect 30850 17747 31406 17781
rect 31868 17747 32424 17781
rect 32886 17747 33442 17781
rect 13330 17587 13886 17621
rect 14348 17587 14904 17621
rect 15366 17587 15922 17621
rect 16384 17587 16940 17621
rect 18634 17019 19190 17053
rect 19652 17019 20208 17053
rect 20670 17019 21226 17053
rect 21688 17019 22244 17053
rect 22706 17019 23262 17053
rect 23724 17019 24280 17053
rect 24742 17019 25298 17053
rect 25760 17019 26316 17053
rect 26778 17019 27334 17053
rect 27796 17019 28352 17053
rect 28814 17019 29370 17053
rect 29832 17019 30388 17053
rect 30850 17019 31406 17053
rect 31868 17019 32424 17053
rect 32886 17019 33442 17053
rect -12070 16173 -11970 16207
rect -11812 16173 -11712 16207
rect -11554 16173 -11454 16207
rect -11296 16173 -11196 16207
rect -11038 16173 -10938 16207
rect -10780 16173 -10680 16207
rect -12070 15645 -11970 15679
rect -11812 15645 -11712 15679
rect -11554 15645 -11454 15679
rect -11296 15645 -11196 15679
rect -11038 15645 -10938 15679
rect -10780 15645 -10680 15679
rect -9470 16173 -9370 16207
rect -9212 16173 -9112 16207
rect -8954 16173 -8854 16207
rect -8696 16173 -8596 16207
rect -8438 16173 -8338 16207
rect -8180 16173 -8080 16207
rect -9470 15645 -9370 15679
rect -9212 15645 -9112 15679
rect -8954 15645 -8854 15679
rect -8696 15645 -8596 15679
rect -8438 15645 -8338 15679
rect -8180 15645 -8080 15679
rect -10234 15461 -10200 15495
rect -7634 15461 -7600 15495
rect -7184 15461 -7150 15495
rect -12070 15240 -11970 15274
rect -11812 15240 -11712 15274
rect -11554 15240 -11454 15274
rect -11296 15240 -11196 15274
rect -11038 15240 -10938 15274
rect -10780 15240 -10680 15274
rect -12070 14930 -11970 14964
rect -11812 14930 -11712 14964
rect -11554 14930 -11454 14964
rect -11296 14930 -11196 14964
rect -11038 14930 -10938 14964
rect -10780 14930 -10680 14964
rect -9470 15240 -9370 15274
rect -9212 15240 -9112 15274
rect -8954 15240 -8854 15274
rect -8696 15240 -8596 15274
rect -8438 15240 -8338 15274
rect -8180 15240 -8080 15274
rect -9470 14930 -9370 14964
rect -9212 14930 -9112 14964
rect -8954 14930 -8854 14964
rect -8696 14930 -8596 14964
rect -8438 14930 -8338 14964
rect -8180 14930 -8080 14964
rect 13742 14542 14298 14576
rect 14760 14542 15316 14576
rect 15778 14542 16334 14576
rect 16796 14542 17352 14576
rect 17814 14542 18370 14576
rect 18832 14542 19388 14576
rect 19850 14542 20406 14576
rect 20868 14542 21424 14576
rect 21886 14542 22442 14576
rect 22904 14542 23460 14576
rect 23922 14542 24478 14576
rect 24940 14542 25496 14576
rect 25958 14542 26514 14576
rect 26976 14542 27532 14576
rect 27994 14542 28550 14576
rect 29012 14542 29568 14576
rect 30030 14542 30586 14576
rect 31048 14542 31604 14576
rect 32066 14542 32622 14576
rect 33084 14542 33640 14576
rect 1976 14066 2532 14100
rect 2994 14066 3550 14100
rect 4012 14066 4568 14100
rect 5030 14066 5586 14100
rect 6048 14066 6604 14100
rect 7066 14066 7622 14100
rect 8084 14066 8640 14100
rect 9102 14066 9658 14100
rect 10120 14066 10676 14100
rect 13742 13832 14298 13866
rect 14760 13832 15316 13866
rect 15778 13832 16334 13866
rect 16796 13832 17352 13866
rect 17814 13832 18370 13866
rect 18832 13832 19388 13866
rect 19850 13832 20406 13866
rect 20868 13832 21424 13866
rect 21886 13832 22442 13866
rect 22904 13832 23460 13866
rect 23922 13832 24478 13866
rect 24940 13832 25496 13866
rect 25958 13832 26514 13866
rect 26976 13832 27532 13866
rect 27994 13832 28550 13866
rect 29012 13832 29568 13866
rect 30030 13832 30586 13866
rect 31048 13832 31604 13866
rect 32066 13832 32622 13866
rect 33084 13832 33640 13866
rect 13742 13724 14298 13758
rect 14760 13724 15316 13758
rect 15778 13724 16334 13758
rect 16796 13724 17352 13758
rect 17814 13724 18370 13758
rect 18832 13724 19388 13758
rect 19850 13724 20406 13758
rect 20868 13724 21424 13758
rect 21886 13724 22442 13758
rect 22904 13724 23460 13758
rect 23922 13724 24478 13758
rect 24940 13724 25496 13758
rect 25958 13724 26514 13758
rect 26976 13724 27532 13758
rect 27994 13724 28550 13758
rect 29012 13724 29568 13758
rect 30030 13724 30586 13758
rect 31048 13724 31604 13758
rect 32066 13724 32622 13758
rect 33084 13724 33640 13758
rect 1976 13356 2532 13390
rect 2994 13356 3550 13390
rect 1976 13248 2532 13282
rect 4012 13356 4568 13390
rect 2994 13248 3550 13282
rect 5030 13356 5586 13390
rect 4012 13248 4568 13282
rect 6048 13356 6604 13390
rect 5030 13248 5586 13282
rect 7066 13356 7622 13390
rect 6048 13248 6604 13282
rect 8084 13356 8640 13390
rect 7066 13248 7622 13282
rect 9102 13356 9658 13390
rect 8084 13248 8640 13282
rect 10120 13356 10676 13390
rect 9102 13248 9658 13282
rect 10120 13248 10676 13282
rect 13742 13014 14298 13048
rect 14760 13014 15316 13048
rect 15778 13014 16334 13048
rect 16796 13014 17352 13048
rect 17814 13014 18370 13048
rect 18832 13014 19388 13048
rect 19850 13014 20406 13048
rect 20868 13014 21424 13048
rect 21886 13014 22442 13048
rect 22904 13014 23460 13048
rect 23922 13014 24478 13048
rect 24940 13014 25496 13048
rect 25958 13014 26514 13048
rect 26976 13014 27532 13048
rect 27994 13014 28550 13048
rect 29012 13014 29568 13048
rect 30030 13014 30586 13048
rect 31048 13014 31604 13048
rect 32066 13014 32622 13048
rect 33084 13014 33640 13048
rect 1976 12538 2532 12572
rect 2994 12538 3550 12572
rect 1976 12430 2532 12464
rect 4012 12538 4568 12572
rect 2994 12430 3550 12464
rect 5030 12538 5586 12572
rect 4012 12430 4568 12464
rect 6048 12538 6604 12572
rect 5030 12430 5586 12464
rect 7066 12538 7622 12572
rect 6048 12430 6604 12464
rect 8084 12538 8640 12572
rect 7066 12430 7622 12464
rect 9102 12538 9658 12572
rect 8084 12430 8640 12464
rect 10120 12538 10676 12572
rect 9102 12430 9658 12464
rect 10120 12430 10676 12464
rect 13742 12346 14298 12380
rect 14760 12346 15316 12380
rect 15778 12346 16334 12380
rect 16796 12346 17352 12380
rect 17814 12346 18370 12380
rect 18832 12346 19388 12380
rect 19850 12346 20406 12380
rect 20868 12346 21424 12380
rect 21886 12346 22442 12380
rect 22904 12346 23460 12380
rect 23922 12346 24478 12380
rect 24940 12346 25496 12380
rect 25958 12346 26514 12380
rect 26976 12346 27532 12380
rect 27994 12346 28550 12380
rect 29012 12346 29568 12380
rect 30030 12346 30586 12380
rect 31048 12346 31604 12380
rect 32066 12346 32622 12380
rect 33084 12346 33640 12380
rect 1976 11720 2532 11754
rect 2994 11720 3550 11754
rect 1976 11612 2532 11646
rect 4012 11720 4568 11754
rect 2994 11612 3550 11646
rect 5030 11720 5586 11754
rect 4012 11612 4568 11646
rect 6048 11720 6604 11754
rect 5030 11612 5586 11646
rect 7066 11720 7622 11754
rect 6048 11612 6604 11646
rect 8084 11720 8640 11754
rect 7066 11612 7622 11646
rect 9102 11720 9658 11754
rect 8084 11612 8640 11646
rect 10120 11720 10676 11754
rect 9102 11612 9658 11646
rect 10120 11612 10676 11646
rect 13742 11636 14298 11670
rect 14760 11636 15316 11670
rect 15778 11636 16334 11670
rect 16796 11636 17352 11670
rect 17814 11636 18370 11670
rect 18832 11636 19388 11670
rect 19850 11636 20406 11670
rect 20868 11636 21424 11670
rect 21886 11636 22442 11670
rect 22904 11636 23460 11670
rect 23922 11636 24478 11670
rect 24940 11636 25496 11670
rect 25958 11636 26514 11670
rect 26976 11636 27532 11670
rect 27994 11636 28550 11670
rect 29012 11636 29568 11670
rect 30030 11636 30586 11670
rect 31048 11636 31604 11670
rect 32066 11636 32622 11670
rect 33084 11636 33640 11670
rect 13742 11114 14298 11148
rect 14760 11114 15316 11148
rect 15778 11114 16334 11148
rect 16796 11114 17352 11148
rect 17814 11114 18370 11148
rect 18832 11114 19388 11148
rect 19850 11114 20406 11148
rect 20868 11114 21424 11148
rect 21886 11114 22442 11148
rect 22904 11114 23460 11148
rect 23922 11114 24478 11148
rect 24940 11114 25496 11148
rect 25958 11114 26514 11148
rect 26976 11114 27532 11148
rect 27994 11114 28550 11148
rect 29012 11114 29568 11148
rect 30030 11114 30586 11148
rect 31048 11114 31604 11148
rect 32066 11114 32622 11148
rect 33084 11114 33640 11148
rect 1976 10902 2532 10936
rect 2994 10902 3550 10936
rect 1976 10794 2532 10828
rect 4012 10902 4568 10936
rect 2994 10794 3550 10828
rect 5030 10902 5586 10936
rect 4012 10794 4568 10828
rect 6048 10902 6604 10936
rect 5030 10794 5586 10828
rect 7066 10902 7622 10936
rect 6048 10794 6604 10828
rect 8084 10902 8640 10936
rect 7066 10794 7622 10828
rect 9102 10902 9658 10936
rect 8084 10794 8640 10828
rect 10120 10902 10676 10936
rect 9102 10794 9658 10828
rect 10120 10794 10676 10828
rect 13742 10404 14298 10438
rect 14760 10404 15316 10438
rect 15778 10404 16334 10438
rect 16796 10404 17352 10438
rect 17814 10404 18370 10438
rect 18832 10404 19388 10438
rect 19850 10404 20406 10438
rect 20868 10404 21424 10438
rect 21886 10404 22442 10438
rect 22904 10404 23460 10438
rect 23922 10404 24478 10438
rect 24940 10404 25496 10438
rect 25958 10404 26514 10438
rect 26976 10404 27532 10438
rect 27994 10404 28550 10438
rect 29012 10404 29568 10438
rect 30030 10404 30586 10438
rect 31048 10404 31604 10438
rect 32066 10404 32622 10438
rect 33084 10404 33640 10438
rect 1976 10084 2532 10118
rect 2994 10084 3550 10118
rect 1976 9976 2532 10010
rect 4012 10084 4568 10118
rect 2994 9976 3550 10010
rect 5030 10084 5586 10118
rect 4012 9976 4568 10010
rect 6048 10084 6604 10118
rect 5030 9976 5586 10010
rect 7066 10084 7622 10118
rect 6048 9976 6604 10010
rect 8084 10084 8640 10118
rect 7066 9976 7622 10010
rect 9102 10084 9658 10118
rect 8084 9976 8640 10010
rect 10120 10084 10676 10118
rect 9102 9976 9658 10010
rect 10120 9976 10676 10010
rect 13740 9880 14296 9914
rect 14758 9880 15314 9914
rect 15776 9880 16332 9914
rect 16794 9880 17350 9914
rect 17812 9880 18368 9914
rect 18830 9880 19386 9914
rect 19848 9880 20404 9914
rect 20866 9880 21422 9914
rect 21884 9880 22440 9914
rect 22902 9880 23458 9914
rect 23920 9880 24476 9914
rect 24938 9880 25494 9914
rect 25956 9880 26512 9914
rect 26974 9880 27530 9914
rect 27992 9880 28548 9914
rect 29010 9880 29566 9914
rect 30028 9880 30584 9914
rect 31046 9880 31602 9914
rect 32064 9880 32620 9914
rect 33082 9880 33638 9914
rect 1976 9266 2532 9300
rect 2994 9266 3550 9300
rect 1976 9158 2532 9192
rect 4012 9266 4568 9300
rect 2994 9158 3550 9192
rect 5030 9266 5586 9300
rect 4012 9158 4568 9192
rect 6048 9266 6604 9300
rect 5030 9158 5586 9192
rect 7066 9266 7622 9300
rect 6048 9158 6604 9192
rect 8084 9266 8640 9300
rect 7066 9158 7622 9192
rect 9102 9266 9658 9300
rect 8084 9158 8640 9192
rect 10120 9266 10676 9300
rect 9102 9158 9658 9192
rect 10120 9158 10676 9192
rect 13740 9170 14296 9204
rect 14758 9170 15314 9204
rect 15776 9170 16332 9204
rect 16794 9170 17350 9204
rect 17812 9170 18368 9204
rect 18830 9170 19386 9204
rect 19848 9170 20404 9204
rect 20866 9170 21422 9204
rect 21884 9170 22440 9204
rect 22902 9170 23458 9204
rect 23920 9170 24476 9204
rect 24938 9170 25494 9204
rect 25956 9170 26512 9204
rect 26974 9170 27530 9204
rect 27992 9170 28548 9204
rect 29010 9170 29566 9204
rect 30028 9170 30584 9204
rect 31046 9170 31602 9204
rect 32064 9170 32620 9204
rect 33082 9170 33638 9204
rect 13740 8646 14296 8680
rect 14758 8646 15314 8680
rect 15776 8646 16332 8680
rect 16794 8646 17350 8680
rect 17812 8646 18368 8680
rect 18830 8646 19386 8680
rect 19848 8646 20404 8680
rect 20866 8646 21422 8680
rect 21884 8646 22440 8680
rect 22902 8646 23458 8680
rect 23920 8646 24476 8680
rect 24938 8646 25494 8680
rect 25956 8646 26512 8680
rect 26974 8646 27530 8680
rect 27992 8646 28548 8680
rect 29010 8646 29566 8680
rect 30028 8646 30584 8680
rect 31046 8646 31602 8680
rect 32064 8646 32620 8680
rect 33082 8646 33638 8680
rect 1976 8448 2532 8482
rect 2994 8448 3550 8482
rect 1976 8340 2532 8374
rect 4012 8448 4568 8482
rect 2994 8340 3550 8374
rect 5030 8448 5586 8482
rect 4012 8340 4568 8374
rect 6048 8448 6604 8482
rect 5030 8340 5586 8374
rect 7066 8448 7622 8482
rect 6048 8340 6604 8374
rect 8084 8448 8640 8482
rect 7066 8340 7622 8374
rect 9102 8448 9658 8482
rect 8084 8340 8640 8374
rect 10120 8448 10676 8482
rect 9102 8340 9658 8374
rect 10120 8340 10676 8374
rect 13740 7936 14296 7970
rect 14758 7936 15314 7970
rect 15776 7936 16332 7970
rect 16794 7936 17350 7970
rect 17812 7936 18368 7970
rect 18830 7936 19386 7970
rect 19848 7936 20404 7970
rect 20866 7936 21422 7970
rect 21884 7936 22440 7970
rect 22902 7936 23458 7970
rect 23920 7936 24476 7970
rect 24938 7936 25494 7970
rect 25956 7936 26512 7970
rect 26974 7936 27530 7970
rect 27992 7936 28548 7970
rect 29010 7936 29566 7970
rect 30028 7936 30584 7970
rect 31046 7936 31602 7970
rect 32064 7936 32620 7970
rect 33082 7936 33638 7970
rect 1976 7630 2532 7664
rect 2994 7630 3550 7664
rect 4012 7630 4568 7664
rect 5030 7630 5586 7664
rect 6048 7630 6604 7664
rect 7066 7630 7622 7664
rect 8084 7630 8640 7664
rect 9102 7630 9658 7664
rect 10120 7630 10676 7664
rect 13740 7414 14296 7448
rect 14758 7414 15314 7448
rect 15776 7414 16332 7448
rect 16794 7414 17350 7448
rect 17812 7414 18368 7448
rect 18830 7414 19386 7448
rect 19848 7414 20404 7448
rect 20866 7414 21422 7448
rect 21884 7414 22440 7448
rect 22902 7414 23458 7448
rect 23920 7414 24476 7448
rect 24938 7414 25494 7448
rect 25956 7414 26512 7448
rect 26974 7414 27530 7448
rect 27992 7414 28548 7448
rect 29010 7414 29566 7448
rect 30028 7414 30584 7448
rect 31046 7414 31602 7448
rect 32064 7414 32620 7448
rect 33082 7414 33638 7448
rect 13740 6704 14296 6738
rect 14758 6704 15314 6738
rect 15776 6704 16332 6738
rect 16794 6704 17350 6738
rect 17812 6704 18368 6738
rect 18830 6704 19386 6738
rect 19848 6704 20404 6738
rect 20866 6704 21422 6738
rect 21884 6704 22440 6738
rect 22902 6704 23458 6738
rect 23920 6704 24476 6738
rect 24938 6704 25494 6738
rect 25956 6704 26512 6738
rect 26974 6704 27530 6738
rect 27992 6704 28548 6738
rect 29010 6704 29566 6738
rect 30028 6704 30584 6738
rect 31046 6704 31602 6738
rect 32064 6704 32620 6738
rect 33082 6704 33638 6738
rect 652 6316 1208 6350
rect 1670 6316 2226 6350
rect 2688 6316 3244 6350
rect 3706 6316 4262 6350
rect 4724 6316 5280 6350
rect 5742 6316 6298 6350
rect 6760 6316 7316 6350
rect 7778 6316 8334 6350
rect 8796 6316 9352 6350
rect 9814 6316 10370 6350
rect 10832 6316 11388 6350
rect 13740 6180 14296 6214
rect 14758 6180 15314 6214
rect 15776 6180 16332 6214
rect 16794 6180 17350 6214
rect 17812 6180 18368 6214
rect 18830 6180 19386 6214
rect 19848 6180 20404 6214
rect 20866 6180 21422 6214
rect 21884 6180 22440 6214
rect 22902 6180 23458 6214
rect 23920 6180 24476 6214
rect 24938 6180 25494 6214
rect 25956 6180 26512 6214
rect 26974 6180 27530 6214
rect 27992 6180 28548 6214
rect 29010 6180 29566 6214
rect 30028 6180 30584 6214
rect 31046 6180 31602 6214
rect 32064 6180 32620 6214
rect 33082 6180 33638 6214
rect 652 5606 1208 5640
rect 1670 5606 2226 5640
rect 2688 5606 3244 5640
rect 3706 5606 4262 5640
rect 4724 5606 5280 5640
rect 5742 5606 6298 5640
rect 6760 5606 7316 5640
rect 7778 5606 8334 5640
rect 8796 5606 9352 5640
rect 9814 5606 10370 5640
rect 10832 5606 11388 5640
rect 13740 5470 14296 5504
rect 14758 5470 15314 5504
rect 15776 5470 16332 5504
rect 16794 5470 17350 5504
rect 17812 5470 18368 5504
rect 18830 5470 19386 5504
rect 19848 5470 20404 5504
rect 20866 5470 21422 5504
rect 21884 5470 22440 5504
rect 22902 5470 23458 5504
rect 23920 5470 24476 5504
rect 24938 5470 25494 5504
rect 25956 5470 26512 5504
rect 26974 5470 27530 5504
rect 27992 5470 28548 5504
rect 29010 5470 29566 5504
rect 30028 5470 30584 5504
rect 31046 5470 31602 5504
rect 32064 5470 32620 5504
rect 33082 5470 33638 5504
rect 652 5204 1208 5238
rect 1670 5204 2226 5238
rect 2688 5204 3244 5238
rect 3706 5204 4262 5238
rect 4724 5204 5280 5238
rect 5742 5204 6298 5238
rect 6760 5204 7316 5238
rect 7778 5204 8334 5238
rect 8796 5204 9352 5238
rect 9814 5204 10370 5238
rect 10832 5204 11388 5238
rect 13740 4946 14296 4980
rect 14758 4946 15314 4980
rect 15776 4946 16332 4980
rect 16794 4946 17350 4980
rect 17812 4946 18368 4980
rect 18830 4946 19386 4980
rect 19848 4946 20404 4980
rect 20866 4946 21422 4980
rect 21884 4946 22440 4980
rect 22902 4946 23458 4980
rect 23920 4946 24476 4980
rect 24938 4946 25494 4980
rect 25956 4946 26512 4980
rect 26974 4946 27530 4980
rect 27992 4946 28548 4980
rect 29010 4946 29566 4980
rect 30028 4946 30584 4980
rect 31046 4946 31602 4980
rect 32064 4946 32620 4980
rect 33082 4946 33638 4980
rect 652 4494 1208 4528
rect 1670 4494 2226 4528
rect 2688 4494 3244 4528
rect 3706 4494 4262 4528
rect 4724 4494 5280 4528
rect 5742 4494 6298 4528
rect 6760 4494 7316 4528
rect 7778 4494 8334 4528
rect 8796 4494 9352 4528
rect 9814 4494 10370 4528
rect 10832 4494 11388 4528
rect 13740 4236 14296 4270
rect 14758 4236 15314 4270
rect 15776 4236 16332 4270
rect 16794 4236 17350 4270
rect 17812 4236 18368 4270
rect 18830 4236 19386 4270
rect 19848 4236 20404 4270
rect 20866 4236 21422 4270
rect 21884 4236 22440 4270
rect 22902 4236 23458 4270
rect 23920 4236 24476 4270
rect 24938 4236 25494 4270
rect 25956 4236 26512 4270
rect 26974 4236 27530 4270
rect 27992 4236 28548 4270
rect 29010 4236 29566 4270
rect 30028 4236 30584 4270
rect 31046 4236 31602 4270
rect 32064 4236 32620 4270
rect 33082 4236 33638 4270
rect 652 4092 1208 4126
rect 1670 4092 2226 4126
rect 2688 4092 3244 4126
rect 3706 4092 4262 4126
rect 4724 4092 5280 4126
rect 5742 4092 6298 4126
rect 6760 4092 7316 4126
rect 7778 4092 8334 4126
rect 8796 4092 9352 4126
rect 9814 4092 10370 4126
rect 10832 4092 11388 4126
rect 13740 3714 14296 3748
rect 14758 3714 15314 3748
rect 15776 3714 16332 3748
rect 16794 3714 17350 3748
rect 17812 3714 18368 3748
rect 18830 3714 19386 3748
rect 19848 3714 20404 3748
rect 20866 3714 21422 3748
rect 21884 3714 22440 3748
rect 22902 3714 23458 3748
rect 23920 3714 24476 3748
rect 24938 3714 25494 3748
rect 25956 3714 26512 3748
rect 26974 3714 27530 3748
rect 27992 3714 28548 3748
rect 29010 3714 29566 3748
rect 30028 3714 30584 3748
rect 31046 3714 31602 3748
rect 32064 3714 32620 3748
rect 33082 3714 33638 3748
rect 652 3382 1208 3416
rect 1670 3382 2226 3416
rect 2688 3382 3244 3416
rect 3706 3382 4262 3416
rect 4724 3382 5280 3416
rect 5742 3382 6298 3416
rect 6760 3382 7316 3416
rect 7778 3382 8334 3416
rect 8796 3382 9352 3416
rect 9814 3382 10370 3416
rect 10832 3382 11388 3416
rect 652 2980 1208 3014
rect 1670 2980 2226 3014
rect 2688 2980 3244 3014
rect 3706 2980 4262 3014
rect 4724 2980 5280 3014
rect 5742 2980 6298 3014
rect 6760 2980 7316 3014
rect 7778 2980 8334 3014
rect 8796 2980 9352 3014
rect 9814 2980 10370 3014
rect 10832 2980 11388 3014
rect 13740 3004 14296 3038
rect 14758 3004 15314 3038
rect 15776 3004 16332 3038
rect 16794 3004 17350 3038
rect 17812 3004 18368 3038
rect 18830 3004 19386 3038
rect 19848 3004 20404 3038
rect 20866 3004 21422 3038
rect 21884 3004 22440 3038
rect 22902 3004 23458 3038
rect 23920 3004 24476 3038
rect 24938 3004 25494 3038
rect 25956 3004 26512 3038
rect 26974 3004 27530 3038
rect 27992 3004 28548 3038
rect 29010 3004 29566 3038
rect 30028 3004 30584 3038
rect 31046 3004 31602 3038
rect 32064 3004 32620 3038
rect 33082 3004 33638 3038
rect 13740 2480 14296 2514
rect 14758 2480 15314 2514
rect 15776 2480 16332 2514
rect 16794 2480 17350 2514
rect 17812 2480 18368 2514
rect 18830 2480 19386 2514
rect 19848 2480 20404 2514
rect 20866 2480 21422 2514
rect 21884 2480 22440 2514
rect 22902 2480 23458 2514
rect 23920 2480 24476 2514
rect 24938 2480 25494 2514
rect 25956 2480 26512 2514
rect 26974 2480 27530 2514
rect 27992 2480 28548 2514
rect 29010 2480 29566 2514
rect 30028 2480 30584 2514
rect 31046 2480 31602 2514
rect 32064 2480 32620 2514
rect 33082 2480 33638 2514
rect 652 2270 1208 2304
rect 1670 2270 2226 2304
rect 2688 2270 3244 2304
rect 3706 2270 4262 2304
rect 4724 2270 5280 2304
rect 5742 2270 6298 2304
rect 6760 2270 7316 2304
rect 7778 2270 8334 2304
rect 8796 2270 9352 2304
rect 9814 2270 10370 2304
rect 10832 2270 11388 2304
rect 13740 1770 14296 1804
rect 14758 1770 15314 1804
rect 15776 1770 16332 1804
rect 16794 1770 17350 1804
rect 17812 1770 18368 1804
rect 18830 1770 19386 1804
rect 19848 1770 20404 1804
rect 20866 1770 21422 1804
rect 21884 1770 22440 1804
rect 22902 1770 23458 1804
rect 23920 1770 24476 1804
rect 24938 1770 25494 1804
rect 25956 1770 26512 1804
rect 26974 1770 27530 1804
rect 27992 1770 28548 1804
rect 29010 1770 29566 1804
rect 30028 1770 30584 1804
rect 31046 1770 31602 1804
rect 32064 1770 32620 1804
rect 33082 1770 33638 1804
rect 1110 1438 1666 1472
rect 2128 1438 2684 1472
rect 3146 1438 3702 1472
rect 4164 1438 4720 1472
rect 5182 1438 5738 1472
rect 6200 1438 6756 1472
rect 7218 1438 7774 1472
rect 8236 1438 8792 1472
rect 9254 1438 9810 1472
rect 10272 1438 10828 1472
rect 13740 1248 14296 1282
rect 14758 1248 15314 1282
rect 15776 1248 16332 1282
rect 16794 1248 17350 1282
rect 17812 1248 18368 1282
rect 18830 1248 19386 1282
rect 19848 1248 20404 1282
rect 20866 1248 21422 1282
rect 21884 1248 22440 1282
rect 22902 1248 23458 1282
rect 23920 1248 24476 1282
rect 24938 1248 25494 1282
rect 25956 1248 26512 1282
rect 26974 1248 27530 1282
rect 27992 1248 28548 1282
rect 29010 1248 29566 1282
rect 30028 1248 30584 1282
rect 31046 1248 31602 1282
rect 32064 1248 32620 1282
rect 33082 1248 33638 1282
rect 1110 728 1666 762
rect 2128 728 2684 762
rect 3146 728 3702 762
rect 4164 728 4720 762
rect 5182 728 5738 762
rect 6200 728 6756 762
rect 7218 728 7774 762
rect 8236 728 8792 762
rect 9254 728 9810 762
rect 10272 728 10828 762
rect 13740 538 14296 572
rect 14758 538 15314 572
rect 15776 538 16332 572
rect 16794 538 17350 572
rect 17812 538 18368 572
rect 18830 538 19386 572
rect 19848 538 20404 572
rect 20866 538 21422 572
rect 21884 538 22440 572
rect 22902 538 23458 572
rect 23920 538 24476 572
rect 24938 538 25494 572
rect 25956 538 26512 572
rect 26974 538 27530 572
rect 27992 538 28548 572
rect 29010 538 29566 572
rect 30028 538 30584 572
rect 31046 538 31602 572
rect 32064 538 32620 572
rect 33082 538 33638 572
<< locali >>
rect 11290 30700 11390 30862
rect 35634 30700 35734 30862
rect 17880 28318 17970 28348
rect 17880 28284 17908 28318
rect 17942 28284 17970 28318
rect 17880 28256 17970 28284
rect 18898 28318 18988 28348
rect 18898 28284 18926 28318
rect 18960 28284 18988 28318
rect 18898 28256 18988 28284
rect 19916 28318 20006 28348
rect 19916 28284 19944 28318
rect 19978 28284 20006 28318
rect 19916 28256 20006 28284
rect 20934 28318 21024 28348
rect 20934 28284 20962 28318
rect 20996 28284 21024 28318
rect 20934 28256 21024 28284
rect 21952 28318 22042 28348
rect 21952 28284 21980 28318
rect 22014 28284 22042 28318
rect 21952 28256 22042 28284
rect 22970 28318 23060 28348
rect 22970 28284 22998 28318
rect 23032 28284 23060 28318
rect 22970 28256 23060 28284
rect 23988 28318 24078 28348
rect 23988 28284 24016 28318
rect 24050 28284 24078 28318
rect 23988 28256 24078 28284
rect 25006 28318 25096 28348
rect 25006 28284 25034 28318
rect 25068 28284 25096 28318
rect 25006 28256 25096 28284
rect 26024 28318 26114 28348
rect 26024 28284 26052 28318
rect 26086 28284 26114 28318
rect 26024 28256 26114 28284
rect 27042 28318 27132 28348
rect 27042 28284 27070 28318
rect 27104 28284 27132 28318
rect 27042 28256 27132 28284
rect 28060 28318 28150 28348
rect 28060 28284 28088 28318
rect 28122 28284 28150 28318
rect 28060 28256 28150 28284
rect 29078 28318 29168 28348
rect 29078 28284 29106 28318
rect 29140 28284 29168 28318
rect 29078 28256 29168 28284
rect 30096 28318 30186 28348
rect 30096 28284 30124 28318
rect 30158 28284 30186 28318
rect 30096 28256 30186 28284
rect 31114 28318 31204 28348
rect 31114 28284 31142 28318
rect 31176 28284 31204 28318
rect 31114 28256 31204 28284
rect 32132 28318 32222 28348
rect 32132 28284 32160 28318
rect 32194 28284 32222 28318
rect 32132 28256 32222 28284
rect 33150 28318 33240 28348
rect 33150 28284 33178 28318
rect 33212 28284 33240 28318
rect 33150 28256 33240 28284
rect 17632 28061 17648 28095
rect 18204 28061 18220 28095
rect 18650 28061 18666 28095
rect 19222 28061 19238 28095
rect 19668 28061 19684 28095
rect 20240 28061 20256 28095
rect 20686 28061 20702 28095
rect 21258 28061 21274 28095
rect 21704 28061 21720 28095
rect 22276 28061 22292 28095
rect 22722 28061 22738 28095
rect 23294 28061 23310 28095
rect 23740 28061 23756 28095
rect 24312 28061 24328 28095
rect 24758 28061 24774 28095
rect 25330 28061 25346 28095
rect 25776 28061 25792 28095
rect 26348 28061 26364 28095
rect 26794 28061 26810 28095
rect 27366 28061 27382 28095
rect 27812 28061 27828 28095
rect 28384 28061 28400 28095
rect 28830 28061 28846 28095
rect 29402 28061 29418 28095
rect 29848 28061 29864 28095
rect 30420 28061 30436 28095
rect 30866 28061 30882 28095
rect 31438 28061 31454 28095
rect 31884 28061 31900 28095
rect 32456 28061 32472 28095
rect 32902 28061 32918 28095
rect 33474 28061 33490 28095
rect 17400 28002 17434 28018
rect 17400 27410 17434 27426
rect 18418 28002 18452 28018
rect 18418 27410 18452 27426
rect 19436 28002 19470 28018
rect 19436 27410 19470 27426
rect 20454 28002 20488 28018
rect 20454 27410 20488 27426
rect 21472 28002 21506 28018
rect 21472 27410 21506 27426
rect 22490 28002 22524 28018
rect 22490 27410 22524 27426
rect 23508 28002 23542 28018
rect 23508 27410 23542 27426
rect 24526 28002 24560 28018
rect 24526 27410 24560 27426
rect 25544 28002 25578 28018
rect 25544 27410 25578 27426
rect 26562 28002 26596 28018
rect 26562 27410 26596 27426
rect 27580 28002 27614 28018
rect 27580 27410 27614 27426
rect 28598 28002 28632 28018
rect 28598 27410 28632 27426
rect 29616 28002 29650 28018
rect 29616 27410 29650 27426
rect 30634 28002 30668 28018
rect 30634 27410 30668 27426
rect 31652 28002 31686 28018
rect 31652 27410 31686 27426
rect 32670 28002 32704 28018
rect 32670 27410 32704 27426
rect 33688 28002 33722 28018
rect 33688 27410 33722 27426
rect 17632 27333 17648 27367
rect 18204 27333 18220 27367
rect 18650 27333 18666 27367
rect 19222 27333 19238 27367
rect 19668 27333 19684 27367
rect 20240 27333 20256 27367
rect 20686 27333 20702 27367
rect 21258 27333 21274 27367
rect 21704 27333 21720 27367
rect 22276 27333 22292 27367
rect 22722 27333 22738 27367
rect 23294 27333 23310 27367
rect 23740 27333 23756 27367
rect 24312 27333 24328 27367
rect 24758 27333 24774 27367
rect 25330 27333 25346 27367
rect 25776 27333 25792 27367
rect 26348 27333 26364 27367
rect 26794 27333 26810 27367
rect 27366 27333 27382 27367
rect 27812 27333 27828 27367
rect 28384 27333 28400 27367
rect 28830 27333 28846 27367
rect 29402 27333 29418 27367
rect 29848 27333 29864 27367
rect 30420 27333 30436 27367
rect 30866 27333 30882 27367
rect 31438 27333 31454 27367
rect 31884 27333 31900 27367
rect 32456 27333 32472 27367
rect 32902 27333 32918 27367
rect 33474 27333 33490 27367
rect 17902 27164 17992 27194
rect 17902 27130 17930 27164
rect 17964 27130 17992 27164
rect 17902 27102 17992 27130
rect 18920 27164 19010 27194
rect 18920 27130 18948 27164
rect 18982 27130 19010 27164
rect 18920 27102 19010 27130
rect 19938 27164 20028 27194
rect 19938 27130 19966 27164
rect 20000 27130 20028 27164
rect 19938 27102 20028 27130
rect 20956 27164 21046 27194
rect 20956 27130 20984 27164
rect 21018 27130 21046 27164
rect 20956 27102 21046 27130
rect 21974 27164 22064 27194
rect 21974 27130 22002 27164
rect 22036 27130 22064 27164
rect 21974 27102 22064 27130
rect 22992 27164 23082 27194
rect 22992 27130 23020 27164
rect 23054 27130 23082 27164
rect 22992 27102 23082 27130
rect 24010 27164 24100 27194
rect 24010 27130 24038 27164
rect 24072 27130 24100 27164
rect 24010 27102 24100 27130
rect 25028 27164 25118 27194
rect 25028 27130 25056 27164
rect 25090 27130 25118 27164
rect 25028 27102 25118 27130
rect 26046 27164 26136 27194
rect 26046 27130 26074 27164
rect 26108 27130 26136 27164
rect 26046 27102 26136 27130
rect 27064 27164 27154 27194
rect 27064 27130 27092 27164
rect 27126 27130 27154 27164
rect 27064 27102 27154 27130
rect 28082 27164 28172 27194
rect 28082 27130 28110 27164
rect 28144 27130 28172 27164
rect 28082 27102 28172 27130
rect 29100 27164 29190 27194
rect 29100 27130 29128 27164
rect 29162 27130 29190 27164
rect 29100 27102 29190 27130
rect 30118 27164 30208 27194
rect 30118 27130 30146 27164
rect 30180 27130 30208 27164
rect 30118 27102 30208 27130
rect 31136 27164 31226 27194
rect 31136 27130 31164 27164
rect 31198 27130 31226 27164
rect 31136 27102 31226 27130
rect 32154 27164 32244 27194
rect 32154 27130 32182 27164
rect 32216 27130 32244 27164
rect 32154 27102 32244 27130
rect 33172 27164 33262 27194
rect 33172 27130 33200 27164
rect 33234 27130 33262 27164
rect 33172 27102 33262 27130
rect 17632 26925 17648 26959
rect 18204 26925 18220 26959
rect 18650 26925 18666 26959
rect 19222 26925 19238 26959
rect 19668 26925 19684 26959
rect 20240 26925 20256 26959
rect 20686 26925 20702 26959
rect 21258 26925 21274 26959
rect 21704 26925 21720 26959
rect 22276 26925 22292 26959
rect 22722 26925 22738 26959
rect 23294 26925 23310 26959
rect 23740 26925 23756 26959
rect 24312 26925 24328 26959
rect 24758 26925 24774 26959
rect 25330 26925 25346 26959
rect 25776 26925 25792 26959
rect 26348 26925 26364 26959
rect 26794 26925 26810 26959
rect 27366 26925 27382 26959
rect 27812 26925 27828 26959
rect 28384 26925 28400 26959
rect 28830 26925 28846 26959
rect 29402 26925 29418 26959
rect 29848 26925 29864 26959
rect 30420 26925 30436 26959
rect 30866 26925 30882 26959
rect 31438 26925 31454 26959
rect 31884 26925 31900 26959
rect 32456 26925 32472 26959
rect 32902 26925 32918 26959
rect 33474 26925 33490 26959
rect 17400 26866 17434 26882
rect 17400 26274 17434 26290
rect 18418 26866 18452 26882
rect 18418 26274 18452 26290
rect 19436 26866 19470 26882
rect 19436 26274 19470 26290
rect 20454 26866 20488 26882
rect 20454 26274 20488 26290
rect 21472 26866 21506 26882
rect 21472 26274 21506 26290
rect 22490 26866 22524 26882
rect 22490 26274 22524 26290
rect 23508 26866 23542 26882
rect 23508 26274 23542 26290
rect 24526 26866 24560 26882
rect 24526 26274 24560 26290
rect 25544 26866 25578 26882
rect 25544 26274 25578 26290
rect 26562 26866 26596 26882
rect 26562 26274 26596 26290
rect 27580 26866 27614 26882
rect 27580 26274 27614 26290
rect 28598 26866 28632 26882
rect 28598 26274 28632 26290
rect 29616 26866 29650 26882
rect 29616 26274 29650 26290
rect 30634 26866 30668 26882
rect 30634 26274 30668 26290
rect 31652 26866 31686 26882
rect 31652 26274 31686 26290
rect 32670 26866 32704 26882
rect 32670 26274 32704 26290
rect 33688 26866 33722 26882
rect 33688 26274 33722 26290
rect 17632 26197 17648 26231
rect 18204 26197 18220 26231
rect 18650 26197 18666 26231
rect 19222 26197 19238 26231
rect 19668 26197 19684 26231
rect 20240 26197 20256 26231
rect 20686 26197 20702 26231
rect 21258 26197 21274 26231
rect 21704 26197 21720 26231
rect 22276 26197 22292 26231
rect 22722 26197 22738 26231
rect 23294 26197 23310 26231
rect 23740 26197 23756 26231
rect 24312 26197 24328 26231
rect 24758 26197 24774 26231
rect 25330 26197 25346 26231
rect 25776 26197 25792 26231
rect 26348 26197 26364 26231
rect 26794 26197 26810 26231
rect 27366 26197 27382 26231
rect 27812 26197 27828 26231
rect 28384 26197 28400 26231
rect 28830 26197 28846 26231
rect 29402 26197 29418 26231
rect 29848 26197 29864 26231
rect 30420 26197 30436 26231
rect 30866 26197 30882 26231
rect 31438 26197 31454 26231
rect 31884 26197 31900 26231
rect 32456 26197 32472 26231
rect 32902 26197 32918 26231
rect 33474 26197 33490 26231
rect 17880 26032 17970 26062
rect 17880 25998 17908 26032
rect 17942 25998 17970 26032
rect 17880 25970 17970 25998
rect 18898 26032 18988 26062
rect 18898 25998 18926 26032
rect 18960 25998 18988 26032
rect 18898 25970 18988 25998
rect 19916 26032 20006 26062
rect 19916 25998 19944 26032
rect 19978 25998 20006 26032
rect 19916 25970 20006 25998
rect 20934 26032 21024 26062
rect 20934 25998 20962 26032
rect 20996 25998 21024 26032
rect 20934 25970 21024 25998
rect 21952 26032 22042 26062
rect 21952 25998 21980 26032
rect 22014 25998 22042 26032
rect 21952 25970 22042 25998
rect 22970 26032 23060 26062
rect 22970 25998 22998 26032
rect 23032 25998 23060 26032
rect 22970 25970 23060 25998
rect 23988 26032 24078 26062
rect 23988 25998 24016 26032
rect 24050 25998 24078 26032
rect 23988 25970 24078 25998
rect 25006 26032 25096 26062
rect 25006 25998 25034 26032
rect 25068 25998 25096 26032
rect 25006 25970 25096 25998
rect 26024 26032 26114 26062
rect 26024 25998 26052 26032
rect 26086 25998 26114 26032
rect 26024 25970 26114 25998
rect 27042 26032 27132 26062
rect 27042 25998 27070 26032
rect 27104 25998 27132 26032
rect 27042 25970 27132 25998
rect 28060 26032 28150 26062
rect 28060 25998 28088 26032
rect 28122 25998 28150 26032
rect 28060 25970 28150 25998
rect 29078 26032 29168 26062
rect 29078 25998 29106 26032
rect 29140 25998 29168 26032
rect 29078 25970 29168 25998
rect 30096 26032 30186 26062
rect 30096 25998 30124 26032
rect 30158 25998 30186 26032
rect 30096 25970 30186 25998
rect 31114 26032 31204 26062
rect 31114 25998 31142 26032
rect 31176 25998 31204 26032
rect 31114 25970 31204 25998
rect 32132 26032 32222 26062
rect 32132 25998 32160 26032
rect 32194 25998 32222 26032
rect 32132 25970 32222 25998
rect 33150 26032 33240 26062
rect 33150 25998 33178 26032
rect 33212 25998 33240 26032
rect 33150 25970 33240 25998
rect 17632 25789 17648 25823
rect 18204 25789 18220 25823
rect 18650 25789 18666 25823
rect 19222 25789 19238 25823
rect 19668 25789 19684 25823
rect 20240 25789 20256 25823
rect 20686 25789 20702 25823
rect 21258 25789 21274 25823
rect 21704 25789 21720 25823
rect 22276 25789 22292 25823
rect 22722 25789 22738 25823
rect 23294 25789 23310 25823
rect 23740 25789 23756 25823
rect 24312 25789 24328 25823
rect 24758 25789 24774 25823
rect 25330 25789 25346 25823
rect 25776 25789 25792 25823
rect 26348 25789 26364 25823
rect 26794 25789 26810 25823
rect 27366 25789 27382 25823
rect 27812 25789 27828 25823
rect 28384 25789 28400 25823
rect 28830 25789 28846 25823
rect 29402 25789 29418 25823
rect 29848 25789 29864 25823
rect 30420 25789 30436 25823
rect 30866 25789 30882 25823
rect 31438 25789 31454 25823
rect 31884 25789 31900 25823
rect 32456 25789 32472 25823
rect 32902 25789 32918 25823
rect 33474 25789 33490 25823
rect 17400 25730 17434 25746
rect 17400 25138 17434 25154
rect 18418 25730 18452 25746
rect 18418 25138 18452 25154
rect 19436 25730 19470 25746
rect 19436 25138 19470 25154
rect 20454 25730 20488 25746
rect 20454 25138 20488 25154
rect 21472 25730 21506 25746
rect 21472 25138 21506 25154
rect 22490 25730 22524 25746
rect 22490 25138 22524 25154
rect 23508 25730 23542 25746
rect 23508 25138 23542 25154
rect 24526 25730 24560 25746
rect 24526 25138 24560 25154
rect 25544 25730 25578 25746
rect 25544 25138 25578 25154
rect 26562 25730 26596 25746
rect 26562 25138 26596 25154
rect 27580 25730 27614 25746
rect 27580 25138 27614 25154
rect 28598 25730 28632 25746
rect 28598 25138 28632 25154
rect 29616 25730 29650 25746
rect 29616 25138 29650 25154
rect 30634 25730 30668 25746
rect 30634 25138 30668 25154
rect 31652 25730 31686 25746
rect 31652 25138 31686 25154
rect 32670 25730 32704 25746
rect 32670 25138 32704 25154
rect 33688 25730 33722 25746
rect 33688 25138 33722 25154
rect 17632 25061 17648 25095
rect 18204 25061 18220 25095
rect 18650 25061 18666 25095
rect 19222 25061 19238 25095
rect 19668 25061 19684 25095
rect 20240 25061 20256 25095
rect 20686 25061 20702 25095
rect 21258 25061 21274 25095
rect 21704 25061 21720 25095
rect 22276 25061 22292 25095
rect 22722 25061 22738 25095
rect 23294 25061 23310 25095
rect 23740 25061 23756 25095
rect 24312 25061 24328 25095
rect 24758 25061 24774 25095
rect 25330 25061 25346 25095
rect 25776 25061 25792 25095
rect 26348 25061 26364 25095
rect 26794 25061 26810 25095
rect 27366 25061 27382 25095
rect 27812 25061 27828 25095
rect 28384 25061 28400 25095
rect 28830 25061 28846 25095
rect 29402 25061 29418 25095
rect 29848 25061 29864 25095
rect 30420 25061 30436 25095
rect 30866 25061 30882 25095
rect 31438 25061 31454 25095
rect 31884 25061 31900 25095
rect 32456 25061 32472 25095
rect 32902 25061 32918 25095
rect 33474 25061 33490 25095
rect 17880 24650 17970 24680
rect 17880 24616 17908 24650
rect 17942 24616 17970 24650
rect 17880 24588 17970 24616
rect 18898 24650 18988 24680
rect 18898 24616 18926 24650
rect 18960 24616 18988 24650
rect 18898 24588 18988 24616
rect 19916 24650 20006 24680
rect 19916 24616 19944 24650
rect 19978 24616 20006 24650
rect 19916 24588 20006 24616
rect 20934 24650 21024 24680
rect 20934 24616 20962 24650
rect 20996 24616 21024 24650
rect 20934 24588 21024 24616
rect 21952 24650 22042 24680
rect 21952 24616 21980 24650
rect 22014 24616 22042 24650
rect 21952 24588 22042 24616
rect 22970 24650 23060 24680
rect 22970 24616 22998 24650
rect 23032 24616 23060 24650
rect 22970 24588 23060 24616
rect 23988 24650 24078 24680
rect 23988 24616 24016 24650
rect 24050 24616 24078 24650
rect 23988 24588 24078 24616
rect 25006 24650 25096 24680
rect 25006 24616 25034 24650
rect 25068 24616 25096 24650
rect 25006 24588 25096 24616
rect 26024 24650 26114 24680
rect 26024 24616 26052 24650
rect 26086 24616 26114 24650
rect 26024 24588 26114 24616
rect 27042 24650 27132 24680
rect 27042 24616 27070 24650
rect 27104 24616 27132 24650
rect 27042 24588 27132 24616
rect 28060 24650 28150 24680
rect 28060 24616 28088 24650
rect 28122 24616 28150 24650
rect 28060 24588 28150 24616
rect 29078 24650 29168 24680
rect 29078 24616 29106 24650
rect 29140 24616 29168 24650
rect 29078 24588 29168 24616
rect 30096 24650 30186 24680
rect 30096 24616 30124 24650
rect 30158 24616 30186 24650
rect 30096 24588 30186 24616
rect 31114 24650 31204 24680
rect 31114 24616 31142 24650
rect 31176 24616 31204 24650
rect 31114 24588 31204 24616
rect 32132 24650 32222 24680
rect 32132 24616 32160 24650
rect 32194 24616 32222 24650
rect 32132 24588 32222 24616
rect 33150 24650 33240 24680
rect 33150 24616 33178 24650
rect 33212 24616 33240 24650
rect 33150 24588 33240 24616
rect 18826 24151 18842 24185
rect 19398 24151 19414 24185
rect 19844 24151 19860 24185
rect 20416 24151 20432 24185
rect 20862 24151 20878 24185
rect 21434 24151 21450 24185
rect 21880 24151 21896 24185
rect 22452 24151 22468 24185
rect 22898 24151 22914 24185
rect 23470 24151 23486 24185
rect 23916 24151 23932 24185
rect 24488 24151 24504 24185
rect 24934 24151 24950 24185
rect 25506 24151 25522 24185
rect 25952 24151 25968 24185
rect 26524 24151 26540 24185
rect 26970 24151 26986 24185
rect 27542 24151 27558 24185
rect 27988 24151 28004 24185
rect 28560 24151 28576 24185
rect 29006 24151 29022 24185
rect 29578 24151 29594 24185
rect 30024 24151 30040 24185
rect 30596 24151 30612 24185
rect 31042 24151 31058 24185
rect 31614 24151 31630 24185
rect 32060 24151 32076 24185
rect 32632 24151 32648 24185
rect 18594 24092 18628 24108
rect 18594 23500 18628 23516
rect 19612 24092 19646 24108
rect 19612 23500 19646 23516
rect 20630 24092 20664 24108
rect 20630 23500 20664 23516
rect 21648 24092 21682 24108
rect 21648 23500 21682 23516
rect 22666 24092 22700 24108
rect 22666 23500 22700 23516
rect 23684 24092 23718 24108
rect 23684 23500 23718 23516
rect 24702 24092 24736 24108
rect 24702 23500 24736 23516
rect 25720 24092 25754 24108
rect 25720 23500 25754 23516
rect 26738 24092 26772 24108
rect 26738 23500 26772 23516
rect 27756 24092 27790 24108
rect 27756 23500 27790 23516
rect 28774 24092 28808 24108
rect 28774 23500 28808 23516
rect 29792 24092 29826 24108
rect 29792 23500 29826 23516
rect 30810 24092 30844 24108
rect 30810 23500 30844 23516
rect 31828 24092 31862 24108
rect 31828 23500 31862 23516
rect 32846 24092 32880 24108
rect 32846 23500 32880 23516
rect 18826 23423 18842 23457
rect 19398 23423 19414 23457
rect 19844 23423 19860 23457
rect 20416 23423 20432 23457
rect 20862 23423 20878 23457
rect 21434 23423 21450 23457
rect 21880 23423 21896 23457
rect 22452 23423 22468 23457
rect 22898 23423 22914 23457
rect 23470 23423 23486 23457
rect 23916 23423 23932 23457
rect 24488 23423 24504 23457
rect 24934 23423 24950 23457
rect 25506 23423 25522 23457
rect 25952 23423 25968 23457
rect 26524 23423 26540 23457
rect 26970 23423 26986 23457
rect 27542 23423 27558 23457
rect 27988 23423 28004 23457
rect 28560 23423 28576 23457
rect 29006 23423 29022 23457
rect 29578 23423 29594 23457
rect 30024 23423 30040 23457
rect 30596 23423 30612 23457
rect 31042 23423 31058 23457
rect 31614 23423 31630 23457
rect 32060 23423 32076 23457
rect 32632 23423 32648 23457
rect 18568 23302 18658 23332
rect 18568 23268 18596 23302
rect 18630 23268 18658 23302
rect 18568 23240 18658 23268
rect 19586 23302 19676 23332
rect 19586 23268 19614 23302
rect 19648 23268 19676 23302
rect 19586 23240 19676 23268
rect 20604 23302 20694 23332
rect 20604 23268 20632 23302
rect 20666 23268 20694 23302
rect 20604 23240 20694 23268
rect 21622 23302 21712 23332
rect 21622 23268 21650 23302
rect 21684 23268 21712 23302
rect 21622 23240 21712 23268
rect 22640 23302 22730 23332
rect 22640 23268 22668 23302
rect 22702 23268 22730 23302
rect 22640 23240 22730 23268
rect 23658 23302 23748 23332
rect 23658 23268 23686 23302
rect 23720 23268 23748 23302
rect 23658 23240 23748 23268
rect 24676 23302 24766 23332
rect 24676 23268 24704 23302
rect 24738 23268 24766 23302
rect 24676 23240 24766 23268
rect 25694 23302 25784 23332
rect 25694 23268 25722 23302
rect 25756 23268 25784 23302
rect 25694 23240 25784 23268
rect 26712 23302 26802 23332
rect 26712 23268 26740 23302
rect 26774 23268 26802 23302
rect 26712 23240 26802 23268
rect 27730 23302 27820 23332
rect 27730 23268 27758 23302
rect 27792 23268 27820 23302
rect 27730 23240 27820 23268
rect 28748 23302 28838 23332
rect 28748 23268 28776 23302
rect 28810 23268 28838 23302
rect 28748 23240 28838 23268
rect 29766 23302 29856 23332
rect 29766 23268 29794 23302
rect 29828 23268 29856 23302
rect 29766 23240 29856 23268
rect 30784 23302 30874 23332
rect 30784 23268 30812 23302
rect 30846 23268 30874 23302
rect 30784 23240 30874 23268
rect 31802 23302 31892 23332
rect 31802 23268 31830 23302
rect 31864 23268 31892 23302
rect 31802 23240 31892 23268
rect 32820 23302 32910 23332
rect 32820 23268 32848 23302
rect 32882 23268 32910 23302
rect 32820 23240 32910 23268
rect 18826 23119 18842 23153
rect 19398 23119 19414 23153
rect 19844 23119 19860 23153
rect 20416 23119 20432 23153
rect 20862 23119 20878 23153
rect 21434 23119 21450 23153
rect 21880 23119 21896 23153
rect 22452 23119 22468 23153
rect 22898 23119 22914 23153
rect 23470 23119 23486 23153
rect 23916 23119 23932 23153
rect 24488 23119 24504 23153
rect 24934 23119 24950 23153
rect 25506 23119 25522 23153
rect 25952 23119 25968 23153
rect 26524 23119 26540 23153
rect 26970 23119 26986 23153
rect 27542 23119 27558 23153
rect 27988 23119 28004 23153
rect 28560 23119 28576 23153
rect 29006 23119 29022 23153
rect 29578 23119 29594 23153
rect 30024 23119 30040 23153
rect 30596 23119 30612 23153
rect 31042 23119 31058 23153
rect 31614 23119 31630 23153
rect 32060 23119 32076 23153
rect 32632 23119 32648 23153
rect 18594 23060 18628 23076
rect 18594 22468 18628 22484
rect 19612 23060 19646 23076
rect 19612 22468 19646 22484
rect 20630 23060 20664 23076
rect 20630 22468 20664 22484
rect 21648 23060 21682 23076
rect 21648 22468 21682 22484
rect 22666 23060 22700 23076
rect 22666 22468 22700 22484
rect 23684 23060 23718 23076
rect 23684 22468 23718 22484
rect 24702 23060 24736 23076
rect 24702 22468 24736 22484
rect 25720 23060 25754 23076
rect 25720 22468 25754 22484
rect 26738 23060 26772 23076
rect 26738 22468 26772 22484
rect 27756 23060 27790 23076
rect 27756 22468 27790 22484
rect 28774 23060 28808 23076
rect 28774 22468 28808 22484
rect 29792 23060 29826 23076
rect 29792 22468 29826 22484
rect 30810 23060 30844 23076
rect 30810 22468 30844 22484
rect 31828 23060 31862 23076
rect 31828 22468 31862 22484
rect 32846 23060 32880 23076
rect 32846 22468 32880 22484
rect 18826 22391 18842 22425
rect 19398 22391 19414 22425
rect 19844 22391 19860 22425
rect 20416 22391 20432 22425
rect 20862 22391 20878 22425
rect 21434 22391 21450 22425
rect 21880 22391 21896 22425
rect 22452 22391 22468 22425
rect 22898 22391 22914 22425
rect 23470 22391 23486 22425
rect 23916 22391 23932 22425
rect 24488 22391 24504 22425
rect 24934 22391 24950 22425
rect 25506 22391 25522 22425
rect 25952 22391 25968 22425
rect 26524 22391 26540 22425
rect 26970 22391 26986 22425
rect 27542 22391 27558 22425
rect 27988 22391 28004 22425
rect 28560 22391 28576 22425
rect 29006 22391 29022 22425
rect 29578 22391 29594 22425
rect 30024 22391 30040 22425
rect 30596 22391 30612 22425
rect 31042 22391 31058 22425
rect 31614 22391 31630 22425
rect 32060 22391 32076 22425
rect 32632 22391 32648 22425
rect 18174 22024 18264 22054
rect 18174 21990 18202 22024
rect 18236 21990 18264 22024
rect 18174 21962 18264 21990
rect 19192 22024 19282 22054
rect 19192 21990 19220 22024
rect 19254 21990 19282 22024
rect 19192 21962 19282 21990
rect 20210 22024 20300 22054
rect 20210 21990 20238 22024
rect 20272 21990 20300 22024
rect 20210 21962 20300 21990
rect 21228 22024 21318 22054
rect 21228 21990 21256 22024
rect 21290 21990 21318 22024
rect 21228 21962 21318 21990
rect 22246 22024 22336 22054
rect 22246 21990 22274 22024
rect 22308 21990 22336 22024
rect 22246 21962 22336 21990
rect 23264 22024 23354 22054
rect 23264 21990 23292 22024
rect 23326 21990 23354 22024
rect 23264 21962 23354 21990
rect 24282 22024 24372 22054
rect 24282 21990 24310 22024
rect 24344 21990 24372 22024
rect 24282 21962 24372 21990
rect 25300 22024 25390 22054
rect 25300 21990 25328 22024
rect 25362 21990 25390 22024
rect 25300 21962 25390 21990
rect 26318 22024 26408 22054
rect 26318 21990 26346 22024
rect 26380 21990 26408 22024
rect 26318 21962 26408 21990
rect 27336 22024 27426 22054
rect 27336 21990 27364 22024
rect 27398 21990 27426 22024
rect 27336 21962 27426 21990
rect 28354 22024 28444 22054
rect 28354 21990 28382 22024
rect 28416 21990 28444 22024
rect 28354 21962 28444 21990
rect 29372 22024 29462 22054
rect 29372 21990 29400 22024
rect 29434 21990 29462 22024
rect 29372 21962 29462 21990
rect 30390 22024 30480 22054
rect 30390 21990 30418 22024
rect 30452 21990 30480 22024
rect 30390 21962 30480 21990
rect 31408 22024 31498 22054
rect 31408 21990 31436 22024
rect 31470 21990 31498 22024
rect 31408 21962 31498 21990
rect 32426 22024 32516 22054
rect 32426 21990 32454 22024
rect 32488 21990 32516 22024
rect 32426 21962 32516 21990
rect 33444 22024 33534 22054
rect 33444 21990 33472 22024
rect 33506 21990 33534 22024
rect 33444 21962 33534 21990
rect 13576 21714 13666 21744
rect 13576 21680 13604 21714
rect 13638 21680 13666 21714
rect 13576 21652 13666 21680
rect 14594 21714 14684 21744
rect 14594 21680 14622 21714
rect 14656 21680 14684 21714
rect 14594 21652 14684 21680
rect 15612 21714 15702 21744
rect 15612 21680 15640 21714
rect 15674 21680 15702 21714
rect 15612 21652 15702 21680
rect 16630 21714 16720 21744
rect 16630 21680 16658 21714
rect 16692 21680 16720 21714
rect 16630 21652 16720 21680
rect 18618 21515 18634 21549
rect 19190 21515 19206 21549
rect 19636 21515 19652 21549
rect 20208 21515 20224 21549
rect 20654 21515 20670 21549
rect 21226 21515 21242 21549
rect 21672 21515 21688 21549
rect 22244 21515 22260 21549
rect 22690 21515 22706 21549
rect 23262 21515 23278 21549
rect 23708 21515 23724 21549
rect 24280 21515 24296 21549
rect 24726 21515 24742 21549
rect 25298 21515 25314 21549
rect 25744 21515 25760 21549
rect 26316 21515 26332 21549
rect 26762 21515 26778 21549
rect 27334 21515 27350 21549
rect 27780 21515 27796 21549
rect 28352 21515 28368 21549
rect 28798 21515 28814 21549
rect 29370 21515 29386 21549
rect 29816 21515 29832 21549
rect 30388 21515 30404 21549
rect 30834 21515 30850 21549
rect 31406 21515 31422 21549
rect 31852 21515 31868 21549
rect 32424 21515 32440 21549
rect 32870 21515 32886 21549
rect 33442 21515 33458 21549
rect 18386 21456 18420 21472
rect 13314 21411 13330 21445
rect 13886 21411 13902 21445
rect 14332 21411 14348 21445
rect 14904 21411 14920 21445
rect 15350 21411 15366 21445
rect 15922 21411 15938 21445
rect 16368 21411 16384 21445
rect 16940 21411 16956 21445
rect 13082 21352 13116 21368
rect 13082 20760 13116 20776
rect 14100 21352 14134 21368
rect 14100 20760 14134 20776
rect 15118 21352 15152 21368
rect 15118 20760 15152 20776
rect 16136 21352 16170 21368
rect 16136 20760 16170 20776
rect 17154 21352 17188 21368
rect 18386 20864 18420 20880
rect 19404 21456 19438 21472
rect 19404 20864 19438 20880
rect 20422 21456 20456 21472
rect 20422 20864 20456 20880
rect 21440 21456 21474 21472
rect 21440 20864 21474 20880
rect 22458 21456 22492 21472
rect 22458 20864 22492 20880
rect 23476 21456 23510 21472
rect 23476 20864 23510 20880
rect 24494 21456 24528 21472
rect 24494 20864 24528 20880
rect 25512 21456 25546 21472
rect 25512 20864 25546 20880
rect 26530 21456 26564 21472
rect 26530 20864 26564 20880
rect 27548 21456 27582 21472
rect 27548 20864 27582 20880
rect 28566 21456 28600 21472
rect 28566 20864 28600 20880
rect 29584 21456 29618 21472
rect 29584 20864 29618 20880
rect 30602 21456 30636 21472
rect 30602 20864 30636 20880
rect 31620 21456 31654 21472
rect 31620 20864 31654 20880
rect 32638 21456 32672 21472
rect 32638 20864 32672 20880
rect 33656 21456 33690 21472
rect 33656 20864 33690 20880
rect 18618 20787 18634 20821
rect 19190 20787 19206 20821
rect 19636 20787 19652 20821
rect 20208 20787 20224 20821
rect 20654 20787 20670 20821
rect 21226 20787 21242 20821
rect 21672 20787 21688 20821
rect 22244 20787 22260 20821
rect 22690 20787 22706 20821
rect 23262 20787 23278 20821
rect 23708 20787 23724 20821
rect 24280 20787 24296 20821
rect 24726 20787 24742 20821
rect 25298 20787 25314 20821
rect 25744 20787 25760 20821
rect 26316 20787 26332 20821
rect 26762 20787 26778 20821
rect 27334 20787 27350 20821
rect 27780 20787 27796 20821
rect 28352 20787 28368 20821
rect 28798 20787 28814 20821
rect 29370 20787 29386 20821
rect 29816 20787 29832 20821
rect 30388 20787 30404 20821
rect 30834 20787 30850 20821
rect 31406 20787 31422 20821
rect 31852 20787 31868 20821
rect 32424 20787 32440 20821
rect 32870 20787 32886 20821
rect 33442 20787 33458 20821
rect 17154 20760 17188 20776
rect 13314 20683 13330 20717
rect 13886 20683 13902 20717
rect 14332 20683 14348 20717
rect 14904 20683 14920 20717
rect 15350 20683 15366 20717
rect 15922 20683 15938 20717
rect 16368 20683 16384 20717
rect 16940 20683 16956 20717
rect 13052 20560 13142 20590
rect 13052 20526 13080 20560
rect 13114 20526 13142 20560
rect 13052 20498 13142 20526
rect 14070 20560 14160 20590
rect 14070 20526 14098 20560
rect 14132 20526 14160 20560
rect 14070 20498 14160 20526
rect 15088 20560 15178 20590
rect 15088 20526 15116 20560
rect 15150 20526 15178 20560
rect 15088 20498 15178 20526
rect 16106 20560 16196 20590
rect 16106 20526 16134 20560
rect 16168 20526 16196 20560
rect 16106 20498 16196 20526
rect 18264 20576 18354 20606
rect 18264 20542 18292 20576
rect 18326 20542 18354 20576
rect 18264 20514 18354 20542
rect 19282 20576 19372 20606
rect 19282 20542 19310 20576
rect 19344 20542 19372 20576
rect 19282 20514 19372 20542
rect 20300 20576 20390 20606
rect 20300 20542 20328 20576
rect 20362 20542 20390 20576
rect 20300 20514 20390 20542
rect 21318 20576 21408 20606
rect 21318 20542 21346 20576
rect 21380 20542 21408 20576
rect 21318 20514 21408 20542
rect 22336 20576 22426 20606
rect 22336 20542 22364 20576
rect 22398 20542 22426 20576
rect 22336 20514 22426 20542
rect 23354 20576 23444 20606
rect 23354 20542 23382 20576
rect 23416 20542 23444 20576
rect 23354 20514 23444 20542
rect 24372 20576 24462 20606
rect 24372 20542 24400 20576
rect 24434 20542 24462 20576
rect 24372 20514 24462 20542
rect 25390 20576 25480 20606
rect 25390 20542 25418 20576
rect 25452 20542 25480 20576
rect 25390 20514 25480 20542
rect 26408 20576 26498 20606
rect 26408 20542 26436 20576
rect 26470 20542 26498 20576
rect 26408 20514 26498 20542
rect 27426 20576 27516 20606
rect 27426 20542 27454 20576
rect 27488 20542 27516 20576
rect 27426 20514 27516 20542
rect 28444 20576 28534 20606
rect 28444 20542 28472 20576
rect 28506 20542 28534 20576
rect 28444 20514 28534 20542
rect 29462 20576 29552 20606
rect 29462 20542 29490 20576
rect 29524 20542 29552 20576
rect 29462 20514 29552 20542
rect 30480 20576 30570 20606
rect 30480 20542 30508 20576
rect 30542 20542 30570 20576
rect 30480 20514 30570 20542
rect 31498 20576 31588 20606
rect 31498 20542 31526 20576
rect 31560 20542 31588 20576
rect 31498 20514 31588 20542
rect 32516 20576 32606 20606
rect 32516 20542 32544 20576
rect 32578 20542 32606 20576
rect 32516 20514 32606 20542
rect 33534 20576 33624 20606
rect 33534 20542 33562 20576
rect 33596 20542 33624 20576
rect 33534 20514 33624 20542
rect 13314 20379 13330 20413
rect 13886 20379 13902 20413
rect 14332 20379 14348 20413
rect 14904 20379 14920 20413
rect 15350 20379 15366 20413
rect 15922 20379 15938 20413
rect 16368 20379 16384 20413
rect 16940 20379 16956 20413
rect 13082 20320 13116 20336
rect 13082 19728 13116 19744
rect 14100 20320 14134 20336
rect 14100 19728 14134 19744
rect 15118 20320 15152 20336
rect 15118 19728 15152 19744
rect 16136 20320 16170 20336
rect 16136 19728 16170 19744
rect 17154 20320 17188 20336
rect 18618 20259 18634 20293
rect 19190 20259 19206 20293
rect 19636 20259 19652 20293
rect 20208 20259 20224 20293
rect 20654 20259 20670 20293
rect 21226 20259 21242 20293
rect 21672 20259 21688 20293
rect 22244 20259 22260 20293
rect 22690 20259 22706 20293
rect 23262 20259 23278 20293
rect 23708 20259 23724 20293
rect 24280 20259 24296 20293
rect 24726 20259 24742 20293
rect 25298 20259 25314 20293
rect 25744 20259 25760 20293
rect 26316 20259 26332 20293
rect 26762 20259 26778 20293
rect 27334 20259 27350 20293
rect 27780 20259 27796 20293
rect 28352 20259 28368 20293
rect 28798 20259 28814 20293
rect 29370 20259 29386 20293
rect 29816 20259 29832 20293
rect 30388 20259 30404 20293
rect 30834 20259 30850 20293
rect 31406 20259 31422 20293
rect 31852 20259 31868 20293
rect 32424 20259 32440 20293
rect 32870 20259 32886 20293
rect 33442 20259 33458 20293
rect 17154 19728 17188 19744
rect 18386 20200 18420 20216
rect 13314 19651 13330 19685
rect 13886 19651 13902 19685
rect 14332 19651 14348 19685
rect 14904 19651 14920 19685
rect 15350 19651 15366 19685
rect 15922 19651 15938 19685
rect 16368 19651 16384 19685
rect 16940 19651 16956 19685
rect 18386 19608 18420 19624
rect 19404 20200 19438 20216
rect 19404 19608 19438 19624
rect 20422 20200 20456 20216
rect 20422 19608 20456 19624
rect 21440 20200 21474 20216
rect 21440 19608 21474 19624
rect 22458 20200 22492 20216
rect 22458 19608 22492 19624
rect 23476 20200 23510 20216
rect 23476 19608 23510 19624
rect 24494 20200 24528 20216
rect 24494 19608 24528 19624
rect 25512 20200 25546 20216
rect 25512 19608 25546 19624
rect 26530 20200 26564 20216
rect 26530 19608 26564 19624
rect 27548 20200 27582 20216
rect 27548 19608 27582 19624
rect 28566 20200 28600 20216
rect 28566 19608 28600 19624
rect 29584 20200 29618 20216
rect 29584 19608 29618 19624
rect 30602 20200 30636 20216
rect 30602 19608 30636 19624
rect 31620 20200 31654 20216
rect 31620 19608 31654 19624
rect 32638 20200 32672 20216
rect 32638 19608 32672 19624
rect 33656 20200 33690 20216
rect 33656 19608 33690 19624
rect 13062 19532 13152 19562
rect 13062 19498 13090 19532
rect 13124 19498 13152 19532
rect 13062 19470 13152 19498
rect 14080 19532 14170 19562
rect 14080 19498 14108 19532
rect 14142 19498 14170 19532
rect 14080 19470 14170 19498
rect 15098 19532 15188 19562
rect 15098 19498 15126 19532
rect 15160 19498 15188 19532
rect 15098 19470 15188 19498
rect 16116 19532 16206 19562
rect 16116 19498 16144 19532
rect 16178 19498 16206 19532
rect 18618 19531 18634 19565
rect 19190 19531 19206 19565
rect 19636 19531 19652 19565
rect 20208 19531 20224 19565
rect 20654 19531 20670 19565
rect 21226 19531 21242 19565
rect 21672 19531 21688 19565
rect 22244 19531 22260 19565
rect 22690 19531 22706 19565
rect 23262 19531 23278 19565
rect 23708 19531 23724 19565
rect 24280 19531 24296 19565
rect 24726 19531 24742 19565
rect 25298 19531 25314 19565
rect 25744 19531 25760 19565
rect 26316 19531 26332 19565
rect 26762 19531 26778 19565
rect 27334 19531 27350 19565
rect 27780 19531 27796 19565
rect 28352 19531 28368 19565
rect 28798 19531 28814 19565
rect 29370 19531 29386 19565
rect 29816 19531 29832 19565
rect 30388 19531 30404 19565
rect 30834 19531 30850 19565
rect 31406 19531 31422 19565
rect 31852 19531 31868 19565
rect 32424 19531 32440 19565
rect 32870 19531 32886 19565
rect 33442 19531 33458 19565
rect 16116 19470 16206 19498
rect 13314 19347 13330 19381
rect 13886 19347 13902 19381
rect 14332 19347 14348 19381
rect 14904 19347 14920 19381
rect 15350 19347 15366 19381
rect 15922 19347 15938 19381
rect 16368 19347 16384 19381
rect 16940 19347 16956 19381
rect 18288 19308 18378 19338
rect 13082 19288 13116 19304
rect 13082 18696 13116 18712
rect 14100 19288 14134 19304
rect 14100 18696 14134 18712
rect 15118 19288 15152 19304
rect 15118 18696 15152 18712
rect 16136 19288 16170 19304
rect 16136 18696 16170 18712
rect 17154 19288 17188 19304
rect 18288 19274 18316 19308
rect 18350 19274 18378 19308
rect 18288 19246 18378 19274
rect 19306 19308 19396 19338
rect 19306 19274 19334 19308
rect 19368 19274 19396 19308
rect 19306 19246 19396 19274
rect 20324 19308 20414 19338
rect 20324 19274 20352 19308
rect 20386 19274 20414 19308
rect 20324 19246 20414 19274
rect 21342 19308 21432 19338
rect 21342 19274 21370 19308
rect 21404 19274 21432 19308
rect 21342 19246 21432 19274
rect 22360 19308 22450 19338
rect 22360 19274 22388 19308
rect 22422 19274 22450 19308
rect 22360 19246 22450 19274
rect 23378 19308 23468 19338
rect 23378 19274 23406 19308
rect 23440 19274 23468 19308
rect 23378 19246 23468 19274
rect 24396 19308 24486 19338
rect 24396 19274 24424 19308
rect 24458 19274 24486 19308
rect 24396 19246 24486 19274
rect 25414 19308 25504 19338
rect 25414 19274 25442 19308
rect 25476 19274 25504 19308
rect 25414 19246 25504 19274
rect 26432 19308 26522 19338
rect 26432 19274 26460 19308
rect 26494 19274 26522 19308
rect 26432 19246 26522 19274
rect 27450 19308 27540 19338
rect 27450 19274 27478 19308
rect 27512 19274 27540 19308
rect 27450 19246 27540 19274
rect 28468 19308 28558 19338
rect 28468 19274 28496 19308
rect 28530 19274 28558 19308
rect 28468 19246 28558 19274
rect 29486 19308 29576 19338
rect 29486 19274 29514 19308
rect 29548 19274 29576 19308
rect 29486 19246 29576 19274
rect 30504 19308 30594 19338
rect 30504 19274 30532 19308
rect 30566 19274 30594 19308
rect 30504 19246 30594 19274
rect 31522 19308 31612 19338
rect 31522 19274 31550 19308
rect 31584 19274 31612 19308
rect 31522 19246 31612 19274
rect 32540 19308 32630 19338
rect 32540 19274 32568 19308
rect 32602 19274 32630 19308
rect 32540 19246 32630 19274
rect 33558 19308 33648 19338
rect 33558 19274 33586 19308
rect 33620 19274 33648 19308
rect 33558 19246 33648 19274
rect 18618 19003 18634 19037
rect 19190 19003 19206 19037
rect 19636 19003 19652 19037
rect 20208 19003 20224 19037
rect 20654 19003 20670 19037
rect 21226 19003 21242 19037
rect 21672 19003 21688 19037
rect 22244 19003 22260 19037
rect 22690 19003 22706 19037
rect 23262 19003 23278 19037
rect 23708 19003 23724 19037
rect 24280 19003 24296 19037
rect 24726 19003 24742 19037
rect 25298 19003 25314 19037
rect 25744 19003 25760 19037
rect 26316 19003 26332 19037
rect 26762 19003 26778 19037
rect 27334 19003 27350 19037
rect 27780 19003 27796 19037
rect 28352 19003 28368 19037
rect 28798 19003 28814 19037
rect 29370 19003 29386 19037
rect 29816 19003 29832 19037
rect 30388 19003 30404 19037
rect 30834 19003 30850 19037
rect 31406 19003 31422 19037
rect 31852 19003 31868 19037
rect 32424 19003 32440 19037
rect 32870 19003 32886 19037
rect 33442 19003 33458 19037
rect 17154 18696 17188 18712
rect 18386 18944 18420 18960
rect 13314 18619 13330 18653
rect 13886 18619 13902 18653
rect 14332 18619 14348 18653
rect 14904 18619 14920 18653
rect 15350 18619 15366 18653
rect 15922 18619 15938 18653
rect 16368 18619 16384 18653
rect 16940 18619 16956 18653
rect 13052 18504 13142 18534
rect 13052 18470 13080 18504
rect 13114 18470 13142 18504
rect 13052 18442 13142 18470
rect 14070 18504 14160 18534
rect 14070 18470 14098 18504
rect 14132 18470 14160 18504
rect 14070 18442 14160 18470
rect 15088 18504 15178 18534
rect 15088 18470 15116 18504
rect 15150 18470 15178 18504
rect 15088 18442 15178 18470
rect 16106 18504 16196 18534
rect 16106 18470 16134 18504
rect 16168 18470 16196 18504
rect 16106 18442 16196 18470
rect 18386 18352 18420 18368
rect 19404 18944 19438 18960
rect 19404 18352 19438 18368
rect 20422 18944 20456 18960
rect 20422 18352 20456 18368
rect 21440 18944 21474 18960
rect 21440 18352 21474 18368
rect 22458 18944 22492 18960
rect 22458 18352 22492 18368
rect 23476 18944 23510 18960
rect 23476 18352 23510 18368
rect 24494 18944 24528 18960
rect 24494 18352 24528 18368
rect 25512 18944 25546 18960
rect 25512 18352 25546 18368
rect 26530 18944 26564 18960
rect 26530 18352 26564 18368
rect 27548 18944 27582 18960
rect 27548 18352 27582 18368
rect 28566 18944 28600 18960
rect 28566 18352 28600 18368
rect 29584 18944 29618 18960
rect 29584 18352 29618 18368
rect 30602 18944 30636 18960
rect 30602 18352 30636 18368
rect 31620 18944 31654 18960
rect 31620 18352 31654 18368
rect 32638 18944 32672 18960
rect 32638 18352 32672 18368
rect 33656 18944 33690 18960
rect 33656 18352 33690 18368
rect 13314 18315 13330 18349
rect 13886 18315 13902 18349
rect 14332 18315 14348 18349
rect 14904 18315 14920 18349
rect 15350 18315 15366 18349
rect 15922 18315 15938 18349
rect 16368 18315 16384 18349
rect 16940 18315 16956 18349
rect 18618 18275 18634 18309
rect 19190 18275 19206 18309
rect 19636 18275 19652 18309
rect 20208 18275 20224 18309
rect 20654 18275 20670 18309
rect 21226 18275 21242 18309
rect 21672 18275 21688 18309
rect 22244 18275 22260 18309
rect 22690 18275 22706 18309
rect 23262 18275 23278 18309
rect 23708 18275 23724 18309
rect 24280 18275 24296 18309
rect 24726 18275 24742 18309
rect 25298 18275 25314 18309
rect 25744 18275 25760 18309
rect 26316 18275 26332 18309
rect 26762 18275 26778 18309
rect 27334 18275 27350 18309
rect 27780 18275 27796 18309
rect 28352 18275 28368 18309
rect 28798 18275 28814 18309
rect 29370 18275 29386 18309
rect 29816 18275 29832 18309
rect 30388 18275 30404 18309
rect 30834 18275 30850 18309
rect 31406 18275 31422 18309
rect 31852 18275 31868 18309
rect 32424 18275 32440 18309
rect 32870 18275 32886 18309
rect 33442 18275 33458 18309
rect 13082 18256 13116 18272
rect 13082 17664 13116 17680
rect 14100 18256 14134 18272
rect 14100 17664 14134 17680
rect 15118 18256 15152 18272
rect 15118 17664 15152 17680
rect 16136 18256 16170 18272
rect 16136 17664 16170 17680
rect 17154 18256 17188 18272
rect 18152 18064 18242 18094
rect 18152 18030 18180 18064
rect 18214 18030 18242 18064
rect 18152 18002 18242 18030
rect 19170 18064 19260 18094
rect 19170 18030 19198 18064
rect 19232 18030 19260 18064
rect 19170 18002 19260 18030
rect 20188 18064 20278 18094
rect 20188 18030 20216 18064
rect 20250 18030 20278 18064
rect 20188 18002 20278 18030
rect 21206 18064 21296 18094
rect 21206 18030 21234 18064
rect 21268 18030 21296 18064
rect 21206 18002 21296 18030
rect 22224 18064 22314 18094
rect 22224 18030 22252 18064
rect 22286 18030 22314 18064
rect 22224 18002 22314 18030
rect 23242 18064 23332 18094
rect 23242 18030 23270 18064
rect 23304 18030 23332 18064
rect 23242 18002 23332 18030
rect 24260 18064 24350 18094
rect 24260 18030 24288 18064
rect 24322 18030 24350 18064
rect 24260 18002 24350 18030
rect 25278 18064 25368 18094
rect 25278 18030 25306 18064
rect 25340 18030 25368 18064
rect 25278 18002 25368 18030
rect 26296 18064 26386 18094
rect 26296 18030 26324 18064
rect 26358 18030 26386 18064
rect 26296 18002 26386 18030
rect 27314 18064 27404 18094
rect 27314 18030 27342 18064
rect 27376 18030 27404 18064
rect 27314 18002 27404 18030
rect 28332 18064 28422 18094
rect 28332 18030 28360 18064
rect 28394 18030 28422 18064
rect 28332 18002 28422 18030
rect 29350 18064 29440 18094
rect 29350 18030 29378 18064
rect 29412 18030 29440 18064
rect 29350 18002 29440 18030
rect 30368 18064 30458 18094
rect 30368 18030 30396 18064
rect 30430 18030 30458 18064
rect 30368 18002 30458 18030
rect 31386 18064 31476 18094
rect 31386 18030 31414 18064
rect 31448 18030 31476 18064
rect 31386 18002 31476 18030
rect 32404 18064 32494 18094
rect 32404 18030 32432 18064
rect 32466 18030 32494 18064
rect 32404 18002 32494 18030
rect 33422 18064 33512 18094
rect 33422 18030 33450 18064
rect 33484 18030 33512 18064
rect 33422 18002 33512 18030
rect 18618 17747 18634 17781
rect 19190 17747 19206 17781
rect 19636 17747 19652 17781
rect 20208 17747 20224 17781
rect 20654 17747 20670 17781
rect 21226 17747 21242 17781
rect 21672 17747 21688 17781
rect 22244 17747 22260 17781
rect 22690 17747 22706 17781
rect 23262 17747 23278 17781
rect 23708 17747 23724 17781
rect 24280 17747 24296 17781
rect 24726 17747 24742 17781
rect 25298 17747 25314 17781
rect 25744 17747 25760 17781
rect 26316 17747 26332 17781
rect 26762 17747 26778 17781
rect 27334 17747 27350 17781
rect 27780 17747 27796 17781
rect 28352 17747 28368 17781
rect 28798 17747 28814 17781
rect 29370 17747 29386 17781
rect 29816 17747 29832 17781
rect 30388 17747 30404 17781
rect 30834 17747 30850 17781
rect 31406 17747 31422 17781
rect 31852 17747 31868 17781
rect 32424 17747 32440 17781
rect 32870 17747 32886 17781
rect 33442 17747 33458 17781
rect 17154 17664 17188 17680
rect 18386 17688 18420 17704
rect 13314 17587 13330 17621
rect 13886 17587 13902 17621
rect 14332 17587 14348 17621
rect 14904 17587 14920 17621
rect 15350 17587 15366 17621
rect 15922 17587 15938 17621
rect 16368 17587 16384 17621
rect 16940 17587 16956 17621
rect 13576 17352 13666 17382
rect 13576 17318 13604 17352
rect 13638 17318 13666 17352
rect 13576 17290 13666 17318
rect 14594 17352 14684 17382
rect 14594 17318 14622 17352
rect 14656 17318 14684 17352
rect 14594 17290 14684 17318
rect 15612 17352 15702 17382
rect 15612 17318 15640 17352
rect 15674 17318 15702 17352
rect 15612 17290 15702 17318
rect 16630 17352 16720 17382
rect 16630 17318 16658 17352
rect 16692 17318 16720 17352
rect 16630 17290 16720 17318
rect 18386 17096 18420 17112
rect 19404 17688 19438 17704
rect 19404 17096 19438 17112
rect 20422 17688 20456 17704
rect 20422 17096 20456 17112
rect 21440 17688 21474 17704
rect 21440 17096 21474 17112
rect 22458 17688 22492 17704
rect 22458 17096 22492 17112
rect 23476 17688 23510 17704
rect 23476 17096 23510 17112
rect 24494 17688 24528 17704
rect 24494 17096 24528 17112
rect 25512 17688 25546 17704
rect 25512 17096 25546 17112
rect 26530 17688 26564 17704
rect 26530 17096 26564 17112
rect 27548 17688 27582 17704
rect 27548 17096 27582 17112
rect 28566 17688 28600 17704
rect 28566 17096 28600 17112
rect 29584 17688 29618 17704
rect 29584 17096 29618 17112
rect 30602 17688 30636 17704
rect 30602 17096 30636 17112
rect 31620 17688 31654 17704
rect 31620 17096 31654 17112
rect 32638 17688 32672 17704
rect 32638 17096 32672 17112
rect 33656 17688 33690 17704
rect 33656 17096 33690 17112
rect 18618 17019 18634 17053
rect 19190 17019 19206 17053
rect 19636 17019 19652 17053
rect 20208 17019 20224 17053
rect 20654 17019 20670 17053
rect 21226 17019 21242 17053
rect 21672 17019 21688 17053
rect 22244 17019 22260 17053
rect 22690 17019 22706 17053
rect 23262 17019 23278 17053
rect 23708 17019 23724 17053
rect 24280 17019 24296 17053
rect 24726 17019 24742 17053
rect 25298 17019 25314 17053
rect 25744 17019 25760 17053
rect 26316 17019 26332 17053
rect 26762 17019 26778 17053
rect 27334 17019 27350 17053
rect 27780 17019 27796 17053
rect 28352 17019 28368 17053
rect 28798 17019 28814 17053
rect 29370 17019 29386 17053
rect 29816 17019 29832 17053
rect 30388 17019 30404 17053
rect 30834 17019 30850 17053
rect 31406 17019 31422 17053
rect 31852 17019 31868 17053
rect 32424 17019 32440 17053
rect 32870 17019 32886 17053
rect 33442 17019 33458 17053
rect -12280 16276 -12234 16309
rect -10540 16276 -10470 16309
rect -12280 16275 -12184 16276
rect -10566 16275 -10470 16276
rect -12280 16213 -12246 16275
rect -10504 16214 -10470 16275
rect -12086 16173 -12070 16207
rect -11970 16173 -11954 16207
rect -11828 16173 -11812 16207
rect -11712 16173 -11696 16207
rect -11570 16173 -11554 16207
rect -11454 16173 -11438 16207
rect -11312 16173 -11296 16207
rect -11196 16173 -11180 16207
rect -11054 16173 -11038 16207
rect -10938 16173 -10922 16207
rect -10796 16173 -10780 16207
rect -10680 16173 -10664 16207
rect -12166 16114 -12132 16130
rect -12166 15722 -12132 15738
rect -11908 16114 -11874 16130
rect -11908 15722 -11874 15738
rect -11650 16114 -11616 16130
rect -11650 15722 -11616 15738
rect -11392 16114 -11358 16130
rect -11392 15722 -11358 15738
rect -11134 16114 -11100 16130
rect -11134 15722 -11100 15738
rect -10876 16114 -10842 16130
rect -10876 15722 -10842 15738
rect -10618 16114 -10584 16130
rect -10618 15722 -10584 15738
rect -12086 15645 -12070 15679
rect -11970 15645 -11954 15679
rect -11828 15645 -11812 15679
rect -11712 15645 -11696 15679
rect -11570 15645 -11554 15679
rect -11454 15645 -11438 15679
rect -11312 15645 -11296 15679
rect -11196 15645 -11180 15679
rect -11054 15645 -11038 15679
rect -10938 15645 -10922 15679
rect -10796 15645 -10780 15679
rect -10680 15645 -10664 15679
rect -12280 15577 -12246 15639
rect -9680 16276 -9634 16309
rect -7940 16276 -7870 16309
rect -9680 16275 -9584 16276
rect -7966 16275 -7870 16276
rect -9680 16213 -9646 16275
rect -7904 16214 -7870 16275
rect -10396 15773 -10367 15807
rect -10333 15773 -10275 15807
rect -10241 15773 -10183 15807
rect -10149 15773 -10120 15807
rect -10504 15577 -10470 15638
rect -12280 15576 -12184 15577
rect -12280 15543 -12234 15576
rect -10540 15544 -10470 15577
rect -10566 15543 -10470 15544
rect -10330 15731 -10264 15739
rect -10330 15697 -10314 15731
rect -10280 15697 -10264 15731
rect -10330 15663 -10264 15697
rect -10330 15629 -10314 15663
rect -10280 15629 -10264 15663
rect -10330 15595 -10264 15629
rect -10330 15561 -10314 15595
rect -10280 15561 -10264 15595
rect -10330 15543 -10264 15561
rect -10230 15731 -10188 15773
rect -10196 15697 -10188 15731
rect -10230 15663 -10188 15697
rect -10196 15629 -10188 15663
rect -9486 16173 -9470 16207
rect -9370 16173 -9354 16207
rect -9228 16173 -9212 16207
rect -9112 16173 -9096 16207
rect -8970 16173 -8954 16207
rect -8854 16173 -8838 16207
rect -8712 16173 -8696 16207
rect -8596 16173 -8580 16207
rect -8454 16173 -8438 16207
rect -8338 16173 -8322 16207
rect -8196 16173 -8180 16207
rect -8080 16173 -8064 16207
rect -9566 16114 -9532 16130
rect -9566 15722 -9532 15738
rect -9308 16114 -9274 16130
rect -9308 15722 -9274 15738
rect -9050 16114 -9016 16130
rect -9050 15722 -9016 15738
rect -8792 16114 -8758 16130
rect -8792 15722 -8758 15738
rect -8534 16114 -8500 16130
rect -8534 15722 -8500 15738
rect -8276 16114 -8242 16130
rect -8276 15722 -8242 15738
rect -8018 16114 -7984 16130
rect -8018 15722 -7984 15738
rect -9486 15645 -9470 15679
rect -9370 15645 -9354 15679
rect -9228 15645 -9212 15679
rect -9112 15645 -9096 15679
rect -8970 15645 -8954 15679
rect -8854 15645 -8838 15679
rect -8712 15645 -8696 15679
rect -8596 15645 -8580 15679
rect -8454 15645 -8438 15679
rect -8338 15645 -8322 15679
rect -8196 15645 -8180 15679
rect -8080 15645 -8064 15679
rect -10230 15595 -10188 15629
rect -10196 15561 -10188 15595
rect -10230 15545 -10188 15561
rect -9680 15577 -9646 15639
rect 11290 16192 11390 16354
rect 35634 16192 35734 16354
rect -7796 15773 -7767 15807
rect -7733 15773 -7675 15807
rect -7641 15773 -7583 15807
rect -7549 15773 -7520 15807
rect -7346 15773 -7317 15807
rect -7283 15773 -7225 15807
rect -7191 15773 -7133 15807
rect -7099 15773 -7070 15807
rect -7904 15577 -7870 15638
rect -9680 15576 -9584 15577
rect -9680 15543 -9634 15576
rect -7940 15544 -7870 15577
rect -7966 15543 -7870 15544
rect -7730 15731 -7664 15739
rect -7730 15697 -7714 15731
rect -7680 15697 -7664 15731
rect -7730 15663 -7664 15697
rect -7730 15629 -7714 15663
rect -7680 15629 -7664 15663
rect -7730 15595 -7664 15629
rect -7730 15561 -7714 15595
rect -7680 15561 -7664 15595
rect -7730 15543 -7664 15561
rect -7630 15731 -7588 15773
rect -7596 15697 -7588 15731
rect -7630 15663 -7588 15697
rect -7596 15629 -7588 15663
rect -7630 15595 -7588 15629
rect -7596 15561 -7588 15595
rect -7630 15545 -7588 15561
rect -7280 15731 -7214 15739
rect -7280 15697 -7264 15731
rect -7230 15697 -7214 15731
rect -7280 15663 -7214 15697
rect -7280 15629 -7264 15663
rect -7230 15629 -7214 15663
rect -7280 15595 -7214 15629
rect -7280 15561 -7264 15595
rect -7230 15561 -7214 15595
rect -7280 15543 -7214 15561
rect -7180 15731 -7138 15773
rect -7146 15697 -7138 15731
rect -7180 15663 -7138 15697
rect -7146 15629 -7138 15663
rect -7180 15595 -7138 15629
rect -7146 15561 -7138 15595
rect -7180 15545 -7138 15561
rect -10330 15484 -10284 15543
rect -10289 15436 -10284 15484
rect -10250 15506 -10184 15509
rect -10250 15495 -10233 15506
rect -10250 15461 -10234 15495
rect -10187 15466 -10184 15506
rect -7730 15484 -7684 15543
rect -10200 15461 -10184 15466
rect -7689 15436 -7684 15484
rect -7650 15506 -7584 15509
rect -7280 15506 -7234 15543
rect -7650 15495 -7633 15506
rect -7650 15461 -7634 15495
rect -7587 15466 -7584 15506
rect -7600 15461 -7584 15466
rect -7240 15458 -7234 15506
rect -7200 15461 -7184 15509
rect -7136 15462 -7134 15509
rect -7150 15461 -7134 15462
rect -10330 15423 -10284 15436
rect -10330 15411 -10264 15423
rect -10330 15377 -10314 15411
rect -10280 15377 -10264 15411
rect -12280 15342 -12210 15376
rect -10540 15342 -10470 15376
rect -12280 15280 -12246 15342
rect -10504 15280 -10470 15342
rect -10330 15343 -10264 15377
rect -10330 15309 -10314 15343
rect -10280 15309 -10264 15343
rect -10330 15297 -10264 15309
rect -10230 15411 -10184 15427
rect -10196 15377 -10184 15411
rect -7730 15423 -7684 15436
rect -7730 15411 -7664 15423
rect -10230 15343 -10184 15377
rect -7730 15377 -7714 15411
rect -7680 15377 -7664 15411
rect -10196 15309 -10184 15343
rect -12086 15240 -12070 15274
rect -11970 15240 -11954 15274
rect -11828 15240 -11812 15274
rect -11712 15240 -11696 15274
rect -11570 15240 -11554 15274
rect -11454 15240 -11438 15274
rect -11312 15240 -11296 15274
rect -11196 15240 -11180 15274
rect -11054 15240 -11038 15274
rect -10938 15240 -10922 15274
rect -10796 15240 -10780 15274
rect -10680 15240 -10664 15274
rect -12166 15190 -12132 15206
rect -12166 14998 -12132 15014
rect -11908 15190 -11874 15206
rect -11908 14998 -11874 15014
rect -11650 15190 -11616 15206
rect -11650 14998 -11616 15014
rect -11392 15190 -11358 15206
rect -11392 14998 -11358 15014
rect -11134 15190 -11100 15206
rect -11134 14998 -11100 15014
rect -10876 15190 -10842 15206
rect -10876 14998 -10842 15014
rect -10618 15190 -10584 15206
rect -10618 14998 -10584 15014
rect -12086 14930 -12070 14964
rect -11970 14930 -11954 14964
rect -11828 14930 -11812 14964
rect -11712 14930 -11696 14964
rect -11570 14930 -11554 14964
rect -11454 14930 -11438 14964
rect -11312 14930 -11296 14964
rect -11196 14930 -11180 14964
rect -11054 14930 -11038 14964
rect -10938 14930 -10922 14964
rect -10796 14930 -10780 14964
rect -10680 14930 -10664 14964
rect -10230 15263 -10184 15309
rect -9680 15342 -9610 15376
rect -7940 15342 -7870 15376
rect -9680 15280 -9646 15342
rect -7904 15280 -7870 15342
rect -7730 15343 -7664 15377
rect -7730 15309 -7714 15343
rect -7680 15309 -7664 15343
rect -7730 15297 -7664 15309
rect -7630 15411 -7584 15427
rect -7596 15377 -7584 15411
rect -7630 15343 -7584 15377
rect -7596 15309 -7584 15343
rect -10396 15229 -10367 15263
rect -10333 15229 -10275 15263
rect -10241 15229 -10183 15263
rect -10149 15229 -10120 15263
rect -9486 15240 -9470 15274
rect -9370 15240 -9354 15274
rect -9228 15240 -9212 15274
rect -9112 15240 -9096 15274
rect -8970 15240 -8954 15274
rect -8854 15240 -8838 15274
rect -8712 15240 -8696 15274
rect -8596 15240 -8580 15274
rect -8454 15240 -8438 15274
rect -8338 15240 -8322 15274
rect -8196 15240 -8180 15274
rect -8080 15240 -8064 15274
rect -9566 15190 -9532 15206
rect -9566 14998 -9532 15014
rect -9308 15190 -9274 15206
rect -9308 14998 -9274 15014
rect -9050 15190 -9016 15206
rect -9050 14998 -9016 15014
rect -8792 15190 -8758 15206
rect -8792 14998 -8758 15014
rect -8534 15190 -8500 15206
rect -8534 14998 -8500 15014
rect -8276 15190 -8242 15206
rect -8276 14998 -8242 15014
rect -8018 15190 -7984 15206
rect -8018 14998 -7984 15014
rect -9486 14930 -9470 14964
rect -9370 14930 -9354 14964
rect -9228 14930 -9212 14964
rect -9112 14930 -9096 14964
rect -8970 14930 -8954 14964
rect -8854 14930 -8838 14964
rect -8712 14930 -8696 14964
rect -8596 14930 -8580 14964
rect -8454 14930 -8438 14964
rect -8338 14930 -8322 14964
rect -8196 14930 -8180 14964
rect -8080 14930 -8064 14964
rect -7630 15263 -7584 15309
rect -7280 15423 -7234 15458
rect -7280 15411 -7214 15423
rect -7280 15377 -7264 15411
rect -7230 15377 -7214 15411
rect -7280 15343 -7214 15377
rect -7280 15309 -7264 15343
rect -7230 15309 -7214 15343
rect -7280 15297 -7214 15309
rect -7180 15411 -7134 15427
rect -7146 15377 -7134 15411
rect -7180 15343 -7134 15377
rect -7146 15309 -7134 15343
rect -7180 15263 -7134 15309
rect -7796 15229 -7767 15263
rect -7733 15229 -7675 15263
rect -7641 15229 -7583 15263
rect -7549 15229 -7520 15263
rect -7346 15229 -7317 15263
rect -7283 15229 -7225 15263
rect -7191 15229 -7133 15263
rect -7099 15229 -7070 15263
rect -1410 15200 -1310 15362
rect -12280 14862 -12246 14924
rect -10504 14862 -10470 14924
rect -12280 14828 -12212 14862
rect -10538 14828 -10470 14862
rect -9680 14862 -9646 14924
rect -7904 14862 -7870 14924
rect -9680 14828 -9612 14862
rect -7938 14828 -7870 14862
rect 35734 15200 35834 15362
rect 13998 14756 14080 14780
rect 13998 14722 14022 14756
rect 14056 14722 14080 14756
rect 13998 14698 14080 14722
rect 15016 14756 15098 14780
rect 15016 14722 15040 14756
rect 15074 14722 15098 14756
rect 15016 14698 15098 14722
rect 16034 14756 16116 14780
rect 16034 14722 16058 14756
rect 16092 14722 16116 14756
rect 16034 14698 16116 14722
rect 17052 14756 17134 14780
rect 17052 14722 17076 14756
rect 17110 14722 17134 14756
rect 17052 14698 17134 14722
rect 18070 14756 18152 14780
rect 18070 14722 18094 14756
rect 18128 14722 18152 14756
rect 18070 14698 18152 14722
rect 19088 14756 19170 14780
rect 19088 14722 19112 14756
rect 19146 14722 19170 14756
rect 19088 14698 19170 14722
rect 20106 14756 20188 14780
rect 20106 14722 20130 14756
rect 20164 14722 20188 14756
rect 20106 14698 20188 14722
rect 21124 14756 21206 14780
rect 21124 14722 21148 14756
rect 21182 14722 21206 14756
rect 21124 14698 21206 14722
rect 22142 14756 22224 14780
rect 22142 14722 22166 14756
rect 22200 14722 22224 14756
rect 22142 14698 22224 14722
rect 23160 14756 23242 14780
rect 23160 14722 23184 14756
rect 23218 14722 23242 14756
rect 23160 14698 23242 14722
rect 24178 14756 24260 14780
rect 24178 14722 24202 14756
rect 24236 14722 24260 14756
rect 24178 14698 24260 14722
rect 25196 14756 25278 14780
rect 25196 14722 25220 14756
rect 25254 14722 25278 14756
rect 25196 14698 25278 14722
rect 26214 14756 26296 14780
rect 26214 14722 26238 14756
rect 26272 14722 26296 14756
rect 26214 14698 26296 14722
rect 27232 14756 27314 14780
rect 27232 14722 27256 14756
rect 27290 14722 27314 14756
rect 27232 14698 27314 14722
rect 28250 14756 28332 14780
rect 28250 14722 28274 14756
rect 28308 14722 28332 14756
rect 28250 14698 28332 14722
rect 29268 14756 29350 14780
rect 29268 14722 29292 14756
rect 29326 14722 29350 14756
rect 29268 14698 29350 14722
rect 30286 14756 30368 14780
rect 30286 14722 30310 14756
rect 30344 14722 30368 14756
rect 30286 14698 30368 14722
rect 31304 14756 31386 14780
rect 31304 14722 31328 14756
rect 31362 14722 31386 14756
rect 31304 14698 31386 14722
rect 32322 14756 32404 14780
rect 32322 14722 32346 14756
rect 32380 14722 32404 14756
rect 32322 14698 32404 14722
rect 33340 14756 33422 14780
rect 33340 14722 33364 14756
rect 33398 14722 33422 14756
rect 33340 14698 33422 14722
rect 13726 14542 13742 14576
rect 14298 14542 14314 14576
rect 14744 14542 14760 14576
rect 15316 14542 15332 14576
rect 15762 14542 15778 14576
rect 16334 14542 16350 14576
rect 16780 14542 16796 14576
rect 17352 14542 17368 14576
rect 17798 14542 17814 14576
rect 18370 14542 18386 14576
rect 18816 14542 18832 14576
rect 19388 14542 19404 14576
rect 19834 14542 19850 14576
rect 20406 14542 20422 14576
rect 20852 14542 20868 14576
rect 21424 14542 21440 14576
rect 21870 14542 21886 14576
rect 22442 14542 22458 14576
rect 22888 14542 22904 14576
rect 23460 14542 23476 14576
rect 23906 14542 23922 14576
rect 24478 14542 24494 14576
rect 24924 14542 24940 14576
rect 25496 14542 25512 14576
rect 25942 14542 25958 14576
rect 26514 14542 26530 14576
rect 26960 14542 26976 14576
rect 27532 14542 27548 14576
rect 27978 14542 27994 14576
rect 28550 14542 28566 14576
rect 28996 14542 29012 14576
rect 29568 14542 29584 14576
rect 30014 14542 30030 14576
rect 30586 14542 30602 14576
rect 31032 14542 31048 14576
rect 31604 14542 31620 14576
rect 32050 14542 32066 14576
rect 32622 14542 32638 14576
rect 33068 14542 33084 14576
rect 33640 14542 33656 14576
rect 13494 14492 13528 14508
rect 1704 14154 1786 14178
rect 1704 14120 1728 14154
rect 1762 14120 1786 14154
rect 1704 14096 1786 14120
rect 2722 14154 2804 14178
rect 2722 14120 2746 14154
rect 2780 14120 2804 14154
rect 1960 14066 1976 14100
rect 2532 14066 2548 14100
rect 2722 14096 2804 14120
rect 3740 14154 3822 14178
rect 3740 14120 3764 14154
rect 3798 14120 3822 14154
rect 2978 14066 2994 14100
rect 3550 14066 3566 14100
rect 3740 14096 3822 14120
rect 4758 14154 4840 14178
rect 4758 14120 4782 14154
rect 4816 14120 4840 14154
rect 3996 14066 4012 14100
rect 4568 14066 4584 14100
rect 4758 14096 4840 14120
rect 5776 14154 5858 14178
rect 5776 14120 5800 14154
rect 5834 14120 5858 14154
rect 5014 14066 5030 14100
rect 5586 14066 5602 14100
rect 5776 14096 5858 14120
rect 6794 14154 6876 14178
rect 6794 14120 6818 14154
rect 6852 14120 6876 14154
rect 6032 14066 6048 14100
rect 6604 14066 6620 14100
rect 6794 14096 6876 14120
rect 7812 14154 7894 14178
rect 7812 14120 7836 14154
rect 7870 14120 7894 14154
rect 7050 14066 7066 14100
rect 7622 14066 7638 14100
rect 7812 14096 7894 14120
rect 8830 14154 8912 14178
rect 8830 14120 8854 14154
rect 8888 14120 8912 14154
rect 8068 14066 8084 14100
rect 8640 14066 8656 14100
rect 8830 14096 8912 14120
rect 9848 14154 9930 14178
rect 9848 14120 9872 14154
rect 9906 14120 9930 14154
rect 9086 14066 9102 14100
rect 9658 14066 9674 14100
rect 9848 14096 9930 14120
rect 10876 14154 10958 14178
rect 10876 14120 10900 14154
rect 10934 14120 10958 14154
rect 10104 14066 10120 14100
rect 10676 14066 10692 14100
rect 10876 14096 10958 14120
rect 1728 14016 1762 14032
rect 1728 13424 1762 13440
rect 2746 14016 2780 14032
rect 2746 13424 2780 13440
rect 3764 14016 3798 14032
rect 3764 13424 3798 13440
rect 4782 14016 4816 14032
rect 4782 13424 4816 13440
rect 5800 14016 5834 14032
rect 5800 13424 5834 13440
rect 6818 14016 6852 14032
rect 6818 13424 6852 13440
rect 7836 14016 7870 14032
rect 7836 13424 7870 13440
rect 8854 14016 8888 14032
rect 8854 13424 8888 13440
rect 9872 14016 9906 14032
rect 9872 13424 9906 13440
rect 10890 14016 10924 14032
rect 13494 13900 13528 13916
rect 14512 14492 14546 14508
rect 14512 13900 14546 13916
rect 15530 14492 15564 14508
rect 15530 13900 15564 13916
rect 16548 14492 16582 14508
rect 16548 13900 16582 13916
rect 17566 14492 17600 14508
rect 17566 13900 17600 13916
rect 18584 14492 18618 14508
rect 18584 13900 18618 13916
rect 19602 14492 19636 14508
rect 19602 13900 19636 13916
rect 20620 14492 20654 14508
rect 20620 13900 20654 13916
rect 21638 14492 21672 14508
rect 21638 13900 21672 13916
rect 22656 14492 22690 14508
rect 22656 13900 22690 13916
rect 23674 14492 23708 14508
rect 23674 13900 23708 13916
rect 24692 14492 24726 14508
rect 24692 13900 24726 13916
rect 25710 14492 25744 14508
rect 25710 13900 25744 13916
rect 26728 14492 26762 14508
rect 26728 13900 26762 13916
rect 27746 14492 27780 14508
rect 27746 13900 27780 13916
rect 28764 14492 28798 14508
rect 28764 13900 28798 13916
rect 29782 14492 29816 14508
rect 29782 13900 29816 13916
rect 30800 14492 30834 14508
rect 30800 13900 30834 13916
rect 31818 14492 31852 14508
rect 31818 13900 31852 13916
rect 32836 14492 32870 14508
rect 32836 13900 32870 13916
rect 33854 14492 33888 14508
rect 33854 13900 33888 13916
rect 13726 13832 13742 13866
rect 14298 13832 14314 13866
rect 14744 13832 14760 13866
rect 15316 13832 15332 13866
rect 15762 13832 15778 13866
rect 16334 13832 16350 13866
rect 16780 13832 16796 13866
rect 17352 13832 17368 13866
rect 17798 13832 17814 13866
rect 18370 13832 18386 13866
rect 18816 13832 18832 13866
rect 19388 13832 19404 13866
rect 19834 13832 19850 13866
rect 20406 13832 20422 13866
rect 20852 13832 20868 13866
rect 21424 13832 21440 13866
rect 21870 13832 21886 13866
rect 22442 13832 22458 13866
rect 22888 13832 22904 13866
rect 23460 13832 23476 13866
rect 23906 13832 23922 13866
rect 24478 13832 24494 13866
rect 24924 13832 24940 13866
rect 25496 13832 25512 13866
rect 25942 13832 25958 13866
rect 26514 13832 26530 13866
rect 26960 13832 26976 13866
rect 27532 13832 27548 13866
rect 27978 13832 27994 13866
rect 28550 13832 28566 13866
rect 28996 13832 29012 13866
rect 29568 13832 29584 13866
rect 30014 13832 30030 13866
rect 30586 13832 30602 13866
rect 31032 13832 31048 13866
rect 31604 13832 31620 13866
rect 32050 13832 32066 13866
rect 32622 13832 32638 13866
rect 33068 13832 33084 13866
rect 33640 13832 33656 13866
rect 13726 13724 13742 13758
rect 14298 13724 14314 13758
rect 14744 13724 14760 13758
rect 15316 13724 15332 13758
rect 15762 13724 15778 13758
rect 16334 13724 16350 13758
rect 16780 13724 16796 13758
rect 17352 13724 17368 13758
rect 17798 13724 17814 13758
rect 18370 13724 18386 13758
rect 18816 13724 18832 13758
rect 19388 13724 19404 13758
rect 19834 13724 19850 13758
rect 20406 13724 20422 13758
rect 20852 13724 20868 13758
rect 21424 13724 21440 13758
rect 21870 13724 21886 13758
rect 22442 13724 22458 13758
rect 22888 13724 22904 13758
rect 23460 13724 23476 13758
rect 23906 13724 23922 13758
rect 24478 13724 24494 13758
rect 24924 13724 24940 13758
rect 25496 13724 25512 13758
rect 25942 13724 25958 13758
rect 26514 13724 26530 13758
rect 26960 13724 26976 13758
rect 27532 13724 27548 13758
rect 27978 13724 27994 13758
rect 28550 13724 28566 13758
rect 28996 13724 29012 13758
rect 29568 13724 29584 13758
rect 30014 13724 30030 13758
rect 30586 13724 30602 13758
rect 31032 13724 31048 13758
rect 31604 13724 31620 13758
rect 32050 13724 32066 13758
rect 32622 13724 32638 13758
rect 33068 13724 33084 13758
rect 33640 13724 33656 13758
rect 10890 13424 10924 13440
rect 13494 13674 13528 13690
rect 1704 13336 1786 13360
rect 1960 13356 1976 13390
rect 2532 13356 2548 13390
rect 1704 13302 1728 13336
rect 1762 13302 1786 13336
rect 1704 13278 1786 13302
rect 2722 13336 2804 13360
rect 2978 13356 2994 13390
rect 3550 13356 3566 13390
rect 2722 13302 2746 13336
rect 2780 13302 2804 13336
rect 1960 13248 1976 13282
rect 2532 13248 2548 13282
rect 2722 13278 2804 13302
rect 3740 13336 3822 13360
rect 3996 13356 4012 13390
rect 4568 13356 4584 13390
rect 3740 13302 3764 13336
rect 3798 13302 3822 13336
rect 2978 13248 2994 13282
rect 3550 13248 3566 13282
rect 3740 13278 3822 13302
rect 4758 13336 4840 13360
rect 5014 13356 5030 13390
rect 5586 13356 5602 13390
rect 4758 13302 4782 13336
rect 4816 13302 4840 13336
rect 3996 13248 4012 13282
rect 4568 13248 4584 13282
rect 4758 13278 4840 13302
rect 5776 13336 5858 13360
rect 6032 13356 6048 13390
rect 6604 13356 6620 13390
rect 5776 13302 5800 13336
rect 5834 13302 5858 13336
rect 5014 13248 5030 13282
rect 5586 13248 5602 13282
rect 5776 13278 5858 13302
rect 6794 13336 6876 13360
rect 7050 13356 7066 13390
rect 7622 13356 7638 13390
rect 6794 13302 6818 13336
rect 6852 13302 6876 13336
rect 6032 13248 6048 13282
rect 6604 13248 6620 13282
rect 6794 13278 6876 13302
rect 7812 13336 7894 13360
rect 8068 13356 8084 13390
rect 8640 13356 8656 13390
rect 7812 13302 7836 13336
rect 7870 13302 7894 13336
rect 7050 13248 7066 13282
rect 7622 13248 7638 13282
rect 7812 13278 7894 13302
rect 8830 13336 8912 13360
rect 9086 13356 9102 13390
rect 9658 13356 9674 13390
rect 8830 13302 8854 13336
rect 8888 13302 8912 13336
rect 8068 13248 8084 13282
rect 8640 13248 8656 13282
rect 8830 13278 8912 13302
rect 9848 13336 9930 13360
rect 10104 13356 10120 13390
rect 10676 13356 10692 13390
rect 9848 13302 9872 13336
rect 9906 13302 9930 13336
rect 9086 13248 9102 13282
rect 9658 13248 9674 13282
rect 9848 13278 9930 13302
rect 10876 13336 10958 13360
rect 10876 13302 10900 13336
rect 10934 13302 10958 13336
rect 10104 13248 10120 13282
rect 10676 13248 10692 13282
rect 10876 13278 10958 13302
rect 7320 13246 7380 13248
rect 1728 13198 1762 13214
rect 1728 12606 1762 12622
rect 2746 13198 2780 13214
rect 2746 12606 2780 12622
rect 3764 13198 3798 13214
rect 3764 12606 3798 12622
rect 4782 13198 4816 13214
rect 4782 12606 4816 12622
rect 5800 13198 5834 13214
rect 5800 12606 5834 12622
rect 6818 13198 6852 13214
rect 6818 12606 6852 12622
rect 7836 13198 7870 13214
rect 7836 12606 7870 12622
rect 8854 13198 8888 13214
rect 8854 12606 8888 12622
rect 9872 13198 9906 13214
rect 9872 12606 9906 12622
rect 10890 13198 10924 13214
rect 13494 13082 13528 13098
rect 14512 13674 14546 13690
rect 14512 13082 14546 13098
rect 15530 13674 15564 13690
rect 15530 13082 15564 13098
rect 16548 13674 16582 13690
rect 16548 13082 16582 13098
rect 17566 13674 17600 13690
rect 17566 13082 17600 13098
rect 18584 13674 18618 13690
rect 18584 13082 18618 13098
rect 19602 13674 19636 13690
rect 19602 13082 19636 13098
rect 20620 13674 20654 13690
rect 20620 13082 20654 13098
rect 21638 13674 21672 13690
rect 21638 13082 21672 13098
rect 22656 13674 22690 13690
rect 22656 13082 22690 13098
rect 23674 13674 23708 13690
rect 23674 13082 23708 13098
rect 24692 13674 24726 13690
rect 24692 13082 24726 13098
rect 25710 13674 25744 13690
rect 25710 13082 25744 13098
rect 26728 13674 26762 13690
rect 26728 13082 26762 13098
rect 27746 13674 27780 13690
rect 27746 13082 27780 13098
rect 28764 13674 28798 13690
rect 28764 13082 28798 13098
rect 29782 13674 29816 13690
rect 29782 13082 29816 13098
rect 30800 13674 30834 13690
rect 30800 13082 30834 13098
rect 31818 13674 31852 13690
rect 31818 13082 31852 13098
rect 32836 13674 32870 13690
rect 32836 13082 32870 13098
rect 33854 13674 33888 13690
rect 33854 13082 33888 13098
rect 13726 13014 13742 13048
rect 14298 13014 14314 13048
rect 14744 13014 14760 13048
rect 15316 13014 15332 13048
rect 15762 13014 15778 13048
rect 16334 13014 16350 13048
rect 16780 13014 16796 13048
rect 17352 13014 17368 13048
rect 17798 13014 17814 13048
rect 18370 13014 18386 13048
rect 18816 13014 18832 13048
rect 19388 13014 19404 13048
rect 19834 13014 19850 13048
rect 20406 13014 20422 13048
rect 20852 13014 20868 13048
rect 21424 13014 21440 13048
rect 21870 13014 21886 13048
rect 22442 13014 22458 13048
rect 22888 13014 22904 13048
rect 23460 13014 23476 13048
rect 23906 13014 23922 13048
rect 24478 13014 24494 13048
rect 24924 13014 24940 13048
rect 25496 13014 25512 13048
rect 25942 13014 25958 13048
rect 26514 13014 26530 13048
rect 26960 13014 26976 13048
rect 27532 13014 27548 13048
rect 27978 13014 27994 13048
rect 28550 13014 28566 13048
rect 28996 13014 29012 13048
rect 29568 13014 29584 13048
rect 30014 13014 30030 13048
rect 30586 13014 30602 13048
rect 31032 13014 31048 13048
rect 31604 13014 31620 13048
rect 32050 13014 32066 13048
rect 32622 13014 32638 13048
rect 33068 13014 33084 13048
rect 33640 13014 33656 13048
rect 14010 12730 14092 12754
rect 14010 12696 14034 12730
rect 14068 12696 14092 12730
rect 14010 12672 14092 12696
rect 15028 12730 15110 12754
rect 15028 12696 15052 12730
rect 15086 12696 15110 12730
rect 15028 12672 15110 12696
rect 16046 12730 16128 12754
rect 16046 12696 16070 12730
rect 16104 12696 16128 12730
rect 16046 12672 16128 12696
rect 17064 12730 17146 12754
rect 17064 12696 17088 12730
rect 17122 12696 17146 12730
rect 17064 12672 17146 12696
rect 18082 12730 18164 12754
rect 18082 12696 18106 12730
rect 18140 12696 18164 12730
rect 18082 12672 18164 12696
rect 19100 12730 19182 12754
rect 19100 12696 19124 12730
rect 19158 12696 19182 12730
rect 19100 12672 19182 12696
rect 20118 12730 20200 12754
rect 20118 12696 20142 12730
rect 20176 12696 20200 12730
rect 20118 12672 20200 12696
rect 21136 12730 21218 12754
rect 21136 12696 21160 12730
rect 21194 12696 21218 12730
rect 21136 12672 21218 12696
rect 22154 12730 22236 12754
rect 22154 12696 22178 12730
rect 22212 12696 22236 12730
rect 22154 12672 22236 12696
rect 23172 12730 23254 12754
rect 23172 12696 23196 12730
rect 23230 12696 23254 12730
rect 23172 12672 23254 12696
rect 24190 12730 24272 12754
rect 24190 12696 24214 12730
rect 24248 12696 24272 12730
rect 24190 12672 24272 12696
rect 25208 12730 25290 12754
rect 25208 12696 25232 12730
rect 25266 12696 25290 12730
rect 25208 12672 25290 12696
rect 26226 12730 26308 12754
rect 26226 12696 26250 12730
rect 26284 12696 26308 12730
rect 26226 12672 26308 12696
rect 27244 12730 27326 12754
rect 27244 12696 27268 12730
rect 27302 12696 27326 12730
rect 27244 12672 27326 12696
rect 28262 12730 28344 12754
rect 28262 12696 28286 12730
rect 28320 12696 28344 12730
rect 28262 12672 28344 12696
rect 29280 12730 29362 12754
rect 29280 12696 29304 12730
rect 29338 12696 29362 12730
rect 29280 12672 29362 12696
rect 30298 12730 30380 12754
rect 30298 12696 30322 12730
rect 30356 12696 30380 12730
rect 30298 12672 30380 12696
rect 31316 12730 31398 12754
rect 31316 12696 31340 12730
rect 31374 12696 31398 12730
rect 31316 12672 31398 12696
rect 32334 12730 32416 12754
rect 32334 12696 32358 12730
rect 32392 12696 32416 12730
rect 32334 12672 32416 12696
rect 33352 12730 33434 12754
rect 33352 12696 33376 12730
rect 33410 12696 33434 12730
rect 33352 12672 33434 12696
rect 10890 12606 10924 12622
rect 3252 12572 3312 12574
rect 4266 12572 4326 12574
rect 8340 12572 8400 12574
rect 9356 12572 9416 12574
rect 1704 12518 1786 12542
rect 1960 12538 1976 12572
rect 2532 12538 2548 12572
rect 1704 12484 1728 12518
rect 1762 12484 1786 12518
rect 1704 12460 1786 12484
rect 2722 12518 2804 12542
rect 2978 12538 2994 12572
rect 3550 12538 3566 12572
rect 2722 12484 2746 12518
rect 2780 12484 2804 12518
rect 1960 12430 1976 12464
rect 2532 12430 2548 12464
rect 2722 12460 2804 12484
rect 3740 12518 3822 12542
rect 3996 12538 4012 12572
rect 4568 12538 4584 12572
rect 3740 12484 3764 12518
rect 3798 12484 3822 12518
rect 2978 12430 2994 12464
rect 3550 12430 3566 12464
rect 3740 12460 3822 12484
rect 4758 12518 4840 12542
rect 5014 12538 5030 12572
rect 5586 12538 5602 12572
rect 4758 12484 4782 12518
rect 4816 12484 4840 12518
rect 3996 12430 4012 12464
rect 4568 12430 4584 12464
rect 4758 12460 4840 12484
rect 5776 12518 5858 12542
rect 6032 12538 6048 12572
rect 6604 12538 6620 12572
rect 5776 12484 5800 12518
rect 5834 12484 5858 12518
rect 5014 12430 5030 12464
rect 5586 12430 5602 12464
rect 5776 12460 5858 12484
rect 6794 12518 6876 12542
rect 7050 12538 7066 12572
rect 7622 12538 7638 12572
rect 6794 12484 6818 12518
rect 6852 12484 6876 12518
rect 6032 12430 6048 12464
rect 6604 12430 6620 12464
rect 6794 12460 6876 12484
rect 7812 12518 7894 12542
rect 8068 12538 8084 12572
rect 8640 12538 8656 12572
rect 7812 12484 7836 12518
rect 7870 12484 7894 12518
rect 7050 12430 7066 12464
rect 7622 12430 7638 12464
rect 7812 12460 7894 12484
rect 8830 12518 8912 12542
rect 9086 12538 9102 12572
rect 9658 12538 9674 12572
rect 8830 12484 8854 12518
rect 8888 12484 8912 12518
rect 8068 12430 8084 12464
rect 8640 12430 8656 12464
rect 8830 12460 8912 12484
rect 9848 12518 9930 12542
rect 10104 12538 10120 12572
rect 10676 12538 10692 12572
rect 9848 12484 9872 12518
rect 9906 12484 9930 12518
rect 9086 12430 9102 12464
rect 9658 12430 9674 12464
rect 9848 12460 9930 12484
rect 10876 12518 10958 12542
rect 10876 12484 10900 12518
rect 10934 12484 10958 12518
rect 10104 12430 10120 12464
rect 10676 12430 10692 12464
rect 10876 12460 10958 12484
rect 1728 12380 1762 12396
rect 1728 11788 1762 11804
rect 2746 12380 2780 12396
rect 2746 11788 2780 11804
rect 3764 12380 3798 12396
rect 3764 11788 3798 11804
rect 4782 12380 4816 12396
rect 4782 11788 4816 11804
rect 5800 12380 5834 12396
rect 5800 11788 5834 11804
rect 6818 12380 6852 12396
rect 6818 11788 6852 11804
rect 7836 12380 7870 12396
rect 7836 11788 7870 11804
rect 8854 12380 8888 12396
rect 8854 11788 8888 11804
rect 9872 12380 9906 12396
rect 9872 11788 9906 11804
rect 10890 12380 10924 12396
rect 13726 12346 13742 12380
rect 14298 12346 14314 12380
rect 14744 12346 14760 12380
rect 15316 12346 15332 12380
rect 15762 12346 15778 12380
rect 16334 12346 16350 12380
rect 16780 12346 16796 12380
rect 17352 12346 17368 12380
rect 17798 12346 17814 12380
rect 18370 12346 18386 12380
rect 18816 12346 18832 12380
rect 19388 12346 19404 12380
rect 19834 12346 19850 12380
rect 20406 12346 20422 12380
rect 20852 12346 20868 12380
rect 21424 12346 21440 12380
rect 21870 12346 21886 12380
rect 22442 12346 22458 12380
rect 22888 12346 22904 12380
rect 23460 12346 23476 12380
rect 23906 12346 23922 12380
rect 24478 12346 24494 12380
rect 24924 12346 24940 12380
rect 25496 12346 25512 12380
rect 25942 12346 25958 12380
rect 26514 12346 26530 12380
rect 26960 12346 26976 12380
rect 27532 12346 27548 12380
rect 27978 12346 27994 12380
rect 28550 12346 28566 12380
rect 28996 12346 29012 12380
rect 29568 12346 29584 12380
rect 30014 12346 30030 12380
rect 30586 12346 30602 12380
rect 31032 12346 31048 12380
rect 31604 12346 31620 12380
rect 32050 12346 32066 12380
rect 32622 12346 32638 12380
rect 33068 12346 33084 12380
rect 33640 12346 33656 12380
rect 23150 12340 23210 12346
rect 10890 11788 10924 11804
rect 13494 12296 13528 12312
rect 3256 11754 3316 11756
rect 4270 11754 4330 11756
rect 8344 11754 8404 11756
rect 9360 11754 9420 11756
rect 1704 11700 1786 11724
rect 1960 11720 1976 11754
rect 2532 11720 2548 11754
rect 1704 11666 1728 11700
rect 1762 11666 1786 11700
rect 1704 11642 1786 11666
rect 2722 11700 2804 11724
rect 2978 11720 2994 11754
rect 3550 11720 3566 11754
rect 2722 11666 2746 11700
rect 2780 11666 2804 11700
rect 1960 11612 1976 11646
rect 2532 11612 2548 11646
rect 2722 11642 2804 11666
rect 3740 11700 3822 11724
rect 3996 11720 4012 11754
rect 4568 11720 4584 11754
rect 3740 11666 3764 11700
rect 3798 11666 3822 11700
rect 2978 11612 2994 11646
rect 3550 11612 3566 11646
rect 3740 11642 3822 11666
rect 4758 11700 4840 11724
rect 5014 11720 5030 11754
rect 5586 11720 5602 11754
rect 4758 11666 4782 11700
rect 4816 11666 4840 11700
rect 3996 11612 4012 11646
rect 4568 11612 4584 11646
rect 4758 11642 4840 11666
rect 5776 11700 5858 11724
rect 6032 11720 6048 11754
rect 6604 11720 6620 11754
rect 5776 11666 5800 11700
rect 5834 11666 5858 11700
rect 5014 11612 5030 11646
rect 5586 11612 5602 11646
rect 5776 11642 5858 11666
rect 6794 11700 6876 11724
rect 7050 11720 7066 11754
rect 7622 11720 7638 11754
rect 6794 11666 6818 11700
rect 6852 11666 6876 11700
rect 6032 11612 6048 11646
rect 6604 11612 6620 11646
rect 6794 11642 6876 11666
rect 7812 11700 7894 11724
rect 8068 11720 8084 11754
rect 8640 11720 8656 11754
rect 7812 11666 7836 11700
rect 7870 11666 7894 11700
rect 7050 11612 7066 11646
rect 7622 11612 7638 11646
rect 7812 11642 7894 11666
rect 8830 11700 8912 11724
rect 9086 11720 9102 11754
rect 9658 11720 9674 11754
rect 8830 11666 8854 11700
rect 8888 11666 8912 11700
rect 8068 11612 8084 11646
rect 8640 11612 8656 11646
rect 8830 11642 8912 11666
rect 9848 11700 9930 11724
rect 10104 11720 10120 11754
rect 10676 11720 10692 11754
rect 9848 11666 9872 11700
rect 9906 11666 9930 11700
rect 9086 11612 9102 11646
rect 9658 11612 9674 11646
rect 9848 11642 9930 11666
rect 10876 11700 10958 11724
rect 13494 11704 13528 11720
rect 14512 12296 14546 12312
rect 14512 11704 14546 11720
rect 15530 12296 15564 12312
rect 15530 11704 15564 11720
rect 16548 12296 16582 12312
rect 16548 11704 16582 11720
rect 17566 12296 17600 12312
rect 17566 11704 17600 11720
rect 18584 12296 18618 12312
rect 18584 11704 18618 11720
rect 19602 12296 19636 12312
rect 19602 11704 19636 11720
rect 20620 12296 20654 12312
rect 20620 11704 20654 11720
rect 21638 12296 21672 12312
rect 21638 11704 21672 11720
rect 22656 12296 22690 12312
rect 22656 11704 22690 11720
rect 23674 12296 23708 12312
rect 23674 11704 23708 11720
rect 24692 12296 24726 12312
rect 24692 11704 24726 11720
rect 25710 12296 25744 12312
rect 25710 11704 25744 11720
rect 26728 12296 26762 12312
rect 26728 11704 26762 11720
rect 27746 12296 27780 12312
rect 27746 11704 27780 11720
rect 28764 12296 28798 12312
rect 28764 11704 28798 11720
rect 29782 12296 29816 12312
rect 29782 11704 29816 11720
rect 30800 12296 30834 12312
rect 30800 11704 30834 11720
rect 31818 12296 31852 12312
rect 31818 11704 31852 11720
rect 32836 12296 32870 12312
rect 32836 11704 32870 11720
rect 33854 12296 33888 12312
rect 33854 11704 33888 11720
rect 10876 11666 10900 11700
rect 10934 11666 10958 11700
rect 19078 11670 19138 11676
rect 21114 11670 21174 11676
rect 22134 11670 22194 11676
rect 27206 11670 27266 11676
rect 10104 11612 10120 11646
rect 10676 11612 10692 11646
rect 10876 11642 10958 11666
rect 13726 11636 13742 11670
rect 14298 11636 14314 11670
rect 14744 11636 14760 11670
rect 15316 11636 15332 11670
rect 15762 11636 15778 11670
rect 16334 11636 16350 11670
rect 16780 11636 16796 11670
rect 17352 11636 17368 11670
rect 17798 11636 17814 11670
rect 18370 11636 18386 11670
rect 18816 11636 18832 11670
rect 19388 11636 19404 11670
rect 19834 11636 19850 11670
rect 20406 11636 20422 11670
rect 20852 11636 20868 11670
rect 21424 11636 21440 11670
rect 21870 11636 21886 11670
rect 22442 11636 22458 11670
rect 22888 11636 22904 11670
rect 23460 11636 23476 11670
rect 23906 11636 23922 11670
rect 24478 11636 24494 11670
rect 24924 11636 24940 11670
rect 25496 11636 25512 11670
rect 25942 11636 25958 11670
rect 26514 11636 26530 11670
rect 26960 11636 26976 11670
rect 27532 11636 27548 11670
rect 27978 11636 27994 11670
rect 28550 11636 28566 11670
rect 28996 11636 29012 11670
rect 29568 11636 29584 11670
rect 30014 11636 30030 11670
rect 30586 11636 30602 11670
rect 31032 11636 31048 11670
rect 31604 11636 31620 11670
rect 32050 11636 32066 11670
rect 32622 11636 32638 11670
rect 33068 11636 33084 11670
rect 33640 11636 33656 11670
rect 1728 11562 1762 11578
rect 1728 10970 1762 10986
rect 2746 11562 2780 11578
rect 2746 10970 2780 10986
rect 3764 11562 3798 11578
rect 3764 10970 3798 10986
rect 4782 11562 4816 11578
rect 4782 10970 4816 10986
rect 5800 11562 5834 11578
rect 5800 10970 5834 10986
rect 6818 11562 6852 11578
rect 6818 10970 6852 10986
rect 7836 11562 7870 11578
rect 7836 10970 7870 10986
rect 8854 11562 8888 11578
rect 8854 10970 8888 10986
rect 9872 11562 9906 11578
rect 9872 10970 9906 10986
rect 10890 11562 10924 11578
rect 13998 11424 14080 11448
rect 13998 11390 14022 11424
rect 14056 11390 14080 11424
rect 13998 11366 14080 11390
rect 15016 11424 15098 11448
rect 15016 11390 15040 11424
rect 15074 11390 15098 11424
rect 15016 11366 15098 11390
rect 16034 11424 16116 11448
rect 16034 11390 16058 11424
rect 16092 11390 16116 11424
rect 16034 11366 16116 11390
rect 17052 11424 17134 11448
rect 17052 11390 17076 11424
rect 17110 11390 17134 11424
rect 17052 11366 17134 11390
rect 18070 11424 18152 11448
rect 18070 11390 18094 11424
rect 18128 11390 18152 11424
rect 18070 11366 18152 11390
rect 19088 11424 19170 11448
rect 19088 11390 19112 11424
rect 19146 11390 19170 11424
rect 19088 11366 19170 11390
rect 20106 11424 20188 11448
rect 20106 11390 20130 11424
rect 20164 11390 20188 11424
rect 20106 11366 20188 11390
rect 21124 11424 21206 11448
rect 21124 11390 21148 11424
rect 21182 11390 21206 11424
rect 21124 11366 21206 11390
rect 22142 11424 22224 11448
rect 22142 11390 22166 11424
rect 22200 11390 22224 11424
rect 22142 11366 22224 11390
rect 23160 11424 23242 11448
rect 23160 11390 23184 11424
rect 23218 11390 23242 11424
rect 23160 11366 23242 11390
rect 24178 11424 24260 11448
rect 24178 11390 24202 11424
rect 24236 11390 24260 11424
rect 24178 11366 24260 11390
rect 25196 11424 25278 11448
rect 25196 11390 25220 11424
rect 25254 11390 25278 11424
rect 25196 11366 25278 11390
rect 26214 11424 26296 11448
rect 26214 11390 26238 11424
rect 26272 11390 26296 11424
rect 26214 11366 26296 11390
rect 27232 11424 27314 11448
rect 27232 11390 27256 11424
rect 27290 11390 27314 11424
rect 27232 11366 27314 11390
rect 28250 11424 28332 11448
rect 28250 11390 28274 11424
rect 28308 11390 28332 11424
rect 28250 11366 28332 11390
rect 29268 11424 29350 11448
rect 29268 11390 29292 11424
rect 29326 11390 29350 11424
rect 29268 11366 29350 11390
rect 30286 11424 30368 11448
rect 30286 11390 30310 11424
rect 30344 11390 30368 11424
rect 30286 11366 30368 11390
rect 31304 11424 31386 11448
rect 31304 11390 31328 11424
rect 31362 11390 31386 11424
rect 31304 11366 31386 11390
rect 32322 11424 32404 11448
rect 32322 11390 32346 11424
rect 32380 11390 32404 11424
rect 32322 11366 32404 11390
rect 33340 11424 33422 11448
rect 33340 11390 33364 11424
rect 33398 11390 33422 11424
rect 33340 11366 33422 11390
rect 13726 11114 13742 11148
rect 14298 11114 14314 11148
rect 14744 11114 14760 11148
rect 15316 11114 15332 11148
rect 15762 11114 15778 11148
rect 16334 11114 16350 11148
rect 16780 11114 16796 11148
rect 17352 11114 17368 11148
rect 17798 11114 17814 11148
rect 18370 11114 18386 11148
rect 18816 11114 18832 11148
rect 19388 11114 19404 11148
rect 19834 11114 19850 11148
rect 20406 11114 20422 11148
rect 20852 11114 20868 11148
rect 21424 11114 21440 11148
rect 21870 11114 21886 11148
rect 22442 11114 22458 11148
rect 22888 11114 22904 11148
rect 23460 11114 23476 11148
rect 23906 11114 23922 11148
rect 24478 11114 24494 11148
rect 24924 11114 24940 11148
rect 25496 11114 25512 11148
rect 25942 11114 25958 11148
rect 26514 11114 26530 11148
rect 26960 11114 26976 11148
rect 27532 11114 27548 11148
rect 27978 11114 27994 11148
rect 28550 11114 28566 11148
rect 28996 11114 29012 11148
rect 29568 11114 29584 11148
rect 30014 11114 30030 11148
rect 30586 11114 30602 11148
rect 31032 11114 31048 11148
rect 31604 11114 31620 11148
rect 32050 11114 32066 11148
rect 32622 11114 32638 11148
rect 33068 11114 33084 11148
rect 33640 11114 33656 11148
rect 15012 11110 15072 11114
rect 16028 11110 16088 11114
rect 20104 11106 20164 11114
rect 24170 11110 24230 11114
rect 26204 11110 26264 11114
rect 32316 11110 32376 11114
rect 10890 10970 10924 10986
rect 13494 11064 13528 11080
rect 1704 10882 1786 10906
rect 1960 10902 1976 10936
rect 2532 10902 2548 10936
rect 1704 10848 1728 10882
rect 1762 10848 1786 10882
rect 1704 10824 1786 10848
rect 2722 10882 2804 10906
rect 2978 10902 2994 10936
rect 3550 10902 3566 10936
rect 2722 10848 2746 10882
rect 2780 10848 2804 10882
rect 1960 10794 1976 10828
rect 2532 10794 2548 10828
rect 2722 10824 2804 10848
rect 3740 10882 3822 10906
rect 3996 10902 4012 10936
rect 4568 10902 4584 10936
rect 3740 10848 3764 10882
rect 3798 10848 3822 10882
rect 2978 10794 2994 10828
rect 3550 10794 3566 10828
rect 3740 10824 3822 10848
rect 4758 10882 4840 10906
rect 5014 10902 5030 10936
rect 5586 10902 5602 10936
rect 4758 10848 4782 10882
rect 4816 10848 4840 10882
rect 3996 10794 4012 10828
rect 4568 10794 4584 10828
rect 4758 10824 4840 10848
rect 5776 10882 5858 10906
rect 6032 10902 6048 10936
rect 6604 10902 6620 10936
rect 5776 10848 5800 10882
rect 5834 10848 5858 10882
rect 5014 10794 5030 10828
rect 5586 10794 5602 10828
rect 5776 10824 5858 10848
rect 6794 10882 6876 10906
rect 7050 10902 7066 10936
rect 7622 10902 7638 10936
rect 6794 10848 6818 10882
rect 6852 10848 6876 10882
rect 6032 10794 6048 10828
rect 6604 10794 6620 10828
rect 6794 10824 6876 10848
rect 7812 10882 7894 10906
rect 8068 10902 8084 10936
rect 8640 10902 8656 10936
rect 7812 10848 7836 10882
rect 7870 10848 7894 10882
rect 7050 10794 7066 10828
rect 7622 10794 7638 10828
rect 7812 10824 7894 10848
rect 8830 10882 8912 10906
rect 9086 10902 9102 10936
rect 9658 10902 9674 10936
rect 8830 10848 8854 10882
rect 8888 10848 8912 10882
rect 8068 10794 8084 10828
rect 8640 10794 8656 10828
rect 8830 10824 8912 10848
rect 9848 10882 9930 10906
rect 10104 10902 10120 10936
rect 10676 10902 10692 10936
rect 9848 10848 9872 10882
rect 9906 10848 9930 10882
rect 9086 10794 9102 10828
rect 9658 10794 9674 10828
rect 9848 10824 9930 10848
rect 10876 10882 10958 10906
rect 10876 10848 10900 10882
rect 10934 10848 10958 10882
rect 10104 10794 10120 10828
rect 10676 10794 10692 10828
rect 10876 10824 10958 10848
rect 7316 10792 7376 10794
rect 1728 10744 1762 10760
rect 1728 10152 1762 10168
rect 2746 10744 2780 10760
rect 2746 10152 2780 10168
rect 3764 10744 3798 10760
rect 3764 10152 3798 10168
rect 4782 10744 4816 10760
rect 4782 10152 4816 10168
rect 5800 10744 5834 10760
rect 5800 10152 5834 10168
rect 6818 10744 6852 10760
rect 6818 10152 6852 10168
rect 7836 10744 7870 10760
rect 7836 10152 7870 10168
rect 8854 10744 8888 10760
rect 8854 10152 8888 10168
rect 9872 10744 9906 10760
rect 9872 10152 9906 10168
rect 10890 10744 10924 10760
rect 13494 10472 13528 10488
rect 14512 11064 14546 11080
rect 14512 10472 14546 10488
rect 15530 11064 15564 11080
rect 15530 10472 15564 10488
rect 16548 11064 16582 11080
rect 16548 10472 16582 10488
rect 17566 11064 17600 11080
rect 17566 10472 17600 10488
rect 18584 11064 18618 11080
rect 18584 10472 18618 10488
rect 19602 11064 19636 11080
rect 19602 10472 19636 10488
rect 20620 11064 20654 11080
rect 20620 10472 20654 10488
rect 21638 11064 21672 11080
rect 21638 10472 21672 10488
rect 22656 11064 22690 11080
rect 22656 10472 22690 10488
rect 23674 11064 23708 11080
rect 23674 10472 23708 10488
rect 24692 11064 24726 11080
rect 24692 10472 24726 10488
rect 25710 11064 25744 11080
rect 25710 10472 25744 10488
rect 26728 11064 26762 11080
rect 26728 10472 26762 10488
rect 27746 11064 27780 11080
rect 27746 10472 27780 10488
rect 28764 11064 28798 11080
rect 28764 10472 28798 10488
rect 29782 11064 29816 11080
rect 29782 10472 29816 10488
rect 30800 11064 30834 11080
rect 30800 10472 30834 10488
rect 31818 11064 31852 11080
rect 31818 10472 31852 10488
rect 32836 11064 32870 11080
rect 32836 10472 32870 10488
rect 33854 11064 33888 11080
rect 33888 10488 33894 10536
rect 33854 10472 33888 10488
rect 17038 10438 17098 10440
rect 13726 10404 13742 10438
rect 14298 10404 14314 10438
rect 14744 10404 14760 10438
rect 15316 10404 15332 10438
rect 15762 10404 15778 10438
rect 16334 10404 16350 10438
rect 16780 10404 16796 10438
rect 17352 10404 17368 10438
rect 17798 10404 17814 10438
rect 18370 10404 18386 10438
rect 18816 10404 18832 10438
rect 19388 10404 19404 10438
rect 19834 10404 19850 10438
rect 20406 10404 20422 10438
rect 20852 10404 20868 10438
rect 21424 10404 21440 10438
rect 21870 10404 21886 10438
rect 22442 10404 22458 10438
rect 22888 10404 22904 10438
rect 23460 10404 23476 10438
rect 23906 10404 23922 10438
rect 24478 10404 24494 10438
rect 24924 10404 24940 10438
rect 25496 10404 25512 10438
rect 25942 10404 25958 10438
rect 26514 10404 26530 10438
rect 26960 10404 26976 10438
rect 27532 10404 27548 10438
rect 27978 10404 27994 10438
rect 28550 10404 28566 10438
rect 28996 10404 29012 10438
rect 29568 10404 29584 10438
rect 30014 10404 30030 10438
rect 30586 10404 30602 10438
rect 31032 10404 31048 10438
rect 31604 10404 31620 10438
rect 32050 10404 32066 10438
rect 32622 10404 32638 10438
rect 33068 10404 33084 10438
rect 33640 10404 33656 10438
rect 19072 10400 19132 10404
rect 28230 10390 28290 10404
rect 29264 10390 29324 10404
rect 10890 10152 10924 10168
rect 13986 10188 14068 10212
rect 13986 10154 14010 10188
rect 14044 10154 14068 10188
rect 13986 10130 14068 10154
rect 15004 10188 15086 10212
rect 15004 10154 15028 10188
rect 15062 10154 15086 10188
rect 15004 10130 15086 10154
rect 16022 10188 16104 10212
rect 16022 10154 16046 10188
rect 16080 10154 16104 10188
rect 16022 10130 16104 10154
rect 17040 10188 17122 10212
rect 17040 10154 17064 10188
rect 17098 10154 17122 10188
rect 17040 10130 17122 10154
rect 18058 10188 18140 10212
rect 18058 10154 18082 10188
rect 18116 10154 18140 10188
rect 18058 10130 18140 10154
rect 19076 10188 19158 10212
rect 19076 10154 19100 10188
rect 19134 10154 19158 10188
rect 19076 10130 19158 10154
rect 20094 10188 20176 10212
rect 20094 10154 20118 10188
rect 20152 10154 20176 10188
rect 20094 10130 20176 10154
rect 21112 10188 21194 10212
rect 21112 10154 21136 10188
rect 21170 10154 21194 10188
rect 21112 10130 21194 10154
rect 22130 10188 22212 10212
rect 22130 10154 22154 10188
rect 22188 10154 22212 10188
rect 22130 10130 22212 10154
rect 23148 10188 23230 10212
rect 23148 10154 23172 10188
rect 23206 10154 23230 10188
rect 23148 10130 23230 10154
rect 24166 10188 24248 10212
rect 24166 10154 24190 10188
rect 24224 10154 24248 10188
rect 24166 10130 24248 10154
rect 25184 10188 25266 10212
rect 25184 10154 25208 10188
rect 25242 10154 25266 10188
rect 25184 10130 25266 10154
rect 26202 10188 26284 10212
rect 26202 10154 26226 10188
rect 26260 10154 26284 10188
rect 26202 10130 26284 10154
rect 27220 10188 27302 10212
rect 27220 10154 27244 10188
rect 27278 10154 27302 10188
rect 27220 10130 27302 10154
rect 28238 10188 28320 10212
rect 28238 10154 28262 10188
rect 28296 10154 28320 10188
rect 28238 10130 28320 10154
rect 29256 10188 29338 10212
rect 29256 10154 29280 10188
rect 29314 10154 29338 10188
rect 29256 10130 29338 10154
rect 30274 10188 30356 10212
rect 30274 10154 30298 10188
rect 30332 10154 30356 10188
rect 30274 10130 30356 10154
rect 31292 10188 31374 10212
rect 31292 10154 31316 10188
rect 31350 10154 31374 10188
rect 31292 10130 31374 10154
rect 32310 10188 32392 10212
rect 32310 10154 32334 10188
rect 32368 10154 32392 10188
rect 32310 10130 32392 10154
rect 33328 10188 33410 10212
rect 33328 10154 33352 10188
rect 33386 10154 33410 10188
rect 33328 10130 33410 10154
rect 3242 10118 3302 10120
rect 4256 10118 4316 10120
rect 8330 10118 8390 10120
rect 9346 10118 9406 10120
rect 1704 10064 1786 10088
rect 1960 10084 1976 10118
rect 2532 10084 2548 10118
rect 1704 10030 1728 10064
rect 1762 10030 1786 10064
rect 1704 10006 1786 10030
rect 2722 10064 2804 10088
rect 2978 10084 2994 10118
rect 3550 10084 3566 10118
rect 2722 10030 2746 10064
rect 2780 10030 2804 10064
rect 1960 9976 1976 10010
rect 2532 9976 2548 10010
rect 2722 10006 2804 10030
rect 3740 10064 3822 10088
rect 3996 10084 4012 10118
rect 4568 10084 4584 10118
rect 3740 10030 3764 10064
rect 3798 10030 3822 10064
rect 2978 9976 2994 10010
rect 3550 9976 3566 10010
rect 3740 10006 3822 10030
rect 4758 10064 4840 10088
rect 5014 10084 5030 10118
rect 5586 10084 5602 10118
rect 4758 10030 4782 10064
rect 4816 10030 4840 10064
rect 3996 9976 4012 10010
rect 4568 9976 4584 10010
rect 4758 10006 4840 10030
rect 5776 10064 5858 10088
rect 6032 10084 6048 10118
rect 6604 10084 6620 10118
rect 5776 10030 5800 10064
rect 5834 10030 5858 10064
rect 5014 9976 5030 10010
rect 5586 9976 5602 10010
rect 5776 10006 5858 10030
rect 6794 10064 6876 10088
rect 7050 10084 7066 10118
rect 7622 10084 7638 10118
rect 6794 10030 6818 10064
rect 6852 10030 6876 10064
rect 6032 9976 6048 10010
rect 6604 9976 6620 10010
rect 6794 10006 6876 10030
rect 7812 10064 7894 10088
rect 8068 10084 8084 10118
rect 8640 10084 8656 10118
rect 7812 10030 7836 10064
rect 7870 10030 7894 10064
rect 7050 9976 7066 10010
rect 7622 9976 7638 10010
rect 7812 10006 7894 10030
rect 8830 10064 8912 10088
rect 9086 10084 9102 10118
rect 9658 10084 9674 10118
rect 8830 10030 8854 10064
rect 8888 10030 8912 10064
rect 8068 9976 8084 10010
rect 8640 9976 8656 10010
rect 8830 10006 8912 10030
rect 9848 10064 9930 10088
rect 10104 10084 10120 10118
rect 10676 10084 10692 10118
rect 9848 10030 9872 10064
rect 9906 10030 9930 10064
rect 9086 9976 9102 10010
rect 9658 9976 9674 10010
rect 9848 10006 9930 10030
rect 10876 10064 10958 10088
rect 10876 10030 10900 10064
rect 10934 10030 10958 10064
rect 10104 9976 10120 10010
rect 10676 9976 10692 10010
rect 10876 10006 10958 10030
rect 1728 9926 1762 9942
rect 1728 9334 1762 9350
rect 2746 9926 2780 9942
rect 2746 9334 2780 9350
rect 3764 9926 3798 9942
rect 3764 9334 3798 9350
rect 4782 9926 4816 9942
rect 4782 9334 4816 9350
rect 5800 9926 5834 9942
rect 5800 9334 5834 9350
rect 6818 9926 6852 9942
rect 6818 9334 6852 9350
rect 7836 9926 7870 9942
rect 7836 9334 7870 9350
rect 8854 9926 8888 9942
rect 8854 9334 8888 9350
rect 9872 9926 9906 9942
rect 9872 9334 9906 9350
rect 10890 9926 10924 9942
rect 13724 9880 13740 9914
rect 14296 9880 14312 9914
rect 14742 9880 14758 9914
rect 15314 9880 15330 9914
rect 15760 9880 15776 9914
rect 16332 9880 16348 9914
rect 16778 9880 16794 9914
rect 17350 9880 17366 9914
rect 17796 9880 17812 9914
rect 18368 9880 18384 9914
rect 18814 9880 18830 9914
rect 19386 9880 19402 9914
rect 19832 9880 19848 9914
rect 20404 9880 20420 9914
rect 20850 9880 20866 9914
rect 21422 9880 21438 9914
rect 21868 9880 21884 9914
rect 22440 9880 22456 9914
rect 22886 9880 22902 9914
rect 23458 9880 23474 9914
rect 23904 9880 23920 9914
rect 24476 9880 24492 9914
rect 24922 9880 24938 9914
rect 25494 9880 25510 9914
rect 25940 9880 25956 9914
rect 26512 9880 26528 9914
rect 26958 9880 26974 9914
rect 27530 9880 27546 9914
rect 27976 9880 27992 9914
rect 28548 9880 28564 9914
rect 28994 9880 29010 9914
rect 29566 9880 29582 9914
rect 30012 9880 30028 9914
rect 30584 9880 30600 9914
rect 31030 9880 31046 9914
rect 31602 9880 31618 9914
rect 32048 9880 32064 9914
rect 32620 9880 32636 9914
rect 33066 9880 33082 9914
rect 33638 9880 33654 9914
rect 16034 9876 16094 9880
rect 10890 9334 10924 9350
rect 13492 9830 13526 9846
rect 3246 9300 3306 9302
rect 4260 9300 4320 9302
rect 8334 9300 8394 9302
rect 9350 9300 9410 9302
rect 1704 9246 1786 9270
rect 1960 9266 1976 9300
rect 2532 9266 2548 9300
rect 1704 9212 1728 9246
rect 1762 9212 1786 9246
rect 1704 9188 1786 9212
rect 2722 9246 2804 9270
rect 2978 9266 2994 9300
rect 3550 9266 3566 9300
rect 2722 9212 2746 9246
rect 2780 9212 2804 9246
rect 1960 9158 1976 9192
rect 2532 9158 2548 9192
rect 2722 9188 2804 9212
rect 3740 9246 3822 9270
rect 3996 9266 4012 9300
rect 4568 9266 4584 9300
rect 3740 9212 3764 9246
rect 3798 9212 3822 9246
rect 2978 9158 2994 9192
rect 3550 9158 3566 9192
rect 3740 9188 3822 9212
rect 4758 9246 4840 9270
rect 5014 9266 5030 9300
rect 5586 9266 5602 9300
rect 4758 9212 4782 9246
rect 4816 9212 4840 9246
rect 3996 9158 4012 9192
rect 4568 9158 4584 9192
rect 4758 9188 4840 9212
rect 5776 9246 5858 9270
rect 6032 9266 6048 9300
rect 6604 9266 6620 9300
rect 5776 9212 5800 9246
rect 5834 9212 5858 9246
rect 5014 9158 5030 9192
rect 5586 9158 5602 9192
rect 5776 9188 5858 9212
rect 6794 9246 6876 9270
rect 7050 9266 7066 9300
rect 7622 9266 7638 9300
rect 6794 9212 6818 9246
rect 6852 9212 6876 9246
rect 6032 9158 6048 9192
rect 6604 9158 6620 9192
rect 6794 9188 6876 9212
rect 7812 9246 7894 9270
rect 8068 9266 8084 9300
rect 8640 9266 8656 9300
rect 7812 9212 7836 9246
rect 7870 9212 7894 9246
rect 7050 9158 7066 9192
rect 7622 9158 7638 9192
rect 7812 9188 7894 9212
rect 8830 9246 8912 9270
rect 9086 9266 9102 9300
rect 9658 9266 9674 9300
rect 8830 9212 8854 9246
rect 8888 9212 8912 9246
rect 8068 9158 8084 9192
rect 8640 9158 8656 9192
rect 8830 9188 8912 9212
rect 9848 9246 9930 9270
rect 10104 9266 10120 9300
rect 10676 9266 10692 9300
rect 9848 9212 9872 9246
rect 9906 9212 9930 9246
rect 9086 9158 9102 9192
rect 9658 9158 9674 9192
rect 9848 9188 9930 9212
rect 10876 9246 10958 9270
rect 10876 9212 10900 9246
rect 10934 9212 10958 9246
rect 13492 9238 13526 9254
rect 14510 9830 14544 9846
rect 14510 9238 14544 9254
rect 15528 9830 15562 9846
rect 15528 9238 15562 9254
rect 16546 9830 16580 9846
rect 16546 9238 16580 9254
rect 17564 9830 17598 9846
rect 17564 9238 17598 9254
rect 18582 9830 18616 9846
rect 18582 9238 18616 9254
rect 19600 9830 19634 9846
rect 19600 9238 19634 9254
rect 20618 9830 20652 9846
rect 20618 9238 20652 9254
rect 21636 9830 21670 9846
rect 21636 9238 21670 9254
rect 22654 9830 22688 9846
rect 22654 9238 22688 9254
rect 23672 9830 23706 9846
rect 23672 9238 23706 9254
rect 24690 9830 24724 9846
rect 24690 9238 24724 9254
rect 25708 9830 25742 9846
rect 25708 9238 25742 9254
rect 26726 9830 26760 9846
rect 26726 9238 26760 9254
rect 27744 9830 27778 9846
rect 27744 9238 27778 9254
rect 28762 9830 28796 9846
rect 28762 9238 28796 9254
rect 29780 9830 29814 9846
rect 29780 9238 29814 9254
rect 30798 9830 30832 9846
rect 30798 9238 30832 9254
rect 31816 9830 31850 9846
rect 31816 9238 31850 9254
rect 32834 9830 32868 9846
rect 32834 9238 32868 9254
rect 33852 9830 33886 9846
rect 33852 9238 33886 9254
rect 10104 9158 10120 9192
rect 10676 9158 10692 9192
rect 10876 9188 10958 9212
rect 21102 9204 21162 9208
rect 22130 9204 22190 9206
rect 24174 9204 24234 9208
rect 13724 9170 13740 9204
rect 14296 9170 14312 9204
rect 14742 9170 14758 9204
rect 15314 9170 15330 9204
rect 15760 9170 15776 9204
rect 16332 9170 16348 9204
rect 16778 9170 16794 9204
rect 17350 9170 17366 9204
rect 17796 9170 17812 9204
rect 18368 9170 18384 9204
rect 18814 9170 18830 9204
rect 19386 9170 19402 9204
rect 19832 9170 19848 9204
rect 20404 9170 20420 9204
rect 20850 9170 20866 9204
rect 21422 9170 21438 9204
rect 21868 9170 21884 9204
rect 22440 9170 22456 9204
rect 22886 9170 22902 9204
rect 23458 9170 23474 9204
rect 23904 9170 23920 9204
rect 24476 9170 24492 9204
rect 24922 9170 24938 9204
rect 25494 9170 25510 9204
rect 25940 9170 25956 9204
rect 26512 9170 26528 9204
rect 26958 9170 26974 9204
rect 27530 9170 27546 9204
rect 27976 9170 27992 9204
rect 28548 9170 28564 9204
rect 28994 9170 29010 9204
rect 29566 9170 29582 9204
rect 30012 9170 30028 9204
rect 30584 9170 30600 9204
rect 31030 9170 31046 9204
rect 31602 9170 31618 9204
rect 32048 9170 32064 9204
rect 32620 9170 32636 9204
rect 33066 9170 33082 9204
rect 33638 9170 33654 9204
rect 1728 9108 1762 9124
rect 1728 8516 1762 8532
rect 2746 9108 2780 9124
rect 2746 8516 2780 8532
rect 3764 9108 3798 9124
rect 3764 8516 3798 8532
rect 4782 9108 4816 9124
rect 4782 8516 4816 8532
rect 5800 9108 5834 9124
rect 5800 8516 5834 8532
rect 6818 9108 6852 9124
rect 6818 8516 6852 8532
rect 7836 9108 7870 9124
rect 7836 8516 7870 8532
rect 8854 9108 8888 9124
rect 8854 8516 8888 8532
rect 9872 9108 9906 9124
rect 9872 8516 9906 8532
rect 10890 9108 10924 9124
rect 13986 8964 14068 8988
rect 13986 8930 14010 8964
rect 14044 8930 14068 8964
rect 13986 8906 14068 8930
rect 15004 8964 15086 8988
rect 15004 8930 15028 8964
rect 15062 8930 15086 8964
rect 15004 8906 15086 8930
rect 16022 8964 16104 8988
rect 16022 8930 16046 8964
rect 16080 8930 16104 8964
rect 16022 8906 16104 8930
rect 17040 8964 17122 8988
rect 17040 8930 17064 8964
rect 17098 8930 17122 8964
rect 17040 8906 17122 8930
rect 18058 8964 18140 8988
rect 18058 8930 18082 8964
rect 18116 8930 18140 8964
rect 18058 8906 18140 8930
rect 19076 8964 19158 8988
rect 19076 8930 19100 8964
rect 19134 8930 19158 8964
rect 19076 8906 19158 8930
rect 20094 8964 20176 8988
rect 20094 8930 20118 8964
rect 20152 8930 20176 8964
rect 20094 8906 20176 8930
rect 21112 8964 21194 8988
rect 21112 8930 21136 8964
rect 21170 8930 21194 8964
rect 21112 8906 21194 8930
rect 22130 8964 22212 8988
rect 22130 8930 22154 8964
rect 22188 8930 22212 8964
rect 22130 8906 22212 8930
rect 23148 8964 23230 8988
rect 23148 8930 23172 8964
rect 23206 8930 23230 8964
rect 23148 8906 23230 8930
rect 24166 8964 24248 8988
rect 24166 8930 24190 8964
rect 24224 8930 24248 8964
rect 24166 8906 24248 8930
rect 25184 8964 25266 8988
rect 25184 8930 25208 8964
rect 25242 8930 25266 8964
rect 25184 8906 25266 8930
rect 26202 8964 26284 8988
rect 26202 8930 26226 8964
rect 26260 8930 26284 8964
rect 26202 8906 26284 8930
rect 27220 8964 27302 8988
rect 27220 8930 27244 8964
rect 27278 8930 27302 8964
rect 27220 8906 27302 8930
rect 28238 8964 28320 8988
rect 28238 8930 28262 8964
rect 28296 8930 28320 8964
rect 28238 8906 28320 8930
rect 29256 8964 29338 8988
rect 29256 8930 29280 8964
rect 29314 8930 29338 8964
rect 29256 8906 29338 8930
rect 30274 8964 30356 8988
rect 30274 8930 30298 8964
rect 30332 8930 30356 8964
rect 30274 8906 30356 8930
rect 31292 8964 31374 8988
rect 31292 8930 31316 8964
rect 31350 8930 31374 8964
rect 31292 8906 31374 8930
rect 32310 8964 32392 8988
rect 32310 8930 32334 8964
rect 32368 8930 32392 8964
rect 32310 8906 32392 8930
rect 33328 8964 33410 8988
rect 33328 8930 33352 8964
rect 33386 8930 33410 8964
rect 33328 8906 33410 8930
rect 13724 8646 13740 8680
rect 14296 8646 14312 8680
rect 14742 8646 14758 8680
rect 15314 8646 15330 8680
rect 15760 8646 15776 8680
rect 16332 8646 16348 8680
rect 16778 8646 16794 8680
rect 17350 8646 17366 8680
rect 17796 8646 17812 8680
rect 18368 8646 18384 8680
rect 18814 8646 18830 8680
rect 19386 8646 19402 8680
rect 19832 8646 19848 8680
rect 20404 8646 20420 8680
rect 20850 8646 20866 8680
rect 21422 8646 21438 8680
rect 21868 8646 21884 8680
rect 22440 8646 22456 8680
rect 22886 8646 22902 8680
rect 23458 8646 23474 8680
rect 23904 8646 23920 8680
rect 24476 8646 24492 8680
rect 24922 8646 24938 8680
rect 25494 8646 25510 8680
rect 25940 8646 25956 8680
rect 26512 8646 26528 8680
rect 26958 8646 26974 8680
rect 27530 8646 27546 8680
rect 27976 8646 27992 8680
rect 28548 8646 28564 8680
rect 28994 8646 29010 8680
rect 29566 8646 29582 8680
rect 30012 8646 30028 8680
rect 30584 8646 30600 8680
rect 31030 8646 31046 8680
rect 31602 8646 31618 8680
rect 32048 8646 32064 8680
rect 32620 8646 32636 8680
rect 33066 8646 33082 8680
rect 33638 8646 33654 8680
rect 10890 8516 10924 8532
rect 13492 8596 13526 8612
rect 2220 8482 2280 8484
rect 3246 8482 3306 8486
rect 4260 8482 4320 8486
rect 5280 8482 5340 8484
rect 6302 8482 6362 8484
rect 8334 8482 8394 8486
rect 9350 8482 9410 8486
rect 10370 8482 10430 8484
rect 1704 8428 1786 8452
rect 1960 8448 1976 8482
rect 2532 8448 2548 8482
rect 1704 8394 1728 8428
rect 1762 8394 1786 8428
rect 1704 8370 1786 8394
rect 2722 8428 2804 8452
rect 2978 8448 2994 8482
rect 3550 8448 3566 8482
rect 2722 8394 2746 8428
rect 2780 8394 2804 8428
rect 1960 8340 1976 8374
rect 2532 8340 2548 8374
rect 2722 8370 2804 8394
rect 3740 8428 3822 8452
rect 3996 8448 4012 8482
rect 4568 8448 4584 8482
rect 3740 8394 3764 8428
rect 3798 8394 3822 8428
rect 2978 8340 2994 8374
rect 3550 8340 3566 8374
rect 3740 8370 3822 8394
rect 4758 8428 4840 8452
rect 5014 8448 5030 8482
rect 5586 8448 5602 8482
rect 4758 8394 4782 8428
rect 4816 8394 4840 8428
rect 3996 8340 4012 8374
rect 4568 8340 4584 8374
rect 4758 8370 4840 8394
rect 5776 8428 5858 8452
rect 6032 8448 6048 8482
rect 6604 8448 6620 8482
rect 5776 8394 5800 8428
rect 5834 8394 5858 8428
rect 5014 8340 5030 8374
rect 5586 8340 5602 8374
rect 5776 8370 5858 8394
rect 6794 8428 6876 8452
rect 7050 8448 7066 8482
rect 7622 8448 7638 8482
rect 6794 8394 6818 8428
rect 6852 8394 6876 8428
rect 6032 8340 6048 8374
rect 6604 8340 6620 8374
rect 6794 8370 6876 8394
rect 7812 8428 7894 8452
rect 8068 8448 8084 8482
rect 8640 8448 8656 8482
rect 7812 8394 7836 8428
rect 7870 8394 7894 8428
rect 7050 8340 7066 8374
rect 7622 8340 7638 8374
rect 7812 8370 7894 8394
rect 8830 8428 8912 8452
rect 9086 8448 9102 8482
rect 9658 8448 9674 8482
rect 8830 8394 8854 8428
rect 8888 8394 8912 8428
rect 8068 8340 8084 8374
rect 8640 8340 8656 8374
rect 8830 8370 8912 8394
rect 9848 8428 9930 8452
rect 10104 8448 10120 8482
rect 10676 8448 10692 8482
rect 9848 8394 9872 8428
rect 9906 8394 9930 8428
rect 9086 8340 9102 8374
rect 9658 8340 9674 8374
rect 9848 8370 9930 8394
rect 10876 8428 10958 8452
rect 10876 8394 10900 8428
rect 10934 8394 10958 8428
rect 10104 8340 10120 8374
rect 10676 8340 10692 8374
rect 10876 8370 10958 8394
rect 1728 8290 1762 8306
rect 1728 7698 1762 7714
rect 2746 8290 2780 8306
rect 2746 7698 2780 7714
rect 3764 8290 3798 8306
rect 3764 7698 3798 7714
rect 4782 8290 4816 8306
rect 4782 7698 4816 7714
rect 5800 8290 5834 8306
rect 5800 7698 5834 7714
rect 6818 8290 6852 8306
rect 6818 7698 6852 7714
rect 7836 8290 7870 8306
rect 7836 7698 7870 7714
rect 8854 8290 8888 8306
rect 8854 7698 8888 7714
rect 9872 8290 9906 8306
rect 9872 7698 9906 7714
rect 10890 8290 10924 8306
rect 13492 8004 13526 8020
rect 14510 8596 14544 8612
rect 14510 8004 14544 8020
rect 15528 8596 15562 8612
rect 15528 8004 15562 8020
rect 16546 8596 16580 8612
rect 16546 8004 16580 8020
rect 17564 8596 17598 8612
rect 17564 8004 17598 8020
rect 18582 8596 18616 8612
rect 18582 8004 18616 8020
rect 19600 8596 19634 8612
rect 19600 8004 19634 8020
rect 20618 8596 20652 8612
rect 20618 8004 20652 8020
rect 21636 8596 21670 8612
rect 21636 8004 21670 8020
rect 22654 8596 22688 8612
rect 22654 8004 22688 8020
rect 23672 8596 23706 8612
rect 23672 8004 23706 8020
rect 24690 8596 24724 8612
rect 24690 8004 24724 8020
rect 25708 8596 25742 8612
rect 25708 8004 25742 8020
rect 26726 8596 26760 8612
rect 26726 8004 26760 8020
rect 27744 8596 27778 8612
rect 27744 8004 27778 8020
rect 28762 8596 28796 8612
rect 28762 8004 28796 8020
rect 29780 8596 29814 8612
rect 29780 8004 29814 8020
rect 30798 8596 30832 8612
rect 30798 8004 30832 8020
rect 31816 8596 31850 8612
rect 31816 8004 31850 8020
rect 32834 8596 32868 8612
rect 32834 8004 32868 8020
rect 33852 8596 33886 8612
rect 33852 8004 33886 8020
rect 13724 7936 13740 7970
rect 14296 7936 14312 7970
rect 14742 7936 14758 7970
rect 15314 7936 15330 7970
rect 15760 7936 15776 7970
rect 16332 7936 16348 7970
rect 16778 7936 16794 7970
rect 17350 7936 17366 7970
rect 17796 7936 17812 7970
rect 18368 7936 18384 7970
rect 18814 7936 18830 7970
rect 19386 7936 19402 7970
rect 19832 7936 19848 7970
rect 20404 7936 20420 7970
rect 20850 7936 20866 7970
rect 21422 7936 21438 7970
rect 21868 7936 21884 7970
rect 22440 7936 22456 7970
rect 22886 7936 22902 7970
rect 23458 7936 23474 7970
rect 23904 7936 23920 7970
rect 24476 7936 24492 7970
rect 24922 7936 24938 7970
rect 25494 7936 25510 7970
rect 25940 7936 25956 7970
rect 26512 7936 26528 7970
rect 26958 7936 26974 7970
rect 27530 7936 27546 7970
rect 27976 7936 27992 7970
rect 28548 7936 28564 7970
rect 28994 7936 29010 7970
rect 29566 7936 29582 7970
rect 30012 7936 30028 7970
rect 30584 7936 30600 7970
rect 31030 7936 31046 7970
rect 31602 7936 31618 7970
rect 32048 7936 32064 7970
rect 32620 7936 32636 7970
rect 33066 7936 33082 7970
rect 33638 7936 33654 7970
rect 10890 7698 10924 7714
rect 13998 7728 14080 7752
rect 13998 7694 14022 7728
rect 14056 7694 14080 7728
rect 13998 7670 14080 7694
rect 15016 7728 15098 7752
rect 15016 7694 15040 7728
rect 15074 7694 15098 7728
rect 15016 7670 15098 7694
rect 16034 7728 16116 7752
rect 16034 7694 16058 7728
rect 16092 7694 16116 7728
rect 16034 7670 16116 7694
rect 17052 7728 17134 7752
rect 17052 7694 17076 7728
rect 17110 7694 17134 7728
rect 17052 7670 17134 7694
rect 18070 7728 18152 7752
rect 18070 7694 18094 7728
rect 18128 7694 18152 7728
rect 18070 7670 18152 7694
rect 19088 7728 19170 7752
rect 19088 7694 19112 7728
rect 19146 7694 19170 7728
rect 19088 7670 19170 7694
rect 20106 7728 20188 7752
rect 20106 7694 20130 7728
rect 20164 7694 20188 7728
rect 20106 7670 20188 7694
rect 21124 7728 21206 7752
rect 21124 7694 21148 7728
rect 21182 7694 21206 7728
rect 21124 7670 21206 7694
rect 22142 7728 22224 7752
rect 22142 7694 22166 7728
rect 22200 7694 22224 7728
rect 22142 7670 22224 7694
rect 23160 7728 23242 7752
rect 23160 7694 23184 7728
rect 23218 7694 23242 7728
rect 23160 7670 23242 7694
rect 24178 7728 24260 7752
rect 24178 7694 24202 7728
rect 24236 7694 24260 7728
rect 24178 7670 24260 7694
rect 25196 7728 25278 7752
rect 25196 7694 25220 7728
rect 25254 7694 25278 7728
rect 25196 7670 25278 7694
rect 26214 7728 26296 7752
rect 26214 7694 26238 7728
rect 26272 7694 26296 7728
rect 26214 7670 26296 7694
rect 27232 7728 27314 7752
rect 27232 7694 27256 7728
rect 27290 7694 27314 7728
rect 27232 7670 27314 7694
rect 28250 7728 28332 7752
rect 28250 7694 28274 7728
rect 28308 7694 28332 7728
rect 28250 7670 28332 7694
rect 29268 7728 29350 7752
rect 29268 7694 29292 7728
rect 29326 7694 29350 7728
rect 29268 7670 29350 7694
rect 30286 7728 30368 7752
rect 30286 7694 30310 7728
rect 30344 7694 30368 7728
rect 30286 7670 30368 7694
rect 31304 7728 31386 7752
rect 31304 7694 31328 7728
rect 31362 7694 31386 7728
rect 31304 7670 31386 7694
rect 32322 7728 32404 7752
rect 32322 7694 32346 7728
rect 32380 7694 32404 7728
rect 32322 7670 32404 7694
rect 33340 7728 33422 7752
rect 33340 7694 33364 7728
rect 33398 7694 33422 7728
rect 33340 7670 33422 7694
rect 1960 7630 1976 7664
rect 2532 7630 2548 7664
rect 2978 7630 2994 7664
rect 3550 7630 3566 7664
rect 3996 7630 4012 7664
rect 4568 7630 4584 7664
rect 5014 7630 5030 7664
rect 5586 7630 5602 7664
rect 6032 7630 6048 7664
rect 6604 7630 6620 7664
rect 7050 7630 7066 7664
rect 7622 7630 7638 7664
rect 8068 7630 8084 7664
rect 8640 7630 8656 7664
rect 9086 7630 9102 7664
rect 9658 7630 9674 7664
rect 10104 7630 10120 7664
rect 10676 7630 10692 7664
rect 1692 7534 1774 7558
rect 1692 7500 1716 7534
rect 1750 7500 1774 7534
rect 1692 7476 1774 7500
rect 2710 7534 2792 7558
rect 2710 7500 2734 7534
rect 2768 7500 2792 7534
rect 2710 7476 2792 7500
rect 3728 7534 3810 7558
rect 3728 7500 3752 7534
rect 3786 7500 3810 7534
rect 3728 7476 3810 7500
rect 4746 7534 4828 7558
rect 4746 7500 4770 7534
rect 4804 7500 4828 7534
rect 4746 7476 4828 7500
rect 5764 7534 5846 7558
rect 5764 7500 5788 7534
rect 5822 7500 5846 7534
rect 5764 7476 5846 7500
rect 6782 7534 6864 7558
rect 6782 7500 6806 7534
rect 6840 7500 6864 7534
rect 6782 7476 6864 7500
rect 7800 7534 7882 7558
rect 7800 7500 7824 7534
rect 7858 7500 7882 7534
rect 7800 7476 7882 7500
rect 8818 7534 8900 7558
rect 8818 7500 8842 7534
rect 8876 7500 8900 7534
rect 8818 7476 8900 7500
rect 9836 7534 9918 7558
rect 9836 7500 9860 7534
rect 9894 7500 9918 7534
rect 9836 7476 9918 7500
rect 10864 7534 10946 7558
rect 10864 7500 10888 7534
rect 10922 7500 10946 7534
rect 10864 7476 10946 7500
rect 13724 7414 13740 7448
rect 14296 7414 14312 7448
rect 14742 7414 14758 7448
rect 15314 7414 15330 7448
rect 15760 7414 15776 7448
rect 16332 7414 16348 7448
rect 16778 7414 16794 7448
rect 17350 7414 17366 7448
rect 17796 7414 17812 7448
rect 18368 7414 18384 7448
rect 18814 7414 18830 7448
rect 19386 7414 19402 7448
rect 19832 7414 19848 7448
rect 20404 7414 20420 7448
rect 20850 7414 20866 7448
rect 21422 7414 21438 7448
rect 21868 7414 21884 7448
rect 22440 7414 22456 7448
rect 22886 7414 22902 7448
rect 23458 7414 23474 7448
rect 23904 7414 23920 7448
rect 24476 7414 24492 7448
rect 24922 7414 24938 7448
rect 25494 7414 25510 7448
rect 25940 7414 25956 7448
rect 26512 7414 26528 7448
rect 26958 7414 26974 7448
rect 27530 7414 27546 7448
rect 27976 7414 27992 7448
rect 28548 7414 28564 7448
rect 28994 7414 29010 7448
rect 29566 7414 29582 7448
rect 30012 7414 30028 7448
rect 30584 7414 30600 7448
rect 31030 7414 31046 7448
rect 31602 7414 31618 7448
rect 32048 7414 32064 7448
rect 32620 7414 32636 7448
rect 33066 7414 33082 7448
rect 33638 7414 33654 7448
rect 13492 7364 13526 7380
rect 13492 6772 13526 6788
rect 14510 7364 14544 7380
rect 14510 6772 14544 6788
rect 15528 7364 15562 7380
rect 15528 6772 15562 6788
rect 16546 7364 16580 7380
rect 16546 6772 16580 6788
rect 17564 7364 17598 7380
rect 17564 6772 17598 6788
rect 18582 7364 18616 7380
rect 18582 6772 18616 6788
rect 19600 7364 19634 7380
rect 19600 6772 19634 6788
rect 20618 7364 20652 7380
rect 20618 6772 20652 6788
rect 21636 7364 21670 7380
rect 21636 6772 21670 6788
rect 22654 7364 22688 7380
rect 22654 6772 22688 6788
rect 23672 7364 23706 7380
rect 23672 6772 23706 6788
rect 24690 7364 24724 7380
rect 24690 6772 24724 6788
rect 25708 7364 25742 7380
rect 25708 6772 25742 6788
rect 26726 7364 26760 7380
rect 26726 6772 26760 6788
rect 27744 7364 27778 7380
rect 27744 6772 27778 6788
rect 28762 7364 28796 7380
rect 28762 6772 28796 6788
rect 29780 7364 29814 7380
rect 29780 6772 29814 6788
rect 30798 7364 30832 7380
rect 30798 6772 30832 6788
rect 31816 7364 31850 7380
rect 31816 6772 31850 6788
rect 32834 7364 32868 7380
rect 32834 6772 32868 6788
rect 33852 7364 33886 7380
rect 33852 6772 33886 6788
rect 22142 6738 22202 6740
rect 24186 6738 24246 6742
rect 32320 6738 32380 6740
rect 13724 6704 13740 6738
rect 14296 6704 14312 6738
rect 14742 6704 14758 6738
rect 15314 6704 15330 6738
rect 15760 6704 15776 6738
rect 16332 6704 16348 6738
rect 16778 6704 16794 6738
rect 17350 6704 17366 6738
rect 17796 6704 17812 6738
rect 18368 6704 18384 6738
rect 18814 6704 18830 6738
rect 19386 6704 19402 6738
rect 19832 6704 19848 6738
rect 20404 6704 20420 6738
rect 20850 6704 20866 6738
rect 21422 6704 21438 6738
rect 21868 6704 21884 6738
rect 22440 6704 22456 6738
rect 22886 6704 22902 6738
rect 23458 6704 23474 6738
rect 23904 6704 23920 6738
rect 24476 6704 24492 6738
rect 24922 6704 24938 6738
rect 25494 6704 25510 6738
rect 25940 6704 25956 6738
rect 26512 6704 26528 6738
rect 26958 6704 26974 6738
rect 27530 6704 27546 6738
rect 27976 6704 27992 6738
rect 28548 6704 28564 6738
rect 28994 6704 29010 6738
rect 29566 6704 29582 6738
rect 30012 6704 30028 6738
rect 30584 6704 30600 6738
rect 31030 6704 31046 6738
rect 31602 6704 31618 6738
rect 32048 6704 32064 6738
rect 32620 6704 32636 6738
rect 33066 6704 33082 6738
rect 33638 6704 33654 6738
rect 896 6586 978 6610
rect 896 6552 920 6586
rect 954 6552 978 6586
rect 896 6528 978 6552
rect 1914 6586 1996 6610
rect 1914 6552 1938 6586
rect 1972 6552 1996 6586
rect 1914 6528 1996 6552
rect 2932 6586 3014 6610
rect 2932 6552 2956 6586
rect 2990 6552 3014 6586
rect 2932 6528 3014 6552
rect 3950 6586 4032 6610
rect 3950 6552 3974 6586
rect 4008 6552 4032 6586
rect 3950 6528 4032 6552
rect 4968 6586 5050 6610
rect 4968 6552 4992 6586
rect 5026 6552 5050 6586
rect 4968 6528 5050 6552
rect 5986 6586 6068 6610
rect 5986 6552 6010 6586
rect 6044 6552 6068 6586
rect 5986 6528 6068 6552
rect 7004 6586 7086 6610
rect 7004 6552 7028 6586
rect 7062 6552 7086 6586
rect 7004 6528 7086 6552
rect 8022 6586 8104 6610
rect 8022 6552 8046 6586
rect 8080 6552 8104 6586
rect 8022 6528 8104 6552
rect 9040 6586 9122 6610
rect 9040 6552 9064 6586
rect 9098 6552 9122 6586
rect 9040 6528 9122 6552
rect 10058 6586 10140 6610
rect 10058 6552 10082 6586
rect 10116 6552 10140 6586
rect 10058 6528 10140 6552
rect 11076 6586 11158 6610
rect 11076 6552 11100 6586
rect 11134 6552 11158 6586
rect 11076 6528 11158 6552
rect 13998 6480 14080 6504
rect 13998 6446 14022 6480
rect 14056 6446 14080 6480
rect 13998 6422 14080 6446
rect 15016 6480 15098 6504
rect 15016 6446 15040 6480
rect 15074 6446 15098 6480
rect 15016 6422 15098 6446
rect 16034 6480 16116 6504
rect 16034 6446 16058 6480
rect 16092 6446 16116 6480
rect 16034 6422 16116 6446
rect 17052 6480 17134 6504
rect 17052 6446 17076 6480
rect 17110 6446 17134 6480
rect 17052 6422 17134 6446
rect 18070 6480 18152 6504
rect 18070 6446 18094 6480
rect 18128 6446 18152 6480
rect 18070 6422 18152 6446
rect 19088 6480 19170 6504
rect 19088 6446 19112 6480
rect 19146 6446 19170 6480
rect 19088 6422 19170 6446
rect 20106 6480 20188 6504
rect 20106 6446 20130 6480
rect 20164 6446 20188 6480
rect 20106 6422 20188 6446
rect 21124 6480 21206 6504
rect 21124 6446 21148 6480
rect 21182 6446 21206 6480
rect 21124 6422 21206 6446
rect 22142 6480 22224 6504
rect 22142 6446 22166 6480
rect 22200 6446 22224 6480
rect 22142 6422 22224 6446
rect 23160 6480 23242 6504
rect 23160 6446 23184 6480
rect 23218 6446 23242 6480
rect 23160 6422 23242 6446
rect 24178 6480 24260 6504
rect 24178 6446 24202 6480
rect 24236 6446 24260 6480
rect 24178 6422 24260 6446
rect 25196 6480 25278 6504
rect 25196 6446 25220 6480
rect 25254 6446 25278 6480
rect 25196 6422 25278 6446
rect 26214 6480 26296 6504
rect 26214 6446 26238 6480
rect 26272 6446 26296 6480
rect 26214 6422 26296 6446
rect 27232 6480 27314 6504
rect 27232 6446 27256 6480
rect 27290 6446 27314 6480
rect 27232 6422 27314 6446
rect 28250 6480 28332 6504
rect 28250 6446 28274 6480
rect 28308 6446 28332 6480
rect 28250 6422 28332 6446
rect 29268 6480 29350 6504
rect 29268 6446 29292 6480
rect 29326 6446 29350 6480
rect 29268 6422 29350 6446
rect 30286 6480 30368 6504
rect 30286 6446 30310 6480
rect 30344 6446 30368 6480
rect 30286 6422 30368 6446
rect 31304 6480 31386 6504
rect 31304 6446 31328 6480
rect 31362 6446 31386 6480
rect 31304 6422 31386 6446
rect 32322 6480 32404 6504
rect 32322 6446 32346 6480
rect 32380 6446 32404 6480
rect 32322 6422 32404 6446
rect 33340 6480 33422 6504
rect 33340 6446 33364 6480
rect 33398 6446 33422 6480
rect 33340 6422 33422 6446
rect 636 6316 652 6350
rect 1208 6316 1224 6350
rect 1654 6316 1670 6350
rect 2226 6316 2242 6350
rect 2672 6316 2688 6350
rect 3244 6316 3260 6350
rect 3690 6316 3706 6350
rect 4262 6316 4278 6350
rect 4708 6316 4724 6350
rect 5280 6316 5296 6350
rect 5726 6316 5742 6350
rect 6298 6316 6314 6350
rect 6744 6316 6760 6350
rect 7316 6316 7332 6350
rect 7762 6316 7778 6350
rect 8334 6316 8350 6350
rect 8780 6316 8796 6350
rect 9352 6316 9368 6350
rect 9798 6316 9814 6350
rect 10370 6316 10386 6350
rect 10816 6316 10832 6350
rect 11388 6316 11404 6350
rect 404 6266 438 6282
rect 404 5674 438 5690
rect 1422 6266 1456 6282
rect 1422 5674 1456 5690
rect 2440 6266 2474 6282
rect 2440 5674 2474 5690
rect 3458 6266 3492 6282
rect 3458 5674 3492 5690
rect 4476 6266 4510 6282
rect 4476 5674 4510 5690
rect 5494 6266 5528 6282
rect 5494 5674 5528 5690
rect 6512 6266 6546 6282
rect 6512 5674 6546 5690
rect 7530 6266 7564 6282
rect 7530 5674 7564 5690
rect 8548 6266 8582 6282
rect 8548 5674 8582 5690
rect 9566 6266 9600 6282
rect 9566 5674 9600 5690
rect 10584 6266 10618 6282
rect 10584 5674 10618 5690
rect 11602 6266 11636 6282
rect 13724 6180 13740 6214
rect 14296 6180 14312 6214
rect 14742 6180 14758 6214
rect 15314 6180 15330 6214
rect 15760 6180 15776 6214
rect 16332 6180 16348 6214
rect 16778 6180 16794 6214
rect 17350 6180 17366 6214
rect 17796 6180 17812 6214
rect 18368 6180 18384 6214
rect 18814 6180 18830 6214
rect 19386 6180 19402 6214
rect 19832 6180 19848 6214
rect 20404 6180 20420 6214
rect 20850 6180 20866 6214
rect 21422 6180 21438 6214
rect 21868 6180 21884 6214
rect 22440 6180 22456 6214
rect 22886 6180 22902 6214
rect 23458 6180 23474 6214
rect 23904 6180 23920 6214
rect 24476 6180 24492 6214
rect 24922 6180 24938 6214
rect 25494 6180 25510 6214
rect 25940 6180 25956 6214
rect 26512 6180 26528 6214
rect 26958 6180 26974 6214
rect 27530 6180 27546 6214
rect 27976 6180 27992 6214
rect 28548 6180 28564 6214
rect 28994 6180 29010 6214
rect 29566 6180 29582 6214
rect 30012 6180 30028 6214
rect 30584 6180 30600 6214
rect 31030 6180 31046 6214
rect 31602 6180 31618 6214
rect 32048 6180 32064 6214
rect 32620 6180 32636 6214
rect 33066 6180 33082 6214
rect 33638 6180 33654 6214
rect 11602 5674 11636 5690
rect 13492 6130 13526 6146
rect 636 5606 652 5640
rect 1208 5606 1224 5640
rect 1654 5606 1670 5640
rect 2226 5606 2242 5640
rect 2672 5606 2688 5640
rect 3244 5606 3260 5640
rect 3690 5606 3706 5640
rect 4262 5606 4278 5640
rect 4708 5606 4724 5640
rect 5280 5606 5296 5640
rect 5726 5606 5742 5640
rect 6298 5606 6314 5640
rect 6744 5606 6760 5640
rect 7316 5606 7332 5640
rect 7762 5606 7778 5640
rect 8334 5606 8350 5640
rect 8780 5606 8796 5640
rect 9352 5606 9368 5640
rect 9798 5606 9814 5640
rect 10370 5606 10386 5640
rect 10816 5606 10832 5640
rect 11388 5606 11404 5640
rect 13492 5538 13526 5554
rect 14510 6130 14544 6146
rect 14510 5538 14544 5554
rect 15528 6130 15562 6146
rect 15528 5538 15562 5554
rect 16546 6130 16580 6146
rect 16546 5538 16580 5554
rect 17564 6130 17598 6146
rect 17564 5538 17598 5554
rect 18582 6130 18616 6146
rect 18582 5538 18616 5554
rect 19600 6130 19634 6146
rect 19600 5538 19634 5554
rect 20618 6130 20652 6146
rect 20618 5538 20652 5554
rect 21636 6130 21670 6146
rect 21636 5538 21670 5554
rect 22654 6130 22688 6146
rect 22654 5538 22688 5554
rect 23672 6130 23706 6146
rect 23672 5538 23706 5554
rect 24690 6130 24724 6146
rect 24690 5538 24724 5554
rect 25708 6130 25742 6146
rect 25708 5538 25742 5554
rect 26726 6130 26760 6146
rect 26726 5538 26760 5554
rect 27744 6130 27778 6146
rect 27744 5538 27778 5554
rect 28762 6130 28796 6146
rect 28762 5538 28796 5554
rect 29780 6130 29814 6146
rect 29780 5538 29814 5554
rect 30798 6130 30832 6146
rect 30798 5538 30832 5554
rect 31816 6130 31850 6146
rect 31816 5538 31850 5554
rect 32834 6130 32868 6146
rect 32834 5538 32868 5554
rect 33852 6130 33886 6146
rect 33852 5538 33886 5554
rect 16018 5504 16078 5508
rect 13724 5470 13740 5504
rect 14296 5470 14312 5504
rect 14742 5470 14758 5504
rect 15314 5470 15330 5504
rect 15760 5470 15776 5504
rect 16332 5470 16348 5504
rect 16778 5470 16794 5504
rect 17350 5470 17366 5504
rect 17796 5470 17812 5504
rect 18368 5470 18384 5504
rect 18814 5470 18830 5504
rect 19386 5470 19402 5504
rect 19832 5470 19848 5504
rect 20404 5470 20420 5504
rect 20850 5470 20866 5504
rect 21422 5470 21438 5504
rect 21868 5470 21884 5504
rect 22440 5470 22456 5504
rect 22886 5470 22902 5504
rect 23458 5470 23474 5504
rect 23904 5470 23920 5504
rect 24476 5470 24492 5504
rect 24922 5470 24938 5504
rect 25494 5470 25510 5504
rect 25940 5470 25956 5504
rect 26512 5470 26528 5504
rect 26958 5470 26974 5504
rect 27530 5470 27546 5504
rect 27976 5470 27992 5504
rect 28548 5470 28564 5504
rect 28994 5470 29010 5504
rect 29566 5470 29582 5504
rect 30012 5470 30028 5504
rect 30584 5470 30600 5504
rect 31030 5470 31046 5504
rect 31602 5470 31618 5504
rect 32048 5470 32064 5504
rect 32620 5470 32636 5504
rect 33066 5470 33082 5504
rect 33638 5470 33654 5504
rect 908 5444 990 5468
rect 908 5410 932 5444
rect 966 5410 990 5444
rect 908 5386 990 5410
rect 1926 5444 2008 5468
rect 1926 5410 1950 5444
rect 1984 5410 2008 5444
rect 1926 5386 2008 5410
rect 2944 5444 3026 5468
rect 2944 5410 2968 5444
rect 3002 5410 3026 5444
rect 2944 5386 3026 5410
rect 3962 5444 4044 5468
rect 3962 5410 3986 5444
rect 4020 5410 4044 5444
rect 3962 5386 4044 5410
rect 4980 5444 5062 5468
rect 4980 5410 5004 5444
rect 5038 5410 5062 5444
rect 4980 5386 5062 5410
rect 5998 5444 6080 5468
rect 5998 5410 6022 5444
rect 6056 5410 6080 5444
rect 5998 5386 6080 5410
rect 7016 5444 7098 5468
rect 7016 5410 7040 5444
rect 7074 5410 7098 5444
rect 7016 5386 7098 5410
rect 8034 5444 8116 5468
rect 8034 5410 8058 5444
rect 8092 5410 8116 5444
rect 8034 5386 8116 5410
rect 9052 5444 9134 5468
rect 9052 5410 9076 5444
rect 9110 5410 9134 5444
rect 9052 5386 9134 5410
rect 10070 5444 10152 5468
rect 10070 5410 10094 5444
rect 10128 5410 10152 5444
rect 10070 5386 10152 5410
rect 11088 5444 11170 5468
rect 11088 5410 11112 5444
rect 11146 5410 11170 5444
rect 11088 5386 11170 5410
rect 13974 5244 14056 5268
rect 636 5204 652 5238
rect 1208 5204 1224 5238
rect 1654 5204 1670 5238
rect 2226 5204 2242 5238
rect 2672 5204 2688 5238
rect 3244 5204 3260 5238
rect 3690 5204 3706 5238
rect 4262 5204 4278 5238
rect 4708 5204 4724 5238
rect 5280 5204 5296 5238
rect 5726 5204 5742 5238
rect 6298 5204 6314 5238
rect 6744 5204 6760 5238
rect 7316 5204 7332 5238
rect 7762 5204 7778 5238
rect 8334 5204 8350 5238
rect 8780 5204 8796 5238
rect 9352 5204 9368 5238
rect 9798 5204 9814 5238
rect 10370 5204 10386 5238
rect 10816 5204 10832 5238
rect 11388 5204 11404 5238
rect 13974 5210 13998 5244
rect 14032 5210 14056 5244
rect 13974 5186 14056 5210
rect 14992 5244 15074 5268
rect 14992 5210 15016 5244
rect 15050 5210 15074 5244
rect 14992 5186 15074 5210
rect 16010 5244 16092 5268
rect 16010 5210 16034 5244
rect 16068 5210 16092 5244
rect 16010 5186 16092 5210
rect 17028 5244 17110 5268
rect 17028 5210 17052 5244
rect 17086 5210 17110 5244
rect 17028 5186 17110 5210
rect 18046 5244 18128 5268
rect 18046 5210 18070 5244
rect 18104 5210 18128 5244
rect 18046 5186 18128 5210
rect 19064 5244 19146 5268
rect 19064 5210 19088 5244
rect 19122 5210 19146 5244
rect 19064 5186 19146 5210
rect 20082 5244 20164 5268
rect 20082 5210 20106 5244
rect 20140 5210 20164 5244
rect 20082 5186 20164 5210
rect 21100 5244 21182 5268
rect 21100 5210 21124 5244
rect 21158 5210 21182 5244
rect 21100 5186 21182 5210
rect 22118 5244 22200 5268
rect 22118 5210 22142 5244
rect 22176 5210 22200 5244
rect 22118 5186 22200 5210
rect 23136 5244 23218 5268
rect 23136 5210 23160 5244
rect 23194 5210 23218 5244
rect 23136 5186 23218 5210
rect 24154 5244 24236 5268
rect 24154 5210 24178 5244
rect 24212 5210 24236 5244
rect 24154 5186 24236 5210
rect 25172 5244 25254 5268
rect 25172 5210 25196 5244
rect 25230 5210 25254 5244
rect 25172 5186 25254 5210
rect 26190 5244 26272 5268
rect 26190 5210 26214 5244
rect 26248 5210 26272 5244
rect 26190 5186 26272 5210
rect 27208 5244 27290 5268
rect 27208 5210 27232 5244
rect 27266 5210 27290 5244
rect 27208 5186 27290 5210
rect 28226 5244 28308 5268
rect 28226 5210 28250 5244
rect 28284 5210 28308 5244
rect 28226 5186 28308 5210
rect 29244 5244 29326 5268
rect 29244 5210 29268 5244
rect 29302 5210 29326 5244
rect 29244 5186 29326 5210
rect 30262 5244 30344 5268
rect 30262 5210 30286 5244
rect 30320 5210 30344 5244
rect 30262 5186 30344 5210
rect 31280 5244 31362 5268
rect 31280 5210 31304 5244
rect 31338 5210 31362 5244
rect 31280 5186 31362 5210
rect 32298 5244 32380 5268
rect 32298 5210 32322 5244
rect 32356 5210 32380 5244
rect 32298 5186 32380 5210
rect 33316 5244 33398 5268
rect 33316 5210 33340 5244
rect 33374 5210 33398 5244
rect 33316 5186 33398 5210
rect 404 5154 438 5170
rect 404 4562 438 4578
rect 1422 5154 1456 5170
rect 1422 4562 1456 4578
rect 2440 5154 2474 5170
rect 2440 4562 2474 4578
rect 3458 5154 3492 5170
rect 3458 4562 3492 4578
rect 4476 5154 4510 5170
rect 4476 4562 4510 4578
rect 5494 5154 5528 5170
rect 5494 4562 5528 4578
rect 6512 5154 6546 5170
rect 6512 4562 6546 4578
rect 7530 5154 7564 5170
rect 7530 4562 7564 4578
rect 8548 5154 8582 5170
rect 8548 4562 8582 4578
rect 9566 5154 9600 5170
rect 9566 4562 9600 4578
rect 10584 5154 10618 5170
rect 10584 4562 10618 4578
rect 11602 5154 11636 5170
rect 13724 4946 13740 4980
rect 14296 4946 14312 4980
rect 14742 4946 14758 4980
rect 15314 4946 15330 4980
rect 15760 4946 15776 4980
rect 16332 4946 16348 4980
rect 16778 4946 16794 4980
rect 17350 4946 17366 4980
rect 17796 4946 17812 4980
rect 18368 4946 18384 4980
rect 18814 4946 18830 4980
rect 19386 4946 19402 4980
rect 19832 4946 19848 4980
rect 20404 4946 20420 4980
rect 20850 4946 20866 4980
rect 21422 4946 21438 4980
rect 21868 4946 21884 4980
rect 22440 4946 22456 4980
rect 22886 4946 22902 4980
rect 23458 4946 23474 4980
rect 23904 4946 23920 4980
rect 24476 4946 24492 4980
rect 24922 4946 24938 4980
rect 25494 4946 25510 4980
rect 25940 4946 25956 4980
rect 26512 4946 26528 4980
rect 26958 4946 26974 4980
rect 27530 4946 27546 4980
rect 27976 4946 27992 4980
rect 28548 4946 28564 4980
rect 28994 4946 29010 4980
rect 29566 4946 29582 4980
rect 30012 4946 30028 4980
rect 30584 4946 30600 4980
rect 31030 4946 31046 4980
rect 31602 4946 31618 4980
rect 32048 4946 32064 4980
rect 32620 4946 32636 4980
rect 33066 4946 33082 4980
rect 33638 4946 33654 4980
rect 11602 4562 11636 4578
rect 13492 4896 13526 4912
rect 636 4494 652 4528
rect 1208 4494 1224 4528
rect 1654 4494 1670 4528
rect 2226 4494 2242 4528
rect 2672 4494 2688 4528
rect 3244 4494 3260 4528
rect 3690 4494 3706 4528
rect 4262 4494 4278 4528
rect 4708 4494 4724 4528
rect 5280 4494 5296 4528
rect 5726 4494 5742 4528
rect 6298 4494 6314 4528
rect 6744 4494 6760 4528
rect 7316 4494 7332 4528
rect 7762 4494 7778 4528
rect 8334 4494 8350 4528
rect 8780 4494 8796 4528
rect 9352 4494 9368 4528
rect 9798 4494 9814 4528
rect 10370 4494 10386 4528
rect 10816 4494 10832 4528
rect 11388 4494 11404 4528
rect 886 4336 968 4360
rect 886 4302 910 4336
rect 944 4302 968 4336
rect 886 4278 968 4302
rect 1904 4336 1986 4360
rect 1904 4302 1928 4336
rect 1962 4302 1986 4336
rect 1904 4278 1986 4302
rect 2922 4336 3004 4360
rect 2922 4302 2946 4336
rect 2980 4302 3004 4336
rect 2922 4278 3004 4302
rect 3940 4336 4022 4360
rect 3940 4302 3964 4336
rect 3998 4302 4022 4336
rect 3940 4278 4022 4302
rect 4958 4336 5040 4360
rect 4958 4302 4982 4336
rect 5016 4302 5040 4336
rect 4958 4278 5040 4302
rect 5976 4336 6058 4360
rect 5976 4302 6000 4336
rect 6034 4302 6058 4336
rect 5976 4278 6058 4302
rect 6994 4336 7076 4360
rect 6994 4302 7018 4336
rect 7052 4302 7076 4336
rect 6994 4278 7076 4302
rect 8012 4336 8094 4360
rect 8012 4302 8036 4336
rect 8070 4302 8094 4336
rect 8012 4278 8094 4302
rect 9030 4336 9112 4360
rect 9030 4302 9054 4336
rect 9088 4302 9112 4336
rect 9030 4278 9112 4302
rect 10048 4336 10130 4360
rect 10048 4302 10072 4336
rect 10106 4302 10130 4336
rect 10048 4278 10130 4302
rect 11066 4336 11148 4360
rect 11066 4302 11090 4336
rect 11124 4302 11148 4336
rect 13492 4304 13526 4320
rect 14510 4896 14544 4912
rect 14510 4304 14544 4320
rect 15528 4896 15562 4912
rect 15528 4304 15562 4320
rect 16546 4896 16580 4912
rect 16546 4304 16580 4320
rect 17564 4896 17598 4912
rect 17564 4304 17598 4320
rect 18582 4896 18616 4912
rect 18582 4304 18616 4320
rect 19600 4896 19634 4912
rect 19600 4304 19634 4320
rect 20618 4896 20652 4912
rect 20618 4304 20652 4320
rect 21636 4896 21670 4912
rect 21636 4304 21670 4320
rect 22654 4896 22688 4912
rect 22654 4304 22688 4320
rect 23672 4896 23706 4912
rect 23672 4304 23706 4320
rect 24690 4896 24724 4912
rect 24690 4304 24724 4320
rect 25708 4896 25742 4912
rect 25708 4304 25742 4320
rect 26726 4896 26760 4912
rect 26726 4304 26760 4320
rect 27744 4896 27778 4912
rect 27744 4304 27778 4320
rect 28762 4896 28796 4912
rect 28762 4304 28796 4320
rect 29780 4896 29814 4912
rect 29780 4304 29814 4320
rect 30798 4896 30832 4912
rect 30798 4304 30832 4320
rect 31816 4896 31850 4912
rect 31816 4304 31850 4320
rect 32834 4896 32868 4912
rect 32834 4304 32868 4320
rect 33852 4896 33886 4912
rect 33852 4304 33886 4320
rect 11066 4278 11148 4302
rect 22142 4270 22202 4272
rect 24186 4270 24246 4274
rect 27224 4270 27284 4274
rect 13724 4236 13740 4270
rect 14296 4236 14312 4270
rect 14742 4236 14758 4270
rect 15314 4236 15330 4270
rect 15760 4236 15776 4270
rect 16332 4236 16348 4270
rect 16778 4236 16794 4270
rect 17350 4236 17366 4270
rect 17796 4236 17812 4270
rect 18368 4236 18384 4270
rect 18814 4236 18830 4270
rect 19386 4236 19402 4270
rect 19832 4236 19848 4270
rect 20404 4236 20420 4270
rect 20850 4236 20866 4270
rect 21422 4236 21438 4270
rect 21868 4236 21884 4270
rect 22440 4236 22456 4270
rect 22886 4236 22902 4270
rect 23458 4236 23474 4270
rect 23904 4236 23920 4270
rect 24476 4236 24492 4270
rect 24922 4236 24938 4270
rect 25494 4236 25510 4270
rect 25940 4236 25956 4270
rect 26512 4236 26528 4270
rect 26958 4236 26974 4270
rect 27530 4236 27546 4270
rect 27976 4236 27992 4270
rect 28548 4236 28564 4270
rect 28994 4236 29010 4270
rect 29566 4236 29582 4270
rect 30012 4236 30028 4270
rect 30584 4236 30600 4270
rect 31030 4236 31046 4270
rect 31602 4236 31618 4270
rect 32048 4236 32064 4270
rect 32620 4236 32636 4270
rect 33066 4236 33082 4270
rect 33638 4236 33654 4270
rect 636 4092 652 4126
rect 1208 4092 1224 4126
rect 1654 4092 1670 4126
rect 2226 4092 2242 4126
rect 2672 4092 2688 4126
rect 3244 4092 3260 4126
rect 3690 4092 3706 4126
rect 4262 4092 4278 4126
rect 4708 4092 4724 4126
rect 5280 4092 5296 4126
rect 5726 4092 5742 4126
rect 6298 4092 6314 4126
rect 6744 4092 6760 4126
rect 7316 4092 7332 4126
rect 7762 4092 7778 4126
rect 8334 4092 8350 4126
rect 8780 4092 8796 4126
rect 9352 4092 9368 4126
rect 9798 4092 9814 4126
rect 10370 4092 10386 4126
rect 10816 4092 10832 4126
rect 11388 4092 11404 4126
rect 404 4042 438 4058
rect 404 3450 438 3466
rect 1422 4042 1456 4058
rect 1422 3450 1456 3466
rect 2440 4042 2474 4058
rect 2440 3450 2474 3466
rect 3458 4042 3492 4058
rect 3458 3450 3492 3466
rect 4476 4042 4510 4058
rect 4476 3450 4510 3466
rect 5494 4042 5528 4058
rect 5494 3450 5528 3466
rect 6512 4042 6546 4058
rect 6512 3450 6546 3466
rect 7530 4042 7564 4058
rect 7530 3450 7564 3466
rect 8548 4042 8582 4058
rect 8548 3450 8582 3466
rect 9566 4042 9600 4058
rect 9566 3450 9600 3466
rect 10584 4042 10618 4058
rect 10584 3450 10618 3466
rect 11602 4042 11636 4058
rect 13986 4020 14068 4044
rect 13986 3986 14010 4020
rect 14044 3986 14068 4020
rect 13986 3962 14068 3986
rect 15004 4020 15086 4044
rect 15004 3986 15028 4020
rect 15062 3986 15086 4020
rect 15004 3962 15086 3986
rect 16022 4020 16104 4044
rect 16022 3986 16046 4020
rect 16080 3986 16104 4020
rect 16022 3962 16104 3986
rect 17040 4020 17122 4044
rect 17040 3986 17064 4020
rect 17098 3986 17122 4020
rect 17040 3962 17122 3986
rect 18058 4020 18140 4044
rect 18058 3986 18082 4020
rect 18116 3986 18140 4020
rect 18058 3962 18140 3986
rect 19076 4020 19158 4044
rect 19076 3986 19100 4020
rect 19134 3986 19158 4020
rect 19076 3962 19158 3986
rect 20094 4020 20176 4044
rect 20094 3986 20118 4020
rect 20152 3986 20176 4020
rect 20094 3962 20176 3986
rect 21112 4020 21194 4044
rect 21112 3986 21136 4020
rect 21170 3986 21194 4020
rect 21112 3962 21194 3986
rect 22130 4020 22212 4044
rect 22130 3986 22154 4020
rect 22188 3986 22212 4020
rect 22130 3962 22212 3986
rect 23148 4020 23230 4044
rect 23148 3986 23172 4020
rect 23206 3986 23230 4020
rect 23148 3962 23230 3986
rect 24166 4020 24248 4044
rect 24166 3986 24190 4020
rect 24224 3986 24248 4020
rect 24166 3962 24248 3986
rect 25184 4020 25266 4044
rect 25184 3986 25208 4020
rect 25242 3986 25266 4020
rect 25184 3962 25266 3986
rect 26202 4020 26284 4044
rect 26202 3986 26226 4020
rect 26260 3986 26284 4020
rect 26202 3962 26284 3986
rect 27220 4020 27302 4044
rect 27220 3986 27244 4020
rect 27278 3986 27302 4020
rect 27220 3962 27302 3986
rect 28238 4020 28320 4044
rect 28238 3986 28262 4020
rect 28296 3986 28320 4020
rect 28238 3962 28320 3986
rect 29256 4020 29338 4044
rect 29256 3986 29280 4020
rect 29314 3986 29338 4020
rect 29256 3962 29338 3986
rect 30274 4020 30356 4044
rect 30274 3986 30298 4020
rect 30332 3986 30356 4020
rect 30274 3962 30356 3986
rect 31292 4020 31374 4044
rect 31292 3986 31316 4020
rect 31350 3986 31374 4020
rect 31292 3962 31374 3986
rect 32310 4020 32392 4044
rect 32310 3986 32334 4020
rect 32368 3986 32392 4020
rect 32310 3962 32392 3986
rect 33328 4020 33410 4044
rect 33328 3986 33352 4020
rect 33386 3986 33410 4020
rect 33328 3962 33410 3986
rect 13724 3714 13740 3748
rect 14296 3714 14312 3748
rect 14742 3714 14758 3748
rect 15314 3714 15330 3748
rect 15760 3714 15776 3748
rect 16332 3714 16348 3748
rect 16778 3714 16794 3748
rect 17350 3714 17366 3748
rect 17796 3714 17812 3748
rect 18368 3714 18384 3748
rect 18814 3714 18830 3748
rect 19386 3714 19402 3748
rect 19832 3714 19848 3748
rect 20404 3714 20420 3748
rect 20850 3714 20866 3748
rect 21422 3714 21438 3748
rect 21868 3714 21884 3748
rect 22440 3714 22456 3748
rect 22886 3714 22902 3748
rect 23458 3714 23474 3748
rect 23904 3714 23920 3748
rect 24476 3714 24492 3748
rect 24922 3714 24938 3748
rect 25494 3714 25510 3748
rect 25940 3714 25956 3748
rect 26512 3714 26528 3748
rect 26958 3714 26974 3748
rect 27530 3714 27546 3748
rect 27976 3714 27992 3748
rect 28548 3714 28564 3748
rect 28994 3714 29010 3748
rect 29566 3714 29582 3748
rect 30012 3714 30028 3748
rect 30584 3714 30600 3748
rect 31030 3714 31046 3748
rect 31602 3714 31618 3748
rect 32048 3714 32064 3748
rect 32620 3714 32636 3748
rect 33066 3714 33082 3748
rect 33638 3714 33654 3748
rect 17046 3712 17106 3714
rect 11602 3450 11636 3466
rect 13492 3664 13526 3680
rect 636 3382 652 3416
rect 1208 3382 1224 3416
rect 1654 3382 1670 3416
rect 2226 3382 2242 3416
rect 2672 3382 2688 3416
rect 3244 3382 3260 3416
rect 3690 3382 3706 3416
rect 4262 3382 4278 3416
rect 4708 3382 4724 3416
rect 5280 3382 5296 3416
rect 5726 3382 5742 3416
rect 6298 3382 6314 3416
rect 6744 3382 6760 3416
rect 7316 3382 7332 3416
rect 7762 3382 7778 3416
rect 8334 3382 8350 3416
rect 8780 3382 8796 3416
rect 9352 3382 9368 3416
rect 9798 3382 9814 3416
rect 10370 3382 10386 3416
rect 10816 3382 10832 3416
rect 11388 3382 11404 3416
rect 886 3230 968 3254
rect 886 3196 910 3230
rect 944 3196 968 3230
rect 886 3172 968 3196
rect 1904 3230 1986 3254
rect 1904 3196 1928 3230
rect 1962 3196 1986 3230
rect 1904 3172 1986 3196
rect 2922 3230 3004 3254
rect 2922 3196 2946 3230
rect 2980 3196 3004 3230
rect 2922 3172 3004 3196
rect 3940 3230 4022 3254
rect 3940 3196 3964 3230
rect 3998 3196 4022 3230
rect 3940 3172 4022 3196
rect 4958 3230 5040 3254
rect 4958 3196 4982 3230
rect 5016 3196 5040 3230
rect 4958 3172 5040 3196
rect 5976 3230 6058 3254
rect 5976 3196 6000 3230
rect 6034 3196 6058 3230
rect 5976 3172 6058 3196
rect 6994 3230 7076 3254
rect 6994 3196 7018 3230
rect 7052 3196 7076 3230
rect 6994 3172 7076 3196
rect 8012 3230 8094 3254
rect 8012 3196 8036 3230
rect 8070 3196 8094 3230
rect 8012 3172 8094 3196
rect 9030 3230 9112 3254
rect 9030 3196 9054 3230
rect 9088 3196 9112 3230
rect 9030 3172 9112 3196
rect 10048 3230 10130 3254
rect 10048 3196 10072 3230
rect 10106 3196 10130 3230
rect 10048 3172 10130 3196
rect 11066 3230 11148 3254
rect 11066 3196 11090 3230
rect 11124 3196 11148 3230
rect 11066 3172 11148 3196
rect 13492 3072 13526 3088
rect 14510 3664 14544 3680
rect 14510 3072 14544 3088
rect 15528 3664 15562 3680
rect 15528 3072 15562 3088
rect 16546 3664 16580 3680
rect 16546 3072 16580 3088
rect 17564 3664 17598 3680
rect 17564 3072 17598 3088
rect 18582 3664 18616 3680
rect 18582 3072 18616 3088
rect 19600 3664 19634 3680
rect 19600 3072 19634 3088
rect 20618 3664 20652 3680
rect 20618 3072 20652 3088
rect 21636 3664 21670 3680
rect 21636 3072 21670 3088
rect 22654 3664 22688 3680
rect 22654 3072 22688 3088
rect 23672 3664 23706 3680
rect 23672 3072 23706 3088
rect 24690 3664 24724 3680
rect 24690 3072 24724 3088
rect 25708 3664 25742 3680
rect 25708 3072 25742 3088
rect 26726 3664 26760 3680
rect 26726 3072 26760 3088
rect 27744 3664 27778 3680
rect 27744 3072 27778 3088
rect 28762 3664 28796 3680
rect 28762 3072 28796 3088
rect 29780 3664 29814 3680
rect 29780 3072 29814 3088
rect 30798 3664 30832 3680
rect 30798 3072 30832 3088
rect 31816 3664 31850 3680
rect 31816 3072 31850 3088
rect 32834 3664 32868 3680
rect 32834 3072 32868 3088
rect 33852 3664 33886 3680
rect 33852 3072 33886 3088
rect 21118 3038 21178 3048
rect 636 2980 652 3014
rect 1208 2980 1224 3014
rect 1654 2980 1670 3014
rect 2226 2980 2242 3014
rect 2672 2980 2688 3014
rect 3244 2980 3260 3014
rect 3690 2980 3706 3014
rect 4262 2980 4278 3014
rect 4708 2980 4724 3014
rect 5280 2980 5296 3014
rect 5726 2980 5742 3014
rect 6298 2980 6314 3014
rect 6744 2980 6760 3014
rect 7316 2980 7332 3014
rect 7762 2980 7778 3014
rect 8334 2980 8350 3014
rect 8780 2980 8796 3014
rect 9352 2980 9368 3014
rect 9798 2980 9814 3014
rect 10370 2980 10386 3014
rect 10816 2980 10832 3014
rect 11388 2980 11404 3014
rect 13724 3004 13740 3038
rect 14296 3004 14312 3038
rect 14742 3004 14758 3038
rect 15314 3004 15330 3038
rect 15760 3004 15776 3038
rect 16332 3004 16348 3038
rect 16778 3004 16794 3038
rect 17350 3004 17366 3038
rect 17796 3004 17812 3038
rect 18368 3004 18384 3038
rect 18814 3004 18830 3038
rect 19386 3004 19402 3038
rect 19832 3004 19848 3038
rect 20404 3004 20420 3038
rect 20850 3004 20866 3038
rect 21422 3004 21438 3038
rect 21868 3004 21884 3038
rect 22440 3004 22456 3038
rect 22886 3004 22902 3038
rect 23458 3004 23474 3038
rect 23904 3004 23920 3038
rect 24476 3004 24492 3038
rect 24922 3004 24938 3038
rect 25494 3004 25510 3038
rect 25940 3004 25956 3038
rect 26512 3004 26528 3038
rect 26958 3004 26974 3038
rect 27530 3004 27546 3038
rect 27976 3004 27992 3038
rect 28548 3004 28564 3038
rect 28994 3004 29010 3038
rect 29566 3004 29582 3038
rect 30012 3004 30028 3038
rect 30584 3004 30600 3038
rect 31030 3004 31046 3038
rect 31602 3004 31618 3038
rect 32048 3004 32064 3038
rect 32620 3004 32636 3038
rect 33066 3004 33082 3038
rect 33638 3004 33654 3038
rect 404 2930 438 2946
rect 404 2338 438 2354
rect 1422 2930 1456 2946
rect 1422 2338 1456 2354
rect 2440 2930 2474 2946
rect 2440 2338 2474 2354
rect 3458 2930 3492 2946
rect 3458 2338 3492 2354
rect 4476 2930 4510 2946
rect 4476 2338 4510 2354
rect 5494 2930 5528 2946
rect 5494 2338 5528 2354
rect 6512 2930 6546 2946
rect 6512 2338 6546 2354
rect 7530 2930 7564 2946
rect 7530 2338 7564 2354
rect 8548 2930 8582 2946
rect 8548 2338 8582 2354
rect 9566 2930 9600 2946
rect 9566 2338 9600 2354
rect 10584 2930 10618 2946
rect 10584 2338 10618 2354
rect 11602 2930 11636 2946
rect 13986 2784 14068 2808
rect 13986 2750 14010 2784
rect 14044 2750 14068 2784
rect 13986 2726 14068 2750
rect 15004 2784 15086 2808
rect 15004 2750 15028 2784
rect 15062 2750 15086 2784
rect 15004 2726 15086 2750
rect 16022 2784 16104 2808
rect 16022 2750 16046 2784
rect 16080 2750 16104 2784
rect 16022 2726 16104 2750
rect 17040 2784 17122 2808
rect 17040 2750 17064 2784
rect 17098 2750 17122 2784
rect 17040 2726 17122 2750
rect 18058 2784 18140 2808
rect 18058 2750 18082 2784
rect 18116 2750 18140 2784
rect 18058 2726 18140 2750
rect 19076 2784 19158 2808
rect 19076 2750 19100 2784
rect 19134 2750 19158 2784
rect 19076 2726 19158 2750
rect 20094 2784 20176 2808
rect 20094 2750 20118 2784
rect 20152 2750 20176 2784
rect 20094 2726 20176 2750
rect 21112 2784 21194 2808
rect 21112 2750 21136 2784
rect 21170 2750 21194 2784
rect 21112 2726 21194 2750
rect 22130 2784 22212 2808
rect 22130 2750 22154 2784
rect 22188 2750 22212 2784
rect 22130 2726 22212 2750
rect 23148 2784 23230 2808
rect 23148 2750 23172 2784
rect 23206 2750 23230 2784
rect 23148 2726 23230 2750
rect 24166 2784 24248 2808
rect 24166 2750 24190 2784
rect 24224 2750 24248 2784
rect 24166 2726 24248 2750
rect 25184 2784 25266 2808
rect 25184 2750 25208 2784
rect 25242 2750 25266 2784
rect 25184 2726 25266 2750
rect 26202 2784 26284 2808
rect 26202 2750 26226 2784
rect 26260 2750 26284 2784
rect 26202 2726 26284 2750
rect 27220 2784 27302 2808
rect 27220 2750 27244 2784
rect 27278 2750 27302 2784
rect 27220 2726 27302 2750
rect 28238 2784 28320 2808
rect 28238 2750 28262 2784
rect 28296 2750 28320 2784
rect 28238 2726 28320 2750
rect 29256 2784 29338 2808
rect 29256 2750 29280 2784
rect 29314 2750 29338 2784
rect 29256 2726 29338 2750
rect 30274 2784 30356 2808
rect 30274 2750 30298 2784
rect 30332 2750 30356 2784
rect 30274 2726 30356 2750
rect 31292 2784 31374 2808
rect 31292 2750 31316 2784
rect 31350 2750 31374 2784
rect 31292 2726 31374 2750
rect 32310 2784 32392 2808
rect 32310 2750 32334 2784
rect 32368 2750 32392 2784
rect 32310 2726 32392 2750
rect 33328 2784 33410 2808
rect 33328 2750 33352 2784
rect 33386 2750 33410 2784
rect 33328 2726 33410 2750
rect 13724 2480 13740 2514
rect 14296 2480 14312 2514
rect 14742 2480 14758 2514
rect 15314 2480 15330 2514
rect 15760 2480 15776 2514
rect 16332 2480 16348 2514
rect 16778 2480 16794 2514
rect 17350 2480 17366 2514
rect 17796 2480 17812 2514
rect 18368 2480 18384 2514
rect 18814 2480 18830 2514
rect 19386 2480 19402 2514
rect 19832 2480 19848 2514
rect 20404 2480 20420 2514
rect 20850 2480 20866 2514
rect 21422 2480 21438 2514
rect 21868 2480 21884 2514
rect 22440 2480 22456 2514
rect 22886 2480 22902 2514
rect 23458 2480 23474 2514
rect 23904 2480 23920 2514
rect 24476 2480 24492 2514
rect 24922 2480 24938 2514
rect 25494 2480 25510 2514
rect 25940 2480 25956 2514
rect 26512 2480 26528 2514
rect 26958 2480 26974 2514
rect 27530 2480 27546 2514
rect 27976 2480 27992 2514
rect 28548 2480 28564 2514
rect 28994 2480 29010 2514
rect 29566 2480 29582 2514
rect 30012 2480 30028 2514
rect 30584 2480 30600 2514
rect 31030 2480 31046 2514
rect 31602 2480 31618 2514
rect 32048 2480 32064 2514
rect 32620 2480 32636 2514
rect 33066 2480 33082 2514
rect 33638 2480 33654 2514
rect 17032 2478 17092 2480
rect 11602 2338 11636 2354
rect 13492 2430 13526 2446
rect 636 2270 652 2304
rect 1208 2270 1224 2304
rect 1654 2270 1670 2304
rect 2226 2270 2242 2304
rect 2672 2270 2688 2304
rect 3244 2270 3260 2304
rect 3690 2270 3706 2304
rect 4262 2270 4278 2304
rect 4708 2270 4724 2304
rect 5280 2270 5296 2304
rect 5726 2270 5742 2304
rect 6298 2270 6314 2304
rect 6744 2270 6760 2304
rect 7316 2270 7332 2304
rect 7762 2270 7778 2304
rect 8334 2270 8350 2304
rect 8780 2270 8796 2304
rect 9352 2270 9368 2304
rect 9798 2270 9814 2304
rect 10370 2270 10386 2304
rect 10816 2270 10832 2304
rect 11388 2270 11404 2304
rect 886 1888 968 1912
rect 886 1854 910 1888
rect 944 1854 968 1888
rect 886 1830 968 1854
rect 1904 1888 1986 1912
rect 1904 1854 1928 1888
rect 1962 1854 1986 1888
rect 1904 1830 1986 1854
rect 2922 1888 3004 1912
rect 2922 1854 2946 1888
rect 2980 1854 3004 1888
rect 2922 1830 3004 1854
rect 3940 1888 4022 1912
rect 3940 1854 3964 1888
rect 3998 1854 4022 1888
rect 3940 1830 4022 1854
rect 4958 1888 5040 1912
rect 4958 1854 4982 1888
rect 5016 1854 5040 1888
rect 4958 1830 5040 1854
rect 5976 1888 6058 1912
rect 5976 1854 6000 1888
rect 6034 1854 6058 1888
rect 5976 1830 6058 1854
rect 6994 1888 7076 1912
rect 6994 1854 7018 1888
rect 7052 1854 7076 1888
rect 6994 1830 7076 1854
rect 8012 1888 8094 1912
rect 8012 1854 8036 1888
rect 8070 1854 8094 1888
rect 8012 1830 8094 1854
rect 9030 1888 9112 1912
rect 9030 1854 9054 1888
rect 9088 1854 9112 1888
rect 9030 1830 9112 1854
rect 10048 1888 10130 1912
rect 10048 1854 10072 1888
rect 10106 1854 10130 1888
rect 10048 1830 10130 1854
rect 11066 1888 11148 1912
rect 11066 1854 11090 1888
rect 11124 1854 11148 1888
rect 11066 1830 11148 1854
rect 13492 1838 13526 1854
rect 14510 2430 14544 2446
rect 14510 1838 14544 1854
rect 15528 2430 15562 2446
rect 15528 1838 15562 1854
rect 16546 2430 16580 2446
rect 16546 1838 16580 1854
rect 17564 2430 17598 2446
rect 17564 1838 17598 1854
rect 18582 2430 18616 2446
rect 18582 1838 18616 1854
rect 19600 2430 19634 2446
rect 19600 1838 19634 1854
rect 20618 2430 20652 2446
rect 20618 1838 20652 1854
rect 21636 2430 21670 2446
rect 21636 1838 21670 1854
rect 22654 2430 22688 2446
rect 22654 1838 22688 1854
rect 23672 2430 23706 2446
rect 23672 1838 23706 1854
rect 24690 2430 24724 2446
rect 24690 1838 24724 1854
rect 25708 2430 25742 2446
rect 25708 1838 25742 1854
rect 26726 2430 26760 2446
rect 26726 1838 26760 1854
rect 27744 2430 27778 2446
rect 27744 1838 27778 1854
rect 28762 2430 28796 2446
rect 28762 1838 28796 1854
rect 29780 2430 29814 2446
rect 29780 1838 29814 1854
rect 30798 2430 30832 2446
rect 30798 1838 30832 1854
rect 31816 2430 31850 2446
rect 31816 1838 31850 1854
rect 32834 2430 32868 2446
rect 32834 1838 32868 1854
rect 33852 2430 33886 2446
rect 33852 1838 33886 1854
rect 15000 1804 15060 1806
rect 21112 1804 21172 1806
rect 23146 1804 23206 1806
rect 27212 1804 27272 1810
rect 31288 1804 31348 1806
rect 32304 1804 32364 1806
rect 13724 1770 13740 1804
rect 14296 1770 14312 1804
rect 14742 1770 14758 1804
rect 15314 1770 15330 1804
rect 15760 1770 15776 1804
rect 16332 1770 16348 1804
rect 16778 1770 16794 1804
rect 17350 1770 17366 1804
rect 17796 1770 17812 1804
rect 18368 1770 18384 1804
rect 18814 1770 18830 1804
rect 19386 1770 19402 1804
rect 19832 1770 19848 1804
rect 20404 1770 20420 1804
rect 20850 1770 20866 1804
rect 21422 1770 21438 1804
rect 21868 1770 21884 1804
rect 22440 1770 22456 1804
rect 22886 1770 22902 1804
rect 23458 1770 23474 1804
rect 23904 1770 23920 1804
rect 24476 1770 24492 1804
rect 24922 1770 24938 1804
rect 25494 1770 25510 1804
rect 25940 1770 25956 1804
rect 26512 1770 26528 1804
rect 26958 1770 26974 1804
rect 27530 1770 27546 1804
rect 27976 1770 27992 1804
rect 28548 1770 28564 1804
rect 28994 1770 29010 1804
rect 29566 1770 29582 1804
rect 30012 1770 30028 1804
rect 30584 1770 30600 1804
rect 31030 1770 31046 1804
rect 31602 1770 31618 1804
rect 32048 1770 32064 1804
rect 32620 1770 32636 1804
rect 33066 1770 33082 1804
rect 33638 1770 33654 1804
rect 13998 1538 14080 1562
rect 13998 1504 14022 1538
rect 14056 1504 14080 1538
rect 13998 1480 14080 1504
rect 15016 1538 15098 1562
rect 15016 1504 15040 1538
rect 15074 1504 15098 1538
rect 15016 1480 15098 1504
rect 16034 1538 16116 1562
rect 16034 1504 16058 1538
rect 16092 1504 16116 1538
rect 16034 1480 16116 1504
rect 17052 1538 17134 1562
rect 17052 1504 17076 1538
rect 17110 1504 17134 1538
rect 17052 1480 17134 1504
rect 18070 1538 18152 1562
rect 18070 1504 18094 1538
rect 18128 1504 18152 1538
rect 18070 1480 18152 1504
rect 19088 1538 19170 1562
rect 19088 1504 19112 1538
rect 19146 1504 19170 1538
rect 19088 1480 19170 1504
rect 20106 1538 20188 1562
rect 20106 1504 20130 1538
rect 20164 1504 20188 1538
rect 20106 1480 20188 1504
rect 21124 1538 21206 1562
rect 21124 1504 21148 1538
rect 21182 1504 21206 1538
rect 21124 1480 21206 1504
rect 22142 1538 22224 1562
rect 22142 1504 22166 1538
rect 22200 1504 22224 1538
rect 22142 1480 22224 1504
rect 23160 1538 23242 1562
rect 23160 1504 23184 1538
rect 23218 1504 23242 1538
rect 23160 1480 23242 1504
rect 24178 1538 24260 1562
rect 24178 1504 24202 1538
rect 24236 1504 24260 1538
rect 24178 1480 24260 1504
rect 25196 1538 25278 1562
rect 25196 1504 25220 1538
rect 25254 1504 25278 1538
rect 25196 1480 25278 1504
rect 26214 1538 26296 1562
rect 26214 1504 26238 1538
rect 26272 1504 26296 1538
rect 26214 1480 26296 1504
rect 27232 1538 27314 1562
rect 27232 1504 27256 1538
rect 27290 1504 27314 1538
rect 27232 1480 27314 1504
rect 28250 1538 28332 1562
rect 28250 1504 28274 1538
rect 28308 1504 28332 1538
rect 28250 1480 28332 1504
rect 29268 1538 29350 1562
rect 29268 1504 29292 1538
rect 29326 1504 29350 1538
rect 29268 1480 29350 1504
rect 30286 1538 30368 1562
rect 30286 1504 30310 1538
rect 30344 1504 30368 1538
rect 30286 1480 30368 1504
rect 31304 1538 31386 1562
rect 31304 1504 31328 1538
rect 31362 1504 31386 1538
rect 31304 1480 31386 1504
rect 32322 1538 32404 1562
rect 32322 1504 32346 1538
rect 32380 1504 32404 1538
rect 32322 1480 32404 1504
rect 33340 1538 33422 1562
rect 33340 1504 33364 1538
rect 33398 1504 33422 1538
rect 33340 1480 33422 1504
rect 1094 1438 1110 1472
rect 1666 1438 1682 1472
rect 2112 1438 2128 1472
rect 2684 1438 2700 1472
rect 3130 1438 3146 1472
rect 3702 1438 3718 1472
rect 4148 1438 4164 1472
rect 4720 1438 4736 1472
rect 5166 1438 5182 1472
rect 5738 1438 5754 1472
rect 6184 1438 6200 1472
rect 6756 1438 6772 1472
rect 7202 1438 7218 1472
rect 7774 1438 7790 1472
rect 8220 1438 8236 1472
rect 8792 1438 8808 1472
rect 9238 1438 9254 1472
rect 9810 1438 9826 1472
rect 10256 1438 10272 1472
rect 10828 1438 10844 1472
rect 862 1388 896 1404
rect 862 796 896 812
rect 1880 1388 1914 1404
rect 1880 796 1914 812
rect 2898 1388 2932 1404
rect 2898 796 2932 812
rect 3916 1388 3950 1404
rect 3916 796 3950 812
rect 4934 1388 4968 1404
rect 4934 796 4968 812
rect 5952 1388 5986 1404
rect 5952 796 5986 812
rect 6970 1388 7004 1404
rect 6970 796 7004 812
rect 7988 1388 8022 1404
rect 7988 796 8022 812
rect 9006 1388 9040 1404
rect 9006 796 9040 812
rect 10024 1388 10058 1404
rect 10024 796 10058 812
rect 11042 1388 11076 1404
rect 13724 1248 13740 1282
rect 14296 1248 14312 1282
rect 14742 1248 14758 1282
rect 15314 1248 15330 1282
rect 15760 1248 15776 1282
rect 16332 1248 16348 1282
rect 16778 1248 16794 1282
rect 17350 1248 17366 1282
rect 17796 1248 17812 1282
rect 18368 1248 18384 1282
rect 18814 1248 18830 1282
rect 19386 1248 19402 1282
rect 19832 1248 19848 1282
rect 20404 1248 20420 1282
rect 20850 1248 20866 1282
rect 21422 1248 21438 1282
rect 21868 1248 21884 1282
rect 22440 1248 22456 1282
rect 22886 1248 22902 1282
rect 23458 1248 23474 1282
rect 23904 1248 23920 1282
rect 24476 1248 24492 1282
rect 24922 1248 24938 1282
rect 25494 1248 25510 1282
rect 25940 1248 25956 1282
rect 26512 1248 26528 1282
rect 26958 1248 26974 1282
rect 27530 1248 27546 1282
rect 27976 1248 27992 1282
rect 28548 1248 28564 1282
rect 28994 1248 29010 1282
rect 29566 1248 29582 1282
rect 30012 1248 30028 1282
rect 30584 1248 30600 1282
rect 31030 1248 31046 1282
rect 31602 1248 31618 1282
rect 32048 1248 32064 1282
rect 32620 1248 32636 1282
rect 33066 1248 33082 1282
rect 33638 1248 33654 1282
rect 11042 796 11076 812
rect 13492 1198 13526 1214
rect 1094 728 1110 762
rect 1666 728 1682 762
rect 2112 728 2128 762
rect 2684 728 2700 762
rect 3130 728 3146 762
rect 3702 728 3718 762
rect 4148 728 4164 762
rect 4720 728 4736 762
rect 5166 728 5182 762
rect 5738 728 5754 762
rect 6184 728 6200 762
rect 6756 728 6772 762
rect 7202 728 7218 762
rect 7774 728 7790 762
rect 8220 728 8236 762
rect 8792 728 8808 762
rect 9238 728 9254 762
rect 9810 728 9826 762
rect 10256 728 10272 762
rect 10828 728 10844 762
rect 13492 606 13526 622
rect 14510 1198 14544 1214
rect 14510 606 14544 622
rect 15528 1198 15562 1214
rect 15528 606 15562 622
rect 16546 1198 16580 1214
rect 16546 606 16580 622
rect 17564 1198 17598 1214
rect 17564 606 17598 622
rect 18582 1198 18616 1214
rect 18582 606 18616 622
rect 19600 1198 19634 1214
rect 19600 606 19634 622
rect 20618 1198 20652 1214
rect 20618 606 20652 622
rect 21636 1198 21670 1214
rect 21636 606 21670 622
rect 22654 1198 22688 1214
rect 22654 606 22688 622
rect 23672 1198 23706 1214
rect 23672 606 23706 622
rect 24690 1198 24724 1214
rect 24690 606 24724 622
rect 25708 1198 25742 1214
rect 25708 606 25742 622
rect 26726 1198 26760 1214
rect 26726 606 26760 622
rect 27744 1198 27778 1214
rect 27744 606 27778 622
rect 28762 1198 28796 1214
rect 28762 606 28796 622
rect 29780 1198 29814 1214
rect 29780 606 29814 622
rect 30798 1198 30832 1214
rect 30798 606 30832 622
rect 31816 1198 31850 1214
rect 31816 606 31850 622
rect 32834 1198 32868 1214
rect 32834 606 32868 622
rect 33852 1198 33886 1214
rect 33852 606 33886 622
rect 13724 538 13740 572
rect 14296 538 14312 572
rect 14742 538 14758 572
rect 15314 538 15330 572
rect 15760 538 15776 572
rect 16332 538 16348 572
rect 16778 538 16794 572
rect 17350 538 17366 572
rect 17796 538 17812 572
rect 18368 538 18384 572
rect 18814 538 18830 572
rect 19386 538 19402 572
rect 19832 538 19848 572
rect 20404 538 20420 572
rect 20850 538 20866 572
rect 21422 538 21438 572
rect 21868 538 21884 572
rect 22440 538 22456 572
rect 22886 538 22902 572
rect 23458 538 23474 572
rect 23904 538 23920 572
rect 24476 538 24492 572
rect 24922 538 24938 572
rect 25494 538 25510 572
rect 25940 538 25956 572
rect 26512 538 26528 572
rect 26958 538 26974 572
rect 27530 538 27546 572
rect 27976 538 27992 572
rect 28548 538 28564 572
rect 28994 538 29010 572
rect 29566 538 29582 572
rect 30012 538 30028 572
rect 30584 538 30600 572
rect 31030 538 31046 572
rect 31602 538 31618 572
rect 32048 538 32064 572
rect 32620 538 32636 572
rect 33066 538 33082 572
rect 33638 538 33654 572
rect 696 442 778 466
rect 696 408 720 442
rect 754 408 778 442
rect 696 384 778 408
rect 1714 442 1796 466
rect 1714 408 1738 442
rect 1772 408 1796 442
rect 1714 384 1796 408
rect 2732 442 2814 466
rect 2732 408 2756 442
rect 2790 408 2814 442
rect 2732 384 2814 408
rect 3750 442 3832 466
rect 3750 408 3774 442
rect 3808 408 3832 442
rect 3750 384 3832 408
rect 4768 442 4850 466
rect 4768 408 4792 442
rect 4826 408 4850 442
rect 4768 384 4850 408
rect 5786 442 5868 466
rect 5786 408 5810 442
rect 5844 408 5868 442
rect 5786 384 5868 408
rect 6804 442 6886 466
rect 6804 408 6828 442
rect 6862 408 6886 442
rect 6804 384 6886 408
rect 7822 442 7904 466
rect 7822 408 7846 442
rect 7880 408 7904 442
rect 7822 384 7904 408
rect 8840 442 8922 466
rect 8840 408 8864 442
rect 8898 408 8922 442
rect 8840 384 8922 408
rect 9858 442 9940 466
rect 9858 408 9882 442
rect 9916 408 9940 442
rect 9858 384 9940 408
rect 10876 442 10958 466
rect 10876 408 10900 442
rect 10934 408 10958 442
rect 10876 384 10958 408
rect 13986 360 14068 384
rect 13986 326 14010 360
rect 14044 326 14068 360
rect 13986 302 14068 326
rect 15004 360 15086 384
rect 15004 326 15028 360
rect 15062 326 15086 360
rect 15004 302 15086 326
rect 16022 360 16104 384
rect 16022 326 16046 360
rect 16080 326 16104 360
rect 16022 302 16104 326
rect 17040 360 17122 384
rect 17040 326 17064 360
rect 17098 326 17122 360
rect 17040 302 17122 326
rect 18058 360 18140 384
rect 18058 326 18082 360
rect 18116 326 18140 360
rect 18058 302 18140 326
rect 19076 360 19158 384
rect 19076 326 19100 360
rect 19134 326 19158 360
rect 19076 302 19158 326
rect 20094 360 20176 384
rect 20094 326 20118 360
rect 20152 326 20176 360
rect 20094 302 20176 326
rect 21112 360 21194 384
rect 21112 326 21136 360
rect 21170 326 21194 360
rect 21112 302 21194 326
rect 22130 360 22212 384
rect 22130 326 22154 360
rect 22188 326 22212 360
rect 22130 302 22212 326
rect 23148 360 23230 384
rect 23148 326 23172 360
rect 23206 326 23230 360
rect 23148 302 23230 326
rect 24166 360 24248 384
rect 24166 326 24190 360
rect 24224 326 24248 360
rect 24166 302 24248 326
rect 25184 360 25266 384
rect 25184 326 25208 360
rect 25242 326 25266 360
rect 25184 302 25266 326
rect 26202 360 26284 384
rect 26202 326 26226 360
rect 26260 326 26284 360
rect 26202 302 26284 326
rect 27220 360 27302 384
rect 27220 326 27244 360
rect 27278 326 27302 360
rect 27220 302 27302 326
rect 28238 360 28320 384
rect 28238 326 28262 360
rect 28296 326 28320 360
rect 28238 302 28320 326
rect 29256 360 29338 384
rect 29256 326 29280 360
rect 29314 326 29338 360
rect 29256 302 29338 326
rect 30274 360 30356 384
rect 30274 326 30298 360
rect 30332 326 30356 360
rect 30274 302 30356 326
rect 31292 360 31374 384
rect 31292 326 31316 360
rect 31350 326 31374 360
rect 31292 302 31374 326
rect 32310 360 32392 384
rect 32310 326 32334 360
rect 32368 326 32392 360
rect 32310 302 32392 326
rect 33328 360 33410 384
rect 33328 326 33352 360
rect 33386 326 33410 360
rect 33328 302 33410 326
rect -1410 -682 -1310 -520
rect 35734 -682 35834 -520
<< viali >>
rect 11390 30762 11452 30862
rect 11452 30762 35572 30862
rect 35572 30762 35634 30862
rect 11290 16812 11390 30242
rect 17694 28061 18158 28095
rect 18712 28061 19176 28095
rect 19730 28061 20194 28095
rect 20748 28061 21212 28095
rect 21766 28061 22230 28095
rect 22784 28061 23248 28095
rect 23802 28061 24266 28095
rect 24820 28061 25284 28095
rect 25838 28061 26302 28095
rect 26856 28061 27320 28095
rect 27874 28061 28338 28095
rect 28892 28061 29356 28095
rect 29910 28061 30374 28095
rect 30928 28061 31392 28095
rect 31946 28061 32410 28095
rect 32964 28061 33428 28095
rect 17400 27426 17434 28002
rect 18418 27426 18452 28002
rect 19436 27426 19470 28002
rect 20454 27426 20488 28002
rect 21472 27426 21506 28002
rect 22490 27426 22524 28002
rect 23508 27426 23542 28002
rect 24526 27426 24560 28002
rect 25544 27426 25578 28002
rect 26562 27426 26596 28002
rect 27580 27426 27614 28002
rect 28598 27426 28632 28002
rect 29616 27426 29650 28002
rect 30634 27426 30668 28002
rect 31652 27426 31686 28002
rect 32670 27426 32704 28002
rect 33688 27426 33722 28002
rect 17694 27333 18158 27367
rect 18712 27333 19176 27367
rect 19730 27333 20194 27367
rect 20748 27333 21212 27367
rect 21766 27333 22230 27367
rect 22784 27333 23248 27367
rect 23802 27333 24266 27367
rect 24820 27333 25284 27367
rect 25838 27333 26302 27367
rect 26856 27333 27320 27367
rect 27874 27333 28338 27367
rect 28892 27333 29356 27367
rect 29910 27333 30374 27367
rect 30928 27333 31392 27367
rect 31946 27333 32410 27367
rect 32964 27333 33428 27367
rect 17694 26925 18158 26959
rect 18712 26925 19176 26959
rect 19730 26925 20194 26959
rect 20748 26925 21212 26959
rect 21766 26925 22230 26959
rect 22784 26925 23248 26959
rect 23802 26925 24266 26959
rect 24820 26925 25284 26959
rect 25838 26925 26302 26959
rect 26856 26925 27320 26959
rect 27874 26925 28338 26959
rect 28892 26925 29356 26959
rect 29910 26925 30374 26959
rect 30928 26925 31392 26959
rect 31946 26925 32410 26959
rect 32964 26925 33428 26959
rect 17400 26290 17434 26866
rect 18418 26290 18452 26866
rect 19436 26290 19470 26866
rect 20454 26290 20488 26866
rect 21472 26290 21506 26866
rect 22490 26290 22524 26866
rect 23508 26290 23542 26866
rect 24526 26290 24560 26866
rect 25544 26290 25578 26866
rect 26562 26290 26596 26866
rect 27580 26290 27614 26866
rect 28598 26290 28632 26866
rect 29616 26290 29650 26866
rect 30634 26290 30668 26866
rect 31652 26290 31686 26866
rect 32670 26290 32704 26866
rect 33688 26290 33722 26866
rect 17694 26197 18158 26231
rect 18712 26197 19176 26231
rect 19730 26197 20194 26231
rect 20748 26197 21212 26231
rect 21766 26197 22230 26231
rect 22784 26197 23248 26231
rect 23802 26197 24266 26231
rect 24820 26197 25284 26231
rect 25838 26197 26302 26231
rect 26856 26197 27320 26231
rect 27874 26197 28338 26231
rect 28892 26197 29356 26231
rect 29910 26197 30374 26231
rect 30928 26197 31392 26231
rect 31946 26197 32410 26231
rect 32964 26197 33428 26231
rect 17694 25789 18158 25823
rect 18712 25789 19176 25823
rect 19730 25789 20194 25823
rect 20748 25789 21212 25823
rect 21766 25789 22230 25823
rect 22784 25789 23248 25823
rect 23802 25789 24266 25823
rect 24820 25789 25284 25823
rect 25838 25789 26302 25823
rect 26856 25789 27320 25823
rect 27874 25789 28338 25823
rect 28892 25789 29356 25823
rect 29910 25789 30374 25823
rect 30928 25789 31392 25823
rect 31946 25789 32410 25823
rect 32964 25789 33428 25823
rect 17400 25154 17434 25730
rect 18418 25154 18452 25730
rect 19436 25154 19470 25730
rect 20454 25154 20488 25730
rect 21472 25154 21506 25730
rect 22490 25154 22524 25730
rect 23508 25154 23542 25730
rect 24526 25154 24560 25730
rect 25544 25154 25578 25730
rect 26562 25154 26596 25730
rect 27580 25154 27614 25730
rect 28598 25154 28632 25730
rect 29616 25154 29650 25730
rect 30634 25154 30668 25730
rect 31652 25154 31686 25730
rect 32670 25154 32704 25730
rect 33688 25154 33722 25730
rect 17694 25061 18158 25095
rect 18712 25061 19176 25095
rect 19730 25061 20194 25095
rect 20748 25061 21212 25095
rect 21766 25061 22230 25095
rect 22784 25061 23248 25095
rect 23802 25061 24266 25095
rect 24820 25061 25284 25095
rect 25838 25061 26302 25095
rect 26856 25061 27320 25095
rect 27874 25061 28338 25095
rect 28892 25061 29356 25095
rect 29910 25061 30374 25095
rect 30928 25061 31392 25095
rect 31946 25061 32410 25095
rect 32964 25061 33428 25095
rect 18888 24151 19352 24185
rect 19906 24151 20370 24185
rect 20924 24151 21388 24185
rect 21942 24151 22406 24185
rect 22960 24151 23424 24185
rect 23978 24151 24442 24185
rect 24996 24151 25460 24185
rect 26014 24151 26478 24185
rect 27032 24151 27496 24185
rect 28050 24151 28514 24185
rect 29068 24151 29532 24185
rect 30086 24151 30550 24185
rect 31104 24151 31568 24185
rect 32122 24151 32586 24185
rect 18594 23516 18628 24092
rect 19612 23516 19646 24092
rect 20630 23516 20664 24092
rect 21648 23516 21682 24092
rect 22666 23516 22700 24092
rect 23684 23516 23718 24092
rect 24702 23516 24736 24092
rect 25720 23516 25754 24092
rect 26738 23516 26772 24092
rect 27756 23516 27790 24092
rect 28774 23516 28808 24092
rect 29792 23516 29826 24092
rect 30810 23516 30844 24092
rect 31828 23516 31862 24092
rect 32846 23516 32880 24092
rect 18888 23423 19352 23457
rect 19906 23423 20370 23457
rect 20924 23423 21388 23457
rect 21942 23423 22406 23457
rect 22960 23423 23424 23457
rect 23978 23423 24442 23457
rect 24996 23423 25460 23457
rect 26014 23423 26478 23457
rect 27032 23423 27496 23457
rect 28050 23423 28514 23457
rect 29068 23423 29532 23457
rect 30086 23423 30550 23457
rect 31104 23423 31568 23457
rect 32122 23423 32586 23457
rect 18888 23119 19352 23153
rect 19906 23119 20370 23153
rect 20924 23119 21388 23153
rect 21942 23119 22406 23153
rect 22960 23119 23424 23153
rect 23978 23119 24442 23153
rect 24996 23119 25460 23153
rect 26014 23119 26478 23153
rect 27032 23119 27496 23153
rect 28050 23119 28514 23153
rect 29068 23119 29532 23153
rect 30086 23119 30550 23153
rect 31104 23119 31568 23153
rect 32122 23119 32586 23153
rect 18594 22484 18628 23060
rect 19612 22484 19646 23060
rect 20630 22484 20664 23060
rect 21648 22484 21682 23060
rect 22666 22484 22700 23060
rect 23684 22484 23718 23060
rect 24702 22484 24736 23060
rect 25720 22484 25754 23060
rect 26738 22484 26772 23060
rect 27756 22484 27790 23060
rect 28774 22484 28808 23060
rect 29792 22484 29826 23060
rect 30810 22484 30844 23060
rect 31828 22484 31862 23060
rect 32846 22484 32880 23060
rect 18888 22391 19352 22425
rect 19906 22391 20370 22425
rect 20924 22391 21388 22425
rect 21942 22391 22406 22425
rect 22960 22391 23424 22425
rect 23978 22391 24442 22425
rect 24996 22391 25460 22425
rect 26014 22391 26478 22425
rect 27032 22391 27496 22425
rect 28050 22391 28514 22425
rect 29068 22391 29532 22425
rect 30086 22391 30550 22425
rect 31104 22391 31568 22425
rect 32122 22391 32586 22425
rect 18680 21515 19144 21549
rect 19698 21515 20162 21549
rect 20716 21515 21180 21549
rect 21734 21515 22198 21549
rect 22752 21515 23216 21549
rect 23770 21515 24234 21549
rect 24788 21515 25252 21549
rect 25806 21515 26270 21549
rect 26824 21515 27288 21549
rect 27842 21515 28306 21549
rect 28860 21515 29324 21549
rect 29878 21515 30342 21549
rect 30896 21515 31360 21549
rect 31914 21515 32378 21549
rect 32932 21515 33396 21549
rect 13376 21411 13840 21445
rect 14394 21411 14858 21445
rect 15412 21411 15876 21445
rect 16430 21411 16894 21445
rect 13082 20776 13116 21352
rect 14100 20776 14134 21352
rect 15118 20776 15152 21352
rect 16136 20776 16170 21352
rect 17154 20776 17188 21352
rect 18386 20880 18420 21456
rect 19404 20880 19438 21456
rect 20422 20880 20456 21456
rect 21440 20880 21474 21456
rect 22458 20880 22492 21456
rect 23476 20880 23510 21456
rect 24494 20880 24528 21456
rect 25512 20880 25546 21456
rect 26530 20880 26564 21456
rect 27548 20880 27582 21456
rect 28566 20880 28600 21456
rect 29584 20880 29618 21456
rect 30602 20880 30636 21456
rect 31620 20880 31654 21456
rect 32638 20880 32672 21456
rect 33656 20880 33690 21456
rect 18680 20787 19144 20821
rect 19698 20787 20162 20821
rect 20716 20787 21180 20821
rect 21734 20787 22198 20821
rect 22752 20787 23216 20821
rect 23770 20787 24234 20821
rect 24788 20787 25252 20821
rect 25806 20787 26270 20821
rect 26824 20787 27288 20821
rect 27842 20787 28306 20821
rect 28860 20787 29324 20821
rect 29878 20787 30342 20821
rect 30896 20787 31360 20821
rect 31914 20787 32378 20821
rect 32932 20787 33396 20821
rect 13376 20683 13840 20717
rect 14394 20683 14858 20717
rect 15412 20683 15876 20717
rect 16430 20683 16894 20717
rect 13376 20379 13840 20413
rect 14394 20379 14858 20413
rect 15412 20379 15876 20413
rect 16430 20379 16894 20413
rect 13082 19744 13116 20320
rect 14100 19744 14134 20320
rect 15118 19744 15152 20320
rect 16136 19744 16170 20320
rect 17154 19744 17188 20320
rect 18680 20259 19144 20293
rect 19698 20259 20162 20293
rect 20716 20259 21180 20293
rect 21734 20259 22198 20293
rect 22752 20259 23216 20293
rect 23770 20259 24234 20293
rect 24788 20259 25252 20293
rect 25806 20259 26270 20293
rect 26824 20259 27288 20293
rect 27842 20259 28306 20293
rect 28860 20259 29324 20293
rect 29878 20259 30342 20293
rect 30896 20259 31360 20293
rect 31914 20259 32378 20293
rect 32932 20259 33396 20293
rect 13376 19651 13840 19685
rect 14394 19651 14858 19685
rect 15412 19651 15876 19685
rect 16430 19651 16894 19685
rect 18386 19624 18420 20200
rect 19404 19624 19438 20200
rect 20422 19624 20456 20200
rect 21440 19624 21474 20200
rect 22458 19624 22492 20200
rect 23476 19624 23510 20200
rect 24494 19624 24528 20200
rect 25512 19624 25546 20200
rect 26530 19624 26564 20200
rect 27548 19624 27582 20200
rect 28566 19624 28600 20200
rect 29584 19624 29618 20200
rect 30602 19624 30636 20200
rect 31620 19624 31654 20200
rect 32638 19624 32672 20200
rect 33656 19624 33690 20200
rect 18680 19531 19144 19565
rect 19698 19531 20162 19565
rect 20716 19531 21180 19565
rect 21734 19531 22198 19565
rect 22752 19531 23216 19565
rect 23770 19531 24234 19565
rect 24788 19531 25252 19565
rect 25806 19531 26270 19565
rect 26824 19531 27288 19565
rect 27842 19531 28306 19565
rect 28860 19531 29324 19565
rect 29878 19531 30342 19565
rect 30896 19531 31360 19565
rect 31914 19531 32378 19565
rect 32932 19531 33396 19565
rect 13376 19347 13840 19381
rect 14394 19347 14858 19381
rect 15412 19347 15876 19381
rect 16430 19347 16894 19381
rect 13082 18712 13116 19288
rect 14100 18712 14134 19288
rect 15118 18712 15152 19288
rect 16136 18712 16170 19288
rect 17154 18712 17188 19288
rect 18680 19003 19144 19037
rect 19698 19003 20162 19037
rect 20716 19003 21180 19037
rect 21734 19003 22198 19037
rect 22752 19003 23216 19037
rect 23770 19003 24234 19037
rect 24788 19003 25252 19037
rect 25806 19003 26270 19037
rect 26824 19003 27288 19037
rect 27842 19003 28306 19037
rect 28860 19003 29324 19037
rect 29878 19003 30342 19037
rect 30896 19003 31360 19037
rect 31914 19003 32378 19037
rect 32932 19003 33396 19037
rect 13376 18619 13840 18653
rect 14394 18619 14858 18653
rect 15412 18619 15876 18653
rect 16430 18619 16894 18653
rect 18386 18368 18420 18944
rect 19404 18368 19438 18944
rect 20422 18368 20456 18944
rect 21440 18368 21474 18944
rect 22458 18368 22492 18944
rect 23476 18368 23510 18944
rect 24494 18368 24528 18944
rect 25512 18368 25546 18944
rect 26530 18368 26564 18944
rect 27548 18368 27582 18944
rect 28566 18368 28600 18944
rect 29584 18368 29618 18944
rect 30602 18368 30636 18944
rect 31620 18368 31654 18944
rect 32638 18368 32672 18944
rect 33656 18368 33690 18944
rect 13376 18315 13840 18349
rect 14394 18315 14858 18349
rect 15412 18315 15876 18349
rect 16430 18315 16894 18349
rect 18680 18275 19144 18309
rect 19698 18275 20162 18309
rect 20716 18275 21180 18309
rect 21734 18275 22198 18309
rect 22752 18275 23216 18309
rect 23770 18275 24234 18309
rect 24788 18275 25252 18309
rect 25806 18275 26270 18309
rect 26824 18275 27288 18309
rect 27842 18275 28306 18309
rect 28860 18275 29324 18309
rect 29878 18275 30342 18309
rect 30896 18275 31360 18309
rect 31914 18275 32378 18309
rect 32932 18275 33396 18309
rect 13082 17680 13116 18256
rect 14100 17680 14134 18256
rect 15118 17680 15152 18256
rect 16136 17680 16170 18256
rect 17154 17680 17188 18256
rect 18680 17747 19144 17781
rect 19698 17747 20162 17781
rect 20716 17747 21180 17781
rect 21734 17747 22198 17781
rect 22752 17747 23216 17781
rect 23770 17747 24234 17781
rect 24788 17747 25252 17781
rect 25806 17747 26270 17781
rect 26824 17747 27288 17781
rect 27842 17747 28306 17781
rect 28860 17747 29324 17781
rect 29878 17747 30342 17781
rect 30896 17747 31360 17781
rect 31914 17747 32378 17781
rect 32932 17747 33396 17781
rect 13376 17587 13840 17621
rect 14394 17587 14858 17621
rect 15412 17587 15876 17621
rect 16430 17587 16894 17621
rect 18386 17112 18420 17688
rect 19404 17112 19438 17688
rect 20422 17112 20456 17688
rect 21440 17112 21474 17688
rect 22458 17112 22492 17688
rect 23476 17112 23510 17688
rect 24494 17112 24528 17688
rect 25512 17112 25546 17688
rect 26530 17112 26564 17688
rect 27548 17112 27582 17688
rect 28566 17112 28600 17688
rect 29584 17112 29618 17688
rect 30602 17112 30636 17688
rect 31620 17112 31654 17688
rect 32638 17112 32672 17688
rect 33656 17112 33690 17688
rect 18680 17019 19144 17053
rect 19698 17019 20162 17053
rect 20716 17019 21180 17053
rect 21734 17019 22198 17053
rect 22752 17019 23216 17053
rect 23770 17019 24234 17053
rect 24788 17019 25252 17053
rect 25806 17019 26270 17053
rect 26824 17019 27288 17053
rect 27842 17019 28306 17053
rect 28860 17019 29324 17053
rect 29878 17019 30342 17053
rect 30896 17019 31360 17053
rect 31914 17019 32378 17053
rect 32932 17019 33396 17053
rect -12234 16309 -12014 16310
rect -10742 16309 -10540 16310
rect -9634 16309 -9414 16310
rect -8142 16309 -7940 16310
rect -12234 16276 -12184 16309
rect -12184 16276 -12014 16309
rect -10742 16276 -10566 16309
rect -10566 16276 -10540 16309
rect -10506 16213 -10470 16214
rect -12282 15640 -12280 16212
rect -12280 15640 -12246 16212
rect -12246 15640 -12244 16212
rect -12062 16173 -11978 16207
rect -11804 16173 -11720 16207
rect -11546 16173 -11462 16207
rect -11288 16173 -11204 16207
rect -11030 16173 -10946 16207
rect -10772 16173 -10688 16207
rect -12166 15738 -12132 16114
rect -11908 15738 -11874 16114
rect -11650 15738 -11616 16114
rect -11392 15738 -11358 16114
rect -11134 15738 -11100 16114
rect -10876 15738 -10842 16114
rect -10618 15738 -10584 16114
rect -12062 15645 -11978 15679
rect -11804 15645 -11720 15679
rect -11546 15645 -11462 15679
rect -11288 15645 -11204 15679
rect -11030 15645 -10946 15679
rect -10772 15645 -10688 15679
rect -10506 15639 -10504 16213
rect -10504 15639 -10470 16213
rect -9634 16276 -9584 16309
rect -9584 16276 -9414 16309
rect -8142 16276 -7966 16309
rect -7966 16276 -7940 16309
rect -7906 16213 -7870 16214
rect -10367 15773 -10333 15807
rect -10275 15773 -10241 15807
rect -10183 15773 -10149 15807
rect -10506 15638 -10470 15639
rect -10742 15577 -10540 15578
rect -12234 15543 -12184 15576
rect -12184 15543 -12014 15576
rect -10742 15544 -10566 15577
rect -10566 15544 -10540 15577
rect -9682 15640 -9680 16212
rect -9680 15640 -9646 16212
rect -9646 15640 -9644 16212
rect -9462 16173 -9378 16207
rect -9204 16173 -9120 16207
rect -8946 16173 -8862 16207
rect -8688 16173 -8604 16207
rect -8430 16173 -8346 16207
rect -8172 16173 -8088 16207
rect -9566 15738 -9532 16114
rect -9308 15738 -9274 16114
rect -9050 15738 -9016 16114
rect -8792 15738 -8758 16114
rect -8534 15738 -8500 16114
rect -8276 15738 -8242 16114
rect -8018 15738 -7984 16114
rect -9462 15645 -9378 15679
rect -9204 15645 -9120 15679
rect -8946 15645 -8862 15679
rect -8688 15645 -8604 15679
rect -8430 15645 -8346 15679
rect -8172 15645 -8088 15679
rect -7906 15639 -7904 16213
rect -7904 15639 -7870 16213
rect 35634 16812 35734 30242
rect 11390 16192 11452 16292
rect 11452 16192 35572 16292
rect 35572 16192 35634 16292
rect -7767 15773 -7733 15807
rect -7675 15773 -7641 15807
rect -7583 15773 -7549 15807
rect -7317 15773 -7283 15807
rect -7225 15773 -7191 15807
rect -7133 15773 -7099 15807
rect -7906 15638 -7870 15639
rect -8142 15577 -7940 15578
rect -9634 15543 -9584 15576
rect -9584 15543 -9414 15576
rect -8142 15544 -7966 15577
rect -7966 15544 -7940 15577
rect -12234 15542 -12014 15543
rect -9634 15542 -9414 15543
rect -10337 15436 -10289 15484
rect -10233 15495 -10187 15506
rect -10233 15466 -10200 15495
rect -10200 15466 -10187 15495
rect -7737 15436 -7689 15484
rect -7633 15495 -7587 15506
rect -7633 15466 -7600 15495
rect -7600 15466 -7587 15495
rect -7288 15458 -7240 15506
rect -7184 15495 -7136 15510
rect -7184 15462 -7150 15495
rect -7150 15462 -7136 15495
rect -12210 15376 -12002 15378
rect -10738 15376 -10540 15380
rect -12210 15342 -12184 15376
rect -12184 15342 -12002 15376
rect -10738 15342 -10566 15376
rect -10566 15342 -10540 15376
rect -12210 15340 -12002 15342
rect -9610 15376 -9402 15378
rect -8138 15376 -7940 15380
rect -12282 14924 -12280 15280
rect -12280 14924 -12246 15280
rect -12062 15240 -11978 15274
rect -11804 15240 -11720 15274
rect -11546 15240 -11462 15274
rect -11288 15240 -11204 15274
rect -11030 15240 -10946 15274
rect -10772 15240 -10688 15274
rect -12166 15014 -12132 15190
rect -11908 15014 -11874 15190
rect -11650 15014 -11616 15190
rect -11392 15014 -11358 15190
rect -11134 15014 -11100 15190
rect -10876 15014 -10842 15190
rect -10618 15014 -10584 15190
rect -12062 14930 -11978 14964
rect -11804 14930 -11720 14964
rect -11546 14930 -11462 14964
rect -11288 14930 -11204 14964
rect -11030 14930 -10946 14964
rect -10772 14930 -10688 14964
rect -10506 14924 -10504 15280
rect -10504 14924 -10470 15280
rect -10470 14924 -10468 15280
rect -9610 15342 -9584 15376
rect -9584 15342 -9402 15376
rect -8138 15342 -7966 15376
rect -7966 15342 -7940 15376
rect -9610 15340 -9402 15342
rect -10367 15229 -10333 15263
rect -10275 15229 -10241 15263
rect -10183 15229 -10149 15263
rect -9682 14924 -9680 15280
rect -9680 14924 -9646 15280
rect -9462 15240 -9378 15274
rect -9204 15240 -9120 15274
rect -8946 15240 -8862 15274
rect -8688 15240 -8604 15274
rect -8430 15240 -8346 15274
rect -8172 15240 -8088 15274
rect -9566 15014 -9532 15190
rect -9308 15014 -9274 15190
rect -9050 15014 -9016 15190
rect -8792 15014 -8758 15190
rect -8534 15014 -8500 15190
rect -8276 15014 -8242 15190
rect -8018 15014 -7984 15190
rect -9462 14930 -9378 14964
rect -9204 14930 -9120 14964
rect -8946 14930 -8862 14964
rect -8688 14930 -8604 14964
rect -8430 14930 -8346 14964
rect -8172 14930 -8088 14964
rect -7906 14924 -7904 15280
rect -7904 14924 -7870 15280
rect -7870 14924 -7868 15280
rect -7767 15229 -7733 15263
rect -7675 15229 -7641 15263
rect -7583 15229 -7549 15263
rect -7317 15229 -7283 15263
rect -7225 15229 -7191 15263
rect -7133 15229 -7099 15263
rect -1310 15262 -1248 15362
rect -1248 15262 35672 15362
rect 35672 15262 35734 15362
rect -12212 14862 -12004 14864
rect -12212 14828 -12184 14862
rect -12184 14828 -12004 14862
rect -10740 14828 -10566 14862
rect -10566 14828 -10538 14862
rect -9612 14862 -9404 14864
rect -9612 14828 -9584 14862
rect -9584 14828 -9404 14862
rect -8140 14828 -7966 14862
rect -7966 14828 -7938 14862
rect -10740 14826 -10538 14828
rect -8140 14826 -7938 14828
rect 13788 14542 14252 14576
rect 14806 14542 15270 14576
rect 15824 14542 16288 14576
rect 16842 14542 17306 14576
rect 17860 14542 18324 14576
rect 18878 14542 19342 14576
rect 19896 14542 20360 14576
rect 20914 14542 21378 14576
rect 21932 14542 22396 14576
rect 22950 14542 23414 14576
rect 23968 14542 24432 14576
rect 24986 14542 25450 14576
rect 26004 14542 26468 14576
rect 27022 14542 27486 14576
rect 28040 14542 28504 14576
rect 29058 14542 29522 14576
rect 30076 14542 30540 14576
rect 31094 14542 31558 14576
rect 32112 14542 32576 14576
rect 33130 14542 33594 14576
rect -1410 210 -1310 14470
rect 2022 14066 2486 14100
rect 3040 14066 3504 14100
rect 4058 14066 4522 14100
rect 5076 14066 5540 14100
rect 6094 14066 6558 14100
rect 7112 14066 7576 14100
rect 8130 14066 8594 14100
rect 9148 14066 9612 14100
rect 10166 14066 10630 14100
rect 1728 13440 1762 14016
rect 2746 13440 2780 14016
rect 3764 13440 3798 14016
rect 4782 13440 4816 14016
rect 5800 13440 5834 14016
rect 6818 13440 6852 14016
rect 7836 13440 7870 14016
rect 8854 13440 8888 14016
rect 9872 13440 9906 14016
rect 10890 13440 10924 14016
rect 13494 13916 13528 14492
rect 14512 13916 14546 14492
rect 15530 13916 15564 14492
rect 16548 13916 16582 14492
rect 17566 13916 17600 14492
rect 18584 13916 18618 14492
rect 19602 13916 19636 14492
rect 20620 13916 20654 14492
rect 21638 13916 21672 14492
rect 22656 13916 22690 14492
rect 23674 13916 23708 14492
rect 24692 13916 24726 14492
rect 25710 13916 25744 14492
rect 26728 13916 26762 14492
rect 27746 13916 27780 14492
rect 28764 13916 28798 14492
rect 29782 13916 29816 14492
rect 30800 13916 30834 14492
rect 31818 13916 31852 14492
rect 32836 13916 32870 14492
rect 33854 13916 33888 14492
rect 13788 13832 14252 13866
rect 14806 13832 15270 13866
rect 15824 13832 16288 13866
rect 16842 13832 17306 13866
rect 17860 13832 18324 13866
rect 18878 13832 19342 13866
rect 19896 13832 20360 13866
rect 20914 13832 21378 13866
rect 21932 13832 22396 13866
rect 22950 13832 23414 13866
rect 23968 13832 24432 13866
rect 24986 13832 25450 13866
rect 26004 13832 26468 13866
rect 27022 13832 27486 13866
rect 28040 13832 28504 13866
rect 29058 13832 29522 13866
rect 30076 13832 30540 13866
rect 31094 13832 31558 13866
rect 32112 13832 32576 13866
rect 33130 13832 33594 13866
rect 13788 13724 14252 13758
rect 14806 13724 15270 13758
rect 15824 13724 16288 13758
rect 16842 13724 17306 13758
rect 17860 13724 18324 13758
rect 18878 13724 19342 13758
rect 19896 13724 20360 13758
rect 20914 13724 21378 13758
rect 21932 13724 22396 13758
rect 22950 13724 23414 13758
rect 23968 13724 24432 13758
rect 24986 13724 25450 13758
rect 26004 13724 26468 13758
rect 27022 13724 27486 13758
rect 28040 13724 28504 13758
rect 29058 13724 29522 13758
rect 30076 13724 30540 13758
rect 31094 13724 31558 13758
rect 32112 13724 32576 13758
rect 33130 13724 33594 13758
rect 2022 13356 2486 13390
rect 3040 13356 3504 13390
rect 2022 13248 2486 13282
rect 4058 13356 4522 13390
rect 3040 13248 3504 13282
rect 5076 13356 5540 13390
rect 4058 13248 4522 13282
rect 6094 13356 6558 13390
rect 5076 13248 5540 13282
rect 7112 13356 7576 13390
rect 6094 13248 6558 13282
rect 8130 13356 8594 13390
rect 7112 13248 7576 13282
rect 9148 13356 9612 13390
rect 8130 13248 8594 13282
rect 10166 13356 10630 13390
rect 9148 13248 9612 13282
rect 10166 13248 10630 13282
rect 1728 12622 1762 13198
rect 2746 12622 2780 13198
rect 3764 12622 3798 13198
rect 4782 12622 4816 13198
rect 5800 12622 5834 13198
rect 6818 12622 6852 13198
rect 7836 12622 7870 13198
rect 8854 12622 8888 13198
rect 9872 12622 9906 13198
rect 10890 12622 10924 13198
rect 13494 13098 13528 13674
rect 14512 13098 14546 13674
rect 15530 13098 15564 13674
rect 16548 13098 16582 13674
rect 17566 13098 17600 13674
rect 18584 13098 18618 13674
rect 19602 13098 19636 13674
rect 20620 13098 20654 13674
rect 21638 13098 21672 13674
rect 22656 13098 22690 13674
rect 23674 13098 23708 13674
rect 24692 13098 24726 13674
rect 25710 13098 25744 13674
rect 26728 13098 26762 13674
rect 27746 13098 27780 13674
rect 28764 13098 28798 13674
rect 29782 13098 29816 13674
rect 30800 13098 30834 13674
rect 31818 13098 31852 13674
rect 32836 13098 32870 13674
rect 33854 13098 33888 13674
rect 13788 13014 14252 13048
rect 14806 13014 15270 13048
rect 15824 13014 16288 13048
rect 16842 13014 17306 13048
rect 17860 13014 18324 13048
rect 18878 13014 19342 13048
rect 19896 13014 20360 13048
rect 20914 13014 21378 13048
rect 21932 13014 22396 13048
rect 22950 13014 23414 13048
rect 23968 13014 24432 13048
rect 24986 13014 25450 13048
rect 26004 13014 26468 13048
rect 27022 13014 27486 13048
rect 28040 13014 28504 13048
rect 29058 13014 29522 13048
rect 30076 13014 30540 13048
rect 31094 13014 31558 13048
rect 32112 13014 32576 13048
rect 33130 13014 33594 13048
rect 2022 12538 2486 12572
rect 3040 12538 3504 12572
rect 2022 12430 2486 12464
rect 4058 12538 4522 12572
rect 3040 12430 3504 12464
rect 5076 12538 5540 12572
rect 4058 12430 4522 12464
rect 6094 12538 6558 12572
rect 5076 12430 5540 12464
rect 7112 12538 7576 12572
rect 6094 12430 6558 12464
rect 8130 12538 8594 12572
rect 7112 12430 7576 12464
rect 9148 12538 9612 12572
rect 8130 12430 8594 12464
rect 10166 12538 10630 12572
rect 9148 12430 9612 12464
rect 10166 12430 10630 12464
rect 1728 11804 1762 12380
rect 2746 11804 2780 12380
rect 3764 11804 3798 12380
rect 4782 11804 4816 12380
rect 5800 11804 5834 12380
rect 6818 11804 6852 12380
rect 7836 11804 7870 12380
rect 8854 11804 8888 12380
rect 9872 11804 9906 12380
rect 10890 11804 10924 12380
rect 13788 12346 14252 12380
rect 14806 12346 15270 12380
rect 15824 12346 16288 12380
rect 16842 12346 17306 12380
rect 17860 12346 18324 12380
rect 18878 12346 19342 12380
rect 19896 12346 20360 12380
rect 20914 12346 21378 12380
rect 21932 12346 22396 12380
rect 22950 12346 23414 12380
rect 23968 12346 24432 12380
rect 24986 12346 25450 12380
rect 26004 12346 26468 12380
rect 27022 12346 27486 12380
rect 28040 12346 28504 12380
rect 29058 12346 29522 12380
rect 30076 12346 30540 12380
rect 31094 12346 31558 12380
rect 32112 12346 32576 12380
rect 33130 12346 33594 12380
rect 2022 11720 2486 11754
rect 3040 11720 3504 11754
rect 2022 11612 2486 11646
rect 4058 11720 4522 11754
rect 3040 11612 3504 11646
rect 5076 11720 5540 11754
rect 4058 11612 4522 11646
rect 6094 11720 6558 11754
rect 5076 11612 5540 11646
rect 7112 11720 7576 11754
rect 6094 11612 6558 11646
rect 8130 11720 8594 11754
rect 7112 11612 7576 11646
rect 9148 11720 9612 11754
rect 8130 11612 8594 11646
rect 10166 11720 10630 11754
rect 9148 11612 9612 11646
rect 13494 11720 13528 12296
rect 14512 11720 14546 12296
rect 15530 11720 15564 12296
rect 16548 11720 16582 12296
rect 17566 11720 17600 12296
rect 18584 11720 18618 12296
rect 19602 11720 19636 12296
rect 20620 11720 20654 12296
rect 21638 11720 21672 12296
rect 22656 11720 22690 12296
rect 23674 11720 23708 12296
rect 24692 11720 24726 12296
rect 25710 11720 25744 12296
rect 26728 11720 26762 12296
rect 27746 11720 27780 12296
rect 28764 11720 28798 12296
rect 29782 11720 29816 12296
rect 30800 11720 30834 12296
rect 31818 11720 31852 12296
rect 32836 11720 32870 12296
rect 33854 11720 33888 12296
rect 10166 11612 10630 11646
rect 13788 11636 14252 11670
rect 14806 11636 15270 11670
rect 15824 11636 16288 11670
rect 16842 11636 17306 11670
rect 17860 11636 18324 11670
rect 18878 11636 19342 11670
rect 19896 11636 20360 11670
rect 20914 11636 21378 11670
rect 21932 11636 22396 11670
rect 22950 11636 23414 11670
rect 23968 11636 24432 11670
rect 24986 11636 25450 11670
rect 26004 11636 26468 11670
rect 27022 11636 27486 11670
rect 28040 11636 28504 11670
rect 29058 11636 29522 11670
rect 30076 11636 30540 11670
rect 31094 11636 31558 11670
rect 32112 11636 32576 11670
rect 33130 11636 33594 11670
rect 1728 10986 1762 11562
rect 2746 10986 2780 11562
rect 3764 10986 3798 11562
rect 4782 10986 4816 11562
rect 5800 10986 5834 11562
rect 6818 10986 6852 11562
rect 7836 10986 7870 11562
rect 8854 10986 8888 11562
rect 9872 10986 9906 11562
rect 10890 10986 10924 11562
rect 13788 11114 14252 11148
rect 14806 11114 15270 11148
rect 15824 11114 16288 11148
rect 16842 11114 17306 11148
rect 17860 11114 18324 11148
rect 18878 11114 19342 11148
rect 19896 11114 20360 11148
rect 20914 11114 21378 11148
rect 21932 11114 22396 11148
rect 22950 11114 23414 11148
rect 23968 11114 24432 11148
rect 24986 11114 25450 11148
rect 26004 11114 26468 11148
rect 27022 11114 27486 11148
rect 28040 11114 28504 11148
rect 29058 11114 29522 11148
rect 30076 11114 30540 11148
rect 31094 11114 31558 11148
rect 32112 11114 32576 11148
rect 33130 11114 33594 11148
rect 2022 10902 2486 10936
rect 3040 10902 3504 10936
rect 2022 10794 2486 10828
rect 4058 10902 4522 10936
rect 3040 10794 3504 10828
rect 5076 10902 5540 10936
rect 4058 10794 4522 10828
rect 6094 10902 6558 10936
rect 5076 10794 5540 10828
rect 7112 10902 7576 10936
rect 6094 10794 6558 10828
rect 8130 10902 8594 10936
rect 7112 10794 7576 10828
rect 9148 10902 9612 10936
rect 8130 10794 8594 10828
rect 10166 10902 10630 10936
rect 9148 10794 9612 10828
rect 10166 10794 10630 10828
rect 1728 10168 1762 10744
rect 2746 10168 2780 10744
rect 3764 10168 3798 10744
rect 4782 10168 4816 10744
rect 5800 10168 5834 10744
rect 6818 10168 6852 10744
rect 7836 10168 7870 10744
rect 8854 10168 8888 10744
rect 9872 10168 9906 10744
rect 10890 10168 10924 10744
rect 13494 10488 13528 11064
rect 14512 10488 14546 11064
rect 15530 10488 15564 11064
rect 16548 10488 16582 11064
rect 17566 10488 17600 11064
rect 18584 10488 18618 11064
rect 19602 10488 19636 11064
rect 20620 10488 20654 11064
rect 21638 10488 21672 11064
rect 22656 10488 22690 11064
rect 23674 10488 23708 11064
rect 24692 10488 24726 11064
rect 25710 10488 25744 11064
rect 26728 10488 26762 11064
rect 27746 10488 27780 11064
rect 28764 10488 28798 11064
rect 29782 10488 29816 11064
rect 30800 10488 30834 11064
rect 31818 10488 31852 11064
rect 32836 10488 32870 11064
rect 33854 10488 33888 11064
rect 13788 10404 14252 10438
rect 14806 10404 15270 10438
rect 15824 10404 16288 10438
rect 16842 10404 17306 10438
rect 17860 10404 18324 10438
rect 18878 10404 19342 10438
rect 19896 10404 20360 10438
rect 20914 10404 21378 10438
rect 21932 10404 22396 10438
rect 22950 10404 23414 10438
rect 23968 10404 24432 10438
rect 24986 10404 25450 10438
rect 26004 10404 26468 10438
rect 27022 10404 27486 10438
rect 28040 10404 28504 10438
rect 29058 10404 29522 10438
rect 30076 10404 30540 10438
rect 31094 10404 31558 10438
rect 32112 10404 32576 10438
rect 33130 10404 33594 10438
rect 2022 10084 2486 10118
rect 3040 10084 3504 10118
rect 2022 9976 2486 10010
rect 4058 10084 4522 10118
rect 3040 9976 3504 10010
rect 5076 10084 5540 10118
rect 4058 9976 4522 10010
rect 6094 10084 6558 10118
rect 5076 9976 5540 10010
rect 7112 10084 7576 10118
rect 6094 9976 6558 10010
rect 8130 10084 8594 10118
rect 7112 9976 7576 10010
rect 9148 10084 9612 10118
rect 8130 9976 8594 10010
rect 10166 10084 10630 10118
rect 9148 9976 9612 10010
rect 10166 9976 10630 10010
rect 1728 9350 1762 9926
rect 2746 9350 2780 9926
rect 3764 9350 3798 9926
rect 4782 9350 4816 9926
rect 5800 9350 5834 9926
rect 6818 9350 6852 9926
rect 7836 9350 7870 9926
rect 8854 9350 8888 9926
rect 9872 9350 9906 9926
rect 10890 9350 10924 9926
rect 13786 9880 14250 9914
rect 14804 9880 15268 9914
rect 15822 9880 16286 9914
rect 16840 9880 17304 9914
rect 17858 9880 18322 9914
rect 18876 9880 19340 9914
rect 19894 9880 20358 9914
rect 20912 9880 21376 9914
rect 21930 9880 22394 9914
rect 22948 9880 23412 9914
rect 23966 9880 24430 9914
rect 24984 9880 25448 9914
rect 26002 9880 26466 9914
rect 27020 9880 27484 9914
rect 28038 9880 28502 9914
rect 29056 9880 29520 9914
rect 30074 9880 30538 9914
rect 31092 9880 31556 9914
rect 32110 9880 32574 9914
rect 33128 9880 33592 9914
rect 2022 9266 2486 9300
rect 3040 9266 3504 9300
rect 2022 9158 2486 9192
rect 4058 9266 4522 9300
rect 3040 9158 3504 9192
rect 5076 9266 5540 9300
rect 4058 9158 4522 9192
rect 6094 9266 6558 9300
rect 5076 9158 5540 9192
rect 7112 9266 7576 9300
rect 6094 9158 6558 9192
rect 8130 9266 8594 9300
rect 7112 9158 7576 9192
rect 9148 9266 9612 9300
rect 8130 9158 8594 9192
rect 10166 9266 10630 9300
rect 9148 9158 9612 9192
rect 13492 9254 13526 9830
rect 14510 9254 14544 9830
rect 15528 9254 15562 9830
rect 16546 9254 16580 9830
rect 17564 9254 17598 9830
rect 18582 9254 18616 9830
rect 19600 9254 19634 9830
rect 20618 9254 20652 9830
rect 21636 9254 21670 9830
rect 22654 9254 22688 9830
rect 23672 9254 23706 9830
rect 24690 9254 24724 9830
rect 25708 9254 25742 9830
rect 26726 9254 26760 9830
rect 27744 9254 27778 9830
rect 28762 9254 28796 9830
rect 29780 9254 29814 9830
rect 30798 9254 30832 9830
rect 31816 9254 31850 9830
rect 32834 9254 32868 9830
rect 33852 9254 33886 9830
rect 10166 9158 10630 9192
rect 13786 9170 14250 9204
rect 14804 9170 15268 9204
rect 15822 9170 16286 9204
rect 16840 9170 17304 9204
rect 17858 9170 18322 9204
rect 18876 9170 19340 9204
rect 19894 9170 20358 9204
rect 20912 9170 21376 9204
rect 21930 9170 22394 9204
rect 22948 9170 23412 9204
rect 23966 9170 24430 9204
rect 24984 9170 25448 9204
rect 26002 9170 26466 9204
rect 27020 9170 27484 9204
rect 28038 9170 28502 9204
rect 29056 9170 29520 9204
rect 30074 9170 30538 9204
rect 31092 9170 31556 9204
rect 32110 9170 32574 9204
rect 33128 9170 33592 9204
rect 1728 8532 1762 9108
rect 2746 8532 2780 9108
rect 3764 8532 3798 9108
rect 4782 8532 4816 9108
rect 5800 8532 5834 9108
rect 6818 8532 6852 9108
rect 7836 8532 7870 9108
rect 8854 8532 8888 9108
rect 9872 8532 9906 9108
rect 10890 8532 10924 9108
rect 13786 8646 14250 8680
rect 14804 8646 15268 8680
rect 15822 8646 16286 8680
rect 16840 8646 17304 8680
rect 17858 8646 18322 8680
rect 18876 8646 19340 8680
rect 19894 8646 20358 8680
rect 20912 8646 21376 8680
rect 21930 8646 22394 8680
rect 22948 8646 23412 8680
rect 23966 8646 24430 8680
rect 24984 8646 25448 8680
rect 26002 8646 26466 8680
rect 27020 8646 27484 8680
rect 28038 8646 28502 8680
rect 29056 8646 29520 8680
rect 30074 8646 30538 8680
rect 31092 8646 31556 8680
rect 32110 8646 32574 8680
rect 33128 8646 33592 8680
rect 2022 8448 2486 8482
rect 3040 8448 3504 8482
rect 2022 8340 2486 8374
rect 4058 8448 4522 8482
rect 3040 8340 3504 8374
rect 5076 8448 5540 8482
rect 4058 8340 4522 8374
rect 6094 8448 6558 8482
rect 5076 8340 5540 8374
rect 7112 8448 7576 8482
rect 6094 8340 6558 8374
rect 8130 8448 8594 8482
rect 7112 8340 7576 8374
rect 9148 8448 9612 8482
rect 8130 8340 8594 8374
rect 10166 8448 10630 8482
rect 9148 8340 9612 8374
rect 10166 8340 10630 8374
rect 1728 7714 1762 8290
rect 2746 7714 2780 8290
rect 3764 7714 3798 8290
rect 4782 7714 4816 8290
rect 5800 7714 5834 8290
rect 6818 7714 6852 8290
rect 7836 7714 7870 8290
rect 8854 7714 8888 8290
rect 9872 7714 9906 8290
rect 10890 7714 10924 8290
rect 13492 8020 13526 8596
rect 14510 8020 14544 8596
rect 15528 8020 15562 8596
rect 16546 8020 16580 8596
rect 17564 8020 17598 8596
rect 18582 8020 18616 8596
rect 19600 8020 19634 8596
rect 20618 8020 20652 8596
rect 21636 8020 21670 8596
rect 22654 8020 22688 8596
rect 23672 8020 23706 8596
rect 24690 8020 24724 8596
rect 25708 8020 25742 8596
rect 26726 8020 26760 8596
rect 27744 8020 27778 8596
rect 28762 8020 28796 8596
rect 29780 8020 29814 8596
rect 30798 8020 30832 8596
rect 31816 8020 31850 8596
rect 32834 8020 32868 8596
rect 33852 8020 33886 8596
rect 13786 7936 14250 7970
rect 14804 7936 15268 7970
rect 15822 7936 16286 7970
rect 16840 7936 17304 7970
rect 17858 7936 18322 7970
rect 18876 7936 19340 7970
rect 19894 7936 20358 7970
rect 20912 7936 21376 7970
rect 21930 7936 22394 7970
rect 22948 7936 23412 7970
rect 23966 7936 24430 7970
rect 24984 7936 25448 7970
rect 26002 7936 26466 7970
rect 27020 7936 27484 7970
rect 28038 7936 28502 7970
rect 29056 7936 29520 7970
rect 30074 7936 30538 7970
rect 31092 7936 31556 7970
rect 32110 7936 32574 7970
rect 33128 7936 33592 7970
rect 2022 7630 2486 7664
rect 3040 7630 3504 7664
rect 4058 7630 4522 7664
rect 5076 7630 5540 7664
rect 6094 7630 6558 7664
rect 7112 7630 7576 7664
rect 8130 7630 8594 7664
rect 9148 7630 9612 7664
rect 10166 7630 10630 7664
rect 13786 7414 14250 7448
rect 14804 7414 15268 7448
rect 15822 7414 16286 7448
rect 16840 7414 17304 7448
rect 17858 7414 18322 7448
rect 18876 7414 19340 7448
rect 19894 7414 20358 7448
rect 20912 7414 21376 7448
rect 21930 7414 22394 7448
rect 22948 7414 23412 7448
rect 23966 7414 24430 7448
rect 24984 7414 25448 7448
rect 26002 7414 26466 7448
rect 27020 7414 27484 7448
rect 28038 7414 28502 7448
rect 29056 7414 29520 7448
rect 30074 7414 30538 7448
rect 31092 7414 31556 7448
rect 32110 7414 32574 7448
rect 33128 7414 33592 7448
rect 13492 6788 13526 7364
rect 14510 6788 14544 7364
rect 15528 6788 15562 7364
rect 16546 6788 16580 7364
rect 17564 6788 17598 7364
rect 18582 6788 18616 7364
rect 19600 6788 19634 7364
rect 20618 6788 20652 7364
rect 21636 6788 21670 7364
rect 22654 6788 22688 7364
rect 23672 6788 23706 7364
rect 24690 6788 24724 7364
rect 25708 6788 25742 7364
rect 26726 6788 26760 7364
rect 27744 6788 27778 7364
rect 28762 6788 28796 7364
rect 29780 6788 29814 7364
rect 30798 6788 30832 7364
rect 31816 6788 31850 7364
rect 32834 6788 32868 7364
rect 33852 6788 33886 7364
rect 13786 6704 14250 6738
rect 14804 6704 15268 6738
rect 15822 6704 16286 6738
rect 16840 6704 17304 6738
rect 17858 6704 18322 6738
rect 18876 6704 19340 6738
rect 19894 6704 20358 6738
rect 20912 6704 21376 6738
rect 21930 6704 22394 6738
rect 22948 6704 23412 6738
rect 23966 6704 24430 6738
rect 24984 6704 25448 6738
rect 26002 6704 26466 6738
rect 27020 6704 27484 6738
rect 28038 6704 28502 6738
rect 29056 6704 29520 6738
rect 30074 6704 30538 6738
rect 31092 6704 31556 6738
rect 32110 6704 32574 6738
rect 33128 6704 33592 6738
rect 698 6316 1162 6350
rect 1716 6316 2180 6350
rect 2734 6316 3198 6350
rect 3752 6316 4216 6350
rect 4770 6316 5234 6350
rect 5788 6316 6252 6350
rect 6806 6316 7270 6350
rect 7824 6316 8288 6350
rect 8842 6316 9306 6350
rect 9860 6316 10324 6350
rect 10878 6316 11342 6350
rect 404 5690 438 6266
rect 1422 5690 1456 6266
rect 2440 5690 2474 6266
rect 3458 5690 3492 6266
rect 4476 5690 4510 6266
rect 5494 5690 5528 6266
rect 6512 5690 6546 6266
rect 7530 5690 7564 6266
rect 8548 5690 8582 6266
rect 9566 5690 9600 6266
rect 10584 5690 10618 6266
rect 11602 5690 11636 6266
rect 13786 6180 14250 6214
rect 14804 6180 15268 6214
rect 15822 6180 16286 6214
rect 16840 6180 17304 6214
rect 17858 6180 18322 6214
rect 18876 6180 19340 6214
rect 19894 6180 20358 6214
rect 20912 6180 21376 6214
rect 21930 6180 22394 6214
rect 22948 6180 23412 6214
rect 23966 6180 24430 6214
rect 24984 6180 25448 6214
rect 26002 6180 26466 6214
rect 27020 6180 27484 6214
rect 28038 6180 28502 6214
rect 29056 6180 29520 6214
rect 30074 6180 30538 6214
rect 31092 6180 31556 6214
rect 32110 6180 32574 6214
rect 33128 6180 33592 6214
rect 698 5606 1162 5640
rect 1716 5606 2180 5640
rect 2734 5606 3198 5640
rect 3752 5606 4216 5640
rect 4770 5606 5234 5640
rect 5788 5606 6252 5640
rect 6806 5606 7270 5640
rect 7824 5606 8288 5640
rect 8842 5606 9306 5640
rect 9860 5606 10324 5640
rect 10878 5606 11342 5640
rect 13492 5554 13526 6130
rect 14510 5554 14544 6130
rect 15528 5554 15562 6130
rect 16546 5554 16580 6130
rect 17564 5554 17598 6130
rect 18582 5554 18616 6130
rect 19600 5554 19634 6130
rect 20618 5554 20652 6130
rect 21636 5554 21670 6130
rect 22654 5554 22688 6130
rect 23672 5554 23706 6130
rect 24690 5554 24724 6130
rect 25708 5554 25742 6130
rect 26726 5554 26760 6130
rect 27744 5554 27778 6130
rect 28762 5554 28796 6130
rect 29780 5554 29814 6130
rect 30798 5554 30832 6130
rect 31816 5554 31850 6130
rect 32834 5554 32868 6130
rect 33852 5554 33886 6130
rect 13786 5470 14250 5504
rect 14804 5470 15268 5504
rect 15822 5470 16286 5504
rect 16840 5470 17304 5504
rect 17858 5470 18322 5504
rect 18876 5470 19340 5504
rect 19894 5470 20358 5504
rect 20912 5470 21376 5504
rect 21930 5470 22394 5504
rect 22948 5470 23412 5504
rect 23966 5470 24430 5504
rect 24984 5470 25448 5504
rect 26002 5470 26466 5504
rect 27020 5470 27484 5504
rect 28038 5470 28502 5504
rect 29056 5470 29520 5504
rect 30074 5470 30538 5504
rect 31092 5470 31556 5504
rect 32110 5470 32574 5504
rect 33128 5470 33592 5504
rect 698 5204 1162 5238
rect 1716 5204 2180 5238
rect 2734 5204 3198 5238
rect 3752 5204 4216 5238
rect 4770 5204 5234 5238
rect 5788 5204 6252 5238
rect 6806 5204 7270 5238
rect 7824 5204 8288 5238
rect 8842 5204 9306 5238
rect 9860 5204 10324 5238
rect 10878 5204 11342 5238
rect 404 4578 438 5154
rect 1422 4578 1456 5154
rect 2440 4578 2474 5154
rect 3458 4578 3492 5154
rect 4476 4578 4510 5154
rect 5494 4578 5528 5154
rect 6512 4578 6546 5154
rect 7530 4578 7564 5154
rect 8548 4578 8582 5154
rect 9566 4578 9600 5154
rect 10584 4578 10618 5154
rect 11602 4578 11636 5154
rect 13786 4946 14250 4980
rect 14804 4946 15268 4980
rect 15822 4946 16286 4980
rect 16840 4946 17304 4980
rect 17858 4946 18322 4980
rect 18876 4946 19340 4980
rect 19894 4946 20358 4980
rect 20912 4946 21376 4980
rect 21930 4946 22394 4980
rect 22948 4946 23412 4980
rect 23966 4946 24430 4980
rect 24984 4946 25448 4980
rect 26002 4946 26466 4980
rect 27020 4946 27484 4980
rect 28038 4946 28502 4980
rect 29056 4946 29520 4980
rect 30074 4946 30538 4980
rect 31092 4946 31556 4980
rect 32110 4946 32574 4980
rect 33128 4946 33592 4980
rect 698 4494 1162 4528
rect 1716 4494 2180 4528
rect 2734 4494 3198 4528
rect 3752 4494 4216 4528
rect 4770 4494 5234 4528
rect 5788 4494 6252 4528
rect 6806 4494 7270 4528
rect 7824 4494 8288 4528
rect 8842 4494 9306 4528
rect 9860 4494 10324 4528
rect 10878 4494 11342 4528
rect 13492 4320 13526 4896
rect 14510 4320 14544 4896
rect 15528 4320 15562 4896
rect 16546 4320 16580 4896
rect 17564 4320 17598 4896
rect 18582 4320 18616 4896
rect 19600 4320 19634 4896
rect 20618 4320 20652 4896
rect 21636 4320 21670 4896
rect 22654 4320 22688 4896
rect 23672 4320 23706 4896
rect 24690 4320 24724 4896
rect 25708 4320 25742 4896
rect 26726 4320 26760 4896
rect 27744 4320 27778 4896
rect 28762 4320 28796 4896
rect 29780 4320 29814 4896
rect 30798 4320 30832 4896
rect 31816 4320 31850 4896
rect 32834 4320 32868 4896
rect 33852 4320 33886 4896
rect 13786 4236 14250 4270
rect 14804 4236 15268 4270
rect 15822 4236 16286 4270
rect 16840 4236 17304 4270
rect 17858 4236 18322 4270
rect 18876 4236 19340 4270
rect 19894 4236 20358 4270
rect 20912 4236 21376 4270
rect 21930 4236 22394 4270
rect 22948 4236 23412 4270
rect 23966 4236 24430 4270
rect 24984 4236 25448 4270
rect 26002 4236 26466 4270
rect 27020 4236 27484 4270
rect 28038 4236 28502 4270
rect 29056 4236 29520 4270
rect 30074 4236 30538 4270
rect 31092 4236 31556 4270
rect 32110 4236 32574 4270
rect 33128 4236 33592 4270
rect 698 4092 1162 4126
rect 1716 4092 2180 4126
rect 2734 4092 3198 4126
rect 3752 4092 4216 4126
rect 4770 4092 5234 4126
rect 5788 4092 6252 4126
rect 6806 4092 7270 4126
rect 7824 4092 8288 4126
rect 8842 4092 9306 4126
rect 9860 4092 10324 4126
rect 10878 4092 11342 4126
rect 404 3466 438 4042
rect 1422 3466 1456 4042
rect 2440 3466 2474 4042
rect 3458 3466 3492 4042
rect 4476 3466 4510 4042
rect 5494 3466 5528 4042
rect 6512 3466 6546 4042
rect 7530 3466 7564 4042
rect 8548 3466 8582 4042
rect 9566 3466 9600 4042
rect 10584 3466 10618 4042
rect 11602 3466 11636 4042
rect 13786 3714 14250 3748
rect 14804 3714 15268 3748
rect 15822 3714 16286 3748
rect 16840 3714 17304 3748
rect 17858 3714 18322 3748
rect 18876 3714 19340 3748
rect 19894 3714 20358 3748
rect 20912 3714 21376 3748
rect 21930 3714 22394 3748
rect 22948 3714 23412 3748
rect 23966 3714 24430 3748
rect 24984 3714 25448 3748
rect 26002 3714 26466 3748
rect 27020 3714 27484 3748
rect 28038 3714 28502 3748
rect 29056 3714 29520 3748
rect 30074 3714 30538 3748
rect 31092 3714 31556 3748
rect 32110 3714 32574 3748
rect 33128 3714 33592 3748
rect 698 3382 1162 3416
rect 1716 3382 2180 3416
rect 2734 3382 3198 3416
rect 3752 3382 4216 3416
rect 4770 3382 5234 3416
rect 5788 3382 6252 3416
rect 6806 3382 7270 3416
rect 7824 3382 8288 3416
rect 8842 3382 9306 3416
rect 9860 3382 10324 3416
rect 10878 3382 11342 3416
rect 13492 3088 13526 3664
rect 14510 3088 14544 3664
rect 15528 3088 15562 3664
rect 16546 3088 16580 3664
rect 17564 3088 17598 3664
rect 18582 3088 18616 3664
rect 19600 3088 19634 3664
rect 20618 3088 20652 3664
rect 21636 3088 21670 3664
rect 22654 3088 22688 3664
rect 23672 3088 23706 3664
rect 24690 3088 24724 3664
rect 25708 3088 25742 3664
rect 26726 3088 26760 3664
rect 27744 3088 27778 3664
rect 28762 3088 28796 3664
rect 29780 3088 29814 3664
rect 30798 3088 30832 3664
rect 31816 3088 31850 3664
rect 32834 3088 32868 3664
rect 33852 3088 33886 3664
rect 698 2980 1162 3014
rect 1716 2980 2180 3014
rect 2734 2980 3198 3014
rect 3752 2980 4216 3014
rect 4770 2980 5234 3014
rect 5788 2980 6252 3014
rect 6806 2980 7270 3014
rect 7824 2980 8288 3014
rect 8842 2980 9306 3014
rect 9860 2980 10324 3014
rect 10878 2980 11342 3014
rect 13786 3004 14250 3038
rect 14804 3004 15268 3038
rect 15822 3004 16286 3038
rect 16840 3004 17304 3038
rect 17858 3004 18322 3038
rect 18876 3004 19340 3038
rect 19894 3004 20358 3038
rect 20912 3004 21376 3038
rect 21930 3004 22394 3038
rect 22948 3004 23412 3038
rect 23966 3004 24430 3038
rect 24984 3004 25448 3038
rect 26002 3004 26466 3038
rect 27020 3004 27484 3038
rect 28038 3004 28502 3038
rect 29056 3004 29520 3038
rect 30074 3004 30538 3038
rect 31092 3004 31556 3038
rect 32110 3004 32574 3038
rect 33128 3004 33592 3038
rect 404 2354 438 2930
rect 1422 2354 1456 2930
rect 2440 2354 2474 2930
rect 3458 2354 3492 2930
rect 4476 2354 4510 2930
rect 5494 2354 5528 2930
rect 6512 2354 6546 2930
rect 7530 2354 7564 2930
rect 8548 2354 8582 2930
rect 9566 2354 9600 2930
rect 10584 2354 10618 2930
rect 11602 2354 11636 2930
rect 13786 2480 14250 2514
rect 14804 2480 15268 2514
rect 15822 2480 16286 2514
rect 16840 2480 17304 2514
rect 17858 2480 18322 2514
rect 18876 2480 19340 2514
rect 19894 2480 20358 2514
rect 20912 2480 21376 2514
rect 21930 2480 22394 2514
rect 22948 2480 23412 2514
rect 23966 2480 24430 2514
rect 24984 2480 25448 2514
rect 26002 2480 26466 2514
rect 27020 2480 27484 2514
rect 28038 2480 28502 2514
rect 29056 2480 29520 2514
rect 30074 2480 30538 2514
rect 31092 2480 31556 2514
rect 32110 2480 32574 2514
rect 33128 2480 33592 2514
rect 698 2270 1162 2304
rect 1716 2270 2180 2304
rect 2734 2270 3198 2304
rect 3752 2270 4216 2304
rect 4770 2270 5234 2304
rect 5788 2270 6252 2304
rect 6806 2270 7270 2304
rect 7824 2270 8288 2304
rect 8842 2270 9306 2304
rect 9860 2270 10324 2304
rect 10878 2270 11342 2304
rect 13492 1854 13526 2430
rect 14510 1854 14544 2430
rect 15528 1854 15562 2430
rect 16546 1854 16580 2430
rect 17564 1854 17598 2430
rect 18582 1854 18616 2430
rect 19600 1854 19634 2430
rect 20618 1854 20652 2430
rect 21636 1854 21670 2430
rect 22654 1854 22688 2430
rect 23672 1854 23706 2430
rect 24690 1854 24724 2430
rect 25708 1854 25742 2430
rect 26726 1854 26760 2430
rect 27744 1854 27778 2430
rect 28762 1854 28796 2430
rect 29780 1854 29814 2430
rect 30798 1854 30832 2430
rect 31816 1854 31850 2430
rect 32834 1854 32868 2430
rect 33852 1854 33886 2430
rect 13786 1770 14250 1804
rect 14804 1770 15268 1804
rect 15822 1770 16286 1804
rect 16840 1770 17304 1804
rect 17858 1770 18322 1804
rect 18876 1770 19340 1804
rect 19894 1770 20358 1804
rect 20912 1770 21376 1804
rect 21930 1770 22394 1804
rect 22948 1770 23412 1804
rect 23966 1770 24430 1804
rect 24984 1770 25448 1804
rect 26002 1770 26466 1804
rect 27020 1770 27484 1804
rect 28038 1770 28502 1804
rect 29056 1770 29520 1804
rect 30074 1770 30538 1804
rect 31092 1770 31556 1804
rect 32110 1770 32574 1804
rect 33128 1770 33592 1804
rect 1156 1438 1620 1472
rect 2174 1438 2638 1472
rect 3192 1438 3656 1472
rect 4210 1438 4674 1472
rect 5228 1438 5692 1472
rect 6246 1438 6710 1472
rect 7264 1438 7728 1472
rect 8282 1438 8746 1472
rect 9300 1438 9764 1472
rect 10318 1438 10782 1472
rect 862 812 896 1388
rect 1880 812 1914 1388
rect 2898 812 2932 1388
rect 3916 812 3950 1388
rect 4934 812 4968 1388
rect 5952 812 5986 1388
rect 6970 812 7004 1388
rect 7988 812 8022 1388
rect 9006 812 9040 1388
rect 10024 812 10058 1388
rect 11042 812 11076 1388
rect 13786 1248 14250 1282
rect 14804 1248 15268 1282
rect 15822 1248 16286 1282
rect 16840 1248 17304 1282
rect 17858 1248 18322 1282
rect 18876 1248 19340 1282
rect 19894 1248 20358 1282
rect 20912 1248 21376 1282
rect 21930 1248 22394 1282
rect 22948 1248 23412 1282
rect 23966 1248 24430 1282
rect 24984 1248 25448 1282
rect 26002 1248 26466 1282
rect 27020 1248 27484 1282
rect 28038 1248 28502 1282
rect 29056 1248 29520 1282
rect 30074 1248 30538 1282
rect 31092 1248 31556 1282
rect 32110 1248 32574 1282
rect 33128 1248 33592 1282
rect 1156 728 1620 762
rect 2174 728 2638 762
rect 3192 728 3656 762
rect 4210 728 4674 762
rect 5228 728 5692 762
rect 6246 728 6710 762
rect 7264 728 7728 762
rect 8282 728 8746 762
rect 9300 728 9764 762
rect 10318 728 10782 762
rect 13492 622 13526 1198
rect 14510 622 14544 1198
rect 15528 622 15562 1198
rect 16546 622 16580 1198
rect 17564 622 17598 1198
rect 18582 622 18616 1198
rect 19600 622 19634 1198
rect 20618 622 20652 1198
rect 21636 622 21670 1198
rect 22654 622 22688 1198
rect 23672 622 23706 1198
rect 24690 622 24724 1198
rect 25708 622 25742 1198
rect 26726 622 26760 1198
rect 27744 622 27778 1198
rect 28762 622 28796 1198
rect 29780 622 29814 1198
rect 30798 622 30832 1198
rect 31816 622 31850 1198
rect 32834 622 32868 1198
rect 33852 622 33886 1198
rect 13786 538 14250 572
rect 14804 538 15268 572
rect 15822 538 16286 572
rect 16840 538 17304 572
rect 17858 538 18322 572
rect 18876 538 19340 572
rect 19894 538 20358 572
rect 20912 538 21376 572
rect 21930 538 22394 572
rect 22948 538 23412 572
rect 23966 538 24430 572
rect 24984 538 25448 572
rect 26002 538 26466 572
rect 27020 538 27484 572
rect 28038 538 28502 572
rect 29056 538 29520 572
rect 30074 538 30538 572
rect 31092 538 31556 572
rect 32110 538 32574 572
rect 33128 538 33592 572
rect 35734 210 35834 14470
rect -1310 -682 -1248 -582
rect -1248 -682 35672 -582
rect 35672 -682 35734 -582
<< metal1 >>
rect 11284 30862 35740 30868
rect 11284 30762 11390 30862
rect 35634 30762 35740 30862
rect 11284 30756 35740 30762
rect -4458 30288 -4398 30294
rect -4458 16436 -4398 30228
rect 11284 30242 11396 30756
rect 11996 30456 12006 30756
rect 35018 30456 35028 30756
rect 11284 16812 11290 30242
rect 11390 16812 11396 30242
rect 14910 30374 31790 30406
rect 14910 30160 14973 30374
rect 31758 30160 31790 30374
rect 14910 30138 14960 30160
rect 15020 30138 15396 30160
rect 15456 30138 15834 30160
rect 15894 30138 16268 30160
rect 16328 30140 31790 30160
rect 35628 30242 35740 30756
rect 16328 30138 19264 30140
rect 19424 28664 19484 30140
rect 21460 28664 21520 30140
rect 21964 28664 22024 30140
rect 22472 28664 22532 30140
rect 22984 28664 23044 30140
rect 23498 28664 23558 30140
rect 25530 28664 25590 30140
rect 27570 28664 27630 30140
rect 28060 28664 28120 30140
rect 28580 28664 28640 30140
rect 29088 28664 29148 30140
rect 29602 28664 29662 30140
rect 31638 28664 31698 30140
rect 19424 28604 31698 28664
rect 18892 28398 18898 28458
rect 18958 28398 18964 28458
rect 17386 28182 18464 28242
rect 17386 28002 17446 28182
rect 17890 28101 17950 28182
rect 17682 28095 18170 28101
rect 17682 28061 17694 28095
rect 18158 28061 18170 28095
rect 17682 28055 18170 28061
rect 17386 27962 17400 28002
rect 17394 27426 17400 27962
rect 17434 27962 17446 28002
rect 18404 28002 18464 28182
rect 18898 28101 18958 28398
rect 19424 28212 19484 28604
rect 19974 28398 19980 28458
rect 20040 28398 20046 28458
rect 20932 28398 20938 28458
rect 20998 28398 21004 28458
rect 19418 28152 19424 28212
rect 19484 28152 19490 28212
rect 18700 28095 19188 28101
rect 18700 28061 18712 28095
rect 19176 28061 19188 28095
rect 18700 28055 19188 28061
rect 18404 27976 18418 28002
rect 17434 27426 17440 27962
rect 18412 27462 18418 27976
rect 17394 27414 17440 27426
rect 18406 27426 18418 27462
rect 18452 27976 18464 28002
rect 19424 28002 19484 28152
rect 19980 28101 20040 28398
rect 20938 28101 20998 28398
rect 21460 28212 21520 28604
rect 21454 28152 21460 28212
rect 21520 28152 21526 28212
rect 19718 28095 20206 28101
rect 19718 28061 19730 28095
rect 20194 28061 20206 28095
rect 19718 28055 20206 28061
rect 20736 28095 21224 28101
rect 20736 28061 20748 28095
rect 21212 28061 21224 28095
rect 20736 28055 21224 28061
rect 20938 28052 20998 28055
rect 19424 27978 19436 28002
rect 18452 27462 18458 27976
rect 19430 27466 19436 27978
rect 18452 27426 18466 27462
rect 17682 27367 18170 27373
rect 17682 27333 17694 27367
rect 18158 27333 18170 27367
rect 17682 27327 18170 27333
rect 18406 27280 18466 27426
rect 19426 27426 19436 27466
rect 19470 27978 19484 28002
rect 20448 28002 20494 28014
rect 19470 27466 19476 27978
rect 19470 27426 19486 27466
rect 20448 27454 20454 28002
rect 18910 27373 18970 27374
rect 18700 27367 19188 27373
rect 18700 27333 18712 27367
rect 19176 27333 19188 27367
rect 18700 27327 19188 27333
rect 17236 27220 17242 27280
rect 17302 27220 17308 27280
rect 18400 27220 18406 27280
rect 18466 27220 18472 27280
rect 17106 27016 17112 27076
rect 17172 27016 17178 27076
rect 15098 24832 15104 24892
rect 15164 24832 15170 24892
rect 12926 21516 14148 21576
rect 12926 19600 12986 21516
rect 13068 21352 13128 21516
rect 13580 21451 13640 21516
rect 13364 21445 13852 21451
rect 13364 21411 13376 21445
rect 13840 21411 13852 21445
rect 13364 21405 13852 21411
rect 13068 21302 13082 21352
rect 13076 20776 13082 21302
rect 13116 21302 13128 21352
rect 14088 21352 14148 21516
rect 14382 21445 14870 21451
rect 14382 21411 14394 21445
rect 14858 21411 14870 21445
rect 14382 21405 14870 21411
rect 13116 20776 13122 21302
rect 14088 21300 14100 21352
rect 13076 20764 13122 20776
rect 14094 20776 14100 21300
rect 14134 21300 14148 21352
rect 15104 21352 15164 24832
rect 17112 24460 17172 27016
rect 17242 24606 17302 27220
rect 18400 27016 18406 27076
rect 18466 27016 18472 27076
rect 17682 26959 18170 26965
rect 17682 26925 17694 26959
rect 18158 26925 18170 26959
rect 17682 26919 18170 26925
rect 17394 26866 17440 26878
rect 17394 26326 17400 26866
rect 17388 26290 17400 26326
rect 17434 26326 17440 26866
rect 18406 26866 18466 27016
rect 18910 26965 18970 27327
rect 18700 26959 19188 26965
rect 18700 26925 18712 26959
rect 19176 26925 19188 26959
rect 18700 26919 19188 26925
rect 18910 26916 18970 26919
rect 18406 26828 18418 26866
rect 17434 26290 17448 26326
rect 18412 26320 18418 26828
rect 17388 26140 17448 26290
rect 18406 26290 18418 26320
rect 18452 26828 18466 26866
rect 19426 26866 19486 27426
rect 20442 27426 20454 27454
rect 20488 27454 20494 28002
rect 21460 28002 21520 28152
rect 21964 28101 22024 28604
rect 21754 28095 22242 28101
rect 21754 28061 21766 28095
rect 22230 28061 22242 28095
rect 21754 28055 22242 28061
rect 21460 27978 21472 28002
rect 21466 27484 21472 27978
rect 20488 27426 20502 27454
rect 19718 27367 20206 27373
rect 19718 27333 19730 27367
rect 20194 27333 20206 27367
rect 19718 27327 20206 27333
rect 20442 27176 20502 27426
rect 21450 27426 21472 27484
rect 21506 27978 21520 28002
rect 22472 28002 22532 28604
rect 22984 28101 23044 28604
rect 23498 28214 23558 28604
rect 23996 28398 24002 28458
rect 24062 28398 24068 28458
rect 25014 28398 25020 28458
rect 25080 28398 25086 28458
rect 23492 28154 23498 28214
rect 23558 28154 23564 28214
rect 22772 28095 23260 28101
rect 22772 28061 22784 28095
rect 23248 28061 23260 28095
rect 22772 28055 23260 28061
rect 21506 27484 21512 27978
rect 22472 27932 22490 28002
rect 21506 27426 21514 27484
rect 20736 27367 21224 27373
rect 20736 27333 20748 27367
rect 21212 27333 21224 27367
rect 20736 27327 21224 27333
rect 20436 27116 20442 27176
rect 20502 27116 20508 27176
rect 19718 26959 20206 26965
rect 19718 26925 19730 26959
rect 20194 26925 20206 26959
rect 19718 26919 20206 26925
rect 20736 26959 21224 26965
rect 20736 26925 20748 26959
rect 21212 26925 21224 26959
rect 20736 26919 21224 26925
rect 18452 26320 18458 26828
rect 19426 26826 19436 26866
rect 18452 26290 18466 26320
rect 19430 26316 19436 26826
rect 17682 26231 18170 26237
rect 17682 26197 17694 26231
rect 18158 26197 18170 26231
rect 17682 26191 18170 26197
rect 17900 26140 17960 26191
rect 18406 26140 18466 26290
rect 19422 26290 19436 26316
rect 19470 26826 19486 26866
rect 20448 26866 20494 26878
rect 19470 26316 19476 26826
rect 19470 26290 19482 26316
rect 20448 26310 20454 26866
rect 18892 26237 18952 26244
rect 18700 26231 19188 26237
rect 18700 26197 18712 26231
rect 19176 26197 19188 26231
rect 18700 26191 19188 26197
rect 17388 26080 18466 26140
rect 18400 25936 18460 25938
rect 17390 25876 18460 25936
rect 17390 25730 17450 25876
rect 17900 25829 17960 25876
rect 17682 25823 18170 25829
rect 17682 25789 17694 25823
rect 18158 25789 18170 25823
rect 17682 25783 18170 25789
rect 17390 25698 17400 25730
rect 17394 25154 17400 25698
rect 17434 25698 17450 25730
rect 18400 25730 18460 25876
rect 18892 25926 18952 26191
rect 18892 25829 18952 25866
rect 19422 26144 19482 26290
rect 20440 26290 20454 26310
rect 20488 26310 20494 26866
rect 21450 26866 21514 27426
rect 22484 27426 22490 27932
rect 22524 27932 22532 28002
rect 23498 28002 23558 28154
rect 24002 28101 24062 28398
rect 25020 28101 25080 28398
rect 25530 28214 25590 28604
rect 26038 28398 26044 28458
rect 26104 28398 26110 28458
rect 27050 28398 27056 28458
rect 27116 28398 27122 28458
rect 25522 28154 25528 28214
rect 25588 28154 25594 28214
rect 23790 28095 24278 28101
rect 23790 28061 23802 28095
rect 24266 28061 24278 28095
rect 23790 28055 24278 28061
rect 24808 28095 25296 28101
rect 24808 28061 24820 28095
rect 25284 28061 25296 28095
rect 24808 28055 25296 28061
rect 23498 27962 23508 28002
rect 22524 27426 22530 27932
rect 23502 27480 23508 27962
rect 22484 27414 22530 27426
rect 23486 27426 23508 27480
rect 23542 27962 23558 28002
rect 24520 28002 24566 28014
rect 23542 27480 23548 27962
rect 23542 27426 23550 27480
rect 24520 27466 24526 28002
rect 21754 27367 22242 27373
rect 21754 27333 21766 27367
rect 22230 27333 22242 27367
rect 21754 27327 22242 27333
rect 22772 27367 23260 27373
rect 22772 27333 22784 27367
rect 23248 27333 23260 27367
rect 22772 27327 23260 27333
rect 22472 27116 22478 27176
rect 22538 27116 22544 27176
rect 21754 26959 22242 26965
rect 21754 26925 21766 26959
rect 22230 26925 22242 26959
rect 21754 26919 22242 26925
rect 21450 26836 21472 26866
rect 21466 26318 21472 26836
rect 20488 26290 20500 26310
rect 19920 26237 19980 26238
rect 19718 26231 20206 26237
rect 19718 26197 19730 26231
rect 20194 26197 20206 26231
rect 19718 26191 20206 26197
rect 19920 26144 19980 26191
rect 20440 26144 20500 26290
rect 21458 26290 21472 26318
rect 21506 26836 21514 26866
rect 22478 26866 22538 27116
rect 22772 26959 23260 26965
rect 22772 26925 22784 26959
rect 23248 26925 23260 26959
rect 22772 26919 23260 26925
rect 21506 26318 21512 26836
rect 22478 26828 22490 26866
rect 22484 26326 22490 26828
rect 21506 26316 21518 26318
rect 21506 26290 21522 26316
rect 20948 26237 21008 26242
rect 20736 26231 21224 26237
rect 20736 26197 20748 26231
rect 21212 26197 21224 26231
rect 20736 26191 21224 26197
rect 20948 26144 21008 26191
rect 19422 26142 21008 26144
rect 21458 26142 21522 26290
rect 22476 26290 22490 26326
rect 22524 26828 22538 26866
rect 23486 26866 23550 27426
rect 24516 27426 24526 27466
rect 24560 27466 24566 28002
rect 25530 28002 25590 28154
rect 26044 28101 26104 28398
rect 27056 28101 27116 28398
rect 27570 28216 27630 28604
rect 27564 28156 27570 28216
rect 27630 28156 27636 28216
rect 25826 28095 26314 28101
rect 25826 28061 25838 28095
rect 26302 28061 26314 28095
rect 25826 28055 26314 28061
rect 26844 28095 27332 28101
rect 26844 28061 26856 28095
rect 27320 28061 27332 28095
rect 26844 28055 27332 28061
rect 25530 27962 25544 28002
rect 25538 27482 25544 27962
rect 24560 27426 24576 27466
rect 24004 27373 24064 27376
rect 23790 27367 24278 27373
rect 23790 27333 23802 27367
rect 24266 27333 24278 27367
rect 23790 27327 24278 27333
rect 24004 26965 24064 27327
rect 24516 27280 24576 27426
rect 25528 27426 25544 27482
rect 25578 27962 25590 28002
rect 26556 28002 26602 28014
rect 25578 27482 25584 27962
rect 25578 27426 25592 27482
rect 26556 27464 26562 28002
rect 25022 27373 25082 27382
rect 24808 27367 25296 27373
rect 24808 27333 24820 27367
rect 25284 27333 25296 27367
rect 24808 27327 25296 27333
rect 24510 27220 24516 27280
rect 24576 27220 24582 27280
rect 24506 27016 24512 27076
rect 24572 27016 24578 27076
rect 23790 26959 24278 26965
rect 23790 26925 23802 26959
rect 24266 26925 24278 26959
rect 23790 26919 24278 26925
rect 24004 26918 24064 26919
rect 23486 26832 23508 26866
rect 22524 26326 22530 26828
rect 23502 26326 23508 26832
rect 22524 26290 22540 26326
rect 21754 26231 22242 26237
rect 21754 26197 21766 26231
rect 22230 26197 22242 26231
rect 21754 26191 22242 26197
rect 19422 26084 20948 26142
rect 18700 25823 19188 25829
rect 18700 25789 18712 25823
rect 19176 25789 19188 25823
rect 18700 25783 19188 25789
rect 18400 25698 18418 25730
rect 17434 25154 17440 25698
rect 18412 25196 18418 25698
rect 17394 25142 17440 25154
rect 18400 25154 18418 25196
rect 18452 25698 18460 25730
rect 19422 25730 19482 26084
rect 21452 26082 21458 26142
rect 21518 26082 21524 26142
rect 20948 26076 21008 26082
rect 20434 25980 20440 26044
rect 20504 25980 20510 26044
rect 19924 25866 19930 25926
rect 19990 25866 19996 25926
rect 20440 25886 20504 25980
rect 19930 25829 19990 25866
rect 19718 25823 20206 25829
rect 19718 25789 19730 25823
rect 20194 25789 20206 25823
rect 19718 25783 20206 25789
rect 18452 25196 18458 25698
rect 19422 25678 19436 25730
rect 18452 25154 18464 25196
rect 19430 25190 19436 25678
rect 17682 25095 18170 25101
rect 17682 25061 17694 25095
rect 18158 25061 18170 25095
rect 17682 25055 18170 25061
rect 18400 24946 18464 25154
rect 19422 25154 19436 25190
rect 19470 25678 19482 25730
rect 20440 25730 20506 25886
rect 20936 25866 20942 25926
rect 21002 25866 21008 25926
rect 20942 25829 21002 25866
rect 20736 25823 21224 25829
rect 20736 25789 20748 25823
rect 21212 25789 21224 25823
rect 20736 25783 21224 25789
rect 20942 25782 21002 25783
rect 20440 25680 20454 25730
rect 19470 25190 19476 25678
rect 19470 25154 19482 25190
rect 20448 25178 20454 25680
rect 18700 25095 19188 25101
rect 18700 25061 18712 25095
rect 19176 25061 19188 25095
rect 18700 25055 19188 25061
rect 17956 24886 18464 24946
rect 17236 24546 17242 24606
rect 17302 24546 17308 24606
rect 17112 24400 17532 24460
rect 17472 21588 17532 24400
rect 17592 22138 17598 22198
rect 17658 22138 17664 22198
rect 16122 21520 17332 21580
rect 17466 21528 17472 21588
rect 17532 21528 17538 21588
rect 15400 21445 15888 21451
rect 15400 21411 15412 21445
rect 15876 21411 15888 21445
rect 15400 21405 15888 21411
rect 14134 20776 14140 21300
rect 14094 20764 14140 20776
rect 15104 20776 15118 21352
rect 15152 20776 15164 21352
rect 16122 21352 16182 21520
rect 16634 21451 16694 21520
rect 16418 21445 16906 21451
rect 16418 21411 16430 21445
rect 16894 21411 16906 21445
rect 16418 21405 16906 21411
rect 16122 21304 16136 21352
rect 13364 20717 13852 20723
rect 13364 20683 13376 20717
rect 13840 20683 13852 20717
rect 13364 20677 13852 20683
rect 14382 20717 14870 20723
rect 14382 20683 14394 20717
rect 14858 20683 14870 20717
rect 14382 20677 14870 20683
rect 14588 20634 14648 20677
rect 14582 20574 14588 20634
rect 14648 20574 14654 20634
rect 14690 20462 14696 20522
rect 14756 20462 14762 20522
rect 14696 20419 14756 20462
rect 13364 20413 13852 20419
rect 13364 20379 13376 20413
rect 13840 20379 13852 20413
rect 13364 20373 13852 20379
rect 14382 20413 14870 20419
rect 14382 20379 14394 20413
rect 14858 20379 14870 20413
rect 14382 20373 14870 20379
rect 13076 20320 13122 20332
rect 13076 19802 13082 20320
rect 13066 19744 13082 19802
rect 13116 19802 13122 20320
rect 14094 20320 14140 20332
rect 13116 19744 13126 19802
rect 14094 19794 14100 20320
rect 12920 19540 12926 19600
rect 12986 19540 12992 19600
rect 12800 18512 12860 18518
rect 12926 18512 12986 19540
rect 13066 19490 13126 19744
rect 14086 19744 14100 19794
rect 14134 19794 14140 20320
rect 15104 20320 15164 20776
rect 16130 20776 16136 21304
rect 16170 21304 16182 21352
rect 17140 21352 17200 21520
rect 17140 21306 17154 21352
rect 16170 20776 16176 21304
rect 16130 20764 16176 20776
rect 17148 20776 17154 21306
rect 17188 21306 17200 21352
rect 17188 20776 17194 21306
rect 17148 20764 17194 20776
rect 15400 20717 15888 20723
rect 15400 20683 15412 20717
rect 15876 20683 15888 20717
rect 15400 20677 15888 20683
rect 16418 20717 16906 20723
rect 16418 20683 16430 20717
rect 16894 20683 16906 20717
rect 16418 20677 16906 20683
rect 15480 20522 15540 20677
rect 15604 20574 15610 20634
rect 15670 20574 15676 20634
rect 15474 20462 15480 20522
rect 15540 20462 15546 20522
rect 15610 20419 15670 20574
rect 15400 20413 15888 20419
rect 15400 20379 15412 20413
rect 15876 20379 15888 20413
rect 15400 20373 15888 20379
rect 16418 20413 16906 20419
rect 16418 20379 16430 20413
rect 16894 20379 16906 20413
rect 16418 20373 16906 20379
rect 14134 19744 14146 19794
rect 13364 19685 13852 19691
rect 13364 19651 13376 19685
rect 13840 19651 13852 19685
rect 13364 19645 13852 19651
rect 13568 19490 13628 19645
rect 14086 19490 14146 19744
rect 15104 19744 15118 20320
rect 15152 19744 15164 20320
rect 16130 20320 16176 20332
rect 16130 19830 16136 20320
rect 14382 19685 14870 19691
rect 14382 19651 14394 19685
rect 14858 19651 14870 19685
rect 14382 19645 14870 19651
rect 13066 19430 14086 19490
rect 14146 19430 14152 19490
rect 13066 19288 13126 19430
rect 13568 19387 13628 19430
rect 13364 19381 13852 19387
rect 13364 19347 13376 19381
rect 13840 19347 13852 19381
rect 13364 19341 13852 19347
rect 13066 19228 13082 19288
rect 13076 18712 13082 19228
rect 13116 19228 13126 19288
rect 14086 19288 14146 19430
rect 14596 19387 14656 19645
rect 14382 19381 14870 19387
rect 14382 19347 14394 19381
rect 14858 19347 14870 19381
rect 14382 19341 14870 19347
rect 13116 18712 13122 19228
rect 14086 19224 14100 19288
rect 13076 18700 13122 18712
rect 14094 18712 14100 19224
rect 14134 19224 14146 19288
rect 15104 19288 15164 19744
rect 16120 19744 16136 19830
rect 16170 19830 16176 20320
rect 17148 20320 17194 20332
rect 16170 19744 16180 19830
rect 17148 19790 17154 20320
rect 15400 19685 15888 19691
rect 15400 19651 15412 19685
rect 15876 19651 15888 19685
rect 15400 19645 15888 19651
rect 15614 19387 15674 19645
rect 16120 19600 16180 19744
rect 17140 19744 17154 19790
rect 17188 19790 17194 20320
rect 17188 19744 17200 19790
rect 16418 19685 16906 19691
rect 16418 19651 16430 19685
rect 16894 19651 16906 19685
rect 16418 19645 16906 19651
rect 16634 19600 16694 19645
rect 17140 19600 17200 19744
rect 16114 19540 16120 19600
rect 16180 19540 17200 19600
rect 15400 19381 15888 19387
rect 15400 19347 15412 19381
rect 15876 19347 15888 19381
rect 15400 19341 15888 19347
rect 14134 18712 14140 19224
rect 14094 18700 14140 18712
rect 15104 18712 15118 19288
rect 15152 18712 15164 19288
rect 16120 19288 16180 19540
rect 16634 19387 16694 19540
rect 16418 19381 16906 19387
rect 16418 19347 16430 19381
rect 16894 19347 16906 19381
rect 16418 19341 16906 19347
rect 16120 19232 16136 19288
rect 13364 18653 13852 18659
rect 13364 18619 13376 18653
rect 13840 18619 13852 18653
rect 13364 18613 13852 18619
rect 14382 18653 14870 18659
rect 14382 18619 14394 18653
rect 14858 18619 14870 18653
rect 14382 18613 14870 18619
rect 14602 18566 14662 18613
rect 12860 18452 14150 18512
rect 14596 18506 14602 18566
rect 14662 18506 14668 18566
rect 12800 18446 12860 18452
rect 13064 18256 13124 18452
rect 13572 18355 13632 18452
rect 13364 18349 13852 18355
rect 13364 18315 13376 18349
rect 13840 18315 13852 18349
rect 13364 18309 13852 18315
rect 13064 18204 13082 18256
rect 13076 17680 13082 18204
rect 13116 18204 13124 18256
rect 14090 18256 14150 18452
rect 14702 18406 14708 18466
rect 14768 18406 14774 18466
rect 14708 18355 14768 18406
rect 14382 18349 14870 18355
rect 14382 18315 14394 18349
rect 14858 18315 14870 18349
rect 14382 18309 14870 18315
rect 14090 18208 14100 18256
rect 13116 17680 13122 18204
rect 13076 17668 13122 17680
rect 14094 17680 14100 18208
rect 14134 18208 14150 18256
rect 15104 18256 15164 18712
rect 16130 18712 16136 19232
rect 16170 19232 16180 19288
rect 17140 19288 17200 19540
rect 17272 19490 17332 21520
rect 17266 19430 17272 19490
rect 17332 19430 17338 19490
rect 17140 19252 17154 19288
rect 16170 18712 16176 19232
rect 16130 18700 16176 18712
rect 17148 18712 17154 19252
rect 17188 19252 17200 19288
rect 17188 18712 17194 19252
rect 17148 18700 17194 18712
rect 15400 18653 15888 18659
rect 15400 18619 15412 18653
rect 15876 18619 15888 18653
rect 15400 18613 15888 18619
rect 16418 18653 16906 18659
rect 16418 18619 16430 18653
rect 16894 18619 16906 18653
rect 16418 18613 16906 18619
rect 15494 18466 15554 18613
rect 15606 18506 15612 18566
rect 15672 18506 15678 18566
rect 17272 18512 17332 19430
rect 17458 19302 17464 19362
rect 17524 19302 17530 19362
rect 15488 18406 15494 18466
rect 15554 18406 15560 18466
rect 15612 18355 15672 18506
rect 16120 18452 17332 18512
rect 15400 18349 15888 18355
rect 15400 18315 15412 18349
rect 15876 18315 15888 18349
rect 15400 18309 15888 18315
rect 14134 17680 14140 18208
rect 15104 18182 15118 18256
rect 14094 17668 14140 17680
rect 15112 17680 15118 18182
rect 15152 18182 15164 18256
rect 16120 18256 16180 18452
rect 16622 18355 16682 18452
rect 16418 18349 16906 18355
rect 16418 18315 16430 18349
rect 16894 18315 16906 18349
rect 16418 18309 16906 18315
rect 16120 18226 16136 18256
rect 15152 17680 15158 18182
rect 16130 17762 16136 18226
rect 15112 17668 15158 17680
rect 16122 17680 16136 17762
rect 16170 18226 16180 18256
rect 17140 18256 17200 18452
rect 16170 17762 16176 18226
rect 17140 18188 17154 18256
rect 16170 17680 16182 17762
rect 15600 17627 15660 17631
rect 13364 17621 13852 17627
rect 13364 17587 13376 17621
rect 13840 17587 13852 17621
rect 13364 17581 13852 17587
rect 14382 17621 14870 17627
rect 14382 17587 14394 17621
rect 14858 17587 14870 17621
rect 14382 17581 14870 17587
rect 15400 17621 15888 17627
rect 15400 17587 15412 17621
rect 15876 17587 15888 17621
rect 15400 17581 15888 17587
rect 12314 17456 12374 17462
rect 14594 17456 14654 17581
rect 12374 17396 14654 17456
rect 12314 17390 12374 17396
rect 12454 17280 12514 17286
rect 15600 17280 15660 17581
rect 12514 17220 15660 17280
rect 12454 17214 12514 17220
rect 13354 17106 13414 17112
rect 16122 17106 16182 17680
rect 17148 17680 17154 18188
rect 17188 18188 17200 18256
rect 17188 17680 17194 18188
rect 17148 17668 17194 17680
rect 16418 17621 16906 17627
rect 16418 17587 16430 17621
rect 16894 17587 16906 17621
rect 16418 17581 16906 17587
rect 13414 17046 16182 17106
rect 13354 17040 13414 17046
rect 12194 16956 12254 16962
rect 17464 16956 17524 19302
rect 17598 18210 17658 22138
rect 17708 21528 17714 21588
rect 17774 21528 17780 21588
rect 17714 19466 17774 21528
rect 17956 20624 18016 24886
rect 18400 24756 18464 24886
rect 18394 24692 18400 24756
rect 18464 24692 18470 24756
rect 18224 24606 18284 24612
rect 18224 21670 18284 24546
rect 18902 24500 18962 25055
rect 19422 25004 19482 25154
rect 20438 25154 20454 25178
rect 20488 25684 20506 25730
rect 21458 25730 21522 26082
rect 21952 25934 22012 26191
rect 22476 26044 22540 26290
rect 23492 26290 23508 26326
rect 23542 26832 23550 26866
rect 24512 26866 24572 27016
rect 25022 26965 25082 27327
rect 24808 26959 25296 26965
rect 24808 26925 24820 26959
rect 25284 26925 25296 26959
rect 24808 26919 25296 26925
rect 24512 26840 24526 26866
rect 23542 26326 23548 26832
rect 23542 26324 23552 26326
rect 23542 26290 23556 26324
rect 22772 26231 23260 26237
rect 22772 26197 22784 26231
rect 23248 26197 23260 26231
rect 22772 26191 23260 26197
rect 22310 25980 22316 26044
rect 22380 25980 22540 26044
rect 22976 25934 23036 26191
rect 23492 26142 23556 26290
rect 24520 26290 24526 26840
rect 24560 26840 24572 26866
rect 25528 26866 25592 27426
rect 26550 27426 26562 27464
rect 26596 27464 26602 28002
rect 27570 28002 27630 28156
rect 28060 28101 28120 28604
rect 28580 28216 28640 28604
rect 28574 28156 28580 28216
rect 28640 28156 28646 28216
rect 27862 28095 28350 28101
rect 27862 28061 27874 28095
rect 28338 28061 28350 28095
rect 27862 28055 28350 28061
rect 27570 27964 27580 28002
rect 27574 27466 27580 27964
rect 26596 27426 26610 27464
rect 26038 27373 26098 27379
rect 25826 27367 26314 27373
rect 25826 27333 25838 27367
rect 26302 27333 26314 27367
rect 25826 27327 26314 27333
rect 26038 26965 26098 27327
rect 26550 27280 26610 27426
rect 27566 27426 27580 27466
rect 27614 27964 27630 28002
rect 28580 28002 28640 28156
rect 29088 28101 29148 28604
rect 29602 28216 29662 28604
rect 30108 28398 30114 28458
rect 30174 28398 30180 28458
rect 31120 28398 31126 28458
rect 31186 28398 31192 28458
rect 29596 28156 29602 28216
rect 29662 28156 29668 28216
rect 28880 28095 29368 28101
rect 28880 28061 28892 28095
rect 29356 28061 29368 28095
rect 28880 28055 29368 28061
rect 29088 28052 29148 28055
rect 27614 27466 27620 27964
rect 28580 27932 28598 28002
rect 27614 27426 27630 27466
rect 27050 27373 27110 27379
rect 26844 27367 27332 27373
rect 26844 27333 26856 27367
rect 27320 27333 27332 27367
rect 26844 27327 27332 27333
rect 26544 27220 26550 27280
rect 26610 27220 26616 27280
rect 27050 27076 27110 27327
rect 26542 27016 26548 27076
rect 26608 27016 26614 27076
rect 27044 27016 27050 27076
rect 27110 27016 27116 27076
rect 25826 26959 26314 26965
rect 25826 26925 25838 26959
rect 26302 26925 26314 26959
rect 25826 26919 26314 26925
rect 26038 26916 26098 26919
rect 24560 26290 24566 26840
rect 25528 26834 25544 26866
rect 25538 26338 25544 26834
rect 24520 26278 24566 26290
rect 25530 26290 25544 26338
rect 25578 26834 25592 26866
rect 26548 26866 26608 27016
rect 27050 26965 27110 27016
rect 26844 26959 27332 26965
rect 26844 26925 26856 26959
rect 27320 26925 27332 26959
rect 26844 26919 27332 26925
rect 27050 26916 27110 26919
rect 26548 26834 26562 26866
rect 25578 26338 25584 26834
rect 25578 26336 25590 26338
rect 25578 26290 25594 26336
rect 26556 26320 26562 26834
rect 24004 26237 24064 26244
rect 23790 26231 24278 26237
rect 23790 26197 23802 26231
rect 24266 26197 24278 26231
rect 23790 26191 24278 26197
rect 24808 26231 25296 26237
rect 24808 26197 24820 26231
rect 25284 26197 25296 26231
rect 24808 26191 25296 26197
rect 23486 26082 23492 26142
rect 23552 26082 23558 26142
rect 21946 25874 21952 25934
rect 22012 25874 22018 25934
rect 22970 25874 22976 25934
rect 23036 25874 23042 25934
rect 21754 25823 22242 25829
rect 21754 25789 21766 25823
rect 22230 25789 22242 25823
rect 21754 25783 22242 25789
rect 22772 25823 23260 25829
rect 22772 25789 22784 25823
rect 23248 25789 23260 25823
rect 22772 25783 23260 25789
rect 20488 25680 20504 25684
rect 21458 25682 21472 25730
rect 20488 25178 20494 25680
rect 21466 25180 21472 25682
rect 20488 25154 20502 25178
rect 19718 25095 20206 25101
rect 19718 25061 19730 25095
rect 20194 25061 20206 25095
rect 19718 25055 20206 25061
rect 19416 24944 19422 25004
rect 19482 24944 19488 25004
rect 19944 24500 20004 25055
rect 20438 24894 20502 25154
rect 21458 25154 21472 25180
rect 21506 25682 21522 25730
rect 22484 25730 22530 25742
rect 21506 25180 21512 25682
rect 22484 25210 22490 25730
rect 21506 25178 21518 25180
rect 21506 25154 21522 25178
rect 20736 25095 21224 25101
rect 20736 25061 20748 25095
rect 21212 25061 21224 25095
rect 20736 25055 21224 25061
rect 20432 24830 20438 24894
rect 20502 24830 20508 24894
rect 20944 24500 21004 25055
rect 21458 25004 21522 25154
rect 22478 25154 22490 25210
rect 22524 25210 22530 25730
rect 23492 25730 23556 26082
rect 24004 25934 24064 26191
rect 23998 25874 24004 25934
rect 24064 25874 24070 25934
rect 24004 25829 24064 25874
rect 25032 25829 25092 26191
rect 25530 26140 25594 26290
rect 26550 26290 26562 26320
rect 26596 26834 26608 26866
rect 27566 26866 27630 27426
rect 28592 27426 28598 27932
rect 28632 27932 28640 28002
rect 29602 28002 29662 28156
rect 30114 28101 30174 28398
rect 31126 28101 31186 28398
rect 31638 28216 31698 28604
rect 32138 28398 32144 28458
rect 32204 28398 32210 28458
rect 31632 28156 31638 28216
rect 31698 28156 31704 28216
rect 29898 28095 30386 28101
rect 29898 28061 29910 28095
rect 30374 28061 30386 28095
rect 29898 28055 30386 28061
rect 30916 28095 31404 28101
rect 30916 28061 30928 28095
rect 31392 28061 31404 28095
rect 30916 28055 31404 28061
rect 29602 27974 29616 28002
rect 28632 27426 28638 27932
rect 29610 27474 29616 27974
rect 28592 27414 28638 27426
rect 29602 27426 29616 27474
rect 29650 27974 29662 28002
rect 30628 28002 30674 28014
rect 29650 27474 29656 27974
rect 29650 27426 29662 27474
rect 30628 27458 30634 28002
rect 27862 27367 28350 27373
rect 27862 27333 27874 27367
rect 28338 27333 28350 27367
rect 27862 27327 28350 27333
rect 28880 27367 29368 27373
rect 28880 27333 28892 27367
rect 29356 27333 29368 27367
rect 28880 27327 29368 27333
rect 28578 27116 28584 27176
rect 28644 27116 28650 27176
rect 28064 27016 28070 27076
rect 28130 27016 28136 27076
rect 28070 26965 28130 27016
rect 27862 26959 28350 26965
rect 27862 26925 27874 26959
rect 28338 26925 28350 26959
rect 27862 26919 28350 26925
rect 26596 26320 26602 26834
rect 27566 26818 27580 26866
rect 27574 26334 27580 26818
rect 26596 26290 26610 26320
rect 26050 26237 26110 26249
rect 25826 26231 26314 26237
rect 25826 26197 25838 26231
rect 26302 26197 26314 26231
rect 25826 26191 26314 26197
rect 25524 26080 25530 26140
rect 25590 26080 25596 26140
rect 23790 25823 24278 25829
rect 23790 25789 23802 25823
rect 24266 25789 24278 25823
rect 23790 25783 24278 25789
rect 24808 25823 25296 25829
rect 24808 25789 24820 25823
rect 25284 25789 25296 25823
rect 24808 25783 25296 25789
rect 25032 25776 25092 25783
rect 23492 25670 23508 25730
rect 22524 25154 22538 25210
rect 23502 25188 23508 25670
rect 21980 25101 22040 25104
rect 21754 25095 22242 25101
rect 21754 25061 21766 25095
rect 22230 25061 22242 25095
rect 21754 25055 22242 25061
rect 21980 25004 22040 25055
rect 22478 25004 22538 25154
rect 23492 25154 23508 25188
rect 23542 25670 23556 25730
rect 24520 25730 24566 25742
rect 23542 25188 23548 25670
rect 23542 25186 23552 25188
rect 24520 25186 24526 25730
rect 23542 25154 23556 25186
rect 22772 25095 23260 25101
rect 22772 25061 22784 25095
rect 23248 25061 23260 25095
rect 22772 25055 23260 25061
rect 21452 24944 21458 25004
rect 21518 24944 21524 25004
rect 21974 24944 21980 25004
rect 22040 24944 22046 25004
rect 22472 24944 22478 25004
rect 22538 24944 22544 25004
rect 22952 25000 23012 25055
rect 23492 25008 23556 25154
rect 24510 25154 24526 25186
rect 24560 25186 24566 25730
rect 25530 25730 25594 26080
rect 26050 25829 26110 26191
rect 26550 26042 26610 26290
rect 27566 26290 27580 26334
rect 27614 26818 27630 26866
rect 28584 26866 28644 27116
rect 29090 27016 29096 27076
rect 29156 27016 29162 27076
rect 29602 27072 29662 27426
rect 30618 27426 30634 27458
rect 30668 27458 30674 28002
rect 31638 28002 31698 28156
rect 32144 28101 32204 28398
rect 32658 28164 33738 28224
rect 31934 28095 32422 28101
rect 31934 28061 31946 28095
rect 32410 28061 32422 28095
rect 31934 28055 32422 28061
rect 31638 27970 31652 28002
rect 31646 27464 31652 27970
rect 30668 27426 30678 27458
rect 29898 27367 30386 27373
rect 29898 27333 29910 27367
rect 30374 27333 30386 27367
rect 29898 27327 30386 27333
rect 30618 27176 30678 27426
rect 31642 27426 31652 27464
rect 31686 27970 31698 28002
rect 32658 28002 32718 28164
rect 33160 28101 33220 28164
rect 32952 28095 33440 28101
rect 32952 28061 32964 28095
rect 33428 28061 33440 28095
rect 32952 28055 33440 28061
rect 32658 27972 32670 28002
rect 31686 27464 31692 27970
rect 32664 27466 32670 27972
rect 31686 27426 31702 27464
rect 30916 27367 31404 27373
rect 30916 27333 30928 27367
rect 31392 27333 31404 27367
rect 30916 27327 31404 27333
rect 30612 27116 30618 27176
rect 30678 27116 30684 27176
rect 31642 27078 31702 27426
rect 32658 27426 32670 27466
rect 32704 27972 32718 28002
rect 33678 28002 33738 28164
rect 32704 27466 32710 27972
rect 33678 27956 33688 28002
rect 32704 27426 32718 27466
rect 32122 27373 32182 27385
rect 31934 27367 32422 27373
rect 31934 27333 31946 27367
rect 32410 27333 32422 27367
rect 31934 27327 32422 27333
rect 31642 27072 31706 27078
rect 29096 26965 29156 27016
rect 29596 27012 29602 27072
rect 29662 27012 29668 27072
rect 30110 27012 30116 27072
rect 30176 27012 30182 27072
rect 30614 27012 30620 27072
rect 30680 27012 30686 27072
rect 31120 27012 31126 27072
rect 31186 27012 31192 27072
rect 31642 27012 31646 27072
rect 28880 26959 29368 26965
rect 28880 26925 28892 26959
rect 29356 26925 29368 26959
rect 28880 26919 29368 26925
rect 28584 26842 28598 26866
rect 27614 26334 27620 26818
rect 27614 26332 27626 26334
rect 27614 26290 27630 26332
rect 27050 26237 27110 26245
rect 26844 26231 27332 26237
rect 26844 26197 26856 26231
rect 27320 26197 27332 26231
rect 26844 26191 27332 26197
rect 26544 25982 26550 26042
rect 26610 25982 26616 26042
rect 27050 25829 27110 26191
rect 27566 26140 27630 26290
rect 28592 26290 28598 26842
rect 28632 26842 28644 26866
rect 29602 26866 29662 27012
rect 30116 26965 30176 27012
rect 29898 26959 30386 26965
rect 29898 26925 29910 26959
rect 30374 26925 30386 26959
rect 29898 26919 30386 26925
rect 28632 26290 28638 26842
rect 29602 26822 29616 26866
rect 29610 26326 29616 26822
rect 28592 26278 28638 26290
rect 29602 26290 29616 26326
rect 29650 26822 29662 26866
rect 30620 26866 30680 27012
rect 31126 26965 31186 27012
rect 31642 27006 31706 27012
rect 30916 26959 31404 26965
rect 30916 26925 30928 26959
rect 31392 26925 31404 26959
rect 30916 26919 31404 26925
rect 30620 26838 30634 26866
rect 29650 26326 29656 26822
rect 30628 26360 30634 26838
rect 29650 26290 29662 26326
rect 27862 26231 28350 26237
rect 27862 26197 27874 26231
rect 28338 26197 28350 26231
rect 27862 26191 28350 26197
rect 28880 26231 29368 26237
rect 28880 26197 28892 26231
rect 29356 26197 29368 26231
rect 28880 26191 29368 26197
rect 29602 26140 29662 26290
rect 30618 26290 30634 26360
rect 30668 26838 30680 26866
rect 31642 26866 31702 27006
rect 32122 26965 32182 27327
rect 32658 27280 32718 27426
rect 33682 27426 33688 27956
rect 33722 27956 33738 28002
rect 33722 27426 33728 27956
rect 33682 27414 33728 27426
rect 32952 27367 33440 27373
rect 32952 27333 32964 27367
rect 33428 27333 33440 27367
rect 32952 27327 33440 27333
rect 32652 27220 32658 27280
rect 32718 27220 32724 27280
rect 33902 27220 33908 27280
rect 33968 27220 33974 27280
rect 32662 27004 33732 27064
rect 31934 26959 32422 26965
rect 31934 26925 31946 26959
rect 32410 26925 32422 26959
rect 31934 26919 32422 26925
rect 30668 26360 30674 26838
rect 31642 26830 31652 26866
rect 30668 26290 30678 26360
rect 31646 26322 31652 26830
rect 29898 26231 30386 26237
rect 29898 26197 29910 26231
rect 30374 26197 30386 26231
rect 29898 26191 30386 26197
rect 30104 26140 30164 26191
rect 27560 26080 27566 26140
rect 27626 26080 27632 26140
rect 28060 26080 28066 26140
rect 28126 26080 28132 26140
rect 28574 26080 28580 26140
rect 28640 26080 28646 26140
rect 29098 26080 29104 26140
rect 29164 26080 29170 26140
rect 29596 26080 29602 26140
rect 29662 26080 29668 26140
rect 30098 26080 30104 26140
rect 30164 26080 30170 26140
rect 30618 26138 30678 26290
rect 31636 26290 31652 26322
rect 31686 26830 31702 26866
rect 32662 26866 32722 27004
rect 33168 26965 33228 27004
rect 32952 26959 33440 26965
rect 32952 26925 32964 26959
rect 33428 26925 33440 26959
rect 32952 26919 33440 26925
rect 32662 26838 32670 26866
rect 31686 26322 31692 26830
rect 31686 26320 31696 26322
rect 32664 26320 32670 26838
rect 31686 26290 31700 26320
rect 31126 26237 31186 26244
rect 30916 26231 31404 26237
rect 30916 26197 30928 26231
rect 31392 26197 31404 26231
rect 30916 26191 31404 26197
rect 31126 26138 31186 26191
rect 31636 26138 31700 26290
rect 32658 26290 32670 26320
rect 32704 26838 32722 26866
rect 33672 26866 33732 27004
rect 32704 26320 32710 26838
rect 33672 26832 33688 26866
rect 32704 26290 32718 26320
rect 32122 26237 32182 26243
rect 31934 26231 32422 26237
rect 31934 26197 31946 26231
rect 32410 26197 32422 26231
rect 31934 26191 32422 26197
rect 25826 25823 26314 25829
rect 25826 25789 25838 25823
rect 26302 25789 26314 25823
rect 25826 25783 26314 25789
rect 26844 25823 27332 25829
rect 26844 25789 26856 25823
rect 27320 25789 27332 25823
rect 26844 25783 27332 25789
rect 27050 25782 27110 25783
rect 25530 25690 25544 25730
rect 25538 25214 25544 25690
rect 24560 25154 24574 25186
rect 23790 25095 24278 25101
rect 23790 25061 23802 25095
rect 24266 25061 24278 25095
rect 23790 25055 24278 25061
rect 18334 24440 18340 24500
rect 18400 24440 18406 24500
rect 18896 24440 18902 24500
rect 18962 24440 18968 24500
rect 19938 24440 19944 24500
rect 20004 24440 20010 24500
rect 20938 24440 20944 24500
rect 21004 24440 21010 24500
rect 18340 21858 18400 24440
rect 22952 24402 23012 24940
rect 23460 25004 23556 25008
rect 23460 25002 23492 25004
rect 23552 24944 23558 25004
rect 23946 24944 23952 25004
rect 24012 24944 24018 25004
rect 23460 24402 23520 24942
rect 23952 24402 24012 24944
rect 24106 24500 24166 25055
rect 24510 24752 24574 25154
rect 25528 25154 25544 25214
rect 25578 25690 25594 25730
rect 26556 25730 26602 25742
rect 25578 25214 25584 25690
rect 25578 25154 25588 25214
rect 26556 25190 26562 25730
rect 24808 25095 25296 25101
rect 24808 25061 24820 25095
rect 25284 25061 25296 25095
rect 24808 25055 25296 25061
rect 24510 24682 24574 24688
rect 24996 25006 25056 25012
rect 24100 24440 24106 24500
rect 24166 24440 24172 24500
rect 24996 24402 25056 24946
rect 25116 24500 25176 25055
rect 25528 25004 25588 25154
rect 26546 25154 26562 25190
rect 26596 25190 26602 25730
rect 27566 25730 27630 26080
rect 28066 25829 28126 26080
rect 27862 25823 28350 25829
rect 27862 25789 27874 25823
rect 28338 25789 28350 25823
rect 27862 25783 28350 25789
rect 27566 25678 27580 25730
rect 27574 25196 27580 25678
rect 26596 25154 26610 25190
rect 25826 25095 26314 25101
rect 25826 25061 25838 25095
rect 26302 25061 26314 25095
rect 25826 25055 26314 25061
rect 25522 24944 25528 25004
rect 25588 24944 25594 25004
rect 26058 24500 26118 25055
rect 26546 24610 26610 25154
rect 27566 25154 27580 25196
rect 27614 25678 27630 25730
rect 28580 25730 28640 26080
rect 29104 25829 29164 26080
rect 28880 25823 29368 25829
rect 28880 25789 28892 25823
rect 29356 25789 29368 25823
rect 28880 25783 29368 25789
rect 27614 25196 27620 25678
rect 28580 25676 28598 25730
rect 28592 25600 28598 25676
rect 27614 25194 27626 25196
rect 27614 25154 27630 25194
rect 26844 25095 27332 25101
rect 26844 25061 26856 25095
rect 27320 25061 27332 25095
rect 26844 25055 27332 25061
rect 27040 25006 27100 25012
rect 27566 25006 27630 25154
rect 28584 25154 28598 25600
rect 28632 25676 28640 25730
rect 29602 25730 29662 26080
rect 30612 26078 30618 26138
rect 30678 26078 30684 26138
rect 31120 26078 31126 26138
rect 31186 26078 31192 26138
rect 31630 26078 31636 26138
rect 31696 26078 31702 26138
rect 30102 25866 30108 25926
rect 30168 25866 30174 25926
rect 31114 25866 31120 25926
rect 31180 25866 31186 25926
rect 30108 25829 30168 25866
rect 31120 25829 31180 25866
rect 29898 25823 30386 25829
rect 29898 25789 29910 25823
rect 30374 25789 30386 25823
rect 29898 25783 30386 25789
rect 30916 25823 31404 25829
rect 30916 25789 30928 25823
rect 31392 25789 31404 25823
rect 30916 25783 31404 25789
rect 29602 25676 29616 25730
rect 28632 25600 28638 25676
rect 28632 25154 28644 25600
rect 29610 25184 29616 25676
rect 28062 25101 28122 25110
rect 27862 25095 28350 25101
rect 27862 25061 27874 25095
rect 28338 25061 28350 25095
rect 27862 25055 28350 25061
rect 26540 24546 26546 24610
rect 26610 24546 26616 24610
rect 25110 24440 25116 24500
rect 25176 24440 25182 24500
rect 26052 24440 26058 24500
rect 26118 24440 26124 24500
rect 27040 24402 27100 24946
rect 27534 25002 27630 25006
rect 27534 25000 27566 25002
rect 27626 24942 27632 25002
rect 28062 24996 28122 25055
rect 28584 25006 28644 25154
rect 29602 25154 29616 25184
rect 29650 25676 29662 25730
rect 30628 25730 30674 25742
rect 29650 25184 29656 25676
rect 30628 25188 30634 25730
rect 29650 25182 29662 25184
rect 29650 25154 29666 25182
rect 29062 25101 29122 25104
rect 28880 25095 29368 25101
rect 28880 25061 28892 25095
rect 29356 25061 29368 25095
rect 28880 25055 29368 25061
rect 27534 24402 27594 24940
rect 28062 24402 28122 24936
rect 28550 25000 28644 25006
rect 28610 24998 28644 25000
rect 28550 24938 28584 24940
rect 28550 24932 28644 24938
rect 29062 24996 29122 25055
rect 29602 25000 29666 25154
rect 30618 25154 30634 25188
rect 30668 25188 30674 25730
rect 31636 25730 31700 26078
rect 32122 25926 32182 26191
rect 32658 26042 32718 26290
rect 33682 26290 33688 26832
rect 33722 26832 33732 26866
rect 33722 26290 33728 26832
rect 33682 26278 33728 26290
rect 32952 26231 33440 26237
rect 32952 26197 32964 26231
rect 33428 26197 33440 26231
rect 32952 26191 33440 26197
rect 32652 25982 32658 26042
rect 32718 25982 32724 26042
rect 32660 25928 32720 25930
rect 32116 25866 32122 25926
rect 32182 25866 32188 25926
rect 32660 25868 33732 25928
rect 32122 25829 32182 25866
rect 31934 25823 32422 25829
rect 31934 25789 31946 25823
rect 32410 25789 32422 25823
rect 31934 25783 32422 25789
rect 32122 25780 32182 25783
rect 31636 25684 31652 25730
rect 30668 25154 30682 25188
rect 31646 25184 31652 25684
rect 29898 25095 30386 25101
rect 29898 25061 29910 25095
rect 30374 25061 30386 25095
rect 29898 25055 30386 25061
rect 29596 24940 29602 25000
rect 29662 24940 29668 25000
rect 28550 24402 28610 24932
rect 29062 24402 29122 24936
rect 30618 24894 30682 25154
rect 31636 25154 31652 25184
rect 31686 25684 31700 25730
rect 32660 25730 32720 25868
rect 33164 25829 33224 25868
rect 32952 25823 33440 25829
rect 32952 25789 32964 25823
rect 33428 25789 33440 25823
rect 32952 25783 33440 25789
rect 32660 25704 32670 25730
rect 31686 25184 31692 25684
rect 32664 25242 32670 25704
rect 31686 25182 31696 25184
rect 31686 25154 31700 25182
rect 30916 25095 31404 25101
rect 30916 25061 30928 25095
rect 31392 25061 31404 25095
rect 30916 25055 31404 25061
rect 31636 25000 31700 25154
rect 32652 25154 32670 25242
rect 32704 25704 32720 25730
rect 33672 25730 33732 25868
rect 32704 25242 32710 25704
rect 33672 25680 33688 25730
rect 32704 25154 32712 25242
rect 31934 25095 32422 25101
rect 31934 25061 31946 25095
rect 32410 25061 32422 25095
rect 31934 25055 32422 25061
rect 31630 24940 31636 25000
rect 31696 24940 31702 25000
rect 30612 24830 30618 24894
rect 30682 24830 30688 24894
rect 32652 24606 32712 25154
rect 33682 25154 33688 25680
rect 33722 25680 33732 25730
rect 33722 25154 33728 25680
rect 33682 25142 33728 25154
rect 32952 25095 33440 25101
rect 32952 25061 32964 25095
rect 33428 25061 33440 25095
rect 32952 25055 33440 25061
rect 33908 24762 33968 27220
rect 33904 24756 33968 24762
rect 33904 24686 33968 24692
rect 32646 24546 32652 24606
rect 32712 24546 32718 24606
rect 20616 24342 30856 24402
rect 18448 24238 18454 24298
rect 18514 24238 18520 24298
rect 18454 22324 18514 24238
rect 18876 24185 19364 24191
rect 18876 24151 18888 24185
rect 19352 24151 19364 24185
rect 18876 24145 19364 24151
rect 19894 24185 20382 24191
rect 19894 24151 19906 24185
rect 20370 24151 20382 24185
rect 19894 24145 20382 24151
rect 18588 24092 18634 24104
rect 18588 23546 18594 24092
rect 18580 23516 18594 23546
rect 18628 23546 18634 24092
rect 19606 24092 19652 24104
rect 18628 23516 18640 23546
rect 19606 23540 19612 24092
rect 18580 23364 18640 23516
rect 19598 23516 19612 23540
rect 19646 23540 19652 24092
rect 20616 24092 20676 24342
rect 21626 24238 21632 24298
rect 21692 24238 21698 24298
rect 20912 24185 21400 24191
rect 20912 24151 20924 24185
rect 21388 24151 21400 24185
rect 20912 24145 21400 24151
rect 19646 23516 19658 23540
rect 18876 23457 19364 23463
rect 18876 23423 18888 23457
rect 19352 23423 19364 23457
rect 18876 23417 19364 23423
rect 19092 23364 19152 23417
rect 19598 23364 19658 23516
rect 20616 23516 20630 24092
rect 20664 23516 20676 24092
rect 21632 24092 21692 24238
rect 21930 24185 22418 24191
rect 21930 24151 21942 24185
rect 22406 24151 22418 24185
rect 21930 24145 22418 24151
rect 21632 24028 21648 24092
rect 19894 23457 20382 23463
rect 19894 23423 19906 23457
rect 20370 23423 20382 23457
rect 19894 23417 20382 23423
rect 18580 23362 19658 23364
rect 18580 23304 19598 23362
rect 19592 23302 19598 23304
rect 19658 23302 19664 23362
rect 20102 23254 20162 23417
rect 20096 23194 20102 23254
rect 20162 23194 20168 23254
rect 20102 23159 20162 23194
rect 18876 23153 19364 23159
rect 18876 23119 18888 23153
rect 19352 23119 19364 23153
rect 18876 23113 19364 23119
rect 19894 23153 20382 23159
rect 19894 23119 19906 23153
rect 20370 23119 20382 23153
rect 19894 23113 20382 23119
rect 18588 23060 18634 23072
rect 18588 22540 18594 23060
rect 18580 22484 18594 22540
rect 18628 22540 18634 23060
rect 19606 23060 19652 23072
rect 18628 22484 18640 22540
rect 19606 22514 19612 23060
rect 18580 22324 18640 22484
rect 19594 22484 19612 22514
rect 19646 22514 19652 23060
rect 20616 23060 20676 23516
rect 21642 23516 21648 24028
rect 21682 24028 21692 24092
rect 22654 24092 22714 24342
rect 22948 24185 23436 24191
rect 22948 24151 22960 24185
rect 23424 24151 23436 24185
rect 22948 24145 23436 24151
rect 23966 24185 24454 24191
rect 23966 24151 23978 24185
rect 24442 24151 24454 24185
rect 23966 24145 24454 24151
rect 21682 23516 21688 24028
rect 21642 23504 21688 23516
rect 22654 23516 22666 24092
rect 22700 23516 22714 24092
rect 23678 24092 23724 24104
rect 23678 23580 23684 24092
rect 21122 23463 21182 23469
rect 20912 23457 21400 23463
rect 20912 23423 20924 23457
rect 21388 23423 21400 23457
rect 20912 23417 21400 23423
rect 21930 23457 22418 23463
rect 21930 23423 21942 23457
rect 22406 23423 22418 23457
rect 21930 23417 22418 23423
rect 21122 23260 21182 23417
rect 21626 23302 21632 23362
rect 21692 23302 21698 23362
rect 21122 23254 21184 23260
rect 21122 23194 21124 23254
rect 21122 23188 21184 23194
rect 21122 23159 21182 23188
rect 20912 23153 21400 23159
rect 20912 23119 20924 23153
rect 21388 23119 21400 23153
rect 20912 23113 21400 23119
rect 19646 22484 19654 22514
rect 18876 22425 19364 22431
rect 18876 22391 18888 22425
rect 19352 22391 19364 22425
rect 18876 22385 19364 22391
rect 19082 22324 19142 22385
rect 19594 22330 19654 22484
rect 20616 22484 20630 23060
rect 20664 22484 20676 23060
rect 21632 23060 21692 23302
rect 22144 23260 22204 23417
rect 22142 23254 22204 23260
rect 22202 23194 22204 23254
rect 22142 23188 22204 23194
rect 22144 23159 22204 23188
rect 21930 23153 22418 23159
rect 21930 23119 21942 23153
rect 22406 23119 22418 23153
rect 21930 23113 22418 23119
rect 22144 23106 22204 23113
rect 21632 23014 21648 23060
rect 19894 22425 20382 22431
rect 19894 22391 19906 22425
rect 20370 22391 20382 22425
rect 19894 22385 20382 22391
rect 19588 22324 19594 22330
rect 18454 22270 19594 22324
rect 19654 22270 19660 22330
rect 18454 22264 19660 22270
rect 20100 22196 20160 22385
rect 20100 22130 20160 22136
rect 20616 21988 20676 22484
rect 21642 22484 21648 23014
rect 21682 23014 21692 23060
rect 22654 23060 22714 23516
rect 23674 23516 23684 23580
rect 23718 23580 23724 24092
rect 24692 24092 24752 24342
rect 25694 24238 25700 24298
rect 25760 24238 25766 24298
rect 24984 24185 25472 24191
rect 24984 24151 24996 24185
rect 25460 24151 25472 24185
rect 24984 24145 25472 24151
rect 23718 23516 23734 23580
rect 22948 23457 23436 23463
rect 22948 23423 22960 23457
rect 23424 23423 23436 23457
rect 22948 23417 23436 23423
rect 23164 23260 23224 23417
rect 23674 23362 23734 23516
rect 24692 23516 24702 24092
rect 24736 23516 24752 24092
rect 25700 24092 25760 24238
rect 26002 24185 26490 24191
rect 26002 24151 26014 24185
rect 26478 24151 26490 24185
rect 26002 24145 26490 24151
rect 25700 24018 25720 24092
rect 24180 23463 24240 23465
rect 23966 23457 24454 23463
rect 23966 23423 23978 23457
rect 24442 23423 24454 23457
rect 23966 23417 24454 23423
rect 23668 23302 23674 23362
rect 23734 23302 23740 23362
rect 23164 23254 23226 23260
rect 23164 23194 23166 23254
rect 23164 23188 23226 23194
rect 24180 23254 24240 23417
rect 23164 23159 23224 23188
rect 24180 23159 24240 23194
rect 22948 23153 23436 23159
rect 22948 23119 22960 23153
rect 23424 23119 23436 23153
rect 22948 23113 23436 23119
rect 23966 23153 24454 23159
rect 23966 23119 23978 23153
rect 24442 23119 24454 23153
rect 23966 23113 24454 23119
rect 21682 22484 21688 23014
rect 21642 22472 21688 22484
rect 22654 22484 22666 23060
rect 22700 22484 22714 23060
rect 23678 23060 23724 23072
rect 23678 22550 23684 23060
rect 21114 22431 21174 22434
rect 20912 22425 21400 22431
rect 20912 22391 20924 22425
rect 21388 22391 21400 22425
rect 20912 22385 21400 22391
rect 21930 22425 22418 22431
rect 21930 22391 21942 22425
rect 22406 22391 22418 22425
rect 21930 22385 22418 22391
rect 21114 22192 21174 22385
rect 22146 22200 22206 22385
rect 22146 22134 22206 22140
rect 21114 22126 21174 22132
rect 22654 21988 22714 22484
rect 23674 22484 23684 22550
rect 23718 22550 23724 23060
rect 24692 23060 24752 23516
rect 25714 23516 25720 24018
rect 25754 23516 25760 24092
rect 25714 23504 25760 23516
rect 26728 24092 26788 24342
rect 27020 24185 27508 24191
rect 27020 24151 27032 24185
rect 27496 24151 27508 24185
rect 27020 24145 27508 24151
rect 28038 24185 28526 24191
rect 28038 24151 28050 24185
rect 28514 24151 28526 24185
rect 28038 24145 28526 24151
rect 26728 23516 26738 24092
rect 26772 23516 26788 24092
rect 27750 24092 27796 24104
rect 27750 23580 27756 24092
rect 24984 23457 25472 23463
rect 24984 23423 24996 23457
rect 25460 23423 25472 23457
rect 24984 23417 25472 23423
rect 26002 23457 26490 23463
rect 26002 23423 26014 23457
rect 26478 23423 26490 23457
rect 26002 23417 26490 23423
rect 25196 23260 25256 23417
rect 25694 23302 25700 23362
rect 25760 23302 25766 23362
rect 25196 23254 25258 23260
rect 25196 23194 25198 23254
rect 25196 23188 25258 23194
rect 25196 23159 25256 23188
rect 24984 23153 25472 23159
rect 24984 23119 24996 23153
rect 25460 23119 25472 23153
rect 24984 23113 25472 23119
rect 23718 22484 23734 22550
rect 22948 22425 23436 22431
rect 22948 22391 22960 22425
rect 23424 22391 23436 22425
rect 22948 22385 23436 22391
rect 23144 22200 23204 22385
rect 23674 22330 23734 22484
rect 24692 22484 24702 23060
rect 24736 22484 24752 23060
rect 25700 23060 25760 23302
rect 26206 23260 26266 23417
rect 26206 23254 26268 23260
rect 26206 23194 26208 23254
rect 26206 23188 26268 23194
rect 26206 23159 26266 23188
rect 26002 23153 26490 23159
rect 26002 23119 26014 23153
rect 26478 23119 26490 23153
rect 26002 23113 26490 23119
rect 25700 22998 25720 23060
rect 25714 22576 25720 22998
rect 24188 22431 24248 22444
rect 23966 22425 24454 22431
rect 23966 22391 23978 22425
rect 24442 22391 24454 22425
rect 23966 22385 24454 22391
rect 23668 22270 23674 22330
rect 23734 22270 23740 22330
rect 23144 22134 23204 22140
rect 24188 22200 24248 22385
rect 24188 22134 24248 22140
rect 24692 21988 24752 22484
rect 25710 22484 25720 22576
rect 25754 22576 25760 23060
rect 26728 23060 26788 23516
rect 27742 23516 27756 23580
rect 27790 23580 27796 24092
rect 28758 24092 28818 24342
rect 29770 24238 29776 24298
rect 29836 24238 29842 24298
rect 29056 24185 29544 24191
rect 29056 24151 29068 24185
rect 29532 24151 29544 24185
rect 29056 24145 29544 24151
rect 28758 23682 28774 24092
rect 28768 23588 28774 23682
rect 27790 23516 27802 23580
rect 27228 23463 27288 23465
rect 27020 23457 27508 23463
rect 27020 23423 27032 23457
rect 27496 23423 27508 23457
rect 27020 23417 27508 23423
rect 27228 23260 27288 23417
rect 27742 23362 27802 23516
rect 28758 23516 28774 23588
rect 28808 23682 28818 24092
rect 29776 24092 29836 24238
rect 30074 24185 30562 24191
rect 30074 24151 30086 24185
rect 30550 24151 30562 24185
rect 30074 24145 30562 24151
rect 29776 24028 29792 24092
rect 28808 23588 28814 23682
rect 28808 23516 28818 23588
rect 28242 23463 28302 23465
rect 28038 23457 28526 23463
rect 28038 23423 28050 23457
rect 28514 23423 28526 23457
rect 28038 23417 28526 23423
rect 27736 23302 27742 23362
rect 27802 23302 27808 23362
rect 28242 23260 28302 23417
rect 27228 23254 27290 23260
rect 27228 23194 27230 23254
rect 27228 23188 27290 23194
rect 28242 23254 28304 23260
rect 28242 23194 28244 23254
rect 28242 23188 28304 23194
rect 27228 23159 27288 23188
rect 28242 23159 28302 23188
rect 27020 23153 27508 23159
rect 27020 23119 27032 23153
rect 27496 23119 27508 23153
rect 27020 23113 27508 23119
rect 28038 23153 28526 23159
rect 28038 23119 28050 23153
rect 28514 23119 28526 23153
rect 28038 23113 28526 23119
rect 25754 22484 25770 22576
rect 25192 22431 25252 22434
rect 24984 22425 25472 22431
rect 24984 22391 24996 22425
rect 25460 22391 25472 22425
rect 24984 22385 25472 22391
rect 25192 22196 25252 22385
rect 25192 22130 25252 22136
rect 25710 22080 25770 22484
rect 26728 22484 26738 23060
rect 26772 22484 26788 23060
rect 27750 23060 27796 23072
rect 27750 22566 27756 23060
rect 26208 22431 26268 22438
rect 26002 22425 26490 22431
rect 26002 22391 26014 22425
rect 26478 22391 26490 22425
rect 26002 22385 26490 22391
rect 26208 22196 26268 22385
rect 26208 22130 26268 22136
rect 25500 22020 25770 22080
rect 20616 21928 24992 21988
rect 25052 21928 25058 21988
rect 18340 21798 22508 21858
rect 18218 21610 18224 21670
rect 18284 21610 18290 21670
rect 19384 21610 19390 21670
rect 19450 21610 19456 21670
rect 17950 20564 17956 20624
rect 18016 20564 18022 20624
rect 17708 19406 17714 19466
rect 17774 19406 17780 19466
rect 17704 19192 17710 19252
rect 17770 19192 17776 19252
rect 17592 18150 17598 18210
rect 17658 18150 17664 18210
rect 12254 16896 17524 16956
rect 12194 16890 12254 16896
rect -12293 16376 -7916 16436
rect -7856 16376 -7850 16436
rect -4464 16376 -4458 16436
rect -4398 16376 -4392 16436
rect -12293 16310 -11988 16376
rect -12293 16276 -12234 16310
rect -12014 16276 -11988 16310
rect -12293 16262 -11988 16276
rect -12293 16212 -12232 16262
rect -12293 16182 -12282 16212
rect -12292 15954 -12282 16182
rect -12293 15894 -12282 15954
rect -12292 15640 -12282 15894
rect -12244 15954 -12232 16212
rect -12182 16114 -12122 16262
rect -12048 16213 -11988 16262
rect -11792 16328 -11732 16329
rect -11016 16328 -10956 16334
rect -11792 16268 -11016 16328
rect -11792 16213 -11732 16268
rect -11534 16213 -11474 16268
rect -11276 16213 -11216 16268
rect -11016 16213 -10956 16268
rect -10760 16310 -10457 16376
rect -10760 16276 -10742 16310
rect -10540 16276 -10457 16310
rect -10760 16262 -10457 16276
rect -10760 16213 -10700 16262
rect -12074 16207 -11966 16213
rect -12074 16173 -12062 16207
rect -11978 16173 -11966 16207
rect -12074 16167 -11966 16173
rect -11816 16207 -11708 16213
rect -11816 16173 -11804 16207
rect -11720 16173 -11708 16207
rect -11816 16167 -11708 16173
rect -11558 16207 -11450 16213
rect -11558 16173 -11546 16207
rect -11462 16173 -11450 16207
rect -11558 16167 -11450 16173
rect -11300 16207 -11192 16213
rect -11300 16173 -11288 16207
rect -11204 16173 -11192 16207
rect -11300 16167 -11192 16173
rect -11042 16207 -10934 16213
rect -11042 16173 -11030 16207
rect -10946 16173 -10934 16207
rect -11042 16167 -10934 16173
rect -10784 16207 -10676 16213
rect -10784 16173 -10772 16207
rect -10688 16173 -10676 16207
rect -10784 16167 -10676 16173
rect -12182 15954 -12166 16114
rect -12244 15894 -12166 15954
rect -12244 15640 -12232 15894
rect -12172 15772 -12166 15894
rect -12292 15590 -12232 15640
rect -12180 15738 -12166 15772
rect -12132 15894 -12122 16114
rect -11914 16114 -11868 16126
rect -12132 15772 -12126 15894
rect -11914 15783 -11908 16114
rect -12132 15738 -12120 15772
rect -12180 15590 -12120 15738
rect -11922 15738 -11908 15783
rect -11874 15783 -11868 16114
rect -11656 16114 -11610 16126
rect -11874 15738 -11862 15783
rect -11656 15758 -11650 16114
rect -12074 15679 -11966 15685
rect -12074 15645 -12062 15679
rect -11978 15645 -11966 15679
rect -12074 15639 -11966 15645
rect -12052 15590 -11992 15639
rect -12293 15576 -11992 15590
rect -12293 15542 -12234 15576
rect -12014 15542 -11992 15576
rect -12293 15530 -11992 15542
rect -11922 15413 -11862 15738
rect -11664 15738 -11650 15758
rect -11616 15758 -11610 16114
rect -11398 16114 -11352 16126
rect -11398 15781 -11392 16114
rect -11616 15738 -11604 15758
rect -11816 15679 -11708 15685
rect -11816 15645 -11804 15679
rect -11720 15645 -11708 15679
rect -11816 15639 -11708 15645
rect -11664 15562 -11604 15738
rect -11406 15738 -11392 15781
rect -11358 15781 -11352 16114
rect -11140 16114 -11094 16126
rect -11358 15738 -11346 15781
rect -11140 15776 -11134 16114
rect -11558 15679 -11450 15685
rect -11558 15645 -11546 15679
rect -11462 15645 -11450 15679
rect -11558 15639 -11450 15645
rect -11670 15502 -11664 15562
rect -11604 15502 -11598 15562
rect -12294 15378 -11990 15388
rect -12294 15340 -12210 15378
rect -12002 15340 -11990 15378
rect -11928 15353 -11922 15413
rect -11862 15353 -11856 15413
rect -12294 15328 -11990 15340
rect -12294 15280 -12234 15328
rect -12294 14924 -12282 15280
rect -12246 14924 -12234 15280
rect -12180 15190 -12120 15328
rect -12050 15280 -11990 15328
rect -12074 15274 -11966 15280
rect -12074 15240 -12062 15274
rect -11978 15240 -11966 15274
rect -12074 15234 -11966 15240
rect -12180 15140 -12166 15190
rect -12172 15053 -12166 15140
rect -12294 14875 -12234 14924
rect -12178 15014 -12166 15053
rect -12132 15140 -12120 15190
rect -11922 15190 -11862 15353
rect -11816 15274 -11708 15280
rect -11816 15240 -11804 15274
rect -11720 15240 -11708 15274
rect -11816 15234 -11708 15240
rect -11922 15153 -11908 15190
rect -12132 15053 -12126 15140
rect -12132 15014 -12118 15053
rect -12178 14875 -12118 15014
rect -11914 15014 -11908 15153
rect -11874 15153 -11862 15190
rect -11664 15220 -11604 15502
rect -11406 15413 -11346 15738
rect -11146 15738 -11134 15776
rect -11100 15776 -11094 16114
rect -10882 16114 -10836 16126
rect -10882 15781 -10876 16114
rect -11100 15738 -11086 15776
rect -11300 15679 -11192 15685
rect -11300 15645 -11288 15679
rect -11204 15645 -11192 15679
rect -11300 15639 -11192 15645
rect -11146 15562 -11086 15738
rect -10888 15738 -10876 15781
rect -10842 15781 -10836 16114
rect -10632 16114 -10572 16262
rect -10632 15896 -10618 16114
rect -10842 15738 -10828 15781
rect -10624 15768 -10618 15896
rect -11042 15679 -10934 15685
rect -11042 15645 -11030 15679
rect -10946 15645 -10934 15679
rect -11042 15639 -10934 15645
rect -11152 15502 -11146 15562
rect -11086 15502 -11080 15562
rect -11412 15353 -11406 15413
rect -11346 15353 -11340 15413
rect -11558 15274 -11450 15280
rect -11558 15240 -11546 15274
rect -11462 15240 -11450 15274
rect -11558 15234 -11450 15240
rect -11664 15190 -11602 15220
rect -11664 15154 -11650 15190
rect -11874 15014 -11868 15153
rect -11914 15002 -11868 15014
rect -11662 15014 -11650 15154
rect -11616 15014 -11602 15190
rect -11406 15190 -11346 15353
rect -11300 15274 -11192 15280
rect -11300 15240 -11288 15274
rect -11204 15240 -11192 15274
rect -11300 15234 -11192 15240
rect -11406 15034 -11392 15190
rect -11662 14974 -11602 15014
rect -11398 15014 -11392 15034
rect -11358 15034 -11346 15190
rect -11146 15190 -11086 15502
rect -10888 15413 -10828 15738
rect -10630 15738 -10618 15768
rect -10584 15956 -10572 16114
rect -10518 16214 -10457 16262
rect -10518 15956 -10506 16214
rect -10584 15896 -10506 15956
rect -10584 15768 -10578 15896
rect -10584 15738 -10570 15768
rect -10784 15679 -10676 15685
rect -10784 15645 -10772 15679
rect -10688 15645 -10676 15679
rect -10784 15639 -10676 15645
rect -10764 15590 -10704 15639
rect -10630 15590 -10570 15738
rect -10518 15638 -10506 15896
rect -10470 16198 -10457 16214
rect -9693 16310 -9388 16376
rect -9693 16276 -9634 16310
rect -9414 16276 -9388 16310
rect -9693 16262 -9388 16276
rect -9693 16212 -9632 16262
rect -10470 15838 -10458 16198
rect -9693 16182 -9682 16212
rect -9692 15954 -9682 16182
rect -9693 15894 -9682 15954
rect -10470 15807 -10120 15838
rect -10470 15773 -10367 15807
rect -10333 15773 -10275 15807
rect -10241 15773 -10183 15807
rect -10149 15773 -10120 15807
rect -10470 15742 -10120 15773
rect -10470 15638 -10458 15742
rect -10518 15590 -10458 15638
rect -9692 15640 -9682 15894
rect -9644 15954 -9632 16212
rect -9582 16114 -9522 16262
rect -9448 16213 -9388 16262
rect -9192 16328 -9132 16329
rect -8416 16328 -8356 16334
rect -9192 16268 -8416 16328
rect -9192 16213 -9132 16268
rect -8934 16213 -8874 16268
rect -8676 16213 -8616 16268
rect -8416 16213 -8356 16268
rect -8160 16310 -7857 16376
rect -8160 16276 -8142 16310
rect -7940 16276 -7857 16310
rect -8160 16262 -7857 16276
rect -8160 16213 -8100 16262
rect -9474 16207 -9366 16213
rect -9474 16173 -9462 16207
rect -9378 16173 -9366 16207
rect -9474 16167 -9366 16173
rect -9216 16207 -9108 16213
rect -9216 16173 -9204 16207
rect -9120 16173 -9108 16207
rect -9216 16167 -9108 16173
rect -8958 16207 -8850 16213
rect -8958 16173 -8946 16207
rect -8862 16173 -8850 16207
rect -8958 16167 -8850 16173
rect -8700 16207 -8592 16213
rect -8700 16173 -8688 16207
rect -8604 16173 -8592 16207
rect -8700 16167 -8592 16173
rect -8442 16207 -8334 16213
rect -8442 16173 -8430 16207
rect -8346 16173 -8334 16207
rect -8442 16167 -8334 16173
rect -8184 16207 -8076 16213
rect -8184 16173 -8172 16207
rect -8088 16173 -8076 16207
rect -8184 16167 -8076 16173
rect -9582 15954 -9566 16114
rect -9644 15894 -9566 15954
rect -9644 15640 -9632 15894
rect -9572 15772 -9566 15894
rect -9692 15590 -9632 15640
rect -9580 15738 -9566 15772
rect -9532 15894 -9522 16114
rect -9314 16114 -9268 16126
rect -9532 15772 -9526 15894
rect -9314 15783 -9308 16114
rect -9532 15738 -9520 15772
rect -9580 15590 -9520 15738
rect -9322 15738 -9308 15783
rect -9274 15783 -9268 16114
rect -9056 16114 -9010 16126
rect -9274 15738 -9262 15783
rect -9056 15758 -9050 16114
rect -9474 15679 -9366 15685
rect -9474 15645 -9462 15679
rect -9378 15645 -9366 15679
rect -9474 15639 -9366 15645
rect -9452 15590 -9392 15639
rect -10764 15578 -10458 15590
rect -10764 15544 -10742 15578
rect -10540 15544 -10458 15578
rect -10764 15530 -10458 15544
rect -9693 15576 -9392 15590
rect -9693 15542 -9634 15576
rect -9414 15542 -9392 15576
rect -9693 15530 -9392 15542
rect -10025 15512 -9965 15518
rect -10245 15506 -10025 15512
rect -10343 15490 -10283 15496
rect -10349 15430 -10343 15490
rect -10283 15430 -10277 15490
rect -10245 15466 -10233 15506
rect -10187 15466 -10025 15506
rect -10245 15452 -10025 15466
rect -10025 15446 -9965 15452
rect -10343 15424 -10283 15430
rect -9322 15413 -9262 15738
rect -9064 15738 -9050 15758
rect -9016 15758 -9010 16114
rect -8798 16114 -8752 16126
rect -8798 15781 -8792 16114
rect -9016 15738 -9004 15758
rect -9216 15679 -9108 15685
rect -9216 15645 -9204 15679
rect -9120 15645 -9108 15679
rect -9216 15639 -9108 15645
rect -9064 15562 -9004 15738
rect -8806 15738 -8792 15781
rect -8758 15781 -8752 16114
rect -8540 16114 -8494 16126
rect -8758 15738 -8746 15781
rect -8540 15776 -8534 16114
rect -8958 15679 -8850 15685
rect -8958 15645 -8946 15679
rect -8862 15645 -8850 15679
rect -8958 15639 -8850 15645
rect -9070 15502 -9064 15562
rect -9004 15502 -8998 15562
rect -11042 15274 -10934 15280
rect -11042 15240 -11030 15274
rect -10946 15240 -10934 15274
rect -11042 15234 -10934 15240
rect -11358 15014 -11352 15034
rect -11398 15002 -11352 15014
rect -11146 15014 -11134 15190
rect -11100 15014 -11086 15190
rect -10888 15190 -10828 15353
rect -10758 15380 -10456 15390
rect -10758 15342 -10738 15380
rect -10540 15342 -10456 15380
rect -10758 15330 -10456 15342
rect -10758 15280 -10698 15330
rect -10784 15274 -10676 15280
rect -10784 15240 -10772 15274
rect -10688 15240 -10676 15274
rect -10784 15234 -10676 15240
rect -10888 15151 -10876 15190
rect -11146 14974 -11086 15014
rect -10882 15014 -10876 15151
rect -10842 15151 -10828 15190
rect -10630 15190 -10570 15330
rect -10842 15014 -10836 15151
rect -10630 15144 -10618 15190
rect -10624 15047 -10618 15144
rect -10882 15002 -10836 15014
rect -10632 15014 -10618 15047
rect -10584 15144 -10570 15190
rect -10516 15294 -10456 15330
rect -9694 15378 -9390 15388
rect -9694 15340 -9610 15378
rect -9402 15340 -9390 15378
rect -9328 15353 -9322 15413
rect -9262 15353 -9256 15413
rect -9694 15328 -9390 15340
rect -10516 15280 -10120 15294
rect -10584 15047 -10578 15144
rect -10584 15014 -10572 15047
rect -12074 14964 -11966 14970
rect -12074 14930 -12062 14964
rect -11978 14930 -11966 14964
rect -12074 14924 -11966 14930
rect -11816 14964 -11708 14970
rect -11816 14930 -11804 14964
rect -11720 14930 -11708 14964
rect -11816 14924 -11708 14930
rect -11558 14964 -11450 14970
rect -11558 14930 -11546 14964
rect -11462 14930 -11450 14964
rect -11558 14924 -11450 14930
rect -11300 14964 -11192 14970
rect -11300 14930 -11288 14964
rect -11204 14930 -11192 14964
rect -11300 14924 -11192 14930
rect -11042 14964 -10934 14970
rect -11042 14930 -11030 14964
rect -10946 14930 -10934 14964
rect -11042 14924 -10934 14930
rect -10784 14964 -10676 14970
rect -10784 14930 -10772 14964
rect -10688 14930 -10676 14964
rect -10784 14924 -10676 14930
rect -12050 14875 -11990 14924
rect -12294 14864 -11990 14875
rect -12294 14828 -12212 14864
rect -12004 14828 -11990 14864
rect -12294 14758 -11990 14828
rect -11792 14865 -11732 14924
rect -11532 14865 -11472 14924
rect -11274 14865 -11214 14924
rect -11018 14865 -10958 14924
rect -10760 14875 -10700 14924
rect -10632 14875 -10572 15014
rect -10516 14924 -10506 15280
rect -10468 15263 -10120 15280
rect -10468 15229 -10367 15263
rect -10333 15229 -10275 15263
rect -10241 15229 -10183 15263
rect -10149 15229 -10120 15263
rect -10468 15198 -10120 15229
rect -9694 15280 -9634 15328
rect -10468 14924 -10456 15198
rect -10516 14875 -10456 14924
rect -11792 14805 -11018 14865
rect -10958 14805 -10952 14865
rect -10760 14862 -10456 14875
rect -10760 14826 -10740 14862
rect -10538 14826 -10456 14862
rect -12293 14740 -11990 14758
rect -10760 14740 -10456 14826
rect -9694 14924 -9682 15280
rect -9646 14924 -9634 15280
rect -9580 15190 -9520 15328
rect -9450 15280 -9390 15328
rect -9474 15274 -9366 15280
rect -9474 15240 -9462 15274
rect -9378 15240 -9366 15274
rect -9474 15234 -9366 15240
rect -9580 15140 -9566 15190
rect -9572 15053 -9566 15140
rect -9694 14875 -9634 14924
rect -9578 15014 -9566 15053
rect -9532 15140 -9520 15190
rect -9322 15190 -9262 15353
rect -9216 15274 -9108 15280
rect -9216 15240 -9204 15274
rect -9120 15240 -9108 15274
rect -9216 15234 -9108 15240
rect -9322 15153 -9308 15190
rect -9532 15053 -9526 15140
rect -9532 15014 -9518 15053
rect -9578 14875 -9518 15014
rect -9314 15014 -9308 15153
rect -9274 15153 -9262 15190
rect -9064 15220 -9004 15502
rect -8806 15413 -8746 15738
rect -8546 15738 -8534 15776
rect -8500 15776 -8494 16114
rect -8282 16114 -8236 16126
rect -8282 15781 -8276 16114
rect -8500 15738 -8486 15776
rect -8700 15679 -8592 15685
rect -8700 15645 -8688 15679
rect -8604 15645 -8592 15679
rect -8700 15639 -8592 15645
rect -8546 15562 -8486 15738
rect -8288 15738 -8276 15781
rect -8242 15781 -8236 16114
rect -8032 16114 -7972 16262
rect -8032 15896 -8018 16114
rect -8242 15738 -8228 15781
rect -8024 15768 -8018 15896
rect -8442 15679 -8334 15685
rect -8442 15645 -8430 15679
rect -8346 15645 -8334 15679
rect -8442 15639 -8334 15645
rect -8552 15502 -8546 15562
rect -8486 15502 -8480 15562
rect -8812 15353 -8806 15413
rect -8746 15353 -8740 15413
rect -8958 15274 -8850 15280
rect -8958 15240 -8946 15274
rect -8862 15240 -8850 15274
rect -8958 15234 -8850 15240
rect -9064 15190 -9002 15220
rect -9064 15154 -9050 15190
rect -9274 15014 -9268 15153
rect -9314 15002 -9268 15014
rect -9062 15014 -9050 15154
rect -9016 15014 -9002 15190
rect -8806 15190 -8746 15353
rect -8700 15274 -8592 15280
rect -8700 15240 -8688 15274
rect -8604 15240 -8592 15274
rect -8700 15234 -8592 15240
rect -8806 15034 -8792 15190
rect -9062 14974 -9002 15014
rect -8798 15014 -8792 15034
rect -8758 15034 -8746 15190
rect -8546 15190 -8486 15502
rect -8288 15413 -8228 15738
rect -8030 15738 -8018 15768
rect -7984 15956 -7972 16114
rect -7918 16214 -7857 16262
rect -7918 15956 -7906 16214
rect -7984 15896 -7906 15956
rect -7984 15768 -7978 15896
rect -7984 15738 -7970 15768
rect -8184 15679 -8076 15685
rect -8184 15645 -8172 15679
rect -8088 15645 -8076 15679
rect -8184 15639 -8076 15645
rect -8164 15590 -8104 15639
rect -8030 15590 -7970 15738
rect -7918 15638 -7906 15896
rect -7870 16198 -7857 16214
rect -3080 16358 8190 16418
rect -7870 15838 -7858 16198
rect -3080 15870 -3014 16358
rect -2786 16162 8190 16358
rect 11284 16298 11396 16812
rect 13248 16694 13308 16700
rect 17710 16694 17770 19192
rect 17956 16952 18016 20564
rect 18086 20466 18092 20526
rect 18152 20466 18158 20526
rect 17950 16892 17956 16952
rect 18016 16892 18022 16952
rect 18092 16822 18152 20466
rect 18224 18002 18284 21610
rect 18668 21549 19156 21555
rect 18668 21515 18680 21549
rect 19144 21515 19156 21549
rect 18668 21509 19156 21515
rect 18380 21456 18426 21468
rect 18380 20916 18386 21456
rect 18372 20880 18386 20916
rect 18420 20916 18426 21456
rect 19390 21456 19450 21610
rect 19686 21549 20174 21555
rect 19686 21515 19698 21549
rect 20162 21515 20174 21549
rect 19686 21509 20174 21515
rect 19390 21430 19404 21456
rect 18420 20880 18432 20916
rect 19398 20904 19404 21430
rect 18372 20722 18432 20880
rect 19388 20880 19404 20904
rect 19438 21430 19450 21456
rect 20406 21456 20466 21798
rect 21420 21610 21426 21670
rect 21486 21610 21492 21670
rect 20704 21549 21192 21555
rect 20704 21515 20716 21549
rect 21180 21515 21192 21549
rect 20704 21509 21192 21515
rect 19438 20904 19444 21430
rect 20406 21410 20422 21456
rect 20416 20904 20422 21410
rect 19438 20880 19448 20904
rect 18668 20821 19156 20827
rect 18668 20787 18680 20821
rect 19144 20787 19156 20821
rect 18668 20781 19156 20787
rect 18886 20722 18946 20781
rect 19388 20722 19448 20880
rect 20408 20880 20422 20904
rect 20456 21410 20466 21456
rect 21426 21456 21486 21610
rect 21928 21606 21934 21670
rect 21998 21606 22004 21670
rect 21934 21555 21998 21606
rect 21722 21549 22210 21555
rect 21722 21515 21734 21549
rect 22198 21515 22210 21549
rect 21722 21509 22210 21515
rect 21426 21432 21440 21456
rect 20456 20904 20462 21410
rect 20456 20880 20468 20904
rect 19686 20821 20174 20827
rect 19686 20787 19698 20821
rect 20162 20787 20174 20821
rect 19686 20781 20174 20787
rect 18372 20662 19448 20722
rect 19878 20420 19938 20781
rect 20408 20722 20468 20880
rect 21434 20880 21440 21432
rect 21474 21432 21486 21456
rect 22448 21456 22508 21798
rect 22952 21555 23012 21928
rect 22740 21549 23228 21555
rect 22740 21515 22752 21549
rect 23216 21515 23228 21549
rect 22740 21509 23228 21515
rect 21474 20880 21480 21432
rect 22448 21402 22458 21456
rect 22452 20908 22458 21402
rect 21434 20868 21480 20880
rect 22444 20880 22458 20908
rect 22492 21402 22508 21456
rect 23460 21456 23520 21928
rect 23952 21555 24012 21928
rect 24990 21555 25050 21928
rect 23758 21549 24246 21555
rect 23758 21515 23770 21549
rect 24234 21515 24246 21549
rect 23758 21509 24246 21515
rect 24776 21549 25264 21555
rect 24776 21515 24788 21549
rect 25252 21515 25264 21549
rect 24776 21509 25264 21515
rect 22492 20908 22498 21402
rect 22492 20880 22504 20908
rect 20704 20821 21192 20827
rect 20704 20787 20716 20821
rect 21180 20787 21192 20821
rect 20704 20781 21192 20787
rect 21722 20821 22210 20827
rect 21722 20787 21734 20821
rect 22198 20787 22210 20821
rect 21722 20781 22210 20787
rect 20402 20662 20408 20722
rect 20468 20662 20474 20722
rect 20916 20668 20976 20781
rect 21922 20668 21982 20781
rect 22444 20722 22504 20880
rect 23460 20880 23476 21456
rect 23510 20880 23520 21456
rect 24488 21456 24534 21468
rect 24488 20904 24494 21456
rect 22740 20821 23228 20827
rect 22740 20787 22752 20821
rect 23216 20787 23228 20821
rect 22740 20781 23228 20787
rect 22954 20726 23014 20781
rect 23460 20726 23520 20880
rect 24480 20880 24494 20904
rect 24528 20904 24534 21456
rect 25500 21456 25560 22020
rect 26728 21988 26788 22484
rect 27742 22484 27756 22566
rect 27790 22566 27796 23060
rect 28758 23060 28818 23516
rect 29786 23516 29792 24028
rect 29826 24028 29836 24092
rect 30796 24092 30856 24342
rect 32966 24238 32972 24298
rect 33032 24238 33038 24298
rect 31092 24185 31580 24191
rect 31092 24151 31104 24185
rect 31568 24151 31580 24185
rect 31092 24145 31580 24151
rect 32110 24185 32598 24191
rect 32110 24151 32122 24185
rect 32586 24151 32598 24185
rect 32110 24145 32598 24151
rect 29826 23516 29832 24028
rect 29786 23504 29832 23516
rect 30796 23516 30810 24092
rect 30844 23516 30856 24092
rect 31822 24092 31868 24104
rect 31822 23592 31828 24092
rect 29274 23463 29334 23465
rect 30284 23463 30344 23465
rect 29056 23457 29544 23463
rect 29056 23423 29068 23457
rect 29532 23423 29544 23457
rect 29056 23417 29544 23423
rect 30074 23457 30562 23463
rect 30074 23423 30086 23457
rect 30550 23423 30562 23457
rect 30074 23417 30562 23423
rect 29274 23260 29334 23417
rect 29772 23302 29778 23362
rect 29838 23302 29844 23362
rect 29274 23254 29336 23260
rect 29274 23194 29276 23254
rect 29274 23188 29336 23194
rect 29274 23159 29334 23188
rect 29056 23153 29544 23159
rect 29056 23119 29068 23153
rect 29532 23119 29544 23153
rect 29056 23113 29544 23119
rect 27790 22484 27802 22566
rect 27020 22425 27508 22431
rect 27020 22391 27032 22425
rect 27496 22391 27508 22425
rect 27020 22385 27508 22391
rect 27212 22196 27272 22385
rect 27742 22330 27802 22484
rect 28758 22484 28774 23060
rect 28808 22484 28818 23060
rect 29778 23060 29838 23302
rect 30284 23260 30344 23417
rect 30284 23254 30346 23260
rect 30284 23194 30286 23254
rect 30284 23188 30346 23194
rect 30284 23159 30344 23188
rect 30074 23153 30562 23159
rect 30074 23119 30086 23153
rect 30550 23119 30562 23153
rect 30074 23113 30562 23119
rect 29778 22992 29792 23060
rect 28038 22425 28526 22431
rect 28038 22391 28050 22425
rect 28514 22391 28526 22425
rect 28038 22385 28526 22391
rect 27736 22270 27742 22330
rect 27802 22270 27808 22330
rect 27212 22130 27272 22136
rect 28244 22200 28304 22385
rect 28244 22134 28304 22140
rect 26002 21728 26008 21792
rect 26072 21728 26078 21792
rect 26008 21670 26072 21728
rect 26728 21698 26788 21928
rect 28758 22088 28818 22484
rect 29786 22484 29792 22992
rect 29826 22992 29838 23060
rect 30796 23060 30856 23516
rect 31814 23516 31828 23592
rect 31862 23592 31868 24092
rect 32840 24092 32886 24104
rect 31862 23516 31874 23592
rect 32840 23542 32846 24092
rect 31092 23457 31580 23463
rect 31092 23423 31104 23457
rect 31568 23423 31580 23457
rect 31092 23417 31580 23423
rect 31306 23260 31366 23417
rect 31814 23364 31874 23516
rect 32830 23516 32846 23542
rect 32880 23542 32886 24092
rect 32880 23516 32890 23542
rect 32110 23457 32598 23463
rect 32110 23423 32122 23457
rect 32586 23423 32598 23457
rect 32110 23417 32598 23423
rect 32336 23364 32396 23417
rect 32830 23364 32890 23516
rect 31814 23362 32890 23364
rect 31808 23302 31814 23362
rect 31874 23304 32890 23362
rect 31874 23302 31880 23304
rect 31306 23254 31368 23260
rect 31306 23194 31308 23254
rect 31306 23188 31368 23194
rect 31306 23159 31366 23188
rect 31092 23153 31580 23159
rect 31092 23119 31104 23153
rect 31568 23119 31580 23153
rect 31092 23113 31580 23119
rect 32110 23153 32598 23159
rect 32110 23119 32122 23153
rect 32586 23119 32598 23153
rect 32110 23113 32598 23119
rect 29826 22484 29832 22992
rect 29786 22472 29832 22484
rect 30796 22484 30810 23060
rect 30844 22484 30856 23060
rect 31822 23060 31868 23072
rect 31822 22560 31828 23060
rect 29260 22431 29320 22434
rect 29056 22425 29544 22431
rect 29056 22391 29068 22425
rect 29532 22391 29544 22425
rect 29056 22385 29544 22391
rect 30074 22425 30562 22431
rect 30074 22391 30086 22425
rect 30550 22391 30562 22425
rect 30074 22385 30562 22391
rect 29260 22196 29320 22385
rect 29260 22130 29320 22136
rect 30288 22196 30348 22385
rect 30288 22130 30348 22136
rect 30796 22088 30856 22484
rect 31810 22484 31828 22560
rect 31862 22560 31868 23060
rect 32840 23060 32886 23072
rect 31862 22484 31870 22560
rect 32840 22556 32846 23060
rect 31308 22431 31368 22434
rect 31092 22425 31580 22431
rect 31092 22391 31104 22425
rect 31568 22391 31580 22425
rect 31092 22385 31580 22391
rect 31308 22196 31368 22385
rect 31810 22334 31870 22484
rect 32830 22484 32846 22556
rect 32880 22556 32886 23060
rect 32880 22484 32890 22556
rect 32110 22425 32598 22431
rect 32110 22391 32122 22425
rect 32586 22391 32598 22425
rect 32110 22385 32598 22391
rect 32298 22334 32358 22385
rect 32830 22334 32890 22484
rect 32972 22334 33032 24238
rect 31808 22330 33032 22334
rect 31804 22270 31810 22330
rect 31870 22274 33032 22330
rect 31870 22270 31876 22274
rect 33760 22138 33766 22198
rect 33826 22138 33832 22198
rect 31308 22130 31368 22136
rect 28758 22028 30856 22088
rect 28758 21698 28818 22028
rect 32620 21912 32626 21972
rect 32686 21912 32692 21972
rect 30066 21728 30072 21792
rect 30136 21728 30142 21792
rect 31090 21728 31096 21792
rect 31160 21728 31166 21792
rect 32102 21728 32108 21792
rect 32172 21728 32178 21792
rect 26004 21606 26010 21670
rect 26074 21606 26080 21670
rect 26728 21638 29122 21698
rect 30072 21674 30136 21728
rect 26008 21555 26072 21606
rect 27040 21555 27100 21638
rect 25794 21549 26282 21555
rect 25794 21515 25806 21549
rect 26270 21515 26282 21549
rect 25794 21509 26282 21515
rect 26812 21549 27300 21555
rect 26812 21515 26824 21549
rect 27288 21515 27300 21549
rect 26812 21509 27300 21515
rect 24528 20880 24540 20904
rect 23758 20821 24246 20827
rect 23758 20787 23770 20821
rect 24234 20787 24246 20821
rect 23758 20781 24246 20787
rect 23974 20726 24034 20781
rect 24480 20726 24540 20880
rect 25500 20880 25512 21456
rect 25546 20880 25560 21456
rect 26524 21456 26570 21468
rect 26524 20958 26530 21456
rect 24776 20821 25264 20827
rect 24776 20787 24788 20821
rect 25252 20787 25264 20821
rect 24776 20781 25264 20787
rect 24984 20726 25044 20781
rect 20408 20526 20468 20662
rect 20916 20608 21982 20668
rect 22438 20662 22444 20722
rect 22504 20662 22510 20722
rect 22780 20664 22786 20724
rect 22846 20664 22852 20724
rect 22954 20666 25044 20726
rect 25500 20724 25560 20880
rect 26518 20880 26530 20958
rect 26564 20958 26570 21456
rect 27534 21456 27594 21638
rect 28062 21555 28122 21638
rect 27830 21549 28318 21555
rect 27830 21515 27842 21549
rect 28306 21515 28318 21549
rect 27830 21509 28318 21515
rect 28062 21508 28122 21509
rect 26564 20880 26578 20958
rect 25794 20821 26282 20827
rect 25794 20787 25806 20821
rect 26270 20787 26282 20821
rect 25794 20781 26282 20787
rect 20402 20466 20408 20526
rect 20468 20466 20474 20526
rect 20916 20420 20976 20608
rect 21422 20468 21428 20528
rect 21488 20468 21494 20528
rect 19388 20356 19394 20416
rect 19454 20356 19460 20416
rect 19878 20360 20976 20420
rect 21428 20416 21488 20468
rect 18668 20293 19156 20299
rect 18668 20259 18680 20293
rect 19144 20259 19156 20293
rect 18668 20253 19156 20259
rect 18380 20200 18426 20212
rect 18380 19660 18386 20200
rect 18376 19624 18386 19660
rect 18420 19660 18426 20200
rect 19394 20200 19454 20356
rect 19878 20299 19938 20360
rect 20916 20299 20976 20360
rect 21422 20356 21428 20416
rect 21488 20356 21494 20416
rect 19686 20293 20174 20299
rect 19686 20259 19698 20293
rect 20162 20259 20174 20293
rect 19686 20253 20174 20259
rect 20704 20293 21192 20299
rect 20704 20259 20716 20293
rect 21180 20259 21192 20293
rect 20704 20253 21192 20259
rect 19394 20174 19404 20200
rect 18420 19624 18436 19660
rect 19398 19648 19404 20174
rect 18376 19466 18436 19624
rect 19392 19624 19404 19648
rect 19438 20174 19454 20200
rect 20416 20200 20462 20212
rect 19438 19648 19444 20174
rect 20416 19650 20422 20200
rect 19438 19624 19452 19648
rect 18668 19565 19156 19571
rect 18668 19531 18680 19565
rect 19144 19531 19156 19565
rect 18668 19525 19156 19531
rect 18890 19466 18950 19525
rect 19392 19466 19452 19624
rect 20410 19624 20422 19650
rect 20456 19650 20462 20200
rect 21428 20200 21488 20356
rect 21922 20299 21982 20608
rect 22786 20410 22846 20664
rect 22444 20350 22846 20410
rect 21722 20293 22210 20299
rect 21722 20259 21734 20293
rect 22198 20259 22210 20293
rect 21722 20253 22210 20259
rect 21428 20178 21440 20200
rect 20456 19624 20470 19650
rect 19872 19571 19932 19572
rect 19686 19565 20174 19571
rect 19686 19531 19698 19565
rect 20162 19531 20174 19565
rect 19686 19525 20174 19531
rect 18376 19406 19452 19466
rect 18376 19252 18436 19406
rect 18370 19192 18376 19252
rect 18436 19192 18442 19252
rect 18374 19082 19450 19142
rect 18374 18944 18434 19082
rect 18888 19043 18948 19082
rect 18668 19037 19156 19043
rect 18668 19003 18680 19037
rect 19144 19003 19156 19037
rect 18668 18997 19156 19003
rect 18374 18910 18386 18944
rect 18380 18368 18386 18910
rect 18420 18910 18434 18944
rect 19390 18944 19450 19082
rect 19872 19043 19932 19525
rect 20410 19362 20470 19624
rect 21434 19624 21440 20178
rect 21474 20178 21488 20200
rect 22444 20200 22504 20350
rect 22740 20293 23228 20299
rect 22740 20259 22752 20293
rect 23216 20259 23228 20293
rect 22740 20253 23228 20259
rect 21474 19624 21480 20178
rect 22444 20142 22458 20200
rect 22452 19654 22458 20142
rect 21434 19612 21480 19624
rect 22446 19624 22458 19654
rect 22492 20142 22504 20200
rect 23460 20200 23520 20666
rect 25494 20664 25500 20724
rect 25560 20664 25566 20724
rect 26518 20528 26578 20880
rect 27534 20880 27548 21456
rect 27582 20880 27594 21456
rect 26812 20821 27300 20827
rect 26812 20787 26824 20821
rect 27288 20787 27300 20821
rect 26812 20781 27300 20787
rect 27028 20726 27088 20781
rect 27534 20726 27594 20880
rect 28550 21456 28610 21638
rect 29062 21555 29122 21638
rect 29566 21610 29572 21670
rect 29632 21610 29638 21670
rect 28848 21549 29336 21555
rect 28848 21515 28860 21549
rect 29324 21515 29336 21549
rect 28848 21509 29336 21515
rect 29062 21502 29122 21509
rect 28550 20880 28566 21456
rect 28600 20880 28610 21456
rect 29572 21456 29632 21610
rect 30072 21555 30136 21610
rect 31096 21555 31160 21728
rect 31600 21610 31606 21670
rect 31666 21610 31672 21670
rect 29866 21549 30354 21555
rect 29866 21515 29878 21549
rect 30342 21515 30354 21549
rect 29866 21509 30354 21515
rect 30884 21549 31372 21555
rect 30884 21515 30896 21549
rect 31360 21515 31372 21549
rect 30884 21509 31372 21515
rect 29572 21428 29584 21456
rect 27830 20821 28318 20827
rect 27830 20787 27842 20821
rect 28306 20787 28318 20821
rect 27830 20781 28318 20787
rect 28054 20726 28114 20781
rect 28550 20726 28610 20880
rect 29578 20880 29584 21428
rect 29618 21428 29632 21456
rect 30596 21456 30642 21468
rect 29618 20880 29624 21428
rect 30596 20904 30602 21456
rect 29578 20868 29624 20880
rect 30588 20880 30602 20904
rect 30636 20904 30642 21456
rect 31606 21456 31666 21610
rect 32108 21555 32172 21728
rect 32626 21674 32686 21912
rect 32626 21614 33702 21674
rect 31902 21549 32390 21555
rect 31902 21515 31914 21549
rect 32378 21515 32390 21549
rect 31902 21509 32390 21515
rect 31606 21432 31620 21456
rect 30636 20880 30648 20904
rect 28848 20821 29336 20827
rect 28848 20787 28860 20821
rect 29324 20787 29336 20821
rect 28848 20781 29336 20787
rect 29866 20821 30354 20827
rect 29866 20787 29878 20821
rect 30342 20787 30354 20821
rect 29866 20781 30354 20787
rect 29066 20726 29126 20781
rect 27028 20666 29126 20726
rect 26512 20468 26518 20528
rect 26578 20468 26584 20528
rect 24478 20354 24484 20414
rect 24544 20354 24550 20414
rect 26512 20354 26518 20414
rect 26578 20354 26584 20414
rect 23758 20293 24246 20299
rect 23758 20259 23770 20293
rect 24234 20259 24246 20293
rect 23758 20253 24246 20259
rect 23460 20156 23476 20200
rect 22492 19654 22498 20142
rect 23470 19654 23476 20156
rect 22492 19624 22506 19654
rect 20910 19571 20970 19572
rect 21916 19571 21976 19572
rect 20704 19565 21192 19571
rect 20704 19531 20716 19565
rect 21180 19531 21192 19565
rect 20704 19525 21192 19531
rect 21722 19565 22210 19571
rect 21722 19531 21734 19565
rect 22198 19531 22210 19565
rect 21722 19525 22210 19531
rect 20410 19296 20470 19302
rect 20404 19098 20410 19158
rect 20470 19098 20476 19158
rect 19686 19037 20174 19043
rect 19686 19003 19698 19037
rect 20162 19003 20174 19037
rect 19686 18997 20174 19003
rect 19390 18922 19404 18944
rect 18420 18368 18426 18910
rect 19398 18396 19404 18922
rect 18380 18356 18426 18368
rect 19392 18368 19404 18396
rect 19438 18922 19450 18944
rect 20410 18944 20470 19098
rect 20910 19043 20970 19525
rect 21916 19043 21976 19525
rect 22446 19362 22506 19624
rect 23462 19624 23476 19654
rect 23510 20156 23520 20200
rect 24484 20200 24544 20354
rect 24776 20293 25264 20299
rect 24776 20259 24788 20293
rect 25252 20259 25264 20293
rect 24776 20253 25264 20259
rect 25794 20293 26282 20299
rect 25794 20259 25806 20293
rect 26270 20259 26282 20293
rect 25794 20253 26282 20259
rect 24484 20172 24494 20200
rect 23510 19654 23516 20156
rect 23510 19624 23522 19654
rect 22740 19565 23228 19571
rect 22740 19531 22752 19565
rect 23216 19531 23228 19565
rect 22740 19525 23228 19531
rect 22966 19470 23026 19525
rect 23462 19470 23522 19624
rect 24488 19624 24494 20172
rect 24528 20172 24544 20200
rect 25506 20200 25552 20212
rect 24528 19624 24534 20172
rect 25506 19648 25512 20200
rect 24488 19612 24534 19624
rect 25500 19624 25512 19648
rect 25546 19648 25552 20200
rect 26518 20200 26578 20354
rect 26812 20293 27300 20299
rect 26812 20259 26824 20293
rect 27288 20259 27300 20293
rect 26812 20253 27300 20259
rect 27830 20293 28318 20299
rect 27830 20259 27842 20293
rect 28306 20259 28318 20293
rect 27830 20253 28318 20259
rect 26518 20170 26530 20200
rect 26524 19652 26530 20170
rect 25546 19624 25560 19648
rect 23758 19565 24246 19571
rect 23758 19531 23770 19565
rect 24234 19531 24246 19565
rect 23758 19525 24246 19531
rect 24776 19565 25264 19571
rect 24776 19531 24788 19565
rect 25252 19531 25264 19565
rect 24776 19525 25264 19531
rect 23978 19470 24038 19525
rect 22966 19410 24038 19470
rect 22440 19302 22446 19362
rect 22506 19302 22512 19362
rect 22438 19200 22444 19260
rect 22504 19200 22510 19260
rect 22444 19158 22504 19200
rect 22438 19098 22444 19158
rect 22504 19098 22510 19158
rect 20704 19037 21192 19043
rect 20704 19003 20716 19037
rect 21180 19003 21192 19037
rect 20704 18997 21192 19003
rect 21722 19037 22210 19043
rect 21722 19003 21734 19037
rect 22198 19003 22210 19037
rect 21722 18997 22210 19003
rect 19438 18396 19444 18922
rect 20410 18920 20422 18944
rect 19438 18368 19452 18396
rect 18668 18309 19156 18315
rect 18668 18275 18680 18309
rect 19144 18275 19156 18309
rect 18668 18269 19156 18275
rect 19392 18210 19452 18368
rect 20416 18368 20422 18920
rect 20456 18920 20470 18944
rect 21434 18944 21480 18956
rect 20456 18368 20462 18920
rect 21434 18392 21440 18944
rect 20416 18356 20462 18368
rect 21428 18368 21440 18392
rect 21474 18392 21480 18944
rect 22444 18944 22504 19098
rect 22740 19037 23228 19043
rect 22740 19003 22752 19037
rect 23216 19003 23228 19037
rect 22740 18997 23228 19003
rect 22444 18916 22458 18944
rect 21474 18368 21488 18392
rect 22452 18387 22458 18916
rect 19884 18315 19944 18322
rect 20922 18315 20982 18322
rect 19686 18309 20174 18315
rect 19686 18275 19698 18309
rect 20162 18275 20174 18309
rect 19686 18269 20174 18275
rect 20704 18309 21192 18315
rect 20704 18275 20716 18309
rect 21180 18275 21192 18309
rect 20704 18269 21192 18275
rect 19386 18150 19392 18210
rect 19452 18150 19458 18210
rect 18218 17942 18224 18002
rect 18284 17942 18290 18002
rect 18374 17844 19450 17904
rect 18374 17688 18434 17844
rect 18888 17787 18948 17844
rect 18668 17781 19156 17787
rect 18668 17747 18680 17781
rect 19144 17747 19156 17781
rect 18668 17741 19156 17747
rect 18374 17650 18386 17688
rect 18380 17112 18386 17650
rect 18420 17650 18434 17688
rect 19390 17688 19450 17844
rect 19884 17787 19944 18269
rect 20400 17840 20406 17900
rect 20466 17840 20472 17900
rect 19686 17781 20174 17787
rect 19686 17747 19698 17781
rect 20162 17747 20174 17781
rect 19686 17741 20174 17747
rect 19390 17662 19404 17688
rect 18420 17112 18426 17650
rect 19398 17138 19404 17662
rect 18380 17100 18426 17112
rect 19388 17112 19404 17138
rect 19438 17662 19450 17688
rect 20406 17688 20466 17840
rect 20922 17787 20982 18269
rect 21428 18210 21488 18368
rect 22446 18368 22458 18387
rect 22492 18916 22504 18944
rect 23462 18944 23522 19410
rect 24474 19406 24480 19466
rect 24540 19406 24546 19466
rect 23758 19037 24246 19043
rect 23758 19003 23770 19037
rect 24234 19003 24246 19037
rect 23758 18997 24246 19003
rect 22492 18387 22498 18916
rect 23462 18906 23476 18944
rect 23470 18402 23476 18906
rect 22492 18368 22506 18387
rect 21928 18315 21988 18322
rect 21722 18309 22210 18315
rect 21722 18275 21734 18309
rect 22198 18275 22210 18309
rect 21722 18269 22210 18275
rect 21422 18150 21428 18210
rect 21488 18150 21494 18210
rect 21428 18102 21488 18150
rect 21422 18042 21428 18102
rect 21488 18042 21494 18102
rect 21928 18052 21988 18269
rect 22446 18218 22506 18368
rect 23460 18368 23476 18402
rect 23510 18906 23522 18944
rect 24480 18944 24540 19406
rect 24982 19304 25042 19525
rect 25500 19466 25560 19624
rect 26518 19624 26530 19652
rect 26564 20170 26578 20200
rect 27542 20200 27588 20212
rect 26564 19652 26570 20170
rect 27542 19652 27548 20200
rect 26564 19624 26578 19652
rect 26012 19571 26072 19578
rect 25794 19565 26282 19571
rect 25794 19531 25806 19565
rect 26270 19531 26282 19565
rect 25794 19525 26282 19531
rect 25494 19406 25500 19466
rect 25560 19406 25566 19466
rect 26012 19304 26072 19525
rect 24982 19244 26072 19304
rect 24982 19043 25042 19244
rect 25494 19100 25500 19160
rect 25560 19100 25566 19160
rect 24776 19037 25264 19043
rect 24776 19003 24788 19037
rect 25252 19003 25264 19037
rect 24776 18997 25264 19003
rect 24982 18992 25042 18997
rect 24480 18920 24494 18944
rect 23510 18402 23516 18906
rect 23510 18368 23520 18402
rect 24488 18398 24494 18920
rect 22740 18309 23228 18315
rect 22740 18275 22752 18309
rect 23216 18275 23228 18309
rect 22740 18269 23228 18275
rect 22964 18218 23024 18269
rect 23460 18218 23520 18368
rect 24482 18368 24494 18398
rect 24528 18920 24540 18944
rect 25500 18944 25560 19100
rect 26012 19043 26072 19244
rect 26518 19160 26578 19624
rect 27536 19624 27548 19652
rect 27582 19652 27588 20200
rect 28550 20200 28610 20666
rect 29568 20354 29574 20414
rect 29634 20354 29640 20414
rect 28848 20293 29336 20299
rect 28848 20259 28860 20293
rect 29324 20259 29336 20293
rect 28848 20253 29336 20259
rect 28550 20180 28566 20200
rect 28560 19652 28566 20180
rect 27582 19624 27596 19652
rect 27024 19571 27084 19578
rect 26812 19565 27300 19571
rect 26812 19531 26824 19565
rect 27288 19531 27300 19565
rect 26812 19525 27300 19531
rect 26512 19100 26518 19160
rect 26578 19100 26584 19160
rect 27024 19043 27084 19525
rect 27536 19466 27596 19624
rect 28550 19624 28566 19652
rect 28600 20180 28610 20200
rect 29574 20200 29634 20354
rect 30074 20299 30134 20781
rect 30588 20722 30648 20880
rect 31614 20880 31620 21432
rect 31654 21432 31666 21456
rect 32626 21456 32686 21614
rect 33140 21555 33200 21614
rect 32920 21549 33408 21555
rect 32920 21515 32932 21549
rect 33396 21515 33408 21549
rect 32920 21509 33408 21515
rect 31654 20880 31660 21432
rect 32626 21420 32638 21456
rect 32632 20908 32638 21420
rect 31614 20868 31660 20880
rect 32624 20880 32638 20908
rect 32672 21420 32686 21456
rect 33642 21456 33702 21614
rect 33642 21432 33656 21456
rect 32672 20908 32678 21420
rect 32672 20880 32684 20908
rect 32104 20827 32164 20833
rect 30884 20821 31372 20827
rect 30884 20787 30896 20821
rect 31360 20787 31372 20821
rect 30884 20781 31372 20787
rect 31902 20821 32390 20827
rect 31902 20787 31914 20821
rect 32378 20787 32390 20821
rect 31902 20781 32390 20787
rect 30582 20662 30588 20722
rect 30648 20662 30654 20722
rect 31098 20299 31158 20781
rect 31602 20354 31608 20414
rect 31668 20354 31674 20414
rect 29866 20293 30354 20299
rect 29866 20259 29878 20293
rect 30342 20259 30354 20293
rect 29866 20253 30354 20259
rect 30884 20293 31372 20299
rect 30884 20259 30896 20293
rect 31360 20259 31372 20293
rect 30884 20253 31372 20259
rect 28600 19652 28606 20180
rect 29574 20172 29584 20200
rect 28600 19624 28610 19652
rect 27830 19565 28318 19571
rect 27830 19531 27842 19565
rect 28306 19531 28318 19565
rect 27830 19525 28318 19531
rect 28054 19468 28114 19525
rect 28550 19468 28610 19624
rect 29578 19624 29584 20172
rect 29618 20172 29634 20200
rect 30596 20200 30642 20212
rect 29618 19624 29624 20172
rect 30596 19660 30602 20200
rect 29578 19612 29624 19624
rect 30586 19624 30602 19660
rect 30636 19660 30642 20200
rect 31608 20200 31668 20354
rect 32104 20299 32164 20781
rect 32624 20722 32684 20880
rect 33650 20880 33656 21432
rect 33690 21432 33702 21456
rect 33690 20880 33696 21432
rect 33650 20868 33696 20880
rect 32920 20821 33408 20827
rect 32920 20787 32932 20821
rect 33396 20787 33408 20821
rect 32920 20781 33408 20787
rect 32618 20662 32624 20722
rect 32684 20662 32690 20722
rect 32626 20360 33702 20420
rect 31902 20293 32390 20299
rect 31902 20259 31914 20293
rect 32378 20259 32390 20293
rect 31902 20253 32390 20259
rect 31608 20176 31620 20200
rect 30636 19624 30646 19660
rect 31614 19652 31620 20176
rect 30068 19571 30128 19572
rect 28848 19565 29336 19571
rect 28848 19531 28860 19565
rect 29324 19531 29336 19565
rect 28848 19525 29336 19531
rect 29866 19565 30354 19571
rect 29866 19531 29878 19565
rect 30342 19531 30354 19565
rect 29866 19525 30354 19531
rect 29066 19468 29126 19525
rect 27530 19406 27536 19466
rect 27596 19406 27602 19466
rect 28054 19408 29126 19468
rect 27528 19100 27534 19160
rect 27594 19100 27600 19160
rect 25794 19037 26282 19043
rect 25794 19003 25806 19037
rect 26270 19003 26282 19037
rect 25794 18997 26282 19003
rect 26812 19037 27300 19043
rect 26812 19003 26824 19037
rect 27288 19003 27300 19037
rect 26812 18997 27300 19003
rect 25500 18922 25512 18944
rect 24528 18398 24534 18920
rect 24528 18368 24542 18398
rect 23758 18309 24246 18315
rect 23758 18275 23770 18309
rect 24234 18275 24246 18309
rect 23758 18269 24246 18275
rect 23976 18218 24036 18269
rect 22440 18158 22446 18218
rect 22506 18158 22512 18218
rect 22964 18158 24036 18218
rect 24242 18158 24248 18218
rect 24308 18158 24314 18218
rect 24482 18212 24542 18368
rect 25506 18368 25512 18922
rect 25546 18922 25560 18944
rect 26524 18944 26570 18956
rect 25546 18368 25552 18922
rect 26524 18394 26530 18944
rect 25506 18356 25552 18368
rect 26518 18368 26530 18394
rect 26564 18394 26570 18944
rect 27534 18944 27594 19100
rect 27830 19037 28318 19043
rect 27830 19003 27842 19037
rect 28306 19003 28318 19037
rect 27830 18997 28318 19003
rect 27534 18918 27548 18944
rect 26564 18368 26578 18394
rect 24776 18309 25264 18315
rect 24776 18275 24788 18309
rect 25252 18275 25264 18309
rect 24776 18269 25264 18275
rect 25794 18309 26282 18315
rect 25794 18275 25806 18309
rect 26270 18275 26282 18309
rect 25794 18269 26282 18275
rect 21928 17992 22704 18052
rect 21928 17787 21988 17992
rect 22434 17840 22440 17900
rect 22500 17840 22506 17900
rect 22644 17888 22704 17992
rect 20704 17781 21192 17787
rect 20704 17747 20716 17781
rect 21180 17747 21192 17781
rect 20704 17741 21192 17747
rect 21722 17781 22210 17787
rect 21722 17747 21734 17781
rect 22198 17747 22210 17781
rect 21722 17741 22210 17747
rect 20406 17662 20422 17688
rect 19438 17138 19444 17662
rect 19438 17112 19448 17138
rect 18668 17053 19156 17059
rect 18668 17019 18680 17053
rect 19144 17019 19156 17053
rect 18668 17013 19156 17019
rect 19388 16952 19448 17112
rect 20416 17112 20422 17662
rect 20456 17662 20466 17688
rect 21434 17688 21480 17700
rect 20456 17112 20462 17662
rect 21434 17134 21440 17688
rect 20416 17100 20462 17112
rect 21424 17112 21440 17134
rect 21474 17134 21480 17688
rect 22440 17688 22500 17840
rect 22638 17828 22644 17888
rect 22704 17828 22710 17888
rect 22740 17781 23228 17787
rect 22740 17747 22752 17781
rect 23216 17747 23228 17781
rect 22740 17741 23228 17747
rect 22440 17658 22458 17688
rect 22452 17148 22458 17658
rect 21474 17112 21484 17134
rect 19686 17053 20174 17059
rect 19686 17019 19698 17053
rect 20162 17019 20174 17053
rect 19686 17013 20174 17019
rect 20704 17053 21192 17059
rect 20704 17019 20716 17053
rect 21180 17019 21192 17053
rect 20704 17013 21192 17019
rect 19382 16892 19388 16952
rect 19448 16892 19454 16952
rect 19896 16838 19956 17013
rect 20920 16838 20980 17013
rect 21424 16952 21484 17112
rect 22446 17112 22458 17148
rect 22492 17658 22500 17688
rect 23460 17688 23520 18158
rect 24248 17948 24308 18158
rect 24476 18152 24482 18212
rect 24542 18152 24548 18212
rect 24978 18090 25038 18269
rect 26006 18090 26066 18269
rect 26518 18212 26578 18368
rect 27542 18368 27548 18918
rect 27582 18918 27594 18944
rect 28550 18944 28610 19408
rect 29564 19302 29570 19362
rect 29630 19302 29636 19362
rect 28848 19037 29336 19043
rect 28848 19003 28860 19037
rect 29324 19003 29336 19037
rect 28848 18997 29336 19003
rect 27582 18368 27588 18918
rect 28550 18914 28566 18944
rect 28560 18400 28566 18914
rect 27542 18356 27588 18368
rect 28548 18368 28566 18400
rect 28600 18914 28610 18944
rect 29570 18944 29630 19302
rect 30068 19043 30128 19525
rect 30432 19420 30438 19480
rect 30498 19420 30504 19480
rect 30438 19160 30498 19420
rect 30586 19370 30646 19624
rect 31606 19624 31620 19652
rect 31654 20176 31668 20200
rect 32626 20200 32686 20360
rect 33140 20299 33200 20360
rect 32920 20293 33408 20299
rect 32920 20259 32932 20293
rect 33396 20259 33408 20293
rect 32920 20253 33408 20259
rect 31654 19652 31660 20176
rect 32626 20166 32638 20200
rect 32632 19664 32638 20166
rect 31654 19624 31666 19652
rect 31092 19571 31152 19572
rect 30884 19565 31372 19571
rect 30884 19531 30896 19565
rect 31360 19531 31372 19565
rect 30884 19525 31372 19531
rect 30580 19310 30586 19370
rect 30646 19310 30652 19370
rect 30432 19100 30438 19160
rect 30498 19100 30504 19160
rect 30584 19102 30590 19162
rect 30650 19102 30656 19162
rect 29866 19037 30354 19043
rect 29866 19003 29878 19037
rect 30342 19003 30354 19037
rect 29866 18997 30354 19003
rect 28600 18400 28606 18914
rect 29570 18912 29584 18944
rect 29578 18400 29584 18912
rect 28600 18368 28608 18400
rect 26812 18309 27300 18315
rect 26812 18275 26824 18309
rect 27288 18275 27300 18309
rect 26812 18269 27300 18275
rect 27830 18309 28318 18315
rect 27830 18275 27842 18309
rect 28306 18275 28318 18309
rect 27830 18269 28318 18275
rect 26512 18152 26518 18212
rect 26578 18152 26584 18212
rect 24978 18030 26066 18090
rect 26510 18042 26516 18102
rect 26576 18042 26582 18102
rect 24248 17888 25556 17948
rect 23758 17781 24246 17787
rect 23758 17747 23770 17781
rect 24234 17747 24246 17781
rect 23758 17741 24246 17747
rect 24776 17781 25264 17787
rect 24776 17747 24788 17781
rect 25252 17747 25264 17781
rect 24776 17741 25264 17747
rect 22492 17148 22498 17658
rect 23460 17630 23476 17688
rect 22492 17112 22506 17148
rect 23470 17144 23476 17630
rect 21722 17053 22210 17059
rect 21722 17019 21734 17053
rect 22198 17019 22210 17053
rect 21722 17013 22210 17019
rect 21418 16892 21424 16952
rect 21484 16892 21490 16952
rect 21926 16838 21986 17013
rect 18086 16762 18092 16822
rect 18152 16762 18158 16822
rect 19896 16778 21986 16838
rect 13244 16634 13248 16694
rect 13308 16634 17770 16694
rect 13248 16628 13308 16634
rect 13128 16576 13188 16582
rect 18092 16576 18152 16762
rect 13188 16516 18152 16576
rect 13128 16510 13188 16516
rect 12682 16458 12742 16464
rect 19896 16458 19956 16778
rect 21926 16568 21986 16778
rect 22446 16682 22506 17112
rect 23460 17112 23476 17144
rect 23510 17630 23520 17688
rect 24488 17688 24534 17700
rect 23510 17144 23516 17630
rect 24488 17156 24494 17688
rect 23510 17112 23520 17144
rect 22740 17053 23228 17059
rect 22740 17019 22752 17053
rect 23216 17019 23228 17053
rect 22740 17013 23228 17019
rect 22964 16958 23024 17013
rect 23460 16958 23520 17112
rect 24482 17112 24494 17156
rect 24528 17156 24534 17688
rect 25496 17688 25556 17888
rect 26006 17888 26066 18030
rect 26006 17787 26066 17828
rect 25794 17781 26282 17787
rect 25794 17747 25806 17781
rect 26270 17747 26282 17781
rect 25794 17741 26282 17747
rect 25496 17636 25512 17688
rect 24528 17112 24542 17156
rect 23758 17053 24246 17059
rect 23758 17019 23770 17053
rect 24234 17019 24246 17053
rect 23758 17013 24246 17019
rect 23976 16958 24036 17013
rect 24482 16958 24542 17112
rect 25506 17112 25512 17636
rect 25546 17636 25556 17688
rect 26516 17688 26576 18042
rect 27022 17888 27082 18269
rect 28052 18216 28112 18269
rect 28548 18216 28608 18368
rect 29572 18368 29584 18400
rect 29618 18912 29630 18944
rect 30590 18944 30650 19102
rect 31092 19043 31152 19525
rect 31606 19260 31666 19624
rect 32626 19624 32638 19664
rect 32672 20166 32686 20200
rect 33642 20200 33702 20360
rect 33642 20178 33656 20200
rect 32672 19664 32678 20166
rect 32672 19624 32686 19664
rect 32098 19571 32158 19578
rect 31902 19565 32390 19571
rect 31902 19531 31914 19565
rect 32378 19531 32390 19565
rect 31902 19525 32390 19531
rect 31600 19200 31606 19260
rect 31666 19200 31672 19260
rect 32098 19043 32158 19525
rect 32626 19370 32686 19624
rect 33650 19624 33656 20178
rect 33690 20178 33702 20200
rect 33690 19624 33696 20178
rect 33650 19612 33696 19624
rect 32920 19565 33408 19571
rect 32920 19531 32932 19565
rect 33396 19531 33408 19565
rect 32920 19525 33408 19531
rect 33766 19370 33826 22138
rect 33908 21970 33968 24686
rect 34196 22270 34202 22330
rect 34262 22270 34268 22330
rect 33908 21904 33968 21910
rect 34044 21610 34050 21670
rect 34110 21610 34116 21670
rect 33884 20468 33890 20528
rect 33950 20468 33956 20528
rect 32620 19310 32626 19370
rect 32686 19310 32692 19370
rect 33760 19310 33766 19370
rect 33826 19310 33832 19370
rect 32618 19102 32624 19162
rect 32684 19102 32690 19162
rect 30884 19037 31372 19043
rect 30884 19003 30896 19037
rect 31360 19003 31372 19037
rect 30884 18997 31372 19003
rect 31902 19037 32390 19043
rect 31902 19003 31914 19037
rect 32378 19003 32390 19037
rect 31902 18997 32390 19003
rect 30590 18924 30602 18944
rect 29618 18400 29624 18912
rect 29618 18368 29632 18400
rect 28848 18309 29336 18315
rect 28848 18275 28860 18309
rect 29324 18275 29336 18309
rect 28848 18269 29336 18275
rect 29064 18216 29124 18269
rect 28052 18156 29124 18216
rect 29572 18214 29632 18368
rect 30596 18368 30602 18924
rect 30636 18924 30650 18944
rect 31614 18944 31660 18956
rect 30636 18368 30642 18924
rect 31614 18396 31620 18944
rect 30596 18356 30642 18368
rect 31608 18368 31620 18396
rect 31654 18396 31660 18944
rect 32624 18944 32684 19102
rect 32920 19037 33408 19043
rect 32920 19003 32932 19037
rect 33396 19003 33408 19037
rect 32920 18997 33408 19003
rect 32624 18920 32638 18944
rect 32632 18404 32638 18920
rect 31654 18368 31668 18396
rect 30080 18315 30140 18322
rect 31104 18315 31164 18322
rect 29866 18309 30354 18315
rect 29866 18275 29878 18309
rect 30342 18275 30354 18309
rect 29866 18269 30354 18275
rect 30884 18309 31372 18315
rect 30884 18275 30896 18309
rect 31360 18275 31372 18309
rect 30884 18269 31372 18275
rect 27022 17822 27082 17828
rect 26812 17781 27300 17787
rect 26812 17747 26824 17781
rect 27288 17747 27300 17781
rect 26812 17741 27300 17747
rect 27830 17781 28318 17787
rect 27830 17747 27842 17781
rect 28306 17747 28318 17781
rect 27830 17741 28318 17747
rect 25546 17112 25552 17636
rect 26516 17624 26530 17688
rect 25506 17100 25552 17112
rect 26524 17112 26530 17624
rect 26564 17624 26576 17688
rect 27542 17688 27588 17700
rect 26564 17112 26570 17624
rect 27542 17140 27548 17688
rect 26524 17100 26570 17112
rect 27534 17112 27548 17140
rect 27582 17140 27588 17688
rect 28548 17688 28608 18156
rect 29566 18154 29572 18214
rect 29632 18154 29638 18214
rect 30080 17894 30140 18269
rect 30080 17888 30142 17894
rect 30080 17828 30082 17888
rect 30588 17840 30594 17900
rect 30654 17840 30660 17900
rect 30080 17822 30142 17828
rect 30080 17787 30140 17822
rect 28848 17781 29336 17787
rect 28848 17747 28860 17781
rect 29324 17747 29336 17781
rect 28848 17741 29336 17747
rect 29866 17781 30354 17787
rect 29866 17747 29878 17781
rect 30342 17747 30354 17781
rect 29866 17741 30354 17747
rect 28548 17650 28566 17688
rect 28560 17142 28566 17650
rect 27582 17112 27594 17140
rect 24776 17053 25264 17059
rect 24776 17019 24788 17053
rect 25252 17019 25264 17053
rect 24776 17013 25264 17019
rect 25794 17053 26282 17059
rect 25794 17019 25806 17053
rect 26270 17019 26282 17053
rect 25794 17013 26282 17019
rect 26812 17053 27300 17059
rect 26812 17019 26824 17053
rect 27288 17019 27300 17053
rect 26812 17013 27300 17019
rect 24992 16958 25052 17013
rect 27018 16958 27078 17013
rect 27534 16958 27594 17112
rect 28548 17112 28566 17142
rect 28600 17650 28608 17688
rect 29578 17688 29624 17700
rect 28600 17142 28606 17650
rect 28600 17112 28608 17142
rect 29578 17138 29584 17688
rect 27830 17053 28318 17059
rect 27830 17019 27842 17053
rect 28306 17019 28318 17053
rect 27830 17013 28318 17019
rect 28052 16958 28112 17013
rect 28548 16958 28608 17112
rect 29576 17112 29584 17138
rect 29618 17138 29624 17688
rect 30594 17688 30654 17840
rect 31104 17787 31164 18269
rect 31608 18214 31668 18368
rect 32624 18368 32638 18404
rect 32672 18920 32684 18944
rect 33650 18944 33696 18956
rect 32672 18404 32678 18920
rect 32672 18368 32684 18404
rect 33650 18392 33656 18944
rect 32110 18315 32170 18328
rect 31902 18309 32390 18315
rect 31902 18275 31914 18309
rect 32378 18275 32390 18309
rect 31902 18269 32390 18275
rect 31602 18154 31608 18214
rect 31668 18154 31674 18214
rect 32110 17787 32170 18269
rect 32624 18210 32684 18368
rect 33640 18368 33656 18392
rect 33690 18392 33696 18944
rect 33690 18368 33700 18392
rect 32920 18309 33408 18315
rect 32920 18275 32932 18309
rect 33396 18275 33408 18309
rect 32920 18269 33408 18275
rect 33138 18210 33198 18269
rect 33640 18210 33700 18368
rect 32624 18150 33700 18210
rect 33766 18102 33826 19310
rect 33890 19162 33950 20468
rect 33884 19102 33890 19162
rect 33950 19102 33956 19162
rect 33760 18042 33766 18102
rect 33826 18042 33832 18102
rect 32622 17840 32628 17900
rect 32688 17840 32694 17900
rect 30884 17781 31372 17787
rect 30884 17747 30896 17781
rect 31360 17747 31372 17781
rect 30884 17741 31372 17747
rect 31902 17781 32390 17787
rect 31902 17747 31914 17781
rect 32378 17747 32390 17781
rect 31902 17741 32390 17747
rect 30594 17662 30602 17688
rect 29618 17112 29636 17138
rect 28848 17053 29336 17059
rect 28848 17019 28860 17053
rect 29324 17019 29336 17053
rect 28848 17013 29336 17019
rect 29064 16958 29124 17013
rect 22964 16898 29124 16958
rect 29576 16952 29636 17112
rect 30596 17112 30602 17662
rect 30636 17662 30654 17688
rect 31614 17688 31660 17700
rect 30636 17112 30642 17662
rect 31614 17134 31620 17688
rect 30596 17100 30642 17112
rect 31612 17112 31620 17134
rect 31654 17134 31660 17688
rect 32628 17688 32688 17840
rect 32920 17781 33408 17787
rect 32920 17747 32932 17781
rect 33396 17747 33408 17781
rect 32920 17741 33408 17747
rect 32628 17658 32638 17688
rect 32632 17150 32638 17658
rect 31654 17112 31672 17134
rect 30084 17059 30144 17066
rect 29866 17053 30354 17059
rect 29866 17019 29878 17053
rect 30342 17019 30354 17053
rect 29866 17013 30354 17019
rect 30884 17053 31372 17059
rect 30884 17019 30896 17053
rect 31360 17019 31372 17053
rect 30884 17013 31372 17019
rect 29570 16892 29576 16952
rect 29636 16892 29642 16952
rect 30084 16840 30144 17013
rect 31104 16840 31164 17013
rect 31612 16952 31672 17112
rect 32626 17112 32638 17150
rect 32672 17658 32688 17688
rect 33650 17688 33696 17700
rect 32672 17150 32678 17658
rect 32672 17112 32686 17150
rect 33650 17138 33656 17688
rect 31902 17053 32390 17059
rect 31902 17019 31914 17053
rect 32378 17019 32390 17053
rect 31902 17013 32390 17019
rect 31606 16892 31612 16952
rect 31672 16892 31678 16952
rect 32106 16840 32166 17013
rect 32626 16956 32686 17112
rect 33642 17112 33656 17138
rect 33690 17138 33696 17688
rect 33690 17112 33702 17138
rect 32920 17053 33408 17059
rect 32920 17019 32932 17053
rect 33396 17019 33408 17053
rect 32920 17013 33408 17019
rect 33140 16956 33200 17013
rect 33642 16956 33702 17112
rect 32626 16896 33702 16956
rect 30084 16780 32166 16840
rect 22440 16622 22446 16682
rect 22506 16622 22512 16682
rect 30084 16568 30144 16780
rect 34050 16682 34110 21610
rect 34202 20414 34262 22270
rect 34196 20354 34202 20414
rect 34262 20354 34268 20414
rect 35628 16812 35634 30242
rect 35734 16812 35740 30242
rect 34044 16622 34050 16682
rect 34110 16622 34116 16682
rect 21926 16508 30144 16568
rect 12742 16398 19956 16458
rect 12682 16392 12742 16398
rect 35628 16298 35740 16812
rect 11284 16292 35740 16298
rect 11284 16192 11390 16292
rect 35634 16192 35740 16292
rect 11284 16186 35740 16192
rect 8046 15870 8190 16162
rect -7870 15807 -7070 15838
rect -7870 15773 -7767 15807
rect -7733 15773 -7675 15807
rect -7641 15773 -7583 15807
rect -7549 15773 -7317 15807
rect -7283 15773 -7225 15807
rect -7191 15773 -7133 15807
rect -7099 15773 -7070 15807
rect -7870 15742 -7070 15773
rect -7870 15638 -7858 15742
rect -7918 15590 -7858 15638
rect -8164 15578 -7858 15590
rect -8164 15544 -8142 15578
rect -7940 15544 -7858 15578
rect -8164 15530 -7858 15544
rect -3080 15562 8190 15870
rect -7425 15512 -7365 15518
rect -7645 15506 -7425 15512
rect -7743 15490 -7683 15496
rect -7749 15430 -7743 15490
rect -7683 15430 -7677 15490
rect -7645 15466 -7633 15506
rect -7587 15466 -7425 15506
rect -7645 15452 -7425 15466
rect -7365 15506 -7228 15512
rect -7365 15458 -7288 15506
rect -7240 15458 -7228 15506
rect -7365 15452 -7228 15458
rect -7196 15510 -7030 15516
rect -7196 15462 -7184 15510
rect -7136 15462 -7030 15510
rect -7196 15456 -7030 15462
rect -7425 15446 -7365 15452
rect -7743 15424 -7683 15430
rect -8442 15274 -8334 15280
rect -8442 15240 -8430 15274
rect -8346 15240 -8334 15274
rect -8442 15234 -8334 15240
rect -8758 15014 -8752 15034
rect -8798 15002 -8752 15014
rect -8546 15014 -8534 15190
rect -8500 15014 -8486 15190
rect -8288 15190 -8228 15353
rect -8158 15380 -7856 15390
rect -8158 15342 -8138 15380
rect -7940 15342 -7856 15380
rect -8158 15330 -7856 15342
rect -8158 15280 -8098 15330
rect -8184 15274 -8076 15280
rect -8184 15240 -8172 15274
rect -8088 15240 -8076 15274
rect -8184 15234 -8076 15240
rect -8288 15151 -8276 15190
rect -8546 14974 -8486 15014
rect -8282 15014 -8276 15151
rect -8242 15151 -8228 15190
rect -8030 15190 -7970 15330
rect -8242 15014 -8236 15151
rect -8030 15144 -8018 15190
rect -8024 15047 -8018 15144
rect -8282 15002 -8236 15014
rect -8032 15014 -8018 15047
rect -7984 15144 -7970 15190
rect -7916 15294 -7856 15330
rect -3080 15368 9272 15562
rect -3080 15362 35840 15368
rect -7916 15280 -7070 15294
rect -7984 15047 -7978 15144
rect -7984 15014 -7972 15047
rect -9474 14964 -9366 14970
rect -9474 14930 -9462 14964
rect -9378 14930 -9366 14964
rect -9474 14924 -9366 14930
rect -9216 14964 -9108 14970
rect -9216 14930 -9204 14964
rect -9120 14930 -9108 14964
rect -9216 14924 -9108 14930
rect -8958 14964 -8850 14970
rect -8958 14930 -8946 14964
rect -8862 14930 -8850 14964
rect -8958 14924 -8850 14930
rect -8700 14964 -8592 14970
rect -8700 14930 -8688 14964
rect -8604 14930 -8592 14964
rect -8700 14924 -8592 14930
rect -8442 14964 -8334 14970
rect -8442 14930 -8430 14964
rect -8346 14930 -8334 14964
rect -8442 14924 -8334 14930
rect -8184 14964 -8076 14970
rect -8184 14930 -8172 14964
rect -8088 14930 -8076 14964
rect -8184 14924 -8076 14930
rect -9450 14875 -9390 14924
rect -9694 14864 -9390 14875
rect -9694 14828 -9612 14864
rect -9404 14828 -9390 14864
rect -9694 14740 -9390 14828
rect -9192 14865 -9132 14924
rect -8932 14865 -8872 14924
rect -8674 14865 -8614 14924
rect -8418 14865 -8358 14924
rect -8160 14875 -8100 14924
rect -8032 14875 -7972 15014
rect -7916 14924 -7906 15280
rect -7868 15263 -7070 15280
rect -7868 15229 -7767 15263
rect -7733 15229 -7675 15263
rect -7641 15229 -7583 15263
rect -7549 15229 -7317 15263
rect -7283 15229 -7225 15263
rect -7191 15229 -7133 15263
rect -7099 15229 -7070 15263
rect -3080 15262 -1310 15362
rect 35734 15262 35840 15362
rect -3080 15256 35840 15262
rect -3080 15240 9270 15256
rect -7868 15198 -7070 15229
rect -7868 14924 -7856 15198
rect -7916 14875 -7856 14924
rect -9192 14805 -8418 14865
rect -8358 14805 -8352 14865
rect -8160 14862 -7856 14875
rect -8160 14826 -8140 14862
rect -7938 14826 -7856 14862
rect -8160 14740 -7856 14826
rect -1416 14740 -1304 15240
rect 12800 15182 12860 15188
rect 13122 15132 13128 15192
rect 13188 15132 13194 15192
rect 13248 15184 13308 15190
rect 12188 14986 12194 15046
rect 12254 14986 12260 15046
rect 12308 14988 12314 15048
rect 12374 14988 12380 15048
rect 12448 15006 12454 15066
rect 12514 15006 12520 15066
rect 12676 15022 12682 15082
rect 12742 15022 12748 15082
rect 12056 14858 12062 14918
rect 12122 14858 12128 14918
rect -12293 14680 -1304 14740
rect -1416 14470 -1304 14680
rect -1416 210 -1410 14470
rect -1310 210 -1304 14470
rect 9344 14260 9350 14320
rect 9410 14260 9416 14320
rect 9350 14216 9410 14260
rect 1716 14156 9410 14216
rect 1716 14016 1776 14156
rect 2226 14106 2286 14156
rect 2010 14100 2498 14106
rect 2010 14066 2022 14100
rect 2486 14066 2498 14100
rect 2010 14060 2498 14066
rect 1716 13986 1728 14016
rect 1722 13458 1728 13986
rect 1712 13440 1728 13458
rect 1762 13986 1776 14016
rect 2732 14016 2792 14156
rect 3234 14106 3294 14156
rect 4262 14106 4322 14156
rect 3028 14100 3516 14106
rect 3028 14066 3040 14100
rect 3504 14066 3516 14100
rect 3028 14060 3516 14066
rect 4046 14100 4534 14106
rect 4046 14066 4058 14100
rect 4522 14066 4534 14100
rect 4046 14060 4534 14066
rect 2732 13992 2746 14016
rect 1762 13458 1768 13986
rect 2740 13462 2746 13992
rect 1762 13440 1772 13458
rect 1712 13198 1772 13440
rect 2732 13440 2746 13462
rect 2780 13992 2792 14016
rect 3758 14016 3804 14028
rect 2780 13462 2786 13992
rect 3758 13464 3764 14016
rect 2780 13440 2792 13462
rect 2010 13390 2498 13396
rect 2010 13356 2022 13390
rect 2486 13356 2498 13390
rect 2010 13350 2498 13356
rect 2226 13288 2286 13350
rect 2010 13282 2498 13288
rect 2010 13248 2022 13282
rect 2486 13248 2498 13282
rect 2010 13242 2498 13248
rect 1712 13168 1728 13198
rect 1722 12644 1728 13168
rect 1714 12622 1728 12644
rect 1762 13168 1772 13198
rect 2732 13198 2792 13440
rect 3752 13440 3764 13464
rect 3798 13464 3804 14016
rect 4770 14016 4830 14156
rect 5276 14106 5336 14156
rect 6290 14106 6350 14156
rect 5064 14100 5552 14106
rect 5064 14066 5076 14100
rect 5540 14066 5552 14100
rect 5064 14060 5552 14066
rect 6082 14100 6570 14106
rect 6082 14066 6094 14100
rect 6558 14066 6570 14100
rect 6082 14060 6570 14066
rect 4770 13978 4782 14016
rect 3798 13440 3812 13464
rect 4776 13460 4782 13978
rect 3028 13390 3516 13396
rect 3028 13356 3040 13390
rect 3504 13356 3516 13390
rect 3028 13350 3516 13356
rect 3230 13288 3290 13350
rect 3028 13282 3516 13288
rect 3028 13248 3040 13282
rect 3504 13248 3516 13282
rect 3028 13242 3516 13248
rect 2732 13172 2746 13198
rect 1762 12644 1768 13168
rect 2740 12648 2746 13172
rect 1762 12622 1774 12644
rect 1714 12380 1774 12622
rect 2734 12622 2746 12648
rect 2780 13172 2792 13198
rect 3752 13198 3812 13440
rect 4770 13440 4782 13460
rect 4816 13978 4830 14016
rect 5794 14016 5840 14028
rect 6806 14016 6866 14156
rect 7322 14106 7382 14156
rect 8328 14106 8388 14156
rect 7100 14100 7588 14106
rect 7100 14066 7112 14100
rect 7576 14066 7588 14100
rect 7100 14060 7588 14066
rect 8118 14100 8606 14106
rect 8118 14066 8130 14100
rect 8594 14066 8606 14100
rect 8118 14060 8606 14066
rect 4816 13460 4822 13978
rect 5794 13468 5800 14016
rect 4816 13440 4830 13460
rect 4046 13390 4534 13396
rect 4046 13356 4058 13390
rect 4522 13356 4534 13390
rect 4046 13350 4534 13356
rect 4260 13288 4320 13350
rect 4046 13282 4534 13288
rect 4046 13248 4058 13282
rect 4522 13248 4534 13282
rect 4046 13242 4534 13248
rect 3752 13174 3764 13198
rect 2780 12648 2786 13172
rect 3758 12650 3764 13174
rect 2780 12622 2794 12648
rect 2010 12572 2498 12578
rect 2010 12538 2022 12572
rect 2486 12538 2498 12572
rect 2010 12532 2498 12538
rect 2226 12470 2286 12532
rect 2010 12464 2498 12470
rect 2010 12430 2022 12464
rect 2486 12430 2498 12464
rect 2010 12424 2498 12430
rect 1714 12354 1728 12380
rect 1722 11816 1728 12354
rect 1714 11804 1728 11816
rect 1762 12354 1774 12380
rect 2734 12380 2794 12622
rect 3754 12622 3764 12650
rect 3798 13174 3812 13198
rect 4770 13198 4830 13440
rect 5790 13440 5800 13468
rect 5834 13468 5840 14016
rect 6804 13982 6818 14016
rect 6806 13970 6818 13982
rect 5834 13440 5850 13468
rect 6812 13460 6818 13970
rect 5064 13390 5552 13396
rect 5064 13356 5076 13390
rect 5540 13356 5552 13390
rect 5064 13350 5552 13356
rect 5262 13288 5322 13350
rect 5064 13282 5552 13288
rect 5064 13248 5076 13282
rect 5540 13248 5552 13282
rect 5064 13242 5552 13248
rect 3798 12650 3804 13174
rect 4770 13170 4782 13198
rect 3798 12622 3814 12650
rect 4776 12646 4782 13170
rect 3028 12572 3516 12578
rect 3028 12538 3040 12572
rect 3504 12538 3516 12572
rect 3028 12532 3516 12538
rect 3242 12470 3302 12532
rect 3028 12464 3516 12470
rect 3028 12430 3040 12464
rect 3504 12430 3516 12464
rect 3028 12424 3516 12430
rect 2734 12358 2746 12380
rect 1762 11816 1768 12354
rect 2740 11820 2746 12358
rect 1762 11804 1774 11816
rect 1714 11562 1774 11804
rect 2734 11804 2746 11820
rect 2780 12358 2794 12380
rect 3754 12380 3814 12622
rect 4772 12622 4782 12646
rect 4816 13170 4830 13198
rect 5790 13198 5850 13440
rect 6802 13440 6818 13460
rect 6852 13970 6866 14016
rect 7830 14016 7876 14028
rect 6852 13460 6858 13970
rect 7830 13460 7836 14016
rect 6852 13440 6862 13460
rect 6082 13390 6570 13396
rect 6082 13356 6094 13390
rect 6558 13356 6570 13390
rect 6082 13350 6570 13356
rect 6292 13288 6352 13350
rect 6082 13282 6570 13288
rect 6082 13248 6094 13282
rect 6558 13248 6570 13282
rect 6082 13242 6570 13248
rect 5790 13178 5800 13198
rect 4816 12646 4822 13170
rect 5794 12654 5800 13178
rect 4816 12622 4832 12646
rect 4046 12572 4534 12578
rect 4046 12538 4058 12572
rect 4522 12538 4534 12572
rect 4046 12532 4534 12538
rect 4260 12470 4320 12532
rect 4046 12464 4534 12470
rect 4046 12430 4058 12464
rect 4522 12430 4534 12464
rect 4046 12424 4534 12430
rect 3754 12360 3764 12380
rect 2780 11820 2786 12358
rect 3758 11822 3764 12360
rect 2780 11804 2794 11820
rect 2010 11754 2498 11760
rect 2010 11720 2022 11754
rect 2486 11720 2498 11754
rect 2010 11714 2498 11720
rect 2220 11652 2280 11714
rect 2010 11646 2498 11652
rect 2010 11612 2022 11646
rect 2486 11612 2498 11646
rect 2010 11606 2498 11612
rect 1714 11526 1728 11562
rect 1722 11004 1728 11526
rect 1714 10986 1728 11004
rect 1762 11526 1774 11562
rect 2734 11562 2794 11804
rect 3754 11804 3764 11822
rect 3798 12360 3814 12380
rect 4772 12380 4832 12622
rect 5792 12622 5800 12654
rect 5834 13178 5850 13198
rect 6802 13198 6862 13440
rect 7824 13440 7836 13460
rect 7870 13460 7876 14016
rect 8840 14016 8900 14156
rect 9350 14106 9410 14156
rect 10870 14126 10876 14186
rect 10936 14126 10942 14186
rect 9136 14100 9624 14106
rect 9136 14066 9148 14100
rect 9612 14066 9624 14100
rect 9136 14060 9624 14066
rect 10154 14100 10642 14106
rect 10154 14066 10166 14100
rect 10630 14066 10642 14100
rect 10154 14060 10642 14066
rect 8840 13980 8854 14016
rect 8848 13460 8854 13980
rect 7870 13440 7884 13460
rect 7100 13390 7588 13396
rect 7100 13356 7112 13390
rect 7576 13356 7588 13390
rect 7100 13350 7588 13356
rect 7308 13288 7368 13350
rect 7100 13282 7588 13288
rect 7100 13248 7112 13282
rect 7576 13248 7588 13282
rect 7100 13242 7588 13248
rect 5834 12654 5840 13178
rect 6802 13170 6818 13198
rect 5834 12622 5852 12654
rect 6812 12646 6818 13170
rect 5064 12572 5552 12578
rect 5064 12538 5076 12572
rect 5540 12538 5552 12572
rect 5064 12532 5552 12538
rect 5262 12470 5322 12532
rect 5064 12464 5552 12470
rect 5064 12430 5076 12464
rect 5540 12430 5552 12464
rect 5064 12424 5552 12430
rect 3798 11822 3804 12360
rect 4772 12356 4782 12380
rect 3798 11804 3814 11822
rect 4776 11818 4782 12356
rect 3028 11754 3516 11760
rect 3028 11720 3040 11754
rect 3504 11720 3516 11754
rect 3028 11714 3516 11720
rect 3242 11652 3302 11714
rect 3028 11646 3516 11652
rect 3028 11612 3040 11646
rect 3504 11612 3516 11646
rect 3028 11606 3516 11612
rect 2734 11530 2746 11562
rect 1762 11004 1768 11526
rect 2740 11008 2746 11530
rect 1762 10986 1774 11004
rect 1714 10744 1774 10986
rect 2734 10986 2746 11008
rect 2780 11530 2794 11562
rect 3754 11562 3814 11804
rect 4772 11804 4782 11818
rect 4816 12356 4832 12380
rect 5792 12380 5852 12622
rect 6804 12622 6818 12646
rect 6852 13170 6862 13198
rect 7824 13198 7884 13440
rect 8844 13440 8854 13460
rect 8888 13980 8900 14016
rect 9866 14016 9912 14028
rect 8888 13460 8894 13980
rect 9866 13464 9872 14016
rect 8888 13440 8904 13460
rect 8118 13390 8606 13396
rect 8118 13356 8130 13390
rect 8594 13356 8606 13390
rect 8118 13350 8606 13356
rect 8330 13288 8390 13350
rect 8118 13282 8606 13288
rect 8118 13248 8130 13282
rect 8594 13248 8606 13282
rect 8118 13242 8606 13248
rect 7824 13170 7836 13198
rect 6852 12646 6858 13170
rect 7830 12646 7836 13170
rect 6852 12622 6864 12646
rect 6082 12572 6570 12578
rect 6082 12538 6094 12572
rect 6558 12538 6570 12572
rect 6082 12532 6570 12538
rect 6292 12470 6352 12532
rect 6082 12464 6570 12470
rect 6082 12430 6094 12464
rect 6558 12430 6570 12464
rect 6082 12424 6570 12430
rect 5792 12364 5800 12380
rect 4816 11818 4822 12356
rect 5794 11826 5800 12364
rect 4816 11804 4832 11818
rect 4046 11754 4534 11760
rect 4046 11720 4058 11754
rect 4522 11720 4534 11754
rect 4046 11714 4534 11720
rect 4254 11652 4314 11714
rect 4046 11646 4534 11652
rect 4046 11612 4058 11646
rect 4522 11612 4534 11646
rect 4046 11606 4534 11612
rect 3754 11532 3764 11562
rect 2780 11008 2786 11530
rect 3758 11010 3764 11532
rect 2780 10986 2794 11008
rect 2010 10936 2498 10942
rect 2010 10902 2022 10936
rect 2486 10902 2498 10936
rect 2010 10896 2498 10902
rect 2218 10834 2278 10896
rect 2010 10828 2498 10834
rect 2010 10794 2022 10828
rect 2486 10794 2498 10828
rect 2010 10788 2498 10794
rect 1714 10714 1728 10744
rect 1722 10184 1728 10714
rect 1714 10168 1728 10184
rect 1762 10714 1774 10744
rect 2734 10744 2794 10986
rect 3754 10986 3764 11010
rect 3798 11532 3814 11562
rect 4772 11562 4832 11804
rect 5792 11804 5800 11826
rect 5834 12364 5852 12380
rect 6804 12380 6864 12622
rect 7826 12622 7836 12646
rect 7870 13170 7884 13198
rect 8844 13198 8904 13440
rect 9860 13440 9872 13464
rect 9906 13464 9912 14016
rect 10876 14016 10936 14126
rect 10876 13980 10890 14016
rect 9906 13440 9920 13464
rect 10884 13460 10890 13980
rect 9136 13390 9624 13396
rect 9136 13356 9148 13390
rect 9612 13356 9624 13390
rect 9136 13350 9624 13356
rect 9342 13288 9402 13350
rect 9136 13282 9624 13288
rect 9136 13248 9148 13282
rect 9612 13248 9624 13282
rect 9136 13242 9624 13248
rect 8844 13170 8854 13198
rect 7870 12646 7876 13170
rect 8848 12646 8854 13170
rect 7870 12622 7886 12646
rect 7100 12572 7588 12578
rect 7100 12538 7112 12572
rect 7576 12538 7588 12572
rect 7100 12532 7588 12538
rect 7308 12470 7368 12532
rect 7100 12464 7588 12470
rect 7100 12430 7112 12464
rect 7576 12430 7588 12464
rect 7100 12424 7588 12430
rect 5834 11826 5840 12364
rect 6804 12356 6818 12380
rect 5834 11804 5852 11826
rect 6812 11818 6818 12356
rect 5064 11754 5552 11760
rect 5064 11720 5076 11754
rect 5540 11720 5552 11754
rect 5064 11714 5552 11720
rect 5256 11652 5316 11714
rect 5064 11646 5552 11652
rect 5064 11612 5076 11646
rect 5540 11612 5552 11646
rect 5064 11606 5552 11612
rect 3798 11010 3804 11532
rect 4772 11528 4782 11562
rect 3798 10986 3814 11010
rect 4776 11006 4782 11528
rect 3028 10936 3516 10942
rect 3028 10902 3040 10936
rect 3504 10902 3516 10936
rect 3028 10896 3516 10902
rect 3236 10834 3296 10896
rect 3028 10828 3516 10834
rect 3028 10794 3040 10828
rect 3504 10794 3516 10828
rect 3028 10788 3516 10794
rect 2734 10718 2746 10744
rect 1762 10184 1768 10714
rect 2740 10188 2746 10718
rect 1762 10168 1774 10184
rect 1714 9926 1774 10168
rect 2734 10168 2746 10188
rect 2780 10718 2794 10744
rect 3754 10744 3814 10986
rect 4772 10986 4782 11006
rect 4816 11528 4832 11562
rect 5792 11562 5852 11804
rect 6804 11804 6818 11818
rect 6852 12356 6864 12380
rect 7826 12380 7886 12622
rect 8846 12622 8854 12646
rect 8888 13170 8904 13198
rect 9860 13198 9920 13440
rect 10882 13440 10890 13460
rect 10924 13980 10936 14016
rect 10924 13460 10930 13980
rect 10924 13440 10942 13460
rect 10154 13390 10642 13396
rect 10154 13356 10166 13390
rect 10630 13356 10642 13390
rect 10154 13350 10642 13356
rect 10362 13288 10422 13350
rect 10154 13282 10642 13288
rect 10154 13248 10166 13282
rect 10630 13248 10642 13282
rect 10154 13242 10642 13248
rect 9860 13174 9872 13198
rect 8888 12646 8894 13170
rect 9866 12650 9872 13174
rect 8888 12622 8906 12646
rect 8118 12572 8606 12578
rect 8118 12538 8130 12572
rect 8594 12538 8606 12572
rect 8118 12532 8606 12538
rect 8330 12470 8390 12532
rect 8118 12464 8606 12470
rect 8118 12430 8130 12464
rect 8594 12430 8606 12464
rect 8118 12424 8606 12430
rect 7826 12356 7836 12380
rect 6852 11818 6858 12356
rect 7830 11818 7836 12356
rect 6852 11804 6864 11818
rect 6082 11754 6570 11760
rect 6082 11720 6094 11754
rect 6558 11720 6570 11754
rect 6082 11714 6570 11720
rect 6286 11652 6346 11714
rect 6082 11646 6570 11652
rect 6082 11612 6094 11646
rect 6558 11612 6570 11646
rect 6082 11606 6570 11612
rect 5792 11536 5800 11562
rect 4816 11006 4822 11528
rect 5794 11014 5800 11536
rect 4816 10986 4832 11006
rect 4046 10936 4534 10942
rect 4046 10902 4058 10936
rect 4522 10902 4534 10936
rect 4046 10896 4534 10902
rect 4252 10834 4312 10896
rect 4046 10828 4534 10834
rect 4046 10794 4058 10828
rect 4522 10794 4534 10828
rect 4046 10788 4534 10794
rect 3754 10720 3764 10744
rect 2780 10188 2786 10718
rect 3758 10190 3764 10720
rect 2780 10168 2794 10188
rect 2010 10118 2498 10124
rect 2010 10084 2022 10118
rect 2486 10084 2498 10118
rect 2010 10078 2498 10084
rect 2220 10016 2280 10078
rect 2010 10010 2498 10016
rect 2010 9976 2022 10010
rect 2486 9976 2498 10010
rect 2010 9970 2498 9976
rect 1714 9894 1728 9926
rect 1722 9372 1728 9894
rect 1714 9350 1728 9372
rect 1762 9894 1774 9926
rect 2734 9926 2794 10168
rect 3754 10168 3764 10190
rect 3798 10720 3814 10744
rect 4772 10744 4832 10986
rect 5792 10986 5800 11014
rect 5834 11536 5852 11562
rect 6804 11562 6864 11804
rect 7826 11804 7836 11818
rect 7870 12356 7886 12380
rect 8846 12380 8906 12622
rect 9862 12622 9872 12650
rect 9906 13174 9920 13198
rect 10882 13198 10942 13440
rect 9906 12650 9912 13174
rect 10882 13170 10890 13198
rect 9906 12622 9922 12650
rect 9136 12572 9624 12578
rect 9136 12538 9148 12572
rect 9612 12538 9624 12572
rect 9136 12532 9624 12538
rect 9342 12470 9402 12532
rect 9136 12464 9624 12470
rect 9136 12430 9148 12464
rect 9612 12430 9624 12464
rect 9136 12424 9624 12430
rect 8846 12356 8854 12380
rect 7870 11818 7876 12356
rect 8848 11818 8854 12356
rect 7870 11804 7886 11818
rect 7100 11754 7588 11760
rect 7100 11720 7112 11754
rect 7576 11720 7588 11754
rect 7100 11714 7588 11720
rect 7302 11652 7362 11714
rect 7100 11646 7588 11652
rect 7100 11612 7112 11646
rect 7576 11612 7588 11646
rect 7100 11606 7588 11612
rect 5834 11014 5840 11536
rect 6804 11528 6818 11562
rect 5834 10986 5852 11014
rect 6812 11006 6818 11528
rect 5064 10936 5552 10942
rect 5064 10902 5076 10936
rect 5540 10902 5552 10936
rect 5064 10896 5552 10902
rect 5254 10834 5314 10896
rect 5064 10828 5552 10834
rect 5064 10794 5076 10828
rect 5540 10794 5552 10828
rect 5064 10788 5552 10794
rect 3798 10190 3804 10720
rect 4772 10716 4782 10744
rect 3798 10168 3814 10190
rect 4776 10186 4782 10716
rect 3028 10118 3516 10124
rect 3028 10084 3040 10118
rect 3504 10084 3516 10118
rect 3028 10078 3516 10084
rect 3234 10016 3294 10078
rect 3028 10010 3516 10016
rect 3028 9976 3040 10010
rect 3504 9976 3516 10010
rect 3028 9970 3516 9976
rect 2734 9898 2746 9926
rect 1762 9372 1768 9894
rect 2740 9376 2746 9898
rect 1762 9350 1774 9372
rect 1714 9108 1774 9350
rect 2734 9350 2746 9376
rect 2780 9898 2794 9926
rect 3754 9926 3814 10168
rect 4772 10168 4782 10186
rect 4816 10716 4832 10744
rect 5792 10744 5852 10986
rect 6804 10986 6818 11006
rect 6852 11528 6864 11562
rect 7826 11562 7886 11804
rect 8846 11804 8854 11818
rect 8888 12356 8906 12380
rect 9862 12380 9922 12622
rect 10884 12622 10890 13170
rect 10924 13170 10942 13198
rect 10924 12646 10930 13170
rect 10924 12622 10944 12646
rect 10154 12572 10642 12578
rect 10154 12538 10166 12572
rect 10630 12538 10642 12572
rect 10154 12532 10642 12538
rect 10362 12470 10422 12532
rect 10154 12464 10642 12470
rect 10154 12430 10166 12464
rect 10630 12430 10642 12464
rect 10154 12424 10642 12430
rect 9862 12360 9872 12380
rect 8888 11818 8894 12356
rect 9866 11822 9872 12360
rect 8888 11804 8906 11818
rect 8118 11754 8606 11760
rect 8118 11720 8130 11754
rect 8594 11720 8606 11754
rect 8118 11714 8606 11720
rect 8324 11652 8384 11714
rect 8118 11646 8606 11652
rect 8118 11612 8130 11646
rect 8594 11612 8606 11646
rect 8118 11606 8606 11612
rect 7826 11528 7836 11562
rect 6852 11006 6858 11528
rect 7830 11006 7836 11528
rect 6852 10986 6864 11006
rect 6082 10936 6570 10942
rect 6082 10902 6094 10936
rect 6558 10902 6570 10936
rect 6082 10896 6570 10902
rect 6284 10834 6344 10896
rect 6082 10828 6570 10834
rect 6082 10794 6094 10828
rect 6558 10794 6570 10828
rect 6082 10788 6570 10794
rect 5792 10724 5800 10744
rect 4816 10186 4822 10716
rect 5794 10194 5800 10724
rect 4816 10168 4832 10186
rect 4046 10118 4534 10124
rect 4046 10084 4058 10118
rect 4522 10084 4534 10118
rect 4046 10078 4534 10084
rect 4254 10016 4314 10078
rect 4046 10010 4534 10016
rect 4046 9976 4058 10010
rect 4522 9976 4534 10010
rect 4046 9970 4534 9976
rect 3754 9900 3764 9926
rect 2780 9376 2786 9898
rect 3758 9378 3764 9900
rect 2780 9350 2794 9376
rect 2010 9300 2498 9306
rect 2010 9266 2022 9300
rect 2486 9266 2498 9300
rect 2010 9260 2498 9266
rect 2222 9198 2282 9260
rect 2010 9192 2498 9198
rect 2010 9158 2022 9192
rect 2486 9158 2498 9192
rect 2010 9152 2498 9158
rect 1714 9082 1728 9108
rect 1722 8554 1728 9082
rect 1714 8532 1728 8554
rect 1762 9082 1774 9108
rect 2734 9108 2794 9350
rect 3754 9350 3764 9378
rect 3798 9900 3814 9926
rect 4772 9926 4832 10168
rect 5792 10168 5800 10194
rect 5834 10724 5852 10744
rect 6804 10744 6864 10986
rect 7826 10986 7836 11006
rect 7870 11528 7886 11562
rect 8846 11562 8906 11804
rect 9862 11804 9872 11822
rect 9906 12360 9922 12380
rect 10884 12380 10944 12622
rect 9906 11822 9912 12360
rect 9906 11804 9922 11822
rect 9136 11754 9624 11760
rect 9136 11720 9148 11754
rect 9612 11720 9624 11754
rect 9136 11714 9624 11720
rect 9336 11652 9396 11714
rect 9136 11646 9624 11652
rect 9136 11612 9148 11646
rect 9612 11612 9624 11646
rect 9136 11606 9624 11612
rect 8846 11528 8854 11562
rect 7870 11006 7876 11528
rect 8848 11006 8854 11528
rect 7870 10986 7886 11006
rect 7100 10936 7588 10942
rect 7100 10902 7112 10936
rect 7576 10902 7588 10936
rect 7100 10896 7588 10902
rect 7300 10834 7360 10896
rect 7100 10828 7588 10834
rect 7100 10794 7112 10828
rect 7576 10794 7588 10828
rect 7100 10788 7588 10794
rect 5834 10194 5840 10724
rect 6804 10716 6818 10744
rect 5834 10168 5852 10194
rect 6812 10186 6818 10716
rect 5064 10118 5552 10124
rect 5064 10084 5076 10118
rect 5540 10084 5552 10118
rect 5064 10078 5552 10084
rect 5256 10016 5316 10078
rect 5064 10010 5552 10016
rect 5064 9976 5076 10010
rect 5540 9976 5552 10010
rect 5064 9970 5552 9976
rect 3798 9378 3804 9900
rect 4772 9896 4782 9926
rect 3798 9350 3814 9378
rect 4776 9374 4782 9896
rect 3028 9300 3516 9306
rect 3028 9266 3040 9300
rect 3504 9266 3516 9300
rect 3028 9260 3516 9266
rect 3236 9198 3296 9260
rect 3028 9192 3516 9198
rect 3028 9158 3040 9192
rect 3504 9158 3516 9192
rect 3028 9152 3516 9158
rect 2734 9086 2746 9108
rect 1762 8554 1768 9082
rect 2740 8558 2746 9086
rect 1762 8532 1774 8554
rect 1714 8290 1774 8532
rect 2734 8532 2746 8558
rect 2780 9086 2794 9108
rect 3754 9108 3814 9350
rect 4772 9350 4782 9374
rect 4816 9896 4832 9926
rect 5792 9926 5852 10168
rect 6804 10168 6818 10186
rect 6852 10716 6864 10744
rect 7826 10744 7886 10986
rect 8846 10986 8854 11006
rect 8888 11528 8906 11562
rect 9862 11562 9922 11804
rect 10884 11804 10890 12380
rect 10924 12356 10944 12380
rect 10924 11818 10930 12356
rect 10924 11804 10944 11818
rect 10154 11754 10642 11760
rect 10154 11720 10166 11754
rect 10630 11720 10642 11754
rect 10154 11714 10642 11720
rect 10356 11652 10416 11714
rect 10154 11646 10642 11652
rect 10154 11612 10166 11646
rect 10630 11612 10642 11646
rect 10154 11606 10642 11612
rect 9862 11532 9872 11562
rect 8888 11006 8894 11528
rect 9866 11010 9872 11532
rect 8888 10986 8906 11006
rect 8118 10936 8606 10942
rect 8118 10902 8130 10936
rect 8594 10902 8606 10936
rect 8118 10896 8606 10902
rect 8322 10834 8382 10896
rect 8118 10828 8606 10834
rect 8118 10794 8130 10828
rect 8594 10794 8606 10828
rect 8118 10788 8606 10794
rect 7826 10716 7836 10744
rect 6852 10186 6858 10716
rect 7830 10186 7836 10716
rect 6852 10168 6864 10186
rect 6082 10118 6570 10124
rect 6082 10084 6094 10118
rect 6558 10084 6570 10118
rect 6082 10078 6570 10084
rect 6286 10016 6346 10078
rect 6082 10010 6570 10016
rect 6082 9976 6094 10010
rect 6558 9976 6570 10010
rect 6082 9970 6570 9976
rect 5792 9904 5800 9926
rect 4816 9374 4822 9896
rect 5794 9382 5800 9904
rect 4816 9350 4832 9374
rect 4046 9300 4534 9306
rect 4046 9266 4058 9300
rect 4522 9266 4534 9300
rect 4046 9260 4534 9266
rect 4256 9198 4316 9260
rect 4046 9192 4534 9198
rect 4046 9158 4058 9192
rect 4522 9158 4534 9192
rect 4046 9152 4534 9158
rect 3754 9088 3764 9108
rect 2780 8558 2786 9086
rect 3758 8560 3764 9088
rect 2780 8532 2794 8558
rect 2010 8482 2498 8488
rect 2010 8448 2022 8482
rect 2486 8448 2498 8482
rect 2010 8442 2498 8448
rect 2224 8380 2284 8442
rect 2010 8374 2498 8380
rect 2010 8340 2022 8374
rect 2486 8340 2498 8374
rect 2010 8334 2498 8340
rect 1714 8264 1728 8290
rect 1722 7714 1728 8264
rect 1762 8264 1774 8290
rect 2734 8290 2794 8532
rect 3754 8532 3764 8560
rect 3798 9088 3814 9108
rect 4772 9108 4832 9350
rect 5792 9350 5800 9382
rect 5834 9904 5852 9926
rect 6804 9926 6864 10168
rect 7826 10168 7836 10186
rect 7870 10716 7886 10744
rect 8846 10744 8906 10986
rect 9862 10986 9872 11010
rect 9906 11532 9922 11562
rect 10884 11562 10944 11804
rect 9906 11010 9912 11532
rect 9906 10986 9922 11010
rect 9136 10936 9624 10942
rect 9136 10902 9148 10936
rect 9612 10902 9624 10936
rect 9136 10896 9624 10902
rect 9334 10834 9394 10896
rect 9136 10828 9624 10834
rect 9136 10794 9148 10828
rect 9612 10794 9624 10828
rect 9136 10788 9624 10794
rect 8846 10716 8854 10744
rect 7870 10186 7876 10716
rect 8848 10186 8854 10716
rect 7870 10168 7886 10186
rect 7100 10118 7588 10124
rect 7100 10084 7112 10118
rect 7576 10084 7588 10118
rect 7100 10078 7588 10084
rect 7302 10016 7362 10078
rect 7100 10010 7588 10016
rect 7100 9976 7112 10010
rect 7576 9976 7588 10010
rect 7100 9970 7588 9976
rect 5834 9382 5840 9904
rect 6804 9896 6818 9926
rect 5834 9350 5852 9382
rect 6812 9374 6818 9896
rect 5064 9300 5552 9306
rect 5064 9266 5076 9300
rect 5540 9266 5552 9300
rect 5064 9260 5552 9266
rect 5258 9198 5318 9260
rect 5064 9192 5552 9198
rect 5064 9158 5076 9192
rect 5540 9158 5552 9192
rect 5064 9152 5552 9158
rect 3798 8560 3804 9088
rect 4772 9084 4782 9108
rect 3798 8532 3814 8560
rect 4776 8556 4782 9084
rect 3028 8482 3516 8488
rect 3028 8448 3040 8482
rect 3504 8448 3516 8482
rect 3028 8442 3516 8448
rect 3238 8380 3298 8442
rect 3028 8374 3516 8380
rect 3028 8340 3040 8374
rect 3504 8340 3516 8374
rect 3028 8334 3516 8340
rect 2734 8268 2746 8290
rect 1762 7714 1768 8264
rect 1722 7702 1768 7714
rect 2740 7714 2746 8268
rect 2780 8268 2794 8290
rect 3754 8290 3814 8532
rect 4772 8532 4782 8556
rect 4816 9084 4832 9108
rect 5792 9108 5852 9350
rect 6804 9350 6818 9374
rect 6852 9896 6864 9926
rect 7826 9926 7886 10168
rect 8846 10168 8854 10186
rect 8888 10716 8906 10744
rect 9862 10744 9922 10986
rect 10884 10986 10890 11562
rect 10924 11528 10944 11562
rect 10924 11006 10930 11528
rect 10924 10986 10944 11006
rect 10154 10936 10642 10942
rect 10154 10902 10166 10936
rect 10630 10902 10642 10936
rect 10154 10896 10642 10902
rect 10354 10834 10414 10896
rect 10154 10828 10642 10834
rect 10154 10794 10166 10828
rect 10630 10794 10642 10828
rect 10154 10788 10642 10794
rect 9862 10720 9872 10744
rect 8888 10186 8894 10716
rect 9866 10190 9872 10720
rect 8888 10168 8906 10186
rect 8118 10118 8606 10124
rect 8118 10084 8130 10118
rect 8594 10084 8606 10118
rect 8118 10078 8606 10084
rect 8324 10016 8384 10078
rect 8118 10010 8606 10016
rect 8118 9976 8130 10010
rect 8594 9976 8606 10010
rect 8118 9970 8606 9976
rect 7826 9896 7836 9926
rect 6852 9374 6858 9896
rect 7830 9374 7836 9896
rect 6852 9350 6864 9374
rect 6082 9300 6570 9306
rect 6082 9266 6094 9300
rect 6558 9266 6570 9300
rect 6082 9260 6570 9266
rect 6288 9198 6348 9260
rect 6082 9192 6570 9198
rect 6082 9158 6094 9192
rect 6558 9158 6570 9192
rect 6082 9152 6570 9158
rect 5792 9092 5800 9108
rect 4816 8556 4822 9084
rect 5794 8564 5800 9092
rect 4816 8532 4832 8556
rect 4046 8482 4534 8488
rect 4046 8448 4058 8482
rect 4522 8448 4534 8482
rect 4046 8442 4534 8448
rect 4258 8380 4318 8442
rect 4046 8374 4534 8380
rect 4046 8340 4058 8374
rect 4522 8340 4534 8374
rect 4046 8334 4534 8340
rect 3754 8270 3764 8290
rect 2780 7714 2786 8268
rect 3758 7760 3764 8270
rect 2740 7702 2786 7714
rect 3748 7714 3764 7760
rect 3798 8270 3814 8290
rect 4772 8290 4832 8532
rect 5792 8532 5800 8564
rect 5834 9092 5852 9108
rect 6804 9108 6864 9350
rect 7826 9350 7836 9374
rect 7870 9896 7886 9926
rect 8846 9926 8906 10168
rect 9862 10168 9872 10190
rect 9906 10720 9922 10744
rect 10884 10744 10944 10986
rect 9906 10190 9912 10720
rect 9906 10168 9922 10190
rect 9136 10118 9624 10124
rect 9136 10084 9148 10118
rect 9612 10084 9624 10118
rect 9136 10078 9624 10084
rect 9336 10016 9396 10078
rect 9136 10010 9624 10016
rect 9136 9976 9148 10010
rect 9612 9976 9624 10010
rect 9136 9970 9624 9976
rect 8846 9896 8854 9926
rect 7870 9374 7876 9896
rect 8848 9374 8854 9896
rect 7870 9350 7886 9374
rect 7100 9300 7588 9306
rect 7100 9266 7112 9300
rect 7576 9266 7588 9300
rect 7100 9260 7588 9266
rect 7304 9198 7364 9260
rect 7100 9192 7588 9198
rect 7100 9158 7112 9192
rect 7576 9158 7588 9192
rect 7100 9152 7588 9158
rect 5834 8564 5840 9092
rect 6804 9084 6818 9108
rect 5834 8532 5852 8564
rect 6812 8556 6818 9084
rect 5064 8482 5552 8488
rect 5064 8448 5076 8482
rect 5540 8448 5552 8482
rect 5064 8442 5552 8448
rect 5260 8380 5320 8442
rect 5064 8374 5552 8380
rect 5064 8340 5076 8374
rect 5540 8340 5552 8374
rect 5064 8334 5552 8340
rect 3798 7760 3804 8270
rect 4772 8266 4782 8290
rect 3798 7714 3808 7760
rect 2010 7664 2498 7670
rect 2010 7630 2022 7664
rect 2486 7630 2498 7664
rect 2010 7624 2498 7630
rect 3028 7664 3516 7670
rect 3028 7630 3040 7664
rect 3504 7630 3516 7664
rect 3028 7624 3516 7630
rect 3748 7540 3808 7714
rect 4776 7714 4782 8266
rect 4816 8266 4832 8290
rect 5792 8290 5852 8532
rect 6804 8532 6818 8556
rect 6852 9084 6864 9108
rect 7826 9108 7886 9350
rect 8846 9350 8854 9374
rect 8888 9896 8906 9926
rect 9862 9926 9922 10168
rect 10884 10168 10890 10744
rect 10924 10716 10944 10744
rect 10924 10186 10930 10716
rect 10924 10168 10944 10186
rect 10154 10118 10642 10124
rect 10154 10084 10166 10118
rect 10630 10084 10642 10118
rect 10154 10078 10642 10084
rect 10356 10016 10416 10078
rect 10154 10010 10642 10016
rect 10154 9976 10166 10010
rect 10630 9976 10642 10010
rect 10154 9970 10642 9976
rect 9862 9900 9872 9926
rect 8888 9374 8894 9896
rect 9866 9378 9872 9900
rect 8888 9350 8906 9374
rect 8118 9300 8606 9306
rect 8118 9266 8130 9300
rect 8594 9266 8606 9300
rect 8118 9260 8606 9266
rect 8326 9198 8386 9260
rect 8118 9192 8606 9198
rect 8118 9158 8130 9192
rect 8594 9158 8606 9192
rect 8118 9152 8606 9158
rect 7826 9084 7836 9108
rect 6852 8556 6858 9084
rect 7830 8556 7836 9084
rect 6852 8532 6864 8556
rect 6082 8482 6570 8488
rect 6082 8448 6094 8482
rect 6558 8448 6570 8482
rect 6082 8442 6570 8448
rect 6290 8380 6350 8442
rect 6082 8374 6570 8380
rect 6082 8340 6094 8374
rect 6558 8340 6570 8374
rect 6082 8334 6570 8340
rect 5792 8274 5800 8290
rect 4816 7714 4822 8266
rect 5794 7762 5800 8274
rect 4776 7702 4822 7714
rect 5786 7714 5800 7762
rect 5834 8274 5852 8290
rect 6804 8290 6864 8532
rect 7826 8532 7836 8556
rect 7870 9084 7886 9108
rect 8846 9108 8906 9350
rect 9862 9350 9872 9378
rect 9906 9900 9922 9926
rect 10884 9926 10944 10168
rect 9906 9378 9912 9900
rect 9906 9350 9922 9378
rect 9136 9300 9624 9306
rect 9136 9266 9148 9300
rect 9612 9266 9624 9300
rect 9136 9260 9624 9266
rect 9338 9198 9398 9260
rect 9136 9192 9624 9198
rect 9136 9158 9148 9192
rect 9612 9158 9624 9192
rect 9136 9152 9624 9158
rect 8846 9084 8854 9108
rect 7870 8556 7876 9084
rect 8848 8556 8854 9084
rect 7870 8532 7886 8556
rect 7100 8482 7588 8488
rect 7100 8448 7112 8482
rect 7576 8448 7588 8482
rect 7100 8442 7588 8448
rect 7306 8380 7366 8442
rect 7100 8374 7588 8380
rect 7100 8340 7112 8374
rect 7576 8340 7588 8374
rect 7100 8334 7588 8340
rect 5834 7762 5840 8274
rect 6804 8266 6818 8290
rect 5834 7714 5846 7762
rect 4046 7664 4534 7670
rect 4046 7630 4058 7664
rect 4522 7630 4534 7664
rect 4046 7624 4534 7630
rect 5064 7664 5552 7670
rect 5064 7630 5076 7664
rect 5540 7630 5552 7664
rect 5064 7624 5552 7630
rect 5786 7540 5846 7714
rect 6812 7714 6818 8266
rect 6852 8266 6864 8290
rect 7826 8290 7886 8532
rect 8846 8532 8854 8556
rect 8888 9084 8906 9108
rect 9862 9108 9922 9350
rect 10884 9350 10890 9926
rect 10924 9896 10944 9926
rect 10924 9374 10930 9896
rect 10924 9350 10944 9374
rect 10154 9300 10642 9306
rect 10154 9266 10166 9300
rect 10630 9266 10642 9300
rect 10154 9260 10642 9266
rect 10358 9198 10418 9260
rect 10154 9192 10642 9198
rect 10154 9158 10166 9192
rect 10630 9158 10642 9192
rect 10154 9152 10642 9158
rect 9862 9088 9872 9108
rect 8888 8556 8894 9084
rect 9866 8560 9872 9088
rect 8888 8532 8906 8556
rect 8118 8482 8606 8488
rect 8118 8448 8130 8482
rect 8594 8448 8606 8482
rect 8118 8442 8606 8448
rect 8328 8380 8388 8442
rect 8118 8374 8606 8380
rect 8118 8340 8130 8374
rect 8594 8340 8606 8374
rect 8118 8334 8606 8340
rect 7826 8266 7836 8290
rect 6852 7714 6858 8266
rect 7830 7758 7836 8266
rect 6812 7702 6858 7714
rect 7822 7714 7836 7758
rect 7870 8266 7886 8290
rect 8846 8290 8906 8532
rect 9862 8532 9872 8560
rect 9906 9088 9922 9108
rect 10884 9108 10944 9350
rect 9906 8560 9912 9088
rect 9906 8532 9922 8560
rect 9136 8482 9624 8488
rect 9136 8448 9148 8482
rect 9612 8448 9624 8482
rect 9136 8442 9624 8448
rect 9340 8380 9400 8442
rect 9136 8374 9624 8380
rect 9136 8340 9148 8374
rect 9612 8340 9624 8374
rect 9136 8334 9624 8340
rect 8846 8266 8854 8290
rect 7870 7758 7876 8266
rect 7870 7714 7882 7758
rect 6082 7664 6570 7670
rect 6082 7630 6094 7664
rect 6558 7630 6570 7664
rect 6082 7624 6570 7630
rect 7100 7664 7588 7670
rect 7100 7630 7112 7664
rect 7576 7630 7588 7664
rect 7100 7624 7588 7630
rect 7822 7540 7882 7714
rect 8848 7714 8854 8266
rect 8888 8266 8906 8290
rect 9862 8290 9922 8532
rect 10884 8532 10890 9108
rect 10924 9084 10944 9108
rect 10924 8556 10930 9084
rect 10924 8532 10944 8556
rect 10154 8482 10642 8488
rect 10154 8448 10166 8482
rect 10630 8448 10642 8482
rect 10154 8442 10642 8448
rect 10360 8380 10420 8442
rect 10154 8374 10642 8380
rect 10154 8340 10166 8374
rect 10630 8340 10642 8374
rect 10154 8334 10642 8340
rect 9862 8270 9872 8290
rect 8888 7714 8894 8266
rect 9866 7756 9872 8270
rect 8848 7702 8894 7714
rect 9858 7714 9872 7756
rect 9906 8270 9922 8290
rect 10884 8290 10944 8532
rect 9906 7756 9912 8270
rect 10884 7768 10890 8290
rect 9906 7714 9918 7756
rect 8118 7664 8606 7670
rect 8118 7630 8130 7664
rect 8594 7630 8606 7664
rect 8118 7624 8606 7630
rect 9136 7664 9624 7670
rect 9136 7630 9148 7664
rect 9612 7630 9624 7664
rect 9136 7624 9624 7630
rect 9858 7540 9918 7714
rect 10878 7714 10890 7768
rect 10924 8266 10944 8290
rect 10924 7768 10930 8266
rect 10924 7714 10938 7768
rect 12062 7718 12122 14858
rect 10154 7664 10642 7670
rect 10154 7630 10166 7664
rect 10630 7630 10642 7664
rect 10154 7624 10642 7630
rect 10372 7540 10432 7624
rect 10878 7540 10938 7714
rect 12056 7658 12062 7718
rect 12122 7658 12128 7718
rect 3748 7480 12042 7540
rect 7508 6732 7514 6792
rect 7574 6732 7580 6792
rect 1404 6646 1464 6652
rect 5478 6586 5484 6646
rect 5544 6586 5550 6646
rect 244 6458 250 6518
rect 310 6458 316 6518
rect 250 4286 310 6458
rect 1404 6454 1464 6586
rect 2922 6458 2928 6518
rect 2988 6458 2994 6518
rect 3954 6458 3960 6518
rect 4020 6458 4026 6518
rect 388 6394 1464 6454
rect 388 6266 448 6394
rect 896 6356 956 6394
rect 686 6350 1174 6356
rect 686 6316 698 6350
rect 1162 6316 1174 6350
rect 686 6310 1174 6316
rect 388 6220 404 6266
rect 398 5690 404 6220
rect 438 6220 448 6266
rect 1404 6266 1464 6394
rect 2928 6356 2988 6458
rect 3960 6356 4020 6458
rect 1704 6350 2192 6356
rect 1704 6316 1716 6350
rect 2180 6316 2192 6350
rect 1704 6310 2192 6316
rect 2722 6350 3210 6356
rect 2722 6316 2734 6350
rect 3198 6316 3210 6350
rect 2722 6310 3210 6316
rect 3740 6350 4228 6356
rect 3740 6316 3752 6350
rect 4216 6316 4228 6350
rect 3740 6310 4228 6316
rect 4758 6350 5246 6356
rect 4758 6316 4770 6350
rect 5234 6316 5246 6350
rect 4758 6310 5246 6316
rect 1404 6226 1422 6266
rect 438 5690 444 6220
rect 398 5678 444 5690
rect 1416 5690 1422 6226
rect 1456 6226 1464 6266
rect 2434 6266 2480 6278
rect 1456 5690 1462 6226
rect 2434 5754 2440 6266
rect 1416 5678 1462 5690
rect 2426 5690 2440 5754
rect 2474 5754 2480 6266
rect 3452 6266 3498 6278
rect 2474 5690 2486 5754
rect 3452 5736 3458 6266
rect 686 5640 1174 5646
rect 686 5606 698 5640
rect 1162 5606 1174 5640
rect 686 5600 1174 5606
rect 1704 5640 2192 5646
rect 1704 5606 1716 5640
rect 2180 5606 2192 5640
rect 1704 5600 2192 5606
rect 1908 5556 1968 5600
rect 1902 5496 1908 5556
rect 1968 5496 1974 5556
rect 1402 5392 1408 5452
rect 1468 5392 1474 5452
rect 1408 5350 1468 5392
rect 388 5290 1468 5350
rect 388 5154 448 5290
rect 892 5244 952 5290
rect 686 5238 1174 5244
rect 686 5204 698 5238
rect 1162 5204 1174 5238
rect 686 5198 1174 5204
rect 388 5108 404 5154
rect 398 4578 404 5108
rect 438 5108 448 5154
rect 1408 5154 1468 5290
rect 2426 5348 2486 5690
rect 3444 5690 3458 5736
rect 3492 5736 3498 6266
rect 4470 6266 4516 6278
rect 4470 5752 4476 6266
rect 3492 5690 3504 5736
rect 2722 5640 3210 5646
rect 2722 5606 2734 5640
rect 3198 5606 3210 5640
rect 2722 5600 3210 5606
rect 2926 5496 2932 5556
rect 2992 5496 2998 5556
rect 1704 5238 2192 5244
rect 1704 5204 1716 5238
rect 2180 5204 2192 5238
rect 1704 5198 2192 5204
rect 438 4578 444 5108
rect 398 4566 444 4578
rect 1408 4578 1422 5154
rect 1456 4578 1468 5154
rect 686 4528 1174 4534
rect 686 4494 698 4528
rect 1162 4494 1174 4528
rect 686 4488 1174 4494
rect 244 4226 250 4286
rect 310 4226 316 4286
rect 250 2160 310 4226
rect 686 4126 1174 4132
rect 686 4092 698 4126
rect 1162 4092 1174 4126
rect 686 4086 1174 4092
rect 398 4042 444 4054
rect 398 3500 404 4042
rect 392 3466 404 3500
rect 438 3500 444 4042
rect 1408 4042 1468 4578
rect 2426 5154 2486 5288
rect 2932 5244 2992 5496
rect 3444 5452 3504 5690
rect 4462 5690 4476 5752
rect 4510 5752 4516 6266
rect 5484 6266 5544 6586
rect 7014 6458 7020 6518
rect 7080 6458 7086 6518
rect 7020 6356 7080 6458
rect 5776 6350 6264 6356
rect 5776 6316 5788 6350
rect 6252 6316 6264 6350
rect 5776 6310 6264 6316
rect 6794 6350 7282 6356
rect 6794 6316 6806 6350
rect 7270 6316 7282 6350
rect 6794 6310 7282 6316
rect 5484 6202 5494 6266
rect 4510 5690 4522 5752
rect 3740 5640 4228 5646
rect 3740 5606 3752 5640
rect 4216 5606 4228 5640
rect 3740 5600 4228 5606
rect 3958 5496 3964 5556
rect 4024 5496 4030 5556
rect 3438 5392 3444 5452
rect 3504 5392 3510 5452
rect 3964 5244 4024 5496
rect 4462 5348 4522 5690
rect 5488 5690 5494 6202
rect 5528 6202 5544 6266
rect 6506 6266 6552 6278
rect 5528 5690 5534 6202
rect 6506 5762 6512 6266
rect 5488 5678 5534 5690
rect 6494 5690 6512 5762
rect 6546 5762 6552 6266
rect 7514 6266 7574 6732
rect 9538 6586 9544 6646
rect 9604 6586 9610 6646
rect 11722 6586 11728 6646
rect 11788 6586 11794 6646
rect 8010 6458 8016 6518
rect 8076 6458 8082 6518
rect 8016 6356 8076 6458
rect 7812 6350 8300 6356
rect 7812 6316 7824 6350
rect 8288 6316 8300 6350
rect 7812 6310 8300 6316
rect 8830 6350 9318 6356
rect 8830 6316 8842 6350
rect 9306 6316 9318 6350
rect 8830 6310 9318 6316
rect 8016 6308 8076 6310
rect 9544 6278 9604 6586
rect 9848 6350 10336 6356
rect 9848 6316 9860 6350
rect 10324 6316 10336 6350
rect 9848 6310 10336 6316
rect 10866 6350 11354 6356
rect 10866 6316 10878 6350
rect 11342 6316 11354 6350
rect 10866 6310 11354 6316
rect 6546 5690 6554 5762
rect 4758 5640 5246 5646
rect 4758 5606 4770 5640
rect 5234 5606 5246 5640
rect 4758 5600 5246 5606
rect 5776 5640 6264 5646
rect 5776 5606 5788 5640
rect 6252 5606 6264 5640
rect 5776 5600 6264 5606
rect 4964 5556 5024 5600
rect 5984 5556 6044 5600
rect 4958 5496 4964 5556
rect 5024 5496 5030 5556
rect 5978 5496 5984 5556
rect 6044 5496 6050 5556
rect 5474 5392 5480 5452
rect 5540 5392 5546 5452
rect 2722 5238 3210 5244
rect 2722 5204 2734 5238
rect 3198 5204 3210 5238
rect 2722 5198 3210 5204
rect 3740 5238 4228 5244
rect 3740 5204 3752 5238
rect 4216 5204 4228 5238
rect 3740 5198 4228 5204
rect 2426 4578 2440 5154
rect 2474 4578 2486 5154
rect 3452 5154 3498 5166
rect 3452 4616 3458 5154
rect 1704 4528 2192 4534
rect 1704 4494 1716 4528
rect 2180 4494 2192 4528
rect 1704 4488 2192 4494
rect 1900 4286 1960 4488
rect 1894 4226 1900 4286
rect 1960 4226 1966 4286
rect 1900 4132 1960 4226
rect 1704 4126 2192 4132
rect 1704 4092 1716 4126
rect 2180 4092 2192 4126
rect 1704 4086 2192 4092
rect 1408 3970 1422 4042
rect 438 3466 452 3500
rect 1416 3496 1422 3970
rect 392 3334 452 3466
rect 1412 3466 1422 3496
rect 1456 3970 1468 4042
rect 2426 4042 2486 4578
rect 3438 4578 3458 4616
rect 3492 4578 3498 5154
rect 2722 4528 3210 4534
rect 2722 4494 2734 4528
rect 3198 4494 3210 4528
rect 2722 4488 3210 4494
rect 3438 4406 3498 4578
rect 4462 5154 4522 5288
rect 4758 5238 5246 5244
rect 4758 5204 4770 5238
rect 5234 5204 5246 5238
rect 4758 5198 5246 5204
rect 4462 4578 4476 5154
rect 4510 4578 4522 5154
rect 3740 4528 4228 4534
rect 3740 4494 3752 4528
rect 4216 4494 4228 4528
rect 3740 4488 4228 4494
rect 3432 4346 3438 4406
rect 3498 4346 3504 4406
rect 2722 4126 3210 4132
rect 2722 4092 2734 4126
rect 3198 4092 3210 4126
rect 2722 4086 3210 4092
rect 1456 3496 1462 3970
rect 1456 3466 1472 3496
rect 686 3416 1174 3422
rect 686 3382 698 3416
rect 1162 3382 1174 3416
rect 686 3376 1174 3382
rect 884 3334 944 3376
rect 1412 3334 1472 3466
rect 2426 3466 2440 4042
rect 2474 3466 2486 4042
rect 3438 4042 3498 4346
rect 3740 4126 4228 4132
rect 3740 4092 3752 4126
rect 4216 4092 4228 4126
rect 3740 4086 4228 4092
rect 3438 3972 3458 4042
rect 1704 3416 2192 3422
rect 1704 3382 1716 3416
rect 2180 3382 2192 3416
rect 1704 3376 2192 3382
rect 392 3274 1472 3334
rect 1412 3234 1472 3274
rect 2426 3342 2486 3466
rect 3452 3466 3458 3972
rect 3492 3466 3498 4042
rect 3452 3454 3498 3466
rect 4462 4042 4522 4578
rect 5480 5154 5540 5392
rect 6494 5348 6554 5690
rect 7514 5690 7530 6266
rect 7564 5690 7574 6266
rect 8542 6266 8588 6278
rect 8542 5752 8548 6266
rect 6794 5640 7282 5646
rect 6794 5606 6806 5640
rect 7270 5606 7282 5640
rect 6794 5600 7282 5606
rect 6998 5496 7004 5556
rect 7064 5496 7070 5556
rect 6488 5288 6494 5348
rect 6554 5288 6560 5348
rect 5776 5238 6264 5244
rect 5776 5204 5788 5238
rect 6252 5204 6264 5238
rect 5776 5198 6264 5204
rect 5480 4578 5494 5154
rect 5528 4578 5540 5154
rect 4758 4528 5246 4534
rect 4758 4494 4770 4528
rect 5234 4494 5246 4528
rect 4758 4488 5246 4494
rect 4970 4286 5030 4488
rect 4964 4226 4970 4286
rect 5030 4226 5036 4286
rect 4970 4132 5030 4226
rect 4758 4126 5246 4132
rect 4758 4092 4770 4126
rect 5234 4092 5246 4126
rect 4758 4086 5246 4092
rect 4462 3466 4476 4042
rect 4510 3466 4522 4042
rect 5480 4042 5540 4578
rect 6494 5154 6554 5288
rect 7004 5244 7064 5496
rect 7514 5452 7574 5690
rect 8528 5690 8548 5752
rect 8582 5690 8588 6266
rect 9544 6266 9606 6278
rect 9544 6234 9566 6266
rect 7812 5640 8300 5646
rect 7812 5606 7824 5640
rect 8288 5606 8300 5640
rect 7812 5600 8300 5606
rect 8014 5556 8074 5562
rect 7508 5392 7514 5452
rect 7574 5392 7580 5452
rect 8014 5244 8074 5496
rect 8528 5348 8588 5690
rect 9560 5690 9566 6234
rect 9600 5690 9606 6266
rect 10578 6266 10624 6278
rect 10578 5724 10584 6266
rect 9560 5678 9606 5690
rect 10572 5690 10584 5724
rect 10618 5724 10624 6266
rect 11596 6266 11642 6278
rect 11596 5744 11602 6266
rect 10618 5690 10632 5724
rect 8830 5640 9318 5646
rect 8830 5606 8842 5640
rect 9306 5606 9318 5640
rect 8830 5600 9318 5606
rect 9848 5640 10336 5646
rect 9848 5606 9860 5640
rect 10324 5606 10336 5640
rect 9848 5600 10336 5606
rect 9028 5556 9088 5600
rect 10046 5556 10106 5600
rect 9022 5496 9028 5556
rect 9088 5496 9094 5556
rect 10046 5490 10106 5496
rect 10572 5462 10632 5690
rect 11588 5690 11602 5744
rect 11636 5744 11642 6266
rect 11636 5690 11648 5744
rect 10866 5640 11354 5646
rect 10866 5606 10878 5640
rect 11342 5606 11354 5640
rect 10866 5600 11354 5606
rect 11076 5462 11136 5600
rect 11588 5462 11648 5690
rect 9544 5392 9550 5452
rect 9610 5392 9616 5452
rect 10572 5402 11648 5462
rect 6794 5238 7282 5244
rect 6794 5204 6806 5238
rect 7270 5204 7282 5238
rect 6794 5198 7282 5204
rect 7812 5238 8300 5244
rect 7812 5204 7824 5238
rect 8288 5204 8300 5238
rect 7812 5198 8300 5204
rect 6494 4578 6512 5154
rect 6546 4578 6554 5154
rect 7524 5154 7570 5166
rect 7524 4634 7530 5154
rect 5776 4528 6264 4534
rect 5776 4494 5788 4528
rect 6252 4494 6264 4528
rect 5776 4488 6264 4494
rect 5978 4286 6038 4488
rect 5972 4226 5978 4286
rect 6038 4226 6044 4286
rect 5978 4132 6038 4226
rect 5776 4126 6264 4132
rect 5776 4092 5788 4126
rect 6252 4092 6264 4126
rect 5776 4086 6264 4092
rect 5480 3936 5494 4042
rect 5488 3528 5494 3936
rect 2722 3416 3210 3422
rect 2722 3382 2734 3416
rect 3198 3382 3210 3416
rect 2722 3376 3210 3382
rect 3740 3416 4228 3422
rect 3740 3382 3752 3416
rect 4216 3382 4228 3416
rect 3740 3376 4228 3382
rect 1406 3174 1412 3234
rect 1472 3174 1478 3234
rect 1900 3062 1906 3122
rect 1966 3062 1972 3122
rect 1906 3020 1966 3062
rect 686 3014 1174 3020
rect 686 2980 698 3014
rect 1162 2980 1174 3014
rect 686 2974 1174 2980
rect 1704 3014 2192 3020
rect 1704 2980 1716 3014
rect 2180 2980 2192 3014
rect 1704 2974 2192 2980
rect 398 2930 444 2942
rect 398 2396 404 2930
rect 388 2354 404 2396
rect 438 2396 444 2930
rect 1416 2930 1462 2942
rect 438 2354 448 2396
rect 1416 2390 1422 2930
rect 388 2210 448 2354
rect 1406 2354 1422 2390
rect 1456 2390 1462 2930
rect 2426 2930 2486 3282
rect 2930 3122 2990 3376
rect 3442 3174 3448 3234
rect 3508 3174 3514 3234
rect 2924 3062 2930 3122
rect 2990 3062 2996 3122
rect 2722 3014 3210 3020
rect 2722 2980 2734 3014
rect 3198 2980 3210 3014
rect 2722 2974 3210 2980
rect 2426 2828 2440 2930
rect 1456 2354 1466 2390
rect 686 2304 1174 2310
rect 686 2270 698 2304
rect 1162 2270 1174 2304
rect 686 2264 1174 2270
rect 892 2210 952 2264
rect 1406 2210 1466 2354
rect 2434 2354 2440 2828
rect 2474 2828 2486 2930
rect 3448 2930 3508 3174
rect 3962 3122 4022 3376
rect 4462 3342 4522 3466
rect 5484 3466 5494 3528
rect 5528 3936 5540 4042
rect 6494 4042 6554 4578
rect 7514 4578 7530 4634
rect 7564 4634 7570 5154
rect 8528 5154 8588 5288
rect 8830 5238 9318 5244
rect 8830 5204 8842 5238
rect 9306 5204 9318 5238
rect 8830 5198 9318 5204
rect 7564 4578 7574 4634
rect 6794 4528 7282 4534
rect 6794 4494 6806 4528
rect 7270 4494 7282 4528
rect 6794 4488 7282 4494
rect 7514 4406 7574 4578
rect 8528 4578 8548 5154
rect 8582 4578 8588 5154
rect 7812 4528 8300 4534
rect 7812 4494 7824 4528
rect 8288 4494 8300 4528
rect 7812 4488 8300 4494
rect 7508 4346 7514 4406
rect 7574 4346 7580 4406
rect 6794 4126 7282 4132
rect 6794 4092 6806 4126
rect 7270 4092 7282 4126
rect 6794 4086 7282 4092
rect 5528 3528 5534 3936
rect 5528 3466 5544 3528
rect 4758 3416 5246 3422
rect 4758 3382 4770 3416
rect 5234 3382 5246 3416
rect 4758 3376 5246 3382
rect 3956 3062 3962 3122
rect 4022 3062 4028 3122
rect 3740 3014 4228 3020
rect 3740 2980 3752 3014
rect 4216 2980 4228 3014
rect 3740 2974 4228 2980
rect 3448 2890 3458 2930
rect 2474 2354 2480 2828
rect 2434 2342 2480 2354
rect 3452 2354 3458 2890
rect 3492 2890 3508 2930
rect 4462 2930 4522 3282
rect 5484 3234 5544 3466
rect 6494 3466 6512 4042
rect 6546 3466 6554 4042
rect 7514 4042 7574 4346
rect 7812 4126 8300 4132
rect 7812 4092 7824 4126
rect 8288 4092 8300 4126
rect 7812 4086 8300 4092
rect 7514 4000 7530 4042
rect 5776 3416 6264 3422
rect 5776 3382 5788 3416
rect 6252 3382 6264 3416
rect 5776 3376 6264 3382
rect 6494 3342 6554 3466
rect 7524 3466 7530 4000
rect 7564 4000 7574 4042
rect 8528 4042 8588 4578
rect 9550 5154 9610 5392
rect 10572 5348 10632 5402
rect 9848 5238 10336 5244
rect 9848 5204 9860 5238
rect 10324 5204 10336 5238
rect 9848 5198 10336 5204
rect 9550 4578 9566 5154
rect 9600 4578 9610 5154
rect 8830 4528 9318 4534
rect 8830 4494 8842 4528
rect 9306 4494 9318 4528
rect 8830 4488 9318 4494
rect 9040 4286 9100 4488
rect 9034 4226 9040 4286
rect 9100 4226 9106 4286
rect 9040 4132 9100 4226
rect 8830 4126 9318 4132
rect 8830 4092 8842 4126
rect 9306 4092 9318 4126
rect 8830 4086 9318 4092
rect 7564 3466 7570 4000
rect 7524 3454 7570 3466
rect 8528 3466 8548 4042
rect 8582 3466 8588 4042
rect 9550 4042 9610 4578
rect 10572 5154 10632 5288
rect 11076 5244 11136 5402
rect 10866 5238 11354 5244
rect 10866 5204 10878 5238
rect 11342 5204 11354 5238
rect 10866 5198 11354 5204
rect 10572 4578 10584 5154
rect 10618 4578 10632 5154
rect 9848 4528 10336 4534
rect 9848 4494 9860 4528
rect 10324 4494 10336 4528
rect 9848 4488 10336 4494
rect 10066 4286 10126 4488
rect 10572 4342 10632 4578
rect 11588 5154 11648 5402
rect 11588 4578 11602 5154
rect 11636 4578 11648 5154
rect 10866 4528 11354 4534
rect 10866 4494 10878 4528
rect 11342 4494 11354 4528
rect 10866 4488 11354 4494
rect 11072 4342 11132 4488
rect 11588 4342 11648 4578
rect 11728 4406 11788 6586
rect 11842 5496 11848 5556
rect 11908 5496 11914 5556
rect 11722 4346 11728 4406
rect 11788 4346 11794 4406
rect 10060 4226 10066 4286
rect 10126 4226 10132 4286
rect 10572 4282 11648 4342
rect 10066 4132 10126 4226
rect 9848 4126 10336 4132
rect 9848 4092 9860 4126
rect 10324 4092 10336 4126
rect 9848 4086 10336 4092
rect 9550 3986 9566 4042
rect 9560 3512 9566 3986
rect 6794 3416 7282 3422
rect 6794 3382 6806 3416
rect 7270 3382 7282 3416
rect 6794 3376 7282 3382
rect 7812 3416 8300 3422
rect 7812 3382 7824 3416
rect 8288 3382 8300 3416
rect 7812 3376 8300 3382
rect 5478 3174 5484 3234
rect 5544 3174 5550 3234
rect 4956 3062 4962 3122
rect 5022 3062 5028 3122
rect 5976 3062 5982 3122
rect 6042 3062 6048 3122
rect 4962 3020 5022 3062
rect 5982 3020 6042 3062
rect 4758 3014 5246 3020
rect 4758 2980 4770 3014
rect 5234 2980 5246 3014
rect 4758 2974 5246 2980
rect 5776 3014 6264 3020
rect 5776 2980 5788 3014
rect 6252 2980 6264 3014
rect 5776 2974 6264 2980
rect 4462 2892 4476 2930
rect 3492 2354 3498 2890
rect 3452 2342 3498 2354
rect 4470 2354 4476 2892
rect 4510 2892 4522 2930
rect 5488 2930 5534 2942
rect 4510 2354 4516 2892
rect 5488 2414 5494 2930
rect 4470 2342 4516 2354
rect 5486 2354 5494 2414
rect 5528 2414 5534 2930
rect 6494 2930 6554 3282
rect 7002 3122 7062 3376
rect 7512 3174 7518 3234
rect 7578 3174 7584 3234
rect 6996 3062 7002 3122
rect 7062 3062 7068 3122
rect 6794 3014 7282 3020
rect 6794 2980 6806 3014
rect 7270 2980 7282 3014
rect 6794 2974 7282 2980
rect 6494 2870 6512 2930
rect 5528 2354 5546 2414
rect 1704 2304 2192 2310
rect 1704 2270 1716 2304
rect 2180 2270 2192 2304
rect 1704 2264 2192 2270
rect 2722 2304 3210 2310
rect 2722 2270 2734 2304
rect 3198 2270 3210 2304
rect 2722 2264 3210 2270
rect 3740 2304 4228 2310
rect 3740 2270 3752 2304
rect 4216 2270 4228 2304
rect 3740 2264 4228 2270
rect 4758 2304 5246 2310
rect 4758 2270 4770 2304
rect 5234 2270 5246 2304
rect 4758 2264 5246 2270
rect 244 2100 250 2160
rect 310 2100 316 2160
rect 388 2150 1466 2210
rect 2920 2160 2980 2264
rect 3952 2160 4012 2264
rect 1406 2030 1466 2150
rect 2914 2100 2920 2160
rect 2980 2100 2986 2160
rect 3946 2100 3952 2160
rect 4012 2100 4018 2160
rect 5486 2030 5546 2354
rect 6506 2354 6512 2870
rect 6546 2870 6554 2930
rect 7518 2930 7578 3174
rect 8012 3122 8072 3376
rect 8012 3056 8072 3062
rect 8528 3342 8588 3466
rect 9554 3466 9566 3512
rect 9600 3986 9610 4042
rect 10572 4042 10632 4282
rect 11072 4132 11132 4282
rect 10866 4126 11354 4132
rect 10866 4092 10878 4126
rect 11342 4092 11354 4126
rect 10866 4086 11354 4092
rect 9600 3512 9606 3986
rect 9600 3466 9614 3512
rect 8830 3416 9318 3422
rect 8830 3382 8842 3416
rect 9306 3382 9318 3416
rect 8830 3376 9318 3382
rect 7812 3014 8300 3020
rect 7812 2980 7824 3014
rect 8288 2980 8300 3014
rect 7812 2974 8300 2980
rect 7518 2884 7530 2930
rect 6546 2354 6552 2870
rect 6506 2342 6552 2354
rect 7524 2354 7530 2884
rect 7564 2884 7578 2930
rect 8528 2930 8588 3282
rect 9554 3234 9614 3466
rect 10572 3466 10584 4042
rect 10618 3466 10632 4042
rect 9848 3416 10336 3422
rect 9848 3382 9860 3416
rect 10324 3382 10336 3416
rect 9848 3376 10336 3382
rect 10572 3342 10632 3466
rect 11588 4042 11648 4282
rect 11588 3466 11602 4042
rect 11636 3466 11648 4042
rect 10866 3416 11354 3422
rect 10866 3382 10878 3416
rect 11342 3382 11354 3416
rect 10866 3376 11354 3382
rect 10566 3282 10572 3342
rect 10632 3282 10638 3342
rect 9548 3174 9554 3234
rect 9614 3174 9620 3234
rect 10572 3230 10632 3282
rect 11080 3230 11140 3376
rect 11588 3230 11648 3466
rect 10572 3170 11648 3230
rect 10044 3122 10104 3128
rect 9020 3062 9026 3122
rect 9086 3062 9092 3122
rect 9026 3020 9086 3062
rect 10044 3020 10104 3062
rect 8830 3014 9318 3020
rect 8830 2980 8842 3014
rect 9306 2980 9318 3014
rect 8830 2974 9318 2980
rect 9848 3014 10336 3020
rect 9848 2980 9860 3014
rect 10324 2980 10336 3014
rect 9848 2974 10336 2980
rect 8528 2888 8548 2930
rect 7564 2354 7570 2884
rect 7524 2342 7570 2354
rect 8542 2354 8548 2888
rect 8582 2354 8588 2930
rect 9560 2930 9606 2942
rect 9560 2382 9566 2930
rect 8542 2342 8588 2354
rect 9546 2354 9566 2382
rect 9600 2354 9606 2930
rect 10572 2930 10632 3170
rect 11080 3020 11140 3170
rect 10866 3014 11354 3020
rect 10866 2980 10878 3014
rect 11342 2980 11354 3014
rect 10866 2974 11354 2980
rect 10572 2866 10584 2930
rect 5776 2304 6264 2310
rect 5776 2270 5788 2304
rect 6252 2270 6264 2304
rect 5776 2264 6264 2270
rect 6794 2304 7282 2310
rect 6794 2270 6806 2304
rect 7270 2270 7282 2304
rect 6794 2264 7282 2270
rect 7812 2304 8300 2310
rect 7812 2270 7824 2304
rect 8288 2270 8300 2304
rect 7812 2264 8300 2270
rect 8830 2304 9318 2310
rect 8830 2270 8842 2304
rect 9306 2270 9318 2304
rect 8830 2264 9318 2270
rect 7012 2160 7072 2264
rect 8008 2160 8068 2264
rect 7006 2100 7012 2160
rect 7072 2100 7078 2160
rect 8002 2100 8008 2160
rect 8068 2100 8074 2160
rect 9546 2030 9606 2354
rect 10578 2354 10584 2866
rect 10618 2866 10632 2930
rect 11588 2930 11648 3170
rect 11588 2888 11602 2930
rect 10618 2354 10624 2866
rect 10578 2342 10624 2354
rect 11596 2354 11602 2888
rect 11636 2888 11648 2930
rect 11636 2354 11642 2888
rect 11596 2342 11642 2354
rect 9848 2304 10336 2310
rect 9848 2270 9860 2304
rect 10324 2270 10336 2304
rect 9848 2264 10336 2270
rect 10866 2304 11354 2310
rect 10866 2270 10878 2304
rect 11342 2270 11354 2304
rect 10866 2264 11354 2270
rect 11728 2030 11788 4346
rect 11848 3122 11908 5496
rect 11842 3062 11848 3122
rect 11908 3062 11914 3122
rect 5480 1970 5486 2030
rect 5546 1970 5552 2030
rect 9540 1970 9546 2030
rect 9606 1970 9612 2030
rect 11722 1970 11728 2030
rect 11788 1970 11794 2030
rect 1406 1964 1466 1970
rect 664 1564 11084 1624
rect 848 1388 908 1564
rect 1348 1478 1408 1564
rect 1144 1472 1632 1478
rect 1144 1438 1156 1472
rect 1620 1438 1632 1472
rect 1144 1432 1632 1438
rect 848 1354 862 1388
rect 856 812 862 1354
rect 896 1354 908 1388
rect 1870 1388 1930 1564
rect 2368 1478 2428 1564
rect 3402 1478 3462 1564
rect 4424 1478 4484 1564
rect 5414 1478 5474 1564
rect 2162 1472 2650 1478
rect 2162 1438 2174 1472
rect 2638 1438 2650 1472
rect 2162 1432 2650 1438
rect 3180 1472 3668 1478
rect 3180 1438 3192 1472
rect 3656 1438 3668 1472
rect 3180 1432 3668 1438
rect 4198 1472 4686 1478
rect 4198 1438 4210 1472
rect 4674 1438 4686 1472
rect 4198 1432 4686 1438
rect 5216 1472 5704 1478
rect 5216 1438 5228 1472
rect 5692 1438 5704 1472
rect 5216 1432 5704 1438
rect 896 812 902 1354
rect 1870 1344 1880 1388
rect 856 800 902 812
rect 1874 812 1880 1344
rect 1914 1344 1930 1388
rect 2892 1388 2938 1400
rect 1914 812 1920 1344
rect 2892 870 2898 1388
rect 1874 800 1920 812
rect 2884 812 2898 870
rect 2932 870 2938 1388
rect 3910 1388 3956 1400
rect 2932 812 2944 870
rect 3910 846 3916 1388
rect 1144 762 1632 768
rect 1144 728 1156 762
rect 1620 728 1632 762
rect 1144 722 1632 728
rect 2162 762 2650 768
rect 2162 728 2174 762
rect 2638 728 2650 762
rect 2162 722 2650 728
rect 2884 664 2944 812
rect 3902 812 3916 846
rect 3950 846 3956 1388
rect 4928 1388 4974 1400
rect 4928 858 4934 1388
rect 3950 812 3962 846
rect 3180 762 3668 768
rect 3180 728 3192 762
rect 3656 728 3668 762
rect 3180 722 3668 728
rect 2878 604 2884 664
rect 2944 604 2950 664
rect -1416 -576 -1304 210
rect 2884 110 2944 604
rect 3902 552 3962 812
rect 4922 812 4934 858
rect 4968 858 4974 1388
rect 5938 1388 5998 1564
rect 6448 1478 6508 1564
rect 7438 1478 7498 1564
rect 8470 1478 8530 1564
rect 9474 1478 9534 1564
rect 6234 1472 6722 1478
rect 6234 1438 6246 1472
rect 6710 1438 6722 1472
rect 6234 1432 6722 1438
rect 7252 1472 7740 1478
rect 7252 1438 7264 1472
rect 7728 1438 7740 1472
rect 7252 1432 7740 1438
rect 8270 1472 8758 1478
rect 8270 1438 8282 1472
rect 8746 1438 8758 1472
rect 8270 1432 8758 1438
rect 9288 1472 9776 1478
rect 9288 1438 9300 1472
rect 9764 1438 9776 1472
rect 9288 1432 9776 1438
rect 6448 1430 6508 1432
rect 8470 1430 8530 1432
rect 5938 1346 5952 1388
rect 4968 812 4982 858
rect 4198 762 4686 768
rect 4198 728 4210 762
rect 4674 728 4686 762
rect 4198 722 4686 728
rect 4922 664 4982 812
rect 5946 812 5952 1346
rect 5986 1346 5998 1388
rect 6964 1388 7010 1400
rect 5986 812 5992 1346
rect 6964 858 6970 1388
rect 5946 800 5992 812
rect 6958 812 6970 858
rect 7004 858 7010 1388
rect 7982 1388 8028 1400
rect 7004 812 7018 858
rect 7982 850 7988 1388
rect 5216 762 5704 768
rect 5216 728 5228 762
rect 5692 728 5704 762
rect 5216 722 5704 728
rect 6234 762 6722 768
rect 6234 728 6246 762
rect 6710 728 6722 762
rect 6234 722 6722 728
rect 6958 664 7018 812
rect 7976 812 7988 850
rect 8022 850 8028 1388
rect 9000 1388 9046 1400
rect 8022 812 8036 850
rect 9000 844 9006 1388
rect 7252 762 7740 768
rect 7252 728 7264 762
rect 7728 728 7740 762
rect 7252 722 7740 728
rect 4916 604 4922 664
rect 4982 604 4988 664
rect 6952 604 6958 664
rect 7018 604 7024 664
rect 3896 492 3902 552
rect 3962 492 3968 552
rect 4922 110 4982 604
rect 6958 110 7018 604
rect 7976 552 8036 812
rect 8994 812 9006 844
rect 9040 844 9046 1388
rect 10014 1388 10074 1564
rect 10494 1478 10554 1564
rect 10306 1472 10794 1478
rect 10306 1438 10318 1472
rect 10782 1438 10794 1472
rect 10306 1432 10794 1438
rect 10014 1320 10024 1388
rect 9040 812 9054 844
rect 8270 762 8758 768
rect 8270 728 8282 762
rect 8746 728 8758 762
rect 8270 722 8758 728
rect 8994 664 9054 812
rect 10018 812 10024 1320
rect 10058 1320 10074 1388
rect 11024 1388 11084 1564
rect 11024 1348 11042 1388
rect 10058 812 10064 1320
rect 10018 800 10064 812
rect 11036 812 11042 1348
rect 11076 1348 11084 1388
rect 11076 812 11082 1348
rect 11036 800 11082 812
rect 9288 762 9776 768
rect 9288 728 9300 762
rect 9764 728 9776 762
rect 9288 722 9776 728
rect 10306 762 10794 768
rect 10306 728 10318 762
rect 10782 728 10794 762
rect 10306 722 10794 728
rect 8988 604 8994 664
rect 9054 604 9060 664
rect 7970 492 7976 552
rect 8036 492 8042 552
rect 8994 110 9054 604
rect 11982 552 12042 7480
rect 12194 6646 12254 14986
rect 12188 6586 12194 6646
rect 12254 6586 12260 6646
rect 12314 6518 12374 14988
rect 12308 6458 12314 6518
rect 12374 6458 12380 6518
rect 12454 5556 12514 15006
rect 12566 14868 12572 14928
rect 12632 14868 12638 14928
rect 12572 8800 12632 14868
rect 12682 14186 12742 15022
rect 12676 14126 12682 14186
rect 12742 14126 12748 14186
rect 12800 11266 12860 15122
rect 13128 14320 13188 15132
rect 13122 14260 13128 14320
rect 13188 14260 13194 14320
rect 12918 12902 12924 12962
rect 12984 12902 12990 12962
rect 12798 11260 12860 11266
rect 12858 11200 12860 11260
rect 12798 11194 12860 11200
rect 12566 8740 12572 8800
rect 12632 8740 12638 8800
rect 12448 5496 12454 5556
rect 12514 5496 12520 5556
rect 12800 5198 12860 11194
rect 12924 10266 12984 12902
rect 13130 12566 13136 12626
rect 13196 12566 13202 12626
rect 13026 11306 13032 11366
rect 13092 11306 13098 11366
rect 12918 10206 12924 10266
rect 12984 10206 12990 10266
rect 13032 5348 13092 11306
rect 13136 10030 13196 12566
rect 13248 10144 13308 15124
rect 13354 15048 13414 15054
rect 13354 12504 13414 14988
rect 24160 14692 24166 14698
rect 13480 14638 24166 14692
rect 24226 14692 24232 14698
rect 29264 14692 29270 14698
rect 24226 14638 29270 14692
rect 29330 14692 29336 14698
rect 33330 14692 33390 14698
rect 29330 14638 33330 14692
rect 13480 14632 33330 14638
rect 33390 14632 33902 14692
rect 13480 14492 13540 14632
rect 14002 14582 14062 14632
rect 15012 14582 15072 14632
rect 13776 14576 14264 14582
rect 13776 14542 13788 14576
rect 14252 14542 14264 14576
rect 13776 14536 14264 14542
rect 14794 14576 15282 14582
rect 14794 14542 14806 14576
rect 15270 14542 15282 14576
rect 14794 14536 15282 14542
rect 15012 14530 15072 14536
rect 13480 13916 13494 14492
rect 13528 13916 13540 14492
rect 14506 14492 14552 14504
rect 14506 13950 14512 14492
rect 13480 13674 13540 13916
rect 14498 13916 14512 13950
rect 14546 13950 14552 14492
rect 15518 14492 15578 14632
rect 16042 14582 16102 14632
rect 17054 14582 17114 14632
rect 15812 14576 16300 14582
rect 15812 14542 15824 14576
rect 16288 14542 16300 14576
rect 15812 14536 16300 14542
rect 16830 14576 17318 14582
rect 16830 14542 16842 14576
rect 17306 14542 17318 14576
rect 16830 14536 17318 14542
rect 17054 14530 17114 14536
rect 14546 13916 14558 13950
rect 13776 13866 14264 13872
rect 13776 13832 13788 13866
rect 14252 13832 14264 13866
rect 13776 13826 14264 13832
rect 13992 13764 14052 13826
rect 13776 13758 14264 13764
rect 13776 13724 13788 13758
rect 14252 13724 14264 13758
rect 13776 13718 14264 13724
rect 13992 13712 14052 13718
rect 13480 13098 13494 13674
rect 13528 13098 13540 13674
rect 13480 12626 13540 13098
rect 14498 13674 14558 13916
rect 15518 13916 15530 14492
rect 15564 13916 15578 14492
rect 16542 14492 16588 14504
rect 16542 13962 16548 14492
rect 14998 13872 15058 13874
rect 14794 13866 15282 13872
rect 14794 13832 14806 13866
rect 15270 13832 15282 13866
rect 14794 13826 15282 13832
rect 14998 13764 15058 13826
rect 14794 13758 15282 13764
rect 14794 13724 14806 13758
rect 15270 13724 15282 13758
rect 14794 13718 15282 13724
rect 14498 13098 14512 13674
rect 14546 13098 14558 13674
rect 15518 13674 15578 13916
rect 16532 13916 16548 13962
rect 16582 13962 16588 14492
rect 17550 14492 17610 14632
rect 18066 14582 18126 14632
rect 19066 14582 19126 14632
rect 17848 14576 18336 14582
rect 17848 14542 17860 14576
rect 18324 14542 18336 14576
rect 17848 14536 18336 14542
rect 18866 14576 19354 14582
rect 18866 14542 18878 14576
rect 19342 14542 19354 14576
rect 18866 14536 19354 14542
rect 16582 13916 16592 13962
rect 16010 13872 16070 13880
rect 15812 13866 16300 13872
rect 15812 13832 15824 13866
rect 16288 13832 16300 13866
rect 15812 13826 16300 13832
rect 16010 13764 16070 13826
rect 15812 13758 16300 13764
rect 15812 13724 15824 13758
rect 16288 13724 16300 13758
rect 15812 13718 16300 13724
rect 15518 13616 15530 13674
rect 13776 13048 14264 13054
rect 13776 13014 13788 13048
rect 14252 13014 14264 13048
rect 13776 13008 14264 13014
rect 14498 12962 14558 13098
rect 15524 13098 15530 13616
rect 15564 13616 15578 13674
rect 16532 13674 16592 13916
rect 17550 13916 17566 14492
rect 17600 13916 17610 14492
rect 18578 14492 18624 14504
rect 18578 13956 18584 14492
rect 16830 13866 17318 13872
rect 16830 13832 16842 13866
rect 17306 13832 17318 13866
rect 16830 13826 17318 13832
rect 17032 13764 17092 13826
rect 16830 13758 17318 13764
rect 16830 13724 16842 13758
rect 17306 13724 17318 13758
rect 16830 13718 17318 13724
rect 17032 13712 17092 13718
rect 15564 13098 15570 13616
rect 15524 13086 15570 13098
rect 16532 13098 16548 13674
rect 16582 13098 16592 13674
rect 17550 13674 17610 13916
rect 18568 13916 18584 13956
rect 18618 13956 18624 14492
rect 19588 14492 19648 14632
rect 20100 14582 20160 14632
rect 21112 14582 21172 14632
rect 19884 14576 20372 14582
rect 19884 14542 19896 14576
rect 20360 14542 20372 14576
rect 19884 14536 20372 14542
rect 20902 14576 21390 14582
rect 20902 14542 20914 14576
rect 21378 14542 21390 14576
rect 20902 14536 21390 14542
rect 18618 13916 18628 13956
rect 17848 13866 18336 13872
rect 17848 13832 17860 13866
rect 18324 13832 18336 13866
rect 17848 13826 18336 13832
rect 18044 13764 18104 13826
rect 17848 13758 18336 13764
rect 17848 13724 17860 13758
rect 18324 13724 18336 13758
rect 17848 13718 18336 13724
rect 18044 13712 18104 13718
rect 17550 13612 17566 13674
rect 14794 13048 15282 13054
rect 14794 13014 14806 13048
rect 15270 13014 15282 13048
rect 14794 13008 15282 13014
rect 15812 13048 16300 13054
rect 15812 13014 15824 13048
rect 16288 13014 16300 13048
rect 15812 13008 16300 13014
rect 16532 12960 16592 13098
rect 17560 13098 17566 13612
rect 17600 13612 17610 13674
rect 18568 13674 18628 13916
rect 19588 13916 19602 14492
rect 19636 13916 19648 14492
rect 20614 14492 20660 14504
rect 20614 13956 20620 14492
rect 18866 13866 19354 13872
rect 18866 13832 18878 13866
rect 19342 13832 19354 13866
rect 18866 13826 19354 13832
rect 19074 13764 19134 13826
rect 18866 13758 19354 13764
rect 18866 13724 18878 13758
rect 19342 13724 19354 13758
rect 18866 13718 19354 13724
rect 19074 13712 19134 13718
rect 17600 13098 17606 13612
rect 17560 13086 17606 13098
rect 18568 13098 18584 13674
rect 18618 13098 18628 13674
rect 19588 13674 19648 13916
rect 20606 13916 20620 13956
rect 20654 13956 20660 14492
rect 21624 14492 21684 14632
rect 22136 14582 22196 14632
rect 23148 14582 23208 14632
rect 21920 14576 22408 14582
rect 21920 14542 21932 14576
rect 22396 14542 22408 14576
rect 21920 14536 22408 14542
rect 22938 14576 23426 14582
rect 22938 14542 22950 14576
rect 23414 14542 23426 14576
rect 22938 14536 23426 14542
rect 20654 13916 20666 13956
rect 20080 13872 20140 13874
rect 19884 13866 20372 13872
rect 19884 13832 19896 13866
rect 20360 13832 20372 13866
rect 19884 13826 20372 13832
rect 20080 13764 20140 13826
rect 19884 13758 20372 13764
rect 19884 13724 19896 13758
rect 20360 13724 20372 13758
rect 19884 13718 20372 13724
rect 19588 13632 19602 13674
rect 16830 13048 17318 13054
rect 16830 13014 16842 13048
rect 17306 13014 17318 13048
rect 16830 13008 17318 13014
rect 17848 13048 18336 13054
rect 17848 13014 17860 13048
rect 18324 13014 18336 13048
rect 17848 13008 18336 13014
rect 18568 12960 18628 13098
rect 19596 13098 19602 13632
rect 19636 13632 19648 13674
rect 20606 13674 20666 13916
rect 21624 13916 21638 14492
rect 21672 13916 21684 14492
rect 22650 14492 22696 14504
rect 22650 13962 22656 14492
rect 21102 13872 21162 13874
rect 20902 13866 21390 13872
rect 20902 13832 20914 13866
rect 21378 13832 21390 13866
rect 20902 13826 21390 13832
rect 21102 13764 21162 13826
rect 20902 13758 21390 13764
rect 20902 13724 20914 13758
rect 21378 13724 21390 13758
rect 20902 13718 21390 13724
rect 19636 13098 19642 13632
rect 19596 13086 19642 13098
rect 20606 13098 20620 13674
rect 20654 13098 20666 13674
rect 21624 13674 21684 13916
rect 22644 13916 22656 13962
rect 22690 13962 22696 14492
rect 23656 14492 23716 14632
rect 24170 14582 24230 14632
rect 25182 14582 25242 14632
rect 23956 14576 24444 14582
rect 23956 14542 23968 14576
rect 24432 14542 24444 14576
rect 23956 14536 24444 14542
rect 24974 14576 25462 14582
rect 24974 14542 24986 14576
rect 25450 14542 25462 14576
rect 24974 14536 25462 14542
rect 25182 14530 25242 14536
rect 22690 13916 22704 13962
rect 21920 13866 22408 13872
rect 21920 13832 21932 13866
rect 22396 13832 22408 13866
rect 21920 13826 22408 13832
rect 22126 13764 22186 13826
rect 21920 13758 22408 13764
rect 21920 13724 21932 13758
rect 22396 13724 22408 13758
rect 21920 13718 22408 13724
rect 22126 13712 22186 13718
rect 21624 13624 21638 13674
rect 18866 13048 19354 13054
rect 18866 13014 18878 13048
rect 19342 13014 19354 13048
rect 18866 13008 19354 13014
rect 19884 13048 20372 13054
rect 19884 13014 19896 13048
rect 20360 13014 20372 13048
rect 19884 13008 20372 13014
rect 20606 12960 20666 13098
rect 21632 13098 21638 13624
rect 21672 13624 21684 13674
rect 22644 13674 22704 13916
rect 23656 13916 23674 14492
rect 23708 13916 23716 14492
rect 24686 14492 24732 14504
rect 24686 13962 24692 14492
rect 23132 13872 23192 13874
rect 22938 13866 23426 13872
rect 22938 13832 22950 13866
rect 23414 13832 23426 13866
rect 22938 13826 23426 13832
rect 23132 13764 23192 13826
rect 22938 13758 23426 13764
rect 22938 13724 22950 13758
rect 23414 13724 23426 13758
rect 22938 13718 23426 13724
rect 21672 13098 21678 13624
rect 21632 13086 21678 13098
rect 22644 13098 22656 13674
rect 22690 13098 22704 13674
rect 23656 13674 23716 13916
rect 24678 13916 24692 13962
rect 24726 13962 24732 14492
rect 25694 14492 25754 14632
rect 26206 14582 26266 14632
rect 27224 14582 27284 14632
rect 25992 14576 26480 14582
rect 25992 14542 26004 14576
rect 26468 14542 26480 14576
rect 25992 14536 26480 14542
rect 27010 14576 27498 14582
rect 27010 14542 27022 14576
rect 27486 14542 27498 14576
rect 27010 14536 27498 14542
rect 26206 14530 26266 14536
rect 24726 13916 24738 13962
rect 24156 13872 24216 13880
rect 23956 13866 24444 13872
rect 23956 13832 23968 13866
rect 24432 13832 24444 13866
rect 23956 13826 24444 13832
rect 24156 13764 24216 13826
rect 23956 13758 24444 13764
rect 23956 13724 23968 13758
rect 24432 13724 24444 13758
rect 23956 13718 24444 13724
rect 23656 13626 23674 13674
rect 20902 13048 21390 13054
rect 20902 13014 20914 13048
rect 21378 13014 21390 13048
rect 20902 13008 21390 13014
rect 21920 13048 22408 13054
rect 21920 13014 21932 13048
rect 22396 13014 22408 13048
rect 21920 13008 22408 13014
rect 22644 12960 22704 13098
rect 23668 13098 23674 13626
rect 23708 13626 23716 13674
rect 24678 13674 24738 13916
rect 25694 13916 25710 14492
rect 25744 13916 25754 14492
rect 26722 14492 26768 14504
rect 26722 13962 26728 14492
rect 25178 13872 25238 13874
rect 24974 13866 25462 13872
rect 24974 13832 24986 13866
rect 25450 13832 25462 13866
rect 24974 13826 25462 13832
rect 25178 13764 25238 13826
rect 24974 13758 25462 13764
rect 24974 13724 24986 13758
rect 25450 13724 25462 13758
rect 24974 13718 25462 13724
rect 23708 13098 23714 13626
rect 23668 13086 23714 13098
rect 24678 13098 24692 13674
rect 24726 13098 24738 13674
rect 25694 13674 25754 13916
rect 26714 13916 26728 13962
rect 26762 13962 26768 14492
rect 27730 14492 27790 14632
rect 28246 14582 28306 14632
rect 29270 14582 29330 14632
rect 28028 14576 28516 14582
rect 28028 14542 28040 14576
rect 28504 14542 28516 14576
rect 28028 14536 28516 14542
rect 29046 14576 29534 14582
rect 29046 14542 29058 14576
rect 29522 14542 29534 14576
rect 29046 14536 29534 14542
rect 26762 13916 26774 13962
rect 26190 13872 26250 13874
rect 25992 13866 26480 13872
rect 25992 13832 26004 13866
rect 26468 13832 26480 13866
rect 25992 13826 26480 13832
rect 26190 13764 26250 13826
rect 25992 13758 26480 13764
rect 25992 13724 26004 13758
rect 26468 13724 26480 13758
rect 25992 13718 26480 13724
rect 25694 13624 25710 13674
rect 22938 13048 23426 13054
rect 22938 13014 22950 13048
rect 23414 13014 23426 13048
rect 22938 13008 23426 13014
rect 23956 13048 24444 13054
rect 23956 13014 23968 13048
rect 24432 13014 24444 13048
rect 23956 13008 24444 13014
rect 24678 12960 24738 13098
rect 25704 13098 25710 13624
rect 25744 13624 25754 13674
rect 26714 13674 26774 13916
rect 27730 13916 27746 14492
rect 27780 13916 27790 14492
rect 28758 14492 28804 14504
rect 28758 13986 28764 14492
rect 27010 13866 27498 13872
rect 27010 13832 27022 13866
rect 27486 13832 27498 13866
rect 27010 13826 27498 13832
rect 27202 13764 27262 13826
rect 27010 13758 27498 13764
rect 27010 13724 27022 13758
rect 27486 13724 27498 13758
rect 27010 13718 27498 13724
rect 27202 13712 27262 13718
rect 25744 13098 25750 13624
rect 25704 13086 25750 13098
rect 26714 13098 26728 13674
rect 26762 13098 26774 13674
rect 27730 13674 27790 13916
rect 28752 13916 28764 13986
rect 28798 13986 28804 14492
rect 29766 14492 29826 14632
rect 30288 14582 30348 14632
rect 31300 14582 31360 14632
rect 30064 14576 30552 14582
rect 30064 14542 30076 14576
rect 30540 14542 30552 14576
rect 30064 14536 30552 14542
rect 31082 14576 31570 14582
rect 31082 14542 31094 14576
rect 31558 14542 31570 14576
rect 31082 14536 31570 14542
rect 28798 13916 28812 13986
rect 28226 13872 28286 13880
rect 28028 13866 28516 13872
rect 28028 13832 28040 13866
rect 28504 13832 28516 13866
rect 28028 13826 28516 13832
rect 28226 13764 28286 13826
rect 28028 13758 28516 13764
rect 28028 13724 28040 13758
rect 28504 13724 28516 13758
rect 28028 13718 28516 13724
rect 27730 13650 27746 13674
rect 24974 13048 25462 13054
rect 24974 13014 24986 13048
rect 25450 13014 25462 13048
rect 24974 13008 25462 13014
rect 25992 13048 26480 13054
rect 25992 13014 26004 13048
rect 26468 13014 26480 13048
rect 25992 13008 26480 13014
rect 26714 12960 26774 13098
rect 27740 13098 27746 13650
rect 27780 13650 27790 13674
rect 28752 13674 28812 13916
rect 29766 13916 29782 14492
rect 29816 13916 29826 14492
rect 30794 14492 30840 14504
rect 30794 14026 30800 14492
rect 29046 13866 29534 13872
rect 29046 13832 29058 13866
rect 29522 13832 29534 13866
rect 29046 13826 29534 13832
rect 29248 13764 29308 13826
rect 29046 13758 29534 13764
rect 29046 13724 29058 13758
rect 29522 13724 29534 13758
rect 29046 13718 29534 13724
rect 29248 13706 29308 13718
rect 27780 13098 27786 13650
rect 27740 13086 27786 13098
rect 28752 13098 28764 13674
rect 28798 13098 28812 13674
rect 29766 13674 29826 13916
rect 30786 13916 30800 14026
rect 30834 14026 30840 14492
rect 31804 14492 31864 14632
rect 32310 14582 32370 14632
rect 33328 14626 33390 14632
rect 33328 14582 33388 14626
rect 32100 14576 32588 14582
rect 32100 14542 32112 14576
rect 32576 14542 32588 14576
rect 32100 14536 32588 14542
rect 33118 14576 33606 14582
rect 33118 14542 33130 14576
rect 33594 14542 33606 14576
rect 33118 14536 33606 14542
rect 30834 13916 30846 14026
rect 30266 13872 30326 13874
rect 30064 13866 30552 13872
rect 30064 13832 30076 13866
rect 30540 13832 30552 13866
rect 30064 13826 30552 13832
rect 30266 13764 30326 13826
rect 30064 13758 30552 13764
rect 30064 13724 30076 13758
rect 30540 13724 30552 13758
rect 30064 13718 30552 13724
rect 29766 13632 29782 13674
rect 27010 13048 27498 13054
rect 27010 13014 27022 13048
rect 27486 13014 27498 13048
rect 27010 13008 27498 13014
rect 28028 13048 28516 13054
rect 28028 13014 28040 13048
rect 28504 13014 28516 13048
rect 28028 13008 28516 13014
rect 28752 12960 28812 13098
rect 29776 13098 29782 13632
rect 29816 13632 29826 13674
rect 30786 13674 30846 13916
rect 31804 13916 31818 14492
rect 31852 13916 31864 14492
rect 32830 14492 32876 14504
rect 32830 13976 32836 14492
rect 31296 13872 31356 13886
rect 31082 13866 31570 13872
rect 31082 13832 31094 13866
rect 31558 13832 31570 13866
rect 31082 13826 31570 13832
rect 31296 13764 31356 13826
rect 31082 13758 31570 13764
rect 31082 13724 31094 13758
rect 31558 13724 31570 13758
rect 31082 13718 31570 13724
rect 29816 13098 29822 13632
rect 29776 13086 29822 13098
rect 30786 13098 30800 13674
rect 30834 13098 30846 13674
rect 31804 13674 31864 13916
rect 32822 13916 32836 13976
rect 32870 13976 32876 14492
rect 33842 14492 33902 14632
rect 32870 13916 32882 13976
rect 32308 13872 32368 13886
rect 32100 13866 32588 13872
rect 32100 13832 32112 13866
rect 32576 13832 32588 13866
rect 32100 13826 32588 13832
rect 32308 13764 32368 13826
rect 32100 13758 32588 13764
rect 32100 13724 32112 13758
rect 32576 13724 32588 13758
rect 32100 13718 32588 13724
rect 31804 13632 31818 13674
rect 29046 13048 29534 13054
rect 29046 13014 29058 13048
rect 29522 13014 29534 13048
rect 29046 13008 29534 13014
rect 30064 13048 30552 13054
rect 30064 13014 30076 13048
rect 30540 13014 30552 13048
rect 30064 13008 30552 13014
rect 30786 12960 30846 13098
rect 31812 13098 31818 13632
rect 31852 13632 31864 13674
rect 32822 13674 32882 13916
rect 33842 13916 33854 14492
rect 33888 13916 33902 14492
rect 33118 13866 33606 13872
rect 33118 13832 33130 13866
rect 33594 13832 33606 13866
rect 33118 13826 33606 13832
rect 33308 13764 33368 13826
rect 33842 13824 33902 13916
rect 35728 14470 35840 15256
rect 33842 13764 34622 13824
rect 33118 13758 33606 13764
rect 33118 13724 33130 13758
rect 33594 13724 33606 13758
rect 33118 13718 33606 13724
rect 33308 13712 33368 13718
rect 31852 13098 31858 13632
rect 31812 13086 31858 13098
rect 32822 13098 32836 13674
rect 32870 13098 32882 13674
rect 33842 13674 33902 13764
rect 33842 13624 33854 13674
rect 31082 13048 31570 13054
rect 31082 13014 31094 13048
rect 31558 13014 31570 13048
rect 31082 13008 31570 13014
rect 32100 13048 32588 13054
rect 32100 13014 32112 13048
rect 32576 13014 32588 13048
rect 32100 13008 32588 13014
rect 32822 12960 32882 13098
rect 33848 13098 33854 13624
rect 33888 13624 33902 13674
rect 33888 13098 33894 13624
rect 33848 13086 33894 13098
rect 33118 13048 33606 13054
rect 33118 13014 33130 13048
rect 33594 13014 33606 13048
rect 33118 13008 33606 13014
rect 14558 12902 34500 12960
rect 14498 12900 34500 12902
rect 14498 12896 14558 12900
rect 15506 12686 15512 12746
rect 15572 12686 15578 12746
rect 17546 12686 17552 12746
rect 17612 12686 17618 12746
rect 19586 12686 19592 12746
rect 19652 12686 19658 12746
rect 21616 12686 21622 12746
rect 21682 12686 21688 12746
rect 23656 12686 23662 12746
rect 23722 12686 23728 12746
rect 25688 12686 25694 12746
rect 25754 12686 25760 12746
rect 27728 12686 27734 12746
rect 27794 12686 27800 12746
rect 29764 12686 29770 12746
rect 29830 12686 29836 12746
rect 31798 12686 31804 12746
rect 31864 12686 31870 12746
rect 13474 12566 13480 12626
rect 13540 12566 13546 12626
rect 14998 12560 15004 12620
rect 15064 12560 15070 12620
rect 13348 12444 13354 12504
rect 13414 12444 13420 12504
rect 13354 10370 13414 12444
rect 15004 12386 15064 12560
rect 13776 12380 14264 12386
rect 13776 12346 13788 12380
rect 14252 12346 14264 12380
rect 13776 12340 14264 12346
rect 14794 12380 15282 12386
rect 14794 12346 14806 12380
rect 15270 12346 15282 12380
rect 14794 12340 15282 12346
rect 13488 12296 13534 12308
rect 14506 12296 14552 12308
rect 15512 12296 15572 12686
rect 16018 12620 16078 12626
rect 16018 12386 16078 12560
rect 17040 12620 17100 12626
rect 17040 12386 17100 12560
rect 15812 12380 16300 12386
rect 15812 12346 15824 12380
rect 16288 12346 16300 12380
rect 15812 12340 16300 12346
rect 16830 12380 17318 12386
rect 16830 12346 16842 12380
rect 17306 12346 17318 12380
rect 16830 12340 17318 12346
rect 16542 12296 16588 12308
rect 13480 12262 13494 12296
rect 13488 11770 13494 12262
rect 13480 11720 13494 11770
rect 13528 12262 13540 12296
rect 13528 11770 13534 12262
rect 14498 12248 14512 12296
rect 13528 11720 13540 11770
rect 14506 11756 14512 12248
rect 13480 11582 13540 11720
rect 14498 11720 14512 11756
rect 14546 12248 14558 12296
rect 14546 11756 14552 12248
rect 15512 12228 15530 12296
rect 15524 11784 15530 12228
rect 14546 11720 14558 11756
rect 13776 11670 14264 11676
rect 13776 11636 13788 11670
rect 14252 11636 14264 11670
rect 13776 11630 14264 11636
rect 13982 11582 14042 11630
rect 14498 11582 14558 11720
rect 15516 11720 15530 11784
rect 15564 12264 15576 12296
rect 15564 12228 15572 12264
rect 15564 11784 15570 12228
rect 15564 11720 15576 11784
rect 16542 11766 16548 12296
rect 16538 11748 16548 11766
rect 16536 11720 16548 11748
rect 16582 11766 16588 12296
rect 17552 12296 17612 12686
rect 18054 12620 18114 12626
rect 18052 12560 18054 12566
rect 19080 12620 19140 12626
rect 18052 12554 18114 12560
rect 19078 12560 19080 12566
rect 19078 12554 19140 12560
rect 18052 12386 18112 12554
rect 18562 12444 18568 12504
rect 18628 12444 18634 12504
rect 17848 12380 18336 12386
rect 17848 12346 17860 12380
rect 18324 12346 18336 12380
rect 17848 12340 18336 12346
rect 17552 12242 17566 12296
rect 17560 11792 17566 12242
rect 17556 11768 17566 11792
rect 16582 11720 16598 11766
rect 17554 11720 17566 11768
rect 17600 12242 17612 12296
rect 18568 12296 18628 12444
rect 19078 12386 19138 12554
rect 18866 12380 19354 12386
rect 18866 12346 18878 12380
rect 19342 12346 19354 12380
rect 18866 12340 19354 12346
rect 18568 12254 18584 12296
rect 17600 11792 17606 12242
rect 18578 11796 18584 12254
rect 17600 11720 17616 11792
rect 18568 11720 18584 11796
rect 18618 12254 18628 12296
rect 19592 12296 19652 12686
rect 20092 12620 20152 12626
rect 20092 12386 20152 12560
rect 21128 12620 21188 12626
rect 21128 12386 21188 12560
rect 19884 12380 20372 12386
rect 19884 12346 19896 12380
rect 20360 12346 20372 12380
rect 19884 12340 20372 12346
rect 20902 12380 21390 12386
rect 20902 12346 20914 12380
rect 21378 12346 21390 12380
rect 20902 12340 21390 12346
rect 20614 12296 20660 12308
rect 21622 12296 21682 12686
rect 22134 12620 22194 12626
rect 23142 12560 23148 12620
rect 23208 12560 23214 12620
rect 22134 12386 22194 12560
rect 23148 12386 23208 12560
rect 21920 12380 22408 12386
rect 21920 12346 21932 12380
rect 22396 12346 22408 12380
rect 21920 12340 22408 12346
rect 22938 12380 23426 12386
rect 22938 12346 22950 12380
rect 23414 12346 23426 12380
rect 22938 12340 23426 12346
rect 18618 11796 18624 12254
rect 19592 12222 19602 12296
rect 18618 11780 18628 11796
rect 18618 11720 18632 11780
rect 19596 11776 19602 12222
rect 19588 11720 19602 11776
rect 19636 12222 19652 12296
rect 20608 12246 20620 12296
rect 19636 11776 19642 12222
rect 20614 11784 20620 12246
rect 19636 11720 19648 11776
rect 20608 11756 20620 11784
rect 20606 11720 20620 11756
rect 20654 12246 20668 12296
rect 20654 11784 20660 12246
rect 21622 12228 21638 12296
rect 21632 11796 21638 12228
rect 20654 11720 20668 11784
rect 14794 11670 15282 11676
rect 14794 11636 14806 11670
rect 15270 11636 15282 11670
rect 14794 11630 15282 11636
rect 13480 11522 14558 11582
rect 14498 11366 14558 11522
rect 15008 11472 15068 11630
rect 15516 11582 15576 11720
rect 15812 11670 16300 11676
rect 15812 11636 15824 11670
rect 16288 11636 16300 11670
rect 15812 11630 16300 11636
rect 15510 11522 15516 11582
rect 15576 11522 15582 11582
rect 15002 11412 15008 11472
rect 15068 11412 15074 11472
rect 14492 11306 14498 11366
rect 14558 11306 14564 11366
rect 13478 11200 13484 11260
rect 13544 11200 13550 11260
rect 13976 11200 13982 11260
rect 14042 11200 14048 11260
rect 14488 11200 14494 11260
rect 14554 11200 14560 11260
rect 13484 11064 13544 11200
rect 13982 11154 14042 11200
rect 13776 11148 14264 11154
rect 13776 11114 13788 11148
rect 14252 11114 14264 11148
rect 13776 11108 14264 11114
rect 13484 11024 13494 11064
rect 13488 10488 13494 11024
rect 13528 11024 13544 11064
rect 14494 11064 14554 11200
rect 15008 11154 15068 11412
rect 14794 11148 15282 11154
rect 14794 11114 14806 11148
rect 15270 11114 15282 11148
rect 14794 11108 15282 11114
rect 13528 10488 13534 11024
rect 14494 11018 14512 11064
rect 13488 10476 13534 10488
rect 14506 10488 14512 11018
rect 14546 11018 14554 11064
rect 15516 11064 15576 11522
rect 16030 11472 16090 11630
rect 16024 11412 16030 11472
rect 16090 11412 16096 11472
rect 16030 11154 16090 11412
rect 16538 11366 16598 11720
rect 16830 11670 17318 11676
rect 16830 11636 16842 11670
rect 17306 11636 17318 11670
rect 16830 11630 17318 11636
rect 17044 11472 17104 11630
rect 17556 11582 17616 11720
rect 18578 11708 18624 11720
rect 17848 11670 18336 11676
rect 17848 11636 17860 11670
rect 18324 11636 18336 11670
rect 17848 11630 18336 11636
rect 18866 11670 19354 11676
rect 18866 11636 18878 11670
rect 19342 11636 19354 11670
rect 18866 11630 19354 11636
rect 17550 11522 17556 11582
rect 17616 11522 17622 11582
rect 17038 11412 17044 11472
rect 17104 11412 17110 11472
rect 16532 11306 16538 11366
rect 16598 11306 16604 11366
rect 17044 11154 17104 11412
rect 15812 11148 16300 11154
rect 15812 11114 15824 11148
rect 16288 11114 16300 11148
rect 15812 11108 16300 11114
rect 16830 11148 17318 11154
rect 16830 11114 16842 11148
rect 17306 11114 17318 11148
rect 16830 11108 17318 11114
rect 16542 11064 16588 11076
rect 17556 11064 17616 11522
rect 18058 11472 18118 11630
rect 19076 11472 19136 11630
rect 19588 11582 19648 11720
rect 19884 11670 20372 11676
rect 19884 11636 19896 11670
rect 20360 11636 20372 11670
rect 19884 11630 20372 11636
rect 19582 11522 19588 11582
rect 19648 11522 19654 11582
rect 18052 11412 18058 11472
rect 18118 11412 18124 11472
rect 19070 11412 19076 11472
rect 19136 11412 19142 11472
rect 18058 11154 18118 11412
rect 18562 11306 18568 11366
rect 18628 11306 18634 11366
rect 17848 11148 18336 11154
rect 17848 11114 17860 11148
rect 18324 11114 18336 11148
rect 17848 11108 18336 11114
rect 15516 11026 15530 11064
rect 14546 10488 14552 11018
rect 15524 10546 15530 11026
rect 14506 10476 14552 10488
rect 15510 10488 15530 10546
rect 15564 11026 15576 11064
rect 15564 10488 15570 11026
rect 16536 11012 16548 11064
rect 16542 10508 16548 11012
rect 13776 10438 14264 10444
rect 13776 10404 13788 10438
rect 14252 10404 14264 10438
rect 13776 10398 14264 10404
rect 14794 10438 15282 10444
rect 14794 10404 14806 10438
rect 15270 10404 15282 10438
rect 14794 10398 15282 10404
rect 13348 10310 13354 10370
rect 13414 10310 13420 10370
rect 15510 10266 15570 10488
rect 16532 10488 16548 10508
rect 16582 11012 16596 11064
rect 16582 10508 16588 11012
rect 17554 11000 17566 11064
rect 17560 10552 17566 11000
rect 16582 10488 16592 10508
rect 15812 10438 16300 10444
rect 15812 10404 15824 10438
rect 16288 10404 16300 10438
rect 15812 10398 16300 10404
rect 13472 10206 13478 10266
rect 13538 10206 13544 10266
rect 14992 10206 14998 10266
rect 15058 10206 15064 10266
rect 15504 10206 15510 10266
rect 15570 10206 15576 10266
rect 13242 10084 13248 10144
rect 13308 10084 13314 10144
rect 13130 9970 13136 10030
rect 13196 9970 13202 10030
rect 13248 8902 13308 10084
rect 13478 9830 13538 10206
rect 13978 9970 13984 10030
rect 14044 9970 14050 10030
rect 13984 9920 14044 9970
rect 14998 9920 15058 10206
rect 15510 9972 15516 10032
rect 15576 9972 15582 10032
rect 13774 9914 14262 9920
rect 13774 9880 13786 9914
rect 14250 9880 14262 9914
rect 13774 9874 14262 9880
rect 14792 9914 15280 9920
rect 14792 9880 14804 9914
rect 15268 9880 15280 9914
rect 14792 9874 15280 9880
rect 14504 9830 14550 9842
rect 15516 9830 15576 9972
rect 16014 9920 16074 10398
rect 16532 10370 16592 10488
rect 17546 10488 17566 10552
rect 17600 11030 17616 11064
rect 18568 11064 18628 11306
rect 19076 11154 19136 11412
rect 18866 11148 19354 11154
rect 18866 11114 18878 11148
rect 19342 11114 19354 11148
rect 18866 11108 19354 11114
rect 19588 11064 19648 11522
rect 20102 11472 20162 11630
rect 20608 11512 20668 11720
rect 21620 11720 21638 11796
rect 21672 12228 21682 12296
rect 22650 12296 22696 12308
rect 21672 11796 21678 12228
rect 21672 11720 21680 11796
rect 22650 11782 22656 12296
rect 22644 11780 22656 11782
rect 20902 11670 21390 11676
rect 20902 11636 20914 11670
rect 21378 11636 21390 11670
rect 20902 11630 21390 11636
rect 20096 11412 20102 11472
rect 20162 11412 20168 11472
rect 20608 11452 20834 11512
rect 21122 11472 21182 11630
rect 21620 11582 21680 11720
rect 22642 11720 22656 11780
rect 22690 11782 22696 12296
rect 23662 12296 23722 12686
rect 24164 12620 24224 12626
rect 24164 12386 24224 12560
rect 25172 12620 25232 12626
rect 25232 12560 25234 12566
rect 25172 12554 25234 12560
rect 25174 12386 25234 12554
rect 23956 12380 24444 12386
rect 23956 12346 23968 12380
rect 24432 12346 24444 12380
rect 23956 12340 24444 12346
rect 24974 12380 25462 12386
rect 24974 12346 24986 12380
rect 25450 12346 25462 12380
rect 24974 12340 25462 12346
rect 24686 12296 24732 12308
rect 25694 12296 25754 12686
rect 26188 12620 26248 12626
rect 27212 12620 27272 12626
rect 26248 12560 26250 12566
rect 26188 12554 26250 12560
rect 26190 12386 26250 12554
rect 27212 12386 27272 12560
rect 25992 12380 26480 12386
rect 25992 12346 26004 12380
rect 26468 12346 26480 12380
rect 25992 12340 26480 12346
rect 27010 12380 27498 12386
rect 27010 12346 27022 12380
rect 27486 12346 27498 12380
rect 27010 12340 27498 12346
rect 26722 12296 26768 12308
rect 27734 12296 27794 12686
rect 28234 12620 28294 12626
rect 29256 12620 29316 12626
rect 28234 12386 28294 12560
rect 29254 12560 29256 12566
rect 29254 12554 29316 12560
rect 28750 12444 28756 12504
rect 28816 12444 28822 12504
rect 28028 12380 28516 12386
rect 28028 12346 28040 12380
rect 28504 12346 28516 12380
rect 28028 12340 28516 12346
rect 23662 12228 23674 12296
rect 23668 11786 23674 12228
rect 22690 11720 22704 11782
rect 23656 11720 23674 11786
rect 23708 12228 23722 12296
rect 24676 12262 24692 12296
rect 23708 11786 23714 12228
rect 23708 11720 23716 11786
rect 24686 11768 24692 12262
rect 21920 11670 22408 11676
rect 21920 11636 21932 11670
rect 22396 11636 22408 11670
rect 21920 11630 22408 11636
rect 21614 11522 21620 11582
rect 21680 11522 21686 11582
rect 20102 11154 20162 11412
rect 20602 11306 20608 11366
rect 20668 11306 20674 11366
rect 19884 11148 20372 11154
rect 19884 11114 19896 11148
rect 20360 11114 20372 11148
rect 19884 11108 20372 11114
rect 20608 11064 20668 11306
rect 20774 11260 20834 11452
rect 21116 11412 21122 11472
rect 21182 11412 21188 11472
rect 20768 11200 20774 11260
rect 20834 11200 20840 11260
rect 21122 11154 21182 11412
rect 20902 11148 21390 11154
rect 20902 11114 20914 11148
rect 21378 11114 21390 11148
rect 20902 11108 21390 11114
rect 17600 11000 17614 11030
rect 18568 11020 18584 11064
rect 17600 10488 17606 11000
rect 16830 10438 17318 10444
rect 16830 10404 16842 10438
rect 17306 10404 17318 10438
rect 16830 10398 17318 10404
rect 16526 10310 16532 10370
rect 16592 10310 16598 10370
rect 16528 10206 16534 10266
rect 16594 10206 16600 10266
rect 15810 9914 16298 9920
rect 15810 9880 15822 9914
rect 16286 9880 16298 9914
rect 15810 9874 16298 9880
rect 13478 9774 13492 9830
rect 13486 9254 13492 9774
rect 13526 9774 13538 9830
rect 14498 9798 14510 9830
rect 13526 9254 13532 9774
rect 14504 9298 14510 9798
rect 13486 9242 13532 9254
rect 14498 9254 14510 9298
rect 14544 9798 14558 9830
rect 15516 9804 15528 9830
rect 14544 9298 14550 9798
rect 14544 9254 14558 9298
rect 13774 9204 14262 9210
rect 13774 9170 13786 9204
rect 14250 9170 14262 9204
rect 13774 9164 14262 9170
rect 14498 9102 14558 9254
rect 15522 9254 15528 9804
rect 15562 9804 15576 9830
rect 16534 9830 16594 10206
rect 17034 9920 17094 10398
rect 17546 10266 17606 10488
rect 18578 10488 18584 11020
rect 18618 11030 18630 11064
rect 18618 11020 18628 11030
rect 19588 11022 19602 11064
rect 18618 10488 18624 11020
rect 19596 10530 19602 11022
rect 19588 10488 19602 10530
rect 19636 11022 19648 11064
rect 19636 10530 19642 11022
rect 20604 11002 20620 11064
rect 19636 10488 19648 10530
rect 20614 10488 20620 11002
rect 20654 11024 20668 11064
rect 21620 11064 21680 11522
rect 22142 11472 22202 11630
rect 22136 11412 22142 11472
rect 22202 11412 22208 11472
rect 22142 11154 22202 11412
rect 22642 11366 22702 11720
rect 22938 11670 23426 11676
rect 22938 11636 22950 11670
rect 23414 11636 23426 11670
rect 22938 11630 23426 11636
rect 23144 11472 23204 11630
rect 23656 11582 23716 11720
rect 24678 11720 24692 11768
rect 24726 12262 24736 12296
rect 24726 11768 24732 12262
rect 25694 12242 25710 12296
rect 25704 11780 25710 12242
rect 24726 11720 24738 11768
rect 23956 11670 24444 11676
rect 23956 11636 23968 11670
rect 24432 11636 24444 11670
rect 23956 11630 24444 11636
rect 23650 11522 23656 11582
rect 23716 11522 23722 11582
rect 23138 11412 23144 11472
rect 23204 11412 23210 11472
rect 22636 11306 22642 11366
rect 22702 11306 22708 11366
rect 22636 11200 22642 11260
rect 22702 11200 22708 11260
rect 21920 11148 22408 11154
rect 21920 11114 21932 11148
rect 22396 11114 22408 11148
rect 21920 11108 22408 11114
rect 22642 11064 22702 11200
rect 23144 11154 23204 11412
rect 22938 11148 23426 11154
rect 22938 11114 22950 11148
rect 23414 11114 23426 11148
rect 22938 11108 23426 11114
rect 23656 11064 23716 11522
rect 24170 11472 24230 11630
rect 24164 11412 24170 11472
rect 24230 11412 24236 11472
rect 24170 11154 24230 11412
rect 24678 11366 24738 11720
rect 25692 11720 25710 11780
rect 25744 12242 25754 12296
rect 26714 12256 26728 12296
rect 25744 11780 25750 12242
rect 26722 11786 26728 12256
rect 25744 11720 25752 11780
rect 26718 11760 26728 11786
rect 24974 11670 25462 11676
rect 24974 11636 24986 11670
rect 25450 11636 25462 11670
rect 24974 11630 25462 11636
rect 25188 11472 25248 11630
rect 25692 11582 25752 11720
rect 26716 11720 26728 11760
rect 26762 12256 26774 12296
rect 26762 11786 26768 12256
rect 27734 12242 27746 12296
rect 26762 11720 26778 11786
rect 27740 11770 27746 12242
rect 27730 11720 27746 11770
rect 27780 12242 27794 12296
rect 28756 12296 28816 12444
rect 29254 12386 29314 12554
rect 29046 12380 29534 12386
rect 29046 12346 29058 12380
rect 29522 12346 29534 12380
rect 29046 12340 29534 12346
rect 27780 11770 27786 12242
rect 28756 12232 28764 12296
rect 28758 11776 28764 12232
rect 27780 11720 27790 11770
rect 28750 11720 28764 11776
rect 28798 12232 28816 12296
rect 29770 12296 29830 12686
rect 30274 12620 30334 12626
rect 31288 12620 31348 12626
rect 30334 12560 30336 12566
rect 30274 12554 30336 12560
rect 31348 12560 31350 12566
rect 31288 12554 31350 12560
rect 30276 12386 30336 12554
rect 31290 12386 31350 12554
rect 30064 12380 30552 12386
rect 30064 12346 30076 12380
rect 30540 12346 30552 12380
rect 30064 12340 30552 12346
rect 31082 12380 31570 12386
rect 31082 12346 31094 12380
rect 31558 12346 31570 12380
rect 31082 12340 31570 12346
rect 30794 12296 30840 12308
rect 31804 12296 31864 12686
rect 32312 12620 32372 12626
rect 32310 12560 32312 12566
rect 32310 12554 32372 12560
rect 32310 12386 32370 12554
rect 32822 12444 32828 12504
rect 32888 12444 32894 12504
rect 33954 12444 33960 12504
rect 34020 12444 34026 12504
rect 32100 12380 32588 12386
rect 32100 12346 32112 12380
rect 32576 12346 32588 12380
rect 32100 12340 32588 12346
rect 32828 12296 32888 12444
rect 33118 12380 33606 12386
rect 33118 12346 33130 12380
rect 33594 12346 33606 12380
rect 33118 12340 33606 12346
rect 29770 12236 29782 12296
rect 28798 11776 28804 12232
rect 28798 11774 28810 11776
rect 28798 11720 28812 11774
rect 29776 11756 29782 12236
rect 29768 11720 29782 11756
rect 29816 12236 29830 12296
rect 30786 12256 30800 12296
rect 29816 11756 29822 12236
rect 30794 11776 30800 12256
rect 29816 11720 29828 11756
rect 25992 11670 26480 11676
rect 25992 11636 26004 11670
rect 26468 11636 26480 11670
rect 25992 11630 26480 11636
rect 25686 11522 25692 11582
rect 25752 11522 25758 11582
rect 25182 11412 25188 11472
rect 25248 11412 25254 11472
rect 24672 11306 24678 11366
rect 24738 11306 24744 11366
rect 24674 11200 24680 11260
rect 24740 11200 24746 11260
rect 23956 11148 24444 11154
rect 23956 11114 23968 11148
rect 24432 11114 24444 11148
rect 23956 11108 24444 11114
rect 24680 11064 24740 11200
rect 25188 11154 25248 11412
rect 24974 11148 25462 11154
rect 24974 11114 24986 11148
rect 25450 11114 25462 11148
rect 24974 11108 25462 11114
rect 25692 11064 25752 11522
rect 26196 11472 26256 11630
rect 26716 11504 26776 11720
rect 27208 11676 27268 11678
rect 27010 11670 27498 11676
rect 27010 11636 27022 11670
rect 27486 11636 27498 11670
rect 27010 11630 27498 11636
rect 26190 11412 26196 11472
rect 26256 11412 26262 11472
rect 26560 11444 26776 11504
rect 27208 11472 27268 11630
rect 27730 11582 27790 11720
rect 28758 11708 28804 11720
rect 28240 11676 28300 11678
rect 28028 11670 28516 11676
rect 28028 11636 28040 11670
rect 28504 11636 28516 11670
rect 28028 11630 28516 11636
rect 29046 11670 29534 11676
rect 29046 11636 29058 11670
rect 29522 11636 29534 11670
rect 29046 11630 29534 11636
rect 27724 11522 27730 11582
rect 27790 11522 27796 11582
rect 26196 11154 26256 11412
rect 26560 11260 26620 11444
rect 27202 11412 27208 11472
rect 27268 11412 27274 11472
rect 26708 11306 26714 11366
rect 26774 11306 26780 11366
rect 26554 11200 26560 11260
rect 26620 11200 26626 11260
rect 25992 11148 26480 11154
rect 25992 11114 26004 11148
rect 26468 11114 26480 11148
rect 25992 11108 26480 11114
rect 20654 11002 20664 11024
rect 21620 11008 21638 11064
rect 20654 10488 20660 11002
rect 21632 10530 21638 11008
rect 18578 10476 18624 10488
rect 19596 10476 19642 10488
rect 20614 10476 20660 10488
rect 21624 10488 21638 10530
rect 21672 11008 21680 11064
rect 22640 11012 22656 11064
rect 21672 10530 21678 11008
rect 21672 10488 21684 10530
rect 17848 10438 18336 10444
rect 17848 10404 17860 10438
rect 18324 10404 18336 10438
rect 17848 10398 18336 10404
rect 18866 10438 19354 10444
rect 18866 10404 18878 10438
rect 19342 10404 19354 10438
rect 18866 10398 19354 10404
rect 19884 10438 20372 10444
rect 19884 10404 19896 10438
rect 20360 10404 20372 10438
rect 19884 10398 20372 10404
rect 20902 10438 21390 10444
rect 20902 10404 20914 10438
rect 21378 10404 21390 10438
rect 20902 10398 21390 10404
rect 17540 10206 17546 10266
rect 17606 10206 17612 10266
rect 17546 9972 17552 10032
rect 17612 9972 17618 10032
rect 16828 9914 17316 9920
rect 16828 9880 16840 9914
rect 17304 9880 17316 9914
rect 16828 9874 17316 9880
rect 15562 9254 15568 9804
rect 16534 9798 16546 9830
rect 16540 9294 16546 9798
rect 15522 9242 15568 9254
rect 16532 9254 16546 9294
rect 16580 9798 16594 9830
rect 17552 9830 17612 9972
rect 18046 9920 18106 10398
rect 18560 10206 18566 10266
rect 18626 10206 18632 10266
rect 17846 9914 18334 9920
rect 17846 9880 17858 9914
rect 18322 9880 18334 9914
rect 17846 9874 18334 9880
rect 17552 9800 17564 9830
rect 16580 9294 16586 9798
rect 16580 9254 16592 9294
rect 14792 9204 15280 9210
rect 14792 9170 14804 9204
rect 15268 9170 15280 9204
rect 14792 9164 15280 9170
rect 15810 9204 16298 9210
rect 15810 9170 15822 9204
rect 16286 9170 16298 9204
rect 15810 9164 16298 9170
rect 13354 9042 13360 9102
rect 13420 9042 13426 9102
rect 14492 9042 14498 9102
rect 14558 9042 14564 9102
rect 13242 8842 13248 8902
rect 13308 8842 13314 8902
rect 13136 8740 13142 8800
rect 13202 8740 13208 8800
rect 13026 5288 13032 5348
rect 13092 5288 13098 5348
rect 13142 5310 13202 8740
rect 13248 7666 13308 8842
rect 13242 7606 13248 7666
rect 13308 7606 13314 7666
rect 12794 5138 12800 5198
rect 12860 5138 12866 5198
rect 13032 1612 13092 5288
rect 13136 5250 13142 5310
rect 13202 5250 13208 5310
rect 13142 2820 13202 5250
rect 13248 2946 13308 7606
rect 13360 6328 13420 9042
rect 14490 8842 14496 8902
rect 14556 8842 14562 8902
rect 14496 8798 14556 8842
rect 13480 8738 14556 8798
rect 13480 8736 14044 8738
rect 13480 8596 13540 8736
rect 13984 8686 14044 8736
rect 13774 8680 14262 8686
rect 13774 8646 13786 8680
rect 14250 8646 14262 8680
rect 13774 8640 14262 8646
rect 13480 8564 13492 8596
rect 13486 8020 13492 8564
rect 13526 8564 13540 8596
rect 14496 8596 14556 8738
rect 15000 8686 15060 9164
rect 15508 8962 15514 9022
rect 15574 8962 15580 9022
rect 14792 8680 15280 8686
rect 14792 8646 14804 8680
rect 15268 8646 15280 8680
rect 14792 8640 15280 8646
rect 13526 8020 13532 8564
rect 14496 8560 14510 8596
rect 13486 8008 13532 8020
rect 14504 8020 14510 8560
rect 14544 8560 14556 8596
rect 15514 8596 15574 8962
rect 16028 8908 16088 9164
rect 16532 9126 16592 9254
rect 17558 9254 17564 9800
rect 17598 9800 17612 9830
rect 18566 9830 18626 10206
rect 19072 9920 19132 10398
rect 19582 10310 19588 10370
rect 19648 10310 19654 10370
rect 18864 9914 19352 9920
rect 18864 9880 18876 9914
rect 19340 9880 19352 9914
rect 18864 9874 19352 9880
rect 17598 9254 17604 9800
rect 18566 9786 18582 9830
rect 18576 9304 18582 9786
rect 17558 9242 17604 9254
rect 18568 9254 18582 9304
rect 18616 9786 18626 9830
rect 19588 9830 19648 10310
rect 21624 10266 21684 10488
rect 22650 10488 22656 11012
rect 22690 11020 22704 11064
rect 22690 11012 22700 11020
rect 23656 11016 23674 11064
rect 22690 10488 22696 11012
rect 23668 10536 23674 11016
rect 22650 10476 22696 10488
rect 23662 10488 23674 10536
rect 23708 11016 23716 11064
rect 24676 11024 24692 11064
rect 23708 10536 23714 11016
rect 23708 10488 23722 10536
rect 21920 10438 22408 10444
rect 21920 10404 21932 10438
rect 22396 10404 22408 10438
rect 21920 10398 22408 10404
rect 22938 10438 23426 10444
rect 22938 10404 22950 10438
rect 23414 10404 23426 10438
rect 22938 10398 23426 10404
rect 23662 10266 23722 10488
rect 24686 10488 24692 11024
rect 24726 11026 24742 11064
rect 24726 11024 24740 11026
rect 24726 10488 24732 11024
rect 25692 11018 25710 11064
rect 25704 10542 25710 11018
rect 25692 10488 25710 10542
rect 25744 11018 25752 11064
rect 26714 11064 26774 11306
rect 27208 11154 27268 11412
rect 27010 11148 27498 11154
rect 27010 11114 27022 11148
rect 27486 11114 27498 11148
rect 27010 11108 27498 11114
rect 27730 11064 27790 11522
rect 28240 11472 28300 11630
rect 29254 11472 29314 11630
rect 29768 11582 29828 11720
rect 30784 11720 30800 11776
rect 30834 12256 30846 12296
rect 30834 11776 30840 12256
rect 30834 11720 30844 11776
rect 30064 11670 30552 11676
rect 30064 11636 30076 11670
rect 30540 11636 30552 11670
rect 30064 11630 30552 11636
rect 29762 11522 29768 11582
rect 29828 11522 29834 11582
rect 28234 11412 28240 11472
rect 28300 11412 28306 11472
rect 29248 11412 29254 11472
rect 29314 11412 29320 11472
rect 28240 11154 28300 11412
rect 28748 11306 28754 11366
rect 28814 11306 28820 11366
rect 28028 11148 28516 11154
rect 28028 11114 28040 11148
rect 28504 11114 28516 11148
rect 28028 11108 28516 11114
rect 28754 11064 28814 11306
rect 29254 11154 29314 11412
rect 29046 11148 29534 11154
rect 29046 11114 29058 11148
rect 29522 11114 29534 11148
rect 29046 11108 29534 11114
rect 25744 10542 25750 11018
rect 26714 11012 26728 11064
rect 25744 10488 25752 10542
rect 26722 10488 26728 11012
rect 26762 11022 26778 11064
rect 26762 11012 26774 11022
rect 26762 10488 26768 11012
rect 24686 10476 24732 10488
rect 25704 10476 25750 10488
rect 26722 10476 26768 10488
rect 27730 10488 27746 11064
rect 27780 10488 27790 11064
rect 28750 11022 28764 11064
rect 28754 11002 28764 11022
rect 23956 10438 24444 10444
rect 23956 10404 23968 10438
rect 24432 10404 24444 10438
rect 23956 10398 24444 10404
rect 24974 10438 25462 10444
rect 24974 10404 24986 10438
rect 25450 10404 25462 10438
rect 24974 10398 25462 10404
rect 25992 10438 26480 10444
rect 25992 10404 26004 10438
rect 26468 10404 26480 10438
rect 25992 10398 26480 10404
rect 27010 10438 27498 10444
rect 27010 10404 27022 10438
rect 27486 10404 27498 10438
rect 27010 10398 27498 10404
rect 25688 10310 25694 10370
rect 25754 10310 25760 10370
rect 21618 10206 21624 10266
rect 21684 10206 21690 10266
rect 23656 10206 23662 10266
rect 23722 10206 23728 10266
rect 20602 10084 20608 10144
rect 20668 10084 20674 10144
rect 22636 10084 22642 10144
rect 22702 10084 22708 10144
rect 24666 10084 24672 10144
rect 24732 10084 24738 10144
rect 19882 9914 20370 9920
rect 19882 9880 19894 9914
rect 20358 9880 20370 9914
rect 19882 9874 20370 9880
rect 18616 9304 18622 9786
rect 19588 9768 19600 9830
rect 18616 9254 18628 9304
rect 19594 9290 19600 9768
rect 16828 9204 17316 9210
rect 16828 9170 16840 9204
rect 17304 9170 17316 9204
rect 16828 9164 17316 9170
rect 17846 9204 18334 9210
rect 17846 9170 17858 9204
rect 18322 9170 18334 9204
rect 17846 9164 18334 9170
rect 16526 9066 16532 9126
rect 16592 9066 16598 9126
rect 16022 8848 16028 8908
rect 16088 8848 16094 8908
rect 16028 8686 16088 8848
rect 15810 8680 16298 8686
rect 15810 8646 15822 8680
rect 16286 8646 16298 8680
rect 15810 8640 16298 8646
rect 14544 8020 14550 8560
rect 15514 8554 15528 8596
rect 15522 8078 15528 8554
rect 14504 8008 14550 8020
rect 15516 8020 15528 8078
rect 15562 8554 15574 8596
rect 16532 8596 16592 9066
rect 17030 8914 17090 9164
rect 17548 8962 17554 9022
rect 17614 8962 17620 9022
rect 17030 8908 17092 8914
rect 17030 8848 17032 8908
rect 17030 8842 17092 8848
rect 17030 8686 17090 8842
rect 16828 8680 17316 8686
rect 16828 8646 16840 8680
rect 17304 8646 17316 8680
rect 16828 8640 17316 8646
rect 15562 8078 15568 8554
rect 16532 8552 16546 8596
rect 15562 8020 15576 8078
rect 16540 8068 16546 8552
rect 13774 7970 14262 7976
rect 13774 7936 13786 7970
rect 14250 7936 14262 7970
rect 13774 7930 14262 7936
rect 14792 7970 15280 7976
rect 14792 7936 14804 7970
rect 15268 7936 15280 7970
rect 14792 7930 15280 7936
rect 14490 7810 14496 7870
rect 14556 7810 14562 7870
rect 13774 7448 14262 7454
rect 13774 7414 13786 7448
rect 14250 7414 14262 7448
rect 13774 7408 14262 7414
rect 13486 7364 13532 7376
rect 13486 6834 13492 7364
rect 13476 6788 13492 6834
rect 13526 6834 13532 7364
rect 14496 7364 14556 7810
rect 15002 7768 15062 7930
rect 14996 7708 15002 7768
rect 15062 7708 15068 7768
rect 15516 7566 15576 8020
rect 16534 8020 16546 8068
rect 16580 8552 16592 8596
rect 17554 8596 17614 8962
rect 18046 8914 18106 9164
rect 18568 9126 18628 9254
rect 19586 9254 19600 9290
rect 19634 9768 19648 9830
rect 20608 9830 20668 10084
rect 20900 9914 21388 9920
rect 20900 9880 20912 9914
rect 21376 9880 21388 9914
rect 20900 9874 21388 9880
rect 21918 9914 22406 9920
rect 21918 9880 21930 9914
rect 22394 9880 22406 9914
rect 21918 9874 22406 9880
rect 20608 9774 20618 9830
rect 19634 9290 19640 9768
rect 19634 9254 19646 9290
rect 18864 9204 19352 9210
rect 18864 9170 18876 9204
rect 19340 9170 19352 9204
rect 18864 9164 19352 9170
rect 18562 9066 18568 9126
rect 18628 9066 18634 9126
rect 18044 8908 18106 8914
rect 18104 8848 18106 8908
rect 18044 8842 18106 8848
rect 18046 8686 18106 8842
rect 17846 8680 18334 8686
rect 17846 8646 17858 8680
rect 18322 8646 18334 8680
rect 17846 8640 18334 8646
rect 17554 8554 17564 8596
rect 16580 8068 16586 8552
rect 16580 8020 16594 8068
rect 15810 7970 16298 7976
rect 15810 7936 15822 7970
rect 16286 7936 16298 7970
rect 15810 7930 16298 7936
rect 16534 7870 16594 8020
rect 17558 8020 17564 8554
rect 17598 8554 17614 8596
rect 18568 8596 18628 9066
rect 19064 8908 19124 9164
rect 19586 9022 19646 9254
rect 20612 9254 20618 9774
rect 20652 9774 20668 9830
rect 21630 9830 21676 9842
rect 20652 9254 20658 9774
rect 21630 9284 21636 9830
rect 20612 9242 20658 9254
rect 21620 9254 21636 9284
rect 21670 9284 21676 9830
rect 22642 9830 22702 10084
rect 22936 9914 23424 9920
rect 22936 9880 22948 9914
rect 23412 9880 23424 9914
rect 22936 9874 23424 9880
rect 23954 9914 24442 9920
rect 23954 9880 23966 9914
rect 24430 9880 24442 9914
rect 23954 9874 24442 9880
rect 22642 9780 22654 9830
rect 21670 9254 21680 9284
rect 19882 9204 20370 9210
rect 19882 9170 19894 9204
rect 20358 9170 20370 9204
rect 19882 9164 20370 9170
rect 20900 9204 21388 9210
rect 20900 9170 20912 9204
rect 21376 9170 21388 9204
rect 20900 9164 21388 9170
rect 19580 8962 19586 9022
rect 19646 8962 19652 9022
rect 20076 8966 20136 9164
rect 21118 8966 21178 9164
rect 21620 9022 21680 9254
rect 22648 9254 22654 9780
rect 22688 9780 22702 9830
rect 23666 9830 23712 9842
rect 22688 9254 22694 9780
rect 23666 9296 23672 9830
rect 22648 9242 22694 9254
rect 23660 9254 23672 9296
rect 23706 9296 23712 9830
rect 24672 9830 24732 10084
rect 24972 9914 25460 9920
rect 24972 9880 24984 9914
rect 25448 9880 25460 9914
rect 24972 9874 25460 9880
rect 24672 9786 24690 9830
rect 23706 9254 23720 9296
rect 21918 9204 22406 9210
rect 21918 9170 21930 9204
rect 22394 9170 22406 9204
rect 21918 9164 22406 9170
rect 22936 9204 23424 9210
rect 22936 9170 22948 9204
rect 23412 9170 23424 9204
rect 22936 9164 23424 9170
rect 19580 8850 19586 8910
rect 19646 8850 19652 8910
rect 20076 8906 21178 8966
rect 21614 8962 21620 9022
rect 21680 8962 21686 9022
rect 19064 8686 19124 8848
rect 18864 8680 19352 8686
rect 18864 8646 18876 8680
rect 19340 8646 19352 8680
rect 18864 8640 19352 8646
rect 17598 8020 17604 8554
rect 18568 8548 18582 8596
rect 18576 8070 18582 8548
rect 17558 8008 17604 8020
rect 18570 8020 18582 8070
rect 18616 8548 18628 8596
rect 19586 8596 19646 8850
rect 20076 8686 20136 8906
rect 20598 8740 20604 8800
rect 20664 8740 20670 8800
rect 19882 8680 20370 8686
rect 19882 8646 19894 8680
rect 20358 8646 20370 8680
rect 19882 8640 20370 8646
rect 18616 8070 18622 8548
rect 19586 8538 19600 8596
rect 18616 8020 18630 8070
rect 16828 7970 17316 7976
rect 16828 7936 16840 7970
rect 17304 7936 17316 7970
rect 16828 7930 17316 7936
rect 17846 7970 18334 7976
rect 17846 7936 17858 7970
rect 18322 7936 18334 7970
rect 17846 7930 18334 7936
rect 16528 7810 16534 7870
rect 16594 7810 16600 7870
rect 16526 7606 16532 7666
rect 16592 7606 16598 7666
rect 17040 7660 17100 7930
rect 18062 7660 18122 7930
rect 18570 7870 18630 8020
rect 19594 8020 19600 8538
rect 19634 8538 19646 8596
rect 20604 8596 20664 8740
rect 21118 8686 21178 8906
rect 21616 8850 21622 8910
rect 21682 8850 21688 8910
rect 20900 8680 21388 8686
rect 20900 8646 20912 8680
rect 21376 8646 21388 8680
rect 20900 8640 21388 8646
rect 20604 8550 20618 8596
rect 19634 8020 19640 8538
rect 19594 8008 19640 8020
rect 20612 8020 20618 8550
rect 20652 8550 20664 8596
rect 21622 8596 21682 8850
rect 22118 8686 22178 9164
rect 22632 8740 22638 8800
rect 22698 8740 22704 8800
rect 21918 8680 22406 8686
rect 21918 8646 21930 8680
rect 22394 8646 22406 8680
rect 21918 8640 22406 8646
rect 20652 8020 20658 8550
rect 21622 8528 21636 8596
rect 20612 8008 20658 8020
rect 21630 8020 21636 8528
rect 21670 8528 21682 8596
rect 22638 8596 22698 8740
rect 23152 8686 23212 9164
rect 23660 9022 23720 9254
rect 24684 9254 24690 9786
rect 24724 9786 24732 9830
rect 25694 9830 25754 10310
rect 26216 9920 26276 10398
rect 26706 10206 26712 10266
rect 26772 10206 26778 10266
rect 25990 9914 26478 9920
rect 25990 9880 26002 9914
rect 26466 9880 26478 9914
rect 25990 9874 26478 9880
rect 24724 9254 24730 9786
rect 25694 9778 25708 9830
rect 25702 9306 25708 9778
rect 24684 9242 24730 9254
rect 25694 9254 25708 9306
rect 25742 9778 25754 9830
rect 26712 9830 26772 10206
rect 27218 9920 27278 10398
rect 27730 10266 27790 10488
rect 28758 10488 28764 11002
rect 28798 11002 28814 11064
rect 29768 11064 29828 11522
rect 30272 11472 30332 11630
rect 30266 11412 30272 11472
rect 30332 11412 30338 11472
rect 30272 11154 30332 11412
rect 30784 11366 30844 11720
rect 31804 11720 31818 12296
rect 31852 12264 31866 12296
rect 32824 12268 32836 12296
rect 31852 11720 31864 12264
rect 32828 12232 32836 12268
rect 32830 11780 32836 12232
rect 31082 11670 31570 11676
rect 31082 11636 31094 11670
rect 31558 11636 31570 11670
rect 31082 11630 31570 11636
rect 31296 11472 31356 11630
rect 31804 11582 31864 11720
rect 32824 11720 32836 11780
rect 32870 12232 32888 12296
rect 33848 12296 33894 12308
rect 32870 11780 32876 12232
rect 32870 11720 32884 11780
rect 33848 11768 33854 12296
rect 32100 11670 32588 11676
rect 32100 11636 32112 11670
rect 32576 11636 32588 11670
rect 32100 11630 32588 11636
rect 31798 11522 31804 11582
rect 31864 11522 31870 11582
rect 31290 11412 31296 11472
rect 31356 11412 31362 11472
rect 30778 11306 30784 11366
rect 30844 11306 30850 11366
rect 30778 11202 30784 11262
rect 30844 11202 30850 11262
rect 30064 11148 30552 11154
rect 30064 11114 30076 11148
rect 30540 11114 30552 11148
rect 30064 11108 30552 11114
rect 30264 11096 30324 11108
rect 30784 11064 30844 11202
rect 31296 11154 31356 11412
rect 31082 11148 31570 11154
rect 31082 11114 31094 11148
rect 31558 11114 31570 11148
rect 31082 11108 31570 11114
rect 29768 11006 29782 11064
rect 28798 10488 28804 11002
rect 29776 10536 29782 11006
rect 28758 10476 28804 10488
rect 29766 10488 29782 10536
rect 29816 11006 29828 11064
rect 30782 11018 30800 11064
rect 29816 10536 29822 11006
rect 30784 10990 30800 11018
rect 30794 10542 30800 10990
rect 29816 10488 29826 10536
rect 28028 10438 28516 10444
rect 28028 10404 28040 10438
rect 28504 10404 28516 10438
rect 28028 10398 28516 10404
rect 29046 10438 29534 10444
rect 29046 10404 29058 10438
rect 29522 10404 29534 10438
rect 29046 10398 29534 10404
rect 27724 10206 27730 10266
rect 27790 10206 27796 10266
rect 28230 9920 28290 10398
rect 28744 10206 28750 10266
rect 28810 10206 28816 10266
rect 27008 9914 27496 9920
rect 27008 9880 27020 9914
rect 27484 9880 27496 9914
rect 27008 9874 27496 9880
rect 28026 9914 28514 9920
rect 28026 9880 28038 9914
rect 28502 9880 28514 9914
rect 28026 9874 28514 9880
rect 26712 9782 26726 9830
rect 25742 9306 25748 9778
rect 25742 9254 25754 9306
rect 26720 9286 26726 9782
rect 23954 9204 24442 9210
rect 23954 9170 23966 9204
rect 24430 9170 24442 9204
rect 23954 9164 24442 9170
rect 24972 9204 25460 9210
rect 24972 9170 24984 9204
rect 25448 9170 25460 9204
rect 24972 9164 25460 9170
rect 23654 8962 23660 9022
rect 23720 8962 23726 9022
rect 24174 8966 24234 9164
rect 25182 8966 25242 9164
rect 25694 9022 25754 9254
rect 26712 9254 26726 9286
rect 26760 9782 26772 9830
rect 27738 9830 27784 9842
rect 26760 9286 26766 9782
rect 27738 9290 27744 9830
rect 26760 9254 26772 9286
rect 25990 9204 26478 9210
rect 25990 9170 26002 9204
rect 26466 9170 26478 9204
rect 25990 9164 26478 9170
rect 23652 8850 23658 8910
rect 23718 8850 23724 8910
rect 24174 8906 25242 8966
rect 25688 8962 25694 9022
rect 25754 8962 25760 9022
rect 25884 8958 25890 9018
rect 25950 8958 25956 9018
rect 22936 8680 23424 8686
rect 22936 8646 22948 8680
rect 23412 8646 23424 8680
rect 22936 8640 23424 8646
rect 22638 8548 22654 8596
rect 21670 8020 21676 8528
rect 21630 8008 21676 8020
rect 22648 8020 22654 8548
rect 22688 8548 22698 8596
rect 23658 8596 23718 8850
rect 24174 8686 24234 8906
rect 24672 8740 24678 8800
rect 24738 8740 24744 8800
rect 23954 8680 24442 8686
rect 23954 8646 23966 8680
rect 24430 8646 24442 8680
rect 23954 8640 24442 8646
rect 22688 8020 22694 8548
rect 23658 8546 23672 8596
rect 22648 8008 22694 8020
rect 23666 8020 23672 8546
rect 23706 8546 23718 8596
rect 24678 8596 24738 8740
rect 25182 8686 25242 8906
rect 25688 8850 25694 8910
rect 25754 8850 25760 8910
rect 24972 8680 25460 8686
rect 24972 8646 24984 8680
rect 25448 8646 25460 8680
rect 24972 8640 25460 8646
rect 24678 8558 24690 8596
rect 23706 8020 23712 8546
rect 24684 8066 24690 8558
rect 23666 8008 23712 8020
rect 24678 8020 24690 8066
rect 24724 8558 24738 8596
rect 25694 8596 25754 8850
rect 25890 8800 25950 8958
rect 26184 8802 26244 9164
rect 26712 9126 26772 9254
rect 27728 9254 27744 9290
rect 27778 9290 27784 9830
rect 28750 9830 28810 10206
rect 29264 9920 29324 10398
rect 29766 10266 29826 10488
rect 30788 10488 30800 10542
rect 30834 10990 30844 11064
rect 31804 11064 31864 11522
rect 32316 11472 32376 11630
rect 32824 11572 32884 11720
rect 33840 11720 33854 11768
rect 33888 11768 33894 12296
rect 33888 11720 33900 11768
rect 33118 11670 33606 11676
rect 33118 11636 33130 11670
rect 33594 11636 33606 11670
rect 33118 11630 33606 11636
rect 33334 11572 33394 11630
rect 33840 11572 33900 11720
rect 33960 11572 34020 12444
rect 32824 11512 34020 11572
rect 32310 11412 32316 11472
rect 32376 11412 32382 11472
rect 32316 11154 32376 11412
rect 32818 11306 32824 11366
rect 32884 11306 32890 11366
rect 32824 11264 32884 11306
rect 32824 11204 33902 11264
rect 33960 11262 34020 11512
rect 32100 11148 32588 11154
rect 32100 11114 32112 11148
rect 32576 11114 32588 11148
rect 32100 11108 32588 11114
rect 31804 11038 31818 11064
rect 30834 10542 30840 10990
rect 31812 10546 31818 11038
rect 30834 10488 30848 10542
rect 30064 10438 30552 10444
rect 30064 10404 30076 10438
rect 30540 10404 30552 10438
rect 30064 10398 30552 10404
rect 30788 10370 30848 10488
rect 31802 10488 31818 10546
rect 31852 11038 31864 11064
rect 32824 11064 32884 11204
rect 33310 11154 33370 11204
rect 33118 11148 33606 11154
rect 33118 11114 33130 11148
rect 33594 11114 33606 11148
rect 33118 11108 33606 11114
rect 33842 11064 33902 11204
rect 33954 11202 33960 11262
rect 34020 11202 34026 11262
rect 31852 10546 31858 11038
rect 32824 11008 32836 11064
rect 31852 10488 31862 10546
rect 31082 10438 31570 10444
rect 31082 10404 31094 10438
rect 31558 10404 31570 10438
rect 31082 10398 31570 10404
rect 30782 10310 30788 10370
rect 30848 10310 30854 10370
rect 31802 10266 31862 10488
rect 32830 10488 32836 11008
rect 32870 11008 32884 11064
rect 33838 11028 33854 11064
rect 33842 11022 33854 11028
rect 32870 10488 32876 11008
rect 33848 10532 33854 11022
rect 32830 10476 32876 10488
rect 33844 10488 33854 10532
rect 33888 11022 33902 11064
rect 33888 10532 33894 11022
rect 33888 10488 33904 10532
rect 32100 10438 32588 10444
rect 32100 10404 32112 10438
rect 32576 10404 32588 10438
rect 32100 10398 32588 10404
rect 33118 10438 33606 10444
rect 33118 10404 33130 10438
rect 33594 10404 33606 10438
rect 33118 10398 33606 10404
rect 29760 10206 29766 10266
rect 29826 10206 29832 10266
rect 31796 10206 31802 10266
rect 31862 10206 31868 10266
rect 32292 9920 32352 10398
rect 33844 10362 33904 10488
rect 33844 10302 34134 10362
rect 33330 9996 33898 10056
rect 33330 9920 33390 9996
rect 29044 9914 29532 9920
rect 29044 9880 29056 9914
rect 29520 9880 29532 9914
rect 29044 9874 29532 9880
rect 30062 9914 30550 9920
rect 30062 9880 30074 9914
rect 30538 9880 30550 9914
rect 30062 9874 30550 9880
rect 31080 9914 31568 9920
rect 31080 9880 31092 9914
rect 31556 9880 31568 9914
rect 31080 9874 31568 9880
rect 32098 9914 32586 9920
rect 32098 9880 32110 9914
rect 32574 9880 32586 9914
rect 32098 9874 32586 9880
rect 33116 9914 33604 9920
rect 33116 9880 33128 9914
rect 33592 9880 33604 9914
rect 33116 9874 33604 9880
rect 28750 9772 28762 9830
rect 28756 9300 28762 9772
rect 27778 9254 27788 9290
rect 27008 9204 27496 9210
rect 27008 9170 27020 9204
rect 27484 9170 27496 9204
rect 27008 9164 27496 9170
rect 26706 9066 26712 9126
rect 26772 9066 26778 9126
rect 25884 8740 25890 8800
rect 25950 8740 25956 8800
rect 26178 8742 26184 8802
rect 26244 8742 26250 8802
rect 26184 8686 26244 8742
rect 25990 8680 26478 8686
rect 25990 8646 26002 8680
rect 26466 8646 26478 8680
rect 25990 8640 26478 8646
rect 24724 8066 24730 8558
rect 25694 8552 25708 8596
rect 24724 8020 24738 8066
rect 18864 7970 19352 7976
rect 18864 7936 18876 7970
rect 19340 7936 19352 7970
rect 18864 7930 19352 7936
rect 19882 7970 20370 7976
rect 19882 7936 19894 7970
rect 20358 7936 20370 7970
rect 19882 7930 20370 7936
rect 20900 7970 21388 7976
rect 20900 7936 20912 7970
rect 21376 7936 21388 7970
rect 20900 7930 21388 7936
rect 21918 7970 22406 7976
rect 21918 7936 21930 7970
rect 22394 7936 22406 7970
rect 21918 7930 22406 7936
rect 22936 7970 23424 7976
rect 22936 7936 22948 7970
rect 23412 7936 23424 7970
rect 22936 7930 23424 7936
rect 23954 7970 24442 7976
rect 23954 7936 23966 7970
rect 24430 7936 24442 7970
rect 23954 7930 24442 7936
rect 18564 7810 18570 7870
rect 18630 7810 18636 7870
rect 15510 7506 15516 7566
rect 15576 7506 15582 7566
rect 14792 7448 15280 7454
rect 14792 7414 14804 7448
rect 15268 7414 15280 7448
rect 14792 7408 15280 7414
rect 14496 7326 14510 7364
rect 13526 6788 13536 6834
rect 14504 6830 14510 7326
rect 13476 6626 13536 6788
rect 14494 6788 14510 6830
rect 14544 7326 14556 7364
rect 15516 7364 15576 7506
rect 15810 7448 16298 7454
rect 15810 7414 15822 7448
rect 16286 7414 16298 7448
rect 15810 7408 16298 7414
rect 14544 6830 14550 7326
rect 15516 7324 15528 7364
rect 14544 6788 14554 6830
rect 13774 6738 14262 6744
rect 13774 6704 13786 6738
rect 14250 6704 14262 6738
rect 13774 6698 14262 6704
rect 13988 6626 14048 6698
rect 14494 6626 14554 6788
rect 15522 6788 15528 7324
rect 15562 7324 15576 7364
rect 16532 7364 16592 7606
rect 17034 7600 17040 7660
rect 17100 7600 17106 7660
rect 18056 7600 18062 7660
rect 18122 7600 18128 7660
rect 17544 7506 17550 7566
rect 17610 7506 17616 7566
rect 16828 7448 17316 7454
rect 16828 7414 16840 7448
rect 17304 7414 17316 7448
rect 16828 7408 17316 7414
rect 15562 6788 15568 7324
rect 16532 7312 16546 7364
rect 15522 6776 15568 6788
rect 16540 6788 16546 7312
rect 16580 7312 16592 7364
rect 17550 7364 17610 7506
rect 18062 7454 18122 7600
rect 17846 7448 18334 7454
rect 17846 7414 17858 7448
rect 18322 7414 18334 7448
rect 17846 7408 18334 7414
rect 17550 7320 17564 7364
rect 16580 6788 16586 7312
rect 17558 6824 17564 7320
rect 16540 6776 16586 6788
rect 17550 6788 17564 6824
rect 17598 7320 17610 7364
rect 18570 7364 18630 7810
rect 19076 7660 19136 7930
rect 20094 7768 20154 7930
rect 21114 7880 21174 7930
rect 22114 7880 22174 7930
rect 23152 7880 23212 7930
rect 24180 7880 24240 7930
rect 20596 7810 20602 7870
rect 20662 7810 20668 7870
rect 21114 7820 24240 7880
rect 20088 7708 20094 7768
rect 20154 7708 20160 7768
rect 19070 7600 19076 7660
rect 19136 7600 19142 7660
rect 20088 7600 20094 7660
rect 20154 7600 20160 7660
rect 19076 7454 19136 7600
rect 19580 7506 19586 7566
rect 19646 7506 19652 7566
rect 18864 7448 19352 7454
rect 18864 7414 18876 7448
rect 19340 7414 19352 7448
rect 18864 7408 19352 7414
rect 17598 6824 17604 7320
rect 17598 6788 17610 6824
rect 14792 6738 15280 6744
rect 14792 6704 14804 6738
rect 15268 6704 15280 6738
rect 14792 6698 15280 6704
rect 15810 6738 16298 6744
rect 15810 6704 15822 6738
rect 16286 6704 16298 6738
rect 15810 6698 16298 6704
rect 16828 6738 17316 6744
rect 16828 6704 16840 6738
rect 17304 6704 17316 6738
rect 16828 6698 17316 6704
rect 14998 6642 15058 6698
rect 13476 6566 14554 6626
rect 14992 6582 14998 6642
rect 15058 6582 15064 6642
rect 15902 6582 15908 6642
rect 15968 6582 15974 6642
rect 14992 6366 14998 6426
rect 15058 6366 15064 6426
rect 14998 6360 15060 6366
rect 13360 6322 13422 6328
rect 13360 6262 13362 6322
rect 13360 6256 13422 6262
rect 13360 4078 13420 6256
rect 15000 6220 15060 6360
rect 15908 6220 15968 6582
rect 16036 6426 16096 6698
rect 16904 6582 16910 6642
rect 16970 6582 16976 6642
rect 16036 6360 16096 6366
rect 16910 6220 16970 6582
rect 17050 6426 17110 6698
rect 17550 6540 17610 6788
rect 18570 6788 18582 7364
rect 18616 6788 18630 7364
rect 19586 7364 19646 7506
rect 20094 7454 20154 7600
rect 19882 7448 20370 7454
rect 19882 7414 19894 7448
rect 20358 7414 20370 7448
rect 19882 7408 20370 7414
rect 19586 7328 19600 7364
rect 17846 6738 18334 6744
rect 17846 6704 17858 6738
rect 18322 6704 18334 6738
rect 17846 6698 18334 6704
rect 18062 6642 18122 6698
rect 18056 6582 18062 6642
rect 18122 6582 18128 6642
rect 17544 6480 17550 6540
rect 17610 6480 17616 6540
rect 17044 6366 17050 6426
rect 17110 6366 17116 6426
rect 18062 6220 18122 6582
rect 13774 6214 14262 6220
rect 13774 6180 13786 6214
rect 14250 6180 14262 6214
rect 13774 6174 14262 6180
rect 14792 6214 15280 6220
rect 14792 6180 14804 6214
rect 15268 6180 15280 6214
rect 14792 6174 15280 6180
rect 15810 6214 16298 6220
rect 15810 6180 15822 6214
rect 16286 6180 16298 6214
rect 15810 6174 16298 6180
rect 16828 6214 17316 6220
rect 16828 6180 16840 6214
rect 17304 6180 17316 6214
rect 16828 6174 17316 6180
rect 17846 6214 18334 6220
rect 17846 6180 17858 6214
rect 18322 6180 18334 6214
rect 17846 6174 18334 6180
rect 13486 6130 13532 6142
rect 13486 5592 13492 6130
rect 13480 5554 13492 5592
rect 13526 5592 13532 6130
rect 14504 6130 14550 6142
rect 14504 5592 14510 6130
rect 13526 5554 13540 5592
rect 13480 5424 13540 5554
rect 14498 5554 14510 5592
rect 14544 5592 14550 6130
rect 15522 6130 15568 6142
rect 15522 5604 15528 6130
rect 14544 5554 14558 5592
rect 13774 5504 14262 5510
rect 13774 5470 13786 5504
rect 14250 5470 14262 5504
rect 13774 5464 14262 5470
rect 13978 5424 14038 5464
rect 14498 5424 14558 5554
rect 15514 5554 15528 5604
rect 15562 5604 15568 6130
rect 16540 6130 16586 6142
rect 16540 5612 16546 6130
rect 15562 5554 15574 5604
rect 14792 5504 15280 5510
rect 14792 5470 14804 5504
rect 15268 5470 15280 5504
rect 14792 5464 15280 5470
rect 13480 5364 14558 5424
rect 14498 5310 14558 5364
rect 14990 5354 14996 5414
rect 15056 5354 15062 5414
rect 14492 5250 14498 5310
rect 14558 5250 14564 5310
rect 14488 5040 14494 5100
rect 14554 5040 14560 5100
rect 13774 4980 14262 4986
rect 13774 4946 13786 4980
rect 14250 4946 14262 4980
rect 13774 4940 14262 4946
rect 13486 4896 13532 4908
rect 13486 4354 13492 4896
rect 13476 4320 13492 4354
rect 13526 4354 13532 4896
rect 14494 4896 14554 5040
rect 14996 4986 15056 5354
rect 15514 5198 15574 5554
rect 16532 5554 16546 5612
rect 16580 5612 16586 6130
rect 17558 6130 17604 6142
rect 16580 5554 16592 5612
rect 17558 5600 17564 6130
rect 15810 5504 16298 5510
rect 15810 5470 15822 5504
rect 16286 5470 16298 5504
rect 15810 5464 16298 5470
rect 16004 5414 16064 5464
rect 15998 5354 16004 5414
rect 16064 5354 16070 5414
rect 15508 5138 15514 5198
rect 15574 5138 15580 5198
rect 16532 5100 16592 5554
rect 17552 5554 17564 5600
rect 17598 5600 17604 6130
rect 18570 6130 18630 6788
rect 19594 6788 19600 7328
rect 19634 7328 19646 7364
rect 20602 7364 20662 7810
rect 21108 7600 21114 7660
rect 21174 7600 21180 7660
rect 24180 7644 24240 7820
rect 24678 7754 24738 8020
rect 25702 8020 25708 8552
rect 25742 8552 25754 8596
rect 26712 8596 26772 9066
rect 27214 8808 27274 9164
rect 27728 8910 27788 9254
rect 28748 9254 28762 9300
rect 28796 9772 28810 9830
rect 29774 9830 29820 9842
rect 28796 9300 28802 9772
rect 29774 9310 29780 9830
rect 28796 9254 28808 9300
rect 28026 9204 28514 9210
rect 28026 9170 28038 9204
rect 28502 9170 28514 9204
rect 28026 9164 28514 9170
rect 27722 8850 27728 8910
rect 27788 8850 27794 8910
rect 27212 8802 27274 8808
rect 27272 8742 27274 8802
rect 27212 8736 27274 8742
rect 27724 8736 27730 8796
rect 27790 8736 27796 8796
rect 27214 8686 27274 8736
rect 27008 8680 27496 8686
rect 27008 8646 27020 8680
rect 27484 8646 27496 8680
rect 27008 8640 27496 8646
rect 26712 8552 26726 8596
rect 25742 8020 25748 8552
rect 25702 8008 25748 8020
rect 26720 8020 26726 8552
rect 26760 8552 26772 8596
rect 27730 8596 27790 8736
rect 28238 8686 28298 9164
rect 28748 9126 28808 9254
rect 29766 9254 29780 9310
rect 29814 9310 29820 9830
rect 30792 9830 30838 9842
rect 29814 9254 29826 9310
rect 30792 9298 30798 9830
rect 29044 9204 29532 9210
rect 29044 9170 29056 9204
rect 29520 9170 29532 9204
rect 29044 9164 29532 9170
rect 28742 9066 28748 9126
rect 28808 9066 28814 9126
rect 28026 8680 28514 8686
rect 28026 8646 28038 8680
rect 28502 8646 28514 8680
rect 28026 8640 28514 8646
rect 27730 8566 27744 8596
rect 26760 8020 26766 8552
rect 27738 8060 27744 8566
rect 26720 8008 26766 8020
rect 27730 8020 27744 8060
rect 27778 8566 27790 8596
rect 28748 8596 28808 9066
rect 29264 8686 29324 9164
rect 29766 8910 29826 9254
rect 30782 9254 30798 9298
rect 30832 9298 30838 9830
rect 31810 9830 31856 9842
rect 31810 9298 31816 9830
rect 30832 9254 30842 9298
rect 30062 9204 30550 9210
rect 30062 9170 30074 9204
rect 30538 9170 30550 9204
rect 30062 9164 30550 9170
rect 29760 8850 29766 8910
rect 29826 8850 29832 8910
rect 30272 8860 30332 9164
rect 30782 9018 30842 9254
rect 31806 9254 31816 9298
rect 31850 9298 31856 9830
rect 32828 9830 32874 9842
rect 32828 9304 32834 9830
rect 31850 9254 31866 9298
rect 31080 9204 31568 9210
rect 31080 9170 31092 9204
rect 31556 9170 31568 9204
rect 31080 9164 31568 9170
rect 31288 9020 31348 9164
rect 30776 8958 30782 9018
rect 30842 8958 30848 9018
rect 31286 9014 31348 9020
rect 31346 8954 31348 9014
rect 31286 8948 31348 8954
rect 31288 8860 31348 8948
rect 31806 8910 31866 9254
rect 32822 9254 32834 9304
rect 32868 9304 32874 9830
rect 33838 9830 33898 9996
rect 33940 9972 33946 10032
rect 34006 9972 34012 10032
rect 34074 10014 34134 10302
rect 33838 9802 33852 9830
rect 33846 9312 33852 9802
rect 32868 9254 32882 9304
rect 32098 9204 32586 9210
rect 32098 9170 32110 9204
rect 32574 9170 32586 9204
rect 32098 9164 32586 9170
rect 30272 8800 31348 8860
rect 31800 8850 31806 8910
rect 31866 8850 31872 8910
rect 29760 8736 29766 8796
rect 29826 8736 29832 8796
rect 29044 8680 29532 8686
rect 29044 8646 29056 8680
rect 29520 8646 29532 8680
rect 29044 8640 29532 8646
rect 27778 8060 27784 8566
rect 28748 8556 28762 8596
rect 27778 8020 27790 8060
rect 28756 8054 28762 8556
rect 24972 7970 25460 7976
rect 24972 7936 24984 7970
rect 25448 7936 25460 7970
rect 24972 7930 25460 7936
rect 25990 7970 26478 7976
rect 25990 7936 26002 7970
rect 26466 7936 26478 7970
rect 25990 7930 26478 7936
rect 27008 7970 27496 7976
rect 27008 7936 27020 7970
rect 27484 7936 27496 7970
rect 27008 7930 27496 7936
rect 25184 7882 25244 7930
rect 24672 7694 24678 7754
rect 24738 7694 24744 7754
rect 25184 7644 25244 7822
rect 21114 7454 21174 7600
rect 24180 7584 25244 7644
rect 26708 7496 26714 7556
rect 26774 7496 26780 7556
rect 20900 7448 21388 7454
rect 20900 7414 20912 7448
rect 21376 7414 21388 7448
rect 20900 7408 21388 7414
rect 21918 7448 22406 7454
rect 21918 7414 21930 7448
rect 22394 7414 22406 7448
rect 21918 7408 22406 7414
rect 22936 7448 23424 7454
rect 22936 7414 22948 7448
rect 23412 7414 23424 7448
rect 22936 7408 23424 7414
rect 23954 7448 24442 7454
rect 23954 7414 23966 7448
rect 24430 7414 24442 7448
rect 23954 7408 24442 7414
rect 24972 7448 25460 7454
rect 24972 7414 24984 7448
rect 25448 7414 25460 7448
rect 24972 7408 25460 7414
rect 25990 7448 26478 7454
rect 25990 7414 26002 7448
rect 26466 7414 26478 7448
rect 25990 7408 26478 7414
rect 19634 6788 19640 7328
rect 20602 7326 20618 7364
rect 19594 6776 19640 6788
rect 20612 6788 20618 7326
rect 20652 7326 20662 7364
rect 21630 7364 21676 7376
rect 20652 6788 20658 7326
rect 21630 6830 21636 7364
rect 20612 6776 20658 6788
rect 21622 6788 21636 6830
rect 21670 6830 21676 7364
rect 22648 7364 22694 7376
rect 21670 6788 21682 6830
rect 22648 6826 22654 7364
rect 18864 6738 19352 6744
rect 18864 6704 18876 6738
rect 19340 6704 19352 6738
rect 18864 6698 19352 6704
rect 19882 6738 20370 6744
rect 19882 6704 19894 6738
rect 20358 6704 20370 6738
rect 19882 6698 20370 6704
rect 20900 6738 21388 6744
rect 20900 6704 20912 6738
rect 21376 6704 21388 6738
rect 20900 6698 21388 6704
rect 19072 6642 19132 6698
rect 20078 6642 20138 6698
rect 21122 6642 21182 6698
rect 21622 6648 21682 6788
rect 22642 6788 22654 6826
rect 22688 6826 22694 7364
rect 23666 7364 23712 7376
rect 22688 6788 22702 6826
rect 23666 6820 23672 7364
rect 21918 6738 22406 6744
rect 21918 6704 21930 6738
rect 22394 6704 22406 6738
rect 21918 6698 22406 6704
rect 19066 6582 19072 6642
rect 19132 6582 19138 6642
rect 20072 6582 20078 6642
rect 20138 6582 20144 6642
rect 21116 6582 21122 6642
rect 21182 6582 21188 6642
rect 21616 6588 21622 6648
rect 21682 6588 21688 6648
rect 19072 6220 19132 6582
rect 20070 6366 20076 6426
rect 20136 6366 20142 6426
rect 21110 6366 21116 6426
rect 21176 6366 21182 6426
rect 20076 6220 20136 6366
rect 20594 6262 20600 6322
rect 20660 6262 20666 6322
rect 18864 6214 19352 6220
rect 18864 6180 18876 6214
rect 19340 6180 19352 6214
rect 18864 6174 19352 6180
rect 19882 6214 20370 6220
rect 19882 6180 19894 6214
rect 20358 6180 20370 6214
rect 19882 6174 20370 6180
rect 18570 6048 18582 6130
rect 18576 5600 18582 6048
rect 17598 5554 17612 5600
rect 16828 5504 17316 5510
rect 16828 5470 16840 5504
rect 17304 5470 17316 5504
rect 16828 5464 17316 5470
rect 17018 5414 17078 5464
rect 17012 5354 17018 5414
rect 17078 5354 17084 5414
rect 17552 5198 17612 5554
rect 18572 5554 18582 5600
rect 18616 6048 18630 6130
rect 19594 6130 19640 6142
rect 18616 5600 18622 6048
rect 18616 5554 18632 5600
rect 19594 5598 19600 6130
rect 17846 5504 18334 5510
rect 17846 5470 17858 5504
rect 18322 5470 18334 5504
rect 17846 5464 18334 5470
rect 18056 5414 18116 5464
rect 18050 5354 18056 5414
rect 18116 5354 18122 5414
rect 17546 5138 17552 5198
rect 17612 5138 17618 5198
rect 16526 5040 16532 5100
rect 16592 5040 16598 5100
rect 18056 4986 18116 5354
rect 18572 5100 18632 5554
rect 19590 5554 19600 5598
rect 19634 5598 19640 6130
rect 20600 6130 20660 6262
rect 21116 6220 21176 6366
rect 20900 6214 21388 6220
rect 20900 6180 20912 6214
rect 21376 6180 21388 6214
rect 20900 6174 21388 6180
rect 20600 6066 20618 6130
rect 19634 5554 19650 5598
rect 18864 5504 19352 5510
rect 18864 5470 18876 5504
rect 19340 5470 19352 5504
rect 18864 5464 19352 5470
rect 19074 5414 19134 5464
rect 19590 5420 19650 5554
rect 20612 5554 20618 6066
rect 20652 6066 20660 6130
rect 21622 6130 21682 6588
rect 22130 6426 22190 6698
rect 22124 6366 22130 6426
rect 22190 6366 22196 6426
rect 22130 6220 22190 6366
rect 22642 6322 22702 6788
rect 23658 6788 23672 6820
rect 23706 6820 23712 7364
rect 24684 7364 24730 7376
rect 24684 6822 24690 7364
rect 23706 6788 23718 6820
rect 22936 6738 23424 6744
rect 22936 6704 22948 6738
rect 23412 6704 23424 6738
rect 22936 6698 23424 6704
rect 23138 6426 23198 6698
rect 23658 6648 23718 6788
rect 24680 6788 24690 6822
rect 24724 6822 24730 7364
rect 25702 7364 25748 7376
rect 24724 6788 24740 6822
rect 25702 6820 25708 7364
rect 23954 6738 24442 6744
rect 23954 6704 23966 6738
rect 24430 6704 24442 6738
rect 23954 6698 24442 6704
rect 23652 6588 23658 6648
rect 23718 6588 23724 6648
rect 24182 6426 24242 6698
rect 23132 6366 23138 6426
rect 23198 6366 23204 6426
rect 24176 6366 24182 6426
rect 24242 6366 24248 6426
rect 22636 6262 22642 6322
rect 22702 6262 22708 6322
rect 21918 6214 22406 6220
rect 21918 6180 21930 6214
rect 22394 6180 22406 6214
rect 21918 6174 22406 6180
rect 21622 6094 21636 6130
rect 20652 5554 20658 6066
rect 21630 5612 21636 6094
rect 20612 5542 20658 5554
rect 21626 5554 21636 5612
rect 21670 6094 21682 6130
rect 22642 6130 22702 6262
rect 23138 6220 23198 6366
rect 24182 6220 24242 6366
rect 24680 6322 24740 6788
rect 25694 6788 25708 6820
rect 25742 6820 25748 7364
rect 26714 7364 26774 7496
rect 27008 7448 27496 7454
rect 27008 7414 27020 7448
rect 27484 7414 27496 7448
rect 27008 7408 27496 7414
rect 25742 6788 25754 6820
rect 24972 6738 25460 6744
rect 24972 6704 24984 6738
rect 25448 6704 25460 6738
rect 24972 6698 25460 6704
rect 25172 6426 25232 6698
rect 25694 6648 25754 6788
rect 26714 6788 26726 7364
rect 26760 6788 26774 7364
rect 27730 7364 27790 8020
rect 28750 8020 28762 8054
rect 28796 8556 28808 8596
rect 29766 8596 29826 8736
rect 30272 8686 30332 8800
rect 31288 8686 31348 8800
rect 31798 8736 31804 8796
rect 31864 8736 31870 8796
rect 30062 8680 30550 8686
rect 30062 8646 30074 8680
rect 30538 8646 30550 8680
rect 30062 8640 30550 8646
rect 31080 8680 31568 8686
rect 31080 8646 31092 8680
rect 31556 8646 31568 8680
rect 31080 8640 31568 8646
rect 28796 8054 28802 8556
rect 29766 8554 29780 8596
rect 28796 8020 28810 8054
rect 28026 7970 28514 7976
rect 28026 7936 28038 7970
rect 28502 7936 28514 7970
rect 28026 7930 28514 7936
rect 28226 7660 28286 7930
rect 28220 7600 28226 7660
rect 28286 7600 28292 7660
rect 28226 7454 28286 7600
rect 28026 7448 28514 7454
rect 28026 7414 28038 7448
rect 28502 7414 28514 7448
rect 28026 7408 28514 7414
rect 27730 7324 27744 7364
rect 27738 6820 27744 7324
rect 25990 6738 26478 6744
rect 25990 6704 26002 6738
rect 26466 6704 26478 6738
rect 25990 6698 26478 6704
rect 25688 6588 25694 6648
rect 25754 6588 25760 6648
rect 26190 6426 26250 6698
rect 25166 6366 25172 6426
rect 25232 6366 25238 6426
rect 26184 6366 26190 6426
rect 26250 6366 26256 6426
rect 24674 6262 24680 6322
rect 24740 6262 24746 6322
rect 22936 6214 23424 6220
rect 22936 6180 22948 6214
rect 23412 6180 23424 6214
rect 22936 6174 23424 6180
rect 23954 6214 24442 6220
rect 23954 6180 23966 6214
rect 24430 6180 24442 6214
rect 23954 6174 24442 6180
rect 21670 5612 21676 6094
rect 22642 6092 22654 6130
rect 21670 5554 21686 5612
rect 19882 5504 20370 5510
rect 19882 5470 19894 5504
rect 20358 5470 20370 5504
rect 19882 5464 20370 5470
rect 20900 5504 21388 5510
rect 20900 5470 20912 5504
rect 21376 5470 21388 5504
rect 20900 5464 21388 5470
rect 21626 5420 21686 5554
rect 22648 5554 22654 6092
rect 22688 6092 22702 6130
rect 23666 6130 23712 6142
rect 22688 5554 22694 6092
rect 23666 5604 23672 6130
rect 22648 5542 22694 5554
rect 23658 5554 23672 5604
rect 23706 5604 23712 6130
rect 24680 6130 24740 6262
rect 25172 6220 25232 6366
rect 26714 6322 26774 6788
rect 27732 6788 27744 6820
rect 27778 7324 27790 7364
rect 28750 7364 28810 8020
rect 29774 8020 29780 8554
rect 29814 8554 29826 8596
rect 30792 8596 30838 8608
rect 29814 8020 29820 8554
rect 30792 8078 30798 8596
rect 29774 8008 29820 8020
rect 30784 8020 30798 8078
rect 30832 8078 30838 8596
rect 31804 8596 31864 8736
rect 32306 8686 32366 9164
rect 32822 9126 32882 9254
rect 33840 9254 33852 9312
rect 33886 9802 33898 9830
rect 33886 9312 33892 9802
rect 33886 9254 33900 9312
rect 33116 9204 33604 9210
rect 33116 9170 33128 9204
rect 33592 9170 33604 9204
rect 33116 9164 33604 9170
rect 33840 9144 33900 9254
rect 32816 9066 32822 9126
rect 32882 9066 32888 9126
rect 33834 9084 33840 9144
rect 33900 9084 33906 9144
rect 32822 8848 32882 9066
rect 32822 8788 33896 8848
rect 33946 8796 34006 9972
rect 34068 9954 34074 10014
rect 34134 9954 34140 10014
rect 34440 9014 34500 12900
rect 34434 8954 34440 9014
rect 34500 8954 34506 9014
rect 34184 8850 34190 8910
rect 34250 8850 34256 8910
rect 32098 8680 32586 8686
rect 32098 8646 32110 8680
rect 32574 8646 32586 8680
rect 32098 8640 32586 8646
rect 31804 8554 31816 8596
rect 30832 8020 30844 8078
rect 29256 7976 29316 7978
rect 29044 7970 29532 7976
rect 29044 7936 29056 7970
rect 29520 7936 29532 7970
rect 29044 7930 29532 7936
rect 30062 7970 30550 7976
rect 30062 7936 30074 7970
rect 30538 7936 30550 7970
rect 30062 7930 30550 7936
rect 29256 7660 29316 7930
rect 30278 7882 30338 7930
rect 30272 7822 30278 7882
rect 30338 7822 30344 7882
rect 30410 7826 30416 7886
rect 30476 7826 30482 7886
rect 30416 7660 30476 7826
rect 30784 7660 30844 8020
rect 31810 8020 31816 8554
rect 31850 8554 31864 8596
rect 32822 8596 32882 8788
rect 33326 8686 33386 8788
rect 33116 8680 33604 8686
rect 33116 8646 33128 8680
rect 33592 8646 33604 8680
rect 33116 8640 33604 8646
rect 32822 8562 32834 8596
rect 31850 8020 31856 8554
rect 32828 8060 32834 8562
rect 31810 8008 31856 8020
rect 32822 8020 32834 8060
rect 32868 8562 32882 8596
rect 33836 8596 33896 8788
rect 33940 8736 33946 8796
rect 34006 8736 34012 8796
rect 33836 8572 33852 8596
rect 32868 8060 32874 8562
rect 32868 8020 32882 8060
rect 31080 7970 31568 7976
rect 31080 7936 31092 7970
rect 31556 7936 31568 7970
rect 31080 7930 31568 7936
rect 32098 7970 32586 7976
rect 32098 7936 32110 7970
rect 32574 7936 32586 7970
rect 32098 7930 32586 7936
rect 32304 7886 32364 7930
rect 31292 7826 31298 7886
rect 31358 7826 31364 7886
rect 32298 7826 32304 7886
rect 32364 7826 32370 7886
rect 32822 7882 32882 8020
rect 33846 8020 33852 8572
rect 33886 8572 33896 8596
rect 33886 8020 33892 8572
rect 33846 8008 33892 8020
rect 33116 7970 33604 7976
rect 33116 7936 33128 7970
rect 33592 7936 33604 7970
rect 33116 7930 33604 7936
rect 29250 7600 29256 7660
rect 29316 7600 29322 7660
rect 30410 7600 30416 7660
rect 30476 7600 30482 7660
rect 30778 7600 30784 7660
rect 30844 7600 30850 7660
rect 29256 7454 29316 7600
rect 30416 7454 30476 7600
rect 30784 7556 30844 7600
rect 30778 7496 30784 7556
rect 30844 7496 30850 7556
rect 31298 7454 31358 7826
rect 32816 7822 32822 7882
rect 32882 7822 32888 7882
rect 32816 7694 32822 7754
rect 32882 7694 32888 7754
rect 31794 7498 31800 7558
rect 31860 7498 31866 7558
rect 29044 7448 29532 7454
rect 29044 7414 29056 7448
rect 29520 7414 29532 7448
rect 29044 7408 29532 7414
rect 30062 7448 30550 7454
rect 30062 7414 30074 7448
rect 30538 7414 30550 7448
rect 30062 7408 30550 7414
rect 31080 7448 31568 7454
rect 31080 7414 31092 7448
rect 31556 7414 31568 7448
rect 31080 7408 31568 7414
rect 31298 7406 31358 7408
rect 27778 6820 27784 7324
rect 28750 7318 28762 7364
rect 28756 6832 28762 7318
rect 27778 6788 27792 6820
rect 27008 6738 27496 6744
rect 27008 6704 27020 6738
rect 27484 6704 27496 6738
rect 27008 6698 27496 6704
rect 27224 6426 27284 6698
rect 27732 6648 27792 6788
rect 28748 6788 28762 6832
rect 28796 7318 28810 7364
rect 29774 7364 29820 7376
rect 28796 6832 28802 7318
rect 28796 6788 28808 6832
rect 29774 6828 29780 7364
rect 28026 6738 28514 6744
rect 28026 6704 28038 6738
rect 28502 6704 28514 6738
rect 28026 6698 28514 6704
rect 27726 6588 27732 6648
rect 27792 6588 27798 6648
rect 27718 6480 27724 6540
rect 27784 6480 27790 6540
rect 27218 6366 27224 6426
rect 27284 6366 27290 6426
rect 26708 6262 26714 6322
rect 26774 6262 26780 6322
rect 27220 6258 27226 6318
rect 27286 6258 27292 6318
rect 27226 6220 27286 6258
rect 24972 6214 25460 6220
rect 24972 6180 24984 6214
rect 25448 6180 25460 6214
rect 24972 6174 25460 6180
rect 25990 6214 26478 6220
rect 25990 6180 26002 6214
rect 26466 6180 26478 6214
rect 25990 6174 26478 6180
rect 27008 6214 27496 6220
rect 27008 6180 27020 6214
rect 27484 6180 27496 6214
rect 27008 6174 27496 6180
rect 24680 6094 24690 6130
rect 23706 5554 23718 5604
rect 21918 5504 22406 5510
rect 21918 5470 21930 5504
rect 22394 5470 22406 5504
rect 21918 5464 22406 5470
rect 22936 5504 23424 5510
rect 22936 5470 22948 5504
rect 23412 5470 23424 5504
rect 22936 5464 23424 5470
rect 23658 5420 23718 5554
rect 24684 5554 24690 6094
rect 24724 6094 24740 6130
rect 25702 6130 25748 6142
rect 24724 5554 24730 6094
rect 25702 5616 25708 6130
rect 24684 5542 24730 5554
rect 25692 5554 25708 5616
rect 25742 5616 25748 6130
rect 26720 6130 26766 6142
rect 25742 5554 25752 5616
rect 26720 5596 26726 6130
rect 23954 5504 24442 5510
rect 23954 5470 23966 5504
rect 24430 5470 24442 5504
rect 23954 5464 24442 5470
rect 24972 5504 25460 5510
rect 24972 5470 24984 5504
rect 25448 5470 25460 5504
rect 24972 5464 25460 5470
rect 25692 5420 25752 5554
rect 26714 5554 26726 5596
rect 26760 5596 26766 6130
rect 27724 6130 27784 6480
rect 28248 6318 28308 6698
rect 28748 6324 28808 6788
rect 29768 6788 29780 6828
rect 29814 6828 29820 7364
rect 30792 7364 30838 7376
rect 30792 6832 30798 7364
rect 29814 6788 29828 6828
rect 29044 6738 29532 6744
rect 29044 6704 29056 6738
rect 29520 6704 29532 6738
rect 29044 6698 29532 6704
rect 28242 6258 28248 6318
rect 28308 6258 28314 6318
rect 28742 6264 28748 6324
rect 28808 6264 28814 6324
rect 28248 6220 28308 6258
rect 28026 6214 28514 6220
rect 28026 6180 28038 6214
rect 28502 6180 28514 6214
rect 28026 6174 28514 6180
rect 27724 6094 27744 6130
rect 26760 5554 26774 5596
rect 25990 5504 26478 5510
rect 25990 5470 26002 5504
rect 26466 5470 26478 5504
rect 25990 5464 26478 5470
rect 19068 5354 19074 5414
rect 19134 5354 19140 5414
rect 19584 5360 19590 5420
rect 19650 5360 19656 5420
rect 23652 5360 23658 5420
rect 23718 5360 23724 5420
rect 25686 5360 25692 5420
rect 25752 5360 25758 5420
rect 18566 5040 18572 5100
rect 18632 5040 18638 5100
rect 14792 4980 15280 4986
rect 14792 4946 14804 4980
rect 15268 4946 15280 4980
rect 14792 4940 15280 4946
rect 15810 4980 16298 4986
rect 15810 4946 15822 4980
rect 16286 4946 16298 4980
rect 15810 4940 16298 4946
rect 16828 4980 17316 4986
rect 16828 4946 16840 4980
rect 17304 4946 17316 4980
rect 16828 4940 17316 4946
rect 17846 4980 18334 4986
rect 17846 4946 17858 4980
rect 18322 4946 18334 4980
rect 17846 4940 18334 4946
rect 14494 4842 14510 4896
rect 13526 4320 13536 4354
rect 14504 4350 14510 4842
rect 13476 4188 13536 4320
rect 14500 4320 14510 4350
rect 14544 4842 14554 4896
rect 15522 4896 15568 4908
rect 14544 4350 14550 4842
rect 15522 4366 15528 4896
rect 14544 4320 14560 4350
rect 13774 4270 14262 4276
rect 13774 4236 13786 4270
rect 14250 4236 14262 4270
rect 13774 4230 14262 4236
rect 13996 4188 14056 4230
rect 14500 4188 14560 4320
rect 15514 4320 15528 4366
rect 15562 4366 15568 4896
rect 16540 4896 16586 4908
rect 15562 4320 15574 4366
rect 16540 4350 16546 4896
rect 14792 4270 15280 4276
rect 14792 4236 14804 4270
rect 15268 4236 15280 4270
rect 14792 4230 15280 4236
rect 13476 4128 14560 4188
rect 13354 4018 13360 4078
rect 13420 4018 13426 4078
rect 14500 3982 14560 4128
rect 13476 3922 14560 3982
rect 13476 3664 13536 3922
rect 13988 3754 14048 3922
rect 14500 3862 14560 3922
rect 14494 3802 14500 3862
rect 14560 3802 14566 3862
rect 13774 3748 14262 3754
rect 13774 3714 13786 3748
rect 14250 3714 14262 3748
rect 13774 3708 14262 3714
rect 13476 3628 13492 3664
rect 13486 3088 13492 3628
rect 13526 3628 13536 3664
rect 14500 3664 14560 3802
rect 14992 3754 15052 4230
rect 15514 4176 15574 4320
rect 16532 4320 16546 4350
rect 16580 4350 16586 4896
rect 17558 4896 17604 4908
rect 17558 4362 17564 4896
rect 16580 4320 16592 4350
rect 15810 4270 16298 4276
rect 15810 4236 15822 4270
rect 16286 4236 16298 4270
rect 15810 4230 16298 4236
rect 15508 4116 15514 4176
rect 15574 4116 15580 4176
rect 15512 3922 15518 3982
rect 15578 3922 15584 3982
rect 14792 3748 15280 3754
rect 14792 3714 14804 3748
rect 15268 3714 15280 3748
rect 14792 3708 15280 3714
rect 13526 3088 13532 3628
rect 14500 3624 14510 3664
rect 13486 3076 13532 3088
rect 14504 3088 14510 3624
rect 14544 3624 14560 3664
rect 15518 3664 15578 3922
rect 16012 3918 16072 4230
rect 16532 4078 16592 4320
rect 17550 4320 17564 4362
rect 17598 4362 17604 4896
rect 18572 4896 18632 5040
rect 19074 4986 19134 5354
rect 18864 4980 19352 4986
rect 18864 4946 18876 4980
rect 19340 4946 19352 4980
rect 18864 4940 19352 4946
rect 18572 4866 18582 4896
rect 18576 4384 18582 4866
rect 17598 4320 17610 4362
rect 16828 4270 17316 4276
rect 16828 4236 16840 4270
rect 17304 4236 17316 4270
rect 16828 4230 17316 4236
rect 16526 4018 16532 4078
rect 16592 4018 16598 4078
rect 17046 3918 17106 4230
rect 17550 4176 17610 4320
rect 18568 4320 18582 4384
rect 18616 4866 18632 4896
rect 19590 4896 19650 5360
rect 21626 5354 21686 5360
rect 22636 5250 22642 5310
rect 22702 5250 22708 5310
rect 24672 5250 24678 5310
rect 24738 5250 24744 5310
rect 21618 5138 21624 5198
rect 21684 5138 21690 5198
rect 20602 5040 20608 5100
rect 20668 5040 20674 5100
rect 19882 4980 20370 4986
rect 19882 4946 19894 4980
rect 20358 4946 20370 4980
rect 19882 4940 20370 4946
rect 18616 4384 18622 4866
rect 19590 4854 19600 4896
rect 18616 4320 18628 4384
rect 19594 4360 19600 4854
rect 17846 4270 18334 4276
rect 17846 4236 17858 4270
rect 18322 4236 18334 4270
rect 17846 4230 18334 4236
rect 17544 4116 17550 4176
rect 17610 4116 17616 4176
rect 18056 4078 18116 4230
rect 18050 4018 18056 4078
rect 18116 4018 18122 4078
rect 17548 3922 17554 3982
rect 17614 3922 17620 3982
rect 16012 3858 17106 3918
rect 16012 3754 16072 3858
rect 17046 3754 17106 3858
rect 15810 3748 16298 3754
rect 15810 3714 15822 3748
rect 16286 3714 16298 3748
rect 15810 3708 16298 3714
rect 16828 3748 17316 3754
rect 16828 3714 16840 3748
rect 17304 3714 17316 3748
rect 16828 3708 17316 3714
rect 14544 3088 14550 3624
rect 15518 3620 15528 3664
rect 14504 3076 14550 3088
rect 15522 3088 15528 3620
rect 15562 3620 15578 3664
rect 16540 3664 16586 3676
rect 15562 3088 15568 3620
rect 16540 3130 16546 3664
rect 15522 3076 15568 3088
rect 16532 3088 16546 3130
rect 16580 3130 16586 3664
rect 17554 3664 17614 3922
rect 18056 3754 18116 4018
rect 18568 3862 18628 4320
rect 19588 4320 19600 4360
rect 19634 4854 19650 4896
rect 20608 4896 20668 5040
rect 20900 4980 21388 4986
rect 20900 4946 20912 4980
rect 21376 4946 21388 4980
rect 20900 4940 21388 4946
rect 20608 4860 20618 4896
rect 19634 4360 19640 4854
rect 19634 4320 19648 4360
rect 20612 4354 20618 4860
rect 18864 4270 19352 4276
rect 18864 4236 18876 4270
rect 19340 4236 19352 4270
rect 18864 4230 19352 4236
rect 19078 4078 19138 4230
rect 19588 4176 19648 4320
rect 20602 4320 20618 4354
rect 20652 4860 20668 4896
rect 21624 4896 21684 5138
rect 21918 4980 22406 4986
rect 21918 4946 21930 4980
rect 22394 4946 22406 4980
rect 21918 4940 22406 4946
rect 21624 4870 21636 4896
rect 20652 4354 20658 4860
rect 21630 4376 21636 4870
rect 20652 4320 20662 4354
rect 19882 4270 20370 4276
rect 19882 4236 19894 4270
rect 20358 4236 20370 4270
rect 19882 4230 20370 4236
rect 19582 4116 19588 4176
rect 19648 4116 19654 4176
rect 20102 4084 20162 4230
rect 18562 3802 18568 3862
rect 18628 3802 18634 3862
rect 17846 3748 18334 3754
rect 17846 3714 17858 3748
rect 18322 3714 18334 3748
rect 17846 3708 18334 3714
rect 17554 3612 17564 3664
rect 16580 3088 16592 3130
rect 13774 3038 14262 3044
rect 13774 3004 13786 3038
rect 14250 3004 14262 3038
rect 13774 2998 14262 3004
rect 14792 3038 15280 3044
rect 14792 3004 14804 3038
rect 15268 3004 15280 3038
rect 14792 2998 15280 3004
rect 15810 3038 16298 3044
rect 15810 3004 15822 3038
rect 16286 3004 16298 3038
rect 15810 2998 16298 3004
rect 13242 2886 13248 2946
rect 13308 2886 13314 2946
rect 13136 2760 13142 2820
rect 13202 2760 13208 2820
rect 13476 2580 14556 2640
rect 13476 2430 13536 2580
rect 13984 2520 14044 2580
rect 13774 2514 14262 2520
rect 13774 2480 13786 2514
rect 14250 2480 14262 2514
rect 13774 2474 14262 2480
rect 13476 2374 13492 2430
rect 13486 1854 13492 2374
rect 13526 2374 13536 2430
rect 14496 2430 14556 2580
rect 14994 2520 15054 2998
rect 16532 2820 16592 3088
rect 17558 3088 17564 3612
rect 17598 3612 17614 3664
rect 18568 3664 18628 3802
rect 19078 3754 19138 4018
rect 20100 4078 20162 4084
rect 20160 4018 20162 4078
rect 20100 4012 20162 4018
rect 19576 3922 19582 3982
rect 19642 3922 19648 3982
rect 18864 3748 19352 3754
rect 18864 3714 18876 3748
rect 19340 3714 19352 3748
rect 18864 3708 19352 3714
rect 18568 3624 18582 3664
rect 17598 3088 17604 3612
rect 18576 3142 18582 3624
rect 17558 3076 17604 3088
rect 18570 3088 18582 3142
rect 18616 3624 18628 3664
rect 19582 3664 19642 3922
rect 20102 3754 20162 4012
rect 20602 3862 20662 4320
rect 21620 4320 21636 4376
rect 21670 4870 21684 4896
rect 22642 4896 22702 5250
rect 22936 4980 23424 4986
rect 22936 4946 22948 4980
rect 23412 4946 23424 4980
rect 22936 4940 23424 4946
rect 23954 4980 24442 4986
rect 23954 4946 23966 4980
rect 24430 4946 24442 4980
rect 23954 4940 24442 4946
rect 21670 4376 21676 4870
rect 22642 4864 22654 4896
rect 21670 4320 21680 4376
rect 20900 4270 21388 4276
rect 20900 4236 20912 4270
rect 21376 4236 21388 4270
rect 20900 4230 21388 4236
rect 21104 4078 21164 4230
rect 21450 4196 21510 4202
rect 21620 4196 21680 4320
rect 22648 4320 22654 4864
rect 22688 4864 22702 4896
rect 23666 4896 23712 4908
rect 22688 4320 22694 4864
rect 23666 4390 23672 4896
rect 22648 4308 22694 4320
rect 23662 4320 23672 4390
rect 23706 4390 23712 4896
rect 24678 4896 24738 5250
rect 26220 5212 26280 5464
rect 26714 5422 26774 5554
rect 27738 5554 27744 6094
rect 27778 5554 27784 6130
rect 28748 6130 28808 6264
rect 29226 6220 29286 6698
rect 29768 6648 29828 6788
rect 30782 6788 30798 6832
rect 30832 6832 30838 7364
rect 31800 7364 31860 7498
rect 32098 7448 32586 7454
rect 32098 7414 32110 7448
rect 32574 7414 32586 7448
rect 32098 7408 32586 7414
rect 31800 7314 31816 7364
rect 30832 6788 30842 6832
rect 31810 6816 31816 7314
rect 30062 6738 30550 6744
rect 30062 6704 30074 6738
rect 30538 6704 30550 6738
rect 30062 6698 30550 6704
rect 29762 6588 29768 6648
rect 29828 6588 29834 6648
rect 29758 6480 29764 6540
rect 29824 6480 29830 6540
rect 29044 6214 29532 6220
rect 29044 6180 29056 6214
rect 29520 6180 29532 6214
rect 29044 6174 29532 6180
rect 28748 6036 28762 6130
rect 28756 5596 28762 6036
rect 27738 5542 27784 5554
rect 28748 5554 28762 5596
rect 28796 6036 28808 6130
rect 29764 6130 29824 6480
rect 30250 6366 30256 6426
rect 30316 6366 30322 6426
rect 30256 6220 30316 6366
rect 30782 6324 30842 6788
rect 31806 6788 31816 6816
rect 31850 7314 31860 7364
rect 32822 7364 32882 7694
rect 33116 7448 33604 7454
rect 33116 7414 33128 7448
rect 33592 7414 33604 7448
rect 33116 7408 33604 7414
rect 31850 6816 31856 7314
rect 32822 7312 32834 7364
rect 32828 6816 32834 7312
rect 31850 6788 31866 6816
rect 31080 6738 31568 6744
rect 31080 6704 31092 6738
rect 31556 6704 31568 6738
rect 31080 6698 31568 6704
rect 31806 6648 31866 6788
rect 32822 6788 32834 6816
rect 32868 7312 32882 7364
rect 33846 7364 33892 7376
rect 32868 6816 32874 7312
rect 33846 6822 33852 7364
rect 32868 6788 32882 6816
rect 32098 6738 32586 6744
rect 32098 6704 32110 6738
rect 32574 6704 32586 6738
rect 32098 6698 32586 6704
rect 31800 6588 31806 6648
rect 31866 6588 31872 6648
rect 31796 6480 31802 6540
rect 31862 6480 31868 6540
rect 31288 6366 31294 6426
rect 31354 6366 31360 6426
rect 30776 6264 30782 6324
rect 30842 6264 30848 6324
rect 31294 6220 31354 6366
rect 30062 6214 30550 6220
rect 30062 6180 30074 6214
rect 30538 6180 30550 6214
rect 30062 6174 30550 6180
rect 31080 6214 31568 6220
rect 31080 6180 31092 6214
rect 31556 6180 31568 6214
rect 31080 6174 31568 6180
rect 29764 6064 29780 6130
rect 28796 5596 28802 6036
rect 28796 5554 28808 5596
rect 27008 5504 27496 5510
rect 27008 5470 27020 5504
rect 27484 5470 27496 5504
rect 27008 5464 27496 5470
rect 28026 5504 28514 5510
rect 28026 5470 28038 5504
rect 28502 5470 28514 5504
rect 28026 5464 28514 5470
rect 26708 5362 26714 5422
rect 26774 5362 26780 5422
rect 27062 5362 27068 5422
rect 27128 5362 27134 5422
rect 26704 5250 26710 5310
rect 26770 5250 26776 5310
rect 26214 5152 26220 5212
rect 26280 5152 26286 5212
rect 24972 4980 25460 4986
rect 24972 4946 24984 4980
rect 25448 4946 25460 4980
rect 24972 4940 25460 4946
rect 25990 4980 26478 4986
rect 25990 4946 26002 4980
rect 26466 4946 26478 4980
rect 25990 4940 26478 4946
rect 24678 4858 24690 4896
rect 23706 4320 23722 4390
rect 21918 4270 22406 4276
rect 21918 4236 21930 4270
rect 22394 4236 22406 4270
rect 21918 4230 22406 4236
rect 22936 4270 23424 4276
rect 22936 4236 22948 4270
rect 23412 4236 23424 4270
rect 22936 4230 23424 4236
rect 21614 4136 21620 4196
rect 21680 4136 21686 4196
rect 21098 4018 21104 4078
rect 21164 4018 21170 4078
rect 20596 3802 20602 3862
rect 20662 3802 20668 3862
rect 19882 3748 20370 3754
rect 19882 3714 19894 3748
rect 20358 3714 20370 3748
rect 19882 3708 20370 3714
rect 18616 3142 18622 3624
rect 19582 3604 19600 3664
rect 18616 3088 18630 3142
rect 16828 3038 17316 3044
rect 16828 3004 16840 3038
rect 17304 3004 17316 3038
rect 16828 2998 17316 3004
rect 17846 3038 18334 3044
rect 17846 3004 17858 3038
rect 18322 3004 18334 3038
rect 17846 2998 18334 3004
rect 17052 2832 17112 2998
rect 16526 2760 16532 2820
rect 16592 2760 16598 2820
rect 17046 2772 17052 2832
rect 17112 2772 17118 2832
rect 15508 2658 15514 2718
rect 15574 2658 15580 2718
rect 17544 2658 17550 2718
rect 17610 2658 17616 2718
rect 14792 2514 15280 2520
rect 14792 2480 14804 2514
rect 15268 2480 15280 2514
rect 14792 2474 15280 2480
rect 13526 1854 13532 2374
rect 13486 1842 13532 1854
rect 14496 1854 14510 2430
rect 14544 1854 14556 2430
rect 15514 2430 15574 2658
rect 16526 2554 16532 2614
rect 16592 2554 16598 2614
rect 15810 2514 16298 2520
rect 15810 2480 15822 2514
rect 16286 2480 16298 2514
rect 15810 2474 16298 2480
rect 15514 2370 15528 2430
rect 15522 1890 15528 2370
rect 13774 1804 14262 1810
rect 13774 1770 13786 1804
rect 14250 1770 14262 1804
rect 13774 1764 14262 1770
rect 13354 1656 13360 1716
rect 13420 1656 13426 1716
rect 13026 1552 13032 1612
rect 13092 1552 13098 1612
rect 13360 1386 13420 1656
rect 14496 1612 14556 1854
rect 15516 1854 15528 1890
rect 15562 2370 15574 2430
rect 16532 2430 16592 2554
rect 16828 2514 17316 2520
rect 16828 2480 16840 2514
rect 17304 2480 17316 2514
rect 16828 2474 17316 2480
rect 16532 2376 16546 2430
rect 15562 1890 15568 2370
rect 16540 1894 16546 2376
rect 15562 1854 15576 1890
rect 14792 1804 15280 1810
rect 14792 1770 14804 1804
rect 15268 1770 15280 1804
rect 14792 1764 15280 1770
rect 14490 1552 14496 1612
rect 14556 1552 14562 1612
rect 15004 1506 15064 1764
rect 14998 1446 15004 1506
rect 15064 1446 15070 1506
rect 13360 1326 14560 1386
rect 11976 492 11982 552
rect 12042 492 12048 552
rect 13360 474 13420 1326
rect 13480 1198 13540 1326
rect 13966 1288 14026 1326
rect 13774 1282 14262 1288
rect 13774 1248 13786 1282
rect 14250 1248 14262 1282
rect 13774 1242 14262 1248
rect 13480 1126 13492 1198
rect 13486 622 13492 1126
rect 13526 1126 13540 1198
rect 14500 1198 14560 1326
rect 15004 1288 15064 1446
rect 15516 1396 15576 1854
rect 16530 1854 16546 1894
rect 16580 2376 16592 2430
rect 17550 2430 17610 2658
rect 18052 2520 18112 2998
rect 18570 2718 18630 3088
rect 19594 3088 19600 3604
rect 19634 3604 19642 3664
rect 20602 3664 20662 3802
rect 21104 3754 21164 4018
rect 21450 3982 21510 4136
rect 21444 3922 21450 3982
rect 21510 3922 21516 3982
rect 21620 3928 21626 3988
rect 21686 3928 21692 3988
rect 20900 3748 21388 3754
rect 20900 3714 20912 3748
rect 21376 3714 21388 3748
rect 20900 3708 21388 3714
rect 20602 3624 20618 3664
rect 19634 3088 19640 3604
rect 20612 3154 20618 3624
rect 19594 3076 19640 3088
rect 20606 3088 20618 3154
rect 20652 3624 20662 3664
rect 21626 3664 21686 3928
rect 22142 3926 22202 4230
rect 23156 4090 23216 4230
rect 23662 4196 23722 4320
rect 24684 4320 24690 4858
rect 24724 4858 24738 4896
rect 25702 4896 25748 4908
rect 24724 4320 24730 4858
rect 25702 4390 25708 4896
rect 24684 4308 24730 4320
rect 25694 4320 25708 4390
rect 25742 4390 25748 4896
rect 26710 4896 26770 5250
rect 27068 5104 27128 5362
rect 27258 5212 27318 5464
rect 28234 5212 28294 5464
rect 27252 5152 27258 5212
rect 27318 5152 27324 5212
rect 28228 5152 28234 5212
rect 28294 5152 28300 5212
rect 28748 5100 28808 5554
rect 29774 5554 29780 6064
rect 29814 6064 29824 6130
rect 30792 6130 30838 6142
rect 29814 5554 29820 6064
rect 30792 5598 30798 6130
rect 29774 5542 29820 5554
rect 30786 5554 30798 5598
rect 30832 5598 30838 6130
rect 31802 6130 31862 6480
rect 32320 6426 32380 6698
rect 32822 6606 32882 6788
rect 33836 6788 33852 6822
rect 33886 6822 33892 7364
rect 33886 6788 33896 6822
rect 33116 6738 33604 6744
rect 33116 6704 33128 6738
rect 33592 6704 33604 6738
rect 33116 6698 33604 6704
rect 33330 6606 33390 6698
rect 33836 6606 33896 6788
rect 32822 6546 33896 6606
rect 32314 6366 32320 6426
rect 32380 6366 32386 6426
rect 32818 6264 32824 6324
rect 32884 6264 32890 6324
rect 32098 6214 32586 6220
rect 32098 6180 32110 6214
rect 32574 6180 32586 6214
rect 32098 6174 32586 6180
rect 31802 6078 31816 6130
rect 31810 5604 31816 6078
rect 30832 5554 30846 5598
rect 29044 5504 29532 5510
rect 29044 5470 29056 5504
rect 29520 5470 29532 5504
rect 29044 5464 29532 5470
rect 30062 5504 30550 5510
rect 30062 5470 30074 5504
rect 30538 5470 30550 5504
rect 30062 5464 30550 5470
rect 29250 5212 29310 5464
rect 30786 5422 30846 5554
rect 31804 5554 31816 5604
rect 31850 6078 31862 6130
rect 32824 6130 32884 6264
rect 33116 6214 33604 6220
rect 33116 6180 33128 6214
rect 33592 6180 33604 6214
rect 33116 6174 33604 6180
rect 32824 6096 32834 6130
rect 31850 5604 31856 6078
rect 31850 5554 31864 5604
rect 32828 5598 32834 6096
rect 31080 5504 31568 5510
rect 31080 5470 31092 5504
rect 31556 5470 31568 5504
rect 31080 5464 31568 5470
rect 30780 5362 30786 5422
rect 30846 5362 30852 5422
rect 29244 5152 29250 5212
rect 29310 5152 29316 5212
rect 31270 5152 31276 5212
rect 31336 5152 31342 5212
rect 27068 5038 27128 5044
rect 28742 5040 28748 5100
rect 28808 5040 28814 5100
rect 30778 5040 30784 5100
rect 30844 5040 30850 5100
rect 27008 4980 27496 4986
rect 27008 4946 27020 4980
rect 27484 4946 27496 4980
rect 27008 4940 27496 4946
rect 28026 4980 28514 4986
rect 28026 4946 28038 4980
rect 28502 4946 28514 4980
rect 28026 4940 28514 4946
rect 26710 4854 26726 4896
rect 25742 4320 25754 4390
rect 23954 4270 24442 4276
rect 23954 4236 23966 4270
rect 24430 4236 24442 4270
rect 23954 4230 24442 4236
rect 24972 4270 25460 4276
rect 24972 4236 24984 4270
rect 25448 4236 25460 4270
rect 24972 4230 25460 4236
rect 23656 4136 23662 4196
rect 23722 4136 23728 4196
rect 24178 4090 24238 4230
rect 25192 4090 25252 4230
rect 25694 4196 25754 4320
rect 26720 4320 26726 4854
rect 26760 4854 26770 4896
rect 27738 4896 27784 4908
rect 26760 4320 26766 4854
rect 27738 4356 27744 4896
rect 26720 4308 26766 4320
rect 27734 4320 27744 4356
rect 27778 4356 27784 4896
rect 28748 4896 28808 5040
rect 29044 4980 29532 4986
rect 29044 4946 29056 4980
rect 29520 4946 29532 4980
rect 29044 4940 29532 4946
rect 30062 4980 30550 4986
rect 30062 4946 30074 4980
rect 30538 4946 30550 4980
rect 30062 4940 30550 4946
rect 28748 4858 28762 4896
rect 28756 4372 28762 4858
rect 27778 4320 27794 4356
rect 25990 4270 26478 4276
rect 25990 4236 26002 4270
rect 26466 4236 26478 4270
rect 25990 4230 26478 4236
rect 27008 4270 27496 4276
rect 27008 4236 27020 4270
rect 27484 4236 27496 4270
rect 27008 4230 27496 4236
rect 25688 4136 25694 4196
rect 25754 4136 25760 4196
rect 26194 4190 26254 4230
rect 27220 4190 27280 4230
rect 27734 4196 27794 4320
rect 28752 4320 28762 4372
rect 28796 4858 28808 4896
rect 29774 4896 29820 4908
rect 28796 4372 28802 4858
rect 28796 4320 28812 4372
rect 29774 4364 29780 4896
rect 28026 4270 28514 4276
rect 28026 4236 28038 4270
rect 28502 4236 28514 4270
rect 28026 4230 28514 4236
rect 26194 4130 27280 4190
rect 27728 4136 27734 4196
rect 27794 4136 27800 4196
rect 26194 4090 26254 4130
rect 23156 4030 26254 4090
rect 26706 4038 26712 4098
rect 26772 4038 26778 4098
rect 23156 3926 23216 4030
rect 23648 3928 23654 3988
rect 23714 3928 23720 3988
rect 22142 3866 23216 3926
rect 22142 3754 22202 3866
rect 23156 3754 23216 3866
rect 21918 3748 22406 3754
rect 21918 3714 21930 3748
rect 22394 3714 22406 3748
rect 21918 3708 22406 3714
rect 22936 3748 23424 3754
rect 22936 3714 22948 3748
rect 23412 3714 23424 3748
rect 22936 3708 23424 3714
rect 20652 3154 20658 3624
rect 21626 3620 21636 3664
rect 20652 3088 20666 3154
rect 21630 3146 21636 3620
rect 18864 3038 19352 3044
rect 18864 3004 18876 3038
rect 19340 3004 19352 3038
rect 18864 2998 19352 3004
rect 19882 3038 20370 3044
rect 19882 3004 19894 3038
rect 20358 3004 20370 3038
rect 19882 2998 20370 3004
rect 18564 2658 18570 2718
rect 18630 2658 18636 2718
rect 19074 2520 19134 2998
rect 19580 2658 19586 2718
rect 19646 2658 19652 2718
rect 17846 2514 18334 2520
rect 17846 2480 17858 2514
rect 18322 2480 18334 2514
rect 17846 2474 18334 2480
rect 18864 2514 19352 2520
rect 18864 2480 18876 2514
rect 19340 2480 19352 2514
rect 18864 2474 19352 2480
rect 17550 2380 17564 2430
rect 16580 1894 16586 2376
rect 16580 1854 16590 1894
rect 17558 1878 17564 2380
rect 15810 1804 16298 1810
rect 15810 1770 15822 1804
rect 16286 1770 16298 1804
rect 15810 1764 16298 1770
rect 16024 1506 16084 1764
rect 16530 1716 16590 1854
rect 17552 1854 17564 1878
rect 17598 2380 17610 2430
rect 18576 2430 18622 2442
rect 17598 1878 17604 2380
rect 17598 1854 17612 1878
rect 18576 1868 18582 2430
rect 16828 1804 17316 1810
rect 16828 1770 16840 1804
rect 17304 1770 17316 1804
rect 16828 1764 17316 1770
rect 16524 1656 16530 1716
rect 16590 1656 16596 1716
rect 16530 1552 16536 1612
rect 16596 1552 16602 1612
rect 16018 1446 16024 1506
rect 16084 1446 16090 1506
rect 15510 1336 15516 1396
rect 15576 1336 15582 1396
rect 14792 1282 15280 1288
rect 14792 1248 14804 1282
rect 15268 1248 15280 1282
rect 14792 1242 15280 1248
rect 13526 622 13532 1126
rect 14500 1122 14510 1198
rect 14504 670 14510 1122
rect 13486 610 13532 622
rect 14496 622 14510 670
rect 14544 1122 14560 1198
rect 15516 1198 15576 1336
rect 16024 1288 16084 1446
rect 15810 1282 16298 1288
rect 15810 1248 15822 1282
rect 16286 1248 16298 1282
rect 15810 1242 16298 1248
rect 14544 670 14550 1122
rect 14544 622 14556 670
rect 13774 572 14262 578
rect 13774 538 13786 572
rect 14250 538 14262 572
rect 13774 532 14262 538
rect 14496 474 14556 622
rect 15516 622 15528 1198
rect 15562 622 15576 1198
rect 16536 1198 16596 1552
rect 17048 1506 17108 1764
rect 17042 1446 17048 1506
rect 17108 1446 17114 1506
rect 17048 1288 17108 1446
rect 17552 1396 17612 1854
rect 18566 1854 18582 1868
rect 18616 1868 18622 2430
rect 19586 2430 19646 2658
rect 20086 2520 20146 2998
rect 20606 2718 20666 3088
rect 21618 3088 21636 3146
rect 21670 3620 21686 3664
rect 22648 3664 22694 3676
rect 21670 3146 21676 3620
rect 21670 3088 21678 3146
rect 22648 3140 22654 3664
rect 20900 3038 21388 3044
rect 20900 3004 20912 3038
rect 21376 3004 21388 3038
rect 20900 2998 21388 3004
rect 20600 2658 20606 2718
rect 20666 2658 20672 2718
rect 21116 2520 21176 2998
rect 21618 2886 21678 3088
rect 22636 3088 22654 3140
rect 22688 3140 22694 3664
rect 23654 3664 23714 3928
rect 24178 3754 24238 4030
rect 25192 3754 25252 4030
rect 25692 3928 25698 3988
rect 25758 3928 25764 3988
rect 23954 3748 24442 3754
rect 23954 3714 23966 3748
rect 24430 3714 24442 3748
rect 23954 3708 24442 3714
rect 24972 3748 25460 3754
rect 24972 3714 24984 3748
rect 25448 3714 25460 3748
rect 24972 3708 25460 3714
rect 23654 3620 23672 3664
rect 22688 3088 22696 3140
rect 21918 3038 22406 3044
rect 21918 3004 21930 3038
rect 22394 3004 22406 3038
rect 21918 2998 22406 3004
rect 21468 2826 21678 2886
rect 22132 2832 22192 2998
rect 22636 2946 22696 3088
rect 23666 3088 23672 3620
rect 23706 3620 23714 3664
rect 24684 3664 24730 3676
rect 23706 3088 23712 3620
rect 24684 3140 24690 3664
rect 23666 3076 23712 3088
rect 24678 3088 24690 3140
rect 24724 3140 24730 3664
rect 25698 3664 25758 3928
rect 26194 3754 26254 4030
rect 25990 3748 26478 3754
rect 25990 3714 26002 3748
rect 26466 3714 26478 3748
rect 25990 3708 26478 3714
rect 25698 3616 25708 3664
rect 24724 3088 24738 3140
rect 22936 3038 23424 3044
rect 22936 3004 22948 3038
rect 23412 3004 23424 3038
rect 22936 2998 23424 3004
rect 23954 3038 24442 3044
rect 23954 3004 23966 3038
rect 24430 3004 24442 3038
rect 23954 2998 24442 3004
rect 24678 2946 24738 3088
rect 25702 3088 25708 3616
rect 25742 3616 25758 3664
rect 26712 3664 26772 4038
rect 27220 3754 27280 4130
rect 27720 3928 27726 3988
rect 27786 3928 27792 3988
rect 27008 3748 27496 3754
rect 27008 3714 27020 3748
rect 27484 3714 27496 3748
rect 27008 3708 27496 3714
rect 26712 3628 26726 3664
rect 25742 3088 25748 3616
rect 26720 3132 26726 3628
rect 25702 3076 25748 3088
rect 26714 3088 26726 3132
rect 26760 3628 26772 3664
rect 27726 3664 27786 3928
rect 28240 3754 28300 4230
rect 28752 3862 28812 4320
rect 29764 4320 29780 4364
rect 29814 4364 29820 4896
rect 30784 4896 30844 5040
rect 31276 4986 31336 5152
rect 31080 4980 31568 4986
rect 31080 4946 31092 4980
rect 31556 4946 31568 4980
rect 31080 4940 31568 4946
rect 30784 4838 30798 4896
rect 29814 4320 29824 4364
rect 30792 4360 30798 4838
rect 29044 4270 29532 4276
rect 29044 4236 29056 4270
rect 29520 4236 29532 4270
rect 29044 4230 29532 4236
rect 28746 3802 28752 3862
rect 28812 3802 28818 3862
rect 28026 3748 28514 3754
rect 28026 3714 28038 3748
rect 28502 3714 28514 3748
rect 28026 3708 28514 3714
rect 26760 3132 26766 3628
rect 27726 3616 27744 3664
rect 26760 3088 26774 3132
rect 27738 3128 27744 3616
rect 24972 3038 25460 3044
rect 24972 3004 24984 3038
rect 25448 3004 25460 3038
rect 24972 2998 25460 3004
rect 25990 3038 26478 3044
rect 25990 3004 26002 3038
rect 26466 3004 26478 3038
rect 25990 2998 26478 3004
rect 26714 2946 26774 3088
rect 27728 3088 27744 3128
rect 27778 3616 27786 3664
rect 28752 3664 28812 3802
rect 29256 3754 29316 4230
rect 29764 3988 29824 4320
rect 30782 4320 30798 4360
rect 30832 4838 30844 4896
rect 31804 4896 31864 5554
rect 32820 5554 32834 5598
rect 32868 6096 32884 6130
rect 33846 6130 33892 6142
rect 32868 5598 32874 6096
rect 32868 5554 32880 5598
rect 33846 5584 33852 6130
rect 32098 5504 32586 5510
rect 32098 5470 32110 5504
rect 32574 5470 32586 5504
rect 32098 5464 32586 5470
rect 32306 5212 32366 5464
rect 32820 5372 32880 5554
rect 33836 5554 33852 5584
rect 33886 5584 33892 6130
rect 33886 5554 33896 5584
rect 33116 5504 33604 5510
rect 33116 5470 33128 5504
rect 33592 5470 33604 5504
rect 33116 5464 33604 5470
rect 33326 5372 33386 5464
rect 33836 5372 33896 5554
rect 32820 5312 33896 5372
rect 32300 5152 32306 5212
rect 32366 5152 32372 5212
rect 32820 5100 32880 5312
rect 32814 5040 32820 5100
rect 32880 5040 32886 5100
rect 32098 4980 32586 4986
rect 32098 4946 32110 4980
rect 32574 4946 32586 4980
rect 32098 4940 32586 4946
rect 33116 4980 33604 4986
rect 33116 4946 33128 4980
rect 33592 4946 33604 4980
rect 33116 4940 33604 4946
rect 31804 4854 31816 4896
rect 30832 4360 30838 4838
rect 31810 4374 31816 4854
rect 30832 4320 30842 4360
rect 30062 4270 30550 4276
rect 30062 4236 30074 4270
rect 30538 4236 30550 4270
rect 30062 4230 30550 4236
rect 29758 3928 29764 3988
rect 29824 3928 29830 3988
rect 30290 3754 30350 4230
rect 30782 3862 30842 4320
rect 31804 4320 31816 4374
rect 31850 4854 31864 4896
rect 32828 4896 32874 4908
rect 31850 4374 31856 4854
rect 31850 4320 31864 4374
rect 32828 4366 32834 4896
rect 31080 4270 31568 4276
rect 31080 4236 31092 4270
rect 31556 4236 31568 4270
rect 31080 4230 31568 4236
rect 31308 3864 31368 4230
rect 31804 3988 31864 4320
rect 32818 4320 32834 4366
rect 32868 4366 32874 4896
rect 33846 4896 33892 4908
rect 32868 4320 32878 4366
rect 33846 4348 33852 4896
rect 32098 4270 32586 4276
rect 32098 4236 32110 4270
rect 32574 4236 32586 4270
rect 32098 4230 32586 4236
rect 32322 3992 32382 4230
rect 32818 4194 32878 4320
rect 33838 4320 33852 4348
rect 33886 4348 33892 4896
rect 33886 4320 33898 4348
rect 33116 4270 33604 4276
rect 33116 4236 33128 4270
rect 33592 4236 33604 4270
rect 33116 4230 33604 4236
rect 33324 4196 33384 4230
rect 33838 4196 33898 4320
rect 33324 4194 33898 4196
rect 32818 4134 33898 4194
rect 32818 4098 32878 4134
rect 32812 4038 32818 4098
rect 32878 4038 32884 4098
rect 31798 3928 31804 3988
rect 31864 3928 31870 3988
rect 32316 3932 32322 3992
rect 32382 3932 32388 3992
rect 33828 3932 33834 3992
rect 33894 3932 33900 3992
rect 30776 3802 30782 3862
rect 30842 3802 30848 3862
rect 29044 3748 29532 3754
rect 29044 3714 29056 3748
rect 29520 3714 29532 3748
rect 29044 3708 29532 3714
rect 30062 3748 30550 3754
rect 30062 3714 30074 3748
rect 30538 3714 30550 3748
rect 30062 3708 30550 3714
rect 28752 3618 28762 3664
rect 27778 3128 27784 3616
rect 28756 3148 28762 3618
rect 27778 3088 27788 3128
rect 27008 3038 27496 3044
rect 27008 3004 27020 3038
rect 27484 3004 27496 3038
rect 27008 2998 27496 3004
rect 22630 2886 22636 2946
rect 22696 2886 22702 2946
rect 24672 2886 24678 2946
rect 24738 2886 24744 2946
rect 26708 2886 26714 2946
rect 26774 2886 26780 2946
rect 27220 2836 27280 2998
rect 27728 2938 27788 3088
rect 28750 3088 28762 3148
rect 28796 3618 28812 3664
rect 29774 3664 29820 3676
rect 28796 3148 28802 3618
rect 28796 3088 28810 3148
rect 29774 3132 29780 3664
rect 28026 3038 28514 3044
rect 28026 3004 28038 3038
rect 28502 3004 28514 3038
rect 28026 2998 28514 3004
rect 27728 2878 27934 2938
rect 21468 2614 21528 2826
rect 22126 2772 22132 2832
rect 22192 2772 22198 2832
rect 27214 2776 27220 2836
rect 27280 2776 27286 2836
rect 21618 2658 21624 2718
rect 21684 2658 21690 2718
rect 23648 2658 23654 2718
rect 23714 2658 23720 2718
rect 25686 2658 25692 2718
rect 25752 2658 25758 2718
rect 27722 2658 27728 2718
rect 27788 2658 27794 2718
rect 21462 2554 21468 2614
rect 21528 2554 21534 2614
rect 19882 2514 20370 2520
rect 19882 2480 19894 2514
rect 20358 2480 20370 2514
rect 19882 2474 20370 2480
rect 20900 2514 21388 2520
rect 20900 2480 20912 2514
rect 21376 2480 21388 2514
rect 20900 2474 21388 2480
rect 19586 1948 19600 2430
rect 19594 1874 19600 1948
rect 18616 1854 18626 1868
rect 17846 1804 18334 1810
rect 17846 1770 17858 1804
rect 18322 1770 18334 1804
rect 17846 1764 18334 1770
rect 18066 1506 18126 1764
rect 18566 1612 18626 1854
rect 19590 1854 19600 1874
rect 19634 1948 19646 2430
rect 20612 2430 20658 2442
rect 19634 1874 19640 1948
rect 20612 1880 20618 2430
rect 19634 1854 19650 1874
rect 18864 1804 19352 1810
rect 18864 1770 18876 1804
rect 19340 1770 19352 1804
rect 18864 1764 19352 1770
rect 18560 1552 18566 1612
rect 18626 1552 18632 1612
rect 19080 1506 19140 1764
rect 18060 1446 18066 1506
rect 18126 1446 18132 1506
rect 19074 1446 19080 1506
rect 19140 1446 19146 1506
rect 17546 1336 17552 1396
rect 17612 1336 17618 1396
rect 16828 1282 17316 1288
rect 16828 1248 16840 1282
rect 17304 1248 17316 1282
rect 16828 1242 17316 1248
rect 16536 1184 16546 1198
rect 14792 572 15280 578
rect 14792 538 14804 572
rect 15268 538 15280 572
rect 14792 532 15280 538
rect 13354 414 13360 474
rect 13420 414 13426 474
rect 14490 414 14496 474
rect 14556 414 14562 474
rect 15008 366 15068 532
rect 15002 306 15008 366
rect 15068 306 15074 366
rect 15516 110 15576 622
rect 16540 622 16546 1184
rect 16580 1184 16596 1198
rect 17552 1198 17612 1336
rect 18066 1288 18126 1446
rect 19080 1288 19140 1446
rect 19590 1396 19650 1854
rect 20606 1854 20618 1880
rect 20652 1880 20658 2430
rect 21624 2430 21684 2658
rect 21918 2514 22406 2520
rect 21918 2480 21930 2514
rect 22394 2480 22406 2514
rect 21918 2474 22406 2480
rect 22936 2514 23424 2520
rect 22936 2480 22948 2514
rect 23412 2480 23424 2514
rect 22936 2474 23424 2480
rect 22648 2430 22694 2442
rect 23654 2430 23714 2658
rect 23954 2514 24442 2520
rect 23954 2480 23966 2514
rect 24430 2480 24442 2514
rect 23954 2474 24442 2480
rect 24972 2514 25460 2520
rect 24972 2480 24984 2514
rect 25448 2480 25460 2514
rect 24972 2474 25460 2480
rect 24684 2430 24730 2442
rect 25692 2430 25752 2658
rect 25990 2514 26478 2520
rect 25990 2480 26002 2514
rect 26466 2480 26478 2514
rect 25990 2474 26478 2480
rect 27008 2514 27496 2520
rect 27008 2480 27020 2514
rect 27484 2480 27496 2514
rect 27008 2474 27496 2480
rect 21624 2374 21636 2430
rect 20652 1854 20666 1880
rect 21630 1878 21636 2374
rect 19882 1804 20370 1810
rect 19882 1770 19894 1804
rect 20358 1770 20370 1804
rect 19882 1764 20370 1770
rect 20112 1506 20172 1764
rect 20606 1612 20666 1854
rect 21628 1854 21636 1878
rect 21670 2374 21684 2430
rect 22642 2394 22654 2430
rect 21670 1878 21676 2374
rect 22648 1906 22654 2394
rect 21670 1854 21688 1878
rect 20900 1804 21388 1810
rect 20900 1770 20912 1804
rect 21376 1770 21388 1804
rect 20900 1764 21388 1770
rect 20754 1658 20760 1718
rect 20820 1658 20826 1718
rect 20600 1552 20606 1612
rect 20666 1552 20672 1612
rect 20106 1446 20112 1506
rect 20172 1446 20178 1506
rect 20760 1474 20820 1658
rect 21124 1506 21184 1764
rect 19584 1336 19590 1396
rect 19650 1336 19656 1396
rect 17846 1282 18334 1288
rect 17846 1248 17858 1282
rect 18322 1248 18334 1282
rect 17846 1242 18334 1248
rect 18864 1282 19352 1288
rect 18864 1248 18876 1282
rect 19340 1248 19352 1282
rect 18864 1242 19352 1248
rect 16580 622 16586 1184
rect 16540 610 16586 622
rect 17552 622 17564 1198
rect 17598 622 17612 1198
rect 18576 1198 18622 1210
rect 18576 664 18582 1198
rect 15810 572 16298 578
rect 15810 538 15822 572
rect 16286 538 16298 572
rect 15810 532 16298 538
rect 16828 572 17316 578
rect 16828 538 16840 572
rect 17304 538 17316 572
rect 16828 532 17316 538
rect 16022 366 16082 532
rect 16022 300 16082 306
rect 17044 366 17104 532
rect 17044 300 17104 306
rect 17552 110 17612 622
rect 18566 622 18582 664
rect 18616 664 18622 1198
rect 19590 1198 19650 1336
rect 20112 1288 20172 1446
rect 20604 1414 20820 1474
rect 21118 1446 21124 1506
rect 21184 1446 21190 1506
rect 19882 1282 20370 1288
rect 19882 1248 19894 1282
rect 20358 1248 20370 1282
rect 19882 1242 20370 1248
rect 18616 622 18626 664
rect 17846 572 18334 578
rect 17846 538 17858 572
rect 18322 538 18334 572
rect 17846 532 18334 538
rect 18056 372 18116 532
rect 18566 474 18626 622
rect 19590 622 19600 1198
rect 19634 622 19650 1198
rect 20604 1198 20664 1414
rect 21124 1288 21184 1446
rect 21628 1396 21688 1854
rect 22638 1854 22654 1906
rect 22688 2394 22702 2430
rect 22688 1906 22694 2394
rect 23654 2380 23672 2430
rect 22688 1854 22698 1906
rect 23666 1884 23672 2380
rect 21918 1804 22406 1810
rect 21918 1770 21930 1804
rect 22394 1770 22406 1804
rect 21918 1764 22406 1770
rect 22132 1506 22192 1764
rect 22638 1718 22698 1854
rect 23664 1854 23672 1884
rect 23706 2380 23714 2430
rect 24678 2398 24690 2430
rect 23706 1884 23712 2380
rect 24684 1894 24690 2398
rect 23706 1854 23724 1884
rect 22936 1804 23424 1810
rect 22936 1770 22948 1804
rect 23412 1770 23424 1804
rect 22936 1764 23424 1770
rect 22632 1658 22638 1718
rect 22698 1658 22704 1718
rect 22636 1552 22642 1612
rect 22702 1552 22708 1612
rect 22126 1446 22132 1506
rect 22192 1446 22198 1506
rect 21622 1336 21628 1396
rect 21688 1336 21694 1396
rect 20900 1282 21388 1288
rect 20900 1248 20912 1282
rect 21376 1248 21388 1282
rect 20900 1242 21388 1248
rect 20604 1172 20618 1198
rect 18864 572 19352 578
rect 18864 538 18876 572
rect 19340 538 19352 572
rect 18864 532 19352 538
rect 18560 414 18566 474
rect 18626 414 18632 474
rect 19082 372 19142 532
rect 18056 366 18118 372
rect 18056 360 18058 366
rect 19082 366 19144 372
rect 19082 360 19084 366
rect 18058 300 18118 306
rect 19084 300 19144 306
rect 19590 110 19650 622
rect 20612 622 20618 1172
rect 20652 1172 20664 1198
rect 21628 1198 21688 1336
rect 22132 1288 22192 1446
rect 21918 1282 22406 1288
rect 21918 1248 21930 1282
rect 22394 1248 22406 1282
rect 21918 1242 22406 1248
rect 20652 622 20658 1172
rect 20612 610 20658 622
rect 21628 622 21636 1198
rect 21670 622 21688 1198
rect 22642 1198 22702 1552
rect 23150 1506 23210 1764
rect 23144 1446 23150 1506
rect 23210 1446 23216 1506
rect 23150 1288 23210 1446
rect 23664 1396 23724 1854
rect 24676 1854 24690 1894
rect 24724 2398 24738 2430
rect 24724 1894 24730 2398
rect 25692 2386 25708 2430
rect 24724 1854 24736 1894
rect 25702 1878 25708 2386
rect 23954 1804 24442 1810
rect 23954 1770 23966 1804
rect 24430 1770 24442 1804
rect 23954 1764 24442 1770
rect 24176 1506 24236 1764
rect 24676 1718 24736 1854
rect 25700 1854 25708 1878
rect 25742 2386 25752 2430
rect 26720 2430 26766 2442
rect 25742 1878 25748 2386
rect 26720 1900 26726 2430
rect 25742 1854 25760 1878
rect 24972 1804 25460 1810
rect 24972 1770 24984 1804
rect 25448 1770 25460 1804
rect 24972 1764 25460 1770
rect 24670 1658 24676 1718
rect 24736 1658 24742 1718
rect 24672 1552 24678 1612
rect 24738 1552 24744 1612
rect 24170 1446 24176 1506
rect 24236 1446 24242 1506
rect 23658 1336 23664 1396
rect 23724 1336 23730 1396
rect 22936 1282 23424 1288
rect 22936 1248 22948 1282
rect 23412 1248 23424 1282
rect 22936 1242 23424 1248
rect 22642 1172 22654 1198
rect 19882 572 20370 578
rect 19882 538 19894 572
rect 20358 538 20370 572
rect 19882 532 20370 538
rect 20900 572 21388 578
rect 20900 538 20912 572
rect 21376 538 21388 572
rect 20900 532 21388 538
rect 20096 366 20156 532
rect 20096 300 20156 306
rect 21132 366 21192 532
rect 21132 300 21192 306
rect 21628 110 21688 622
rect 22648 622 22654 1172
rect 22688 1172 22702 1198
rect 23664 1198 23724 1336
rect 24176 1288 24236 1446
rect 23954 1282 24442 1288
rect 23954 1248 23966 1282
rect 24430 1248 24442 1282
rect 23954 1242 24442 1248
rect 22688 622 22694 1172
rect 22648 610 22694 622
rect 23664 622 23672 1198
rect 23706 622 23724 1198
rect 24678 1198 24738 1552
rect 25178 1506 25238 1764
rect 25172 1446 25178 1506
rect 25238 1446 25244 1506
rect 25178 1288 25238 1446
rect 25700 1396 25760 1854
rect 26712 1854 26726 1900
rect 26760 1900 26766 2430
rect 27728 2430 27788 2658
rect 27874 2614 27934 2878
rect 27868 2554 27874 2614
rect 27934 2554 27940 2614
rect 28238 2520 28298 2998
rect 28750 2718 28810 3088
rect 29768 3088 29780 3132
rect 29814 3132 29820 3664
rect 30782 3664 30842 3802
rect 31308 3754 31368 3804
rect 32322 3754 32382 3932
rect 32816 3804 32822 3864
rect 32882 3804 32888 3864
rect 31080 3748 31568 3754
rect 31080 3714 31092 3748
rect 31556 3714 31568 3748
rect 31080 3708 31568 3714
rect 32098 3748 32586 3754
rect 32098 3714 32110 3748
rect 32574 3714 32586 3748
rect 32098 3708 32586 3714
rect 30782 3618 30798 3664
rect 30792 3136 30798 3618
rect 29814 3088 29828 3132
rect 29044 3038 29532 3044
rect 29044 3004 29056 3038
rect 29520 3004 29532 3038
rect 29044 2998 29532 3004
rect 28744 2658 28750 2718
rect 28810 2658 28816 2718
rect 29258 2520 29318 2998
rect 29768 2946 29828 3088
rect 30784 3088 30798 3136
rect 30832 3618 30842 3664
rect 31810 3664 31856 3676
rect 32822 3664 32882 3804
rect 33116 3748 33604 3754
rect 33116 3714 33128 3748
rect 33592 3714 33604 3748
rect 33116 3708 33604 3714
rect 30832 3136 30838 3618
rect 30832 3088 30844 3136
rect 31810 3132 31816 3664
rect 30062 3038 30550 3044
rect 30062 3004 30074 3038
rect 30538 3004 30550 3038
rect 30062 2998 30550 3004
rect 29762 2886 29768 2946
rect 29828 2886 29834 2946
rect 29764 2658 29770 2718
rect 29830 2658 29836 2718
rect 28026 2514 28514 2520
rect 28026 2480 28038 2514
rect 28502 2480 28514 2514
rect 28026 2474 28514 2480
rect 29044 2514 29532 2520
rect 29044 2480 29056 2514
rect 29520 2480 29532 2514
rect 29044 2474 29532 2480
rect 27728 2386 27744 2430
rect 26760 1854 26772 1900
rect 27738 1880 27744 2386
rect 25990 1804 26478 1810
rect 25990 1770 26002 1804
rect 26466 1770 26478 1804
rect 25990 1764 26478 1770
rect 26198 1506 26258 1764
rect 26540 1658 26546 1718
rect 26606 1658 26612 1718
rect 26192 1446 26198 1506
rect 26258 1446 26264 1506
rect 26546 1466 26606 1658
rect 26712 1612 26772 1854
rect 27732 1854 27744 1880
rect 27778 2386 27788 2430
rect 28756 2430 28802 2442
rect 27778 1880 27784 2386
rect 28756 1894 28762 2430
rect 27778 1854 27792 1880
rect 27008 1804 27496 1810
rect 27008 1770 27020 1804
rect 27484 1770 27496 1804
rect 27008 1764 27496 1770
rect 26706 1552 26712 1612
rect 26772 1552 26778 1612
rect 27218 1506 27278 1764
rect 25694 1336 25700 1396
rect 25760 1336 25766 1396
rect 24972 1282 25460 1288
rect 24972 1248 24984 1282
rect 25448 1248 25460 1282
rect 24972 1242 25460 1248
rect 24678 1162 24690 1198
rect 21918 572 22406 578
rect 21918 538 21930 572
rect 22394 538 22406 572
rect 21918 532 22406 538
rect 22936 572 23424 578
rect 22936 538 22948 572
rect 23412 538 23424 572
rect 22936 532 23424 538
rect 22138 366 22198 532
rect 23152 366 23212 532
rect 23146 306 23152 366
rect 23212 306 23218 366
rect 22138 300 22198 306
rect 23664 110 23724 622
rect 24684 622 24690 1162
rect 24724 1162 24738 1198
rect 25700 1198 25760 1336
rect 26198 1288 26258 1446
rect 26546 1406 26772 1466
rect 27212 1446 27218 1506
rect 27278 1446 27284 1506
rect 25990 1282 26478 1288
rect 25990 1248 26002 1282
rect 26466 1248 26478 1282
rect 25990 1242 26478 1248
rect 24724 622 24730 1162
rect 24684 610 24730 622
rect 25700 622 25708 1198
rect 25742 622 25760 1198
rect 26712 1198 26772 1406
rect 27218 1288 27278 1446
rect 27732 1396 27792 1854
rect 28752 1854 28762 1894
rect 28796 1894 28802 2430
rect 29770 2430 29830 2658
rect 30272 2520 30332 2998
rect 30784 2718 30844 3088
rect 31800 3088 31816 3132
rect 31850 3132 31856 3664
rect 32820 3630 32834 3664
rect 32822 3620 32834 3630
rect 31850 3088 31860 3132
rect 31080 3038 31568 3044
rect 31080 3004 31092 3038
rect 31556 3004 31568 3038
rect 31080 2998 31568 3004
rect 30778 2658 30784 2718
rect 30844 2658 30850 2718
rect 30778 2554 30784 2614
rect 30844 2554 30850 2614
rect 30062 2514 30550 2520
rect 30062 2480 30074 2514
rect 30538 2480 30550 2514
rect 30062 2474 30550 2480
rect 30280 2470 30340 2474
rect 29770 2364 29780 2430
rect 29774 1900 29780 2364
rect 28796 1854 28812 1894
rect 28026 1804 28514 1810
rect 28026 1770 28038 1804
rect 28502 1770 28514 1804
rect 28026 1764 28514 1770
rect 28244 1506 28304 1764
rect 28752 1612 28812 1854
rect 29764 1854 29780 1900
rect 29814 2364 29830 2430
rect 30784 2430 30844 2554
rect 31308 2520 31368 2998
rect 31800 2946 31860 3088
rect 32828 3088 32834 3620
rect 32868 3620 32882 3664
rect 33834 3664 33894 3932
rect 32868 3088 32874 3620
rect 33834 3610 33852 3664
rect 32828 3076 32874 3088
rect 33846 3088 33852 3610
rect 33886 3626 33898 3664
rect 33886 3610 33894 3626
rect 33886 3088 33892 3610
rect 33846 3076 33892 3088
rect 32098 3038 32586 3044
rect 32098 3004 32110 3038
rect 32574 3004 32586 3038
rect 32098 2998 32586 3004
rect 33116 3038 33604 3044
rect 33116 3004 33128 3038
rect 33592 3004 33604 3038
rect 33116 2998 33604 3004
rect 31794 2886 31800 2946
rect 31860 2886 31866 2946
rect 32320 2836 32380 2998
rect 33328 2836 33388 2998
rect 33946 2946 34006 8736
rect 34068 7822 34074 7882
rect 34134 7822 34140 7882
rect 34074 6324 34134 7822
rect 34190 7558 34250 8850
rect 34306 7600 34312 7660
rect 34372 7600 34378 7660
rect 34184 7498 34190 7558
rect 34250 7498 34256 7558
rect 34068 6264 34074 6324
rect 34134 6264 34140 6324
rect 34064 5362 34070 5422
rect 34130 5362 34136 5422
rect 34070 4098 34130 5362
rect 34190 4196 34250 7498
rect 34184 4136 34190 4196
rect 34250 4136 34256 4196
rect 34064 4038 34070 4098
rect 34130 4038 34136 4098
rect 33940 2886 33946 2946
rect 34006 2886 34012 2946
rect 32314 2776 32320 2836
rect 32380 2776 32386 2836
rect 33322 2776 33328 2836
rect 33388 2776 33394 2836
rect 34190 2720 34250 4136
rect 34312 3864 34372 7600
rect 34440 6432 34500 8954
rect 34438 6426 34500 6432
rect 34498 6366 34500 6426
rect 34438 6360 34500 6366
rect 34440 3992 34500 6360
rect 34434 3932 34440 3992
rect 34500 3932 34506 3992
rect 34306 3804 34312 3864
rect 34372 3804 34378 3864
rect 34562 2836 34622 13764
rect 34668 9954 34674 10014
rect 34734 9954 34740 10014
rect 34556 2776 34562 2836
rect 34622 2776 34628 2836
rect 31800 2658 31806 2718
rect 31866 2658 31872 2718
rect 32822 2660 34250 2720
rect 31080 2514 31568 2520
rect 31080 2480 31092 2514
rect 31556 2480 31568 2514
rect 31080 2474 31568 2480
rect 30784 2384 30798 2430
rect 29814 1900 29820 2364
rect 29814 1854 29824 1900
rect 29044 1804 29532 1810
rect 29044 1770 29056 1804
rect 29520 1770 29532 1804
rect 29044 1764 29532 1770
rect 28746 1552 28752 1612
rect 28812 1552 28818 1612
rect 29262 1506 29322 1764
rect 28238 1446 28244 1506
rect 28304 1446 28310 1506
rect 29256 1446 29262 1506
rect 29322 1446 29328 1506
rect 27726 1336 27732 1396
rect 27792 1336 27798 1396
rect 27008 1282 27496 1288
rect 27008 1248 27020 1282
rect 27484 1248 27496 1282
rect 27008 1242 27496 1248
rect 26712 1162 26726 1198
rect 23954 572 24442 578
rect 23954 538 23966 572
rect 24430 538 24442 572
rect 23954 532 24442 538
rect 24972 572 25460 578
rect 24972 538 24984 572
rect 25448 538 25460 572
rect 24972 532 25460 538
rect 24168 366 24228 532
rect 25178 372 25238 532
rect 24168 300 24228 306
rect 25176 366 25238 372
rect 25236 360 25238 366
rect 25176 300 25236 306
rect 25700 110 25760 622
rect 26720 622 26726 1162
rect 26760 1162 26772 1198
rect 27732 1198 27792 1336
rect 28244 1288 28304 1446
rect 29262 1288 29322 1446
rect 29764 1396 29824 1854
rect 30792 1854 30798 2384
rect 30832 2384 30844 2430
rect 31806 2430 31866 2658
rect 32098 2514 32586 2520
rect 32098 2480 32110 2514
rect 32574 2480 32586 2514
rect 32098 2474 32586 2480
rect 30832 1854 30838 2384
rect 31806 2370 31816 2430
rect 31810 1878 31816 2370
rect 30792 1842 30838 1854
rect 31804 1854 31816 1878
rect 31850 2370 31866 2430
rect 32822 2430 32882 2660
rect 33320 2520 33380 2660
rect 33116 2514 33604 2520
rect 33116 2480 33128 2514
rect 33592 2480 33604 2514
rect 33116 2474 33604 2480
rect 31850 1878 31856 2370
rect 31850 1854 31864 1878
rect 30062 1804 30550 1810
rect 30062 1770 30074 1804
rect 30538 1770 30550 1804
rect 30062 1764 30550 1770
rect 31080 1804 31568 1810
rect 31080 1770 31092 1804
rect 31556 1770 31568 1804
rect 31080 1764 31568 1770
rect 30276 1506 30336 1764
rect 30776 1552 30782 1612
rect 30842 1552 30848 1612
rect 30270 1446 30276 1506
rect 30336 1446 30342 1506
rect 29758 1336 29764 1396
rect 29824 1336 29830 1396
rect 28026 1282 28514 1288
rect 28026 1248 28038 1282
rect 28502 1248 28514 1282
rect 28026 1242 28514 1248
rect 29044 1282 29532 1288
rect 29044 1248 29056 1282
rect 29520 1248 29532 1282
rect 29044 1242 29532 1248
rect 26760 622 26766 1162
rect 26720 610 26766 622
rect 27732 622 27744 1198
rect 27778 622 27792 1198
rect 28756 1198 28802 1210
rect 28756 674 28762 1198
rect 27216 578 27276 580
rect 25990 572 26478 578
rect 25990 538 26002 572
rect 26466 538 26478 572
rect 25990 532 26478 538
rect 27008 572 27496 578
rect 27008 538 27020 572
rect 27484 538 27496 572
rect 27008 532 27496 538
rect 26194 372 26254 532
rect 26192 366 26254 372
rect 26252 360 26254 366
rect 27216 366 27276 532
rect 26192 300 26252 306
rect 27216 300 27276 306
rect 27732 110 27792 622
rect 28746 622 28762 674
rect 28796 674 28802 1198
rect 29764 1198 29824 1336
rect 30276 1288 30336 1446
rect 30062 1282 30550 1288
rect 30062 1248 30074 1282
rect 30538 1248 30550 1282
rect 30062 1242 30550 1248
rect 28796 622 28806 674
rect 28026 572 28514 578
rect 28026 538 28038 572
rect 28502 538 28514 572
rect 28026 532 28514 538
rect 28238 366 28298 532
rect 28746 474 28806 622
rect 29764 622 29780 1198
rect 29814 622 29824 1198
rect 30782 1198 30842 1552
rect 31290 1506 31350 1764
rect 31284 1446 31290 1506
rect 31350 1446 31356 1506
rect 31290 1288 31350 1446
rect 31804 1396 31864 1854
rect 32822 1854 32834 2430
rect 32868 1854 32882 2430
rect 33836 2430 33896 2660
rect 33960 2554 33966 2614
rect 34026 2554 34032 2614
rect 33836 2376 33852 2430
rect 32098 1804 32586 1810
rect 32098 1770 32110 1804
rect 32574 1770 32586 1804
rect 32098 1764 32586 1770
rect 32312 1506 32372 1764
rect 32822 1718 32882 1854
rect 33846 1854 33852 2376
rect 33886 2376 33896 2430
rect 33886 1854 33892 2376
rect 33846 1842 33892 1854
rect 33116 1804 33604 1810
rect 33116 1770 33128 1804
rect 33592 1770 33604 1804
rect 33116 1764 33604 1770
rect 32816 1658 32822 1718
rect 32882 1658 32888 1718
rect 32816 1552 32822 1612
rect 32882 1552 32888 1612
rect 32306 1446 32312 1506
rect 32372 1446 32378 1506
rect 31798 1336 31804 1396
rect 31864 1336 31870 1396
rect 31080 1282 31568 1288
rect 31080 1248 31092 1282
rect 31556 1248 31568 1282
rect 31080 1242 31568 1248
rect 30782 1154 30798 1198
rect 29044 572 29532 578
rect 29044 538 29056 572
rect 29520 538 29532 572
rect 29044 532 29532 538
rect 28740 414 28746 474
rect 28806 414 28812 474
rect 29258 372 29318 532
rect 29258 366 29320 372
rect 29258 360 29260 366
rect 28238 300 28298 306
rect 29260 300 29320 306
rect 29764 110 29824 622
rect 30792 622 30798 1154
rect 30832 1154 30842 1198
rect 31804 1198 31864 1336
rect 32312 1288 32372 1446
rect 32822 1396 32882 1552
rect 32822 1336 33900 1396
rect 32098 1282 32586 1288
rect 32098 1248 32110 1282
rect 32574 1248 32586 1282
rect 32098 1242 32586 1248
rect 30832 622 30838 1154
rect 30792 610 30838 622
rect 31804 622 31816 1198
rect 31850 622 31864 1198
rect 32822 1198 32882 1336
rect 33338 1288 33398 1336
rect 33116 1282 33604 1288
rect 33116 1248 33128 1282
rect 33592 1248 33604 1282
rect 33116 1242 33604 1248
rect 32822 1190 32834 1198
rect 30280 578 30340 580
rect 30062 572 30550 578
rect 30062 538 30074 572
rect 30538 538 30550 572
rect 30062 532 30550 538
rect 31080 572 31568 578
rect 31080 538 31092 572
rect 31556 538 31568 572
rect 31080 532 31568 538
rect 30280 372 30340 532
rect 31294 372 31354 532
rect 30278 366 30340 372
rect 30338 360 30340 366
rect 31292 366 31354 372
rect 30278 300 30338 306
rect 31352 360 31354 366
rect 31292 300 31352 306
rect 31804 110 31864 622
rect 32828 622 32834 1190
rect 32868 1190 32882 1198
rect 33840 1198 33900 1336
rect 32868 622 32874 1190
rect 33840 1180 33852 1198
rect 32828 610 32874 622
rect 33846 622 33852 1180
rect 33886 1180 33900 1198
rect 33886 622 33892 1180
rect 33846 610 33892 622
rect 32314 578 32374 580
rect 32098 572 32586 578
rect 32098 538 32110 572
rect 32574 538 32586 572
rect 32098 532 32586 538
rect 33116 572 33604 578
rect 33116 538 33128 572
rect 33592 538 33604 572
rect 33116 532 33604 538
rect 32314 372 32374 532
rect 33966 474 34026 2554
rect 34674 1612 34734 9954
rect 34668 1552 34674 1612
rect 34734 1552 34740 1612
rect 33960 414 33966 474
rect 34026 414 34032 474
rect 32314 366 32376 372
rect 32314 360 32316 366
rect 32316 300 32376 306
rect 35728 210 35734 14470
rect 35834 210 35840 14470
rect 2794 64 2944 110
rect 2990 64 6164 110
rect 6224 64 12616 110
rect 12676 64 34718 110
rect 34778 64 34880 110
rect 2794 -90 2840 64
rect 34840 -90 34880 64
rect 2794 -136 34880 -90
rect -704 -576 -694 -276
rect 35118 -576 35128 -276
rect 35728 -576 35840 210
rect -1416 -582 35840 -576
rect -1416 -682 -1310 -582
rect 35734 -682 35840 -582
rect -1416 -688 35840 -682
<< via1 >>
rect -4458 30228 -4398 30288
rect 11396 30456 11996 30756
rect 35028 30456 35628 30756
rect 14973 30160 31758 30374
rect 18898 28398 18958 28458
rect 19980 28398 20040 28458
rect 20938 28398 20998 28458
rect 19424 28152 19484 28212
rect 21460 28152 21520 28212
rect 17242 27220 17302 27280
rect 18406 27220 18466 27280
rect 17112 27016 17172 27076
rect 15104 24832 15164 24892
rect 18406 27016 18466 27076
rect 24002 28398 24062 28458
rect 25020 28398 25080 28458
rect 23498 28154 23558 28214
rect 20442 27116 20502 27176
rect 18892 25866 18952 25926
rect 26044 28398 26104 28458
rect 27056 28398 27116 28458
rect 25528 28154 25588 28214
rect 22478 27116 22538 27176
rect 27570 28156 27630 28216
rect 24516 27220 24576 27280
rect 24512 27016 24572 27076
rect 20948 26082 21008 26142
rect 21458 26082 21518 26142
rect 20440 25980 20504 26044
rect 19930 25866 19990 25926
rect 20942 25866 21002 25926
rect 17242 24546 17302 24606
rect 17598 22138 17658 22198
rect 17472 21528 17532 21588
rect 14588 20574 14648 20634
rect 14696 20462 14756 20522
rect 12926 19540 12986 19600
rect 15610 20574 15670 20634
rect 15480 20462 15540 20522
rect 14086 19430 14146 19490
rect 16120 19540 16180 19600
rect 12800 18452 12860 18512
rect 14602 18506 14662 18566
rect 14708 18406 14768 18466
rect 17272 19430 17332 19490
rect 15612 18506 15672 18566
rect 17464 19302 17524 19362
rect 15494 18406 15554 18466
rect 12314 17396 12374 17456
rect 12454 17220 12514 17280
rect 13354 17046 13414 17106
rect 17714 21528 17774 21588
rect 18400 24692 18464 24756
rect 18224 24546 18284 24606
rect 22316 25980 22380 26044
rect 28580 28156 28640 28216
rect 30114 28398 30174 28458
rect 31126 28398 31186 28458
rect 29602 28156 29662 28216
rect 26550 27220 26610 27280
rect 26548 27016 26608 27076
rect 27050 27016 27110 27076
rect 23492 26082 23552 26142
rect 21952 25874 22012 25934
rect 22976 25874 23036 25934
rect 19422 24944 19482 25004
rect 20438 24830 20502 24894
rect 24004 25874 24064 25934
rect 32144 28398 32204 28458
rect 31638 28156 31698 28216
rect 28584 27116 28644 27176
rect 28070 27016 28130 27076
rect 25530 26080 25590 26140
rect 21458 24944 21518 25004
rect 21980 24944 22040 25004
rect 22478 24944 22538 25004
rect 29096 27016 29156 27076
rect 30618 27116 30678 27176
rect 29602 27012 29662 27072
rect 30116 27012 30176 27072
rect 30620 27012 30680 27072
rect 31126 27012 31186 27072
rect 31646 27012 31706 27072
rect 26550 25982 26610 26042
rect 32658 27220 32718 27280
rect 33908 27220 33968 27280
rect 27566 26080 27626 26140
rect 28066 26080 28126 26140
rect 28580 26080 28640 26140
rect 29104 26080 29164 26140
rect 29602 26080 29662 26140
rect 30104 26080 30164 26140
rect 22952 24940 23012 25000
rect 18340 24440 18400 24500
rect 18902 24440 18962 24500
rect 19944 24440 20004 24500
rect 20944 24440 21004 24500
rect 23492 25002 23552 25004
rect 23460 24944 23552 25002
rect 23952 24944 24012 25004
rect 23460 24942 23520 24944
rect 24510 24688 24574 24752
rect 24996 24946 25056 25006
rect 24106 24440 24166 24500
rect 25528 24944 25588 25004
rect 30618 26078 30678 26138
rect 31126 26078 31186 26138
rect 31636 26078 31696 26138
rect 30108 25866 30168 25926
rect 31120 25866 31180 25926
rect 27040 24946 27100 25006
rect 26546 24546 26610 24610
rect 25116 24440 25176 24500
rect 26058 24440 26118 24500
rect 27566 25000 27626 25002
rect 27534 24942 27626 25000
rect 27534 24940 27594 24942
rect 28062 24936 28122 24996
rect 28550 24998 28610 25000
rect 28550 24940 28644 24998
rect 28584 24938 28644 24940
rect 32658 25982 32718 26042
rect 32122 25866 32182 25926
rect 29062 24936 29122 24996
rect 29602 24940 29662 25000
rect 31636 24940 31696 25000
rect 30618 24830 30682 24894
rect 33904 24692 33968 24756
rect 32652 24546 32712 24606
rect 18454 24238 18514 24298
rect 21632 24238 21692 24298
rect 19598 23302 19658 23362
rect 20102 23194 20162 23254
rect 21632 23302 21692 23362
rect 21124 23194 21184 23254
rect 22142 23194 22202 23254
rect 19594 22270 19654 22330
rect 20100 22136 20160 22196
rect 25700 24238 25760 24298
rect 23674 23302 23734 23362
rect 23166 23194 23226 23254
rect 24180 23194 24240 23254
rect 21114 22132 21174 22192
rect 22146 22140 22206 22200
rect 25700 23302 25760 23362
rect 25198 23194 25258 23254
rect 26208 23194 26268 23254
rect 23674 22270 23734 22330
rect 23144 22140 23204 22200
rect 24188 22140 24248 22200
rect 29776 24238 29836 24298
rect 27742 23302 27802 23362
rect 27230 23194 27290 23254
rect 28244 23194 28304 23254
rect 25192 22136 25252 22196
rect 26208 22136 26268 22196
rect 24992 21928 25052 21988
rect 18224 21610 18284 21670
rect 19390 21610 19450 21670
rect 17956 20564 18016 20624
rect 17714 19406 17774 19466
rect 17710 19192 17770 19252
rect 17598 18150 17658 18210
rect 12194 16896 12254 16956
rect -7916 16376 -7856 16436
rect -4458 16376 -4398 16436
rect -11016 16268 -10956 16328
rect -11664 15502 -11604 15562
rect -11922 15353 -11862 15413
rect -11146 15502 -11086 15562
rect -11406 15353 -11346 15413
rect -8416 16268 -8356 16328
rect -10343 15484 -10283 15490
rect -10343 15436 -10337 15484
rect -10337 15436 -10289 15484
rect -10289 15436 -10283 15484
rect -10343 15430 -10283 15436
rect -10025 15452 -9965 15512
rect -9064 15502 -9004 15562
rect -10888 15353 -10828 15413
rect -9322 15353 -9262 15413
rect -11018 14805 -10958 14865
rect -8546 15502 -8486 15562
rect -8806 15353 -8746 15413
rect 18092 20466 18152 20526
rect 17956 16892 18016 16952
rect 21426 21610 21486 21670
rect 21934 21606 21998 21670
rect 20408 20662 20468 20722
rect 32972 24238 33032 24298
rect 29778 23302 29838 23362
rect 29276 23194 29336 23254
rect 30286 23194 30346 23254
rect 27742 22270 27802 22330
rect 27212 22136 27272 22196
rect 28244 22140 28304 22200
rect 26728 21928 26788 21988
rect 26008 21728 26072 21792
rect 31814 23302 31874 23362
rect 31308 23194 31368 23254
rect 29260 22136 29320 22196
rect 30288 22136 30348 22196
rect 31810 22270 31870 22330
rect 31308 22136 31368 22196
rect 33766 22138 33826 22198
rect 32626 21912 32686 21972
rect 30072 21728 30136 21792
rect 31096 21728 31160 21792
rect 32108 21728 32172 21792
rect 26010 21606 26074 21670
rect 22444 20662 22504 20722
rect 22786 20664 22846 20724
rect 20408 20466 20468 20526
rect 21428 20468 21488 20528
rect 19394 20356 19454 20416
rect 21428 20356 21488 20416
rect 18376 19192 18436 19252
rect 25500 20664 25560 20724
rect 29572 21610 29632 21670
rect 31606 21610 31666 21670
rect 26518 20468 26578 20528
rect 24484 20354 24544 20414
rect 26518 20354 26578 20414
rect 20410 19302 20470 19362
rect 20410 19098 20470 19158
rect 22446 19302 22506 19362
rect 22444 19200 22504 19260
rect 22444 19098 22504 19158
rect 19392 18150 19452 18210
rect 18224 17942 18284 18002
rect 20406 17840 20466 17900
rect 24480 19406 24540 19466
rect 21428 18150 21488 18210
rect 21428 18042 21488 18102
rect 25500 19406 25560 19466
rect 25500 19100 25560 19160
rect 29574 20354 29634 20414
rect 26518 19100 26578 19160
rect 30588 20662 30648 20722
rect 31608 20354 31668 20414
rect 32624 20662 32684 20722
rect 27536 19406 27596 19466
rect 27534 19100 27594 19160
rect 22446 18158 22506 18218
rect 24248 18158 24308 18218
rect 22440 17840 22500 17900
rect 22644 17828 22704 17888
rect 19388 16892 19448 16952
rect 24482 18152 24542 18212
rect 29570 19302 29630 19362
rect 30438 19420 30498 19480
rect 30586 19310 30646 19370
rect 30438 19100 30498 19160
rect 30590 19102 30650 19162
rect 26518 18152 26578 18212
rect 26516 18042 26576 18102
rect 21424 16892 21484 16952
rect 18092 16762 18152 16822
rect 13248 16634 13308 16694
rect 13128 16516 13188 16576
rect 26006 17828 26066 17888
rect 31606 19200 31666 19260
rect 34202 22270 34262 22330
rect 33908 21910 33968 21970
rect 34050 21610 34110 21670
rect 33890 20468 33950 20528
rect 32626 19310 32686 19370
rect 33766 19310 33826 19370
rect 32624 19102 32684 19162
rect 27022 17828 27082 17888
rect 29572 18154 29632 18214
rect 30082 17828 30142 17888
rect 30594 17840 30654 17900
rect 31608 18154 31668 18214
rect 33890 19102 33950 19162
rect 33766 18042 33826 18102
rect 32628 17840 32688 17900
rect 29576 16892 29636 16952
rect 31612 16892 31672 16952
rect 22446 16622 22506 16682
rect 34202 20354 34262 20414
rect 34050 16622 34110 16682
rect 12682 16398 12742 16458
rect -2718 15870 8046 16162
rect -7743 15484 -7683 15490
rect -7743 15436 -7737 15484
rect -7737 15436 -7689 15484
rect -7689 15436 -7683 15484
rect -7743 15430 -7683 15436
rect -7425 15452 -7365 15512
rect -8288 15353 -8228 15413
rect -8418 14805 -8358 14865
rect 12800 15122 12860 15182
rect 13128 15132 13188 15192
rect 12194 14986 12254 15046
rect 12314 14988 12374 15048
rect 12454 15006 12514 15066
rect 12682 15022 12742 15082
rect 12062 14858 12122 14918
rect 9350 14260 9410 14320
rect 10876 14126 10936 14186
rect 12062 7658 12122 7718
rect 7514 6732 7574 6792
rect 1404 6586 1464 6646
rect 5484 6586 5544 6646
rect 250 6458 310 6518
rect 2928 6458 2988 6518
rect 3960 6458 4020 6518
rect 1908 5496 1968 5556
rect 1408 5392 1468 5452
rect 2932 5496 2992 5556
rect 2426 5288 2486 5348
rect 250 4226 310 4286
rect 7020 6458 7080 6518
rect 3964 5496 4024 5556
rect 3444 5392 3504 5452
rect 9544 6586 9604 6646
rect 11728 6586 11788 6646
rect 8016 6458 8076 6518
rect 4964 5496 5024 5556
rect 5984 5496 6044 5556
rect 5480 5392 5540 5452
rect 4462 5288 4522 5348
rect 1900 4226 1960 4286
rect 3438 4346 3498 4406
rect 7004 5496 7064 5556
rect 6494 5288 6554 5348
rect 4970 4226 5030 4286
rect 8014 5496 8074 5556
rect 7514 5392 7574 5452
rect 9028 5496 9088 5556
rect 10046 5496 10106 5556
rect 9550 5392 9610 5452
rect 8528 5288 8588 5348
rect 5978 4226 6038 4286
rect 2426 3282 2486 3342
rect 1412 3174 1472 3234
rect 1906 3062 1966 3122
rect 3448 3174 3508 3234
rect 2930 3062 2990 3122
rect 7514 4346 7574 4406
rect 4462 3282 4522 3342
rect 3962 3062 4022 3122
rect 10572 5288 10632 5348
rect 9040 4226 9100 4286
rect 11848 5496 11908 5556
rect 11728 4346 11788 4406
rect 10066 4226 10126 4286
rect 6494 3282 6554 3342
rect 5484 3174 5544 3234
rect 4962 3062 5022 3122
rect 5982 3062 6042 3122
rect 7518 3174 7578 3234
rect 7002 3062 7062 3122
rect 250 2100 310 2160
rect 2920 2100 2980 2160
rect 3952 2100 4012 2160
rect 8012 3062 8072 3122
rect 8528 3282 8588 3342
rect 10572 3282 10632 3342
rect 9554 3174 9614 3234
rect 9026 3062 9086 3122
rect 10044 3062 10104 3122
rect 7012 2100 7072 2160
rect 8008 2100 8068 2160
rect 11848 3062 11908 3122
rect 1406 1970 1466 2030
rect 5486 1970 5546 2030
rect 9546 1970 9606 2030
rect 11728 1970 11788 2030
rect 2884 604 2944 664
rect 4922 604 4982 664
rect 6958 604 7018 664
rect 3902 492 3962 552
rect 8994 604 9054 664
rect 7976 492 8036 552
rect 12194 6586 12254 6646
rect 12314 6458 12374 6518
rect 12572 14868 12632 14928
rect 12682 14126 12742 14186
rect 13248 15124 13308 15184
rect 13128 14260 13188 14320
rect 12924 12902 12984 12962
rect 12798 11200 12858 11260
rect 12572 8740 12632 8800
rect 12454 5496 12514 5556
rect 13136 12566 13196 12626
rect 13032 11306 13092 11366
rect 12924 10206 12984 10266
rect 13354 14988 13414 15048
rect 24166 14638 24226 14698
rect 29270 14638 29330 14698
rect 33330 14632 33390 14692
rect 14498 12902 14558 12962
rect 15512 12686 15572 12746
rect 17552 12686 17612 12746
rect 19592 12686 19652 12746
rect 21622 12686 21682 12746
rect 23662 12686 23722 12746
rect 25694 12686 25754 12746
rect 27734 12686 27794 12746
rect 29770 12686 29830 12746
rect 31804 12686 31864 12746
rect 13480 12566 13540 12626
rect 15004 12560 15064 12620
rect 13354 12444 13414 12504
rect 16018 12560 16078 12620
rect 17040 12560 17100 12620
rect 18054 12560 18114 12620
rect 19080 12560 19140 12620
rect 18568 12444 18628 12504
rect 20092 12560 20152 12620
rect 21128 12560 21188 12620
rect 22134 12560 22194 12620
rect 23148 12560 23208 12620
rect 15516 11522 15576 11582
rect 15008 11412 15068 11472
rect 14498 11306 14558 11366
rect 13484 11200 13544 11260
rect 13982 11200 14042 11260
rect 14494 11200 14554 11260
rect 16030 11412 16090 11472
rect 17556 11522 17616 11582
rect 17044 11412 17104 11472
rect 16538 11306 16598 11366
rect 19588 11522 19648 11582
rect 18058 11412 18118 11472
rect 19076 11412 19136 11472
rect 18568 11306 18628 11366
rect 13354 10310 13414 10370
rect 13478 10206 13538 10266
rect 14998 10206 15058 10266
rect 15510 10206 15570 10266
rect 13248 10084 13308 10144
rect 13136 9970 13196 10030
rect 13984 9970 14044 10030
rect 15516 9972 15576 10032
rect 20102 11412 20162 11472
rect 24164 12560 24224 12620
rect 25172 12560 25232 12620
rect 26188 12560 26248 12620
rect 27212 12560 27272 12620
rect 28234 12560 28294 12620
rect 29256 12560 29316 12620
rect 28756 12444 28816 12504
rect 21620 11522 21680 11582
rect 20608 11306 20668 11366
rect 21122 11412 21182 11472
rect 20774 11200 20834 11260
rect 16532 10310 16592 10370
rect 16534 10206 16594 10266
rect 22142 11412 22202 11472
rect 23656 11522 23716 11582
rect 23144 11412 23204 11472
rect 22642 11306 22702 11366
rect 22642 11200 22702 11260
rect 24170 11412 24230 11472
rect 30274 12560 30334 12620
rect 31288 12560 31348 12620
rect 32312 12560 32372 12620
rect 32828 12444 32888 12504
rect 33960 12444 34020 12504
rect 25692 11522 25752 11582
rect 25188 11412 25248 11472
rect 24678 11306 24738 11366
rect 24680 11200 24740 11260
rect 26196 11412 26256 11472
rect 27730 11522 27790 11582
rect 27208 11412 27268 11472
rect 26714 11306 26774 11366
rect 26560 11200 26620 11260
rect 17546 10206 17606 10266
rect 17552 9972 17612 10032
rect 18566 10206 18626 10266
rect 13360 9042 13420 9102
rect 14498 9042 14558 9102
rect 13248 8842 13308 8902
rect 13142 8740 13202 8800
rect 13032 5288 13092 5348
rect 13248 7606 13308 7666
rect 12800 5138 12860 5198
rect 13142 5250 13202 5310
rect 14496 8842 14556 8902
rect 15514 8962 15574 9022
rect 19588 10310 19648 10370
rect 29768 11522 29828 11582
rect 28240 11412 28300 11472
rect 29254 11412 29314 11472
rect 28754 11306 28814 11366
rect 25694 10310 25754 10370
rect 21624 10206 21684 10266
rect 23662 10206 23722 10266
rect 20608 10084 20668 10144
rect 22642 10084 22702 10144
rect 24672 10084 24732 10144
rect 16532 9066 16592 9126
rect 16028 8848 16088 8908
rect 17554 8962 17614 9022
rect 17032 8848 17092 8908
rect 14496 7810 14556 7870
rect 15002 7708 15062 7768
rect 18568 9066 18628 9126
rect 18044 8848 18104 8908
rect 19586 8962 19646 9022
rect 19064 8848 19124 8908
rect 19586 8850 19646 8910
rect 21620 8962 21680 9022
rect 20604 8740 20664 8800
rect 16534 7810 16594 7870
rect 16532 7606 16592 7666
rect 21622 8850 21682 8910
rect 22638 8740 22698 8800
rect 26712 10206 26772 10266
rect 30272 11412 30332 11472
rect 31804 11522 31864 11582
rect 31296 11412 31356 11472
rect 30784 11306 30844 11366
rect 30784 11202 30844 11262
rect 27730 10206 27790 10266
rect 28750 10206 28810 10266
rect 23660 8962 23720 9022
rect 23658 8850 23718 8910
rect 25694 8962 25754 9022
rect 25890 8958 25950 9018
rect 24678 8740 24738 8800
rect 25694 8850 25754 8910
rect 32316 11412 32376 11472
rect 32824 11306 32884 11366
rect 33960 11202 34020 11262
rect 30788 10310 30848 10370
rect 29766 10206 29826 10266
rect 31802 10206 31862 10266
rect 26712 9066 26772 9126
rect 25890 8740 25950 8800
rect 26184 8742 26244 8802
rect 18570 7810 18630 7870
rect 15516 7506 15576 7566
rect 17040 7600 17100 7660
rect 18062 7600 18122 7660
rect 17550 7506 17610 7566
rect 20602 7810 20662 7870
rect 20094 7708 20154 7768
rect 19076 7600 19136 7660
rect 20094 7600 20154 7660
rect 19586 7506 19646 7566
rect 14998 6582 15058 6642
rect 15908 6582 15968 6642
rect 14998 6366 15058 6426
rect 13362 6262 13422 6322
rect 16910 6582 16970 6642
rect 16036 6366 16096 6426
rect 18062 6582 18122 6642
rect 17550 6480 17610 6540
rect 17050 6366 17110 6426
rect 14996 5354 15056 5414
rect 14498 5250 14558 5310
rect 14494 5040 14554 5100
rect 16004 5354 16064 5414
rect 15514 5138 15574 5198
rect 21114 7600 21174 7660
rect 27728 8850 27788 8910
rect 27212 8742 27272 8802
rect 27730 8736 27790 8796
rect 28748 9066 28808 9126
rect 29766 8850 29826 8910
rect 30782 8958 30842 9018
rect 31286 8954 31346 9014
rect 33946 9972 34006 10032
rect 31806 8850 31866 8910
rect 29766 8736 29826 8796
rect 25184 7822 25244 7882
rect 24678 7694 24738 7754
rect 26714 7496 26774 7556
rect 19072 6582 19132 6642
rect 20078 6582 20138 6642
rect 21122 6582 21182 6642
rect 21622 6588 21682 6648
rect 20076 6366 20136 6426
rect 21116 6366 21176 6426
rect 20600 6262 20660 6322
rect 17018 5354 17078 5414
rect 18056 5354 18116 5414
rect 17552 5138 17612 5198
rect 16532 5040 16592 5100
rect 22130 6366 22190 6426
rect 23658 6588 23718 6648
rect 23138 6366 23198 6426
rect 24182 6366 24242 6426
rect 22642 6262 22702 6322
rect 31804 8736 31864 8796
rect 28226 7600 28286 7660
rect 25694 6588 25754 6648
rect 25172 6366 25232 6426
rect 26190 6366 26250 6426
rect 24680 6262 24740 6322
rect 32822 9066 32882 9126
rect 33840 9084 33900 9144
rect 34074 9954 34134 10014
rect 34440 8954 34500 9014
rect 34190 8850 34250 8910
rect 30278 7822 30338 7882
rect 30416 7826 30476 7886
rect 33946 8736 34006 8796
rect 31298 7826 31358 7886
rect 32304 7826 32364 7886
rect 29256 7600 29316 7660
rect 30416 7600 30476 7660
rect 30784 7600 30844 7660
rect 30784 7496 30844 7556
rect 32822 7822 32882 7882
rect 32822 7694 32882 7754
rect 31800 7498 31860 7558
rect 27732 6588 27792 6648
rect 27724 6480 27784 6540
rect 27224 6366 27284 6426
rect 26714 6262 26774 6322
rect 27226 6258 27286 6318
rect 28248 6258 28308 6318
rect 28748 6264 28808 6324
rect 19074 5354 19134 5414
rect 19590 5360 19650 5420
rect 21626 5360 21686 5420
rect 23658 5360 23718 5420
rect 25692 5360 25752 5420
rect 18572 5040 18632 5100
rect 13360 4018 13420 4078
rect 14500 3802 14560 3862
rect 15514 4116 15574 4176
rect 15518 3922 15578 3982
rect 16532 4018 16592 4078
rect 22642 5250 22702 5310
rect 24678 5250 24738 5310
rect 21624 5138 21684 5198
rect 20608 5040 20668 5100
rect 17550 4116 17610 4176
rect 18056 4018 18116 4078
rect 17554 3922 17614 3982
rect 19588 4116 19648 4176
rect 19078 4018 19138 4078
rect 18568 3802 18628 3862
rect 13248 2886 13308 2946
rect 13142 2760 13202 2820
rect 20100 4018 20160 4078
rect 19582 3922 19642 3982
rect 29768 6588 29828 6648
rect 29764 6480 29824 6540
rect 30256 6366 30316 6426
rect 31806 6588 31866 6648
rect 31802 6480 31862 6540
rect 31294 6366 31354 6426
rect 30782 6264 30842 6324
rect 26714 5362 26774 5422
rect 27068 5362 27128 5422
rect 26710 5250 26770 5310
rect 26220 5152 26280 5212
rect 21450 4136 21510 4196
rect 21620 4136 21680 4196
rect 21104 4018 21164 4078
rect 20602 3802 20662 3862
rect 16532 2760 16592 2820
rect 17052 2772 17112 2832
rect 15514 2658 15574 2718
rect 17550 2658 17610 2718
rect 16532 2554 16592 2614
rect 13360 1656 13420 1716
rect 13032 1552 13092 1612
rect 14496 1552 14556 1612
rect 15004 1446 15064 1506
rect 11982 492 12042 552
rect 21450 3922 21510 3982
rect 21626 3928 21686 3988
rect 27258 5152 27318 5212
rect 28234 5152 28294 5212
rect 27068 5044 27128 5104
rect 32320 6366 32380 6426
rect 32824 6264 32884 6324
rect 30786 5362 30846 5422
rect 29250 5152 29310 5212
rect 31276 5152 31336 5212
rect 28748 5040 28808 5100
rect 30784 5040 30844 5100
rect 23662 4136 23722 4196
rect 25694 4136 25754 4196
rect 27734 4136 27794 4196
rect 26712 4038 26772 4098
rect 23654 3928 23714 3988
rect 18570 2658 18630 2718
rect 19586 2658 19646 2718
rect 16530 1656 16590 1716
rect 16536 1552 16596 1612
rect 16024 1446 16084 1506
rect 15516 1336 15576 1396
rect 17048 1446 17108 1506
rect 20606 2658 20666 2718
rect 25698 3928 25758 3988
rect 27726 3928 27786 3988
rect 28752 3802 28812 3862
rect 32306 5152 32366 5212
rect 32820 5040 32880 5100
rect 29764 3928 29824 3988
rect 32818 4038 32878 4098
rect 31804 3928 31864 3988
rect 32322 3932 32382 3992
rect 33834 3932 33894 3992
rect 30782 3802 30842 3862
rect 31308 3804 31368 3864
rect 22636 2886 22696 2946
rect 24678 2886 24738 2946
rect 26714 2886 26774 2946
rect 22132 2772 22192 2832
rect 27220 2776 27280 2836
rect 21624 2658 21684 2718
rect 23654 2658 23714 2718
rect 25692 2658 25752 2718
rect 27728 2658 27788 2718
rect 21468 2554 21528 2614
rect 18566 1552 18626 1612
rect 18066 1446 18126 1506
rect 19080 1446 19140 1506
rect 17552 1336 17612 1396
rect 13360 414 13420 474
rect 14496 414 14556 474
rect 15008 306 15068 366
rect 20760 1658 20820 1718
rect 20606 1552 20666 1612
rect 20112 1446 20172 1506
rect 19590 1336 19650 1396
rect 16022 306 16082 366
rect 17044 306 17104 366
rect 21124 1446 21184 1506
rect 22638 1658 22698 1718
rect 22642 1552 22702 1612
rect 22132 1446 22192 1506
rect 21628 1336 21688 1396
rect 18566 414 18626 474
rect 18058 306 18118 366
rect 19084 306 19144 366
rect 23150 1446 23210 1506
rect 24676 1658 24736 1718
rect 24678 1552 24738 1612
rect 24176 1446 24236 1506
rect 23664 1336 23724 1396
rect 20096 306 20156 366
rect 21132 306 21192 366
rect 25178 1446 25238 1506
rect 27874 2554 27934 2614
rect 32822 3804 32882 3864
rect 28750 2658 28810 2718
rect 29768 2886 29828 2946
rect 29770 2658 29830 2718
rect 26546 1658 26606 1718
rect 26198 1446 26258 1506
rect 26712 1552 26772 1612
rect 25700 1336 25760 1396
rect 22138 306 22198 366
rect 23152 306 23212 366
rect 27218 1446 27278 1506
rect 30784 2658 30844 2718
rect 30784 2554 30844 2614
rect 31800 2886 31860 2946
rect 34074 7822 34134 7882
rect 34312 7600 34372 7660
rect 34190 7498 34250 7558
rect 34074 6264 34134 6324
rect 34070 5362 34130 5422
rect 34190 4136 34250 4196
rect 34070 4038 34130 4098
rect 33946 2886 34006 2946
rect 32320 2776 32380 2836
rect 33328 2776 33388 2836
rect 34438 6366 34498 6426
rect 34440 3932 34500 3992
rect 34312 3804 34372 3864
rect 34674 9954 34734 10014
rect 34562 2776 34622 2836
rect 31806 2658 31866 2718
rect 28752 1552 28812 1612
rect 28244 1446 28304 1506
rect 29262 1446 29322 1506
rect 27732 1336 27792 1396
rect 24168 306 24228 366
rect 25176 306 25236 366
rect 30782 1552 30842 1612
rect 30276 1446 30336 1506
rect 29764 1336 29824 1396
rect 26192 306 26252 366
rect 27216 306 27276 366
rect 31290 1446 31350 1506
rect 33966 2554 34026 2614
rect 32822 1658 32882 1718
rect 32822 1552 32882 1612
rect 32312 1446 32372 1506
rect 31804 1336 31864 1396
rect 28746 414 28806 474
rect 28238 306 28298 366
rect 29260 306 29320 366
rect 30278 306 30338 366
rect 31292 306 31352 366
rect 34674 1552 34734 1612
rect 33966 414 34026 474
rect 32316 306 32376 366
rect 2840 -90 34840 64
rect -1304 -576 -704 -276
rect 35128 -576 35728 -276
<< metal2 >>
rect 11396 30756 11996 30766
rect 11396 30446 11996 30456
rect 35028 30756 35628 30766
rect 35028 30446 35628 30456
rect 14910 30374 31790 30406
rect -4458 30288 -4398 30297
rect -4464 30228 -4458 30288
rect -4398 30228 -4392 30288
rect -4458 30219 -4398 30228
rect 14910 30160 14973 30374
rect 31758 30160 31790 30374
rect 14910 30140 31790 30160
rect 14910 30138 19264 30140
rect 18898 28458 18958 28464
rect 19980 28458 20040 28464
rect 20938 28458 20998 28464
rect 24002 28458 24062 28464
rect 25020 28458 25080 28464
rect 26044 28458 26104 28464
rect 27056 28458 27116 28464
rect 30114 28458 30174 28464
rect 31126 28458 31186 28464
rect 32144 28458 32204 28464
rect 18958 28398 19980 28458
rect 20040 28398 20938 28458
rect 20998 28398 24002 28458
rect 24062 28398 25020 28458
rect 25080 28398 26044 28458
rect 26104 28398 27056 28458
rect 27116 28398 30114 28458
rect 30174 28398 31126 28458
rect 31186 28398 32144 28458
rect 18898 28392 18958 28398
rect 19980 28392 20040 28398
rect 20938 28392 20998 28398
rect 24002 28392 24062 28398
rect 25020 28392 25080 28398
rect 26044 28392 26104 28398
rect 27056 28392 27116 28398
rect 30114 28392 30174 28398
rect 31126 28392 31186 28398
rect 32144 28392 32204 28398
rect 19424 28212 19484 28218
rect 21460 28212 21520 28218
rect 23498 28214 23558 28220
rect 25528 28214 25588 28220
rect 27570 28216 27630 28222
rect 28580 28216 28640 28222
rect 29602 28216 29662 28222
rect 31638 28216 31698 28222
rect 19484 28152 21460 28212
rect 21520 28154 23498 28212
rect 23558 28154 25528 28214
rect 25588 28156 27570 28214
rect 27630 28156 28580 28216
rect 28640 28156 29602 28216
rect 29662 28156 31638 28216
rect 25588 28154 27768 28156
rect 21520 28152 23680 28154
rect 19424 28146 19484 28152
rect 21460 28146 21520 28152
rect 23498 28148 23558 28152
rect 25528 28148 25588 28154
rect 27570 28150 27630 28154
rect 28580 28150 28640 28156
rect 29602 28150 29662 28156
rect 31638 28150 31698 28156
rect 17242 27280 17302 27286
rect 18406 27280 18466 27286
rect 24516 27280 24576 27286
rect 17302 27220 18406 27280
rect 18466 27220 24516 27280
rect 17242 27214 17302 27220
rect 18406 27214 18466 27220
rect 24516 27214 24576 27220
rect 26550 27280 26610 27286
rect 32658 27280 32718 27286
rect 33908 27280 33968 27286
rect 26610 27220 32658 27280
rect 32718 27220 33908 27280
rect 26550 27214 26610 27220
rect 32658 27214 32718 27220
rect 33908 27214 33968 27220
rect 20442 27176 20502 27182
rect 22478 27176 22538 27182
rect 28584 27176 28644 27182
rect 30618 27176 30678 27182
rect 20502 27116 22478 27176
rect 22538 27168 22956 27176
rect 23172 27168 28584 27176
rect 22538 27122 28584 27168
rect 22538 27118 24972 27122
rect 22538 27116 23946 27118
rect 24184 27116 24972 27118
rect 25188 27116 28584 27122
rect 28644 27116 30618 27176
rect 20442 27110 20502 27116
rect 22478 27110 22538 27116
rect 28584 27110 28644 27116
rect 30618 27110 30678 27116
rect 17112 27076 17172 27082
rect 18406 27076 18466 27082
rect 24512 27076 24572 27082
rect 26548 27076 26608 27082
rect 17172 27016 18406 27076
rect 18466 27016 24512 27076
rect 24572 27016 26548 27076
rect 17112 27010 17172 27016
rect 18406 27010 18466 27016
rect 24512 27010 24572 27016
rect 26548 27010 26608 27016
rect 27050 27076 27110 27082
rect 28070 27076 28130 27082
rect 29096 27076 29156 27082
rect 27110 27016 28070 27076
rect 28130 27016 29096 27076
rect 27050 27010 27110 27016
rect 28070 27010 28130 27016
rect 29096 27010 29156 27016
rect 29602 27072 29662 27078
rect 30116 27072 30176 27078
rect 30620 27072 30680 27078
rect 31126 27072 31186 27078
rect 29662 27012 30116 27072
rect 30176 27012 30620 27072
rect 30680 27012 31126 27072
rect 31186 27012 31646 27072
rect 31706 27012 31712 27072
rect 29602 27006 29662 27012
rect 30116 27006 30176 27012
rect 30620 27006 30680 27012
rect 31126 27006 31186 27012
rect 21458 26142 21518 26148
rect 23492 26142 23552 26148
rect 25530 26142 25590 26146
rect 20942 26082 20948 26142
rect 21008 26082 21458 26142
rect 21518 26082 23492 26142
rect 23552 26140 25734 26142
rect 27566 26140 27626 26146
rect 28066 26140 28126 26146
rect 28580 26140 28640 26146
rect 29104 26140 29164 26146
rect 29602 26140 29662 26146
rect 30104 26140 30164 26146
rect 23552 26082 25530 26140
rect 21458 26076 21518 26082
rect 23492 26076 23552 26082
rect 25590 26080 27566 26140
rect 27626 26080 28066 26140
rect 28126 26080 28580 26140
rect 28640 26080 29104 26140
rect 29164 26080 29602 26140
rect 29662 26080 30104 26140
rect 30164 26138 30472 26140
rect 30618 26138 30678 26144
rect 31126 26138 31186 26144
rect 31636 26138 31696 26144
rect 30164 26080 30618 26138
rect 25530 26074 25590 26080
rect 27566 26074 27626 26080
rect 28066 26074 28126 26080
rect 28580 26074 28640 26080
rect 29104 26074 29164 26080
rect 29501 26078 30016 26080
rect 29602 26074 29662 26078
rect 30104 26074 30164 26080
rect 30266 26078 30618 26080
rect 30678 26078 31126 26138
rect 31186 26078 31636 26138
rect 30618 26072 30678 26078
rect 31126 26072 31186 26078
rect 31636 26072 31696 26078
rect 20440 26044 20504 26050
rect 22316 26044 22380 26050
rect 20504 25980 22316 26044
rect 20440 25974 20504 25980
rect 22316 25974 22380 25980
rect 26550 26042 26610 26048
rect 32658 26042 32718 26048
rect 26610 25982 32658 26042
rect 26550 25976 26610 25982
rect 32658 25976 32718 25982
rect 21952 25934 22012 25940
rect 22976 25934 23036 25940
rect 24004 25934 24064 25940
rect 19930 25926 19990 25932
rect 20942 25926 21002 25932
rect 18886 25866 18892 25926
rect 18952 25866 19930 25926
rect 19990 25866 20942 25926
rect 22012 25874 22976 25934
rect 23036 25874 24004 25934
rect 21952 25868 22012 25874
rect 22976 25868 23036 25874
rect 24004 25868 24064 25874
rect 30108 25926 30168 25932
rect 31120 25926 31180 25932
rect 32122 25926 32182 25932
rect 19930 25860 19990 25866
rect 20942 25860 21002 25866
rect 30168 25866 31120 25926
rect 31180 25866 32122 25926
rect 30108 25860 30168 25866
rect 31120 25860 31180 25866
rect 32122 25860 32182 25866
rect 19422 25004 19482 25010
rect 21458 25004 21518 25010
rect 21980 25004 22040 25010
rect 22478 25004 22538 25010
rect 23492 25004 23552 25010
rect 23952 25004 24012 25010
rect 24990 25004 24996 25006
rect 19482 24944 21458 25004
rect 21518 24944 21980 25004
rect 22040 24944 22478 25004
rect 22538 25002 23492 25004
rect 22538 25000 23460 25002
rect 22538 24944 22952 25000
rect 19422 24938 19482 24944
rect 21458 24938 21518 24944
rect 21980 24938 22040 24944
rect 22478 24938 22538 24944
rect 22946 24940 22952 24944
rect 23012 24944 23460 25000
rect 23552 24944 23952 25004
rect 24012 24946 24996 25004
rect 25056 25004 25062 25006
rect 25528 25004 25588 25010
rect 27034 25004 27040 25006
rect 25056 24946 25528 25004
rect 24012 24944 25528 24946
rect 25588 24946 27040 25004
rect 27100 25004 27106 25006
rect 27100 25002 27412 25004
rect 27566 25002 27626 25008
rect 29602 25002 29662 25006
rect 27100 25000 27566 25002
rect 27626 25000 29790 25002
rect 31636 25000 31696 25006
rect 27100 24946 27534 25000
rect 25588 24944 27534 24946
rect 23012 24940 23018 24944
rect 23454 24942 23460 24944
rect 23520 24942 23552 24944
rect 23492 24938 23552 24942
rect 23952 24938 24012 24944
rect 25528 24938 25588 24944
rect 25672 24942 26998 24944
rect 27204 24942 27534 24944
rect 27626 24996 28550 25000
rect 28610 24998 29602 25000
rect 27626 24942 28062 24996
rect 27528 24940 27534 24942
rect 27594 24940 27626 24942
rect 27566 24936 27626 24940
rect 28056 24936 28062 24942
rect 28122 24942 28550 24996
rect 28122 24936 28128 24942
rect 28544 24940 28550 24942
rect 28644 24996 29602 24998
rect 28644 24942 29062 24996
rect 28578 24938 28584 24940
rect 28644 24938 28650 24942
rect 29056 24936 29062 24942
rect 29122 24942 29602 24996
rect 29122 24936 29128 24942
rect 29662 24940 31636 25000
rect 29602 24934 29662 24940
rect 31636 24934 31696 24940
rect 15104 24894 15164 24898
rect 20438 24894 20502 24900
rect 30618 24894 30682 24900
rect 15102 24892 20438 24894
rect 15102 24832 15104 24892
rect 15164 24832 20438 24892
rect 15102 24830 20438 24832
rect 20502 24830 30618 24894
rect 15104 24826 15164 24830
rect 20438 24824 20502 24830
rect 30618 24824 30682 24830
rect 18400 24756 18464 24762
rect 18464 24752 33904 24756
rect 18464 24692 24510 24752
rect 18400 24686 18464 24692
rect 24504 24688 24510 24692
rect 24574 24692 33904 24752
rect 33968 24692 33974 24756
rect 24574 24688 24580 24692
rect 17242 24606 17302 24612
rect 26546 24610 26610 24616
rect 17302 24546 18224 24606
rect 18284 24546 26546 24606
rect 32652 24606 32712 24612
rect 26610 24546 32652 24606
rect 17242 24540 17302 24546
rect 26546 24540 26610 24546
rect 32652 24540 32712 24546
rect 18340 24500 18400 24506
rect 18902 24500 18962 24506
rect 19944 24500 20004 24506
rect 20944 24500 21004 24506
rect 24106 24500 24166 24506
rect 25116 24500 25176 24506
rect 26058 24500 26118 24506
rect 18400 24440 18902 24500
rect 18962 24440 19944 24500
rect 20004 24440 20944 24500
rect 21004 24440 24106 24500
rect 24166 24440 25116 24500
rect 25176 24440 26058 24500
rect 18340 24434 18400 24440
rect 18902 24434 18962 24440
rect 19944 24434 20004 24440
rect 20944 24434 21004 24440
rect 24106 24434 24166 24440
rect 25116 24434 25176 24440
rect 26058 24434 26118 24440
rect 18454 24298 18514 24304
rect 21632 24298 21692 24304
rect 25700 24298 25760 24304
rect 29776 24298 29836 24304
rect 32972 24298 33032 24304
rect 18514 24238 21632 24298
rect 21692 24238 25700 24298
rect 25760 24238 29776 24298
rect 29836 24238 32972 24298
rect 18454 24232 18514 24238
rect 21632 24232 21692 24238
rect 25700 24232 25760 24238
rect 29776 24232 29836 24238
rect 32972 24232 33032 24238
rect 19598 23362 19658 23368
rect 21632 23362 21692 23368
rect 23674 23362 23734 23368
rect 25700 23362 25760 23368
rect 27742 23362 27802 23368
rect 29778 23362 29838 23368
rect 31814 23362 31874 23368
rect 19658 23302 21632 23362
rect 21692 23302 23674 23362
rect 23734 23302 25700 23362
rect 25760 23302 27742 23362
rect 27802 23302 29778 23362
rect 29838 23302 31814 23362
rect 19598 23296 19658 23302
rect 21632 23296 21692 23302
rect 23674 23296 23734 23302
rect 25700 23296 25760 23302
rect 27742 23296 27802 23302
rect 29778 23296 29838 23302
rect 31814 23296 31874 23302
rect 20102 23254 20162 23260
rect 20162 23194 21124 23254
rect 21184 23194 22142 23254
rect 22202 23194 23166 23254
rect 23226 23194 24180 23254
rect 24240 23194 25198 23254
rect 25258 23194 26208 23254
rect 26268 23194 27230 23254
rect 27290 23194 28244 23254
rect 28304 23194 29276 23254
rect 29336 23194 30286 23254
rect 30346 23194 31308 23254
rect 31368 23194 31374 23254
rect 20102 23188 20162 23194
rect 19594 22330 19654 22336
rect 23674 22330 23734 22336
rect 27742 22330 27802 22336
rect 31810 22330 31870 22336
rect 34202 22330 34262 22336
rect 12062 22270 19594 22330
rect 19654 22270 23674 22330
rect 23734 22270 27742 22330
rect 27802 22270 31810 22330
rect 31870 22270 34202 22330
rect -7916 16436 -7856 16442
rect -4458 16436 -4398 16442
rect -7856 16376 -4458 16436
rect -7916 16370 -7856 16376
rect -4458 16370 -4398 16376
rect -11022 16268 -11016 16328
rect -10956 16268 -10357 16328
rect -8422 16268 -8416 16328
rect -8356 16268 -7757 16328
rect -11664 15562 -11604 15568
rect -11146 15562 -11086 15568
rect -13297 15502 -13288 15562
rect -13228 15502 -11664 15562
rect -11604 15502 -11146 15562
rect -11664 15496 -11604 15502
rect -11146 15496 -11086 15502
rect -10417 15490 -10357 16268
rect -9064 15562 -9004 15568
rect -8546 15562 -8486 15568
rect -10417 15430 -10343 15490
rect -10283 15430 -10277 15490
rect -10031 15452 -10025 15512
rect -9965 15452 -9959 15512
rect -9675 15502 -9666 15562
rect -9606 15502 -9064 15562
rect -9004 15502 -8546 15562
rect -9064 15496 -9004 15502
rect -8546 15496 -8486 15502
rect -7817 15490 -7757 16268
rect -3080 16162 8190 16418
rect -3080 15870 -2718 16162
rect 8134 15870 8190 16162
rect -3080 15562 8190 15870
rect -11922 15413 -11862 15419
rect -11406 15413 -11346 15419
rect -12495 15353 -12486 15413
rect -12426 15353 -11922 15413
rect -11862 15353 -11406 15413
rect -11346 15353 -10888 15413
rect -10828 15353 -10822 15413
rect -11922 15347 -11862 15353
rect -11406 15347 -11346 15353
rect -11018 14865 -10958 14871
rect -10025 14866 -9965 15452
rect -7817 15430 -7743 15490
rect -7683 15430 -7677 15490
rect -7431 15452 -7425 15512
rect -7365 15452 -7359 15512
rect -9322 15413 -9262 15419
rect -8806 15413 -8746 15419
rect -9859 15353 -9850 15413
rect -9790 15353 -9322 15413
rect -9262 15353 -8806 15413
rect -8746 15353 -8288 15413
rect -8228 15353 -8222 15413
rect -9322 15347 -9262 15353
rect -8806 15347 -8746 15353
rect -8418 14866 -8358 14871
rect -7425 14866 -7365 15452
rect -3080 15240 9272 15562
rect -10511 14865 -7365 14866
rect -10958 14806 -8418 14865
rect -10958 14805 -10407 14806
rect -8358 14806 -7365 14865
rect 12062 14918 12122 22270
rect 19594 22264 19654 22270
rect 23674 22264 23734 22270
rect 27742 22264 27802 22270
rect 31810 22264 31870 22270
rect 34202 22264 34262 22270
rect 17598 22198 17658 22204
rect 22140 22198 22146 22200
rect 17658 22196 22146 22198
rect 17658 22138 20100 22196
rect 17598 22132 17658 22138
rect 20094 22136 20100 22138
rect 20160 22192 22146 22196
rect 20160 22138 21114 22192
rect 20160 22136 20166 22138
rect 21108 22132 21114 22138
rect 21174 22140 22146 22192
rect 22206 22198 22212 22200
rect 23138 22198 23144 22200
rect 22206 22140 23144 22198
rect 23204 22198 23210 22200
rect 24182 22198 24188 22200
rect 23204 22140 24188 22198
rect 24248 22198 24254 22200
rect 28238 22198 28244 22200
rect 24248 22196 28244 22198
rect 24248 22140 25192 22196
rect 21174 22138 25192 22140
rect 21174 22132 21180 22138
rect 25186 22136 25192 22138
rect 25252 22138 26208 22196
rect 25252 22136 25258 22138
rect 26202 22136 26208 22138
rect 26268 22138 27212 22196
rect 26268 22136 26274 22138
rect 27206 22136 27212 22138
rect 27272 22140 28244 22196
rect 28304 22198 28310 22200
rect 33766 22198 33826 22204
rect 28304 22196 33766 22198
rect 28304 22140 29260 22196
rect 27272 22138 29260 22140
rect 27272 22136 27278 22138
rect 29254 22136 29260 22138
rect 29320 22138 30288 22196
rect 29320 22136 29326 22138
rect 30282 22136 30288 22138
rect 30348 22138 31308 22196
rect 30348 22136 30354 22138
rect 31302 22136 31308 22138
rect 31368 22138 33766 22196
rect 31368 22136 31374 22138
rect 33766 22132 33826 22138
rect 24992 21988 25052 21994
rect 25052 21928 26728 21988
rect 26788 21928 26794 21988
rect 32626 21974 32686 21978
rect 32624 21972 33968 21974
rect 24992 21922 25052 21928
rect 32624 21912 32626 21972
rect 32686 21970 33968 21972
rect 32686 21912 33908 21970
rect 32624 21910 33908 21912
rect 33968 21910 33974 21970
rect 32626 21906 32686 21910
rect 26008 21792 26072 21798
rect 30072 21792 30136 21798
rect 31096 21792 31160 21798
rect 32108 21792 32172 21798
rect 26072 21728 30072 21792
rect 30136 21728 31096 21792
rect 31160 21728 32108 21792
rect 26008 21722 26072 21728
rect 30072 21722 30136 21728
rect 31096 21722 31160 21728
rect 32108 21722 32172 21728
rect 18224 21670 18284 21676
rect 19390 21670 19450 21676
rect 21426 21670 21486 21676
rect 18284 21610 19390 21670
rect 19450 21610 21426 21670
rect 18224 21604 18284 21610
rect 19390 21604 19450 21610
rect 21426 21604 21486 21610
rect 21934 21670 21998 21676
rect 26010 21670 26074 21676
rect 21998 21606 26010 21670
rect 21934 21600 21998 21606
rect 26010 21600 26074 21606
rect 29572 21670 29632 21676
rect 31606 21670 31666 21676
rect 34050 21670 34110 21676
rect 29632 21610 31606 21670
rect 31666 21610 34050 21670
rect 29572 21604 29632 21610
rect 31606 21604 31666 21610
rect 34050 21604 34110 21610
rect 17472 21588 17532 21594
rect 17714 21588 17774 21594
rect 17532 21528 17714 21588
rect 17472 21522 17532 21528
rect 17714 21522 17774 21528
rect 20408 20722 20468 20728
rect 22444 20722 22504 20728
rect 20468 20662 22444 20722
rect 20408 20656 20468 20662
rect 22444 20656 22504 20662
rect 22786 20724 22846 20730
rect 25500 20724 25560 20730
rect 22846 20664 25500 20724
rect 22786 20658 22846 20664
rect 25500 20658 25560 20664
rect 30588 20722 30648 20728
rect 32624 20722 32684 20728
rect 30648 20662 32624 20722
rect 30588 20656 30648 20662
rect 14588 20634 14648 20640
rect 15610 20634 15670 20640
rect 14648 20574 15610 20634
rect 14588 20568 14648 20574
rect 15610 20568 15670 20574
rect 17956 20624 18016 20630
rect 30696 20624 30756 20662
rect 32624 20656 32684 20662
rect 18016 20564 30756 20624
rect 17956 20558 18016 20564
rect 14696 20522 14756 20528
rect 15480 20522 15540 20528
rect 14756 20462 15480 20522
rect 14696 20456 14756 20462
rect 15480 20456 15540 20462
rect 18092 20526 18152 20532
rect 20408 20526 20468 20532
rect 18152 20466 20408 20526
rect 18092 20460 18152 20466
rect 20408 20460 20468 20466
rect 21428 20528 21488 20534
rect 26518 20528 26578 20534
rect 33890 20528 33950 20534
rect 21488 20468 26518 20528
rect 26578 20468 33890 20528
rect 21428 20462 21488 20468
rect 26518 20462 26578 20468
rect 33890 20462 33950 20468
rect 19394 20416 19454 20422
rect 21428 20416 21488 20422
rect 19454 20356 21428 20416
rect 19394 20350 19454 20356
rect 21428 20350 21488 20356
rect 24484 20414 24544 20420
rect 26518 20414 26578 20420
rect 24544 20354 26518 20414
rect 24484 20348 24544 20354
rect 26518 20348 26578 20354
rect 29574 20414 29634 20420
rect 31608 20416 31668 20420
rect 31540 20414 31668 20416
rect 34202 20414 34262 20420
rect 29634 20354 31608 20414
rect 31668 20354 34202 20414
rect 29574 20348 29634 20354
rect 31540 20352 31668 20354
rect 31608 20348 31668 20352
rect 34202 20348 34262 20354
rect 12926 19600 12986 19606
rect 16120 19600 16180 19606
rect 12986 19540 16120 19600
rect 12926 19534 12986 19540
rect 16120 19534 16180 19540
rect 14086 19490 14146 19496
rect 17272 19490 17332 19496
rect 14146 19430 17272 19490
rect 30438 19480 30498 19486
rect 14086 19424 14146 19430
rect 17272 19424 17332 19430
rect 17714 19466 17774 19472
rect 24480 19466 24540 19472
rect 25500 19466 25560 19472
rect 27536 19466 27596 19472
rect 17774 19406 24480 19466
rect 24540 19406 25500 19466
rect 25560 19406 27536 19466
rect 30498 19420 34860 19480
rect 30438 19414 30498 19420
rect 17714 19400 17774 19406
rect 24480 19400 24540 19406
rect 25500 19400 25560 19406
rect 27536 19400 27596 19406
rect 30586 19370 30646 19376
rect 32626 19370 32686 19376
rect 33766 19370 33826 19376
rect 17464 19362 17524 19368
rect 22446 19362 22506 19368
rect 29570 19362 29630 19368
rect 17524 19302 20410 19362
rect 20470 19302 22446 19362
rect 22506 19302 29570 19362
rect 30646 19310 32626 19370
rect 32686 19310 33766 19370
rect 30586 19304 30646 19310
rect 32626 19304 32686 19310
rect 33766 19304 33826 19310
rect 17464 19296 17524 19302
rect 22446 19296 22506 19302
rect 29570 19296 29630 19302
rect 22444 19260 22504 19266
rect 31606 19260 31666 19266
rect 17710 19252 17770 19258
rect 18376 19252 18436 19258
rect 17770 19192 18376 19252
rect 22504 19200 31606 19260
rect 22444 19194 22504 19200
rect 31606 19194 31666 19200
rect 17710 19186 17770 19192
rect 18376 19186 18436 19192
rect 20410 19158 20470 19164
rect 22444 19158 22504 19164
rect 20470 19098 22444 19158
rect 20410 19092 20470 19098
rect 22444 19092 22504 19098
rect 25500 19160 25560 19166
rect 26518 19160 26578 19166
rect 27534 19160 27594 19166
rect 30438 19160 30498 19166
rect 25560 19100 26518 19160
rect 26578 19100 27534 19160
rect 27594 19100 30438 19160
rect 25500 19094 25560 19100
rect 26518 19094 26578 19100
rect 27534 19094 27594 19100
rect 30438 19094 30498 19100
rect 30590 19162 30650 19168
rect 32624 19162 32684 19168
rect 33890 19162 33950 19168
rect 30650 19102 32624 19162
rect 32684 19102 33890 19162
rect 33950 19102 34732 19162
rect 30590 19096 30650 19102
rect 32624 19096 32684 19102
rect 33890 19096 33950 19102
rect 14602 18566 14662 18572
rect 15612 18566 15672 18572
rect 12794 18452 12800 18512
rect 12860 18452 12866 18512
rect 14662 18506 15612 18566
rect 14602 18500 14662 18506
rect 15612 18500 15672 18506
rect 14708 18466 14768 18472
rect 15494 18466 15554 18472
rect 12308 17396 12314 17456
rect 12374 17396 12380 17456
rect 12188 16896 12194 16956
rect 12254 16896 12260 16956
rect 12194 15046 12254 16896
rect 12194 14980 12254 14986
rect 12314 15048 12374 17396
rect 12448 17220 12454 17280
rect 12514 17220 12520 17280
rect 12454 15066 12514 17220
rect 12676 16398 12682 16458
rect 12742 16398 12748 16458
rect 12682 15082 12742 16398
rect 12800 15182 12860 18452
rect 14768 18406 15494 18466
rect 14708 18400 14768 18406
rect 15494 18400 15554 18406
rect 22446 18218 22506 18224
rect 24248 18218 24308 18224
rect 17598 18210 17658 18216
rect 19392 18210 19452 18216
rect 21428 18210 21488 18216
rect 17658 18150 19392 18210
rect 19452 18150 21428 18210
rect 22506 18158 24248 18218
rect 22446 18152 22506 18158
rect 24248 18152 24308 18158
rect 24482 18212 24542 18218
rect 26518 18212 26578 18218
rect 24542 18152 26518 18212
rect 17598 18144 17658 18150
rect 13348 17046 13354 17106
rect 13414 17046 13420 17106
rect 13242 16634 13248 16694
rect 13308 16634 13314 16694
rect 13122 16516 13128 16576
rect 13188 16516 13194 16576
rect 13128 15192 13188 16516
rect 13248 15600 13308 16634
rect 13231 15591 13321 15600
rect 13231 15492 13321 15501
rect 12794 15122 12800 15182
rect 12860 15122 12866 15182
rect 13248 15184 13308 15492
rect 13128 15126 13188 15132
rect 13242 15124 13248 15184
rect 13308 15124 13314 15184
rect 13354 15048 13414 17046
rect 12682 15016 12742 15022
rect 12454 15000 12514 15006
rect 13348 14988 13354 15048
rect 13414 14988 13420 15048
rect 12314 14982 12374 14988
rect 12572 14928 12632 14934
rect 17826 14928 17886 18150
rect 19392 18144 19452 18150
rect 21428 18144 21488 18150
rect 24482 18146 24542 18152
rect 26518 18146 26578 18152
rect 29572 18214 29632 18220
rect 31608 18214 31668 18220
rect 29632 18154 31608 18214
rect 29572 18148 29632 18154
rect 31608 18148 31668 18154
rect 21428 18102 21488 18108
rect 26516 18102 26576 18108
rect 33766 18102 33826 18108
rect 21488 18042 26516 18102
rect 26576 18042 33766 18102
rect 21428 18036 21488 18042
rect 26516 18036 26576 18042
rect 33766 18036 33826 18042
rect 18224 18002 18284 18008
rect 18284 17942 30808 18002
rect 18224 17936 18284 17942
rect 20406 17900 20466 17906
rect 22440 17900 22500 17906
rect 20466 17840 22440 17900
rect 30594 17900 30654 17906
rect 30748 17900 30808 17942
rect 32628 17900 32688 17906
rect 20406 17834 20466 17840
rect 22440 17834 22500 17840
rect 22644 17888 22704 17894
rect 22704 17828 26006 17888
rect 26066 17828 27022 17888
rect 27082 17828 30082 17888
rect 30142 17828 30148 17888
rect 30654 17840 32628 17900
rect 30594 17834 30654 17840
rect 32628 17834 32688 17840
rect 22644 17822 22704 17828
rect 17956 16952 18016 16958
rect 19388 16952 19448 16958
rect 21424 16952 21484 16958
rect 18016 16892 19388 16952
rect 19448 16892 21424 16952
rect 17956 16886 18016 16892
rect 19388 16886 19448 16892
rect 21424 16886 21484 16892
rect 29576 16952 29636 16958
rect 31612 16952 31672 16958
rect 29636 16892 31612 16952
rect 29576 16886 29636 16892
rect 18092 16822 18152 16828
rect 29706 16822 29766 16892
rect 31612 16886 31672 16892
rect 18152 16762 29766 16822
rect 18092 16756 18152 16762
rect 22446 16682 22506 16688
rect 34050 16682 34110 16688
rect 22506 16622 34050 16682
rect 22446 16616 22506 16622
rect 12632 14868 17886 14928
rect 12572 14862 12632 14868
rect 12062 14852 12122 14858
rect -8358 14805 -7807 14806
rect -11018 14799 -10958 14805
rect -8418 14799 -8358 14805
rect 24166 14698 24226 16622
rect 24166 14632 24226 14638
rect 29270 14698 29330 16622
rect 33330 14692 33390 16622
rect 34050 16616 34110 16622
rect 29270 14632 29330 14638
rect 33324 14632 33330 14692
rect 33390 14632 33396 14692
rect -13105 14576 -13015 14580
rect -9874 14576 -9774 14585
rect -13110 14571 -9874 14576
rect -13110 14481 -13105 14571
rect -13015 14481 -9874 14571
rect -13110 14476 -9874 14481
rect -9774 14476 -9766 14576
rect -13105 14472 -13015 14476
rect -9874 14467 -9774 14476
rect -13499 14354 -13409 14358
rect -9686 14354 -9586 14363
rect -13504 14349 -9686 14354
rect -13504 14259 -13499 14349
rect -13409 14259 -9686 14349
rect -13504 14254 -9686 14259
rect 9350 14320 9410 14326
rect 13128 14320 13188 14326
rect 9410 14260 13128 14320
rect 9350 14254 9410 14260
rect 13128 14254 13188 14260
rect -13499 14250 -13409 14254
rect -9686 14245 -9586 14254
rect 10876 14186 10936 14192
rect 12682 14186 12742 14192
rect 10936 14126 12682 14186
rect 10876 14120 10936 14126
rect 12682 14120 12742 14126
rect 12924 12962 12984 12968
rect 12984 12902 14498 12962
rect 14558 12902 14564 12962
rect 12924 12896 12984 12902
rect 15512 12746 15572 12752
rect 17552 12746 17612 12752
rect 19592 12746 19652 12752
rect 21622 12746 21682 12752
rect 23662 12746 23722 12752
rect 25694 12746 25754 12752
rect 27734 12746 27794 12752
rect 29770 12746 29830 12752
rect 31804 12746 31864 12752
rect 15572 12686 17552 12746
rect 17612 12686 19592 12746
rect 19652 12686 21622 12746
rect 21682 12686 23662 12746
rect 23722 12686 25694 12746
rect 25754 12686 27734 12746
rect 27794 12686 29770 12746
rect 29830 12686 31804 12746
rect 15512 12680 15572 12686
rect 17552 12680 17612 12686
rect 19592 12680 19652 12686
rect 21622 12680 21682 12686
rect 23662 12680 23722 12686
rect 25694 12680 25754 12686
rect 27734 12680 27794 12686
rect 29770 12680 29830 12686
rect 31804 12680 31864 12686
rect 13136 12626 13196 12632
rect 13480 12626 13540 12632
rect 13196 12566 13480 12626
rect 13136 12560 13196 12566
rect 13480 12560 13540 12566
rect 15004 12620 15064 12626
rect 23148 12620 23208 12626
rect 15064 12560 16018 12620
rect 16078 12560 17040 12620
rect 17100 12560 18054 12620
rect 18114 12560 19080 12620
rect 19140 12560 20092 12620
rect 20152 12560 21128 12620
rect 21188 12560 22134 12620
rect 22194 12560 23148 12620
rect 23208 12560 24164 12620
rect 24224 12560 25172 12620
rect 25232 12560 26188 12620
rect 26248 12560 27212 12620
rect 27272 12560 28234 12620
rect 28294 12560 29256 12620
rect 29316 12560 30274 12620
rect 30334 12560 31288 12620
rect 31348 12560 32312 12620
rect 32372 12560 32378 12620
rect 15004 12554 15064 12560
rect 23148 12554 23208 12560
rect 13354 12504 13414 12510
rect 18568 12504 18628 12510
rect 28756 12504 28816 12510
rect 32828 12504 32888 12510
rect 33960 12504 34020 12510
rect 13414 12444 18568 12504
rect 18628 12444 28756 12504
rect 28816 12444 32828 12504
rect 32888 12444 33960 12504
rect 13354 12438 13414 12444
rect 18568 12438 18628 12444
rect 28756 12438 28816 12444
rect 32828 12438 32888 12444
rect 33960 12438 34020 12444
rect 15516 11582 15576 11588
rect 17556 11582 17616 11588
rect 19588 11582 19648 11588
rect 21620 11582 21680 11588
rect 23656 11582 23716 11588
rect 25692 11582 25752 11588
rect 27730 11582 27790 11588
rect 29768 11582 29828 11588
rect 31804 11582 31864 11588
rect 15576 11522 17556 11582
rect 17616 11522 19588 11582
rect 19648 11522 21620 11582
rect 21680 11522 23656 11582
rect 23716 11522 25692 11582
rect 25752 11522 27730 11582
rect 27790 11522 29768 11582
rect 29828 11522 31804 11582
rect 15516 11516 15576 11522
rect 17556 11516 17616 11522
rect 19588 11516 19648 11522
rect 21620 11516 21680 11522
rect 23656 11516 23716 11522
rect 25692 11516 25752 11522
rect 27730 11516 27790 11522
rect 29768 11516 29828 11522
rect 31804 11516 31864 11522
rect 15008 11472 15068 11478
rect 16030 11472 16090 11478
rect 17044 11472 17104 11478
rect 18058 11472 18118 11478
rect 19076 11472 19136 11478
rect 20102 11472 20162 11478
rect 21122 11472 21182 11478
rect 22142 11472 22202 11478
rect 23144 11472 23204 11478
rect 24170 11472 24230 11478
rect 25188 11472 25248 11478
rect 26196 11472 26256 11478
rect 27208 11472 27268 11478
rect 28240 11472 28300 11478
rect 29254 11472 29314 11478
rect 30272 11472 30332 11478
rect 31296 11472 31356 11478
rect 32316 11472 32376 11478
rect 15068 11412 16030 11472
rect 16090 11412 17044 11472
rect 17104 11412 18058 11472
rect 18118 11412 19076 11472
rect 19136 11412 20102 11472
rect 20162 11412 21122 11472
rect 21182 11412 22142 11472
rect 22202 11412 23144 11472
rect 23204 11412 24170 11472
rect 24230 11412 25188 11472
rect 25248 11412 26196 11472
rect 26256 11412 27208 11472
rect 27268 11412 28240 11472
rect 28300 11412 29254 11472
rect 29314 11412 30272 11472
rect 30332 11412 31296 11472
rect 31356 11412 32316 11472
rect 15008 11406 15068 11412
rect 16030 11406 16090 11412
rect 17044 11406 17104 11412
rect 18058 11406 18118 11412
rect 19076 11406 19136 11412
rect 20102 11406 20162 11412
rect 21122 11406 21182 11412
rect 22142 11406 22202 11412
rect 23144 11406 23204 11412
rect 24170 11406 24230 11412
rect 25188 11406 25248 11412
rect 26196 11406 26256 11412
rect 27208 11406 27268 11412
rect 28240 11406 28300 11412
rect 29254 11406 29314 11412
rect 30272 11406 30332 11412
rect 31296 11406 31356 11412
rect 32316 11406 32376 11412
rect 13032 11366 13092 11372
rect 14498 11366 14558 11372
rect 16538 11366 16598 11372
rect 18568 11366 18628 11372
rect 20608 11366 20668 11372
rect 22642 11366 22702 11372
rect 24678 11366 24738 11372
rect 26714 11366 26774 11372
rect 28754 11366 28814 11372
rect 30784 11366 30844 11372
rect 32824 11366 32884 11372
rect 13092 11306 14498 11366
rect 14558 11306 16538 11366
rect 16598 11306 18568 11366
rect 18628 11306 20608 11366
rect 20668 11306 22642 11366
rect 22702 11306 24678 11366
rect 24738 11306 26714 11366
rect 26774 11306 28754 11366
rect 28814 11306 30784 11366
rect 30844 11306 32824 11366
rect 13032 11300 13092 11306
rect 14498 11300 14558 11306
rect 16538 11300 16598 11306
rect 18568 11300 18628 11306
rect 20608 11300 20668 11306
rect 22642 11300 22702 11306
rect 24678 11300 24738 11306
rect 26714 11300 26774 11306
rect 28754 11300 28814 11306
rect 30784 11300 30844 11306
rect 32824 11300 32884 11306
rect 13484 11260 13544 11266
rect 13982 11260 14042 11266
rect 14494 11260 14554 11266
rect 20774 11260 20834 11266
rect 22642 11260 22702 11266
rect 24680 11260 24740 11266
rect 26560 11260 26620 11266
rect 12792 11200 12798 11260
rect 12858 11200 13484 11260
rect 13544 11200 13982 11260
rect 14042 11200 14494 11260
rect 14554 11200 20774 11260
rect 20834 11200 22642 11260
rect 22702 11200 24680 11260
rect 24740 11200 26560 11260
rect 13484 11194 13544 11200
rect 13982 11194 14042 11200
rect 14494 11194 14554 11200
rect 20774 11194 20834 11200
rect 22642 11194 22702 11200
rect 24680 11194 24740 11200
rect 26560 11194 26620 11200
rect 30784 11262 30844 11268
rect 33960 11262 34020 11268
rect 30844 11202 33960 11262
rect 30784 11196 30844 11202
rect 33960 11196 34020 11202
rect -11022 11009 -10932 11014
rect -11026 10929 -11017 11009
rect -10937 10929 -10928 11009
rect -6664 11001 -6578 11006
rect -11022 10869 -10932 10929
rect -6668 10925 -6659 11001
rect -6583 10925 -6574 11001
rect -6664 10871 -6578 10925
rect -11022 10779 -8595 10869
rect -6664 10785 -4371 10871
rect -8685 10703 -8595 10779
rect -8685 10604 -8595 10613
rect -4457 10689 -4371 10785
rect -4457 10594 -4371 10603
rect 13354 10370 13414 10376
rect 16532 10370 16592 10376
rect 19588 10370 19648 10376
rect 25694 10370 25754 10376
rect 30788 10370 30848 10376
rect 13414 10310 16532 10370
rect 16592 10310 19588 10370
rect 19648 10310 25694 10370
rect 25754 10310 30788 10370
rect 13354 10304 13414 10310
rect 16532 10304 16592 10310
rect 19588 10304 19648 10310
rect 25694 10304 25754 10310
rect 30788 10304 30848 10310
rect 12924 10266 12984 10272
rect 13478 10266 13538 10272
rect 14998 10266 15058 10272
rect 12984 10206 13478 10266
rect 13538 10206 14998 10266
rect 12924 10200 12984 10206
rect 13478 10200 13538 10206
rect 14998 10200 15058 10206
rect 15510 10266 15570 10272
rect 16534 10266 16594 10272
rect 17546 10266 17606 10272
rect 18566 10266 18626 10272
rect 21624 10266 21684 10272
rect 23662 10266 23722 10272
rect 26712 10266 26772 10272
rect 27730 10266 27790 10272
rect 28750 10266 28810 10272
rect 29766 10266 29826 10272
rect 31802 10266 31862 10272
rect 15570 10206 16534 10266
rect 16594 10206 17546 10266
rect 17606 10206 18566 10266
rect 18626 10206 21624 10266
rect 21684 10206 23662 10266
rect 23722 10206 26712 10266
rect 26772 10206 27730 10266
rect 27790 10206 28750 10266
rect 28810 10206 29766 10266
rect 29826 10206 31802 10266
rect 15510 10200 15570 10206
rect 16534 10200 16594 10206
rect 17546 10200 17606 10206
rect 18566 10200 18626 10206
rect 21624 10200 21684 10206
rect 23662 10200 23722 10206
rect 26712 10200 26772 10206
rect 27730 10200 27790 10206
rect 28750 10200 28810 10206
rect 29766 10200 29826 10206
rect 31802 10200 31862 10206
rect 13248 10144 13308 10150
rect 20608 10144 20668 10150
rect 22642 10144 22702 10150
rect 24672 10144 24732 10150
rect 34672 10144 34732 19102
rect 13308 10084 20608 10144
rect 20668 10084 22642 10144
rect 22702 10084 24672 10144
rect 24732 10084 34732 10144
rect 13248 10078 13308 10084
rect 20608 10078 20668 10084
rect 22642 10078 22702 10084
rect 24672 10078 24732 10084
rect 13136 10030 13196 10036
rect 13984 10030 14044 10036
rect 13196 9970 13984 10030
rect 13136 9964 13196 9970
rect 13984 9964 14044 9970
rect 15516 10032 15576 10038
rect 17552 10032 17612 10038
rect 33946 10032 34006 10038
rect 15576 9972 17552 10032
rect 17612 9972 33946 10032
rect 15516 9966 15576 9972
rect 17552 9966 17612 9972
rect 33946 9966 34006 9972
rect 34074 10014 34134 10020
rect 34674 10014 34734 10020
rect 34134 9954 34674 10014
rect 34074 9948 34134 9954
rect 34674 9948 34734 9954
rect 33840 9144 33900 9150
rect 34800 9144 34860 19420
rect 16532 9126 16592 9132
rect 18568 9126 18628 9132
rect 26712 9126 26772 9132
rect 28748 9126 28808 9132
rect 32822 9126 32882 9132
rect 13360 9102 13420 9108
rect 14498 9102 14558 9108
rect 13420 9042 14498 9102
rect 14558 9042 15380 9102
rect 16592 9066 18568 9126
rect 18628 9066 26712 9126
rect 26772 9066 28748 9126
rect 28808 9066 32822 9126
rect 33900 9084 34860 9144
rect 33840 9078 33900 9084
rect 16532 9060 16592 9066
rect 18568 9060 18628 9066
rect 26712 9060 26772 9066
rect 28748 9060 28808 9066
rect 32822 9060 32882 9066
rect 13360 9036 13420 9042
rect 14498 9036 14558 9042
rect 13248 8902 13308 8908
rect 14496 8902 14556 8908
rect 13308 8842 14496 8902
rect 15320 8906 15380 9042
rect 15514 9022 15574 9028
rect 17554 9022 17614 9028
rect 19586 9022 19646 9028
rect 21620 9022 21680 9028
rect 23660 9022 23720 9028
rect 25694 9022 25754 9028
rect 15574 8962 17554 9022
rect 17614 8962 19586 9022
rect 19646 8962 21620 9022
rect 21680 8962 23660 9022
rect 23720 8962 25694 9022
rect 15514 8956 15574 8962
rect 17554 8956 17614 8962
rect 19586 8956 19646 8962
rect 21620 8956 21680 8962
rect 23660 8956 23720 8962
rect 25694 8956 25754 8962
rect 25890 9018 25950 9024
rect 30782 9018 30842 9024
rect 25950 8958 30782 9018
rect 34440 9014 34500 9020
rect 25890 8952 25950 8958
rect 30782 8952 30842 8958
rect 31280 8954 31286 9014
rect 31346 8954 34440 9014
rect 34440 8948 34500 8954
rect 16028 8908 16088 8914
rect 19586 8910 19646 8916
rect 21622 8910 21682 8916
rect 23658 8910 23718 8916
rect 25694 8910 25754 8916
rect 27728 8910 27788 8916
rect 29766 8910 29826 8916
rect 31806 8910 31866 8916
rect 34190 8910 34250 8916
rect 15320 8848 16028 8906
rect 16088 8848 17032 8908
rect 17092 8848 18044 8908
rect 18104 8848 19064 8908
rect 19124 8848 19130 8908
rect 19646 8850 21622 8910
rect 21682 8850 23658 8910
rect 23718 8850 25694 8910
rect 25754 8850 27728 8910
rect 27788 8850 29766 8910
rect 29826 8850 31806 8910
rect 31866 8850 34190 8910
rect 15320 8846 16370 8848
rect 16028 8842 16088 8846
rect 19586 8844 19646 8850
rect 21622 8844 21682 8850
rect 23658 8844 23718 8850
rect 25694 8844 25754 8850
rect 27728 8844 27788 8850
rect 29766 8844 29826 8850
rect 31806 8844 31866 8850
rect 34190 8844 34250 8850
rect 13248 8836 13308 8842
rect 14496 8836 14556 8842
rect 12572 8800 12632 8806
rect 13142 8800 13202 8806
rect 20604 8800 20664 8806
rect 22638 8800 22698 8806
rect 24678 8800 24738 8806
rect 25890 8800 25950 8806
rect 12632 8740 13142 8800
rect 13202 8740 20604 8800
rect 20664 8740 22638 8800
rect 22698 8740 24678 8800
rect 24738 8740 25890 8800
rect 12572 8734 12632 8740
rect 13142 8734 13202 8740
rect 20604 8734 20664 8740
rect 22638 8734 22698 8740
rect 24678 8734 24738 8740
rect 25890 8734 25950 8740
rect 26184 8802 26244 8808
rect 26244 8742 27212 8802
rect 27272 8742 27278 8802
rect 27730 8796 27790 8802
rect 29766 8796 29826 8802
rect 31804 8796 31864 8802
rect 33946 8796 34006 8802
rect 26184 8736 26244 8742
rect 27790 8736 29766 8796
rect 29826 8736 31804 8796
rect 31864 8736 33946 8796
rect 27730 8730 27790 8736
rect 29766 8730 29826 8736
rect 31804 8730 31864 8736
rect 33946 8730 34006 8736
rect 30278 7882 30338 7888
rect 14496 7870 14556 7876
rect 16534 7870 16594 7876
rect 18570 7870 18630 7876
rect 20602 7870 20662 7876
rect 14556 7810 16534 7870
rect 16594 7810 18570 7870
rect 18630 7810 20602 7870
rect 25178 7822 25184 7882
rect 25244 7822 30278 7882
rect 30278 7816 30338 7822
rect 30416 7886 30476 7892
rect 31298 7886 31358 7892
rect 32304 7886 32364 7892
rect 30476 7826 31298 7886
rect 31358 7826 32304 7886
rect 30416 7820 30476 7826
rect 31298 7820 31358 7826
rect 32304 7820 32364 7826
rect 32822 7882 32882 7888
rect 34074 7882 34134 7888
rect 32882 7822 34074 7882
rect 32822 7816 32882 7822
rect 34074 7816 34134 7822
rect 14496 7804 14556 7810
rect 16534 7804 16594 7810
rect 18570 7804 18630 7810
rect 20602 7804 20662 7810
rect 15002 7768 15062 7774
rect 20094 7768 20154 7774
rect 12062 7718 12122 7724
rect 15062 7708 20094 7768
rect 15002 7702 15062 7708
rect 20094 7702 20154 7708
rect 24678 7754 24738 7760
rect 32822 7754 32882 7760
rect 24738 7694 32822 7754
rect 24678 7688 24738 7694
rect 32822 7688 32882 7694
rect 7514 6792 7574 6798
rect 12062 6792 12122 7658
rect 13248 7666 13308 7672
rect 16532 7666 16592 7672
rect 13308 7606 16532 7666
rect 13248 7600 13308 7606
rect 16532 7600 16592 7606
rect 17040 7660 17100 7666
rect 18062 7660 18122 7666
rect 19076 7660 19136 7666
rect 20094 7660 20154 7666
rect 21114 7660 21174 7666
rect 28226 7660 28286 7666
rect 29256 7660 29316 7666
rect 30416 7660 30476 7666
rect 17100 7600 18062 7660
rect 18122 7600 19076 7660
rect 19136 7600 20094 7660
rect 20154 7600 21114 7660
rect 21174 7600 28226 7660
rect 28286 7600 29256 7660
rect 29316 7600 30416 7660
rect 17040 7594 17100 7600
rect 18062 7594 18122 7600
rect 19076 7594 19136 7600
rect 20094 7594 20154 7600
rect 21114 7594 21174 7600
rect 28226 7594 28286 7600
rect 29256 7594 29316 7600
rect 30416 7594 30476 7600
rect 30784 7660 30844 7666
rect 34312 7660 34372 7666
rect 30844 7600 34312 7660
rect 30784 7594 30844 7600
rect 34312 7594 34372 7600
rect 15516 7566 15576 7572
rect 17550 7566 17610 7572
rect 19586 7566 19646 7572
rect 15576 7506 17550 7566
rect 17610 7506 19586 7566
rect 15516 7500 15576 7506
rect 17550 7500 17610 7506
rect 19586 7500 19646 7506
rect 26714 7556 26774 7562
rect 30784 7556 30844 7562
rect 26774 7496 30784 7556
rect 26714 7490 26774 7496
rect 30784 7490 30844 7496
rect 31800 7558 31860 7564
rect 34190 7558 34250 7564
rect 31860 7498 34190 7558
rect 31800 7492 31860 7498
rect 34190 7492 34250 7498
rect 7574 6732 12122 6792
rect 7514 6726 7574 6732
rect 5484 6646 5544 6652
rect 9544 6646 9604 6652
rect 11728 6646 11788 6652
rect 12194 6646 12254 6652
rect 21622 6648 21682 6654
rect 23658 6648 23718 6654
rect 25694 6648 25754 6654
rect 27732 6648 27792 6654
rect 1398 6586 1404 6646
rect 1464 6586 5484 6646
rect 5544 6586 9544 6646
rect 9604 6586 11728 6646
rect 11788 6586 12194 6646
rect 5484 6580 5544 6586
rect 9544 6580 9604 6586
rect 11728 6580 11788 6586
rect 12194 6580 12254 6586
rect 14998 6642 15058 6648
rect 15908 6642 15968 6648
rect 16910 6642 16970 6648
rect 18062 6642 18122 6648
rect 19072 6642 19132 6648
rect 20078 6642 20138 6648
rect 21122 6642 21182 6648
rect 15058 6582 15908 6642
rect 15968 6582 16910 6642
rect 16970 6582 18062 6642
rect 18122 6582 19072 6642
rect 19132 6582 20078 6642
rect 20138 6582 21122 6642
rect 21682 6588 23658 6648
rect 23718 6588 25694 6648
rect 25754 6588 27732 6648
rect 21622 6582 21682 6588
rect 23658 6582 23718 6588
rect 25694 6582 25754 6588
rect 27732 6582 27792 6588
rect 29768 6648 29828 6654
rect 31806 6648 31866 6654
rect 29828 6588 31806 6648
rect 29768 6582 29828 6588
rect 31806 6582 31866 6588
rect 14998 6576 15058 6582
rect 15908 6576 15968 6582
rect 16910 6576 16970 6582
rect 18062 6576 18122 6582
rect 19072 6576 19132 6582
rect 20078 6576 20138 6582
rect 21122 6576 21182 6582
rect 17550 6540 17610 6546
rect 27724 6540 27784 6546
rect 29764 6540 29824 6546
rect 31802 6540 31862 6546
rect 250 6518 310 6524
rect 2928 6518 2988 6524
rect 3960 6518 4020 6524
rect 7020 6518 7080 6524
rect 8016 6518 8076 6524
rect 12314 6518 12374 6524
rect -1851 6458 -1842 6518
rect -1782 6458 250 6518
rect 310 6458 2928 6518
rect 2988 6458 3960 6518
rect 4020 6458 7020 6518
rect 7080 6458 8016 6518
rect 8076 6458 12314 6518
rect 17610 6480 27724 6540
rect 27784 6480 29764 6540
rect 29824 6480 31802 6540
rect 17550 6474 17610 6480
rect 27724 6474 27784 6480
rect 29764 6474 29824 6480
rect 31802 6474 31862 6480
rect 250 6452 310 6458
rect 2928 6452 2988 6458
rect 3960 6452 4020 6458
rect 7020 6452 7080 6458
rect 8016 6452 8076 6458
rect 12314 6452 12374 6458
rect 14998 6426 15058 6432
rect 17050 6426 17110 6432
rect 20076 6426 20136 6432
rect 21116 6426 21176 6432
rect 22130 6426 22190 6432
rect 23138 6426 23198 6432
rect 24182 6426 24242 6432
rect 25172 6426 25232 6432
rect 26190 6426 26250 6432
rect 27224 6426 27284 6432
rect 30256 6426 30316 6432
rect 31294 6426 31354 6432
rect 32320 6426 32380 6432
rect 15058 6366 16036 6426
rect 16096 6366 17050 6426
rect 17110 6366 20076 6426
rect 20136 6366 21116 6426
rect 21176 6366 22130 6426
rect 22190 6366 23138 6426
rect 23198 6366 24182 6426
rect 24242 6366 25172 6426
rect 25232 6366 26190 6426
rect 26250 6366 27224 6426
rect 27284 6366 30256 6426
rect 30316 6366 31294 6426
rect 31354 6366 32320 6426
rect 32380 6366 34438 6426
rect 34498 6366 34504 6426
rect 14998 6360 15058 6366
rect 17050 6360 17110 6366
rect 20076 6360 20136 6366
rect 21116 6360 21176 6366
rect 22130 6360 22190 6366
rect 23138 6360 23198 6366
rect 24182 6360 24242 6366
rect 25172 6360 25232 6366
rect 26190 6360 26250 6366
rect 27224 6360 27284 6366
rect 30256 6360 30316 6366
rect 31294 6360 31354 6366
rect 32320 6360 32380 6366
rect 20600 6322 20660 6328
rect 22642 6322 22702 6328
rect 24680 6322 24740 6328
rect 26714 6322 26774 6328
rect 28748 6324 28808 6330
rect 30782 6324 30842 6330
rect 32824 6324 32884 6330
rect 34074 6324 34134 6330
rect 13356 6262 13362 6322
rect 13422 6262 20600 6322
rect 20660 6262 22642 6322
rect 22702 6262 24680 6322
rect 24740 6262 26714 6322
rect 20600 6256 20660 6262
rect 22642 6256 22702 6262
rect 24680 6256 24740 6262
rect 26714 6256 26774 6262
rect 27226 6318 27286 6324
rect 28248 6318 28308 6324
rect 27286 6258 28248 6318
rect 28808 6264 30782 6324
rect 30842 6264 32824 6324
rect 32884 6264 34074 6324
rect 28748 6258 28808 6264
rect 30782 6258 30842 6264
rect 32824 6258 32884 6264
rect 34074 6258 34134 6264
rect 27226 6252 27286 6258
rect 28248 6252 28308 6258
rect -1566 5556 -1506 5565
rect 1908 5556 1968 5562
rect 2932 5556 2992 5562
rect 3964 5556 4024 5562
rect 4964 5556 5024 5562
rect 5984 5556 6044 5562
rect 7004 5556 7064 5562
rect 9028 5556 9088 5562
rect 11848 5556 11908 5562
rect 12454 5556 12514 5562
rect -1506 5496 1908 5556
rect 1968 5496 2932 5556
rect 2992 5496 3964 5556
rect 4024 5496 4964 5556
rect 5024 5496 5984 5556
rect 6044 5496 7004 5556
rect 7064 5496 8014 5556
rect 8074 5496 9028 5556
rect 9088 5496 10046 5556
rect 10106 5496 11848 5556
rect 11908 5496 12454 5556
rect -1566 5487 -1506 5496
rect 1908 5490 1968 5496
rect 2932 5490 2992 5496
rect 3964 5490 4024 5496
rect 4964 5490 5024 5496
rect 5984 5490 6044 5496
rect 7004 5490 7064 5496
rect 9028 5490 9088 5496
rect 11848 5490 11908 5496
rect 12454 5490 12514 5496
rect 1408 5452 1468 5458
rect 3444 5452 3504 5458
rect 5480 5452 5540 5458
rect 7514 5452 7574 5458
rect 9550 5452 9610 5458
rect 1468 5392 3444 5452
rect 3504 5392 5480 5452
rect 5540 5392 7514 5452
rect 7574 5392 9550 5452
rect 19590 5420 19650 5426
rect 23658 5420 23718 5426
rect 25692 5420 25752 5426
rect 1408 5386 1468 5392
rect 3444 5386 3504 5392
rect 5480 5386 5540 5392
rect 7514 5386 7574 5392
rect 9550 5386 9610 5392
rect 14996 5414 15056 5420
rect 16004 5414 16064 5420
rect 17018 5414 17078 5420
rect 18056 5414 18116 5420
rect 19074 5414 19134 5420
rect 15056 5354 16004 5414
rect 16064 5354 17018 5414
rect 17078 5354 18056 5414
rect 18116 5354 19074 5414
rect 19650 5360 21626 5420
rect 21686 5360 23658 5420
rect 23718 5360 25692 5420
rect 19590 5354 19650 5360
rect 23658 5354 23718 5360
rect 25692 5354 25752 5360
rect 26714 5422 26774 5428
rect 27068 5422 27128 5428
rect 26774 5362 27068 5422
rect 26714 5356 26774 5362
rect 27068 5356 27128 5362
rect 30786 5422 30846 5428
rect 34070 5422 34130 5428
rect 30846 5362 34070 5422
rect 30786 5356 30846 5362
rect 34070 5356 34130 5362
rect 6494 5348 6554 5354
rect 13032 5348 13092 5354
rect 14996 5348 15056 5354
rect 16004 5348 16064 5354
rect 17018 5348 17078 5354
rect 18056 5348 18116 5354
rect 19074 5348 19134 5354
rect 2420 5288 2426 5348
rect 2486 5288 4462 5348
rect 4522 5288 6494 5348
rect 6554 5288 8528 5348
rect 8588 5288 10572 5348
rect 10632 5288 13032 5348
rect 6494 5282 6554 5288
rect 13032 5282 13092 5288
rect 13142 5310 13202 5316
rect 14498 5310 14558 5316
rect 22642 5310 22702 5316
rect 24678 5310 24738 5316
rect 26710 5310 26770 5316
rect 13202 5250 14498 5310
rect 14558 5250 22642 5310
rect 22702 5250 24678 5310
rect 24738 5250 26710 5310
rect 13142 5244 13202 5250
rect 14498 5244 14558 5250
rect 22642 5244 22702 5250
rect 24678 5244 24738 5250
rect 26710 5244 26770 5250
rect 26220 5212 26280 5218
rect 27258 5212 27318 5218
rect 28234 5212 28294 5218
rect 29250 5212 29310 5218
rect 31276 5212 31336 5218
rect 32306 5212 32366 5218
rect 12800 5198 12860 5204
rect 15514 5198 15574 5204
rect 17552 5198 17612 5204
rect 21624 5198 21684 5204
rect 12860 5138 15514 5198
rect 15574 5138 17552 5198
rect 17612 5138 21624 5198
rect 26280 5152 27258 5212
rect 27318 5152 28234 5212
rect 28294 5152 29250 5212
rect 29310 5152 31276 5212
rect 31336 5152 32306 5212
rect 26220 5146 26280 5152
rect 27258 5146 27318 5152
rect 28234 5146 28294 5152
rect 29250 5146 29310 5152
rect 31276 5146 31336 5152
rect 32306 5146 32366 5152
rect 12800 5132 12860 5138
rect 15514 5132 15574 5138
rect 17552 5132 17612 5138
rect 21624 5132 21684 5138
rect 14494 5100 14554 5106
rect 16532 5100 16592 5106
rect 18572 5100 18632 5106
rect 20608 5100 20668 5106
rect 26712 5100 26772 5106
rect 27062 5100 27068 5104
rect 14554 5040 16532 5100
rect 16592 5040 18572 5100
rect 18632 5040 20608 5100
rect 20668 5044 27068 5100
rect 27128 5100 27134 5104
rect 28748 5100 28808 5106
rect 30784 5100 30844 5106
rect 32820 5100 32880 5106
rect 27128 5044 28748 5100
rect 20668 5040 28748 5044
rect 28808 5040 30784 5100
rect 30844 5040 32820 5100
rect 14494 5034 14554 5040
rect 16532 5034 16592 5040
rect 18572 5034 18632 5040
rect 20608 5034 20668 5040
rect 26712 5034 26772 5040
rect 28748 5034 28808 5040
rect 30784 5034 30844 5040
rect 32820 5034 32880 5040
rect 3438 4406 3498 4412
rect 7514 4406 7574 4412
rect 11728 4406 11788 4412
rect 3498 4346 7514 4406
rect 7574 4346 11728 4406
rect 3438 4340 3498 4346
rect 7514 4340 7574 4346
rect 11728 4340 11788 4346
rect 250 4286 310 4292
rect 1900 4286 1960 4292
rect 4970 4286 5030 4292
rect 5978 4286 6038 4292
rect 9040 4286 9100 4292
rect 10066 4286 10126 4292
rect 310 4226 1900 4286
rect 1960 4226 4970 4286
rect 5030 4226 5978 4286
rect 6038 4226 9040 4286
rect 9100 4226 10066 4286
rect 250 4220 310 4226
rect 1900 4220 1960 4226
rect 4970 4220 5030 4226
rect 5978 4220 6038 4226
rect 9040 4220 9100 4226
rect 10066 4220 10126 4226
rect 21620 4196 21680 4202
rect 23662 4196 23722 4202
rect 25694 4196 25754 4202
rect 27734 4196 27794 4202
rect 34190 4196 34250 4202
rect 15514 4176 15574 4182
rect 17550 4176 17610 4182
rect 19588 4176 19648 4182
rect 15574 4116 17550 4176
rect 17610 4116 19588 4176
rect 21444 4136 21450 4196
rect 21510 4136 21620 4196
rect 21680 4136 23662 4196
rect 23722 4136 25694 4196
rect 25754 4136 27734 4196
rect 27794 4136 34190 4196
rect 21620 4130 21680 4136
rect 23662 4130 23722 4136
rect 25694 4130 25754 4136
rect 27734 4130 27794 4136
rect 34190 4130 34250 4136
rect 15514 4110 15574 4116
rect 17550 4110 17610 4116
rect 19588 4110 19648 4116
rect 26712 4098 26772 4104
rect 32818 4098 32878 4104
rect 34070 4098 34130 4104
rect 13360 4078 13420 4084
rect 16532 4078 16592 4084
rect 13420 4018 16532 4078
rect 13360 4012 13420 4018
rect 16532 4012 16592 4018
rect 18056 4078 18116 4084
rect 21104 4078 21164 4084
rect 18116 4018 19078 4078
rect 19138 4018 20100 4078
rect 20160 4018 21104 4078
rect 26772 4038 32818 4098
rect 32878 4038 34070 4098
rect 26712 4032 26772 4038
rect 32818 4032 32878 4038
rect 34070 4032 34130 4038
rect 18056 4012 18116 4018
rect 21104 4012 21164 4018
rect 21626 3988 21686 3994
rect 23654 3988 23714 3994
rect 25698 3988 25758 3994
rect 27726 3988 27786 3994
rect 29764 3988 29824 3994
rect 31804 3988 31864 3994
rect 15518 3982 15578 3988
rect 17554 3982 17614 3988
rect 19582 3982 19642 3988
rect 21450 3982 21510 3988
rect 15578 3922 17554 3982
rect 17614 3922 19582 3982
rect 19642 3922 21450 3982
rect 21686 3928 23654 3988
rect 23714 3928 25698 3988
rect 25758 3928 27726 3988
rect 27786 3928 29764 3988
rect 29824 3928 31804 3988
rect 21626 3922 21686 3928
rect 23654 3922 23714 3928
rect 25698 3922 25758 3928
rect 27726 3922 27786 3928
rect 29764 3922 29824 3928
rect 31804 3922 31864 3928
rect 32322 3992 32382 3998
rect 33834 3992 33894 3998
rect 34440 3992 34500 3998
rect 32382 3932 33834 3992
rect 33894 3932 34440 3992
rect 32322 3926 32382 3932
rect 33834 3926 33894 3932
rect 34440 3926 34500 3932
rect 15518 3916 15578 3922
rect 17554 3916 17614 3922
rect 19582 3916 19642 3922
rect 21450 3916 21510 3922
rect 14500 3862 14560 3868
rect 18568 3862 18628 3868
rect 20602 3862 20662 3868
rect 28752 3862 28812 3868
rect 30782 3862 30842 3868
rect 32822 3864 32882 3870
rect 34312 3864 34372 3870
rect 14560 3802 18568 3862
rect 18628 3802 20602 3862
rect 20662 3802 28752 3862
rect 28812 3802 30782 3862
rect 31302 3804 31308 3864
rect 31368 3804 32822 3864
rect 32882 3804 34312 3864
rect 14500 3796 14560 3802
rect 18568 3796 18628 3802
rect 20602 3796 20662 3802
rect 28752 3796 28812 3802
rect 30782 3796 30842 3802
rect 32822 3798 32882 3804
rect 34312 3798 34372 3804
rect -10744 3789 -10642 3794
rect -6568 3791 -6474 3796
rect -10748 3697 -10739 3789
rect -10647 3697 -10638 3789
rect -6572 3707 -6563 3791
rect -6479 3707 -6470 3791
rect -10744 3649 -10642 3697
rect -10744 3547 -8631 3649
rect -8733 3485 -8631 3547
rect -6568 3639 -6474 3707
rect -6568 3545 -4455 3639
rect -8733 3374 -8631 3383
rect -4549 3473 -4455 3545
rect -4549 3370 -4455 3379
rect 10572 3342 10632 3348
rect 2420 3282 2426 3342
rect 2486 3282 4462 3342
rect 4522 3282 6494 3342
rect 6554 3282 8528 3342
rect 8588 3282 10572 3342
rect 10572 3276 10632 3282
rect 1412 3234 1472 3240
rect 3448 3234 3508 3240
rect 5484 3234 5544 3240
rect 7518 3234 7578 3240
rect 9554 3234 9614 3240
rect 1472 3174 3448 3234
rect 3508 3174 5484 3234
rect 5544 3174 7518 3234
rect 7578 3174 9554 3234
rect 1412 3168 1472 3174
rect 3448 3168 3508 3174
rect 5484 3168 5544 3174
rect 7518 3168 7578 3174
rect 9554 3168 9614 3174
rect 1906 3122 1966 3128
rect 2930 3122 2990 3128
rect 3962 3122 4022 3128
rect 4962 3122 5022 3128
rect 5982 3122 6042 3128
rect 7002 3122 7062 3128
rect 9026 3122 9086 3128
rect 11848 3122 11908 3128
rect 1966 3062 2930 3122
rect 2990 3062 3962 3122
rect 4022 3062 4962 3122
rect 5022 3062 5982 3122
rect 6042 3062 7002 3122
rect 7062 3062 8012 3122
rect 8072 3062 9026 3122
rect 9086 3062 10044 3122
rect 10104 3062 11848 3122
rect 1906 3056 1966 3062
rect 2930 3056 2990 3062
rect 3962 3056 4022 3062
rect 4962 3056 5022 3062
rect 5982 3056 6042 3062
rect 7002 3056 7062 3062
rect 9026 3056 9086 3062
rect 11848 3056 11908 3062
rect 13248 2946 13308 2952
rect 22636 2946 22696 2952
rect 24678 2946 24738 2952
rect 26714 2946 26774 2952
rect 13308 2886 22636 2946
rect 22696 2886 24678 2946
rect 24738 2886 26714 2946
rect 13248 2880 13308 2886
rect 22636 2880 22696 2886
rect 24678 2880 24738 2886
rect 26714 2880 26774 2886
rect 29768 2946 29828 2952
rect 31800 2946 31860 2952
rect 33946 2946 34006 2952
rect 29828 2886 31800 2946
rect 31860 2886 33946 2946
rect 29768 2880 29828 2886
rect 31800 2880 31860 2886
rect 33946 2880 34006 2886
rect 17052 2832 17112 2838
rect 22132 2832 22192 2838
rect 13142 2820 13202 2826
rect 16532 2820 16592 2826
rect 13202 2760 16532 2820
rect 17112 2772 22132 2832
rect 17052 2766 17112 2772
rect 22132 2766 22192 2772
rect 27220 2836 27280 2842
rect 32320 2836 32380 2842
rect 27280 2776 32320 2836
rect 27220 2770 27280 2776
rect 32320 2770 32380 2776
rect 33328 2836 33388 2842
rect 34562 2836 34622 2842
rect 33388 2776 34562 2836
rect 33328 2770 33388 2776
rect 34562 2770 34622 2776
rect 13142 2754 13202 2760
rect 16532 2754 16592 2760
rect 15514 2718 15574 2724
rect 17550 2718 17610 2724
rect 18570 2718 18630 2724
rect 19586 2718 19646 2724
rect 20606 2718 20666 2724
rect 21624 2718 21684 2724
rect 23654 2718 23714 2724
rect 25692 2718 25752 2724
rect 27728 2718 27788 2724
rect 28750 2718 28810 2724
rect 29770 2718 29830 2724
rect 30784 2718 30844 2724
rect 31806 2718 31866 2724
rect 15574 2658 17550 2718
rect 17610 2658 18570 2718
rect 18630 2658 19586 2718
rect 19646 2658 20606 2718
rect 20666 2658 21624 2718
rect 21684 2658 23654 2718
rect 23714 2658 25692 2718
rect 25752 2658 27728 2718
rect 27788 2658 28750 2718
rect 28810 2658 29770 2718
rect 29830 2658 30784 2718
rect 30844 2658 31806 2718
rect 15514 2652 15574 2658
rect 17550 2652 17610 2658
rect 18570 2652 18630 2658
rect 19586 2652 19646 2658
rect 20606 2652 20666 2658
rect 21624 2652 21684 2658
rect 23654 2652 23714 2658
rect 25692 2652 25752 2658
rect 27728 2652 27788 2658
rect 28750 2652 28810 2658
rect 29770 2652 29830 2658
rect 30784 2652 30844 2658
rect 31806 2652 31866 2658
rect 16532 2614 16592 2620
rect 21468 2614 21528 2620
rect 27874 2614 27934 2620
rect 30784 2614 30844 2620
rect 33966 2614 34026 2620
rect 16592 2554 21468 2614
rect 21528 2554 27874 2614
rect 27934 2554 30784 2614
rect 30844 2554 33966 2614
rect 16532 2548 16592 2554
rect 21468 2548 21528 2554
rect 27874 2548 27934 2554
rect 30784 2548 30844 2554
rect 33966 2548 34026 2554
rect 250 2160 310 2166
rect 2920 2160 2980 2166
rect 3952 2160 4012 2166
rect 7012 2160 7072 2166
rect 8008 2160 8068 2166
rect 310 2100 2920 2160
rect 2980 2100 3952 2160
rect 4012 2100 7012 2160
rect 7072 2100 8008 2160
rect 250 2094 310 2100
rect 2920 2094 2980 2100
rect 3952 2094 4012 2100
rect 7012 2094 7072 2100
rect 8008 2094 8068 2100
rect 5486 2030 5546 2036
rect 9546 2030 9606 2036
rect 11728 2030 11788 2036
rect 1400 1970 1406 2030
rect 1466 1970 5486 2030
rect 5546 1970 9546 2030
rect 9606 1970 11728 2030
rect 5486 1964 5546 1970
rect 9546 1964 9606 1970
rect 11728 1964 11788 1970
rect 13360 1716 13420 1722
rect 16530 1716 16590 1722
rect 13420 1656 16530 1716
rect 13360 1650 13420 1656
rect 16530 1650 16590 1656
rect 20760 1718 20820 1724
rect 22638 1718 22698 1724
rect 24676 1718 24736 1724
rect 26546 1718 26606 1724
rect 32822 1718 32882 1724
rect 20820 1658 22638 1718
rect 22698 1658 24676 1718
rect 24736 1658 26546 1718
rect 26606 1658 32822 1718
rect 20760 1652 20820 1658
rect 22638 1652 22698 1658
rect 24676 1652 24736 1658
rect 26546 1652 26606 1658
rect 32822 1652 32882 1658
rect 13032 1612 13092 1618
rect 14496 1612 14556 1618
rect 16536 1612 16596 1618
rect 18566 1612 18626 1618
rect 20606 1612 20666 1618
rect 22642 1612 22702 1618
rect 24678 1612 24738 1618
rect 26712 1612 26772 1618
rect 28752 1612 28812 1618
rect 30782 1612 30842 1618
rect 32822 1612 32882 1618
rect 34674 1612 34734 1618
rect 13092 1552 14496 1612
rect 14556 1552 16536 1612
rect 16596 1552 18566 1612
rect 18626 1552 20606 1612
rect 20666 1552 22642 1612
rect 22702 1552 24678 1612
rect 24738 1552 26712 1612
rect 26772 1552 28752 1612
rect 28812 1552 30782 1612
rect 30842 1552 32822 1612
rect 32882 1552 34674 1612
rect 13032 1546 13092 1552
rect 14496 1546 14556 1552
rect 16536 1546 16596 1552
rect 18566 1546 18626 1552
rect 20606 1546 20666 1552
rect 22642 1546 22702 1552
rect 24678 1546 24738 1552
rect 26712 1546 26772 1552
rect 28752 1546 28812 1552
rect 30782 1546 30842 1552
rect 32822 1546 32882 1552
rect 34674 1546 34734 1552
rect 15004 1506 15064 1512
rect 16024 1506 16084 1512
rect 17048 1506 17108 1512
rect 18066 1506 18126 1512
rect 19080 1506 19140 1512
rect 20112 1506 20172 1512
rect 21124 1506 21184 1512
rect 22132 1506 22192 1512
rect 23150 1506 23210 1512
rect 24176 1506 24236 1512
rect 25178 1506 25238 1512
rect 26198 1506 26258 1512
rect 27218 1506 27278 1512
rect 28244 1506 28304 1512
rect 29262 1506 29322 1512
rect 30276 1506 30336 1512
rect 31290 1506 31350 1512
rect 32312 1506 32372 1512
rect 15064 1446 16024 1506
rect 16084 1446 17048 1506
rect 17108 1446 18066 1506
rect 18126 1446 19080 1506
rect 19140 1446 20112 1506
rect 20172 1446 21124 1506
rect 21184 1446 22132 1506
rect 22192 1446 23150 1506
rect 23210 1446 24176 1506
rect 24236 1446 25178 1506
rect 25238 1446 26198 1506
rect 26258 1446 27218 1506
rect 27278 1446 28244 1506
rect 28304 1446 29262 1506
rect 29322 1446 30276 1506
rect 30336 1446 31290 1506
rect 31350 1446 32312 1506
rect 15004 1440 15064 1446
rect 16024 1440 16084 1446
rect 17048 1440 17108 1446
rect 18066 1440 18126 1446
rect 19080 1440 19140 1446
rect 20112 1440 20172 1446
rect 21124 1440 21184 1446
rect 22132 1440 22192 1446
rect 23150 1440 23210 1446
rect 24176 1440 24236 1446
rect 25178 1440 25238 1446
rect 26198 1440 26258 1446
rect 27218 1440 27278 1446
rect 28244 1440 28304 1446
rect 29262 1440 29322 1446
rect 30276 1440 30336 1446
rect 31290 1440 31350 1446
rect 32312 1440 32372 1446
rect 15516 1396 15576 1402
rect 17552 1396 17612 1402
rect 19590 1396 19650 1402
rect 21628 1396 21688 1402
rect 23664 1396 23724 1402
rect 25700 1396 25760 1402
rect 27732 1396 27792 1402
rect 29764 1396 29824 1402
rect 31804 1396 31864 1402
rect 15576 1336 17552 1396
rect 17612 1336 19590 1396
rect 19650 1336 21628 1396
rect 21688 1336 23664 1396
rect 23724 1336 25700 1396
rect 25760 1336 27732 1396
rect 27792 1336 29764 1396
rect 29824 1336 31804 1396
rect 15516 1330 15576 1336
rect 17552 1330 17612 1336
rect 19590 1330 19650 1336
rect 21628 1330 21688 1336
rect 23664 1330 23724 1336
rect 25700 1330 25760 1336
rect 27732 1330 27792 1336
rect 29764 1330 29824 1336
rect 31804 1330 31864 1336
rect 2884 664 2944 670
rect 4922 664 4982 670
rect 6958 664 7018 670
rect 8994 664 9054 670
rect 2944 604 4922 664
rect 4982 604 6958 664
rect 7018 604 8994 664
rect 2884 598 2944 604
rect 4922 598 4982 604
rect 6958 598 7018 604
rect 8994 598 9054 604
rect 3902 552 3962 558
rect 7976 552 8036 558
rect 11982 552 12042 558
rect 3962 492 7976 552
rect 8036 492 11982 552
rect 3902 486 3962 492
rect 7976 486 8036 492
rect 11982 486 12042 492
rect 13360 474 13420 480
rect 14496 474 14556 480
rect 18566 474 18626 480
rect 28746 474 28806 480
rect 33966 474 34026 480
rect 13420 414 14496 474
rect 14556 414 18566 474
rect 18626 414 28746 474
rect 28806 414 33966 474
rect 13360 408 13420 414
rect 14496 408 14556 414
rect 18566 408 18626 414
rect 28746 408 28806 414
rect 33966 408 34026 414
rect 15008 366 15068 372
rect 23152 366 23212 372
rect 15068 306 16022 366
rect 16082 306 17044 366
rect 17104 306 18058 366
rect 18118 306 19084 366
rect 19144 306 20096 366
rect 20156 306 21132 366
rect 21192 306 22138 366
rect 22198 306 23152 366
rect 23212 306 24168 366
rect 24228 306 25176 366
rect 25236 306 26192 366
rect 26252 306 27216 366
rect 27276 306 28238 366
rect 28298 306 29260 366
rect 29320 306 30278 366
rect 30338 306 31292 366
rect 31352 306 32316 366
rect 32376 306 32382 366
rect 15008 300 15068 306
rect 23152 300 23212 306
rect 2794 64 34880 110
rect 2794 -90 2840 64
rect 34840 -90 34880 64
rect 2794 -136 34880 -90
rect -1304 -276 -704 -266
rect -1304 -586 -704 -576
rect 35128 -276 35728 -266
rect 35128 -586 35728 -576
<< via2 >>
rect 11396 30456 11996 30756
rect 35028 30456 35628 30756
rect -4458 30228 -4398 30288
rect 14973 30160 31758 30374
rect -13288 15502 -13228 15562
rect -9666 15502 -9606 15562
rect -2718 15870 8046 16162
rect 8046 15870 8134 16162
rect -12486 15353 -12426 15413
rect -9850 15353 -9790 15413
rect 13231 15501 13321 15591
rect -13105 14481 -13015 14571
rect -9874 14476 -9774 14576
rect -13499 14259 -13409 14349
rect -9686 14254 -9586 14354
rect -11017 10929 -10937 11009
rect -6659 10925 -6583 11001
rect -8685 10613 -8595 10703
rect -4457 10603 -4371 10689
rect -1842 6458 -1782 6518
rect -1566 5496 -1506 5556
rect -10739 3697 -10647 3789
rect -6563 3707 -6479 3791
rect -8733 3383 -8631 3485
rect -4549 3379 -4455 3473
rect 2840 -90 34840 64
rect -1304 -576 -704 -276
rect 35128 -576 35728 -276
<< metal3 >>
rect 11386 30756 12006 30761
rect 11386 30456 11396 30756
rect 11996 30456 12006 30756
rect 11386 30451 12006 30456
rect 35018 30756 35638 30761
rect 35018 30456 35028 30756
rect 35628 30456 35638 30756
rect 35018 30451 35638 30456
rect 14910 30374 31790 30406
rect -4486 30293 -4350 30322
rect -4486 30229 -4463 30293
rect -4393 30229 -4350 30293
rect -4486 30228 -4458 30229
rect -4398 30228 -4350 30229
rect -4486 30192 -4350 30228
rect 14910 30160 14973 30374
rect 31758 30160 31790 30374
rect 14910 30140 31790 30160
rect 14910 30138 19264 30140
rect -4256 29480 10784 29626
rect -4256 29470 9938 29480
rect -4256 28780 -4104 29470
rect -3408 28782 9938 29470
rect 10628 28782 10784 29480
rect -3408 28780 10784 28782
rect -4256 28450 10784 28780
rect -4256 15788 -3074 28450
rect -2786 17250 9120 28190
rect 9484 17250 10784 28450
rect -2786 16162 10784 17250
rect 8134 15870 10784 16162
rect 8046 15788 10784 15870
rect -13310 15562 -13210 15584
rect -13310 15502 -13288 15562
rect -13228 15502 -13210 15562
rect -13504 14349 -13404 14354
rect -13504 14259 -13499 14349
rect -13409 14259 -13404 14349
rect -13504 3497 -13404 14259
rect -13310 5903 -13210 15502
rect -9686 15562 -9586 15580
rect -9686 15502 -9666 15562
rect -9606 15502 -9586 15562
rect -12510 15413 -12410 15434
rect -12510 15353 -12486 15413
rect -12426 15353 -12410 15413
rect -12510 14688 -12410 15353
rect -12510 14582 -12410 14588
rect -9874 15413 -9774 15436
rect -9874 15353 -9850 15413
rect -9790 15353 -9774 15413
rect -9874 14581 -9774 15353
rect -9879 14576 -9769 14581
rect -13110 14571 -13010 14576
rect -13110 14481 -13105 14571
rect -13015 14481 -13010 14571
rect -13110 10725 -13010 14481
rect -9879 14476 -9874 14576
rect -9774 14476 -9769 14576
rect -9879 14471 -9769 14476
rect -9686 14359 -9586 15502
rect -4256 15562 10784 15788
rect 13227 15596 13325 15601
rect 13226 15595 13326 15596
rect -4256 15462 9286 15562
rect 13226 15497 13227 15595
rect 13325 15497 13326 15595
rect 13226 15496 13326 15497
rect 13227 15491 13325 15496
rect -4256 14780 -4102 15462
rect -3768 14780 9286 15462
rect -4256 14624 9286 14780
rect 10952 14470 11052 14476
rect -1600 14370 10952 14470
rect -9691 14354 -9581 14359
rect -9691 14254 -9686 14354
rect -9586 14254 -9581 14354
rect -9691 14249 -9581 14254
rect -11124 14114 -10954 14120
rect -12012 14010 -11124 14012
rect -12572 13944 -11124 14010
rect -8772 14118 -8612 14124
rect -10954 13958 -8772 14012
rect -6398 14122 -6256 14128
rect -8612 13980 -6398 14012
rect -4024 14106 -3862 14112
rect -6256 13980 -4024 14012
rect -8612 13958 -4024 13980
rect -10954 13944 -4024 13958
rect -3862 14010 -2653 14012
rect -3862 13944 -2610 14010
rect -12572 13408 -2610 13944
rect -12572 11918 -11971 13408
rect -10026 13056 -7214 13156
rect -10026 12776 -9896 13056
rect -7314 12776 -7214 13056
rect -12700 11820 -12694 11918
rect -12596 11820 -11971 11918
rect -13115 10627 -13109 10725
rect -13011 10627 -13005 10725
rect -13110 10626 -13010 10627
rect -12572 9826 -11971 11820
rect -11684 11009 -9896 12776
rect -11684 10976 -11017 11009
rect -11022 10929 -11017 10976
rect -10937 10976 -9896 11009
rect -9644 11021 -7856 12776
rect -9644 10976 -9331 11021
rect -10937 10929 -10932 10976
rect -11022 10924 -10932 10929
rect -9337 10923 -9331 10976
rect -9233 10976 -7856 11021
rect -7444 11001 -5656 12776
rect -7444 10976 -6659 11001
rect -9233 10923 -9227 10976
rect -6664 10925 -6659 10976
rect -6583 10976 -5656 11001
rect -5404 11029 -3616 12776
rect -5404 10976 -5191 11029
rect -6583 10925 -6578 10976
rect -5197 10931 -5191 10976
rect -5093 10976 -3616 11029
rect -3213 11908 -2610 13408
rect -1858 12903 -1758 12904
rect -1863 12805 -1857 12903
rect -1759 12805 -1753 12903
rect -3213 11786 -2562 11908
rect -2440 11786 -2434 11908
rect -5093 10931 -5087 10976
rect -5192 10930 -5092 10931
rect -9332 10922 -9232 10923
rect -6664 10920 -6578 10925
rect -8101 10882 -8003 10887
rect -7570 10882 -7470 10888
rect -8102 10881 -7570 10882
rect -8102 10783 -8101 10881
rect -8003 10783 -7570 10881
rect -8102 10782 -7570 10783
rect -3901 10880 -3803 10885
rect -3400 10880 -3300 10886
rect -8101 10777 -8003 10782
rect -7570 10776 -7470 10782
rect -3902 10879 -3400 10880
rect -3902 10781 -3901 10879
rect -3803 10781 -3400 10879
rect -3902 10780 -3400 10781
rect -3901 10775 -3803 10780
rect -3400 10774 -3300 10780
rect -10156 10725 -10056 10726
rect -5956 10725 -5856 10726
rect -10161 10676 -10155 10725
rect -12678 9708 -12672 9826
rect -12554 9708 -11971 9826
rect -13100 8615 -13000 8616
rect -13105 8517 -13099 8615
rect -13001 8517 -12995 8615
rect -13315 5805 -13309 5903
rect -13211 5805 -13205 5903
rect -13310 5804 -13210 5805
rect -13509 3399 -13503 3497
rect -13405 3399 -13399 3497
rect -13504 3398 -13404 3399
rect -13100 1627 -13000 8517
rect -12572 8256 -11971 9708
rect -11684 10627 -10155 10676
rect -10057 10676 -10051 10725
rect -8690 10703 -8590 10708
rect -8690 10676 -8685 10703
rect -10057 10627 -9896 10676
rect -11684 8876 -9896 10627
rect -9644 10613 -8685 10676
rect -8595 10676 -8590 10703
rect -5961 10676 -5955 10725
rect -8595 10613 -7856 10676
rect -9644 8876 -7856 10613
rect -7444 10627 -5955 10676
rect -5857 10676 -5851 10725
rect -4462 10689 -4366 10694
rect -4462 10676 -4457 10689
rect -5857 10627 -5656 10676
rect -7444 8876 -5656 10627
rect -5404 10603 -4457 10676
rect -4371 10676 -4366 10689
rect -4371 10603 -3616 10676
rect -5404 8876 -3616 10603
rect -3213 9850 -2610 11786
rect -3213 9742 -2534 9850
rect -2426 9742 -2420 9850
rect -10102 8616 -10002 8876
rect -7192 8616 -7092 8876
rect -10510 8516 -10504 8616
rect -10404 8516 -7092 8616
rect -3213 8256 -2610 9742
rect -12572 7654 -2610 8256
rect -12572 7652 -2956 7654
rect -11068 7570 -10886 7652
rect -11068 7402 -11061 7570
rect -10893 7402 -10886 7570
rect -8768 7570 -8586 7652
rect -8768 7402 -8761 7570
rect -8593 7402 -8586 7570
rect -6468 7570 -6286 7652
rect -6468 7402 -6461 7570
rect -6293 7402 -6286 7570
rect -4048 7570 -3866 7652
rect -4048 7402 -4041 7570
rect -3873 7402 -3866 7570
rect -11062 7401 -10892 7402
rect -8762 7401 -8592 7402
rect -6462 7401 -6292 7402
rect -4042 7401 -3872 7402
rect -11062 6884 -10892 6890
rect -11950 6780 -11062 6782
rect -12309 6778 -11062 6780
rect -12509 6714 -11062 6778
rect -8762 6884 -8592 6890
rect -10892 6714 -8762 6782
rect -6462 6884 -6292 6890
rect -8592 6714 -6462 6782
rect -4042 6884 -3872 6890
rect -6292 6714 -4042 6782
rect -3872 6778 -2591 6782
rect -3872 6714 -2548 6778
rect -12509 6178 -2548 6714
rect -12509 4688 -11909 6178
rect -11530 5804 -11524 5904
rect -11424 5804 -7198 5904
rect -10006 5546 -9906 5804
rect -7298 5546 -7198 5804
rect -12638 4590 -12632 4688
rect -12534 4590 -11909 4688
rect -12509 2596 -11909 4590
rect -11622 3789 -9834 5546
rect -11622 3746 -10739 3789
rect -10744 3697 -10739 3746
rect -10647 3746 -9834 3789
rect -9582 3797 -7794 5546
rect -9582 3746 -9303 3797
rect -10647 3697 -10642 3746
rect -9309 3699 -9303 3746
rect -9205 3746 -7794 3797
rect -7382 3791 -5594 5546
rect -7382 3746 -6563 3791
rect -9205 3699 -9199 3746
rect -6568 3707 -6563 3746
rect -6479 3746 -5594 3791
rect -5342 3801 -3554 5546
rect -5342 3746 -5083 3801
rect -6479 3707 -6474 3746
rect -6568 3702 -6474 3707
rect -5089 3703 -5083 3746
rect -4985 3746 -3554 3801
rect -3151 4678 -2548 6178
rect -1858 6518 -1758 12805
rect -1600 8863 -1500 14370
rect 10952 14364 11052 14370
rect -1605 8765 -1599 8863
rect -1501 8765 -1495 8863
rect -1600 8764 -1500 8765
rect -1858 6458 -1842 6518
rect -1782 6458 -1758 6518
rect -1858 5665 -1758 6458
rect -1863 5567 -1857 5665
rect -1759 5567 -1753 5665
rect -1858 5566 -1758 5567
rect -1586 5556 -1486 5594
rect -1586 5496 -1566 5556
rect -1506 5496 -1486 5556
rect -3151 4556 -2500 4678
rect -2378 4556 -2372 4678
rect -4985 3703 -4979 3746
rect -5084 3702 -4984 3703
rect -9304 3698 -9204 3699
rect -10744 3692 -10642 3697
rect -8085 3644 -7987 3649
rect -7554 3644 -7454 3650
rect -3845 3644 -3747 3649
rect -3344 3644 -3244 3650
rect -8086 3643 -7554 3644
rect -8086 3545 -8085 3643
rect -7987 3545 -7554 3643
rect -8086 3544 -7554 3545
rect -3846 3643 -3344 3644
rect -3846 3545 -3845 3643
rect -3747 3545 -3344 3643
rect -3846 3544 -3344 3545
rect -8085 3539 -7987 3544
rect -7554 3538 -7454 3544
rect -3845 3539 -3747 3544
rect -3344 3538 -3244 3544
rect -5940 3501 -5840 3502
rect -10180 3497 -10080 3498
rect -10185 3446 -10179 3497
rect -12616 2478 -12610 2596
rect -12492 2478 -11909 2596
rect -13103 1529 -13097 1627
rect -12999 1529 -12993 1627
rect -13100 1528 -13000 1529
rect -12509 1028 -11909 2478
rect -11622 3399 -10179 3446
rect -10081 3446 -10075 3497
rect -8738 3485 -8626 3490
rect -8738 3446 -8733 3485
rect -10081 3399 -9834 3446
rect -11622 1646 -9834 3399
rect -9582 3383 -8733 3446
rect -8631 3446 -8626 3485
rect -5945 3446 -5939 3501
rect -8631 3383 -7794 3446
rect -9582 1646 -7794 3383
rect -7382 3403 -5939 3446
rect -5841 3446 -5835 3501
rect -4554 3473 -4450 3478
rect -4554 3446 -4549 3473
rect -5841 3403 -5594 3446
rect -7382 1646 -5594 3403
rect -5342 3379 -4549 3446
rect -4455 3446 -4450 3473
rect -4455 3379 -3554 3446
rect -5342 1646 -3554 3379
rect -3151 2620 -2548 4556
rect -3151 2512 -2472 2620
rect -2364 2512 -2358 2620
rect -10126 1378 -10026 1646
rect -7176 1378 -7076 1646
rect -10126 1278 -7076 1378
rect -3151 1028 -2548 2512
rect -1586 1625 -1486 5496
rect -1591 1527 -1585 1625
rect -1487 1527 -1481 1625
rect -1586 1526 -1486 1527
rect -12509 484 -2548 1028
rect -12509 422 -11094 484
rect -10918 422 -8682 484
rect -11094 302 -10918 308
rect -8506 422 -6362 484
rect -8682 302 -8506 308
rect -6186 422 -3962 484
rect -6362 302 -6186 308
rect -3786 424 -2548 484
rect -3786 422 -3061 424
rect -3962 302 -3786 308
rect 2794 64 34880 110
rect 2794 -90 2840 64
rect 34840 -90 34880 64
rect 2794 -136 34880 -90
rect -1314 -276 -694 -271
rect -1314 -576 -1304 -276
rect -704 -576 -694 -276
rect -1314 -581 -694 -576
rect 35118 -276 35738 -271
rect 35118 -576 35128 -276
rect 35728 -576 35738 -276
rect 35118 -581 35738 -576
<< via3 >>
rect 11396 30456 11996 30756
rect 35028 30456 35628 30756
rect -4463 30288 -4393 30293
rect -4463 30229 -4458 30288
rect -4458 30229 -4398 30288
rect -4398 30229 -4393 30288
rect 14973 30160 31758 30374
rect -4104 28780 -3408 29470
rect 9938 28782 10628 29480
rect -3074 28190 9484 28450
rect -3074 16162 -2786 28190
rect 9120 17250 9484 28190
rect -3074 15870 -2718 16162
rect -2718 15870 8046 16162
rect -3074 15788 8046 15870
rect -12510 14588 -12410 14688
rect 13227 15591 13325 15595
rect 13227 15501 13231 15591
rect 13231 15501 13321 15591
rect 13321 15501 13325 15591
rect 13227 15497 13325 15501
rect -4102 14780 -3768 15462
rect 10952 14370 11052 14470
rect -11124 13944 -10954 14114
rect -8772 13958 -8612 14118
rect -6398 13980 -6256 14122
rect -4024 13944 -3862 14106
rect -12694 11820 -12596 11918
rect -13109 10627 -13011 10725
rect -9331 10923 -9233 11021
rect -5191 10931 -5093 11029
rect -1857 12805 -1759 12903
rect -2562 11786 -2440 11908
rect -8101 10783 -8003 10881
rect -7570 10782 -7470 10882
rect -3901 10781 -3803 10879
rect -3400 10780 -3300 10880
rect -12672 9708 -12554 9826
rect -13099 8517 -13001 8615
rect -13309 5805 -13211 5903
rect -13503 3399 -13405 3497
rect -10155 10627 -10057 10725
rect -5955 10627 -5857 10725
rect -2534 9742 -2426 9850
rect -10504 8516 -10404 8616
rect -11061 7402 -10893 7570
rect -8761 7402 -8593 7570
rect -6461 7402 -6293 7570
rect -4041 7402 -3873 7570
rect -11062 6714 -10892 6884
rect -8762 6714 -8592 6884
rect -6462 6714 -6292 6884
rect -4042 6714 -3872 6884
rect -11524 5804 -11424 5904
rect -12632 4590 -12534 4688
rect -9303 3699 -9205 3797
rect -5083 3703 -4985 3801
rect -1599 8765 -1501 8863
rect -1857 5567 -1759 5665
rect -2500 4556 -2378 4678
rect -8085 3545 -7987 3643
rect -7554 3544 -7454 3644
rect -3845 3545 -3747 3643
rect -3344 3544 -3244 3644
rect -12610 2478 -12492 2596
rect -13097 1529 -12999 1627
rect -10179 3399 -10081 3497
rect -5939 3403 -5841 3501
rect -2472 2512 -2364 2620
rect -1585 1527 -1487 1625
rect -11094 308 -10918 484
rect -8682 308 -8506 484
rect -6362 308 -6186 484
rect -3962 308 -3786 484
rect 2840 -90 34840 64
rect -1304 -576 -704 -276
rect 35128 -576 35728 -276
<< mimcap >>
rect -3070 29476 3130 29526
rect -3070 29176 2780 29476
rect 3080 29176 3130 29476
rect -3070 29126 3130 29176
rect 3330 29476 9530 29526
rect 3330 29176 9180 29476
rect 9480 29176 9530 29476
rect 3330 29126 9530 29176
rect -4156 28394 -3356 28444
rect -4156 22694 -3706 28394
rect -3406 22694 -3356 28394
rect 9888 28394 10688 28444
rect -2216 27476 2984 27526
rect -2216 22776 2634 27476
rect 2934 22776 2984 27476
rect -2216 22726 2984 22776
rect 3384 27476 8584 27526
rect 3384 22776 8234 27476
rect 8534 22776 8584 27476
rect 3384 22726 8584 22776
rect -4156 22644 -3356 22694
rect 9888 22694 10338 28394
rect 10638 22694 10688 28394
rect 9888 22644 10688 22694
rect -4156 21902 -3356 21952
rect -4156 16202 -3706 21902
rect -3406 16202 -3356 21902
rect -2216 21876 2984 21926
rect -2216 17176 2634 21876
rect 2934 17176 2984 21876
rect -2216 17126 2984 17176
rect 3384 21876 8584 21926
rect 3384 17176 8234 21876
rect 8534 17176 8584 21876
rect 3384 17126 8584 17176
rect 9888 21902 10688 21952
rect -4156 16152 -3356 16202
rect 9888 16202 10338 21902
rect 10638 16202 10688 21902
rect 9888 16152 10688 16202
rect -3570 15476 2630 15526
rect -3570 15176 2280 15476
rect 2580 15176 2630 15476
rect -3570 15126 2630 15176
rect 2830 15476 9030 15526
rect 2830 15176 8680 15476
rect 8980 15176 9030 15476
rect 2830 15126 9030 15176
rect -12289 13870 -9889 13910
rect -12289 13550 -12249 13870
rect -9929 13550 -9889 13870
rect -12289 13510 -9889 13550
rect -9506 13870 -7906 13910
rect -9506 13550 -9466 13870
rect -7946 13550 -7906 13870
rect -9506 13510 -7906 13550
rect -7118 13872 -5518 13912
rect -7118 13552 -7078 13872
rect -5558 13552 -5518 13872
rect -7118 13512 -5518 13552
rect -5135 13872 -2735 13912
rect -5135 13552 -5095 13872
rect -2775 13552 -2735 13872
rect -5135 13512 -2735 13552
rect -12470 12636 -12070 12676
rect -12470 11116 -12430 12636
rect -12110 11116 -12070 12636
rect -12470 11076 -12070 11116
rect -11584 12636 -9984 12676
rect -11584 11116 -11544 12636
rect -10024 11116 -9984 12636
rect -11584 11076 -9984 11116
rect -9544 12636 -7944 12676
rect -9544 11116 -9504 12636
rect -7984 11116 -7944 12636
rect -9544 11076 -7944 11116
rect -7344 12636 -5744 12676
rect -7344 11116 -7304 12636
rect -5784 11116 -5744 12636
rect -7344 11076 -5744 11116
rect -5304 12636 -3704 12676
rect -5304 11116 -5264 12636
rect -3744 11116 -3704 12636
rect -5304 11076 -3704 11116
rect -3114 12638 -2714 12678
rect -3114 11118 -3074 12638
rect -2754 11118 -2714 12638
rect -3114 11078 -2714 11118
rect -12470 10532 -12070 10572
rect -12470 9012 -12430 10532
rect -12110 9012 -12070 10532
rect -12470 8972 -12070 9012
rect -11584 10536 -9984 10576
rect -11584 9016 -11544 10536
rect -10024 9016 -9984 10536
rect -11584 8976 -9984 9016
rect -9544 10536 -7944 10576
rect -9544 9016 -9504 10536
rect -7984 9016 -7944 10536
rect -9544 8976 -7944 9016
rect -7344 10536 -5744 10576
rect -7344 9016 -7304 10536
rect -5784 9016 -5744 10536
rect -7344 8976 -5744 9016
rect -5304 10536 -3704 10576
rect -5304 9016 -5264 10536
rect -3744 9016 -3704 10536
rect -5304 8976 -3704 9016
rect -3114 10534 -2714 10574
rect -3114 9014 -3074 10534
rect -2754 9014 -2714 10534
rect -3114 8974 -2714 9014
rect -12289 8114 -9889 8154
rect -12289 7794 -12249 8114
rect -9929 7794 -9889 8114
rect -12289 7754 -9889 7794
rect -9506 8114 -7906 8154
rect -9506 7794 -9466 8114
rect -7946 7794 -7906 8114
rect -9506 7754 -7906 7794
rect -7118 8116 -5518 8156
rect -7118 7796 -7078 8116
rect -5558 7796 -5518 8116
rect -7118 7756 -5518 7796
rect -5135 8116 -2735 8156
rect -5135 7796 -5095 8116
rect -2775 7796 -2735 8116
rect -5135 7756 -2735 7796
rect -12227 6640 -9827 6680
rect -12227 6320 -12187 6640
rect -9867 6320 -9827 6640
rect -12227 6280 -9827 6320
rect -9444 6640 -7844 6680
rect -9444 6320 -9404 6640
rect -7884 6320 -7844 6640
rect -9444 6280 -7844 6320
rect -7056 6642 -5456 6682
rect -7056 6322 -7016 6642
rect -5496 6322 -5456 6642
rect -7056 6282 -5456 6322
rect -5073 6642 -2673 6682
rect -5073 6322 -5033 6642
rect -2713 6322 -2673 6642
rect -5073 6282 -2673 6322
rect -12408 5406 -12008 5446
rect -12408 3886 -12368 5406
rect -12048 3886 -12008 5406
rect -12408 3846 -12008 3886
rect -11522 5406 -9922 5446
rect -11522 3886 -11482 5406
rect -9962 3886 -9922 5406
rect -11522 3846 -9922 3886
rect -9482 5406 -7882 5446
rect -9482 3886 -9442 5406
rect -7922 3886 -7882 5406
rect -9482 3846 -7882 3886
rect -7282 5406 -5682 5446
rect -7282 3886 -7242 5406
rect -5722 3886 -5682 5406
rect -7282 3846 -5682 3886
rect -5242 5406 -3642 5446
rect -5242 3886 -5202 5406
rect -3682 3886 -3642 5406
rect -5242 3846 -3642 3886
rect -3052 5408 -2652 5448
rect -3052 3888 -3012 5408
rect -2692 3888 -2652 5408
rect -3052 3848 -2652 3888
rect -12408 3302 -12008 3342
rect -12408 1782 -12368 3302
rect -12048 1782 -12008 3302
rect -12408 1742 -12008 1782
rect -11522 3306 -9922 3346
rect -11522 1786 -11482 3306
rect -9962 1786 -9922 3306
rect -11522 1746 -9922 1786
rect -9482 3306 -7882 3346
rect -9482 1786 -9442 3306
rect -7922 1786 -7882 3306
rect -9482 1746 -7882 1786
rect -7282 3306 -5682 3346
rect -7282 1786 -7242 3306
rect -5722 1786 -5682 3306
rect -7282 1746 -5682 1786
rect -5242 3306 -3642 3346
rect -5242 1786 -5202 3306
rect -3682 1786 -3642 3306
rect -5242 1746 -3642 1786
rect -3052 3304 -2652 3344
rect -3052 1784 -3012 3304
rect -2692 1784 -2652 3304
rect -3052 1744 -2652 1784
rect -12227 884 -9827 924
rect -12227 564 -12187 884
rect -9867 564 -9827 884
rect -12227 524 -9827 564
rect -9444 884 -7844 924
rect -9444 564 -9404 884
rect -7884 564 -7844 884
rect -9444 524 -7844 564
rect -7056 886 -5456 926
rect -7056 566 -7016 886
rect -5496 566 -5456 886
rect -7056 526 -5456 566
rect -5073 886 -2673 926
rect -5073 566 -5033 886
rect -2713 566 -2673 886
rect -5073 526 -2673 566
<< mimcapcontact >>
rect 2780 29176 3080 29476
rect 9180 29176 9480 29476
rect -3706 22694 -3406 28394
rect 2634 22776 2934 27476
rect 8234 22776 8534 27476
rect 10338 22694 10638 28394
rect -3706 16202 -3406 21902
rect 2634 17176 2934 21876
rect 8234 17176 8534 21876
rect 10338 16202 10638 21902
rect 2280 15176 2580 15476
rect 8680 15176 8980 15476
rect -12249 13550 -9929 13870
rect -9466 13550 -7946 13870
rect -7078 13552 -5558 13872
rect -5095 13552 -2775 13872
rect -12430 11116 -12110 12636
rect -11544 11116 -10024 12636
rect -9504 11116 -7984 12636
rect -7304 11116 -5784 12636
rect -5264 11116 -3744 12636
rect -3074 11118 -2754 12638
rect -12430 9012 -12110 10532
rect -11544 9016 -10024 10536
rect -9504 9016 -7984 10536
rect -7304 9016 -5784 10536
rect -5264 9016 -3744 10536
rect -3074 9014 -2754 10534
rect -12249 7794 -9929 8114
rect -9466 7794 -7946 8114
rect -7078 7796 -5558 8116
rect -5095 7796 -2775 8116
rect -12187 6320 -9867 6640
rect -9404 6320 -7884 6640
rect -7016 6322 -5496 6642
rect -5033 6322 -2713 6642
rect -12368 3886 -12048 5406
rect -11482 3886 -9962 5406
rect -9442 3886 -7922 5406
rect -7242 3886 -5722 5406
rect -5202 3886 -3682 5406
rect -3012 3888 -2692 5408
rect -12368 1782 -12048 3302
rect -11482 1786 -9962 3306
rect -9442 1786 -7922 3306
rect -7242 1786 -5722 3306
rect -5202 1786 -3682 3306
rect -3012 1784 -2692 3304
rect -12187 564 -9867 884
rect -9404 564 -7884 884
rect -7016 566 -5496 886
rect -5033 566 -2713 886
<< metal4 >>
rect -4928 30756 35912 30940
rect -4928 30456 11396 30756
rect 11996 30456 35028 30756
rect 35628 30456 35912 30756
rect -4928 30374 35912 30456
rect -4928 30293 14973 30374
rect -4928 30229 -4463 30293
rect -4393 30229 14973 30293
rect -4928 30160 14973 30229
rect 31758 30160 35912 30374
rect -4928 30140 35912 30160
rect -4256 29480 10784 29626
rect -4256 29476 9938 29480
rect -4256 29470 2780 29476
rect -4256 28780 -4104 29470
rect -3408 29176 2780 29470
rect 3080 29176 9180 29476
rect 9480 29176 9938 29476
rect -3408 28782 9938 29176
rect 10628 28782 10784 29480
rect -3408 28780 10784 28782
rect -4256 28450 10784 28780
rect -4256 28394 -3074 28450
rect -4256 22694 -3706 28394
rect -3406 22694 -3074 28394
rect 9484 28394 10784 28450
rect -4256 21902 -3074 22694
rect -4256 16202 -3706 21902
rect -3406 16202 -3074 21902
rect -4256 15788 -3074 16202
rect -2316 27476 8684 27626
rect -2316 22776 2634 27476
rect 2934 22776 8234 27476
rect 8534 22776 8684 27476
rect -2316 21876 8684 22776
rect -2316 17176 2634 21876
rect 2934 17176 8234 21876
rect 8534 17176 8684 21876
rect -2316 16724 8684 17176
rect 9484 22694 10338 28394
rect 10638 22694 10784 28394
rect 9484 21902 10784 22694
rect 9484 17104 10338 21902
rect -2316 16627 9585 16724
rect -2316 16626 8684 16627
rect -2586 16162 8190 16244
rect 8078 15788 8190 16162
rect -4256 15702 8190 15788
rect -4254 15562 8190 15702
rect -4254 15476 9190 15562
rect -4254 15462 2280 15476
rect -4254 14780 -4102 15462
rect -3768 15176 2280 15462
rect 2580 15176 8680 15476
rect 8980 15176 9190 15476
rect -3768 14780 9190 15176
rect 9488 15140 9585 16627
rect 9854 16202 10338 17104
rect 10638 16202 10784 21902
rect 9854 15692 10784 16202
rect 11138 15595 13326 15596
rect 11138 15497 13227 15595
rect 13325 15497 13326 15595
rect 11138 15496 13326 15497
rect 11138 15140 11238 15496
rect 9488 15040 11238 15140
rect -12511 14688 -12409 14689
rect -12511 14588 -12510 14688
rect -12410 14588 -12409 14688
rect -4254 14624 9190 14780
rect -12511 14587 -12409 14588
rect -12510 13220 -12410 14587
rect 10952 14471 11052 15040
rect 10951 14470 11053 14471
rect 10951 14370 10952 14470
rect 11052 14370 11053 14470
rect 10951 14369 11053 14370
rect -6399 14122 -6255 14123
rect -8773 14118 -8611 14119
rect -11125 14114 -10953 14115
rect -11125 13944 -11124 14114
rect -10954 13944 -10953 14114
rect -8773 13958 -8772 14118
rect -8612 13958 -8611 14118
rect -6399 13980 -6398 14122
rect -6256 13980 -6255 14122
rect -6399 13979 -6255 13980
rect -4025 14106 -3861 14107
rect -8773 13957 -8611 13958
rect -11125 13943 -10953 13944
rect -11124 13871 -10954 13943
rect -8772 13871 -8612 13957
rect -6398 13873 -6256 13979
rect -4025 13944 -4024 14106
rect -3862 13944 -3861 14106
rect -4025 13943 -3861 13944
rect -4024 13873 -3862 13943
rect -7079 13872 -5557 13873
rect -12250 13870 -9928 13871
rect -12250 13550 -12249 13870
rect -9929 13550 -9928 13870
rect -12250 13549 -9928 13550
rect -9467 13870 -7945 13871
rect -9467 13550 -9466 13870
rect -7946 13550 -7945 13870
rect -7079 13552 -7078 13872
rect -5558 13552 -5557 13872
rect -7079 13551 -5557 13552
rect -5096 13872 -2774 13873
rect -5096 13552 -5095 13872
rect -2775 13552 -2774 13872
rect -5096 13551 -2774 13552
rect -9467 13549 -7945 13550
rect -12510 13120 -10034 13220
rect -10134 12904 -10034 13120
rect -10134 12903 -1758 12904
rect -10134 12805 -1857 12903
rect -1759 12805 -1758 12903
rect -10134 12804 -1758 12805
rect -10134 12637 -10034 12804
rect -12431 12636 -12109 12637
rect -12695 11918 -12595 11919
rect -12431 11918 -12430 12636
rect -12695 11820 -12694 11918
rect -12596 11820 -12430 11918
rect -12695 11819 -12595 11820
rect -12431 11116 -12430 11820
rect -12110 11116 -12109 12636
rect -12431 11115 -12109 11116
rect -11545 12636 -10023 12637
rect -11545 11116 -11544 12636
rect -10024 11116 -10023 12636
rect -11545 11115 -10023 11116
rect -9505 12636 -7983 12637
rect -9505 11116 -9504 12636
rect -7984 11884 -7983 12636
rect -7984 11784 -7706 11884
rect -7984 11116 -7983 11784
rect -9505 11115 -7983 11116
rect -9332 11021 -9232 11022
rect -9332 10923 -9331 11021
rect -9233 10923 -9232 11021
rect -9332 10726 -9232 10923
rect -13110 10725 -9232 10726
rect -13110 10627 -13109 10725
rect -13011 10627 -10155 10725
rect -10057 10627 -9232 10725
rect -13110 10626 -9232 10627
rect -8102 10881 -8002 10882
rect -8102 10783 -8101 10881
rect -8003 10783 -8002 10881
rect -8102 10537 -8002 10783
rect -11545 10536 -10023 10537
rect -12431 10532 -12109 10533
rect -12673 9826 -12553 9827
rect -12431 9826 -12430 10532
rect -12673 9708 -12672 9826
rect -12554 9708 -12430 9826
rect -12673 9707 -12553 9708
rect -12431 9012 -12430 9708
rect -12110 9012 -12109 10532
rect -11545 9016 -11544 10536
rect -10024 9016 -10023 10536
rect -11545 9015 -10023 9016
rect -9505 10536 -7983 10537
rect -9505 9016 -9504 10536
rect -7984 9016 -7983 10536
rect -9505 9015 -7983 9016
rect -12431 9011 -12109 9012
rect -10152 8864 -10052 9015
rect -7806 8864 -7706 11784
rect -7570 10883 -7470 12804
rect -5934 12637 -5834 12804
rect -7305 12636 -5783 12637
rect -7305 11116 -7304 12636
rect -5784 11116 -5783 12636
rect -7305 11115 -5783 11116
rect -5265 12636 -3743 12637
rect -5265 11116 -5264 12636
rect -3744 11884 -3743 12636
rect -3744 11784 -3506 11884
rect -3744 11116 -3743 11784
rect -5265 11115 -3743 11116
rect -5192 11029 -5092 11030
rect -5192 10931 -5191 11029
rect -5093 10931 -5092 11029
rect -7571 10882 -7469 10883
rect -7571 10782 -7570 10882
rect -7470 10782 -7469 10882
rect -7571 10781 -7469 10782
rect -5192 10726 -5092 10931
rect -5956 10725 -5092 10726
rect -5956 10627 -5955 10725
rect -5857 10627 -5092 10725
rect -5956 10626 -5092 10627
rect -3902 10879 -3802 10880
rect -3902 10781 -3901 10879
rect -3803 10781 -3802 10879
rect -3902 10537 -3802 10781
rect -7305 10536 -5783 10537
rect -7305 9016 -7304 10536
rect -5784 9016 -5783 10536
rect -7305 9015 -5783 9016
rect -5265 10536 -3743 10537
rect -5265 9016 -5264 10536
rect -3744 9016 -3743 10536
rect -5265 9015 -3743 9016
rect -5952 8864 -5852 9015
rect -3606 8864 -3506 11784
rect -3400 10881 -3300 12804
rect -3075 12638 -2753 12639
rect -3075 11118 -3074 12638
rect -2754 11908 -2753 12638
rect -2563 11908 -2439 11909
rect -2754 11786 -2562 11908
rect -2440 11786 -2439 11908
rect -2754 11118 -2753 11786
rect -2563 11785 -2439 11786
rect -3075 11117 -2753 11118
rect -3401 10880 -3299 10881
rect -3401 10780 -3400 10880
rect -3300 10780 -3299 10880
rect -3401 10779 -3299 10780
rect -3075 10534 -2753 10535
rect -3075 9014 -3074 10534
rect -2754 9850 -2753 10534
rect -2535 9850 -2425 9851
rect -2754 9742 -2534 9850
rect -2426 9742 -2425 9850
rect -2754 9014 -2753 9742
rect -2535 9741 -2425 9742
rect -3075 9013 -2753 9014
rect -10152 8863 -1500 8864
rect -10152 8765 -1599 8863
rect -1501 8765 -1500 8863
rect -10152 8764 -1500 8765
rect -10505 8616 -10403 8617
rect -13100 8615 -10504 8616
rect -13100 8517 -13099 8615
rect -13001 8517 -10504 8615
rect -13100 8516 -10504 8517
rect -10404 8516 -10403 8616
rect -10505 8515 -10403 8516
rect -7079 8116 -5557 8117
rect -12250 8114 -9928 8115
rect -12250 7794 -12249 8114
rect -9929 7794 -9928 8114
rect -12250 7793 -9928 7794
rect -9467 8114 -7945 8115
rect -9467 7794 -9466 8114
rect -7946 7794 -7945 8114
rect -7079 7796 -7078 8116
rect -5558 7796 -5557 8116
rect -7079 7795 -5557 7796
rect -5096 8116 -2774 8117
rect -5096 7796 -5095 8116
rect -2775 7796 -2774 8116
rect -5096 7795 -2774 7796
rect -9467 7793 -7945 7794
rect -11062 7570 -10892 7793
rect -11062 7402 -11061 7570
rect -10893 7402 -10892 7570
rect -11062 6885 -10892 7402
rect -8762 7570 -8592 7793
rect -8762 7402 -8761 7570
rect -8593 7402 -8592 7570
rect -8762 6885 -8592 7402
rect -6462 7570 -6292 7795
rect -6462 7402 -6461 7570
rect -6293 7402 -6292 7570
rect -6462 6885 -6292 7402
rect -4042 7570 -3872 7795
rect -4042 7402 -4041 7570
rect -3873 7402 -3872 7570
rect -4042 6885 -3872 7402
rect -11063 6884 -10891 6885
rect -11063 6714 -11062 6884
rect -10892 6714 -10891 6884
rect -11063 6713 -10891 6714
rect -8763 6884 -8591 6885
rect -8763 6714 -8762 6884
rect -8592 6714 -8591 6884
rect -8763 6713 -8591 6714
rect -6463 6884 -6291 6885
rect -6463 6714 -6462 6884
rect -6292 6714 -6291 6884
rect -6463 6713 -6291 6714
rect -4043 6884 -3871 6885
rect -4043 6714 -4042 6884
rect -3872 6714 -3871 6884
rect -4043 6713 -3871 6714
rect -11062 6641 -10892 6713
rect -8762 6641 -8592 6713
rect -6462 6643 -6292 6713
rect -4042 6643 -3872 6713
rect -7017 6642 -5495 6643
rect -12188 6640 -9866 6641
rect -12188 6320 -12187 6640
rect -9867 6320 -9866 6640
rect -12188 6319 -9866 6320
rect -9405 6640 -7883 6641
rect -9405 6320 -9404 6640
rect -7884 6320 -7883 6640
rect -7017 6322 -7016 6642
rect -5496 6322 -5495 6642
rect -7017 6321 -5495 6322
rect -5034 6642 -2712 6643
rect -5034 6322 -5033 6642
rect -2713 6322 -2712 6642
rect -5034 6321 -2712 6322
rect -9405 6319 -7883 6320
rect -11525 5904 -11423 5905
rect -13310 5903 -11524 5904
rect -13310 5805 -13309 5903
rect -13211 5805 -11524 5903
rect -13310 5804 -11524 5805
rect -11424 5804 -11423 5904
rect -11525 5803 -11423 5804
rect -10158 5665 -1758 5666
rect -10158 5567 -1857 5665
rect -1759 5567 -1758 5665
rect -10158 5566 -1758 5567
rect -10158 5407 -10058 5566
rect -12369 5406 -12047 5407
rect -12633 4688 -12533 4689
rect -12369 4688 -12368 5406
rect -12633 4590 -12632 4688
rect -12534 4590 -12368 4688
rect -12633 4589 -12533 4590
rect -12369 3886 -12368 4590
rect -12048 3886 -12047 5406
rect -12369 3885 -12047 3886
rect -11483 5406 -9961 5407
rect -11483 3886 -11482 5406
rect -9962 3886 -9961 5406
rect -11483 3885 -9961 3886
rect -9443 5406 -7921 5407
rect -9443 3886 -9442 5406
rect -7922 4646 -7921 5406
rect -7922 4546 -7690 4646
rect -7922 3886 -7921 4546
rect -9443 3885 -7921 3886
rect -9304 3797 -9204 3798
rect -9304 3699 -9303 3797
rect -9205 3699 -9204 3797
rect -9304 3498 -9204 3699
rect -13504 3497 -9204 3498
rect -13504 3399 -13503 3497
rect -13405 3399 -10179 3497
rect -10081 3399 -9204 3497
rect -13504 3398 -9204 3399
rect -8086 3643 -7986 3644
rect -8086 3545 -8085 3643
rect -7987 3545 -7986 3643
rect -8086 3307 -7986 3545
rect -11483 3306 -9961 3307
rect -12369 3302 -12047 3303
rect -12611 2596 -12491 2597
rect -12369 2596 -12368 3302
rect -12611 2478 -12610 2596
rect -12492 2478 -12368 2596
rect -12611 2477 -12491 2478
rect -12369 1782 -12368 2478
rect -12048 1782 -12047 3302
rect -11483 1786 -11482 3306
rect -9962 1786 -9961 3306
rect -11483 1785 -9961 1786
rect -9443 3306 -7921 3307
rect -9443 1786 -9442 3306
rect -7922 1786 -7921 3306
rect -9443 1785 -7921 1786
rect -12369 1781 -12047 1782
rect -10176 1628 -10076 1785
rect -13098 1627 -9512 1628
rect -13098 1529 -13097 1627
rect -12999 1626 -9512 1627
rect -7790 1626 -7690 4546
rect -7554 3645 -7454 5566
rect -5918 5407 -5818 5566
rect -7243 5406 -5721 5407
rect -7243 3886 -7242 5406
rect -5722 3886 -5721 5406
rect -7243 3885 -5721 3886
rect -5203 5406 -3681 5407
rect -5203 3886 -5202 5406
rect -3682 4646 -3681 5406
rect -3682 4546 -3450 4646
rect -3682 3886 -3681 4546
rect -5203 3885 -3681 3886
rect -5084 3801 -4984 3802
rect -5084 3703 -5083 3801
rect -4985 3703 -4984 3801
rect -7555 3644 -7453 3645
rect -7555 3544 -7554 3644
rect -7454 3544 -7453 3644
rect -7555 3543 -7453 3544
rect -5084 3502 -4984 3703
rect -5940 3501 -4984 3502
rect -5940 3403 -5939 3501
rect -5841 3403 -4984 3501
rect -5940 3402 -4984 3403
rect -3846 3643 -3746 3644
rect -3846 3545 -3845 3643
rect -3747 3545 -3746 3643
rect -3846 3307 -3746 3545
rect -7243 3306 -5721 3307
rect -7243 1786 -7242 3306
rect -5722 1786 -5721 3306
rect -7243 1785 -5721 1786
rect -5203 3306 -3681 3307
rect -5203 1786 -5202 3306
rect -3682 1786 -3681 3306
rect -5203 1785 -3681 1786
rect -5936 1626 -5836 1785
rect -3550 1626 -3450 4546
rect -3344 3645 -3244 5566
rect -3013 5408 -2691 5409
rect -3013 3888 -3012 5408
rect -2692 4678 -2691 5408
rect -2501 4678 -2377 4679
rect -2692 4556 -2500 4678
rect -2378 4556 -2377 4678
rect -2692 3888 -2691 4556
rect -2501 4555 -2377 4556
rect -3013 3887 -2691 3888
rect -3345 3644 -3243 3645
rect -3345 3544 -3344 3644
rect -3244 3544 -3243 3644
rect -3345 3543 -3243 3544
rect -3013 3304 -2691 3305
rect -3013 1784 -3012 3304
rect -2692 2620 -2691 3304
rect -2473 2620 -2363 2621
rect -2692 2512 -2472 2620
rect -2364 2512 -2363 2620
rect -2692 1784 -2691 2512
rect -2473 2511 -2363 2512
rect -3013 1783 -2691 1784
rect -12999 1625 -1486 1626
rect -12999 1529 -1585 1625
rect -13098 1528 -1585 1529
rect -10176 1527 -1585 1528
rect -1487 1527 -1486 1625
rect -10176 1526 -1486 1527
rect -7017 886 -5495 887
rect -12188 884 -9866 885
rect -12188 564 -12187 884
rect -9867 564 -9866 884
rect -12188 563 -9866 564
rect -9405 884 -7883 885
rect -9405 564 -9404 884
rect -7884 564 -7883 884
rect -7017 566 -7016 886
rect -5496 566 -5495 886
rect -7017 565 -5495 566
rect -5034 886 -2712 887
rect -5034 566 -5033 886
rect -2713 566 -2712 886
rect -5034 565 -2712 566
rect -9405 563 -7883 564
rect -11094 485 -10918 563
rect -8682 485 -8506 563
rect -6362 485 -6186 565
rect -3962 485 -3786 565
rect -11095 484 -10917 485
rect -11095 308 -11094 484
rect -10918 308 -10917 484
rect -11095 307 -10917 308
rect -8683 484 -8505 485
rect -8683 308 -8682 484
rect -8506 308 -8505 484
rect -8683 307 -8505 308
rect -6363 484 -6185 485
rect -6363 308 -6362 484
rect -6186 308 -6185 484
rect -6363 307 -6185 308
rect -3963 484 -3785 485
rect -3963 308 -3962 484
rect -3786 308 -3785 484
rect -3963 307 -3785 308
rect -11094 140 -10918 307
rect -8682 140 -8506 307
rect -6362 140 -6186 307
rect -3962 140 -3786 307
rect -13514 64 35912 140
rect -13514 -90 2840 64
rect 34840 -90 35912 64
rect -13514 -276 35912 -90
rect -13514 -576 -1304 -276
rect -704 -576 35128 -276
rect 35728 -576 35912 -276
rect -13514 -660 35912 -576
<< via4 >>
rect -4104 28780 -3408 29470
rect 9938 28782 10628 29480
rect -3074 28190 9484 28450
rect -3074 16162 -2786 28190
rect -2786 27986 9120 28190
rect -2786 16162 -2586 27986
rect 9028 17250 9120 27986
rect 9120 17250 9484 28190
rect 9028 17104 9484 17250
rect -3074 15788 8046 16162
rect 8046 15788 8078 16162
rect -4102 14780 -3768 15462
<< mimcap2 >>
rect -3070 29076 2730 29526
rect -3070 28776 -3020 29076
rect 2680 28776 2730 29076
rect -3070 28726 2730 28776
rect 3330 29076 9130 29526
rect 3330 28776 3380 29076
rect 9080 28776 9130 29076
rect 3330 28726 9130 28776
rect -4156 22594 -3756 28444
rect -4156 22294 -4106 22594
rect -3806 22294 -3756 22594
rect -2216 22676 2584 27526
rect -2216 22376 -2166 22676
rect 2534 22376 2584 22676
rect -2216 22326 2584 22376
rect 3384 22676 8184 27526
rect 3384 22376 3434 22676
rect 8134 22376 8184 22676
rect 3384 22326 8184 22376
rect 9888 22594 10288 28444
rect -4156 22244 -3756 22294
rect 9888 22294 9938 22594
rect 10238 22294 10288 22594
rect 9888 22244 10288 22294
rect -4156 16102 -3756 21952
rect -2216 17076 2584 21926
rect -2216 16776 -2166 17076
rect 2534 16776 2584 17076
rect -2216 16726 2584 16776
rect 3384 17076 8184 21926
rect 3384 16776 3434 17076
rect 8134 16776 8184 17076
rect 3384 16726 8184 16776
rect -4156 15802 -4106 16102
rect -3806 15802 -3756 16102
rect -4156 15752 -3756 15802
rect 9888 16102 10288 21952
rect 9888 15816 9938 16102
rect 10238 15816 10288 16102
rect 9888 15752 10288 15816
rect -3570 15076 2230 15526
rect -3570 14776 -3520 15076
rect 2180 14776 2230 15076
rect -3570 14726 2230 14776
rect 2830 15076 8630 15526
rect 2830 14776 2880 15076
rect 8580 14776 8630 15076
rect 2830 14726 8630 14776
<< mimcap2contact >>
rect -3020 28776 2680 29076
rect 3380 28776 9080 29076
rect -4106 22294 -3806 22594
rect -2166 22376 2534 22676
rect 3434 22376 8134 22676
rect 9938 22294 10238 22594
rect -2166 16776 2534 17076
rect 3434 16776 8134 17076
rect -4106 15802 -3806 16102
rect 9938 15816 10238 16102
rect -3520 14776 2180 15076
rect 2880 14776 8580 15076
<< metal5 >>
rect -4256 29480 10784 29626
rect -4256 29470 9938 29480
rect -4256 28780 -4104 29470
rect -3408 29076 9938 29470
rect -3408 28780 -3020 29076
rect -4256 28776 -3020 28780
rect 2680 28776 3380 29076
rect 9080 28782 9938 29076
rect 10628 28782 10784 29480
rect 9080 28776 10784 28782
rect -4256 28450 10784 28776
rect -4256 22594 -3074 28450
rect -4256 22294 -4106 22594
rect -3806 22294 -3074 22594
rect -4256 16102 -3074 22294
rect -2586 22676 9028 27986
rect -2586 22376 -2166 22676
rect 2534 22376 3434 22676
rect 8134 22376 9028 22676
rect -2586 17104 9028 22376
rect 9484 22594 10784 28450
rect 9484 22294 9938 22594
rect 10238 22294 10784 22594
rect 9484 17104 10784 22294
rect -2586 17076 10784 17104
rect -2586 16776 -2166 17076
rect 2534 16776 3434 17076
rect 8134 17022 10784 17076
rect 8134 16776 8186 17022
rect -2586 16162 8186 16776
rect -4256 15802 -4106 16102
rect -3806 15802 -3074 16102
rect -4256 15788 -3074 15802
rect 8078 15788 8186 16162
rect -4256 15558 8186 15788
rect 9840 16102 10784 17022
rect 9840 15816 9938 16102
rect 10238 15816 10784 16102
rect 9840 15776 10784 15816
rect -4256 15462 9084 15558
rect -4256 14780 -4102 15462
rect -3768 15076 9084 15462
rect -3768 14780 -3520 15076
rect -4256 14776 -3520 14780
rect 2180 14776 2880 15076
rect 8580 14776 9084 15076
rect -4256 14624 9084 14776
<< labels >>
flabel metal4 -5616 -342 -5562 -296 1 FreeSans 480 0 0 0 VSS
port 4 n ground bidirectional
flabel metal4 -9816 8794 -9798 8822 1 FreeSans 480 0 0 0 vse
port 6 n
flabel metal4 -9746 12834 -9732 12846 1 FreeSans 480 0 0 0 vip
flabel metal1 704 1582 716 1600 1 FreeSans 480 0 0 0 ibiasn
port 7 n
flabel metal4 -4738 30526 -4712 30558 1 FreeSans 480 0 0 0 VDD
port 3 n power bidirectional
flabel metal1 -7056 15480 -7054 15484 1 FreeSans 480 0 0 0 rst_n
port 8 n
flabel metal1 -7332 15474 -7328 15480 1 FreeSans 480 0 0 0 rst
flabel metal3 -9542 5852 -9520 5872 1 FreeSans 480 0 0 0 vdiffp
port 1 n
flabel metal4 -9702 5600 -9680 5618 1 FreeSans 480 0 0 0 vip
flabel metal4 -9786 1568 -9770 1582 1 FreeSans 480 0 0 0 vim
flabel metal3 -9812 1318 -9800 1332 1 FreeSans 480 0 0 0 vdiffm
port 2 n
flabel metal3 -9752 13102 -9732 13118 1 FreeSans 480 0 0 0 vocm
port 5 n
flabel metal3 -9862 8562 -9854 8578 1 FreeSans 480 0 0 0 vim
flabel metal1 -7485 15474 -7477 15480 1 FreeSans 480 0 0 0 txgate_1/tx
flabel metal1 -9303 15454 -9293 15462 1 FreeSans 480 0 0 0 txgate_1/out
flabel metal1 -9041 15460 -9031 15468 1 FreeSans 480 0 0 0 txgate_1/in
flabel metal1 -8787 16402 -8777 16412 1 FreeSans 480 0 0 0 txgate_1/VDD
flabel metal1 -8789 14712 -8781 14718 1 FreeSans 480 0 0 0 txgate_1/VSS
flabel metal2 -7787 15976 -7777 15984 1 FreeSans 480 0 0 0 txgate_1/txb
flabel locali -7718 15535 -7684 15569 0 FreeSans 340 0 0 0 txgate_1/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -7718 15467 -7684 15501 0 FreeSans 340 0 0 0 txgate_1/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -7626 15467 -7592 15501 0 FreeSans 340 0 0 0 txgate_1/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -7583 15773 -7549 15807 0 FreeSans 200 0 0 0 txgate_1/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -7583 15229 -7549 15263 0 FreeSans 200 0 0 0 txgate_1/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -7583 15229 -7549 15263 0 FreeSans 200 0 0 0 txgate_1/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -7583 15773 -7549 15807 0 FreeSans 200 0 0 0 txgate_1/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -7520 15246 -7520 15246 6 txgate_1/sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 -10085 15474 -10077 15480 1 FreeSans 480 0 0 0 txgate_0/tx
flabel metal1 -11903 15454 -11893 15462 1 FreeSans 480 0 0 0 txgate_0/out
flabel metal1 -11641 15460 -11631 15468 1 FreeSans 480 0 0 0 txgate_0/in
flabel metal1 -11387 16402 -11377 16412 1 FreeSans 480 0 0 0 txgate_0/VDD
flabel metal1 -11389 14712 -11381 14718 1 FreeSans 480 0 0 0 txgate_0/VSS
flabel metal2 -10387 15976 -10377 15984 1 FreeSans 480 0 0 0 txgate_0/txb
flabel locali -10318 15535 -10284 15569 0 FreeSans 340 0 0 0 txgate_0/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -10318 15467 -10284 15501 0 FreeSans 340 0 0 0 txgate_0/sky130_fd_sc_hd__inv_1_0/Y
flabel locali -10226 15467 -10192 15501 0 FreeSans 340 0 0 0 txgate_0/sky130_fd_sc_hd__inv_1_0/A
flabel nwell -10183 15773 -10149 15807 0 FreeSans 200 0 0 0 txgate_0/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -10183 15229 -10149 15263 0 FreeSans 200 0 0 0 txgate_0/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -10183 15229 -10149 15263 0 FreeSans 200 0 0 0 txgate_0/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -10183 15773 -10149 15807 0 FreeSans 200 0 0 0 txgate_0/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -10120 15246 -10120 15246 6 txgate_0/sky130_fd_sc_hd__inv_1_0/inv_1
flabel locali -7268 15535 -7234 15569 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali -7268 15467 -7234 15501 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali -7176 15467 -7142 15501 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/A
flabel nwell -7133 15773 -7099 15807 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -7133 15229 -7099 15263 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -7133 15229 -7099 15263 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -7133 15773 -7099 15807 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -7070 15246 -7070 15246 6 sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 2834 14188 2834 14188 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias1
flabel metal1 4706 7514 4706 7514 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias2
flabel metal1 34092 7222 34116 7252 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/VSS
flabel metal1 34468 8070 34468 8070 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias3
flabel metal1 34212 8276 34212 8276 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascnm
flabel metal1 34348 4044 34348 4044 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias4
flabel metal1 13050 8438 13078 8468 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vtail_cascn
flabel metal1 13368 11780 13400 11820 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascnp
flabel metal1 14234 14642 14324 14672 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M8d
flabel metal1 13156 8178 13194 8214 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vmirror
flabel metal1 33850 9910 33886 9940 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M16d
flabel metal1 266 5000 294 5044 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vip
flabel metal1 11866 5004 11898 5042 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vim
flabel metal1 5710 1574 5806 1610 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/ibiasn
flabel metal1 10860 4300 10908 4324 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vtail_cascn
flabel metal4 -8 -204 18 -182 1 FreeSans 3200 0 0 0 se_fold_casc_wide_swing_ota_0/VSS
flabel metal2 4348 6606 4396 6622 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpp
flabel metal1 1424 4372 1456 4400 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpm
flabel metal4 -792 30450 -766 30544 1 FreeSans 3200 0 0 0 se_fold_casc_wide_swing_ota_0/VDD
flabel metal4 11506 15538 11526 15558 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vo
flabel metal1 33520 18168 33526 18186 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vo
flabel metal1 18410 24990 18442 25022 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M9d
flabel metal1 13844 21532 13916 21562 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascnm
flabel metal1 16568 21540 16610 21562 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascnp
flabel metal1 15122 21502 15148 21540 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vtail_cascp
flabel metal1 14610 17494 14640 17520 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vip
flabel metal1 15618 17490 15648 17524 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vim
flabel metal2 31084 22150 31146 22178 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vmirror
flabel metal1 27122 24354 27174 24380 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/VDD
flabel metal2 21358 23312 21426 23342 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpp
flabel metal2 21582 22280 21634 22314 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpm
flabel metal2 19236 28424 19236 28424 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias1
flabel metal2 20214 28162 20244 28190 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/VDD
flabel metal1 17258 27150 17292 27172 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M7d
flabel metal2 18646 27026 18704 27062 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M13d
flabel metal2 20672 24846 20750 24880 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vtail_cascp
flabel metal1 28422 20680 28458 20708 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/VDD
flabel metal2 22778 16632 22832 16666 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M8d
flabel metal2 23202 21620 23284 21652 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias2
flabel metal2 27752 19110 27814 19140 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M16d
flabel metal2 27344 19422 27408 19454 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M13d
flabel metal1 18236 21460 18276 21494 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M7d
flabel metal2 33306 19322 33368 19354 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vmirror
flabel metal2 31420 19212 31470 19248 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpm
flabel metal2 31472 18164 31564 18196 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vcascpp
flabel metal2 18530 20492 18530 20492 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/vbias1
flabel metal2 18400 16906 18456 16940 1 FreeSans 480 0 0 0 se_fold_casc_wide_swing_ota_0/M9d
<< end >>
