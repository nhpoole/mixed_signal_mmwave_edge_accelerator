magic
tech sky130A
magscale 1 2
timestamp 1622264460
<< metal3 >>
rect -850 15222 849 15250
rect -850 13678 765 15222
rect 829 13678 849 15222
rect -850 13650 849 13678
rect -850 13522 849 13550
rect -850 11978 765 13522
rect 829 11978 849 13522
rect -850 11950 849 11978
rect -850 11822 849 11850
rect -850 10278 765 11822
rect 829 10278 849 11822
rect -850 10250 849 10278
rect -850 10122 849 10150
rect -850 8578 765 10122
rect 829 8578 849 10122
rect -850 8550 849 8578
rect -850 8422 849 8450
rect -850 6878 765 8422
rect 829 6878 849 8422
rect -850 6850 849 6878
rect -850 6722 849 6750
rect -850 5178 765 6722
rect 829 5178 849 6722
rect -850 5150 849 5178
rect -850 5022 849 5050
rect -850 3478 765 5022
rect 829 3478 849 5022
rect -850 3450 849 3478
rect -850 3322 849 3350
rect -850 1778 765 3322
rect 829 1778 849 3322
rect -850 1750 849 1778
rect -850 1622 849 1650
rect -850 78 765 1622
rect 829 78 849 1622
rect -850 50 849 78
rect -850 -78 849 -50
rect -850 -1622 765 -78
rect 829 -1622 849 -78
rect -850 -1650 849 -1622
rect -850 -1778 849 -1750
rect -850 -3322 765 -1778
rect 829 -3322 849 -1778
rect -850 -3350 849 -3322
rect -850 -3478 849 -3450
rect -850 -5022 765 -3478
rect 829 -5022 849 -3478
rect -850 -5050 849 -5022
rect -850 -5178 849 -5150
rect -850 -6722 765 -5178
rect 829 -6722 849 -5178
rect -850 -6750 849 -6722
rect -850 -6878 849 -6850
rect -850 -8422 765 -6878
rect 829 -8422 849 -6878
rect -850 -8450 849 -8422
rect -850 -8578 849 -8550
rect -850 -10122 765 -8578
rect 829 -10122 849 -8578
rect -850 -10150 849 -10122
rect -850 -10278 849 -10250
rect -850 -11822 765 -10278
rect 829 -11822 849 -10278
rect -850 -11850 849 -11822
rect -850 -11978 849 -11950
rect -850 -13522 765 -11978
rect 829 -13522 849 -11978
rect -850 -13550 849 -13522
rect -850 -13678 849 -13650
rect -850 -15222 765 -13678
rect 829 -15222 849 -13678
rect -850 -15250 849 -15222
<< via3 >>
rect 765 13678 829 15222
rect 765 11978 829 13522
rect 765 10278 829 11822
rect 765 8578 829 10122
rect 765 6878 829 8422
rect 765 5178 829 6722
rect 765 3478 829 5022
rect 765 1778 829 3322
rect 765 78 829 1622
rect 765 -1622 829 -78
rect 765 -3322 829 -1778
rect 765 -5022 829 -3478
rect 765 -6722 829 -5178
rect 765 -8422 829 -6878
rect 765 -10122 829 -8578
rect 765 -11822 829 -10278
rect 765 -13522 829 -11978
rect 765 -15222 829 -13678
<< mimcap >>
rect -750 15110 650 15150
rect -750 13790 -710 15110
rect 610 13790 650 15110
rect -750 13750 650 13790
rect -750 13410 650 13450
rect -750 12090 -710 13410
rect 610 12090 650 13410
rect -750 12050 650 12090
rect -750 11710 650 11750
rect -750 10390 -710 11710
rect 610 10390 650 11710
rect -750 10350 650 10390
rect -750 10010 650 10050
rect -750 8690 -710 10010
rect 610 8690 650 10010
rect -750 8650 650 8690
rect -750 8310 650 8350
rect -750 6990 -710 8310
rect 610 6990 650 8310
rect -750 6950 650 6990
rect -750 6610 650 6650
rect -750 5290 -710 6610
rect 610 5290 650 6610
rect -750 5250 650 5290
rect -750 4910 650 4950
rect -750 3590 -710 4910
rect 610 3590 650 4910
rect -750 3550 650 3590
rect -750 3210 650 3250
rect -750 1890 -710 3210
rect 610 1890 650 3210
rect -750 1850 650 1890
rect -750 1510 650 1550
rect -750 190 -710 1510
rect 610 190 650 1510
rect -750 150 650 190
rect -750 -190 650 -150
rect -750 -1510 -710 -190
rect 610 -1510 650 -190
rect -750 -1550 650 -1510
rect -750 -1890 650 -1850
rect -750 -3210 -710 -1890
rect 610 -3210 650 -1890
rect -750 -3250 650 -3210
rect -750 -3590 650 -3550
rect -750 -4910 -710 -3590
rect 610 -4910 650 -3590
rect -750 -4950 650 -4910
rect -750 -5290 650 -5250
rect -750 -6610 -710 -5290
rect 610 -6610 650 -5290
rect -750 -6650 650 -6610
rect -750 -6990 650 -6950
rect -750 -8310 -710 -6990
rect 610 -8310 650 -6990
rect -750 -8350 650 -8310
rect -750 -8690 650 -8650
rect -750 -10010 -710 -8690
rect 610 -10010 650 -8690
rect -750 -10050 650 -10010
rect -750 -10390 650 -10350
rect -750 -11710 -710 -10390
rect 610 -11710 650 -10390
rect -750 -11750 650 -11710
rect -750 -12090 650 -12050
rect -750 -13410 -710 -12090
rect 610 -13410 650 -12090
rect -750 -13450 650 -13410
rect -750 -13790 650 -13750
rect -750 -15110 -710 -13790
rect 610 -15110 650 -13790
rect -750 -15150 650 -15110
<< mimcapcontact >>
rect -710 13790 610 15110
rect -710 12090 610 13410
rect -710 10390 610 11710
rect -710 8690 610 10010
rect -710 6990 610 8310
rect -710 5290 610 6610
rect -710 3590 610 4910
rect -710 1890 610 3210
rect -710 190 610 1510
rect -710 -1510 610 -190
rect -710 -3210 610 -1890
rect -710 -4910 610 -3590
rect -710 -6610 610 -5290
rect -710 -8310 610 -6990
rect -710 -10010 610 -8690
rect -710 -11710 610 -10390
rect -710 -13410 610 -12090
rect -710 -15110 610 -13790
<< metal4 >>
rect 749 15222 845 15238
rect -711 15110 611 15111
rect -711 13790 -710 15110
rect 610 13790 611 15110
rect -711 13789 611 13790
rect 749 13678 765 15222
rect 829 13678 845 15222
rect 749 13662 845 13678
rect 749 13522 845 13538
rect -711 13410 611 13411
rect -711 12090 -710 13410
rect 610 12090 611 13410
rect -711 12089 611 12090
rect 749 11978 765 13522
rect 829 11978 845 13522
rect 749 11962 845 11978
rect 749 11822 845 11838
rect -711 11710 611 11711
rect -711 10390 -710 11710
rect 610 10390 611 11710
rect -711 10389 611 10390
rect 749 10278 765 11822
rect 829 10278 845 11822
rect 749 10262 845 10278
rect 749 10122 845 10138
rect -711 10010 611 10011
rect -711 8690 -710 10010
rect 610 8690 611 10010
rect -711 8689 611 8690
rect 749 8578 765 10122
rect 829 8578 845 10122
rect 749 8562 845 8578
rect 749 8422 845 8438
rect -711 8310 611 8311
rect -711 6990 -710 8310
rect 610 6990 611 8310
rect -711 6989 611 6990
rect 749 6878 765 8422
rect 829 6878 845 8422
rect 749 6862 845 6878
rect 749 6722 845 6738
rect -711 6610 611 6611
rect -711 5290 -710 6610
rect 610 5290 611 6610
rect -711 5289 611 5290
rect 749 5178 765 6722
rect 829 5178 845 6722
rect 749 5162 845 5178
rect 749 5022 845 5038
rect -711 4910 611 4911
rect -711 3590 -710 4910
rect 610 3590 611 4910
rect -711 3589 611 3590
rect 749 3478 765 5022
rect 829 3478 845 5022
rect 749 3462 845 3478
rect 749 3322 845 3338
rect -711 3210 611 3211
rect -711 1890 -710 3210
rect 610 1890 611 3210
rect -711 1889 611 1890
rect 749 1778 765 3322
rect 829 1778 845 3322
rect 749 1762 845 1778
rect 749 1622 845 1638
rect -711 1510 611 1511
rect -711 190 -710 1510
rect 610 190 611 1510
rect -711 189 611 190
rect 749 78 765 1622
rect 829 78 845 1622
rect 749 62 845 78
rect 749 -78 845 -62
rect -711 -190 611 -189
rect -711 -1510 -710 -190
rect 610 -1510 611 -190
rect -711 -1511 611 -1510
rect 749 -1622 765 -78
rect 829 -1622 845 -78
rect 749 -1638 845 -1622
rect 749 -1778 845 -1762
rect -711 -1890 611 -1889
rect -711 -3210 -710 -1890
rect 610 -3210 611 -1890
rect -711 -3211 611 -3210
rect 749 -3322 765 -1778
rect 829 -3322 845 -1778
rect 749 -3338 845 -3322
rect 749 -3478 845 -3462
rect -711 -3590 611 -3589
rect -711 -4910 -710 -3590
rect 610 -4910 611 -3590
rect -711 -4911 611 -4910
rect 749 -5022 765 -3478
rect 829 -5022 845 -3478
rect 749 -5038 845 -5022
rect 749 -5178 845 -5162
rect -711 -5290 611 -5289
rect -711 -6610 -710 -5290
rect 610 -6610 611 -5290
rect -711 -6611 611 -6610
rect 749 -6722 765 -5178
rect 829 -6722 845 -5178
rect 749 -6738 845 -6722
rect 749 -6878 845 -6862
rect -711 -6990 611 -6989
rect -711 -8310 -710 -6990
rect 610 -8310 611 -6990
rect -711 -8311 611 -8310
rect 749 -8422 765 -6878
rect 829 -8422 845 -6878
rect 749 -8438 845 -8422
rect 749 -8578 845 -8562
rect -711 -8690 611 -8689
rect -711 -10010 -710 -8690
rect 610 -10010 611 -8690
rect -711 -10011 611 -10010
rect 749 -10122 765 -8578
rect 829 -10122 845 -8578
rect 749 -10138 845 -10122
rect 749 -10278 845 -10262
rect -711 -10390 611 -10389
rect -711 -11710 -710 -10390
rect 610 -11710 611 -10390
rect -711 -11711 611 -11710
rect 749 -11822 765 -10278
rect 829 -11822 845 -10278
rect 749 -11838 845 -11822
rect 749 -11978 845 -11962
rect -711 -12090 611 -12089
rect -711 -13410 -710 -12090
rect 610 -13410 611 -12090
rect -711 -13411 611 -13410
rect 749 -13522 765 -11978
rect 829 -13522 845 -11978
rect 749 -13538 845 -13522
rect 749 -13678 845 -13662
rect -711 -13790 611 -13789
rect -711 -15110 -710 -13790
rect 610 -15110 611 -13790
rect -711 -15111 611 -15110
rect 749 -15222 765 -13678
rect 829 -15222 845 -13678
rect 749 -15238 845 -15222
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -850 13650 750 15250
string parameters w 7.00 l 7.00 val 103.32 carea 2.00 cperi 0.19 nx 1 ny 18 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
string library sky130
<< end >>
