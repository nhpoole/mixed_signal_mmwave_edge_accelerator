magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -7331 -1960 7331 1960
<< nwell >>
rect -6071 -700 6071 700
<< pmos >>
rect -5977 -600 -5177 600
rect -5119 -600 -4319 600
rect -4261 -600 -3461 600
rect -3403 -600 -2603 600
rect -2545 -600 -1745 600
rect -1687 -600 -887 600
rect -829 -600 -29 600
rect 29 -600 829 600
rect 887 -600 1687 600
rect 1745 -600 2545 600
rect 2603 -600 3403 600
rect 3461 -600 4261 600
rect 4319 -600 5119 600
rect 5177 -600 5977 600
<< pdiff >>
rect -6035 561 -5977 600
rect -6035 527 -6023 561
rect -5989 527 -5977 561
rect -6035 493 -5977 527
rect -6035 459 -6023 493
rect -5989 459 -5977 493
rect -6035 425 -5977 459
rect -6035 391 -6023 425
rect -5989 391 -5977 425
rect -6035 357 -5977 391
rect -6035 323 -6023 357
rect -5989 323 -5977 357
rect -6035 289 -5977 323
rect -6035 255 -6023 289
rect -5989 255 -5977 289
rect -6035 221 -5977 255
rect -6035 187 -6023 221
rect -5989 187 -5977 221
rect -6035 153 -5977 187
rect -6035 119 -6023 153
rect -5989 119 -5977 153
rect -6035 85 -5977 119
rect -6035 51 -6023 85
rect -5989 51 -5977 85
rect -6035 17 -5977 51
rect -6035 -17 -6023 17
rect -5989 -17 -5977 17
rect -6035 -51 -5977 -17
rect -6035 -85 -6023 -51
rect -5989 -85 -5977 -51
rect -6035 -119 -5977 -85
rect -6035 -153 -6023 -119
rect -5989 -153 -5977 -119
rect -6035 -187 -5977 -153
rect -6035 -221 -6023 -187
rect -5989 -221 -5977 -187
rect -6035 -255 -5977 -221
rect -6035 -289 -6023 -255
rect -5989 -289 -5977 -255
rect -6035 -323 -5977 -289
rect -6035 -357 -6023 -323
rect -5989 -357 -5977 -323
rect -6035 -391 -5977 -357
rect -6035 -425 -6023 -391
rect -5989 -425 -5977 -391
rect -6035 -459 -5977 -425
rect -6035 -493 -6023 -459
rect -5989 -493 -5977 -459
rect -6035 -527 -5977 -493
rect -6035 -561 -6023 -527
rect -5989 -561 -5977 -527
rect -6035 -600 -5977 -561
rect -5177 561 -5119 600
rect -5177 527 -5165 561
rect -5131 527 -5119 561
rect -5177 493 -5119 527
rect -5177 459 -5165 493
rect -5131 459 -5119 493
rect -5177 425 -5119 459
rect -5177 391 -5165 425
rect -5131 391 -5119 425
rect -5177 357 -5119 391
rect -5177 323 -5165 357
rect -5131 323 -5119 357
rect -5177 289 -5119 323
rect -5177 255 -5165 289
rect -5131 255 -5119 289
rect -5177 221 -5119 255
rect -5177 187 -5165 221
rect -5131 187 -5119 221
rect -5177 153 -5119 187
rect -5177 119 -5165 153
rect -5131 119 -5119 153
rect -5177 85 -5119 119
rect -5177 51 -5165 85
rect -5131 51 -5119 85
rect -5177 17 -5119 51
rect -5177 -17 -5165 17
rect -5131 -17 -5119 17
rect -5177 -51 -5119 -17
rect -5177 -85 -5165 -51
rect -5131 -85 -5119 -51
rect -5177 -119 -5119 -85
rect -5177 -153 -5165 -119
rect -5131 -153 -5119 -119
rect -5177 -187 -5119 -153
rect -5177 -221 -5165 -187
rect -5131 -221 -5119 -187
rect -5177 -255 -5119 -221
rect -5177 -289 -5165 -255
rect -5131 -289 -5119 -255
rect -5177 -323 -5119 -289
rect -5177 -357 -5165 -323
rect -5131 -357 -5119 -323
rect -5177 -391 -5119 -357
rect -5177 -425 -5165 -391
rect -5131 -425 -5119 -391
rect -5177 -459 -5119 -425
rect -5177 -493 -5165 -459
rect -5131 -493 -5119 -459
rect -5177 -527 -5119 -493
rect -5177 -561 -5165 -527
rect -5131 -561 -5119 -527
rect -5177 -600 -5119 -561
rect -4319 561 -4261 600
rect -4319 527 -4307 561
rect -4273 527 -4261 561
rect -4319 493 -4261 527
rect -4319 459 -4307 493
rect -4273 459 -4261 493
rect -4319 425 -4261 459
rect -4319 391 -4307 425
rect -4273 391 -4261 425
rect -4319 357 -4261 391
rect -4319 323 -4307 357
rect -4273 323 -4261 357
rect -4319 289 -4261 323
rect -4319 255 -4307 289
rect -4273 255 -4261 289
rect -4319 221 -4261 255
rect -4319 187 -4307 221
rect -4273 187 -4261 221
rect -4319 153 -4261 187
rect -4319 119 -4307 153
rect -4273 119 -4261 153
rect -4319 85 -4261 119
rect -4319 51 -4307 85
rect -4273 51 -4261 85
rect -4319 17 -4261 51
rect -4319 -17 -4307 17
rect -4273 -17 -4261 17
rect -4319 -51 -4261 -17
rect -4319 -85 -4307 -51
rect -4273 -85 -4261 -51
rect -4319 -119 -4261 -85
rect -4319 -153 -4307 -119
rect -4273 -153 -4261 -119
rect -4319 -187 -4261 -153
rect -4319 -221 -4307 -187
rect -4273 -221 -4261 -187
rect -4319 -255 -4261 -221
rect -4319 -289 -4307 -255
rect -4273 -289 -4261 -255
rect -4319 -323 -4261 -289
rect -4319 -357 -4307 -323
rect -4273 -357 -4261 -323
rect -4319 -391 -4261 -357
rect -4319 -425 -4307 -391
rect -4273 -425 -4261 -391
rect -4319 -459 -4261 -425
rect -4319 -493 -4307 -459
rect -4273 -493 -4261 -459
rect -4319 -527 -4261 -493
rect -4319 -561 -4307 -527
rect -4273 -561 -4261 -527
rect -4319 -600 -4261 -561
rect -3461 561 -3403 600
rect -3461 527 -3449 561
rect -3415 527 -3403 561
rect -3461 493 -3403 527
rect -3461 459 -3449 493
rect -3415 459 -3403 493
rect -3461 425 -3403 459
rect -3461 391 -3449 425
rect -3415 391 -3403 425
rect -3461 357 -3403 391
rect -3461 323 -3449 357
rect -3415 323 -3403 357
rect -3461 289 -3403 323
rect -3461 255 -3449 289
rect -3415 255 -3403 289
rect -3461 221 -3403 255
rect -3461 187 -3449 221
rect -3415 187 -3403 221
rect -3461 153 -3403 187
rect -3461 119 -3449 153
rect -3415 119 -3403 153
rect -3461 85 -3403 119
rect -3461 51 -3449 85
rect -3415 51 -3403 85
rect -3461 17 -3403 51
rect -3461 -17 -3449 17
rect -3415 -17 -3403 17
rect -3461 -51 -3403 -17
rect -3461 -85 -3449 -51
rect -3415 -85 -3403 -51
rect -3461 -119 -3403 -85
rect -3461 -153 -3449 -119
rect -3415 -153 -3403 -119
rect -3461 -187 -3403 -153
rect -3461 -221 -3449 -187
rect -3415 -221 -3403 -187
rect -3461 -255 -3403 -221
rect -3461 -289 -3449 -255
rect -3415 -289 -3403 -255
rect -3461 -323 -3403 -289
rect -3461 -357 -3449 -323
rect -3415 -357 -3403 -323
rect -3461 -391 -3403 -357
rect -3461 -425 -3449 -391
rect -3415 -425 -3403 -391
rect -3461 -459 -3403 -425
rect -3461 -493 -3449 -459
rect -3415 -493 -3403 -459
rect -3461 -527 -3403 -493
rect -3461 -561 -3449 -527
rect -3415 -561 -3403 -527
rect -3461 -600 -3403 -561
rect -2603 561 -2545 600
rect -2603 527 -2591 561
rect -2557 527 -2545 561
rect -2603 493 -2545 527
rect -2603 459 -2591 493
rect -2557 459 -2545 493
rect -2603 425 -2545 459
rect -2603 391 -2591 425
rect -2557 391 -2545 425
rect -2603 357 -2545 391
rect -2603 323 -2591 357
rect -2557 323 -2545 357
rect -2603 289 -2545 323
rect -2603 255 -2591 289
rect -2557 255 -2545 289
rect -2603 221 -2545 255
rect -2603 187 -2591 221
rect -2557 187 -2545 221
rect -2603 153 -2545 187
rect -2603 119 -2591 153
rect -2557 119 -2545 153
rect -2603 85 -2545 119
rect -2603 51 -2591 85
rect -2557 51 -2545 85
rect -2603 17 -2545 51
rect -2603 -17 -2591 17
rect -2557 -17 -2545 17
rect -2603 -51 -2545 -17
rect -2603 -85 -2591 -51
rect -2557 -85 -2545 -51
rect -2603 -119 -2545 -85
rect -2603 -153 -2591 -119
rect -2557 -153 -2545 -119
rect -2603 -187 -2545 -153
rect -2603 -221 -2591 -187
rect -2557 -221 -2545 -187
rect -2603 -255 -2545 -221
rect -2603 -289 -2591 -255
rect -2557 -289 -2545 -255
rect -2603 -323 -2545 -289
rect -2603 -357 -2591 -323
rect -2557 -357 -2545 -323
rect -2603 -391 -2545 -357
rect -2603 -425 -2591 -391
rect -2557 -425 -2545 -391
rect -2603 -459 -2545 -425
rect -2603 -493 -2591 -459
rect -2557 -493 -2545 -459
rect -2603 -527 -2545 -493
rect -2603 -561 -2591 -527
rect -2557 -561 -2545 -527
rect -2603 -600 -2545 -561
rect -1745 561 -1687 600
rect -1745 527 -1733 561
rect -1699 527 -1687 561
rect -1745 493 -1687 527
rect -1745 459 -1733 493
rect -1699 459 -1687 493
rect -1745 425 -1687 459
rect -1745 391 -1733 425
rect -1699 391 -1687 425
rect -1745 357 -1687 391
rect -1745 323 -1733 357
rect -1699 323 -1687 357
rect -1745 289 -1687 323
rect -1745 255 -1733 289
rect -1699 255 -1687 289
rect -1745 221 -1687 255
rect -1745 187 -1733 221
rect -1699 187 -1687 221
rect -1745 153 -1687 187
rect -1745 119 -1733 153
rect -1699 119 -1687 153
rect -1745 85 -1687 119
rect -1745 51 -1733 85
rect -1699 51 -1687 85
rect -1745 17 -1687 51
rect -1745 -17 -1733 17
rect -1699 -17 -1687 17
rect -1745 -51 -1687 -17
rect -1745 -85 -1733 -51
rect -1699 -85 -1687 -51
rect -1745 -119 -1687 -85
rect -1745 -153 -1733 -119
rect -1699 -153 -1687 -119
rect -1745 -187 -1687 -153
rect -1745 -221 -1733 -187
rect -1699 -221 -1687 -187
rect -1745 -255 -1687 -221
rect -1745 -289 -1733 -255
rect -1699 -289 -1687 -255
rect -1745 -323 -1687 -289
rect -1745 -357 -1733 -323
rect -1699 -357 -1687 -323
rect -1745 -391 -1687 -357
rect -1745 -425 -1733 -391
rect -1699 -425 -1687 -391
rect -1745 -459 -1687 -425
rect -1745 -493 -1733 -459
rect -1699 -493 -1687 -459
rect -1745 -527 -1687 -493
rect -1745 -561 -1733 -527
rect -1699 -561 -1687 -527
rect -1745 -600 -1687 -561
rect -887 561 -829 600
rect -887 527 -875 561
rect -841 527 -829 561
rect -887 493 -829 527
rect -887 459 -875 493
rect -841 459 -829 493
rect -887 425 -829 459
rect -887 391 -875 425
rect -841 391 -829 425
rect -887 357 -829 391
rect -887 323 -875 357
rect -841 323 -829 357
rect -887 289 -829 323
rect -887 255 -875 289
rect -841 255 -829 289
rect -887 221 -829 255
rect -887 187 -875 221
rect -841 187 -829 221
rect -887 153 -829 187
rect -887 119 -875 153
rect -841 119 -829 153
rect -887 85 -829 119
rect -887 51 -875 85
rect -841 51 -829 85
rect -887 17 -829 51
rect -887 -17 -875 17
rect -841 -17 -829 17
rect -887 -51 -829 -17
rect -887 -85 -875 -51
rect -841 -85 -829 -51
rect -887 -119 -829 -85
rect -887 -153 -875 -119
rect -841 -153 -829 -119
rect -887 -187 -829 -153
rect -887 -221 -875 -187
rect -841 -221 -829 -187
rect -887 -255 -829 -221
rect -887 -289 -875 -255
rect -841 -289 -829 -255
rect -887 -323 -829 -289
rect -887 -357 -875 -323
rect -841 -357 -829 -323
rect -887 -391 -829 -357
rect -887 -425 -875 -391
rect -841 -425 -829 -391
rect -887 -459 -829 -425
rect -887 -493 -875 -459
rect -841 -493 -829 -459
rect -887 -527 -829 -493
rect -887 -561 -875 -527
rect -841 -561 -829 -527
rect -887 -600 -829 -561
rect -29 561 29 600
rect -29 527 -17 561
rect 17 527 29 561
rect -29 493 29 527
rect -29 459 -17 493
rect 17 459 29 493
rect -29 425 29 459
rect -29 391 -17 425
rect 17 391 29 425
rect -29 357 29 391
rect -29 323 -17 357
rect 17 323 29 357
rect -29 289 29 323
rect -29 255 -17 289
rect 17 255 29 289
rect -29 221 29 255
rect -29 187 -17 221
rect 17 187 29 221
rect -29 153 29 187
rect -29 119 -17 153
rect 17 119 29 153
rect -29 85 29 119
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -119 29 -85
rect -29 -153 -17 -119
rect 17 -153 29 -119
rect -29 -187 29 -153
rect -29 -221 -17 -187
rect 17 -221 29 -187
rect -29 -255 29 -221
rect -29 -289 -17 -255
rect 17 -289 29 -255
rect -29 -323 29 -289
rect -29 -357 -17 -323
rect 17 -357 29 -323
rect -29 -391 29 -357
rect -29 -425 -17 -391
rect 17 -425 29 -391
rect -29 -459 29 -425
rect -29 -493 -17 -459
rect 17 -493 29 -459
rect -29 -527 29 -493
rect -29 -561 -17 -527
rect 17 -561 29 -527
rect -29 -600 29 -561
rect 829 561 887 600
rect 829 527 841 561
rect 875 527 887 561
rect 829 493 887 527
rect 829 459 841 493
rect 875 459 887 493
rect 829 425 887 459
rect 829 391 841 425
rect 875 391 887 425
rect 829 357 887 391
rect 829 323 841 357
rect 875 323 887 357
rect 829 289 887 323
rect 829 255 841 289
rect 875 255 887 289
rect 829 221 887 255
rect 829 187 841 221
rect 875 187 887 221
rect 829 153 887 187
rect 829 119 841 153
rect 875 119 887 153
rect 829 85 887 119
rect 829 51 841 85
rect 875 51 887 85
rect 829 17 887 51
rect 829 -17 841 17
rect 875 -17 887 17
rect 829 -51 887 -17
rect 829 -85 841 -51
rect 875 -85 887 -51
rect 829 -119 887 -85
rect 829 -153 841 -119
rect 875 -153 887 -119
rect 829 -187 887 -153
rect 829 -221 841 -187
rect 875 -221 887 -187
rect 829 -255 887 -221
rect 829 -289 841 -255
rect 875 -289 887 -255
rect 829 -323 887 -289
rect 829 -357 841 -323
rect 875 -357 887 -323
rect 829 -391 887 -357
rect 829 -425 841 -391
rect 875 -425 887 -391
rect 829 -459 887 -425
rect 829 -493 841 -459
rect 875 -493 887 -459
rect 829 -527 887 -493
rect 829 -561 841 -527
rect 875 -561 887 -527
rect 829 -600 887 -561
rect 1687 561 1745 600
rect 1687 527 1699 561
rect 1733 527 1745 561
rect 1687 493 1745 527
rect 1687 459 1699 493
rect 1733 459 1745 493
rect 1687 425 1745 459
rect 1687 391 1699 425
rect 1733 391 1745 425
rect 1687 357 1745 391
rect 1687 323 1699 357
rect 1733 323 1745 357
rect 1687 289 1745 323
rect 1687 255 1699 289
rect 1733 255 1745 289
rect 1687 221 1745 255
rect 1687 187 1699 221
rect 1733 187 1745 221
rect 1687 153 1745 187
rect 1687 119 1699 153
rect 1733 119 1745 153
rect 1687 85 1745 119
rect 1687 51 1699 85
rect 1733 51 1745 85
rect 1687 17 1745 51
rect 1687 -17 1699 17
rect 1733 -17 1745 17
rect 1687 -51 1745 -17
rect 1687 -85 1699 -51
rect 1733 -85 1745 -51
rect 1687 -119 1745 -85
rect 1687 -153 1699 -119
rect 1733 -153 1745 -119
rect 1687 -187 1745 -153
rect 1687 -221 1699 -187
rect 1733 -221 1745 -187
rect 1687 -255 1745 -221
rect 1687 -289 1699 -255
rect 1733 -289 1745 -255
rect 1687 -323 1745 -289
rect 1687 -357 1699 -323
rect 1733 -357 1745 -323
rect 1687 -391 1745 -357
rect 1687 -425 1699 -391
rect 1733 -425 1745 -391
rect 1687 -459 1745 -425
rect 1687 -493 1699 -459
rect 1733 -493 1745 -459
rect 1687 -527 1745 -493
rect 1687 -561 1699 -527
rect 1733 -561 1745 -527
rect 1687 -600 1745 -561
rect 2545 561 2603 600
rect 2545 527 2557 561
rect 2591 527 2603 561
rect 2545 493 2603 527
rect 2545 459 2557 493
rect 2591 459 2603 493
rect 2545 425 2603 459
rect 2545 391 2557 425
rect 2591 391 2603 425
rect 2545 357 2603 391
rect 2545 323 2557 357
rect 2591 323 2603 357
rect 2545 289 2603 323
rect 2545 255 2557 289
rect 2591 255 2603 289
rect 2545 221 2603 255
rect 2545 187 2557 221
rect 2591 187 2603 221
rect 2545 153 2603 187
rect 2545 119 2557 153
rect 2591 119 2603 153
rect 2545 85 2603 119
rect 2545 51 2557 85
rect 2591 51 2603 85
rect 2545 17 2603 51
rect 2545 -17 2557 17
rect 2591 -17 2603 17
rect 2545 -51 2603 -17
rect 2545 -85 2557 -51
rect 2591 -85 2603 -51
rect 2545 -119 2603 -85
rect 2545 -153 2557 -119
rect 2591 -153 2603 -119
rect 2545 -187 2603 -153
rect 2545 -221 2557 -187
rect 2591 -221 2603 -187
rect 2545 -255 2603 -221
rect 2545 -289 2557 -255
rect 2591 -289 2603 -255
rect 2545 -323 2603 -289
rect 2545 -357 2557 -323
rect 2591 -357 2603 -323
rect 2545 -391 2603 -357
rect 2545 -425 2557 -391
rect 2591 -425 2603 -391
rect 2545 -459 2603 -425
rect 2545 -493 2557 -459
rect 2591 -493 2603 -459
rect 2545 -527 2603 -493
rect 2545 -561 2557 -527
rect 2591 -561 2603 -527
rect 2545 -600 2603 -561
rect 3403 561 3461 600
rect 3403 527 3415 561
rect 3449 527 3461 561
rect 3403 493 3461 527
rect 3403 459 3415 493
rect 3449 459 3461 493
rect 3403 425 3461 459
rect 3403 391 3415 425
rect 3449 391 3461 425
rect 3403 357 3461 391
rect 3403 323 3415 357
rect 3449 323 3461 357
rect 3403 289 3461 323
rect 3403 255 3415 289
rect 3449 255 3461 289
rect 3403 221 3461 255
rect 3403 187 3415 221
rect 3449 187 3461 221
rect 3403 153 3461 187
rect 3403 119 3415 153
rect 3449 119 3461 153
rect 3403 85 3461 119
rect 3403 51 3415 85
rect 3449 51 3461 85
rect 3403 17 3461 51
rect 3403 -17 3415 17
rect 3449 -17 3461 17
rect 3403 -51 3461 -17
rect 3403 -85 3415 -51
rect 3449 -85 3461 -51
rect 3403 -119 3461 -85
rect 3403 -153 3415 -119
rect 3449 -153 3461 -119
rect 3403 -187 3461 -153
rect 3403 -221 3415 -187
rect 3449 -221 3461 -187
rect 3403 -255 3461 -221
rect 3403 -289 3415 -255
rect 3449 -289 3461 -255
rect 3403 -323 3461 -289
rect 3403 -357 3415 -323
rect 3449 -357 3461 -323
rect 3403 -391 3461 -357
rect 3403 -425 3415 -391
rect 3449 -425 3461 -391
rect 3403 -459 3461 -425
rect 3403 -493 3415 -459
rect 3449 -493 3461 -459
rect 3403 -527 3461 -493
rect 3403 -561 3415 -527
rect 3449 -561 3461 -527
rect 3403 -600 3461 -561
rect 4261 561 4319 600
rect 4261 527 4273 561
rect 4307 527 4319 561
rect 4261 493 4319 527
rect 4261 459 4273 493
rect 4307 459 4319 493
rect 4261 425 4319 459
rect 4261 391 4273 425
rect 4307 391 4319 425
rect 4261 357 4319 391
rect 4261 323 4273 357
rect 4307 323 4319 357
rect 4261 289 4319 323
rect 4261 255 4273 289
rect 4307 255 4319 289
rect 4261 221 4319 255
rect 4261 187 4273 221
rect 4307 187 4319 221
rect 4261 153 4319 187
rect 4261 119 4273 153
rect 4307 119 4319 153
rect 4261 85 4319 119
rect 4261 51 4273 85
rect 4307 51 4319 85
rect 4261 17 4319 51
rect 4261 -17 4273 17
rect 4307 -17 4319 17
rect 4261 -51 4319 -17
rect 4261 -85 4273 -51
rect 4307 -85 4319 -51
rect 4261 -119 4319 -85
rect 4261 -153 4273 -119
rect 4307 -153 4319 -119
rect 4261 -187 4319 -153
rect 4261 -221 4273 -187
rect 4307 -221 4319 -187
rect 4261 -255 4319 -221
rect 4261 -289 4273 -255
rect 4307 -289 4319 -255
rect 4261 -323 4319 -289
rect 4261 -357 4273 -323
rect 4307 -357 4319 -323
rect 4261 -391 4319 -357
rect 4261 -425 4273 -391
rect 4307 -425 4319 -391
rect 4261 -459 4319 -425
rect 4261 -493 4273 -459
rect 4307 -493 4319 -459
rect 4261 -527 4319 -493
rect 4261 -561 4273 -527
rect 4307 -561 4319 -527
rect 4261 -600 4319 -561
rect 5119 561 5177 600
rect 5119 527 5131 561
rect 5165 527 5177 561
rect 5119 493 5177 527
rect 5119 459 5131 493
rect 5165 459 5177 493
rect 5119 425 5177 459
rect 5119 391 5131 425
rect 5165 391 5177 425
rect 5119 357 5177 391
rect 5119 323 5131 357
rect 5165 323 5177 357
rect 5119 289 5177 323
rect 5119 255 5131 289
rect 5165 255 5177 289
rect 5119 221 5177 255
rect 5119 187 5131 221
rect 5165 187 5177 221
rect 5119 153 5177 187
rect 5119 119 5131 153
rect 5165 119 5177 153
rect 5119 85 5177 119
rect 5119 51 5131 85
rect 5165 51 5177 85
rect 5119 17 5177 51
rect 5119 -17 5131 17
rect 5165 -17 5177 17
rect 5119 -51 5177 -17
rect 5119 -85 5131 -51
rect 5165 -85 5177 -51
rect 5119 -119 5177 -85
rect 5119 -153 5131 -119
rect 5165 -153 5177 -119
rect 5119 -187 5177 -153
rect 5119 -221 5131 -187
rect 5165 -221 5177 -187
rect 5119 -255 5177 -221
rect 5119 -289 5131 -255
rect 5165 -289 5177 -255
rect 5119 -323 5177 -289
rect 5119 -357 5131 -323
rect 5165 -357 5177 -323
rect 5119 -391 5177 -357
rect 5119 -425 5131 -391
rect 5165 -425 5177 -391
rect 5119 -459 5177 -425
rect 5119 -493 5131 -459
rect 5165 -493 5177 -459
rect 5119 -527 5177 -493
rect 5119 -561 5131 -527
rect 5165 -561 5177 -527
rect 5119 -600 5177 -561
rect 5977 561 6035 600
rect 5977 527 5989 561
rect 6023 527 6035 561
rect 5977 493 6035 527
rect 5977 459 5989 493
rect 6023 459 6035 493
rect 5977 425 6035 459
rect 5977 391 5989 425
rect 6023 391 6035 425
rect 5977 357 6035 391
rect 5977 323 5989 357
rect 6023 323 6035 357
rect 5977 289 6035 323
rect 5977 255 5989 289
rect 6023 255 6035 289
rect 5977 221 6035 255
rect 5977 187 5989 221
rect 6023 187 6035 221
rect 5977 153 6035 187
rect 5977 119 5989 153
rect 6023 119 6035 153
rect 5977 85 6035 119
rect 5977 51 5989 85
rect 6023 51 6035 85
rect 5977 17 6035 51
rect 5977 -17 5989 17
rect 6023 -17 6035 17
rect 5977 -51 6035 -17
rect 5977 -85 5989 -51
rect 6023 -85 6035 -51
rect 5977 -119 6035 -85
rect 5977 -153 5989 -119
rect 6023 -153 6035 -119
rect 5977 -187 6035 -153
rect 5977 -221 5989 -187
rect 6023 -221 6035 -187
rect 5977 -255 6035 -221
rect 5977 -289 5989 -255
rect 6023 -289 6035 -255
rect 5977 -323 6035 -289
rect 5977 -357 5989 -323
rect 6023 -357 6035 -323
rect 5977 -391 6035 -357
rect 5977 -425 5989 -391
rect 6023 -425 6035 -391
rect 5977 -459 6035 -425
rect 5977 -493 5989 -459
rect 6023 -493 6035 -459
rect 5977 -527 6035 -493
rect 5977 -561 5989 -527
rect 6023 -561 6035 -527
rect 5977 -600 6035 -561
<< pdiffc >>
rect -6023 527 -5989 561
rect -6023 459 -5989 493
rect -6023 391 -5989 425
rect -6023 323 -5989 357
rect -6023 255 -5989 289
rect -6023 187 -5989 221
rect -6023 119 -5989 153
rect -6023 51 -5989 85
rect -6023 -17 -5989 17
rect -6023 -85 -5989 -51
rect -6023 -153 -5989 -119
rect -6023 -221 -5989 -187
rect -6023 -289 -5989 -255
rect -6023 -357 -5989 -323
rect -6023 -425 -5989 -391
rect -6023 -493 -5989 -459
rect -6023 -561 -5989 -527
rect -5165 527 -5131 561
rect -5165 459 -5131 493
rect -5165 391 -5131 425
rect -5165 323 -5131 357
rect -5165 255 -5131 289
rect -5165 187 -5131 221
rect -5165 119 -5131 153
rect -5165 51 -5131 85
rect -5165 -17 -5131 17
rect -5165 -85 -5131 -51
rect -5165 -153 -5131 -119
rect -5165 -221 -5131 -187
rect -5165 -289 -5131 -255
rect -5165 -357 -5131 -323
rect -5165 -425 -5131 -391
rect -5165 -493 -5131 -459
rect -5165 -561 -5131 -527
rect -4307 527 -4273 561
rect -4307 459 -4273 493
rect -4307 391 -4273 425
rect -4307 323 -4273 357
rect -4307 255 -4273 289
rect -4307 187 -4273 221
rect -4307 119 -4273 153
rect -4307 51 -4273 85
rect -4307 -17 -4273 17
rect -4307 -85 -4273 -51
rect -4307 -153 -4273 -119
rect -4307 -221 -4273 -187
rect -4307 -289 -4273 -255
rect -4307 -357 -4273 -323
rect -4307 -425 -4273 -391
rect -4307 -493 -4273 -459
rect -4307 -561 -4273 -527
rect -3449 527 -3415 561
rect -3449 459 -3415 493
rect -3449 391 -3415 425
rect -3449 323 -3415 357
rect -3449 255 -3415 289
rect -3449 187 -3415 221
rect -3449 119 -3415 153
rect -3449 51 -3415 85
rect -3449 -17 -3415 17
rect -3449 -85 -3415 -51
rect -3449 -153 -3415 -119
rect -3449 -221 -3415 -187
rect -3449 -289 -3415 -255
rect -3449 -357 -3415 -323
rect -3449 -425 -3415 -391
rect -3449 -493 -3415 -459
rect -3449 -561 -3415 -527
rect -2591 527 -2557 561
rect -2591 459 -2557 493
rect -2591 391 -2557 425
rect -2591 323 -2557 357
rect -2591 255 -2557 289
rect -2591 187 -2557 221
rect -2591 119 -2557 153
rect -2591 51 -2557 85
rect -2591 -17 -2557 17
rect -2591 -85 -2557 -51
rect -2591 -153 -2557 -119
rect -2591 -221 -2557 -187
rect -2591 -289 -2557 -255
rect -2591 -357 -2557 -323
rect -2591 -425 -2557 -391
rect -2591 -493 -2557 -459
rect -2591 -561 -2557 -527
rect -1733 527 -1699 561
rect -1733 459 -1699 493
rect -1733 391 -1699 425
rect -1733 323 -1699 357
rect -1733 255 -1699 289
rect -1733 187 -1699 221
rect -1733 119 -1699 153
rect -1733 51 -1699 85
rect -1733 -17 -1699 17
rect -1733 -85 -1699 -51
rect -1733 -153 -1699 -119
rect -1733 -221 -1699 -187
rect -1733 -289 -1699 -255
rect -1733 -357 -1699 -323
rect -1733 -425 -1699 -391
rect -1733 -493 -1699 -459
rect -1733 -561 -1699 -527
rect -875 527 -841 561
rect -875 459 -841 493
rect -875 391 -841 425
rect -875 323 -841 357
rect -875 255 -841 289
rect -875 187 -841 221
rect -875 119 -841 153
rect -875 51 -841 85
rect -875 -17 -841 17
rect -875 -85 -841 -51
rect -875 -153 -841 -119
rect -875 -221 -841 -187
rect -875 -289 -841 -255
rect -875 -357 -841 -323
rect -875 -425 -841 -391
rect -875 -493 -841 -459
rect -875 -561 -841 -527
rect -17 527 17 561
rect -17 459 17 493
rect -17 391 17 425
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect -17 -425 17 -391
rect -17 -493 17 -459
rect -17 -561 17 -527
rect 841 527 875 561
rect 841 459 875 493
rect 841 391 875 425
rect 841 323 875 357
rect 841 255 875 289
rect 841 187 875 221
rect 841 119 875 153
rect 841 51 875 85
rect 841 -17 875 17
rect 841 -85 875 -51
rect 841 -153 875 -119
rect 841 -221 875 -187
rect 841 -289 875 -255
rect 841 -357 875 -323
rect 841 -425 875 -391
rect 841 -493 875 -459
rect 841 -561 875 -527
rect 1699 527 1733 561
rect 1699 459 1733 493
rect 1699 391 1733 425
rect 1699 323 1733 357
rect 1699 255 1733 289
rect 1699 187 1733 221
rect 1699 119 1733 153
rect 1699 51 1733 85
rect 1699 -17 1733 17
rect 1699 -85 1733 -51
rect 1699 -153 1733 -119
rect 1699 -221 1733 -187
rect 1699 -289 1733 -255
rect 1699 -357 1733 -323
rect 1699 -425 1733 -391
rect 1699 -493 1733 -459
rect 1699 -561 1733 -527
rect 2557 527 2591 561
rect 2557 459 2591 493
rect 2557 391 2591 425
rect 2557 323 2591 357
rect 2557 255 2591 289
rect 2557 187 2591 221
rect 2557 119 2591 153
rect 2557 51 2591 85
rect 2557 -17 2591 17
rect 2557 -85 2591 -51
rect 2557 -153 2591 -119
rect 2557 -221 2591 -187
rect 2557 -289 2591 -255
rect 2557 -357 2591 -323
rect 2557 -425 2591 -391
rect 2557 -493 2591 -459
rect 2557 -561 2591 -527
rect 3415 527 3449 561
rect 3415 459 3449 493
rect 3415 391 3449 425
rect 3415 323 3449 357
rect 3415 255 3449 289
rect 3415 187 3449 221
rect 3415 119 3449 153
rect 3415 51 3449 85
rect 3415 -17 3449 17
rect 3415 -85 3449 -51
rect 3415 -153 3449 -119
rect 3415 -221 3449 -187
rect 3415 -289 3449 -255
rect 3415 -357 3449 -323
rect 3415 -425 3449 -391
rect 3415 -493 3449 -459
rect 3415 -561 3449 -527
rect 4273 527 4307 561
rect 4273 459 4307 493
rect 4273 391 4307 425
rect 4273 323 4307 357
rect 4273 255 4307 289
rect 4273 187 4307 221
rect 4273 119 4307 153
rect 4273 51 4307 85
rect 4273 -17 4307 17
rect 4273 -85 4307 -51
rect 4273 -153 4307 -119
rect 4273 -221 4307 -187
rect 4273 -289 4307 -255
rect 4273 -357 4307 -323
rect 4273 -425 4307 -391
rect 4273 -493 4307 -459
rect 4273 -561 4307 -527
rect 5131 527 5165 561
rect 5131 459 5165 493
rect 5131 391 5165 425
rect 5131 323 5165 357
rect 5131 255 5165 289
rect 5131 187 5165 221
rect 5131 119 5165 153
rect 5131 51 5165 85
rect 5131 -17 5165 17
rect 5131 -85 5165 -51
rect 5131 -153 5165 -119
rect 5131 -221 5165 -187
rect 5131 -289 5165 -255
rect 5131 -357 5165 -323
rect 5131 -425 5165 -391
rect 5131 -493 5165 -459
rect 5131 -561 5165 -527
rect 5989 527 6023 561
rect 5989 459 6023 493
rect 5989 391 6023 425
rect 5989 323 6023 357
rect 5989 255 6023 289
rect 5989 187 6023 221
rect 5989 119 6023 153
rect 5989 51 6023 85
rect 5989 -17 6023 17
rect 5989 -85 6023 -51
rect 5989 -153 6023 -119
rect 5989 -221 6023 -187
rect 5989 -289 6023 -255
rect 5989 -357 6023 -323
rect 5989 -425 6023 -391
rect 5989 -493 6023 -459
rect 5989 -561 6023 -527
<< poly >>
rect -5823 681 -5331 697
rect -5823 664 -5798 681
rect -5977 647 -5798 664
rect -5764 647 -5730 681
rect -5696 647 -5662 681
rect -5628 647 -5594 681
rect -5560 647 -5526 681
rect -5492 647 -5458 681
rect -5424 647 -5390 681
rect -5356 664 -5331 681
rect -4965 681 -4473 697
rect -4965 664 -4940 681
rect -5356 647 -5177 664
rect -5977 600 -5177 647
rect -5119 647 -4940 664
rect -4906 647 -4872 681
rect -4838 647 -4804 681
rect -4770 647 -4736 681
rect -4702 647 -4668 681
rect -4634 647 -4600 681
rect -4566 647 -4532 681
rect -4498 664 -4473 681
rect -4107 681 -3615 697
rect -4107 664 -4082 681
rect -4498 647 -4319 664
rect -5119 600 -4319 647
rect -4261 647 -4082 664
rect -4048 647 -4014 681
rect -3980 647 -3946 681
rect -3912 647 -3878 681
rect -3844 647 -3810 681
rect -3776 647 -3742 681
rect -3708 647 -3674 681
rect -3640 664 -3615 681
rect -3249 681 -2757 697
rect -3249 664 -3224 681
rect -3640 647 -3461 664
rect -4261 600 -3461 647
rect -3403 647 -3224 664
rect -3190 647 -3156 681
rect -3122 647 -3088 681
rect -3054 647 -3020 681
rect -2986 647 -2952 681
rect -2918 647 -2884 681
rect -2850 647 -2816 681
rect -2782 664 -2757 681
rect -2391 681 -1899 697
rect -2391 664 -2366 681
rect -2782 647 -2603 664
rect -3403 600 -2603 647
rect -2545 647 -2366 664
rect -2332 647 -2298 681
rect -2264 647 -2230 681
rect -2196 647 -2162 681
rect -2128 647 -2094 681
rect -2060 647 -2026 681
rect -1992 647 -1958 681
rect -1924 664 -1899 681
rect -1533 681 -1041 697
rect -1533 664 -1508 681
rect -1924 647 -1745 664
rect -2545 600 -1745 647
rect -1687 647 -1508 664
rect -1474 647 -1440 681
rect -1406 647 -1372 681
rect -1338 647 -1304 681
rect -1270 647 -1236 681
rect -1202 647 -1168 681
rect -1134 647 -1100 681
rect -1066 664 -1041 681
rect -675 681 -183 697
rect -675 664 -650 681
rect -1066 647 -887 664
rect -1687 600 -887 647
rect -829 647 -650 664
rect -616 647 -582 681
rect -548 647 -514 681
rect -480 647 -446 681
rect -412 647 -378 681
rect -344 647 -310 681
rect -276 647 -242 681
rect -208 664 -183 681
rect 183 681 675 697
rect 183 664 208 681
rect -208 647 -29 664
rect -829 600 -29 647
rect 29 647 208 664
rect 242 647 276 681
rect 310 647 344 681
rect 378 647 412 681
rect 446 647 480 681
rect 514 647 548 681
rect 582 647 616 681
rect 650 664 675 681
rect 1041 681 1533 697
rect 1041 664 1066 681
rect 650 647 829 664
rect 29 600 829 647
rect 887 647 1066 664
rect 1100 647 1134 681
rect 1168 647 1202 681
rect 1236 647 1270 681
rect 1304 647 1338 681
rect 1372 647 1406 681
rect 1440 647 1474 681
rect 1508 664 1533 681
rect 1899 681 2391 697
rect 1899 664 1924 681
rect 1508 647 1687 664
rect 887 600 1687 647
rect 1745 647 1924 664
rect 1958 647 1992 681
rect 2026 647 2060 681
rect 2094 647 2128 681
rect 2162 647 2196 681
rect 2230 647 2264 681
rect 2298 647 2332 681
rect 2366 664 2391 681
rect 2757 681 3249 697
rect 2757 664 2782 681
rect 2366 647 2545 664
rect 1745 600 2545 647
rect 2603 647 2782 664
rect 2816 647 2850 681
rect 2884 647 2918 681
rect 2952 647 2986 681
rect 3020 647 3054 681
rect 3088 647 3122 681
rect 3156 647 3190 681
rect 3224 664 3249 681
rect 3615 681 4107 697
rect 3615 664 3640 681
rect 3224 647 3403 664
rect 2603 600 3403 647
rect 3461 647 3640 664
rect 3674 647 3708 681
rect 3742 647 3776 681
rect 3810 647 3844 681
rect 3878 647 3912 681
rect 3946 647 3980 681
rect 4014 647 4048 681
rect 4082 664 4107 681
rect 4473 681 4965 697
rect 4473 664 4498 681
rect 4082 647 4261 664
rect 3461 600 4261 647
rect 4319 647 4498 664
rect 4532 647 4566 681
rect 4600 647 4634 681
rect 4668 647 4702 681
rect 4736 647 4770 681
rect 4804 647 4838 681
rect 4872 647 4906 681
rect 4940 664 4965 681
rect 5331 681 5823 697
rect 5331 664 5356 681
rect 4940 647 5119 664
rect 4319 600 5119 647
rect 5177 647 5356 664
rect 5390 647 5424 681
rect 5458 647 5492 681
rect 5526 647 5560 681
rect 5594 647 5628 681
rect 5662 647 5696 681
rect 5730 647 5764 681
rect 5798 664 5823 681
rect 5798 647 5977 664
rect 5177 600 5977 647
rect -5977 -647 -5177 -600
rect -5977 -664 -5798 -647
rect -5823 -681 -5798 -664
rect -5764 -681 -5730 -647
rect -5696 -681 -5662 -647
rect -5628 -681 -5594 -647
rect -5560 -681 -5526 -647
rect -5492 -681 -5458 -647
rect -5424 -681 -5390 -647
rect -5356 -664 -5177 -647
rect -5119 -647 -4319 -600
rect -5119 -664 -4940 -647
rect -5356 -681 -5331 -664
rect -5823 -697 -5331 -681
rect -4965 -681 -4940 -664
rect -4906 -681 -4872 -647
rect -4838 -681 -4804 -647
rect -4770 -681 -4736 -647
rect -4702 -681 -4668 -647
rect -4634 -681 -4600 -647
rect -4566 -681 -4532 -647
rect -4498 -664 -4319 -647
rect -4261 -647 -3461 -600
rect -4261 -664 -4082 -647
rect -4498 -681 -4473 -664
rect -4965 -697 -4473 -681
rect -4107 -681 -4082 -664
rect -4048 -681 -4014 -647
rect -3980 -681 -3946 -647
rect -3912 -681 -3878 -647
rect -3844 -681 -3810 -647
rect -3776 -681 -3742 -647
rect -3708 -681 -3674 -647
rect -3640 -664 -3461 -647
rect -3403 -647 -2603 -600
rect -3403 -664 -3224 -647
rect -3640 -681 -3615 -664
rect -4107 -697 -3615 -681
rect -3249 -681 -3224 -664
rect -3190 -681 -3156 -647
rect -3122 -681 -3088 -647
rect -3054 -681 -3020 -647
rect -2986 -681 -2952 -647
rect -2918 -681 -2884 -647
rect -2850 -681 -2816 -647
rect -2782 -664 -2603 -647
rect -2545 -647 -1745 -600
rect -2545 -664 -2366 -647
rect -2782 -681 -2757 -664
rect -3249 -697 -2757 -681
rect -2391 -681 -2366 -664
rect -2332 -681 -2298 -647
rect -2264 -681 -2230 -647
rect -2196 -681 -2162 -647
rect -2128 -681 -2094 -647
rect -2060 -681 -2026 -647
rect -1992 -681 -1958 -647
rect -1924 -664 -1745 -647
rect -1687 -647 -887 -600
rect -1687 -664 -1508 -647
rect -1924 -681 -1899 -664
rect -2391 -697 -1899 -681
rect -1533 -681 -1508 -664
rect -1474 -681 -1440 -647
rect -1406 -681 -1372 -647
rect -1338 -681 -1304 -647
rect -1270 -681 -1236 -647
rect -1202 -681 -1168 -647
rect -1134 -681 -1100 -647
rect -1066 -664 -887 -647
rect -829 -647 -29 -600
rect -829 -664 -650 -647
rect -1066 -681 -1041 -664
rect -1533 -697 -1041 -681
rect -675 -681 -650 -664
rect -616 -681 -582 -647
rect -548 -681 -514 -647
rect -480 -681 -446 -647
rect -412 -681 -378 -647
rect -344 -681 -310 -647
rect -276 -681 -242 -647
rect -208 -664 -29 -647
rect 29 -647 829 -600
rect 29 -664 208 -647
rect -208 -681 -183 -664
rect -675 -697 -183 -681
rect 183 -681 208 -664
rect 242 -681 276 -647
rect 310 -681 344 -647
rect 378 -681 412 -647
rect 446 -681 480 -647
rect 514 -681 548 -647
rect 582 -681 616 -647
rect 650 -664 829 -647
rect 887 -647 1687 -600
rect 887 -664 1066 -647
rect 650 -681 675 -664
rect 183 -697 675 -681
rect 1041 -681 1066 -664
rect 1100 -681 1134 -647
rect 1168 -681 1202 -647
rect 1236 -681 1270 -647
rect 1304 -681 1338 -647
rect 1372 -681 1406 -647
rect 1440 -681 1474 -647
rect 1508 -664 1687 -647
rect 1745 -647 2545 -600
rect 1745 -664 1924 -647
rect 1508 -681 1533 -664
rect 1041 -697 1533 -681
rect 1899 -681 1924 -664
rect 1958 -681 1992 -647
rect 2026 -681 2060 -647
rect 2094 -681 2128 -647
rect 2162 -681 2196 -647
rect 2230 -681 2264 -647
rect 2298 -681 2332 -647
rect 2366 -664 2545 -647
rect 2603 -647 3403 -600
rect 2603 -664 2782 -647
rect 2366 -681 2391 -664
rect 1899 -697 2391 -681
rect 2757 -681 2782 -664
rect 2816 -681 2850 -647
rect 2884 -681 2918 -647
rect 2952 -681 2986 -647
rect 3020 -681 3054 -647
rect 3088 -681 3122 -647
rect 3156 -681 3190 -647
rect 3224 -664 3403 -647
rect 3461 -647 4261 -600
rect 3461 -664 3640 -647
rect 3224 -681 3249 -664
rect 2757 -697 3249 -681
rect 3615 -681 3640 -664
rect 3674 -681 3708 -647
rect 3742 -681 3776 -647
rect 3810 -681 3844 -647
rect 3878 -681 3912 -647
rect 3946 -681 3980 -647
rect 4014 -681 4048 -647
rect 4082 -664 4261 -647
rect 4319 -647 5119 -600
rect 4319 -664 4498 -647
rect 4082 -681 4107 -664
rect 3615 -697 4107 -681
rect 4473 -681 4498 -664
rect 4532 -681 4566 -647
rect 4600 -681 4634 -647
rect 4668 -681 4702 -647
rect 4736 -681 4770 -647
rect 4804 -681 4838 -647
rect 4872 -681 4906 -647
rect 4940 -664 5119 -647
rect 5177 -647 5977 -600
rect 5177 -664 5356 -647
rect 4940 -681 4965 -664
rect 4473 -697 4965 -681
rect 5331 -681 5356 -664
rect 5390 -681 5424 -647
rect 5458 -681 5492 -647
rect 5526 -681 5560 -647
rect 5594 -681 5628 -647
rect 5662 -681 5696 -647
rect 5730 -681 5764 -647
rect 5798 -664 5977 -647
rect 5798 -681 5823 -664
rect 5331 -697 5823 -681
<< polycont >>
rect -5798 647 -5764 681
rect -5730 647 -5696 681
rect -5662 647 -5628 681
rect -5594 647 -5560 681
rect -5526 647 -5492 681
rect -5458 647 -5424 681
rect -5390 647 -5356 681
rect -4940 647 -4906 681
rect -4872 647 -4838 681
rect -4804 647 -4770 681
rect -4736 647 -4702 681
rect -4668 647 -4634 681
rect -4600 647 -4566 681
rect -4532 647 -4498 681
rect -4082 647 -4048 681
rect -4014 647 -3980 681
rect -3946 647 -3912 681
rect -3878 647 -3844 681
rect -3810 647 -3776 681
rect -3742 647 -3708 681
rect -3674 647 -3640 681
rect -3224 647 -3190 681
rect -3156 647 -3122 681
rect -3088 647 -3054 681
rect -3020 647 -2986 681
rect -2952 647 -2918 681
rect -2884 647 -2850 681
rect -2816 647 -2782 681
rect -2366 647 -2332 681
rect -2298 647 -2264 681
rect -2230 647 -2196 681
rect -2162 647 -2128 681
rect -2094 647 -2060 681
rect -2026 647 -1992 681
rect -1958 647 -1924 681
rect -1508 647 -1474 681
rect -1440 647 -1406 681
rect -1372 647 -1338 681
rect -1304 647 -1270 681
rect -1236 647 -1202 681
rect -1168 647 -1134 681
rect -1100 647 -1066 681
rect -650 647 -616 681
rect -582 647 -548 681
rect -514 647 -480 681
rect -446 647 -412 681
rect -378 647 -344 681
rect -310 647 -276 681
rect -242 647 -208 681
rect 208 647 242 681
rect 276 647 310 681
rect 344 647 378 681
rect 412 647 446 681
rect 480 647 514 681
rect 548 647 582 681
rect 616 647 650 681
rect 1066 647 1100 681
rect 1134 647 1168 681
rect 1202 647 1236 681
rect 1270 647 1304 681
rect 1338 647 1372 681
rect 1406 647 1440 681
rect 1474 647 1508 681
rect 1924 647 1958 681
rect 1992 647 2026 681
rect 2060 647 2094 681
rect 2128 647 2162 681
rect 2196 647 2230 681
rect 2264 647 2298 681
rect 2332 647 2366 681
rect 2782 647 2816 681
rect 2850 647 2884 681
rect 2918 647 2952 681
rect 2986 647 3020 681
rect 3054 647 3088 681
rect 3122 647 3156 681
rect 3190 647 3224 681
rect 3640 647 3674 681
rect 3708 647 3742 681
rect 3776 647 3810 681
rect 3844 647 3878 681
rect 3912 647 3946 681
rect 3980 647 4014 681
rect 4048 647 4082 681
rect 4498 647 4532 681
rect 4566 647 4600 681
rect 4634 647 4668 681
rect 4702 647 4736 681
rect 4770 647 4804 681
rect 4838 647 4872 681
rect 4906 647 4940 681
rect 5356 647 5390 681
rect 5424 647 5458 681
rect 5492 647 5526 681
rect 5560 647 5594 681
rect 5628 647 5662 681
rect 5696 647 5730 681
rect 5764 647 5798 681
rect -5798 -681 -5764 -647
rect -5730 -681 -5696 -647
rect -5662 -681 -5628 -647
rect -5594 -681 -5560 -647
rect -5526 -681 -5492 -647
rect -5458 -681 -5424 -647
rect -5390 -681 -5356 -647
rect -4940 -681 -4906 -647
rect -4872 -681 -4838 -647
rect -4804 -681 -4770 -647
rect -4736 -681 -4702 -647
rect -4668 -681 -4634 -647
rect -4600 -681 -4566 -647
rect -4532 -681 -4498 -647
rect -4082 -681 -4048 -647
rect -4014 -681 -3980 -647
rect -3946 -681 -3912 -647
rect -3878 -681 -3844 -647
rect -3810 -681 -3776 -647
rect -3742 -681 -3708 -647
rect -3674 -681 -3640 -647
rect -3224 -681 -3190 -647
rect -3156 -681 -3122 -647
rect -3088 -681 -3054 -647
rect -3020 -681 -2986 -647
rect -2952 -681 -2918 -647
rect -2884 -681 -2850 -647
rect -2816 -681 -2782 -647
rect -2366 -681 -2332 -647
rect -2298 -681 -2264 -647
rect -2230 -681 -2196 -647
rect -2162 -681 -2128 -647
rect -2094 -681 -2060 -647
rect -2026 -681 -1992 -647
rect -1958 -681 -1924 -647
rect -1508 -681 -1474 -647
rect -1440 -681 -1406 -647
rect -1372 -681 -1338 -647
rect -1304 -681 -1270 -647
rect -1236 -681 -1202 -647
rect -1168 -681 -1134 -647
rect -1100 -681 -1066 -647
rect -650 -681 -616 -647
rect -582 -681 -548 -647
rect -514 -681 -480 -647
rect -446 -681 -412 -647
rect -378 -681 -344 -647
rect -310 -681 -276 -647
rect -242 -681 -208 -647
rect 208 -681 242 -647
rect 276 -681 310 -647
rect 344 -681 378 -647
rect 412 -681 446 -647
rect 480 -681 514 -647
rect 548 -681 582 -647
rect 616 -681 650 -647
rect 1066 -681 1100 -647
rect 1134 -681 1168 -647
rect 1202 -681 1236 -647
rect 1270 -681 1304 -647
rect 1338 -681 1372 -647
rect 1406 -681 1440 -647
rect 1474 -681 1508 -647
rect 1924 -681 1958 -647
rect 1992 -681 2026 -647
rect 2060 -681 2094 -647
rect 2128 -681 2162 -647
rect 2196 -681 2230 -647
rect 2264 -681 2298 -647
rect 2332 -681 2366 -647
rect 2782 -681 2816 -647
rect 2850 -681 2884 -647
rect 2918 -681 2952 -647
rect 2986 -681 3020 -647
rect 3054 -681 3088 -647
rect 3122 -681 3156 -647
rect 3190 -681 3224 -647
rect 3640 -681 3674 -647
rect 3708 -681 3742 -647
rect 3776 -681 3810 -647
rect 3844 -681 3878 -647
rect 3912 -681 3946 -647
rect 3980 -681 4014 -647
rect 4048 -681 4082 -647
rect 4498 -681 4532 -647
rect 4566 -681 4600 -647
rect 4634 -681 4668 -647
rect 4702 -681 4736 -647
rect 4770 -681 4804 -647
rect 4838 -681 4872 -647
rect 4906 -681 4940 -647
rect 5356 -681 5390 -647
rect 5424 -681 5458 -647
rect 5492 -681 5526 -647
rect 5560 -681 5594 -647
rect 5628 -681 5662 -647
rect 5696 -681 5730 -647
rect 5764 -681 5798 -647
<< locali >>
rect -5823 647 -5798 681
rect -5764 647 -5738 681
rect -5696 647 -5666 681
rect -5628 647 -5594 681
rect -5560 647 -5526 681
rect -5488 647 -5458 681
rect -5416 647 -5390 681
rect -5356 647 -5331 681
rect -4965 647 -4940 681
rect -4906 647 -4880 681
rect -4838 647 -4808 681
rect -4770 647 -4736 681
rect -4702 647 -4668 681
rect -4630 647 -4600 681
rect -4558 647 -4532 681
rect -4498 647 -4473 681
rect -4107 647 -4082 681
rect -4048 647 -4022 681
rect -3980 647 -3950 681
rect -3912 647 -3878 681
rect -3844 647 -3810 681
rect -3772 647 -3742 681
rect -3700 647 -3674 681
rect -3640 647 -3615 681
rect -3249 647 -3224 681
rect -3190 647 -3164 681
rect -3122 647 -3092 681
rect -3054 647 -3020 681
rect -2986 647 -2952 681
rect -2914 647 -2884 681
rect -2842 647 -2816 681
rect -2782 647 -2757 681
rect -2391 647 -2366 681
rect -2332 647 -2306 681
rect -2264 647 -2234 681
rect -2196 647 -2162 681
rect -2128 647 -2094 681
rect -2056 647 -2026 681
rect -1984 647 -1958 681
rect -1924 647 -1899 681
rect -1533 647 -1508 681
rect -1474 647 -1448 681
rect -1406 647 -1376 681
rect -1338 647 -1304 681
rect -1270 647 -1236 681
rect -1198 647 -1168 681
rect -1126 647 -1100 681
rect -1066 647 -1041 681
rect -675 647 -650 681
rect -616 647 -590 681
rect -548 647 -518 681
rect -480 647 -446 681
rect -412 647 -378 681
rect -340 647 -310 681
rect -268 647 -242 681
rect -208 647 -183 681
rect 183 647 208 681
rect 242 647 268 681
rect 310 647 340 681
rect 378 647 412 681
rect 446 647 480 681
rect 518 647 548 681
rect 590 647 616 681
rect 650 647 675 681
rect 1041 647 1066 681
rect 1100 647 1126 681
rect 1168 647 1198 681
rect 1236 647 1270 681
rect 1304 647 1338 681
rect 1376 647 1406 681
rect 1448 647 1474 681
rect 1508 647 1533 681
rect 1899 647 1924 681
rect 1958 647 1984 681
rect 2026 647 2056 681
rect 2094 647 2128 681
rect 2162 647 2196 681
rect 2234 647 2264 681
rect 2306 647 2332 681
rect 2366 647 2391 681
rect 2757 647 2782 681
rect 2816 647 2842 681
rect 2884 647 2914 681
rect 2952 647 2986 681
rect 3020 647 3054 681
rect 3092 647 3122 681
rect 3164 647 3190 681
rect 3224 647 3249 681
rect 3615 647 3640 681
rect 3674 647 3700 681
rect 3742 647 3772 681
rect 3810 647 3844 681
rect 3878 647 3912 681
rect 3950 647 3980 681
rect 4022 647 4048 681
rect 4082 647 4107 681
rect 4473 647 4498 681
rect 4532 647 4558 681
rect 4600 647 4630 681
rect 4668 647 4702 681
rect 4736 647 4770 681
rect 4808 647 4838 681
rect 4880 647 4906 681
rect 4940 647 4965 681
rect 5331 647 5356 681
rect 5390 647 5416 681
rect 5458 647 5488 681
rect 5526 647 5560 681
rect 5594 647 5628 681
rect 5666 647 5696 681
rect 5738 647 5764 681
rect 5798 647 5823 681
rect -6023 561 -5989 604
rect -6023 493 -5989 523
rect -6023 425 -5989 451
rect -6023 357 -5989 379
rect -6023 289 -5989 307
rect -6023 221 -5989 235
rect -6023 153 -5989 163
rect -6023 85 -5989 91
rect -6023 17 -5989 19
rect -6023 -19 -5989 -17
rect -6023 -91 -5989 -85
rect -6023 -163 -5989 -153
rect -6023 -235 -5989 -221
rect -6023 -307 -5989 -289
rect -6023 -379 -5989 -357
rect -6023 -451 -5989 -425
rect -6023 -523 -5989 -493
rect -6023 -604 -5989 -561
rect -5165 561 -5131 604
rect -5165 493 -5131 523
rect -5165 425 -5131 451
rect -5165 357 -5131 379
rect -5165 289 -5131 307
rect -5165 221 -5131 235
rect -5165 153 -5131 163
rect -5165 85 -5131 91
rect -5165 17 -5131 19
rect -5165 -19 -5131 -17
rect -5165 -91 -5131 -85
rect -5165 -163 -5131 -153
rect -5165 -235 -5131 -221
rect -5165 -307 -5131 -289
rect -5165 -379 -5131 -357
rect -5165 -451 -5131 -425
rect -5165 -523 -5131 -493
rect -5165 -604 -5131 -561
rect -4307 561 -4273 604
rect -4307 493 -4273 523
rect -4307 425 -4273 451
rect -4307 357 -4273 379
rect -4307 289 -4273 307
rect -4307 221 -4273 235
rect -4307 153 -4273 163
rect -4307 85 -4273 91
rect -4307 17 -4273 19
rect -4307 -19 -4273 -17
rect -4307 -91 -4273 -85
rect -4307 -163 -4273 -153
rect -4307 -235 -4273 -221
rect -4307 -307 -4273 -289
rect -4307 -379 -4273 -357
rect -4307 -451 -4273 -425
rect -4307 -523 -4273 -493
rect -4307 -604 -4273 -561
rect -3449 561 -3415 604
rect -3449 493 -3415 523
rect -3449 425 -3415 451
rect -3449 357 -3415 379
rect -3449 289 -3415 307
rect -3449 221 -3415 235
rect -3449 153 -3415 163
rect -3449 85 -3415 91
rect -3449 17 -3415 19
rect -3449 -19 -3415 -17
rect -3449 -91 -3415 -85
rect -3449 -163 -3415 -153
rect -3449 -235 -3415 -221
rect -3449 -307 -3415 -289
rect -3449 -379 -3415 -357
rect -3449 -451 -3415 -425
rect -3449 -523 -3415 -493
rect -3449 -604 -3415 -561
rect -2591 561 -2557 604
rect -2591 493 -2557 523
rect -2591 425 -2557 451
rect -2591 357 -2557 379
rect -2591 289 -2557 307
rect -2591 221 -2557 235
rect -2591 153 -2557 163
rect -2591 85 -2557 91
rect -2591 17 -2557 19
rect -2591 -19 -2557 -17
rect -2591 -91 -2557 -85
rect -2591 -163 -2557 -153
rect -2591 -235 -2557 -221
rect -2591 -307 -2557 -289
rect -2591 -379 -2557 -357
rect -2591 -451 -2557 -425
rect -2591 -523 -2557 -493
rect -2591 -604 -2557 -561
rect -1733 561 -1699 604
rect -1733 493 -1699 523
rect -1733 425 -1699 451
rect -1733 357 -1699 379
rect -1733 289 -1699 307
rect -1733 221 -1699 235
rect -1733 153 -1699 163
rect -1733 85 -1699 91
rect -1733 17 -1699 19
rect -1733 -19 -1699 -17
rect -1733 -91 -1699 -85
rect -1733 -163 -1699 -153
rect -1733 -235 -1699 -221
rect -1733 -307 -1699 -289
rect -1733 -379 -1699 -357
rect -1733 -451 -1699 -425
rect -1733 -523 -1699 -493
rect -1733 -604 -1699 -561
rect -875 561 -841 604
rect -875 493 -841 523
rect -875 425 -841 451
rect -875 357 -841 379
rect -875 289 -841 307
rect -875 221 -841 235
rect -875 153 -841 163
rect -875 85 -841 91
rect -875 17 -841 19
rect -875 -19 -841 -17
rect -875 -91 -841 -85
rect -875 -163 -841 -153
rect -875 -235 -841 -221
rect -875 -307 -841 -289
rect -875 -379 -841 -357
rect -875 -451 -841 -425
rect -875 -523 -841 -493
rect -875 -604 -841 -561
rect -17 561 17 604
rect -17 493 17 523
rect -17 425 17 451
rect -17 357 17 379
rect -17 289 17 307
rect -17 221 17 235
rect -17 153 17 163
rect -17 85 17 91
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -91 17 -85
rect -17 -163 17 -153
rect -17 -235 17 -221
rect -17 -307 17 -289
rect -17 -379 17 -357
rect -17 -451 17 -425
rect -17 -523 17 -493
rect -17 -604 17 -561
rect 841 561 875 604
rect 841 493 875 523
rect 841 425 875 451
rect 841 357 875 379
rect 841 289 875 307
rect 841 221 875 235
rect 841 153 875 163
rect 841 85 875 91
rect 841 17 875 19
rect 841 -19 875 -17
rect 841 -91 875 -85
rect 841 -163 875 -153
rect 841 -235 875 -221
rect 841 -307 875 -289
rect 841 -379 875 -357
rect 841 -451 875 -425
rect 841 -523 875 -493
rect 841 -604 875 -561
rect 1699 561 1733 604
rect 1699 493 1733 523
rect 1699 425 1733 451
rect 1699 357 1733 379
rect 1699 289 1733 307
rect 1699 221 1733 235
rect 1699 153 1733 163
rect 1699 85 1733 91
rect 1699 17 1733 19
rect 1699 -19 1733 -17
rect 1699 -91 1733 -85
rect 1699 -163 1733 -153
rect 1699 -235 1733 -221
rect 1699 -307 1733 -289
rect 1699 -379 1733 -357
rect 1699 -451 1733 -425
rect 1699 -523 1733 -493
rect 1699 -604 1733 -561
rect 2557 561 2591 604
rect 2557 493 2591 523
rect 2557 425 2591 451
rect 2557 357 2591 379
rect 2557 289 2591 307
rect 2557 221 2591 235
rect 2557 153 2591 163
rect 2557 85 2591 91
rect 2557 17 2591 19
rect 2557 -19 2591 -17
rect 2557 -91 2591 -85
rect 2557 -163 2591 -153
rect 2557 -235 2591 -221
rect 2557 -307 2591 -289
rect 2557 -379 2591 -357
rect 2557 -451 2591 -425
rect 2557 -523 2591 -493
rect 2557 -604 2591 -561
rect 3415 561 3449 604
rect 3415 493 3449 523
rect 3415 425 3449 451
rect 3415 357 3449 379
rect 3415 289 3449 307
rect 3415 221 3449 235
rect 3415 153 3449 163
rect 3415 85 3449 91
rect 3415 17 3449 19
rect 3415 -19 3449 -17
rect 3415 -91 3449 -85
rect 3415 -163 3449 -153
rect 3415 -235 3449 -221
rect 3415 -307 3449 -289
rect 3415 -379 3449 -357
rect 3415 -451 3449 -425
rect 3415 -523 3449 -493
rect 3415 -604 3449 -561
rect 4273 561 4307 604
rect 4273 493 4307 523
rect 4273 425 4307 451
rect 4273 357 4307 379
rect 4273 289 4307 307
rect 4273 221 4307 235
rect 4273 153 4307 163
rect 4273 85 4307 91
rect 4273 17 4307 19
rect 4273 -19 4307 -17
rect 4273 -91 4307 -85
rect 4273 -163 4307 -153
rect 4273 -235 4307 -221
rect 4273 -307 4307 -289
rect 4273 -379 4307 -357
rect 4273 -451 4307 -425
rect 4273 -523 4307 -493
rect 4273 -604 4307 -561
rect 5131 561 5165 604
rect 5131 493 5165 523
rect 5131 425 5165 451
rect 5131 357 5165 379
rect 5131 289 5165 307
rect 5131 221 5165 235
rect 5131 153 5165 163
rect 5131 85 5165 91
rect 5131 17 5165 19
rect 5131 -19 5165 -17
rect 5131 -91 5165 -85
rect 5131 -163 5165 -153
rect 5131 -235 5165 -221
rect 5131 -307 5165 -289
rect 5131 -379 5165 -357
rect 5131 -451 5165 -425
rect 5131 -523 5165 -493
rect 5131 -604 5165 -561
rect 5989 561 6023 604
rect 5989 493 6023 523
rect 5989 425 6023 451
rect 5989 357 6023 379
rect 5989 289 6023 307
rect 5989 221 6023 235
rect 5989 153 6023 163
rect 5989 85 6023 91
rect 5989 17 6023 19
rect 5989 -19 6023 -17
rect 5989 -91 6023 -85
rect 5989 -163 6023 -153
rect 5989 -235 6023 -221
rect 5989 -307 6023 -289
rect 5989 -379 6023 -357
rect 5989 -451 6023 -425
rect 5989 -523 6023 -493
rect 5989 -604 6023 -561
rect -5823 -681 -5798 -647
rect -5764 -681 -5738 -647
rect -5696 -681 -5666 -647
rect -5628 -681 -5594 -647
rect -5560 -681 -5526 -647
rect -5488 -681 -5458 -647
rect -5416 -681 -5390 -647
rect -5356 -681 -5331 -647
rect -4965 -681 -4940 -647
rect -4906 -681 -4880 -647
rect -4838 -681 -4808 -647
rect -4770 -681 -4736 -647
rect -4702 -681 -4668 -647
rect -4630 -681 -4600 -647
rect -4558 -681 -4532 -647
rect -4498 -681 -4473 -647
rect -4107 -681 -4082 -647
rect -4048 -681 -4022 -647
rect -3980 -681 -3950 -647
rect -3912 -681 -3878 -647
rect -3844 -681 -3810 -647
rect -3772 -681 -3742 -647
rect -3700 -681 -3674 -647
rect -3640 -681 -3615 -647
rect -3249 -681 -3224 -647
rect -3190 -681 -3164 -647
rect -3122 -681 -3092 -647
rect -3054 -681 -3020 -647
rect -2986 -681 -2952 -647
rect -2914 -681 -2884 -647
rect -2842 -681 -2816 -647
rect -2782 -681 -2757 -647
rect -2391 -681 -2366 -647
rect -2332 -681 -2306 -647
rect -2264 -681 -2234 -647
rect -2196 -681 -2162 -647
rect -2128 -681 -2094 -647
rect -2056 -681 -2026 -647
rect -1984 -681 -1958 -647
rect -1924 -681 -1899 -647
rect -1533 -681 -1508 -647
rect -1474 -681 -1448 -647
rect -1406 -681 -1376 -647
rect -1338 -681 -1304 -647
rect -1270 -681 -1236 -647
rect -1198 -681 -1168 -647
rect -1126 -681 -1100 -647
rect -1066 -681 -1041 -647
rect -675 -681 -650 -647
rect -616 -681 -590 -647
rect -548 -681 -518 -647
rect -480 -681 -446 -647
rect -412 -681 -378 -647
rect -340 -681 -310 -647
rect -268 -681 -242 -647
rect -208 -681 -183 -647
rect 183 -681 208 -647
rect 242 -681 268 -647
rect 310 -681 340 -647
rect 378 -681 412 -647
rect 446 -681 480 -647
rect 518 -681 548 -647
rect 590 -681 616 -647
rect 650 -681 675 -647
rect 1041 -681 1066 -647
rect 1100 -681 1126 -647
rect 1168 -681 1198 -647
rect 1236 -681 1270 -647
rect 1304 -681 1338 -647
rect 1376 -681 1406 -647
rect 1448 -681 1474 -647
rect 1508 -681 1533 -647
rect 1899 -681 1924 -647
rect 1958 -681 1984 -647
rect 2026 -681 2056 -647
rect 2094 -681 2128 -647
rect 2162 -681 2196 -647
rect 2234 -681 2264 -647
rect 2306 -681 2332 -647
rect 2366 -681 2391 -647
rect 2757 -681 2782 -647
rect 2816 -681 2842 -647
rect 2884 -681 2914 -647
rect 2952 -681 2986 -647
rect 3020 -681 3054 -647
rect 3092 -681 3122 -647
rect 3164 -681 3190 -647
rect 3224 -681 3249 -647
rect 3615 -681 3640 -647
rect 3674 -681 3700 -647
rect 3742 -681 3772 -647
rect 3810 -681 3844 -647
rect 3878 -681 3912 -647
rect 3950 -681 3980 -647
rect 4022 -681 4048 -647
rect 4082 -681 4107 -647
rect 4473 -681 4498 -647
rect 4532 -681 4558 -647
rect 4600 -681 4630 -647
rect 4668 -681 4702 -647
rect 4736 -681 4770 -647
rect 4808 -681 4838 -647
rect 4880 -681 4906 -647
rect 4940 -681 4965 -647
rect 5331 -681 5356 -647
rect 5390 -681 5416 -647
rect 5458 -681 5488 -647
rect 5526 -681 5560 -647
rect 5594 -681 5628 -647
rect 5666 -681 5696 -647
rect 5738 -681 5764 -647
rect 5798 -681 5823 -647
<< viali >>
rect -5738 647 -5730 681
rect -5730 647 -5704 681
rect -5666 647 -5662 681
rect -5662 647 -5632 681
rect -5594 647 -5560 681
rect -5522 647 -5492 681
rect -5492 647 -5488 681
rect -5450 647 -5424 681
rect -5424 647 -5416 681
rect -4880 647 -4872 681
rect -4872 647 -4846 681
rect -4808 647 -4804 681
rect -4804 647 -4774 681
rect -4736 647 -4702 681
rect -4664 647 -4634 681
rect -4634 647 -4630 681
rect -4592 647 -4566 681
rect -4566 647 -4558 681
rect -4022 647 -4014 681
rect -4014 647 -3988 681
rect -3950 647 -3946 681
rect -3946 647 -3916 681
rect -3878 647 -3844 681
rect -3806 647 -3776 681
rect -3776 647 -3772 681
rect -3734 647 -3708 681
rect -3708 647 -3700 681
rect -3164 647 -3156 681
rect -3156 647 -3130 681
rect -3092 647 -3088 681
rect -3088 647 -3058 681
rect -3020 647 -2986 681
rect -2948 647 -2918 681
rect -2918 647 -2914 681
rect -2876 647 -2850 681
rect -2850 647 -2842 681
rect -2306 647 -2298 681
rect -2298 647 -2272 681
rect -2234 647 -2230 681
rect -2230 647 -2200 681
rect -2162 647 -2128 681
rect -2090 647 -2060 681
rect -2060 647 -2056 681
rect -2018 647 -1992 681
rect -1992 647 -1984 681
rect -1448 647 -1440 681
rect -1440 647 -1414 681
rect -1376 647 -1372 681
rect -1372 647 -1342 681
rect -1304 647 -1270 681
rect -1232 647 -1202 681
rect -1202 647 -1198 681
rect -1160 647 -1134 681
rect -1134 647 -1126 681
rect -590 647 -582 681
rect -582 647 -556 681
rect -518 647 -514 681
rect -514 647 -484 681
rect -446 647 -412 681
rect -374 647 -344 681
rect -344 647 -340 681
rect -302 647 -276 681
rect -276 647 -268 681
rect 268 647 276 681
rect 276 647 302 681
rect 340 647 344 681
rect 344 647 374 681
rect 412 647 446 681
rect 484 647 514 681
rect 514 647 518 681
rect 556 647 582 681
rect 582 647 590 681
rect 1126 647 1134 681
rect 1134 647 1160 681
rect 1198 647 1202 681
rect 1202 647 1232 681
rect 1270 647 1304 681
rect 1342 647 1372 681
rect 1372 647 1376 681
rect 1414 647 1440 681
rect 1440 647 1448 681
rect 1984 647 1992 681
rect 1992 647 2018 681
rect 2056 647 2060 681
rect 2060 647 2090 681
rect 2128 647 2162 681
rect 2200 647 2230 681
rect 2230 647 2234 681
rect 2272 647 2298 681
rect 2298 647 2306 681
rect 2842 647 2850 681
rect 2850 647 2876 681
rect 2914 647 2918 681
rect 2918 647 2948 681
rect 2986 647 3020 681
rect 3058 647 3088 681
rect 3088 647 3092 681
rect 3130 647 3156 681
rect 3156 647 3164 681
rect 3700 647 3708 681
rect 3708 647 3734 681
rect 3772 647 3776 681
rect 3776 647 3806 681
rect 3844 647 3878 681
rect 3916 647 3946 681
rect 3946 647 3950 681
rect 3988 647 4014 681
rect 4014 647 4022 681
rect 4558 647 4566 681
rect 4566 647 4592 681
rect 4630 647 4634 681
rect 4634 647 4664 681
rect 4702 647 4736 681
rect 4774 647 4804 681
rect 4804 647 4808 681
rect 4846 647 4872 681
rect 4872 647 4880 681
rect 5416 647 5424 681
rect 5424 647 5450 681
rect 5488 647 5492 681
rect 5492 647 5522 681
rect 5560 647 5594 681
rect 5632 647 5662 681
rect 5662 647 5666 681
rect 5704 647 5730 681
rect 5730 647 5738 681
rect -6023 527 -5989 557
rect -6023 523 -5989 527
rect -6023 459 -5989 485
rect -6023 451 -5989 459
rect -6023 391 -5989 413
rect -6023 379 -5989 391
rect -6023 323 -5989 341
rect -6023 307 -5989 323
rect -6023 255 -5989 269
rect -6023 235 -5989 255
rect -6023 187 -5989 197
rect -6023 163 -5989 187
rect -6023 119 -5989 125
rect -6023 91 -5989 119
rect -6023 51 -5989 53
rect -6023 19 -5989 51
rect -6023 -51 -5989 -19
rect -6023 -53 -5989 -51
rect -6023 -119 -5989 -91
rect -6023 -125 -5989 -119
rect -6023 -187 -5989 -163
rect -6023 -197 -5989 -187
rect -6023 -255 -5989 -235
rect -6023 -269 -5989 -255
rect -6023 -323 -5989 -307
rect -6023 -341 -5989 -323
rect -6023 -391 -5989 -379
rect -6023 -413 -5989 -391
rect -6023 -459 -5989 -451
rect -6023 -485 -5989 -459
rect -6023 -527 -5989 -523
rect -6023 -557 -5989 -527
rect -5165 527 -5131 557
rect -5165 523 -5131 527
rect -5165 459 -5131 485
rect -5165 451 -5131 459
rect -5165 391 -5131 413
rect -5165 379 -5131 391
rect -5165 323 -5131 341
rect -5165 307 -5131 323
rect -5165 255 -5131 269
rect -5165 235 -5131 255
rect -5165 187 -5131 197
rect -5165 163 -5131 187
rect -5165 119 -5131 125
rect -5165 91 -5131 119
rect -5165 51 -5131 53
rect -5165 19 -5131 51
rect -5165 -51 -5131 -19
rect -5165 -53 -5131 -51
rect -5165 -119 -5131 -91
rect -5165 -125 -5131 -119
rect -5165 -187 -5131 -163
rect -5165 -197 -5131 -187
rect -5165 -255 -5131 -235
rect -5165 -269 -5131 -255
rect -5165 -323 -5131 -307
rect -5165 -341 -5131 -323
rect -5165 -391 -5131 -379
rect -5165 -413 -5131 -391
rect -5165 -459 -5131 -451
rect -5165 -485 -5131 -459
rect -5165 -527 -5131 -523
rect -5165 -557 -5131 -527
rect -4307 527 -4273 557
rect -4307 523 -4273 527
rect -4307 459 -4273 485
rect -4307 451 -4273 459
rect -4307 391 -4273 413
rect -4307 379 -4273 391
rect -4307 323 -4273 341
rect -4307 307 -4273 323
rect -4307 255 -4273 269
rect -4307 235 -4273 255
rect -4307 187 -4273 197
rect -4307 163 -4273 187
rect -4307 119 -4273 125
rect -4307 91 -4273 119
rect -4307 51 -4273 53
rect -4307 19 -4273 51
rect -4307 -51 -4273 -19
rect -4307 -53 -4273 -51
rect -4307 -119 -4273 -91
rect -4307 -125 -4273 -119
rect -4307 -187 -4273 -163
rect -4307 -197 -4273 -187
rect -4307 -255 -4273 -235
rect -4307 -269 -4273 -255
rect -4307 -323 -4273 -307
rect -4307 -341 -4273 -323
rect -4307 -391 -4273 -379
rect -4307 -413 -4273 -391
rect -4307 -459 -4273 -451
rect -4307 -485 -4273 -459
rect -4307 -527 -4273 -523
rect -4307 -557 -4273 -527
rect -3449 527 -3415 557
rect -3449 523 -3415 527
rect -3449 459 -3415 485
rect -3449 451 -3415 459
rect -3449 391 -3415 413
rect -3449 379 -3415 391
rect -3449 323 -3415 341
rect -3449 307 -3415 323
rect -3449 255 -3415 269
rect -3449 235 -3415 255
rect -3449 187 -3415 197
rect -3449 163 -3415 187
rect -3449 119 -3415 125
rect -3449 91 -3415 119
rect -3449 51 -3415 53
rect -3449 19 -3415 51
rect -3449 -51 -3415 -19
rect -3449 -53 -3415 -51
rect -3449 -119 -3415 -91
rect -3449 -125 -3415 -119
rect -3449 -187 -3415 -163
rect -3449 -197 -3415 -187
rect -3449 -255 -3415 -235
rect -3449 -269 -3415 -255
rect -3449 -323 -3415 -307
rect -3449 -341 -3415 -323
rect -3449 -391 -3415 -379
rect -3449 -413 -3415 -391
rect -3449 -459 -3415 -451
rect -3449 -485 -3415 -459
rect -3449 -527 -3415 -523
rect -3449 -557 -3415 -527
rect -2591 527 -2557 557
rect -2591 523 -2557 527
rect -2591 459 -2557 485
rect -2591 451 -2557 459
rect -2591 391 -2557 413
rect -2591 379 -2557 391
rect -2591 323 -2557 341
rect -2591 307 -2557 323
rect -2591 255 -2557 269
rect -2591 235 -2557 255
rect -2591 187 -2557 197
rect -2591 163 -2557 187
rect -2591 119 -2557 125
rect -2591 91 -2557 119
rect -2591 51 -2557 53
rect -2591 19 -2557 51
rect -2591 -51 -2557 -19
rect -2591 -53 -2557 -51
rect -2591 -119 -2557 -91
rect -2591 -125 -2557 -119
rect -2591 -187 -2557 -163
rect -2591 -197 -2557 -187
rect -2591 -255 -2557 -235
rect -2591 -269 -2557 -255
rect -2591 -323 -2557 -307
rect -2591 -341 -2557 -323
rect -2591 -391 -2557 -379
rect -2591 -413 -2557 -391
rect -2591 -459 -2557 -451
rect -2591 -485 -2557 -459
rect -2591 -527 -2557 -523
rect -2591 -557 -2557 -527
rect -1733 527 -1699 557
rect -1733 523 -1699 527
rect -1733 459 -1699 485
rect -1733 451 -1699 459
rect -1733 391 -1699 413
rect -1733 379 -1699 391
rect -1733 323 -1699 341
rect -1733 307 -1699 323
rect -1733 255 -1699 269
rect -1733 235 -1699 255
rect -1733 187 -1699 197
rect -1733 163 -1699 187
rect -1733 119 -1699 125
rect -1733 91 -1699 119
rect -1733 51 -1699 53
rect -1733 19 -1699 51
rect -1733 -51 -1699 -19
rect -1733 -53 -1699 -51
rect -1733 -119 -1699 -91
rect -1733 -125 -1699 -119
rect -1733 -187 -1699 -163
rect -1733 -197 -1699 -187
rect -1733 -255 -1699 -235
rect -1733 -269 -1699 -255
rect -1733 -323 -1699 -307
rect -1733 -341 -1699 -323
rect -1733 -391 -1699 -379
rect -1733 -413 -1699 -391
rect -1733 -459 -1699 -451
rect -1733 -485 -1699 -459
rect -1733 -527 -1699 -523
rect -1733 -557 -1699 -527
rect -875 527 -841 557
rect -875 523 -841 527
rect -875 459 -841 485
rect -875 451 -841 459
rect -875 391 -841 413
rect -875 379 -841 391
rect -875 323 -841 341
rect -875 307 -841 323
rect -875 255 -841 269
rect -875 235 -841 255
rect -875 187 -841 197
rect -875 163 -841 187
rect -875 119 -841 125
rect -875 91 -841 119
rect -875 51 -841 53
rect -875 19 -841 51
rect -875 -51 -841 -19
rect -875 -53 -841 -51
rect -875 -119 -841 -91
rect -875 -125 -841 -119
rect -875 -187 -841 -163
rect -875 -197 -841 -187
rect -875 -255 -841 -235
rect -875 -269 -841 -255
rect -875 -323 -841 -307
rect -875 -341 -841 -323
rect -875 -391 -841 -379
rect -875 -413 -841 -391
rect -875 -459 -841 -451
rect -875 -485 -841 -459
rect -875 -527 -841 -523
rect -875 -557 -841 -527
rect -17 527 17 557
rect -17 523 17 527
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect -17 -527 17 -523
rect -17 -557 17 -527
rect 841 527 875 557
rect 841 523 875 527
rect 841 459 875 485
rect 841 451 875 459
rect 841 391 875 413
rect 841 379 875 391
rect 841 323 875 341
rect 841 307 875 323
rect 841 255 875 269
rect 841 235 875 255
rect 841 187 875 197
rect 841 163 875 187
rect 841 119 875 125
rect 841 91 875 119
rect 841 51 875 53
rect 841 19 875 51
rect 841 -51 875 -19
rect 841 -53 875 -51
rect 841 -119 875 -91
rect 841 -125 875 -119
rect 841 -187 875 -163
rect 841 -197 875 -187
rect 841 -255 875 -235
rect 841 -269 875 -255
rect 841 -323 875 -307
rect 841 -341 875 -323
rect 841 -391 875 -379
rect 841 -413 875 -391
rect 841 -459 875 -451
rect 841 -485 875 -459
rect 841 -527 875 -523
rect 841 -557 875 -527
rect 1699 527 1733 557
rect 1699 523 1733 527
rect 1699 459 1733 485
rect 1699 451 1733 459
rect 1699 391 1733 413
rect 1699 379 1733 391
rect 1699 323 1733 341
rect 1699 307 1733 323
rect 1699 255 1733 269
rect 1699 235 1733 255
rect 1699 187 1733 197
rect 1699 163 1733 187
rect 1699 119 1733 125
rect 1699 91 1733 119
rect 1699 51 1733 53
rect 1699 19 1733 51
rect 1699 -51 1733 -19
rect 1699 -53 1733 -51
rect 1699 -119 1733 -91
rect 1699 -125 1733 -119
rect 1699 -187 1733 -163
rect 1699 -197 1733 -187
rect 1699 -255 1733 -235
rect 1699 -269 1733 -255
rect 1699 -323 1733 -307
rect 1699 -341 1733 -323
rect 1699 -391 1733 -379
rect 1699 -413 1733 -391
rect 1699 -459 1733 -451
rect 1699 -485 1733 -459
rect 1699 -527 1733 -523
rect 1699 -557 1733 -527
rect 2557 527 2591 557
rect 2557 523 2591 527
rect 2557 459 2591 485
rect 2557 451 2591 459
rect 2557 391 2591 413
rect 2557 379 2591 391
rect 2557 323 2591 341
rect 2557 307 2591 323
rect 2557 255 2591 269
rect 2557 235 2591 255
rect 2557 187 2591 197
rect 2557 163 2591 187
rect 2557 119 2591 125
rect 2557 91 2591 119
rect 2557 51 2591 53
rect 2557 19 2591 51
rect 2557 -51 2591 -19
rect 2557 -53 2591 -51
rect 2557 -119 2591 -91
rect 2557 -125 2591 -119
rect 2557 -187 2591 -163
rect 2557 -197 2591 -187
rect 2557 -255 2591 -235
rect 2557 -269 2591 -255
rect 2557 -323 2591 -307
rect 2557 -341 2591 -323
rect 2557 -391 2591 -379
rect 2557 -413 2591 -391
rect 2557 -459 2591 -451
rect 2557 -485 2591 -459
rect 2557 -527 2591 -523
rect 2557 -557 2591 -527
rect 3415 527 3449 557
rect 3415 523 3449 527
rect 3415 459 3449 485
rect 3415 451 3449 459
rect 3415 391 3449 413
rect 3415 379 3449 391
rect 3415 323 3449 341
rect 3415 307 3449 323
rect 3415 255 3449 269
rect 3415 235 3449 255
rect 3415 187 3449 197
rect 3415 163 3449 187
rect 3415 119 3449 125
rect 3415 91 3449 119
rect 3415 51 3449 53
rect 3415 19 3449 51
rect 3415 -51 3449 -19
rect 3415 -53 3449 -51
rect 3415 -119 3449 -91
rect 3415 -125 3449 -119
rect 3415 -187 3449 -163
rect 3415 -197 3449 -187
rect 3415 -255 3449 -235
rect 3415 -269 3449 -255
rect 3415 -323 3449 -307
rect 3415 -341 3449 -323
rect 3415 -391 3449 -379
rect 3415 -413 3449 -391
rect 3415 -459 3449 -451
rect 3415 -485 3449 -459
rect 3415 -527 3449 -523
rect 3415 -557 3449 -527
rect 4273 527 4307 557
rect 4273 523 4307 527
rect 4273 459 4307 485
rect 4273 451 4307 459
rect 4273 391 4307 413
rect 4273 379 4307 391
rect 4273 323 4307 341
rect 4273 307 4307 323
rect 4273 255 4307 269
rect 4273 235 4307 255
rect 4273 187 4307 197
rect 4273 163 4307 187
rect 4273 119 4307 125
rect 4273 91 4307 119
rect 4273 51 4307 53
rect 4273 19 4307 51
rect 4273 -51 4307 -19
rect 4273 -53 4307 -51
rect 4273 -119 4307 -91
rect 4273 -125 4307 -119
rect 4273 -187 4307 -163
rect 4273 -197 4307 -187
rect 4273 -255 4307 -235
rect 4273 -269 4307 -255
rect 4273 -323 4307 -307
rect 4273 -341 4307 -323
rect 4273 -391 4307 -379
rect 4273 -413 4307 -391
rect 4273 -459 4307 -451
rect 4273 -485 4307 -459
rect 4273 -527 4307 -523
rect 4273 -557 4307 -527
rect 5131 527 5165 557
rect 5131 523 5165 527
rect 5131 459 5165 485
rect 5131 451 5165 459
rect 5131 391 5165 413
rect 5131 379 5165 391
rect 5131 323 5165 341
rect 5131 307 5165 323
rect 5131 255 5165 269
rect 5131 235 5165 255
rect 5131 187 5165 197
rect 5131 163 5165 187
rect 5131 119 5165 125
rect 5131 91 5165 119
rect 5131 51 5165 53
rect 5131 19 5165 51
rect 5131 -51 5165 -19
rect 5131 -53 5165 -51
rect 5131 -119 5165 -91
rect 5131 -125 5165 -119
rect 5131 -187 5165 -163
rect 5131 -197 5165 -187
rect 5131 -255 5165 -235
rect 5131 -269 5165 -255
rect 5131 -323 5165 -307
rect 5131 -341 5165 -323
rect 5131 -391 5165 -379
rect 5131 -413 5165 -391
rect 5131 -459 5165 -451
rect 5131 -485 5165 -459
rect 5131 -527 5165 -523
rect 5131 -557 5165 -527
rect 5989 527 6023 557
rect 5989 523 6023 527
rect 5989 459 6023 485
rect 5989 451 6023 459
rect 5989 391 6023 413
rect 5989 379 6023 391
rect 5989 323 6023 341
rect 5989 307 6023 323
rect 5989 255 6023 269
rect 5989 235 6023 255
rect 5989 187 6023 197
rect 5989 163 6023 187
rect 5989 119 6023 125
rect 5989 91 6023 119
rect 5989 51 6023 53
rect 5989 19 6023 51
rect 5989 -51 6023 -19
rect 5989 -53 6023 -51
rect 5989 -119 6023 -91
rect 5989 -125 6023 -119
rect 5989 -187 6023 -163
rect 5989 -197 6023 -187
rect 5989 -255 6023 -235
rect 5989 -269 6023 -255
rect 5989 -323 6023 -307
rect 5989 -341 6023 -323
rect 5989 -391 6023 -379
rect 5989 -413 6023 -391
rect 5989 -459 6023 -451
rect 5989 -485 6023 -459
rect 5989 -527 6023 -523
rect 5989 -557 6023 -527
rect -5738 -681 -5730 -647
rect -5730 -681 -5704 -647
rect -5666 -681 -5662 -647
rect -5662 -681 -5632 -647
rect -5594 -681 -5560 -647
rect -5522 -681 -5492 -647
rect -5492 -681 -5488 -647
rect -5450 -681 -5424 -647
rect -5424 -681 -5416 -647
rect -4880 -681 -4872 -647
rect -4872 -681 -4846 -647
rect -4808 -681 -4804 -647
rect -4804 -681 -4774 -647
rect -4736 -681 -4702 -647
rect -4664 -681 -4634 -647
rect -4634 -681 -4630 -647
rect -4592 -681 -4566 -647
rect -4566 -681 -4558 -647
rect -4022 -681 -4014 -647
rect -4014 -681 -3988 -647
rect -3950 -681 -3946 -647
rect -3946 -681 -3916 -647
rect -3878 -681 -3844 -647
rect -3806 -681 -3776 -647
rect -3776 -681 -3772 -647
rect -3734 -681 -3708 -647
rect -3708 -681 -3700 -647
rect -3164 -681 -3156 -647
rect -3156 -681 -3130 -647
rect -3092 -681 -3088 -647
rect -3088 -681 -3058 -647
rect -3020 -681 -2986 -647
rect -2948 -681 -2918 -647
rect -2918 -681 -2914 -647
rect -2876 -681 -2850 -647
rect -2850 -681 -2842 -647
rect -2306 -681 -2298 -647
rect -2298 -681 -2272 -647
rect -2234 -681 -2230 -647
rect -2230 -681 -2200 -647
rect -2162 -681 -2128 -647
rect -2090 -681 -2060 -647
rect -2060 -681 -2056 -647
rect -2018 -681 -1992 -647
rect -1992 -681 -1984 -647
rect -1448 -681 -1440 -647
rect -1440 -681 -1414 -647
rect -1376 -681 -1372 -647
rect -1372 -681 -1342 -647
rect -1304 -681 -1270 -647
rect -1232 -681 -1202 -647
rect -1202 -681 -1198 -647
rect -1160 -681 -1134 -647
rect -1134 -681 -1126 -647
rect -590 -681 -582 -647
rect -582 -681 -556 -647
rect -518 -681 -514 -647
rect -514 -681 -484 -647
rect -446 -681 -412 -647
rect -374 -681 -344 -647
rect -344 -681 -340 -647
rect -302 -681 -276 -647
rect -276 -681 -268 -647
rect 268 -681 276 -647
rect 276 -681 302 -647
rect 340 -681 344 -647
rect 344 -681 374 -647
rect 412 -681 446 -647
rect 484 -681 514 -647
rect 514 -681 518 -647
rect 556 -681 582 -647
rect 582 -681 590 -647
rect 1126 -681 1134 -647
rect 1134 -681 1160 -647
rect 1198 -681 1202 -647
rect 1202 -681 1232 -647
rect 1270 -681 1304 -647
rect 1342 -681 1372 -647
rect 1372 -681 1376 -647
rect 1414 -681 1440 -647
rect 1440 -681 1448 -647
rect 1984 -681 1992 -647
rect 1992 -681 2018 -647
rect 2056 -681 2060 -647
rect 2060 -681 2090 -647
rect 2128 -681 2162 -647
rect 2200 -681 2230 -647
rect 2230 -681 2234 -647
rect 2272 -681 2298 -647
rect 2298 -681 2306 -647
rect 2842 -681 2850 -647
rect 2850 -681 2876 -647
rect 2914 -681 2918 -647
rect 2918 -681 2948 -647
rect 2986 -681 3020 -647
rect 3058 -681 3088 -647
rect 3088 -681 3092 -647
rect 3130 -681 3156 -647
rect 3156 -681 3164 -647
rect 3700 -681 3708 -647
rect 3708 -681 3734 -647
rect 3772 -681 3776 -647
rect 3776 -681 3806 -647
rect 3844 -681 3878 -647
rect 3916 -681 3946 -647
rect 3946 -681 3950 -647
rect 3988 -681 4014 -647
rect 4014 -681 4022 -647
rect 4558 -681 4566 -647
rect 4566 -681 4592 -647
rect 4630 -681 4634 -647
rect 4634 -681 4664 -647
rect 4702 -681 4736 -647
rect 4774 -681 4804 -647
rect 4804 -681 4808 -647
rect 4846 -681 4872 -647
rect 4872 -681 4880 -647
rect 5416 -681 5424 -647
rect 5424 -681 5450 -647
rect 5488 -681 5492 -647
rect 5492 -681 5522 -647
rect 5560 -681 5594 -647
rect 5632 -681 5662 -647
rect 5662 -681 5666 -647
rect 5704 -681 5730 -647
rect 5730 -681 5738 -647
<< metal1 >>
rect -5781 681 -5373 687
rect -5781 647 -5738 681
rect -5704 647 -5666 681
rect -5632 647 -5594 681
rect -5560 647 -5522 681
rect -5488 647 -5450 681
rect -5416 647 -5373 681
rect -5781 641 -5373 647
rect -4923 681 -4515 687
rect -4923 647 -4880 681
rect -4846 647 -4808 681
rect -4774 647 -4736 681
rect -4702 647 -4664 681
rect -4630 647 -4592 681
rect -4558 647 -4515 681
rect -4923 641 -4515 647
rect -4065 681 -3657 687
rect -4065 647 -4022 681
rect -3988 647 -3950 681
rect -3916 647 -3878 681
rect -3844 647 -3806 681
rect -3772 647 -3734 681
rect -3700 647 -3657 681
rect -4065 641 -3657 647
rect -3207 681 -2799 687
rect -3207 647 -3164 681
rect -3130 647 -3092 681
rect -3058 647 -3020 681
rect -2986 647 -2948 681
rect -2914 647 -2876 681
rect -2842 647 -2799 681
rect -3207 641 -2799 647
rect -2349 681 -1941 687
rect -2349 647 -2306 681
rect -2272 647 -2234 681
rect -2200 647 -2162 681
rect -2128 647 -2090 681
rect -2056 647 -2018 681
rect -1984 647 -1941 681
rect -2349 641 -1941 647
rect -1491 681 -1083 687
rect -1491 647 -1448 681
rect -1414 647 -1376 681
rect -1342 647 -1304 681
rect -1270 647 -1232 681
rect -1198 647 -1160 681
rect -1126 647 -1083 681
rect -1491 641 -1083 647
rect -633 681 -225 687
rect -633 647 -590 681
rect -556 647 -518 681
rect -484 647 -446 681
rect -412 647 -374 681
rect -340 647 -302 681
rect -268 647 -225 681
rect -633 641 -225 647
rect 225 681 633 687
rect 225 647 268 681
rect 302 647 340 681
rect 374 647 412 681
rect 446 647 484 681
rect 518 647 556 681
rect 590 647 633 681
rect 225 641 633 647
rect 1083 681 1491 687
rect 1083 647 1126 681
rect 1160 647 1198 681
rect 1232 647 1270 681
rect 1304 647 1342 681
rect 1376 647 1414 681
rect 1448 647 1491 681
rect 1083 641 1491 647
rect 1941 681 2349 687
rect 1941 647 1984 681
rect 2018 647 2056 681
rect 2090 647 2128 681
rect 2162 647 2200 681
rect 2234 647 2272 681
rect 2306 647 2349 681
rect 1941 641 2349 647
rect 2799 681 3207 687
rect 2799 647 2842 681
rect 2876 647 2914 681
rect 2948 647 2986 681
rect 3020 647 3058 681
rect 3092 647 3130 681
rect 3164 647 3207 681
rect 2799 641 3207 647
rect 3657 681 4065 687
rect 3657 647 3700 681
rect 3734 647 3772 681
rect 3806 647 3844 681
rect 3878 647 3916 681
rect 3950 647 3988 681
rect 4022 647 4065 681
rect 3657 641 4065 647
rect 4515 681 4923 687
rect 4515 647 4558 681
rect 4592 647 4630 681
rect 4664 647 4702 681
rect 4736 647 4774 681
rect 4808 647 4846 681
rect 4880 647 4923 681
rect 4515 641 4923 647
rect 5373 681 5781 687
rect 5373 647 5416 681
rect 5450 647 5488 681
rect 5522 647 5560 681
rect 5594 647 5632 681
rect 5666 647 5704 681
rect 5738 647 5781 681
rect 5373 641 5781 647
rect -6029 557 -5983 600
rect -6029 523 -6023 557
rect -5989 523 -5983 557
rect -6029 485 -5983 523
rect -6029 451 -6023 485
rect -5989 451 -5983 485
rect -6029 413 -5983 451
rect -6029 379 -6023 413
rect -5989 379 -5983 413
rect -6029 341 -5983 379
rect -6029 307 -6023 341
rect -5989 307 -5983 341
rect -6029 269 -5983 307
rect -6029 235 -6023 269
rect -5989 235 -5983 269
rect -6029 197 -5983 235
rect -6029 163 -6023 197
rect -5989 163 -5983 197
rect -6029 125 -5983 163
rect -6029 91 -6023 125
rect -5989 91 -5983 125
rect -6029 53 -5983 91
rect -6029 19 -6023 53
rect -5989 19 -5983 53
rect -6029 -19 -5983 19
rect -6029 -53 -6023 -19
rect -5989 -53 -5983 -19
rect -6029 -91 -5983 -53
rect -6029 -125 -6023 -91
rect -5989 -125 -5983 -91
rect -6029 -163 -5983 -125
rect -6029 -197 -6023 -163
rect -5989 -197 -5983 -163
rect -6029 -235 -5983 -197
rect -6029 -269 -6023 -235
rect -5989 -269 -5983 -235
rect -6029 -307 -5983 -269
rect -6029 -341 -6023 -307
rect -5989 -341 -5983 -307
rect -6029 -379 -5983 -341
rect -6029 -413 -6023 -379
rect -5989 -413 -5983 -379
rect -6029 -451 -5983 -413
rect -6029 -485 -6023 -451
rect -5989 -485 -5983 -451
rect -6029 -523 -5983 -485
rect -6029 -557 -6023 -523
rect -5989 -557 -5983 -523
rect -6029 -600 -5983 -557
rect -5171 557 -5125 600
rect -5171 523 -5165 557
rect -5131 523 -5125 557
rect -5171 485 -5125 523
rect -5171 451 -5165 485
rect -5131 451 -5125 485
rect -5171 413 -5125 451
rect -5171 379 -5165 413
rect -5131 379 -5125 413
rect -5171 341 -5125 379
rect -5171 307 -5165 341
rect -5131 307 -5125 341
rect -5171 269 -5125 307
rect -5171 235 -5165 269
rect -5131 235 -5125 269
rect -5171 197 -5125 235
rect -5171 163 -5165 197
rect -5131 163 -5125 197
rect -5171 125 -5125 163
rect -5171 91 -5165 125
rect -5131 91 -5125 125
rect -5171 53 -5125 91
rect -5171 19 -5165 53
rect -5131 19 -5125 53
rect -5171 -19 -5125 19
rect -5171 -53 -5165 -19
rect -5131 -53 -5125 -19
rect -5171 -91 -5125 -53
rect -5171 -125 -5165 -91
rect -5131 -125 -5125 -91
rect -5171 -163 -5125 -125
rect -5171 -197 -5165 -163
rect -5131 -197 -5125 -163
rect -5171 -235 -5125 -197
rect -5171 -269 -5165 -235
rect -5131 -269 -5125 -235
rect -5171 -307 -5125 -269
rect -5171 -341 -5165 -307
rect -5131 -341 -5125 -307
rect -5171 -379 -5125 -341
rect -5171 -413 -5165 -379
rect -5131 -413 -5125 -379
rect -5171 -451 -5125 -413
rect -5171 -485 -5165 -451
rect -5131 -485 -5125 -451
rect -5171 -523 -5125 -485
rect -5171 -557 -5165 -523
rect -5131 -557 -5125 -523
rect -5171 -600 -5125 -557
rect -4313 557 -4267 600
rect -4313 523 -4307 557
rect -4273 523 -4267 557
rect -4313 485 -4267 523
rect -4313 451 -4307 485
rect -4273 451 -4267 485
rect -4313 413 -4267 451
rect -4313 379 -4307 413
rect -4273 379 -4267 413
rect -4313 341 -4267 379
rect -4313 307 -4307 341
rect -4273 307 -4267 341
rect -4313 269 -4267 307
rect -4313 235 -4307 269
rect -4273 235 -4267 269
rect -4313 197 -4267 235
rect -4313 163 -4307 197
rect -4273 163 -4267 197
rect -4313 125 -4267 163
rect -4313 91 -4307 125
rect -4273 91 -4267 125
rect -4313 53 -4267 91
rect -4313 19 -4307 53
rect -4273 19 -4267 53
rect -4313 -19 -4267 19
rect -4313 -53 -4307 -19
rect -4273 -53 -4267 -19
rect -4313 -91 -4267 -53
rect -4313 -125 -4307 -91
rect -4273 -125 -4267 -91
rect -4313 -163 -4267 -125
rect -4313 -197 -4307 -163
rect -4273 -197 -4267 -163
rect -4313 -235 -4267 -197
rect -4313 -269 -4307 -235
rect -4273 -269 -4267 -235
rect -4313 -307 -4267 -269
rect -4313 -341 -4307 -307
rect -4273 -341 -4267 -307
rect -4313 -379 -4267 -341
rect -4313 -413 -4307 -379
rect -4273 -413 -4267 -379
rect -4313 -451 -4267 -413
rect -4313 -485 -4307 -451
rect -4273 -485 -4267 -451
rect -4313 -523 -4267 -485
rect -4313 -557 -4307 -523
rect -4273 -557 -4267 -523
rect -4313 -600 -4267 -557
rect -3455 557 -3409 600
rect -3455 523 -3449 557
rect -3415 523 -3409 557
rect -3455 485 -3409 523
rect -3455 451 -3449 485
rect -3415 451 -3409 485
rect -3455 413 -3409 451
rect -3455 379 -3449 413
rect -3415 379 -3409 413
rect -3455 341 -3409 379
rect -3455 307 -3449 341
rect -3415 307 -3409 341
rect -3455 269 -3409 307
rect -3455 235 -3449 269
rect -3415 235 -3409 269
rect -3455 197 -3409 235
rect -3455 163 -3449 197
rect -3415 163 -3409 197
rect -3455 125 -3409 163
rect -3455 91 -3449 125
rect -3415 91 -3409 125
rect -3455 53 -3409 91
rect -3455 19 -3449 53
rect -3415 19 -3409 53
rect -3455 -19 -3409 19
rect -3455 -53 -3449 -19
rect -3415 -53 -3409 -19
rect -3455 -91 -3409 -53
rect -3455 -125 -3449 -91
rect -3415 -125 -3409 -91
rect -3455 -163 -3409 -125
rect -3455 -197 -3449 -163
rect -3415 -197 -3409 -163
rect -3455 -235 -3409 -197
rect -3455 -269 -3449 -235
rect -3415 -269 -3409 -235
rect -3455 -307 -3409 -269
rect -3455 -341 -3449 -307
rect -3415 -341 -3409 -307
rect -3455 -379 -3409 -341
rect -3455 -413 -3449 -379
rect -3415 -413 -3409 -379
rect -3455 -451 -3409 -413
rect -3455 -485 -3449 -451
rect -3415 -485 -3409 -451
rect -3455 -523 -3409 -485
rect -3455 -557 -3449 -523
rect -3415 -557 -3409 -523
rect -3455 -600 -3409 -557
rect -2597 557 -2551 600
rect -2597 523 -2591 557
rect -2557 523 -2551 557
rect -2597 485 -2551 523
rect -2597 451 -2591 485
rect -2557 451 -2551 485
rect -2597 413 -2551 451
rect -2597 379 -2591 413
rect -2557 379 -2551 413
rect -2597 341 -2551 379
rect -2597 307 -2591 341
rect -2557 307 -2551 341
rect -2597 269 -2551 307
rect -2597 235 -2591 269
rect -2557 235 -2551 269
rect -2597 197 -2551 235
rect -2597 163 -2591 197
rect -2557 163 -2551 197
rect -2597 125 -2551 163
rect -2597 91 -2591 125
rect -2557 91 -2551 125
rect -2597 53 -2551 91
rect -2597 19 -2591 53
rect -2557 19 -2551 53
rect -2597 -19 -2551 19
rect -2597 -53 -2591 -19
rect -2557 -53 -2551 -19
rect -2597 -91 -2551 -53
rect -2597 -125 -2591 -91
rect -2557 -125 -2551 -91
rect -2597 -163 -2551 -125
rect -2597 -197 -2591 -163
rect -2557 -197 -2551 -163
rect -2597 -235 -2551 -197
rect -2597 -269 -2591 -235
rect -2557 -269 -2551 -235
rect -2597 -307 -2551 -269
rect -2597 -341 -2591 -307
rect -2557 -341 -2551 -307
rect -2597 -379 -2551 -341
rect -2597 -413 -2591 -379
rect -2557 -413 -2551 -379
rect -2597 -451 -2551 -413
rect -2597 -485 -2591 -451
rect -2557 -485 -2551 -451
rect -2597 -523 -2551 -485
rect -2597 -557 -2591 -523
rect -2557 -557 -2551 -523
rect -2597 -600 -2551 -557
rect -1739 557 -1693 600
rect -1739 523 -1733 557
rect -1699 523 -1693 557
rect -1739 485 -1693 523
rect -1739 451 -1733 485
rect -1699 451 -1693 485
rect -1739 413 -1693 451
rect -1739 379 -1733 413
rect -1699 379 -1693 413
rect -1739 341 -1693 379
rect -1739 307 -1733 341
rect -1699 307 -1693 341
rect -1739 269 -1693 307
rect -1739 235 -1733 269
rect -1699 235 -1693 269
rect -1739 197 -1693 235
rect -1739 163 -1733 197
rect -1699 163 -1693 197
rect -1739 125 -1693 163
rect -1739 91 -1733 125
rect -1699 91 -1693 125
rect -1739 53 -1693 91
rect -1739 19 -1733 53
rect -1699 19 -1693 53
rect -1739 -19 -1693 19
rect -1739 -53 -1733 -19
rect -1699 -53 -1693 -19
rect -1739 -91 -1693 -53
rect -1739 -125 -1733 -91
rect -1699 -125 -1693 -91
rect -1739 -163 -1693 -125
rect -1739 -197 -1733 -163
rect -1699 -197 -1693 -163
rect -1739 -235 -1693 -197
rect -1739 -269 -1733 -235
rect -1699 -269 -1693 -235
rect -1739 -307 -1693 -269
rect -1739 -341 -1733 -307
rect -1699 -341 -1693 -307
rect -1739 -379 -1693 -341
rect -1739 -413 -1733 -379
rect -1699 -413 -1693 -379
rect -1739 -451 -1693 -413
rect -1739 -485 -1733 -451
rect -1699 -485 -1693 -451
rect -1739 -523 -1693 -485
rect -1739 -557 -1733 -523
rect -1699 -557 -1693 -523
rect -1739 -600 -1693 -557
rect -881 557 -835 600
rect -881 523 -875 557
rect -841 523 -835 557
rect -881 485 -835 523
rect -881 451 -875 485
rect -841 451 -835 485
rect -881 413 -835 451
rect -881 379 -875 413
rect -841 379 -835 413
rect -881 341 -835 379
rect -881 307 -875 341
rect -841 307 -835 341
rect -881 269 -835 307
rect -881 235 -875 269
rect -841 235 -835 269
rect -881 197 -835 235
rect -881 163 -875 197
rect -841 163 -835 197
rect -881 125 -835 163
rect -881 91 -875 125
rect -841 91 -835 125
rect -881 53 -835 91
rect -881 19 -875 53
rect -841 19 -835 53
rect -881 -19 -835 19
rect -881 -53 -875 -19
rect -841 -53 -835 -19
rect -881 -91 -835 -53
rect -881 -125 -875 -91
rect -841 -125 -835 -91
rect -881 -163 -835 -125
rect -881 -197 -875 -163
rect -841 -197 -835 -163
rect -881 -235 -835 -197
rect -881 -269 -875 -235
rect -841 -269 -835 -235
rect -881 -307 -835 -269
rect -881 -341 -875 -307
rect -841 -341 -835 -307
rect -881 -379 -835 -341
rect -881 -413 -875 -379
rect -841 -413 -835 -379
rect -881 -451 -835 -413
rect -881 -485 -875 -451
rect -841 -485 -835 -451
rect -881 -523 -835 -485
rect -881 -557 -875 -523
rect -841 -557 -835 -523
rect -881 -600 -835 -557
rect -23 557 23 600
rect -23 523 -17 557
rect 17 523 23 557
rect -23 485 23 523
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -523 23 -485
rect -23 -557 -17 -523
rect 17 -557 23 -523
rect -23 -600 23 -557
rect 835 557 881 600
rect 835 523 841 557
rect 875 523 881 557
rect 835 485 881 523
rect 835 451 841 485
rect 875 451 881 485
rect 835 413 881 451
rect 835 379 841 413
rect 875 379 881 413
rect 835 341 881 379
rect 835 307 841 341
rect 875 307 881 341
rect 835 269 881 307
rect 835 235 841 269
rect 875 235 881 269
rect 835 197 881 235
rect 835 163 841 197
rect 875 163 881 197
rect 835 125 881 163
rect 835 91 841 125
rect 875 91 881 125
rect 835 53 881 91
rect 835 19 841 53
rect 875 19 881 53
rect 835 -19 881 19
rect 835 -53 841 -19
rect 875 -53 881 -19
rect 835 -91 881 -53
rect 835 -125 841 -91
rect 875 -125 881 -91
rect 835 -163 881 -125
rect 835 -197 841 -163
rect 875 -197 881 -163
rect 835 -235 881 -197
rect 835 -269 841 -235
rect 875 -269 881 -235
rect 835 -307 881 -269
rect 835 -341 841 -307
rect 875 -341 881 -307
rect 835 -379 881 -341
rect 835 -413 841 -379
rect 875 -413 881 -379
rect 835 -451 881 -413
rect 835 -485 841 -451
rect 875 -485 881 -451
rect 835 -523 881 -485
rect 835 -557 841 -523
rect 875 -557 881 -523
rect 835 -600 881 -557
rect 1693 557 1739 600
rect 1693 523 1699 557
rect 1733 523 1739 557
rect 1693 485 1739 523
rect 1693 451 1699 485
rect 1733 451 1739 485
rect 1693 413 1739 451
rect 1693 379 1699 413
rect 1733 379 1739 413
rect 1693 341 1739 379
rect 1693 307 1699 341
rect 1733 307 1739 341
rect 1693 269 1739 307
rect 1693 235 1699 269
rect 1733 235 1739 269
rect 1693 197 1739 235
rect 1693 163 1699 197
rect 1733 163 1739 197
rect 1693 125 1739 163
rect 1693 91 1699 125
rect 1733 91 1739 125
rect 1693 53 1739 91
rect 1693 19 1699 53
rect 1733 19 1739 53
rect 1693 -19 1739 19
rect 1693 -53 1699 -19
rect 1733 -53 1739 -19
rect 1693 -91 1739 -53
rect 1693 -125 1699 -91
rect 1733 -125 1739 -91
rect 1693 -163 1739 -125
rect 1693 -197 1699 -163
rect 1733 -197 1739 -163
rect 1693 -235 1739 -197
rect 1693 -269 1699 -235
rect 1733 -269 1739 -235
rect 1693 -307 1739 -269
rect 1693 -341 1699 -307
rect 1733 -341 1739 -307
rect 1693 -379 1739 -341
rect 1693 -413 1699 -379
rect 1733 -413 1739 -379
rect 1693 -451 1739 -413
rect 1693 -485 1699 -451
rect 1733 -485 1739 -451
rect 1693 -523 1739 -485
rect 1693 -557 1699 -523
rect 1733 -557 1739 -523
rect 1693 -600 1739 -557
rect 2551 557 2597 600
rect 2551 523 2557 557
rect 2591 523 2597 557
rect 2551 485 2597 523
rect 2551 451 2557 485
rect 2591 451 2597 485
rect 2551 413 2597 451
rect 2551 379 2557 413
rect 2591 379 2597 413
rect 2551 341 2597 379
rect 2551 307 2557 341
rect 2591 307 2597 341
rect 2551 269 2597 307
rect 2551 235 2557 269
rect 2591 235 2597 269
rect 2551 197 2597 235
rect 2551 163 2557 197
rect 2591 163 2597 197
rect 2551 125 2597 163
rect 2551 91 2557 125
rect 2591 91 2597 125
rect 2551 53 2597 91
rect 2551 19 2557 53
rect 2591 19 2597 53
rect 2551 -19 2597 19
rect 2551 -53 2557 -19
rect 2591 -53 2597 -19
rect 2551 -91 2597 -53
rect 2551 -125 2557 -91
rect 2591 -125 2597 -91
rect 2551 -163 2597 -125
rect 2551 -197 2557 -163
rect 2591 -197 2597 -163
rect 2551 -235 2597 -197
rect 2551 -269 2557 -235
rect 2591 -269 2597 -235
rect 2551 -307 2597 -269
rect 2551 -341 2557 -307
rect 2591 -341 2597 -307
rect 2551 -379 2597 -341
rect 2551 -413 2557 -379
rect 2591 -413 2597 -379
rect 2551 -451 2597 -413
rect 2551 -485 2557 -451
rect 2591 -485 2597 -451
rect 2551 -523 2597 -485
rect 2551 -557 2557 -523
rect 2591 -557 2597 -523
rect 2551 -600 2597 -557
rect 3409 557 3455 600
rect 3409 523 3415 557
rect 3449 523 3455 557
rect 3409 485 3455 523
rect 3409 451 3415 485
rect 3449 451 3455 485
rect 3409 413 3455 451
rect 3409 379 3415 413
rect 3449 379 3455 413
rect 3409 341 3455 379
rect 3409 307 3415 341
rect 3449 307 3455 341
rect 3409 269 3455 307
rect 3409 235 3415 269
rect 3449 235 3455 269
rect 3409 197 3455 235
rect 3409 163 3415 197
rect 3449 163 3455 197
rect 3409 125 3455 163
rect 3409 91 3415 125
rect 3449 91 3455 125
rect 3409 53 3455 91
rect 3409 19 3415 53
rect 3449 19 3455 53
rect 3409 -19 3455 19
rect 3409 -53 3415 -19
rect 3449 -53 3455 -19
rect 3409 -91 3455 -53
rect 3409 -125 3415 -91
rect 3449 -125 3455 -91
rect 3409 -163 3455 -125
rect 3409 -197 3415 -163
rect 3449 -197 3455 -163
rect 3409 -235 3455 -197
rect 3409 -269 3415 -235
rect 3449 -269 3455 -235
rect 3409 -307 3455 -269
rect 3409 -341 3415 -307
rect 3449 -341 3455 -307
rect 3409 -379 3455 -341
rect 3409 -413 3415 -379
rect 3449 -413 3455 -379
rect 3409 -451 3455 -413
rect 3409 -485 3415 -451
rect 3449 -485 3455 -451
rect 3409 -523 3455 -485
rect 3409 -557 3415 -523
rect 3449 -557 3455 -523
rect 3409 -600 3455 -557
rect 4267 557 4313 600
rect 4267 523 4273 557
rect 4307 523 4313 557
rect 4267 485 4313 523
rect 4267 451 4273 485
rect 4307 451 4313 485
rect 4267 413 4313 451
rect 4267 379 4273 413
rect 4307 379 4313 413
rect 4267 341 4313 379
rect 4267 307 4273 341
rect 4307 307 4313 341
rect 4267 269 4313 307
rect 4267 235 4273 269
rect 4307 235 4313 269
rect 4267 197 4313 235
rect 4267 163 4273 197
rect 4307 163 4313 197
rect 4267 125 4313 163
rect 4267 91 4273 125
rect 4307 91 4313 125
rect 4267 53 4313 91
rect 4267 19 4273 53
rect 4307 19 4313 53
rect 4267 -19 4313 19
rect 4267 -53 4273 -19
rect 4307 -53 4313 -19
rect 4267 -91 4313 -53
rect 4267 -125 4273 -91
rect 4307 -125 4313 -91
rect 4267 -163 4313 -125
rect 4267 -197 4273 -163
rect 4307 -197 4313 -163
rect 4267 -235 4313 -197
rect 4267 -269 4273 -235
rect 4307 -269 4313 -235
rect 4267 -307 4313 -269
rect 4267 -341 4273 -307
rect 4307 -341 4313 -307
rect 4267 -379 4313 -341
rect 4267 -413 4273 -379
rect 4307 -413 4313 -379
rect 4267 -451 4313 -413
rect 4267 -485 4273 -451
rect 4307 -485 4313 -451
rect 4267 -523 4313 -485
rect 4267 -557 4273 -523
rect 4307 -557 4313 -523
rect 4267 -600 4313 -557
rect 5125 557 5171 600
rect 5125 523 5131 557
rect 5165 523 5171 557
rect 5125 485 5171 523
rect 5125 451 5131 485
rect 5165 451 5171 485
rect 5125 413 5171 451
rect 5125 379 5131 413
rect 5165 379 5171 413
rect 5125 341 5171 379
rect 5125 307 5131 341
rect 5165 307 5171 341
rect 5125 269 5171 307
rect 5125 235 5131 269
rect 5165 235 5171 269
rect 5125 197 5171 235
rect 5125 163 5131 197
rect 5165 163 5171 197
rect 5125 125 5171 163
rect 5125 91 5131 125
rect 5165 91 5171 125
rect 5125 53 5171 91
rect 5125 19 5131 53
rect 5165 19 5171 53
rect 5125 -19 5171 19
rect 5125 -53 5131 -19
rect 5165 -53 5171 -19
rect 5125 -91 5171 -53
rect 5125 -125 5131 -91
rect 5165 -125 5171 -91
rect 5125 -163 5171 -125
rect 5125 -197 5131 -163
rect 5165 -197 5171 -163
rect 5125 -235 5171 -197
rect 5125 -269 5131 -235
rect 5165 -269 5171 -235
rect 5125 -307 5171 -269
rect 5125 -341 5131 -307
rect 5165 -341 5171 -307
rect 5125 -379 5171 -341
rect 5125 -413 5131 -379
rect 5165 -413 5171 -379
rect 5125 -451 5171 -413
rect 5125 -485 5131 -451
rect 5165 -485 5171 -451
rect 5125 -523 5171 -485
rect 5125 -557 5131 -523
rect 5165 -557 5171 -523
rect 5125 -600 5171 -557
rect 5983 557 6029 600
rect 5983 523 5989 557
rect 6023 523 6029 557
rect 5983 485 6029 523
rect 5983 451 5989 485
rect 6023 451 6029 485
rect 5983 413 6029 451
rect 5983 379 5989 413
rect 6023 379 6029 413
rect 5983 341 6029 379
rect 5983 307 5989 341
rect 6023 307 6029 341
rect 5983 269 6029 307
rect 5983 235 5989 269
rect 6023 235 6029 269
rect 5983 197 6029 235
rect 5983 163 5989 197
rect 6023 163 6029 197
rect 5983 125 6029 163
rect 5983 91 5989 125
rect 6023 91 6029 125
rect 5983 53 6029 91
rect 5983 19 5989 53
rect 6023 19 6029 53
rect 5983 -19 6029 19
rect 5983 -53 5989 -19
rect 6023 -53 6029 -19
rect 5983 -91 6029 -53
rect 5983 -125 5989 -91
rect 6023 -125 6029 -91
rect 5983 -163 6029 -125
rect 5983 -197 5989 -163
rect 6023 -197 6029 -163
rect 5983 -235 6029 -197
rect 5983 -269 5989 -235
rect 6023 -269 6029 -235
rect 5983 -307 6029 -269
rect 5983 -341 5989 -307
rect 6023 -341 6029 -307
rect 5983 -379 6029 -341
rect 5983 -413 5989 -379
rect 6023 -413 6029 -379
rect 5983 -451 6029 -413
rect 5983 -485 5989 -451
rect 6023 -485 6029 -451
rect 5983 -523 6029 -485
rect 5983 -557 5989 -523
rect 6023 -557 6029 -523
rect 5983 -600 6029 -557
rect -5781 -647 -5373 -641
rect -5781 -681 -5738 -647
rect -5704 -681 -5666 -647
rect -5632 -681 -5594 -647
rect -5560 -681 -5522 -647
rect -5488 -681 -5450 -647
rect -5416 -681 -5373 -647
rect -5781 -687 -5373 -681
rect -4923 -647 -4515 -641
rect -4923 -681 -4880 -647
rect -4846 -681 -4808 -647
rect -4774 -681 -4736 -647
rect -4702 -681 -4664 -647
rect -4630 -681 -4592 -647
rect -4558 -681 -4515 -647
rect -4923 -687 -4515 -681
rect -4065 -647 -3657 -641
rect -4065 -681 -4022 -647
rect -3988 -681 -3950 -647
rect -3916 -681 -3878 -647
rect -3844 -681 -3806 -647
rect -3772 -681 -3734 -647
rect -3700 -681 -3657 -647
rect -4065 -687 -3657 -681
rect -3207 -647 -2799 -641
rect -3207 -681 -3164 -647
rect -3130 -681 -3092 -647
rect -3058 -681 -3020 -647
rect -2986 -681 -2948 -647
rect -2914 -681 -2876 -647
rect -2842 -681 -2799 -647
rect -3207 -687 -2799 -681
rect -2349 -647 -1941 -641
rect -2349 -681 -2306 -647
rect -2272 -681 -2234 -647
rect -2200 -681 -2162 -647
rect -2128 -681 -2090 -647
rect -2056 -681 -2018 -647
rect -1984 -681 -1941 -647
rect -2349 -687 -1941 -681
rect -1491 -647 -1083 -641
rect -1491 -681 -1448 -647
rect -1414 -681 -1376 -647
rect -1342 -681 -1304 -647
rect -1270 -681 -1232 -647
rect -1198 -681 -1160 -647
rect -1126 -681 -1083 -647
rect -1491 -687 -1083 -681
rect -633 -647 -225 -641
rect -633 -681 -590 -647
rect -556 -681 -518 -647
rect -484 -681 -446 -647
rect -412 -681 -374 -647
rect -340 -681 -302 -647
rect -268 -681 -225 -647
rect -633 -687 -225 -681
rect 225 -647 633 -641
rect 225 -681 268 -647
rect 302 -681 340 -647
rect 374 -681 412 -647
rect 446 -681 484 -647
rect 518 -681 556 -647
rect 590 -681 633 -647
rect 225 -687 633 -681
rect 1083 -647 1491 -641
rect 1083 -681 1126 -647
rect 1160 -681 1198 -647
rect 1232 -681 1270 -647
rect 1304 -681 1342 -647
rect 1376 -681 1414 -647
rect 1448 -681 1491 -647
rect 1083 -687 1491 -681
rect 1941 -647 2349 -641
rect 1941 -681 1984 -647
rect 2018 -681 2056 -647
rect 2090 -681 2128 -647
rect 2162 -681 2200 -647
rect 2234 -681 2272 -647
rect 2306 -681 2349 -647
rect 1941 -687 2349 -681
rect 2799 -647 3207 -641
rect 2799 -681 2842 -647
rect 2876 -681 2914 -647
rect 2948 -681 2986 -647
rect 3020 -681 3058 -647
rect 3092 -681 3130 -647
rect 3164 -681 3207 -647
rect 2799 -687 3207 -681
rect 3657 -647 4065 -641
rect 3657 -681 3700 -647
rect 3734 -681 3772 -647
rect 3806 -681 3844 -647
rect 3878 -681 3916 -647
rect 3950 -681 3988 -647
rect 4022 -681 4065 -647
rect 3657 -687 4065 -681
rect 4515 -647 4923 -641
rect 4515 -681 4558 -647
rect 4592 -681 4630 -647
rect 4664 -681 4702 -647
rect 4736 -681 4774 -647
rect 4808 -681 4846 -647
rect 4880 -681 4923 -647
rect 4515 -687 4923 -681
rect 5373 -647 5781 -641
rect 5373 -681 5416 -647
rect 5450 -681 5488 -647
rect 5522 -681 5560 -647
rect 5594 -681 5632 -647
rect 5666 -681 5704 -647
rect 5738 -681 5781 -647
rect 5373 -687 5781 -681
<< end >>
