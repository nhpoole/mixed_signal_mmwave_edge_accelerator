magic
tech sky130A
timestamp 1626486988
<< checkpaint >>
rect -720 -717 720 717
<< metal4 >>
rect -90 59 90 87
rect -90 -59 -59 59
rect 59 -59 90 59
rect -90 -87 90 -59
<< via4 >>
rect -59 -59 59 59
<< metal5 >>
rect -90 59 90 87
rect -90 -59 -59 59
rect 59 -59 90 59
rect -90 -87 90 -59
<< end >>
