magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1804 -1560 1804 1560
<< pwell >>
rect -544 -300 544 300
<< nmoslvt >>
rect -358 -100 -158 100
rect -100 -100 100 100
rect 158 -100 358 100
<< ndiff >>
rect -416 85 -358 100
rect -416 51 -404 85
rect -370 51 -358 85
rect -416 17 -358 51
rect -416 -17 -404 17
rect -370 -17 -358 17
rect -416 -51 -358 -17
rect -416 -85 -404 -51
rect -370 -85 -358 -51
rect -416 -100 -358 -85
rect -158 85 -100 100
rect -158 51 -146 85
rect -112 51 -100 85
rect -158 17 -100 51
rect -158 -17 -146 17
rect -112 -17 -100 17
rect -158 -51 -100 -17
rect -158 -85 -146 -51
rect -112 -85 -100 -51
rect -158 -100 -100 -85
rect 100 85 158 100
rect 100 51 112 85
rect 146 51 158 85
rect 100 17 158 51
rect 100 -17 112 17
rect 146 -17 158 17
rect 100 -51 158 -17
rect 100 -85 112 -51
rect 146 -85 158 -51
rect 100 -100 158 -85
rect 358 85 416 100
rect 358 51 370 85
rect 404 51 416 85
rect 358 17 416 51
rect 358 -17 370 17
rect 404 -17 416 17
rect 358 -51 416 -17
rect 358 -85 370 -51
rect 404 -85 416 -51
rect 358 -100 416 -85
<< ndiffc >>
rect -404 51 -370 85
rect -404 -17 -370 17
rect -404 -85 -370 -51
rect -146 51 -112 85
rect -146 -17 -112 17
rect -146 -85 -112 -51
rect 112 51 146 85
rect 112 -17 146 17
rect 112 -85 146 -51
rect 370 51 404 85
rect 370 -17 404 17
rect 370 -85 404 -51
<< psubdiff >>
rect -518 240 -391 274
rect -357 240 -323 274
rect -289 240 -255 274
rect -221 240 -187 274
rect -153 240 -119 274
rect -85 240 -51 274
rect -17 240 17 274
rect 51 240 85 274
rect 119 240 153 274
rect 187 240 221 274
rect 255 240 289 274
rect 323 240 357 274
rect 391 240 518 274
rect -518 153 -484 240
rect -518 85 -484 119
rect 484 153 518 240
rect -518 17 -484 51
rect -518 -51 -484 -17
rect -518 -119 -484 -85
rect 484 85 518 119
rect 484 17 518 51
rect 484 -51 518 -17
rect -518 -240 -484 -153
rect 484 -119 518 -85
rect 484 -240 518 -153
rect -518 -274 -391 -240
rect -357 -274 -323 -240
rect -289 -274 -255 -240
rect -221 -274 -187 -240
rect -153 -274 -119 -240
rect -85 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 85 -240
rect 119 -274 153 -240
rect 187 -274 221 -240
rect 255 -274 289 -240
rect 323 -274 357 -240
rect 391 -274 518 -240
<< psubdiffcont >>
rect -391 240 -357 274
rect -323 240 -289 274
rect -255 240 -221 274
rect -187 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 187 274
rect 221 240 255 274
rect 289 240 323 274
rect 357 240 391 274
rect -518 119 -484 153
rect 484 119 518 153
rect -518 51 -484 85
rect -518 -17 -484 17
rect -518 -85 -484 -51
rect 484 51 518 85
rect 484 -17 518 17
rect 484 -85 518 -51
rect -518 -153 -484 -119
rect 484 -153 518 -119
rect -391 -274 -357 -240
rect -323 -274 -289 -240
rect -255 -274 -221 -240
rect -187 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 187 -240
rect 221 -274 255 -240
rect 289 -274 323 -240
rect 357 -274 391 -240
<< poly >>
rect -324 172 -192 188
rect -324 155 -275 172
rect -358 138 -275 155
rect -241 155 -192 172
rect -66 172 66 188
rect -66 155 -17 172
rect -241 138 -158 155
rect -358 100 -158 138
rect -100 138 -17 155
rect 17 155 66 172
rect 192 172 324 188
rect 192 155 241 172
rect 17 138 100 155
rect -100 100 100 138
rect 158 138 241 155
rect 275 155 324 172
rect 275 138 358 155
rect 158 100 358 138
rect -358 -138 -158 -100
rect -358 -155 -275 -138
rect -324 -172 -275 -155
rect -241 -155 -158 -138
rect -100 -138 100 -100
rect -100 -155 -17 -138
rect -241 -172 -192 -155
rect -324 -188 -192 -172
rect -66 -172 -17 -155
rect 17 -155 100 -138
rect 158 -138 358 -100
rect 158 -155 241 -138
rect 17 -172 66 -155
rect -66 -188 66 -172
rect 192 -172 241 -155
rect 275 -155 358 -138
rect 275 -172 324 -155
rect 192 -188 324 -172
<< polycont >>
rect -275 138 -241 172
rect -17 138 17 172
rect 241 138 275 172
rect -275 -172 -241 -138
rect -17 -172 17 -138
rect 241 -172 275 -138
<< locali >>
rect -518 240 -391 274
rect -357 240 -323 274
rect -289 240 -255 274
rect -221 240 -187 274
rect -153 240 -119 274
rect -85 240 -51 274
rect -17 240 17 274
rect 51 240 85 274
rect 119 240 153 274
rect 187 240 221 274
rect 255 240 289 274
rect 323 240 357 274
rect 391 240 518 274
rect -518 153 -484 240
rect -324 138 -275 172
rect -241 138 -192 172
rect -66 138 -17 172
rect 17 138 66 172
rect 192 138 241 172
rect 275 138 324 172
rect 484 153 518 240
rect -518 85 -484 119
rect -518 17 -484 51
rect -518 -51 -484 -17
rect -518 -119 -484 -85
rect -404 85 -370 104
rect -404 17 -370 19
rect -404 -19 -370 -17
rect -404 -104 -370 -85
rect -146 85 -112 104
rect -146 17 -112 19
rect -146 -19 -112 -17
rect -146 -104 -112 -85
rect 112 85 146 104
rect 112 17 146 19
rect 112 -19 146 -17
rect 112 -104 146 -85
rect 370 85 404 104
rect 370 17 404 19
rect 370 -19 404 -17
rect 370 -104 404 -85
rect 484 85 518 119
rect 484 17 518 51
rect 484 -51 518 -17
rect 484 -119 518 -85
rect -518 -240 -484 -153
rect -324 -172 -275 -138
rect -241 -172 -192 -138
rect -66 -172 -17 -138
rect 17 -172 66 -138
rect 192 -172 241 -138
rect 275 -172 324 -138
rect 484 -240 518 -153
rect -518 -274 -391 -240
rect -357 -274 -323 -240
rect -289 -274 -255 -240
rect -221 -274 -187 -240
rect -153 -274 -119 -240
rect -85 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 85 -240
rect 119 -274 153 -240
rect 187 -274 221 -240
rect 255 -274 289 -240
rect 323 -274 357 -240
rect 391 -274 518 -240
<< viali >>
rect -275 138 -241 172
rect -17 138 17 172
rect 241 138 275 172
rect -404 51 -370 53
rect -404 19 -370 51
rect -404 -51 -370 -19
rect -404 -53 -370 -51
rect -146 51 -112 53
rect -146 19 -112 51
rect -146 -51 -112 -19
rect -146 -53 -112 -51
rect 112 51 146 53
rect 112 19 146 51
rect 112 -51 146 -19
rect 112 -53 146 -51
rect 370 51 404 53
rect 370 19 404 51
rect 370 -51 404 -19
rect 370 -53 404 -51
rect -275 -172 -241 -138
rect -17 -172 17 -138
rect 241 -172 275 -138
<< metal1 >>
rect -312 172 -204 178
rect -312 138 -275 172
rect -241 138 -204 172
rect -312 132 -204 138
rect -54 172 54 178
rect -54 138 -17 172
rect 17 138 54 172
rect -54 132 54 138
rect 204 172 312 178
rect 204 138 241 172
rect 275 138 312 172
rect 204 132 312 138
rect -410 53 -364 100
rect -410 19 -404 53
rect -370 19 -364 53
rect -410 -19 -364 19
rect -410 -53 -404 -19
rect -370 -53 -364 -19
rect -410 -100 -364 -53
rect -152 53 -106 100
rect -152 19 -146 53
rect -112 19 -106 53
rect -152 -19 -106 19
rect -152 -53 -146 -19
rect -112 -53 -106 -19
rect -152 -100 -106 -53
rect 106 53 152 100
rect 106 19 112 53
rect 146 19 152 53
rect 106 -19 152 19
rect 106 -53 112 -19
rect 146 -53 152 -19
rect 106 -100 152 -53
rect 364 53 410 100
rect 364 19 370 53
rect 404 19 410 53
rect 364 -19 410 19
rect 364 -53 370 -19
rect 404 -53 410 -19
rect 364 -100 410 -53
rect -312 -138 -204 -132
rect -312 -172 -275 -138
rect -241 -172 -204 -138
rect -312 -178 -204 -172
rect -54 -138 54 -132
rect -54 -172 -17 -138
rect 17 -172 54 -138
rect -54 -178 54 -172
rect 204 -138 312 -132
rect 204 -172 241 -138
rect 275 -172 312 -138
rect 204 -178 312 -172
<< properties >>
string FIXED_BBOX -501 -257 501 257
<< end >>
