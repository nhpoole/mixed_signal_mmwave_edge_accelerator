magic
tech sky130A
timestamp 1626065694
<< checkpaint >>
rect -732 -654 732 654
<< metal1 >>
rect -102 13 102 24
rect -102 -13 -93 13
rect -67 -13 -61 13
rect -35 -13 -29 13
rect -3 -13 3 13
rect 29 -13 35 13
rect 61 -13 67 13
rect 93 -13 102 13
rect -102 -24 102 -13
<< via1 >>
rect -93 -13 -67 13
rect -61 -13 -35 13
rect -29 -13 -3 13
rect 3 -13 29 13
rect 35 -13 61 13
rect 67 -13 93 13
<< metal2 >>
rect -102 13 102 24
rect -102 -13 -93 13
rect -67 -13 -61 13
rect -35 -13 -29 13
rect -3 -13 3 13
rect 29 -13 35 13
rect 61 -13 67 13
rect 93 -13 102 13
rect -102 -24 102 -13
<< end >>
