magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< nwell >>
rect -36 538 512 1177
<< poly >>
rect 114 567 144 761
rect 81 501 144 567
rect 114 255 144 501
<< locali >>
rect 0 1103 476 1137
rect 62 910 96 1103
rect 64 501 98 567
rect 166 551 200 976
rect 270 910 304 1103
rect 374 1028 408 1103
rect 166 517 217 551
rect 166 92 200 517
rect 62 17 96 92
rect 270 17 304 92
rect 374 17 408 92
rect 0 -17 476 17
use contact_15  contact_15_0
timestamp 1624494425
transform 1 0 48 0 1 501
box 0 0 66 66
use contact_28  contact_28_0
timestamp 1624494425
transform 1 0 366 0 1 51
box -26 -26 76 108
use contact_27  contact_27_0
timestamp 1624494425
transform 1 0 366 0 1 987
box -59 -43 109 125
use nmos_m2_w0_740_sli_dli_da_p  nmos_m2_w0_740_sli_dli_da_p_0
timestamp 1624494425
transform 1 0 54 0 1 51
box -26 -26 284 204
use pmos_m2_w1_260_sli_dli_da_p  pmos_m2_w1_260_sli_dli_da_p_0
timestamp 1624494425
transform 1 0 54 0 1 817
box -59 -56 317 306
<< labels >>
rlabel locali s 81 534 81 534 4 A
rlabel locali s 200 534 200 534 4 Z
rlabel locali s 238 0 238 0 4 gnd
rlabel locali s 238 1120 238 1120 4 vdd
<< properties >>
string FIXED_BBOX 0 0 476 1120
<< end >>
