magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -2605 -1548 2605 1548
<< pwell >>
rect -1345 -226 1345 226
<< nmos >>
rect -1261 -200 -1061 200
rect -1003 -200 -803 200
rect -745 -200 -545 200
rect -487 -200 -287 200
rect -229 -200 -29 200
rect 29 -200 229 200
rect 287 -200 487 200
rect 545 -200 745 200
rect 803 -200 1003 200
rect 1061 -200 1261 200
<< ndiff >>
rect -1319 187 -1261 200
rect -1319 153 -1307 187
rect -1273 153 -1261 187
rect -1319 119 -1261 153
rect -1319 85 -1307 119
rect -1273 85 -1261 119
rect -1319 51 -1261 85
rect -1319 17 -1307 51
rect -1273 17 -1261 51
rect -1319 -17 -1261 17
rect -1319 -51 -1307 -17
rect -1273 -51 -1261 -17
rect -1319 -85 -1261 -51
rect -1319 -119 -1307 -85
rect -1273 -119 -1261 -85
rect -1319 -153 -1261 -119
rect -1319 -187 -1307 -153
rect -1273 -187 -1261 -153
rect -1319 -200 -1261 -187
rect -1061 187 -1003 200
rect -1061 153 -1049 187
rect -1015 153 -1003 187
rect -1061 119 -1003 153
rect -1061 85 -1049 119
rect -1015 85 -1003 119
rect -1061 51 -1003 85
rect -1061 17 -1049 51
rect -1015 17 -1003 51
rect -1061 -17 -1003 17
rect -1061 -51 -1049 -17
rect -1015 -51 -1003 -17
rect -1061 -85 -1003 -51
rect -1061 -119 -1049 -85
rect -1015 -119 -1003 -85
rect -1061 -153 -1003 -119
rect -1061 -187 -1049 -153
rect -1015 -187 -1003 -153
rect -1061 -200 -1003 -187
rect -803 187 -745 200
rect -803 153 -791 187
rect -757 153 -745 187
rect -803 119 -745 153
rect -803 85 -791 119
rect -757 85 -745 119
rect -803 51 -745 85
rect -803 17 -791 51
rect -757 17 -745 51
rect -803 -17 -745 17
rect -803 -51 -791 -17
rect -757 -51 -745 -17
rect -803 -85 -745 -51
rect -803 -119 -791 -85
rect -757 -119 -745 -85
rect -803 -153 -745 -119
rect -803 -187 -791 -153
rect -757 -187 -745 -153
rect -803 -200 -745 -187
rect -545 187 -487 200
rect -545 153 -533 187
rect -499 153 -487 187
rect -545 119 -487 153
rect -545 85 -533 119
rect -499 85 -487 119
rect -545 51 -487 85
rect -545 17 -533 51
rect -499 17 -487 51
rect -545 -17 -487 17
rect -545 -51 -533 -17
rect -499 -51 -487 -17
rect -545 -85 -487 -51
rect -545 -119 -533 -85
rect -499 -119 -487 -85
rect -545 -153 -487 -119
rect -545 -187 -533 -153
rect -499 -187 -487 -153
rect -545 -200 -487 -187
rect -287 187 -229 200
rect -287 153 -275 187
rect -241 153 -229 187
rect -287 119 -229 153
rect -287 85 -275 119
rect -241 85 -229 119
rect -287 51 -229 85
rect -287 17 -275 51
rect -241 17 -229 51
rect -287 -17 -229 17
rect -287 -51 -275 -17
rect -241 -51 -229 -17
rect -287 -85 -229 -51
rect -287 -119 -275 -85
rect -241 -119 -229 -85
rect -287 -153 -229 -119
rect -287 -187 -275 -153
rect -241 -187 -229 -153
rect -287 -200 -229 -187
rect -29 187 29 200
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -200 29 -187
rect 229 187 287 200
rect 229 153 241 187
rect 275 153 287 187
rect 229 119 287 153
rect 229 85 241 119
rect 275 85 287 119
rect 229 51 287 85
rect 229 17 241 51
rect 275 17 287 51
rect 229 -17 287 17
rect 229 -51 241 -17
rect 275 -51 287 -17
rect 229 -85 287 -51
rect 229 -119 241 -85
rect 275 -119 287 -85
rect 229 -153 287 -119
rect 229 -187 241 -153
rect 275 -187 287 -153
rect 229 -200 287 -187
rect 487 187 545 200
rect 487 153 499 187
rect 533 153 545 187
rect 487 119 545 153
rect 487 85 499 119
rect 533 85 545 119
rect 487 51 545 85
rect 487 17 499 51
rect 533 17 545 51
rect 487 -17 545 17
rect 487 -51 499 -17
rect 533 -51 545 -17
rect 487 -85 545 -51
rect 487 -119 499 -85
rect 533 -119 545 -85
rect 487 -153 545 -119
rect 487 -187 499 -153
rect 533 -187 545 -153
rect 487 -200 545 -187
rect 745 187 803 200
rect 745 153 757 187
rect 791 153 803 187
rect 745 119 803 153
rect 745 85 757 119
rect 791 85 803 119
rect 745 51 803 85
rect 745 17 757 51
rect 791 17 803 51
rect 745 -17 803 17
rect 745 -51 757 -17
rect 791 -51 803 -17
rect 745 -85 803 -51
rect 745 -119 757 -85
rect 791 -119 803 -85
rect 745 -153 803 -119
rect 745 -187 757 -153
rect 791 -187 803 -153
rect 745 -200 803 -187
rect 1003 187 1061 200
rect 1003 153 1015 187
rect 1049 153 1061 187
rect 1003 119 1061 153
rect 1003 85 1015 119
rect 1049 85 1061 119
rect 1003 51 1061 85
rect 1003 17 1015 51
rect 1049 17 1061 51
rect 1003 -17 1061 17
rect 1003 -51 1015 -17
rect 1049 -51 1061 -17
rect 1003 -85 1061 -51
rect 1003 -119 1015 -85
rect 1049 -119 1061 -85
rect 1003 -153 1061 -119
rect 1003 -187 1015 -153
rect 1049 -187 1061 -153
rect 1003 -200 1061 -187
rect 1261 187 1319 200
rect 1261 153 1273 187
rect 1307 153 1319 187
rect 1261 119 1319 153
rect 1261 85 1273 119
rect 1307 85 1319 119
rect 1261 51 1319 85
rect 1261 17 1273 51
rect 1307 17 1319 51
rect 1261 -17 1319 17
rect 1261 -51 1273 -17
rect 1307 -51 1319 -17
rect 1261 -85 1319 -51
rect 1261 -119 1273 -85
rect 1307 -119 1319 -85
rect 1261 -153 1319 -119
rect 1261 -187 1273 -153
rect 1307 -187 1319 -153
rect 1261 -200 1319 -187
<< ndiffc >>
rect -1307 153 -1273 187
rect -1307 85 -1273 119
rect -1307 17 -1273 51
rect -1307 -51 -1273 -17
rect -1307 -119 -1273 -85
rect -1307 -187 -1273 -153
rect -1049 153 -1015 187
rect -1049 85 -1015 119
rect -1049 17 -1015 51
rect -1049 -51 -1015 -17
rect -1049 -119 -1015 -85
rect -1049 -187 -1015 -153
rect -791 153 -757 187
rect -791 85 -757 119
rect -791 17 -757 51
rect -791 -51 -757 -17
rect -791 -119 -757 -85
rect -791 -187 -757 -153
rect -533 153 -499 187
rect -533 85 -499 119
rect -533 17 -499 51
rect -533 -51 -499 -17
rect -533 -119 -499 -85
rect -533 -187 -499 -153
rect -275 153 -241 187
rect -275 85 -241 119
rect -275 17 -241 51
rect -275 -51 -241 -17
rect -275 -119 -241 -85
rect -275 -187 -241 -153
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect 241 153 275 187
rect 241 85 275 119
rect 241 17 275 51
rect 241 -51 275 -17
rect 241 -119 275 -85
rect 241 -187 275 -153
rect 499 153 533 187
rect 499 85 533 119
rect 499 17 533 51
rect 499 -51 533 -17
rect 499 -119 533 -85
rect 499 -187 533 -153
rect 757 153 791 187
rect 757 85 791 119
rect 757 17 791 51
rect 757 -51 791 -17
rect 757 -119 791 -85
rect 757 -187 791 -153
rect 1015 153 1049 187
rect 1015 85 1049 119
rect 1015 17 1049 51
rect 1015 -51 1049 -17
rect 1015 -119 1049 -85
rect 1015 -187 1049 -153
rect 1273 153 1307 187
rect 1273 85 1307 119
rect 1273 17 1307 51
rect 1273 -51 1307 -17
rect 1273 -119 1307 -85
rect 1273 -187 1307 -153
<< poly >>
rect -1227 272 -1095 288
rect -1227 255 -1178 272
rect -1261 238 -1178 255
rect -1144 255 -1095 272
rect -969 272 -837 288
rect -969 255 -920 272
rect -1144 238 -1061 255
rect -1261 200 -1061 238
rect -1003 238 -920 255
rect -886 255 -837 272
rect -711 272 -579 288
rect -711 255 -662 272
rect -886 238 -803 255
rect -1003 200 -803 238
rect -745 238 -662 255
rect -628 255 -579 272
rect -453 272 -321 288
rect -453 255 -404 272
rect -628 238 -545 255
rect -745 200 -545 238
rect -487 238 -404 255
rect -370 255 -321 272
rect -195 272 -63 288
rect -195 255 -146 272
rect -370 238 -287 255
rect -487 200 -287 238
rect -229 238 -146 255
rect -112 255 -63 272
rect 63 272 195 288
rect 63 255 112 272
rect -112 238 -29 255
rect -229 200 -29 238
rect 29 238 112 255
rect 146 255 195 272
rect 321 272 453 288
rect 321 255 370 272
rect 146 238 229 255
rect 29 200 229 238
rect 287 238 370 255
rect 404 255 453 272
rect 579 272 711 288
rect 579 255 628 272
rect 404 238 487 255
rect 287 200 487 238
rect 545 238 628 255
rect 662 255 711 272
rect 837 272 969 288
rect 837 255 886 272
rect 662 238 745 255
rect 545 200 745 238
rect 803 238 886 255
rect 920 255 969 272
rect 1095 272 1227 288
rect 1095 255 1144 272
rect 920 238 1003 255
rect 803 200 1003 238
rect 1061 238 1144 255
rect 1178 255 1227 272
rect 1178 238 1261 255
rect 1061 200 1261 238
rect -1261 -238 -1061 -200
rect -1261 -255 -1178 -238
rect -1227 -272 -1178 -255
rect -1144 -255 -1061 -238
rect -1003 -238 -803 -200
rect -1003 -255 -920 -238
rect -1144 -272 -1095 -255
rect -1227 -288 -1095 -272
rect -969 -272 -920 -255
rect -886 -255 -803 -238
rect -745 -238 -545 -200
rect -745 -255 -662 -238
rect -886 -272 -837 -255
rect -969 -288 -837 -272
rect -711 -272 -662 -255
rect -628 -255 -545 -238
rect -487 -238 -287 -200
rect -487 -255 -404 -238
rect -628 -272 -579 -255
rect -711 -288 -579 -272
rect -453 -272 -404 -255
rect -370 -255 -287 -238
rect -229 -238 -29 -200
rect -229 -255 -146 -238
rect -370 -272 -321 -255
rect -453 -288 -321 -272
rect -195 -272 -146 -255
rect -112 -255 -29 -238
rect 29 -238 229 -200
rect 29 -255 112 -238
rect -112 -272 -63 -255
rect -195 -288 -63 -272
rect 63 -272 112 -255
rect 146 -255 229 -238
rect 287 -238 487 -200
rect 287 -255 370 -238
rect 146 -272 195 -255
rect 63 -288 195 -272
rect 321 -272 370 -255
rect 404 -255 487 -238
rect 545 -238 745 -200
rect 545 -255 628 -238
rect 404 -272 453 -255
rect 321 -288 453 -272
rect 579 -272 628 -255
rect 662 -255 745 -238
rect 803 -238 1003 -200
rect 803 -255 886 -238
rect 662 -272 711 -255
rect 579 -288 711 -272
rect 837 -272 886 -255
rect 920 -255 1003 -238
rect 1061 -238 1261 -200
rect 1061 -255 1144 -238
rect 920 -272 969 -255
rect 837 -288 969 -272
rect 1095 -272 1144 -255
rect 1178 -255 1261 -238
rect 1178 -272 1227 -255
rect 1095 -288 1227 -272
<< polycont >>
rect -1178 238 -1144 272
rect -920 238 -886 272
rect -662 238 -628 272
rect -404 238 -370 272
rect -146 238 -112 272
rect 112 238 146 272
rect 370 238 404 272
rect 628 238 662 272
rect 886 238 920 272
rect 1144 238 1178 272
rect -1178 -272 -1144 -238
rect -920 -272 -886 -238
rect -662 -272 -628 -238
rect -404 -272 -370 -238
rect -146 -272 -112 -238
rect 112 -272 146 -238
rect 370 -272 404 -238
rect 628 -272 662 -238
rect 886 -272 920 -238
rect 1144 -272 1178 -238
<< locali >>
rect -1227 238 -1178 272
rect -1144 238 -1095 272
rect -969 238 -920 272
rect -886 238 -837 272
rect -711 238 -662 272
rect -628 238 -579 272
rect -453 238 -404 272
rect -370 238 -321 272
rect -195 238 -146 272
rect -112 238 -63 272
rect 63 238 112 272
rect 146 238 195 272
rect 321 238 370 272
rect 404 238 453 272
rect 579 238 628 272
rect 662 238 711 272
rect 837 238 886 272
rect 920 238 969 272
rect 1095 238 1144 272
rect 1178 238 1227 272
rect -1307 187 -1273 204
rect -1307 119 -1273 127
rect -1307 51 -1273 55
rect -1307 -55 -1273 -51
rect -1307 -127 -1273 -119
rect -1307 -204 -1273 -187
rect -1049 187 -1015 204
rect -1049 119 -1015 127
rect -1049 51 -1015 55
rect -1049 -55 -1015 -51
rect -1049 -127 -1015 -119
rect -1049 -204 -1015 -187
rect -791 187 -757 204
rect -791 119 -757 127
rect -791 51 -757 55
rect -791 -55 -757 -51
rect -791 -127 -757 -119
rect -791 -204 -757 -187
rect -533 187 -499 204
rect -533 119 -499 127
rect -533 51 -499 55
rect -533 -55 -499 -51
rect -533 -127 -499 -119
rect -533 -204 -499 -187
rect -275 187 -241 204
rect -275 119 -241 127
rect -275 51 -241 55
rect -275 -55 -241 -51
rect -275 -127 -241 -119
rect -275 -204 -241 -187
rect -17 187 17 204
rect -17 119 17 127
rect -17 51 17 55
rect -17 -55 17 -51
rect -17 -127 17 -119
rect -17 -204 17 -187
rect 241 187 275 204
rect 241 119 275 127
rect 241 51 275 55
rect 241 -55 275 -51
rect 241 -127 275 -119
rect 241 -204 275 -187
rect 499 187 533 204
rect 499 119 533 127
rect 499 51 533 55
rect 499 -55 533 -51
rect 499 -127 533 -119
rect 499 -204 533 -187
rect 757 187 791 204
rect 757 119 791 127
rect 757 51 791 55
rect 757 -55 791 -51
rect 757 -127 791 -119
rect 757 -204 791 -187
rect 1015 187 1049 204
rect 1015 119 1049 127
rect 1015 51 1049 55
rect 1015 -55 1049 -51
rect 1015 -127 1049 -119
rect 1015 -204 1049 -187
rect 1273 187 1307 204
rect 1273 119 1307 127
rect 1273 51 1307 55
rect 1273 -55 1307 -51
rect 1273 -127 1307 -119
rect 1273 -204 1307 -187
rect -1227 -272 -1178 -238
rect -1144 -272 -1095 -238
rect -969 -272 -920 -238
rect -886 -272 -837 -238
rect -711 -272 -662 -238
rect -628 -272 -579 -238
rect -453 -272 -404 -238
rect -370 -272 -321 -238
rect -195 -272 -146 -238
rect -112 -272 -63 -238
rect 63 -272 112 -238
rect 146 -272 195 -238
rect 321 -272 370 -238
rect 404 -272 453 -238
rect 579 -272 628 -238
rect 662 -272 711 -238
rect 837 -272 886 -238
rect 920 -272 969 -238
rect 1095 -272 1144 -238
rect 1178 -272 1227 -238
<< viali >>
rect -1178 238 -1144 272
rect -920 238 -886 272
rect -662 238 -628 272
rect -404 238 -370 272
rect -146 238 -112 272
rect 112 238 146 272
rect 370 238 404 272
rect 628 238 662 272
rect 886 238 920 272
rect 1144 238 1178 272
rect -1307 153 -1273 161
rect -1307 127 -1273 153
rect -1307 85 -1273 89
rect -1307 55 -1273 85
rect -1307 -17 -1273 17
rect -1307 -85 -1273 -55
rect -1307 -89 -1273 -85
rect -1307 -153 -1273 -127
rect -1307 -161 -1273 -153
rect -1049 153 -1015 161
rect -1049 127 -1015 153
rect -1049 85 -1015 89
rect -1049 55 -1015 85
rect -1049 -17 -1015 17
rect -1049 -85 -1015 -55
rect -1049 -89 -1015 -85
rect -1049 -153 -1015 -127
rect -1049 -161 -1015 -153
rect -791 153 -757 161
rect -791 127 -757 153
rect -791 85 -757 89
rect -791 55 -757 85
rect -791 -17 -757 17
rect -791 -85 -757 -55
rect -791 -89 -757 -85
rect -791 -153 -757 -127
rect -791 -161 -757 -153
rect -533 153 -499 161
rect -533 127 -499 153
rect -533 85 -499 89
rect -533 55 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -55
rect -533 -89 -499 -85
rect -533 -153 -499 -127
rect -533 -161 -499 -153
rect -275 153 -241 161
rect -275 127 -241 153
rect -275 85 -241 89
rect -275 55 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -55
rect -275 -89 -241 -85
rect -275 -153 -241 -127
rect -275 -161 -241 -153
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect 241 153 275 161
rect 241 127 275 153
rect 241 85 275 89
rect 241 55 275 85
rect 241 -17 275 17
rect 241 -85 275 -55
rect 241 -89 275 -85
rect 241 -153 275 -127
rect 241 -161 275 -153
rect 499 153 533 161
rect 499 127 533 153
rect 499 85 533 89
rect 499 55 533 85
rect 499 -17 533 17
rect 499 -85 533 -55
rect 499 -89 533 -85
rect 499 -153 533 -127
rect 499 -161 533 -153
rect 757 153 791 161
rect 757 127 791 153
rect 757 85 791 89
rect 757 55 791 85
rect 757 -17 791 17
rect 757 -85 791 -55
rect 757 -89 791 -85
rect 757 -153 791 -127
rect 757 -161 791 -153
rect 1015 153 1049 161
rect 1015 127 1049 153
rect 1015 85 1049 89
rect 1015 55 1049 85
rect 1015 -17 1049 17
rect 1015 -85 1049 -55
rect 1015 -89 1049 -85
rect 1015 -153 1049 -127
rect 1015 -161 1049 -153
rect 1273 153 1307 161
rect 1273 127 1307 153
rect 1273 85 1307 89
rect 1273 55 1307 85
rect 1273 -17 1307 17
rect 1273 -85 1307 -55
rect 1273 -89 1307 -85
rect 1273 -153 1307 -127
rect 1273 -161 1307 -153
rect -1178 -272 -1144 -238
rect -920 -272 -886 -238
rect -662 -272 -628 -238
rect -404 -272 -370 -238
rect -146 -272 -112 -238
rect 112 -272 146 -238
rect 370 -272 404 -238
rect 628 -272 662 -238
rect 886 -272 920 -238
rect 1144 -272 1178 -238
<< metal1 >>
rect -1215 272 -1107 278
rect -1215 238 -1178 272
rect -1144 238 -1107 272
rect -1215 232 -1107 238
rect -957 272 -849 278
rect -957 238 -920 272
rect -886 238 -849 272
rect -957 232 -849 238
rect -699 272 -591 278
rect -699 238 -662 272
rect -628 238 -591 272
rect -699 232 -591 238
rect -441 272 -333 278
rect -441 238 -404 272
rect -370 238 -333 272
rect -441 232 -333 238
rect -183 272 -75 278
rect -183 238 -146 272
rect -112 238 -75 272
rect -183 232 -75 238
rect 75 272 183 278
rect 75 238 112 272
rect 146 238 183 272
rect 75 232 183 238
rect 333 272 441 278
rect 333 238 370 272
rect 404 238 441 272
rect 333 232 441 238
rect 591 272 699 278
rect 591 238 628 272
rect 662 238 699 272
rect 591 232 699 238
rect 849 272 957 278
rect 849 238 886 272
rect 920 238 957 272
rect 849 232 957 238
rect 1107 272 1215 278
rect 1107 238 1144 272
rect 1178 238 1215 272
rect 1107 232 1215 238
rect -1313 161 -1267 200
rect -1313 127 -1307 161
rect -1273 127 -1267 161
rect -1313 89 -1267 127
rect -1313 55 -1307 89
rect -1273 55 -1267 89
rect -1313 17 -1267 55
rect -1313 -17 -1307 17
rect -1273 -17 -1267 17
rect -1313 -55 -1267 -17
rect -1313 -89 -1307 -55
rect -1273 -89 -1267 -55
rect -1313 -127 -1267 -89
rect -1313 -161 -1307 -127
rect -1273 -161 -1267 -127
rect -1313 -200 -1267 -161
rect -1055 161 -1009 200
rect -1055 127 -1049 161
rect -1015 127 -1009 161
rect -1055 89 -1009 127
rect -1055 55 -1049 89
rect -1015 55 -1009 89
rect -1055 17 -1009 55
rect -1055 -17 -1049 17
rect -1015 -17 -1009 17
rect -1055 -55 -1009 -17
rect -1055 -89 -1049 -55
rect -1015 -89 -1009 -55
rect -1055 -127 -1009 -89
rect -1055 -161 -1049 -127
rect -1015 -161 -1009 -127
rect -1055 -200 -1009 -161
rect -797 161 -751 200
rect -797 127 -791 161
rect -757 127 -751 161
rect -797 89 -751 127
rect -797 55 -791 89
rect -757 55 -751 89
rect -797 17 -751 55
rect -797 -17 -791 17
rect -757 -17 -751 17
rect -797 -55 -751 -17
rect -797 -89 -791 -55
rect -757 -89 -751 -55
rect -797 -127 -751 -89
rect -797 -161 -791 -127
rect -757 -161 -751 -127
rect -797 -200 -751 -161
rect -539 161 -493 200
rect -539 127 -533 161
rect -499 127 -493 161
rect -539 89 -493 127
rect -539 55 -533 89
rect -499 55 -493 89
rect -539 17 -493 55
rect -539 -17 -533 17
rect -499 -17 -493 17
rect -539 -55 -493 -17
rect -539 -89 -533 -55
rect -499 -89 -493 -55
rect -539 -127 -493 -89
rect -539 -161 -533 -127
rect -499 -161 -493 -127
rect -539 -200 -493 -161
rect -281 161 -235 200
rect -281 127 -275 161
rect -241 127 -235 161
rect -281 89 -235 127
rect -281 55 -275 89
rect -241 55 -235 89
rect -281 17 -235 55
rect -281 -17 -275 17
rect -241 -17 -235 17
rect -281 -55 -235 -17
rect -281 -89 -275 -55
rect -241 -89 -235 -55
rect -281 -127 -235 -89
rect -281 -161 -275 -127
rect -241 -161 -235 -127
rect -281 -200 -235 -161
rect -23 161 23 200
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -200 23 -161
rect 235 161 281 200
rect 235 127 241 161
rect 275 127 281 161
rect 235 89 281 127
rect 235 55 241 89
rect 275 55 281 89
rect 235 17 281 55
rect 235 -17 241 17
rect 275 -17 281 17
rect 235 -55 281 -17
rect 235 -89 241 -55
rect 275 -89 281 -55
rect 235 -127 281 -89
rect 235 -161 241 -127
rect 275 -161 281 -127
rect 235 -200 281 -161
rect 493 161 539 200
rect 493 127 499 161
rect 533 127 539 161
rect 493 89 539 127
rect 493 55 499 89
rect 533 55 539 89
rect 493 17 539 55
rect 493 -17 499 17
rect 533 -17 539 17
rect 493 -55 539 -17
rect 493 -89 499 -55
rect 533 -89 539 -55
rect 493 -127 539 -89
rect 493 -161 499 -127
rect 533 -161 539 -127
rect 493 -200 539 -161
rect 751 161 797 200
rect 751 127 757 161
rect 791 127 797 161
rect 751 89 797 127
rect 751 55 757 89
rect 791 55 797 89
rect 751 17 797 55
rect 751 -17 757 17
rect 791 -17 797 17
rect 751 -55 797 -17
rect 751 -89 757 -55
rect 791 -89 797 -55
rect 751 -127 797 -89
rect 751 -161 757 -127
rect 791 -161 797 -127
rect 751 -200 797 -161
rect 1009 161 1055 200
rect 1009 127 1015 161
rect 1049 127 1055 161
rect 1009 89 1055 127
rect 1009 55 1015 89
rect 1049 55 1055 89
rect 1009 17 1055 55
rect 1009 -17 1015 17
rect 1049 -17 1055 17
rect 1009 -55 1055 -17
rect 1009 -89 1015 -55
rect 1049 -89 1055 -55
rect 1009 -127 1055 -89
rect 1009 -161 1015 -127
rect 1049 -161 1055 -127
rect 1009 -200 1055 -161
rect 1267 161 1313 200
rect 1267 127 1273 161
rect 1307 127 1313 161
rect 1267 89 1313 127
rect 1267 55 1273 89
rect 1307 55 1313 89
rect 1267 17 1313 55
rect 1267 -17 1273 17
rect 1307 -17 1313 17
rect 1267 -55 1313 -17
rect 1267 -89 1273 -55
rect 1307 -89 1313 -55
rect 1267 -127 1313 -89
rect 1267 -161 1273 -127
rect 1307 -161 1313 -127
rect 1267 -200 1313 -161
rect -1215 -238 -1107 -232
rect -1215 -272 -1178 -238
rect -1144 -272 -1107 -238
rect -1215 -278 -1107 -272
rect -957 -238 -849 -232
rect -957 -272 -920 -238
rect -886 -272 -849 -238
rect -957 -278 -849 -272
rect -699 -238 -591 -232
rect -699 -272 -662 -238
rect -628 -272 -591 -238
rect -699 -278 -591 -272
rect -441 -238 -333 -232
rect -441 -272 -404 -238
rect -370 -272 -333 -238
rect -441 -278 -333 -272
rect -183 -238 -75 -232
rect -183 -272 -146 -238
rect -112 -272 -75 -238
rect -183 -278 -75 -272
rect 75 -238 183 -232
rect 75 -272 112 -238
rect 146 -272 183 -238
rect 75 -278 183 -272
rect 333 -238 441 -232
rect 333 -272 370 -238
rect 404 -272 441 -238
rect 333 -278 441 -272
rect 591 -238 699 -232
rect 591 -272 628 -238
rect 662 -272 699 -238
rect 591 -278 699 -272
rect 849 -238 957 -232
rect 849 -272 886 -238
rect 920 -272 957 -238
rect 849 -278 957 -272
rect 1107 -238 1215 -232
rect 1107 -272 1144 -238
rect 1178 -272 1215 -238
rect 1107 -278 1215 -272
<< end >>
