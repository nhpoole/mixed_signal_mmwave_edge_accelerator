magic
tech sky130A
timestamp 1622079218
<< viali >>
rect 859 104 883 128
rect 40 58 64 82
rect 163 43 187 67
rect 717 -2 741 22
<< metal1 >>
rect -77 196 32 244
rect 853 128 996 131
rect 853 104 859 128
rect 883 104 996 128
rect 853 101 996 104
rect -33 82 70 85
rect -33 58 40 82
rect 64 58 70 82
rect -33 55 70 58
rect 157 67 193 70
rect 157 43 163 67
rect 187 43 193 67
rect 157 40 193 43
rect 157 30 190 40
rect -82 0 190 30
rect 711 22 939 25
rect 711 -2 717 22
rect 741 -2 939 22
rect 711 -5 939 -2
rect -67 -76 30 -28
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_0
timestamp 1620951057
transform 1 0 24 0 1 -52
box -19 -24 893 296
<< labels >>
flabel metal1 -13 64 -10 68 1 FreeSans 240 0 0 0 CLK
flabel metal1 -63 10 -60 14 1 FreeSans 240 0 0 0 D
flabel metal1 -30 -53 -28 -50 1 FreeSans 240 0 0 0 VSS
flabel metal1 -45 218 -44 220 1 FreeSans 240 0 0 0 VDD
flabel metal1 966 113 968 115 1 FreeSans 240 0 0 0 QB
flabel metal1 920 11 921 12 1 FreeSans 240 0 0 0 Q
<< end >>
