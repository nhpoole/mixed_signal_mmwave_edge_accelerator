magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1296 -1309 3632 2727
<< metal1 >>
rect 552 1388 616 1440
rect 1720 1388 1784 1440
rect 552 -26 616 26
rect 1720 -26 1784 26
<< metal2 >>
rect 137 538 203 590
rect 369 0 397 1414
rect 556 1390 612 1438
rect 1082 609 1148 661
rect 1305 538 1371 590
rect 556 -24 612 24
rect 1537 0 1565 1414
rect 1724 1390 1780 1438
rect 2250 609 2316 661
rect 1724 -24 1780 24
<< metal3 >>
rect 535 1365 633 1463
rect 1703 1365 1801 1463
rect 0 278 2336 338
rect 535 -49 633 49
rect 1703 -49 1801 49
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_1
timestamp 1626486988
transform 1 0 0 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_0
timestamp 1626486988
transform 1 0 1168 0 1 0
box -36 -43 1204 1467
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_5
timestamp 1626486988
transform 1 0 551 0 1 1377
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_4
timestamp 1626486988
transform 1 0 551 0 1 -37
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_3
timestamp 1626486988
transform 1 0 1719 0 1 1377
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_2
timestamp 1626486988
transform 1 0 1719 0 1 -37
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1626486988
transform 1 0 363 0 1 271
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1626486988
transform 1 0 1531 0 1 271
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_3
timestamp 1626486988
transform 1 0 552 0 1 1382
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1626486988
transform 1 0 552 0 1 -32
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1626486988
transform 1 0 1720 0 1 1382
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1626486988
transform 1 0 1720 0 1 -32
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_3
timestamp 1626486988
transform 1 0 555 0 1 1381
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_2
timestamp 1626486988
transform 1 0 555 0 1 -33
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1
timestamp 1626486988
transform 1 0 1723 0 1 1381
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_0
timestamp 1626486988
transform 1 0 1723 0 1 -33
box 0 0 58 66
<< labels >>
rlabel metal3 s 535 1365 633 1463 4 vdd
rlabel metal3 s 1703 1365 1801 1463 4 vdd
rlabel metal3 s 535 -49 633 49 4 gnd
rlabel metal3 s 1703 -49 1801 49 4 gnd
rlabel metal3 s 0 278 2336 338 4 clk
rlabel metal2 s 137 538 203 590 4 din_0
rlabel metal2 s 1082 609 1148 661 4 dout_0
rlabel metal2 s 1305 538 1371 590 4 din_1
rlabel metal2 s 2250 609 2316 661 4 dout_1
<< properties >>
string FIXED_BBOX 0 0 2336 1414
<< end >>
