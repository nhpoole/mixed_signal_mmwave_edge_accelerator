* Stimulus file.

.param Itail_filt=0.1u Ibias_filt=0.1u Ccomp_filt=0p vcmdes=1 vcmdes_filt=1.1 vincm=1.1 vsig=0 vdd=1.8
+   Wp=16 Wn=2 Wpcm=64 Wncm=4 Wbias=1 Lbias_diff=4.8 Lbias_se=6.4 nfactorL=1 nfactorW=6 K=1 K2=0.5
+   Cacc=1n Rhpf=10meg Kcap=10000 Rbase=100 Cfilt=5p Cmult=1p

vdd VDD GND 'vdd'
vin vin GND sin('vdd/2' '0.2*vdd/2' 50 0)
vincm vincm GND 'vincm'
vocm vocm GND 'vcmdes'
vgc0 gain_ctrl_0 GND 0
vgc1 gain_ctrl_1 GND 0
*e1 vbuf 0 vcap vbuf 10000

.ic v(net6)='vcmdes'
.ic v(net3)='vcmdes'
*.options savecurrents
.save all @r8[i] @r9[i] @r10[i] @r11[i] @c17[i] @c21[i] @c16[i] @c19[i]
*.save vin vhpf votap votam vop vom vcm vip vim
.tran 10u 200m

.control
run
write input_amplifier_tran.raw
quit
.endc
