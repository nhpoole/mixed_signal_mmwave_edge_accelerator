magic
tech sky130A
magscale 1 2
timestamp 1621829047
<< nwell >>
rect -2355 -700 2355 700
<< pmoshvt >>
rect -2261 -600 -1861 600
rect -1803 -600 -1403 600
rect -1345 -600 -945 600
rect -887 -600 -487 600
rect -429 -600 -29 600
rect 29 -600 429 600
rect 487 -600 887 600
rect 945 -600 1345 600
rect 1403 -600 1803 600
rect 1861 -600 2261 600
<< pdiff >>
rect -2319 588 -2261 600
rect -2319 -588 -2307 588
rect -2273 -588 -2261 588
rect -2319 -600 -2261 -588
rect -1861 588 -1803 600
rect -1861 -588 -1849 588
rect -1815 -588 -1803 588
rect -1861 -600 -1803 -588
rect -1403 588 -1345 600
rect -1403 -588 -1391 588
rect -1357 -588 -1345 588
rect -1403 -600 -1345 -588
rect -945 588 -887 600
rect -945 -588 -933 588
rect -899 -588 -887 588
rect -945 -600 -887 -588
rect -487 588 -429 600
rect -487 -588 -475 588
rect -441 -588 -429 588
rect -487 -600 -429 -588
rect -29 588 29 600
rect -29 -588 -17 588
rect 17 -588 29 588
rect -29 -600 29 -588
rect 429 588 487 600
rect 429 -588 441 588
rect 475 -588 487 588
rect 429 -600 487 -588
rect 887 588 945 600
rect 887 -588 899 588
rect 933 -588 945 588
rect 887 -600 945 -588
rect 1345 588 1403 600
rect 1345 -588 1357 588
rect 1391 -588 1403 588
rect 1345 -600 1403 -588
rect 1803 588 1861 600
rect 1803 -588 1815 588
rect 1849 -588 1861 588
rect 1803 -600 1861 -588
rect 2261 588 2319 600
rect 2261 -588 2273 588
rect 2307 -588 2319 588
rect 2261 -600 2319 -588
<< pdiffc >>
rect -2307 -588 -2273 588
rect -1849 -588 -1815 588
rect -1391 -588 -1357 588
rect -933 -588 -899 588
rect -475 -588 -441 588
rect -17 -588 17 588
rect 441 -588 475 588
rect 899 -588 933 588
rect 1357 -588 1391 588
rect 1815 -588 1849 588
rect 2273 -588 2307 588
<< poly >>
rect -2187 681 -1935 697
rect -2187 664 -2171 681
rect -2261 647 -2171 664
rect -1951 664 -1935 681
rect -1729 681 -1477 697
rect -1729 664 -1713 681
rect -1951 647 -1861 664
rect -2261 600 -1861 647
rect -1803 647 -1713 664
rect -1493 664 -1477 681
rect -1271 681 -1019 697
rect -1271 664 -1255 681
rect -1493 647 -1403 664
rect -1803 600 -1403 647
rect -1345 647 -1255 664
rect -1035 664 -1019 681
rect -813 681 -561 697
rect -813 664 -797 681
rect -1035 647 -945 664
rect -1345 600 -945 647
rect -887 647 -797 664
rect -577 664 -561 681
rect -355 681 -103 697
rect -355 664 -339 681
rect -577 647 -487 664
rect -887 600 -487 647
rect -429 647 -339 664
rect -119 664 -103 681
rect 103 681 355 697
rect 103 664 119 681
rect -119 647 -29 664
rect -429 600 -29 647
rect 29 647 119 664
rect 339 664 355 681
rect 561 681 813 697
rect 561 664 577 681
rect 339 647 429 664
rect 29 600 429 647
rect 487 647 577 664
rect 797 664 813 681
rect 1019 681 1271 697
rect 1019 664 1035 681
rect 797 647 887 664
rect 487 600 887 647
rect 945 647 1035 664
rect 1255 664 1271 681
rect 1477 681 1729 697
rect 1477 664 1493 681
rect 1255 647 1345 664
rect 945 600 1345 647
rect 1403 647 1493 664
rect 1713 664 1729 681
rect 1935 681 2187 697
rect 1935 664 1951 681
rect 1713 647 1803 664
rect 1403 600 1803 647
rect 1861 647 1951 664
rect 2171 664 2187 681
rect 2171 647 2261 664
rect 1861 600 2261 647
rect -2261 -647 -1861 -600
rect -2261 -664 -2171 -647
rect -2187 -681 -2171 -664
rect -1951 -664 -1861 -647
rect -1803 -647 -1403 -600
rect -1803 -664 -1713 -647
rect -1951 -681 -1935 -664
rect -2187 -697 -1935 -681
rect -1729 -681 -1713 -664
rect -1493 -664 -1403 -647
rect -1345 -647 -945 -600
rect -1345 -664 -1255 -647
rect -1493 -681 -1477 -664
rect -1729 -697 -1477 -681
rect -1271 -681 -1255 -664
rect -1035 -664 -945 -647
rect -887 -647 -487 -600
rect -887 -664 -797 -647
rect -1035 -681 -1019 -664
rect -1271 -697 -1019 -681
rect -813 -681 -797 -664
rect -577 -664 -487 -647
rect -429 -647 -29 -600
rect -429 -664 -339 -647
rect -577 -681 -561 -664
rect -813 -697 -561 -681
rect -355 -681 -339 -664
rect -119 -664 -29 -647
rect 29 -647 429 -600
rect 29 -664 119 -647
rect -119 -681 -103 -664
rect -355 -697 -103 -681
rect 103 -681 119 -664
rect 339 -664 429 -647
rect 487 -647 887 -600
rect 487 -664 577 -647
rect 339 -681 355 -664
rect 103 -697 355 -681
rect 561 -681 577 -664
rect 797 -664 887 -647
rect 945 -647 1345 -600
rect 945 -664 1035 -647
rect 797 -681 813 -664
rect 561 -697 813 -681
rect 1019 -681 1035 -664
rect 1255 -664 1345 -647
rect 1403 -647 1803 -600
rect 1403 -664 1493 -647
rect 1255 -681 1271 -664
rect 1019 -697 1271 -681
rect 1477 -681 1493 -664
rect 1713 -664 1803 -647
rect 1861 -647 2261 -600
rect 1861 -664 1951 -647
rect 1713 -681 1729 -664
rect 1477 -697 1729 -681
rect 1935 -681 1951 -664
rect 2171 -664 2261 -647
rect 2171 -681 2187 -664
rect 1935 -697 2187 -681
<< polycont >>
rect -2171 647 -1951 681
rect -1713 647 -1493 681
rect -1255 647 -1035 681
rect -797 647 -577 681
rect -339 647 -119 681
rect 119 647 339 681
rect 577 647 797 681
rect 1035 647 1255 681
rect 1493 647 1713 681
rect 1951 647 2171 681
rect -2171 -681 -1951 -647
rect -1713 -681 -1493 -647
rect -1255 -681 -1035 -647
rect -797 -681 -577 -647
rect -339 -681 -119 -647
rect 119 -681 339 -647
rect 577 -681 797 -647
rect 1035 -681 1255 -647
rect 1493 -681 1713 -647
rect 1951 -681 2171 -647
<< locali >>
rect -2187 647 -2171 681
rect -1951 647 -1935 681
rect -1729 647 -1713 681
rect -1493 647 -1477 681
rect -1271 647 -1255 681
rect -1035 647 -1019 681
rect -813 647 -797 681
rect -577 647 -561 681
rect -355 647 -339 681
rect -119 647 -103 681
rect 103 647 119 681
rect 339 647 355 681
rect 561 647 577 681
rect 797 647 813 681
rect 1019 647 1035 681
rect 1255 647 1271 681
rect 1477 647 1493 681
rect 1713 647 1729 681
rect 1935 647 1951 681
rect 2171 647 2187 681
rect -2307 588 -2273 604
rect -2307 -604 -2273 -588
rect -1849 588 -1815 604
rect -1849 -604 -1815 -588
rect -1391 588 -1357 604
rect -1391 -604 -1357 -588
rect -933 588 -899 604
rect -933 -604 -899 -588
rect -475 588 -441 604
rect -475 -604 -441 -588
rect -17 588 17 604
rect -17 -604 17 -588
rect 441 588 475 604
rect 441 -604 475 -588
rect 899 588 933 604
rect 899 -604 933 -588
rect 1357 588 1391 604
rect 1357 -604 1391 -588
rect 1815 588 1849 604
rect 1815 -604 1849 -588
rect 2273 588 2307 604
rect 2273 -604 2307 -588
rect -2187 -681 -2171 -647
rect -1951 -681 -1935 -647
rect -1729 -681 -1713 -647
rect -1493 -681 -1477 -647
rect -1271 -681 -1255 -647
rect -1035 -681 -1019 -647
rect -813 -681 -797 -647
rect -577 -681 -561 -647
rect -355 -681 -339 -647
rect -119 -681 -103 -647
rect 103 -681 119 -647
rect 339 -681 355 -647
rect 561 -681 577 -647
rect 797 -681 813 -647
rect 1019 -681 1035 -647
rect 1255 -681 1271 -647
rect 1477 -681 1493 -647
rect 1713 -681 1729 -647
rect 1935 -681 1951 -647
rect 2171 -681 2187 -647
<< viali >>
rect -2153 647 -1969 681
rect -1695 647 -1511 681
rect -1237 647 -1053 681
rect -779 647 -595 681
rect -321 647 -137 681
rect 137 647 321 681
rect 595 647 779 681
rect 1053 647 1237 681
rect 1511 647 1695 681
rect 1969 647 2153 681
rect -2307 -588 -2273 588
rect -1849 -588 -1815 588
rect -1391 -588 -1357 588
rect -933 -588 -899 588
rect -475 -588 -441 588
rect -17 -588 17 588
rect 441 -588 475 588
rect 899 -588 933 588
rect 1357 -588 1391 588
rect 1815 -588 1849 588
rect 2273 -588 2307 588
rect -2153 -681 -1969 -647
rect -1695 -681 -1511 -647
rect -1237 -681 -1053 -647
rect -779 -681 -595 -647
rect -321 -681 -137 -647
rect 137 -681 321 -647
rect 595 -681 779 -647
rect 1053 -681 1237 -647
rect 1511 -681 1695 -647
rect 1969 -681 2153 -647
<< metal1 >>
rect -2165 681 -1957 687
rect -2165 647 -2153 681
rect -1969 647 -1957 681
rect -2165 641 -1957 647
rect -1707 681 -1499 687
rect -1707 647 -1695 681
rect -1511 647 -1499 681
rect -1707 641 -1499 647
rect -1249 681 -1041 687
rect -1249 647 -1237 681
rect -1053 647 -1041 681
rect -1249 641 -1041 647
rect -791 681 -583 687
rect -791 647 -779 681
rect -595 647 -583 681
rect -791 641 -583 647
rect -333 681 -125 687
rect -333 647 -321 681
rect -137 647 -125 681
rect -333 641 -125 647
rect 125 681 333 687
rect 125 647 137 681
rect 321 647 333 681
rect 125 641 333 647
rect 583 681 791 687
rect 583 647 595 681
rect 779 647 791 681
rect 583 641 791 647
rect 1041 681 1249 687
rect 1041 647 1053 681
rect 1237 647 1249 681
rect 1041 641 1249 647
rect 1499 681 1707 687
rect 1499 647 1511 681
rect 1695 647 1707 681
rect 1499 641 1707 647
rect 1957 681 2165 687
rect 1957 647 1969 681
rect 2153 647 2165 681
rect 1957 641 2165 647
rect -2313 588 -2267 600
rect -2313 -588 -2307 588
rect -2273 -588 -2267 588
rect -2313 -600 -2267 -588
rect -1855 588 -1809 600
rect -1855 -588 -1849 588
rect -1815 -588 -1809 588
rect -1855 -600 -1809 -588
rect -1397 588 -1351 600
rect -1397 -588 -1391 588
rect -1357 -588 -1351 588
rect -1397 -600 -1351 -588
rect -939 588 -893 600
rect -939 -588 -933 588
rect -899 -588 -893 588
rect -939 -600 -893 -588
rect -481 588 -435 600
rect -481 -588 -475 588
rect -441 -588 -435 588
rect -481 -600 -435 -588
rect -23 588 23 600
rect -23 -588 -17 588
rect 17 -588 23 588
rect -23 -600 23 -588
rect 435 588 481 600
rect 435 -588 441 588
rect 475 -588 481 588
rect 435 -600 481 -588
rect 893 588 939 600
rect 893 -588 899 588
rect 933 -588 939 588
rect 893 -600 939 -588
rect 1351 588 1397 600
rect 1351 -588 1357 588
rect 1391 -588 1397 588
rect 1351 -600 1397 -588
rect 1809 588 1855 600
rect 1809 -588 1815 588
rect 1849 -588 1855 588
rect 1809 -600 1855 -588
rect 2267 588 2313 600
rect 2267 -588 2273 588
rect 2307 -588 2313 588
rect 2267 -600 2313 -588
rect -2165 -647 -1957 -641
rect -2165 -681 -2153 -647
rect -1969 -681 -1957 -647
rect -2165 -687 -1957 -681
rect -1707 -647 -1499 -641
rect -1707 -681 -1695 -647
rect -1511 -681 -1499 -647
rect -1707 -687 -1499 -681
rect -1249 -647 -1041 -641
rect -1249 -681 -1237 -647
rect -1053 -681 -1041 -647
rect -1249 -687 -1041 -681
rect -791 -647 -583 -641
rect -791 -681 -779 -647
rect -595 -681 -583 -647
rect -791 -687 -583 -681
rect -333 -647 -125 -641
rect -333 -681 -321 -647
rect -137 -681 -125 -647
rect -333 -687 -125 -681
rect 125 -647 333 -641
rect 125 -681 137 -647
rect 321 -681 333 -647
rect 125 -687 333 -681
rect 583 -647 791 -641
rect 583 -681 595 -647
rect 779 -681 791 -647
rect 583 -687 791 -681
rect 1041 -647 1249 -641
rect 1041 -681 1053 -647
rect 1237 -681 1249 -647
rect 1041 -687 1249 -681
rect 1499 -647 1707 -641
rect 1499 -681 1511 -647
rect 1695 -681 1707 -647
rect 1499 -687 1707 -681
rect 1957 -647 2165 -641
rect 1957 -681 1969 -647
rect 2153 -681 2165 -647
rect 1957 -687 2165 -681
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_hvt
string parameters w 6 l 2 m 1 nf 10 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
