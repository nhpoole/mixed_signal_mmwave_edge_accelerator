magic
tech sky130A
timestamp 1626065694
<< checkpaint >>
rect -505 -521 870 848
<< nwell >>
rect 125 109 240 218
<< nsubdiff >>
rect 160 172 201 185
rect 160 155 172 172
rect 189 155 201 172
rect 160 143 201 155
<< nsubdiffcont >>
rect 172 155 189 172
<< locali >>
rect 158 172 203 187
rect 158 155 172 172
rect 189 155 203 172
rect 158 141 203 155
<< end >>
