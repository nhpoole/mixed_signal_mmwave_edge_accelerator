magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1286 -1286 1436 1358
<< pwell >>
rect -26 -26 176 98
<< scnmos >>
rect 60 0 90 72
<< ndiff >>
rect 0 0 60 72
rect 90 0 150 72
<< poly >>
rect 60 72 90 98
rect 60 -26 90 0
<< locali >>
rect 8 3 42 69
rect 108 3 142 69
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_11  sky130_sram_2kbyte_1rw1r_32x512_8_contact_11_1
timestamp 1626065694
transform 1 0 0 0 1 3
box -26 -22 76 88
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_11  sky130_sram_2kbyte_1rw1r_32x512_8_contact_11_0
timestamp 1626065694
transform 1 0 100 0 1 3
box -26 -22 76 88
<< labels >>
rlabel locali s 25 36 25 36 4 S
rlabel locali s 125 36 125 36 4 D
rlabel poly s 75 36 75 36 4 G
<< properties >>
string FIXED_BBOX -25 -26 175 98
<< end >>
