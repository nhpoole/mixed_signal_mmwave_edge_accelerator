magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< nwell >>
rect 1756 0 3264 490
<< poly >>
rect 77 155 136 185
rect 1588 155 1784 185
<< locali >>
rect 60 137 94 203
rect 829 103 3246 137
<< metal1 >>
rect 848 0 876 395
rect 2496 0 2524 395
use nmos_m1_w7_000_sli_dli_da_p  nmos_m1_w7_000_sli_dli_da_p_0
timestamp 1624494425
transform 0 1 162 -1 0 245
box -26 -26 176 1426
use pmos_m1_w7_000_sli_dli_da_p  pmos_m1_w7_000_sli_dli_da_p_0
timestamp 1624494425
transform 0 1 1810 -1 0 245
box -59 -54 209 1454
use contact_14  contact_14_0
timestamp 1624494425
transform 1 0 837 0 1 354
box -26 -26 76 108
use contact_7  contact_7_0
timestamp 1624494425
transform 1 0 2481 0 1 187
box 0 0 58 66
use contact_7  contact_7_1
timestamp 1624494425
transform 1 0 833 0 1 187
box 0 0 58 66
use contact_15  contact_15_0
timestamp 1624494425
transform 1 0 44 0 1 137
box 0 0 66 66
use contact_7  contact_7_2
timestamp 1624494425
transform 1 0 833 0 1 362
box 0 0 58 66
use contact_7  contact_7_3
timestamp 1624494425
transform 1 0 2481 0 1 362
box 0 0 58 66
use contact_13  contact_13_0
timestamp 1624494425
transform 1 0 2485 0 1 354
box -59 -43 109 125
<< labels >>
rlabel locali s 77 170 77 170 4 A
rlabel locali s 2037 120 2037 120 4 Z
rlabel metal1 s 848 0 876 395 4 gnd
rlabel metal1 s 2496 0 2524 395 4 vdd
<< properties >>
string FIXED_BBOX 0 0 3246 395
<< end >>
