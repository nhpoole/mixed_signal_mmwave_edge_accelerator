magic
tech sky130A
magscale 1 2
timestamp 1620694387
<< nmoslvt >>
rect -5570 -300 -4610 300
rect -4552 -300 -3592 300
rect -3534 -300 -2574 300
rect -2516 -300 -1556 300
rect -1498 -300 -538 300
rect -480 -300 480 300
rect 538 -300 1498 300
rect 1556 -300 2516 300
rect 2574 -300 3534 300
rect 3592 -300 4552 300
rect 4610 -300 5570 300
<< ndiff >>
rect -5628 288 -5570 300
rect -5628 -288 -5616 288
rect -5582 -288 -5570 288
rect -5628 -300 -5570 -288
rect -4610 288 -4552 300
rect -4610 -288 -4598 288
rect -4564 -288 -4552 288
rect -4610 -300 -4552 -288
rect -3592 288 -3534 300
rect -3592 -288 -3580 288
rect -3546 -288 -3534 288
rect -3592 -300 -3534 -288
rect -2574 288 -2516 300
rect -2574 -288 -2562 288
rect -2528 -288 -2516 288
rect -2574 -300 -2516 -288
rect -1556 288 -1498 300
rect -1556 -288 -1544 288
rect -1510 -288 -1498 288
rect -1556 -300 -1498 -288
rect -538 288 -480 300
rect -538 -288 -526 288
rect -492 -288 -480 288
rect -538 -300 -480 -288
rect 480 288 538 300
rect 480 -288 492 288
rect 526 -288 538 288
rect 480 -300 538 -288
rect 1498 288 1556 300
rect 1498 -288 1510 288
rect 1544 -288 1556 288
rect 1498 -300 1556 -288
rect 2516 288 2574 300
rect 2516 -288 2528 288
rect 2562 -288 2574 288
rect 2516 -300 2574 -288
rect 3534 288 3592 300
rect 3534 -288 3546 288
rect 3580 -288 3592 288
rect 3534 -300 3592 -288
rect 4552 288 4610 300
rect 4552 -288 4564 288
rect 4598 -288 4610 288
rect 4552 -300 4610 -288
rect 5570 288 5628 300
rect 5570 -288 5582 288
rect 5616 -288 5628 288
rect 5570 -300 5628 -288
<< ndiffc >>
rect -5616 -288 -5582 288
rect -4598 -288 -4564 288
rect -3580 -288 -3546 288
rect -2562 -288 -2528 288
rect -1544 -288 -1510 288
rect -526 -288 -492 288
rect 492 -288 526 288
rect 1510 -288 1544 288
rect 2528 -288 2562 288
rect 3546 -288 3580 288
rect 4564 -288 4598 288
rect 5582 -288 5616 288
<< poly >>
rect -5384 372 -4796 388
rect -5384 355 -5368 372
rect -5570 338 -5368 355
rect -4812 355 -4796 372
rect -4366 372 -3778 388
rect -4366 355 -4350 372
rect -4812 338 -4610 355
rect -5570 300 -4610 338
rect -4552 338 -4350 355
rect -3794 355 -3778 372
rect -3348 372 -2760 388
rect -3348 355 -3332 372
rect -3794 338 -3592 355
rect -4552 300 -3592 338
rect -3534 338 -3332 355
rect -2776 355 -2760 372
rect -2330 372 -1742 388
rect -2330 355 -2314 372
rect -2776 338 -2574 355
rect -3534 300 -2574 338
rect -2516 338 -2314 355
rect -1758 355 -1742 372
rect -1312 372 -724 388
rect -1312 355 -1296 372
rect -1758 338 -1556 355
rect -2516 300 -1556 338
rect -1498 338 -1296 355
rect -740 355 -724 372
rect -294 372 294 388
rect -294 355 -278 372
rect -740 338 -538 355
rect -1498 300 -538 338
rect -480 338 -278 355
rect 278 355 294 372
rect 724 372 1312 388
rect 724 355 740 372
rect 278 338 480 355
rect -480 300 480 338
rect 538 338 740 355
rect 1296 355 1312 372
rect 1742 372 2330 388
rect 1742 355 1758 372
rect 1296 338 1498 355
rect 538 300 1498 338
rect 1556 338 1758 355
rect 2314 355 2330 372
rect 2760 372 3348 388
rect 2760 355 2776 372
rect 2314 338 2516 355
rect 1556 300 2516 338
rect 2574 338 2776 355
rect 3332 355 3348 372
rect 3778 372 4366 388
rect 3778 355 3794 372
rect 3332 338 3534 355
rect 2574 300 3534 338
rect 3592 338 3794 355
rect 4350 355 4366 372
rect 4796 372 5384 388
rect 4796 355 4812 372
rect 4350 338 4552 355
rect 3592 300 4552 338
rect 4610 338 4812 355
rect 5368 355 5384 372
rect 5368 338 5570 355
rect 4610 300 5570 338
rect -5570 -338 -4610 -300
rect -5570 -355 -5368 -338
rect -5384 -372 -5368 -355
rect -4812 -355 -4610 -338
rect -4552 -338 -3592 -300
rect -4552 -355 -4350 -338
rect -4812 -372 -4796 -355
rect -5384 -388 -4796 -372
rect -4366 -372 -4350 -355
rect -3794 -355 -3592 -338
rect -3534 -338 -2574 -300
rect -3534 -355 -3332 -338
rect -3794 -372 -3778 -355
rect -4366 -388 -3778 -372
rect -3348 -372 -3332 -355
rect -2776 -355 -2574 -338
rect -2516 -338 -1556 -300
rect -2516 -355 -2314 -338
rect -2776 -372 -2760 -355
rect -3348 -388 -2760 -372
rect -2330 -372 -2314 -355
rect -1758 -355 -1556 -338
rect -1498 -338 -538 -300
rect -1498 -355 -1296 -338
rect -1758 -372 -1742 -355
rect -2330 -388 -1742 -372
rect -1312 -372 -1296 -355
rect -740 -355 -538 -338
rect -480 -338 480 -300
rect -480 -355 -278 -338
rect -740 -372 -724 -355
rect -1312 -388 -724 -372
rect -294 -372 -278 -355
rect 278 -355 480 -338
rect 538 -338 1498 -300
rect 538 -355 740 -338
rect 278 -372 294 -355
rect -294 -388 294 -372
rect 724 -372 740 -355
rect 1296 -355 1498 -338
rect 1556 -338 2516 -300
rect 1556 -355 1758 -338
rect 1296 -372 1312 -355
rect 724 -388 1312 -372
rect 1742 -372 1758 -355
rect 2314 -355 2516 -338
rect 2574 -338 3534 -300
rect 2574 -355 2776 -338
rect 2314 -372 2330 -355
rect 1742 -388 2330 -372
rect 2760 -372 2776 -355
rect 3332 -355 3534 -338
rect 3592 -338 4552 -300
rect 3592 -355 3794 -338
rect 3332 -372 3348 -355
rect 2760 -388 3348 -372
rect 3778 -372 3794 -355
rect 4350 -355 4552 -338
rect 4610 -338 5570 -300
rect 4610 -355 4812 -338
rect 4350 -372 4366 -355
rect 3778 -388 4366 -372
rect 4796 -372 4812 -355
rect 5368 -355 5570 -338
rect 5368 -372 5384 -355
rect 4796 -388 5384 -372
<< polycont >>
rect -5368 338 -4812 372
rect -4350 338 -3794 372
rect -3332 338 -2776 372
rect -2314 338 -1758 372
rect -1296 338 -740 372
rect -278 338 278 372
rect 740 338 1296 372
rect 1758 338 2314 372
rect 2776 338 3332 372
rect 3794 338 4350 372
rect 4812 338 5368 372
rect -5368 -372 -4812 -338
rect -4350 -372 -3794 -338
rect -3332 -372 -2776 -338
rect -2314 -372 -1758 -338
rect -1296 -372 -740 -338
rect -278 -372 278 -338
rect 740 -372 1296 -338
rect 1758 -372 2314 -338
rect 2776 -372 3332 -338
rect 3794 -372 4350 -338
rect 4812 -372 5368 -338
<< locali >>
rect -5384 338 -5368 372
rect -4812 338 -4796 372
rect -4366 338 -4350 372
rect -3794 338 -3778 372
rect -3348 338 -3332 372
rect -2776 338 -2760 372
rect -2330 338 -2314 372
rect -1758 338 -1742 372
rect -1312 338 -1296 372
rect -740 338 -724 372
rect -294 338 -278 372
rect 278 338 294 372
rect 724 338 740 372
rect 1296 338 1312 372
rect 1742 338 1758 372
rect 2314 338 2330 372
rect 2760 338 2776 372
rect 3332 338 3348 372
rect 3778 338 3794 372
rect 4350 338 4366 372
rect 4796 338 4812 372
rect 5368 338 5384 372
rect -5616 288 -5582 304
rect -5616 -304 -5582 -288
rect -4598 288 -4564 304
rect -4598 -304 -4564 -288
rect -3580 288 -3546 304
rect -3580 -304 -3546 -288
rect -2562 288 -2528 304
rect -2562 -304 -2528 -288
rect -1544 288 -1510 304
rect -1544 -304 -1510 -288
rect -526 288 -492 304
rect -526 -304 -492 -288
rect 492 288 526 304
rect 492 -304 526 -288
rect 1510 288 1544 304
rect 1510 -304 1544 -288
rect 2528 288 2562 304
rect 2528 -304 2562 -288
rect 3546 288 3580 304
rect 3546 -304 3580 -288
rect 4564 288 4598 304
rect 4564 -304 4598 -288
rect 5582 288 5616 304
rect 5582 -304 5616 -288
rect -5384 -372 -5368 -338
rect -4812 -372 -4796 -338
rect -4366 -372 -4350 -338
rect -3794 -372 -3778 -338
rect -3348 -372 -3332 -338
rect -2776 -372 -2760 -338
rect -2330 -372 -2314 -338
rect -1758 -372 -1742 -338
rect -1312 -372 -1296 -338
rect -740 -372 -724 -338
rect -294 -372 -278 -338
rect 278 -372 294 -338
rect 724 -372 740 -338
rect 1296 -372 1312 -338
rect 1742 -372 1758 -338
rect 2314 -372 2330 -338
rect 2760 -372 2776 -338
rect 3332 -372 3348 -338
rect 3778 -372 3794 -338
rect 4350 -372 4366 -338
rect 4796 -372 4812 -338
rect 5368 -372 5384 -338
<< viali >>
rect -5322 338 -4858 372
rect -4304 338 -3840 372
rect -3286 338 -2822 372
rect -2268 338 -1804 372
rect -1250 338 -786 372
rect -232 338 232 372
rect 786 338 1250 372
rect 1804 338 2268 372
rect 2822 338 3286 372
rect 3840 338 4304 372
rect 4858 338 5322 372
rect -5616 -288 -5582 288
rect -4598 -288 -4564 288
rect -3580 -288 -3546 288
rect -2562 -288 -2528 288
rect -1544 -288 -1510 288
rect -526 -288 -492 288
rect 492 -288 526 288
rect 1510 -288 1544 288
rect 2528 -288 2562 288
rect 3546 -288 3580 288
rect 4564 -288 4598 288
rect 5582 -288 5616 288
rect -5322 -372 -4858 -338
rect -4304 -372 -3840 -338
rect -3286 -372 -2822 -338
rect -2268 -372 -1804 -338
rect -1250 -372 -786 -338
rect -232 -372 232 -338
rect 786 -372 1250 -338
rect 1804 -372 2268 -338
rect 2822 -372 3286 -338
rect 3840 -372 4304 -338
rect 4858 -372 5322 -338
<< metal1 >>
rect -5334 372 -4846 378
rect -5334 338 -5322 372
rect -4858 338 -4846 372
rect -5334 332 -4846 338
rect -4316 372 -3828 378
rect -4316 338 -4304 372
rect -3840 338 -3828 372
rect -4316 332 -3828 338
rect -3298 372 -2810 378
rect -3298 338 -3286 372
rect -2822 338 -2810 372
rect -3298 332 -2810 338
rect -2280 372 -1792 378
rect -2280 338 -2268 372
rect -1804 338 -1792 372
rect -2280 332 -1792 338
rect -1262 372 -774 378
rect -1262 338 -1250 372
rect -786 338 -774 372
rect -1262 332 -774 338
rect -244 372 244 378
rect -244 338 -232 372
rect 232 338 244 372
rect -244 332 244 338
rect 774 372 1262 378
rect 774 338 786 372
rect 1250 338 1262 372
rect 774 332 1262 338
rect 1792 372 2280 378
rect 1792 338 1804 372
rect 2268 338 2280 372
rect 1792 332 2280 338
rect 2810 372 3298 378
rect 2810 338 2822 372
rect 3286 338 3298 372
rect 2810 332 3298 338
rect 3828 372 4316 378
rect 3828 338 3840 372
rect 4304 338 4316 372
rect 3828 332 4316 338
rect 4846 372 5334 378
rect 4846 338 4858 372
rect 5322 338 5334 372
rect 4846 332 5334 338
rect -5622 288 -5576 300
rect -5622 -288 -5616 288
rect -5582 -288 -5576 288
rect -5622 -300 -5576 -288
rect -4604 288 -4558 300
rect -4604 -288 -4598 288
rect -4564 -288 -4558 288
rect -4604 -300 -4558 -288
rect -3586 288 -3540 300
rect -3586 -288 -3580 288
rect -3546 -288 -3540 288
rect -3586 -300 -3540 -288
rect -2568 288 -2522 300
rect -2568 -288 -2562 288
rect -2528 -288 -2522 288
rect -2568 -300 -2522 -288
rect -1550 288 -1504 300
rect -1550 -288 -1544 288
rect -1510 -288 -1504 288
rect -1550 -300 -1504 -288
rect -532 288 -486 300
rect -532 -288 -526 288
rect -492 -288 -486 288
rect -532 -300 -486 -288
rect 486 288 532 300
rect 486 -288 492 288
rect 526 -288 532 288
rect 486 -300 532 -288
rect 1504 288 1550 300
rect 1504 -288 1510 288
rect 1544 -288 1550 288
rect 1504 -300 1550 -288
rect 2522 288 2568 300
rect 2522 -288 2528 288
rect 2562 -288 2568 288
rect 2522 -300 2568 -288
rect 3540 288 3586 300
rect 3540 -288 3546 288
rect 3580 -288 3586 288
rect 3540 -300 3586 -288
rect 4558 288 4604 300
rect 4558 -288 4564 288
rect 4598 -288 4604 288
rect 4558 -300 4604 -288
rect 5576 288 5622 300
rect 5576 -288 5582 288
rect 5616 -288 5622 288
rect 5576 -300 5622 -288
rect -5334 -338 -4846 -332
rect -5334 -372 -5322 -338
rect -4858 -372 -4846 -338
rect -5334 -378 -4846 -372
rect -4316 -338 -3828 -332
rect -4316 -372 -4304 -338
rect -3840 -372 -3828 -338
rect -4316 -378 -3828 -372
rect -3298 -338 -2810 -332
rect -3298 -372 -3286 -338
rect -2822 -372 -2810 -338
rect -3298 -378 -2810 -372
rect -2280 -338 -1792 -332
rect -2280 -372 -2268 -338
rect -1804 -372 -1792 -338
rect -2280 -378 -1792 -372
rect -1262 -338 -774 -332
rect -1262 -372 -1250 -338
rect -786 -372 -774 -338
rect -1262 -378 -774 -372
rect -244 -338 244 -332
rect -244 -372 -232 -338
rect 232 -372 244 -338
rect -244 -378 244 -372
rect 774 -338 1262 -332
rect 774 -372 786 -338
rect 1250 -372 1262 -338
rect 774 -378 1262 -372
rect 1792 -338 2280 -332
rect 1792 -372 1804 -338
rect 2268 -372 2280 -338
rect 1792 -378 2280 -372
rect 2810 -338 3298 -332
rect 2810 -372 2822 -338
rect 3286 -372 3298 -338
rect 2810 -378 3298 -372
rect 3828 -338 4316 -332
rect 3828 -372 3840 -338
rect 4304 -372 4316 -338
rect 3828 -378 4316 -372
rect 4846 -338 5334 -332
rect 4846 -372 4858 -338
rect 5322 -372 5334 -338
rect 4846 -378 5334 -372
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string parameters w 3 l 4.8 m 1 nf 11 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
