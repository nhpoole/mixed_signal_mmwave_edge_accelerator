magic
tech sky130A
timestamp 1626065694
<< checkpaint >>
rect -701 -701 701 701
<< via4 >>
rect -59 -59 59 59
<< metal5 >>
rect -71 59 71 71
rect -71 -59 -59 59
rect 59 -59 71 59
rect -71 -71 71 -59
<< end >>
