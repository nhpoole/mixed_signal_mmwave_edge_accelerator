magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -17828 -2138 78210 32088
<< nwell >>
rect 36584 12390 38738 14006
<< nsubdiff >>
rect 36718 13937 38682 13970
rect 36718 13903 36901 13937
rect 36935 13903 36969 13937
rect 37003 13903 37037 13937
rect 37071 13903 37105 13937
rect 37139 13903 37173 13937
rect 37207 13903 37241 13937
rect 37275 13903 37309 13937
rect 37343 13903 37377 13937
rect 37411 13903 37445 13937
rect 37479 13903 37513 13937
rect 37547 13903 37581 13937
rect 37615 13903 37649 13937
rect 37683 13903 37717 13937
rect 37751 13903 37785 13937
rect 37819 13903 37853 13937
rect 37887 13903 37921 13937
rect 37955 13903 37989 13937
rect 38023 13903 38057 13937
rect 38091 13903 38125 13937
rect 38159 13903 38193 13937
rect 38227 13903 38261 13937
rect 38295 13903 38329 13937
rect 38363 13903 38397 13937
rect 38431 13903 38465 13937
rect 38499 13903 38682 13937
rect 36718 13870 38682 13903
rect 36718 13793 36818 13870
rect 36718 13759 36751 13793
rect 36785 13759 36818 13793
rect 36718 13725 36818 13759
rect 36718 13691 36751 13725
rect 36785 13691 36818 13725
rect 36718 13657 36818 13691
rect 36718 13623 36751 13657
rect 36785 13623 36818 13657
rect 36718 13589 36818 13623
rect 36718 13555 36751 13589
rect 36785 13555 36818 13589
rect 36718 13521 36818 13555
rect 36718 13487 36751 13521
rect 36785 13487 36818 13521
rect 36718 13453 36818 13487
rect 36718 13419 36751 13453
rect 36785 13419 36818 13453
rect 36718 13385 36818 13419
rect 36718 13351 36751 13385
rect 36785 13351 36818 13385
rect 36718 13317 36818 13351
rect 36718 13283 36751 13317
rect 36785 13283 36818 13317
rect 36718 13249 36818 13283
rect 36718 13215 36751 13249
rect 36785 13215 36818 13249
rect 36718 13181 36818 13215
rect 36718 13147 36751 13181
rect 36785 13147 36818 13181
rect 36718 13113 36818 13147
rect 36718 13079 36751 13113
rect 36785 13079 36818 13113
rect 36718 13045 36818 13079
rect 36718 13011 36751 13045
rect 36785 13011 36818 13045
rect 36718 12977 36818 13011
rect 36718 12943 36751 12977
rect 36785 12943 36818 12977
rect 36718 12909 36818 12943
rect 36718 12875 36751 12909
rect 36785 12875 36818 12909
rect 36718 12841 36818 12875
rect 36718 12807 36751 12841
rect 36785 12807 36818 12841
rect 36718 12773 36818 12807
rect 36718 12739 36751 12773
rect 36785 12739 36818 12773
rect 36718 12705 36818 12739
rect 36718 12671 36751 12705
rect 36785 12671 36818 12705
rect 36718 12637 36818 12671
rect 36718 12603 36751 12637
rect 36785 12603 36818 12637
rect 36718 12526 36818 12603
rect 38582 13793 38682 13870
rect 38582 13759 38615 13793
rect 38649 13759 38682 13793
rect 38582 13725 38682 13759
rect 38582 13691 38615 13725
rect 38649 13691 38682 13725
rect 38582 13657 38682 13691
rect 38582 13623 38615 13657
rect 38649 13623 38682 13657
rect 38582 13589 38682 13623
rect 38582 13555 38615 13589
rect 38649 13555 38682 13589
rect 38582 13521 38682 13555
rect 38582 13487 38615 13521
rect 38649 13487 38682 13521
rect 38582 13453 38682 13487
rect 38582 13419 38615 13453
rect 38649 13419 38682 13453
rect 38582 13385 38682 13419
rect 38582 13351 38615 13385
rect 38649 13351 38682 13385
rect 38582 13317 38682 13351
rect 38582 13283 38615 13317
rect 38649 13283 38682 13317
rect 38582 13249 38682 13283
rect 38582 13215 38615 13249
rect 38649 13215 38682 13249
rect 38582 13181 38682 13215
rect 38582 13147 38615 13181
rect 38649 13147 38682 13181
rect 38582 13113 38682 13147
rect 38582 13079 38615 13113
rect 38649 13079 38682 13113
rect 38582 13045 38682 13079
rect 38582 13011 38615 13045
rect 38649 13011 38682 13045
rect 38582 12977 38682 13011
rect 38582 12943 38615 12977
rect 38649 12943 38682 12977
rect 38582 12909 38682 12943
rect 38582 12875 38615 12909
rect 38649 12875 38682 12909
rect 38582 12841 38682 12875
rect 38582 12807 38615 12841
rect 38649 12807 38682 12841
rect 38582 12773 38682 12807
rect 38582 12739 38615 12773
rect 38649 12739 38682 12773
rect 38582 12705 38682 12739
rect 38582 12671 38615 12705
rect 38649 12671 38682 12705
rect 38582 12637 38682 12671
rect 38582 12603 38615 12637
rect 38649 12603 38682 12637
rect 38582 12526 38682 12603
rect 36718 12493 38682 12526
rect 36718 12459 36901 12493
rect 36935 12459 36969 12493
rect 37003 12459 37037 12493
rect 37071 12459 37105 12493
rect 37139 12459 37173 12493
rect 37207 12459 37241 12493
rect 37275 12459 37309 12493
rect 37343 12459 37377 12493
rect 37411 12459 37445 12493
rect 37479 12459 37513 12493
rect 37547 12459 37581 12493
rect 37615 12459 37649 12493
rect 37683 12459 37717 12493
rect 37751 12459 37785 12493
rect 37819 12459 37853 12493
rect 37887 12459 37921 12493
rect 37955 12459 37989 12493
rect 38023 12459 38057 12493
rect 38091 12459 38125 12493
rect 38159 12459 38193 12493
rect 38227 12459 38261 12493
rect 38295 12459 38329 12493
rect 38363 12459 38397 12493
rect 38431 12459 38465 12493
rect 38499 12459 38682 12493
rect 36718 12426 38682 12459
<< nsubdiffcont >>
rect 36901 13903 36935 13937
rect 36969 13903 37003 13937
rect 37037 13903 37071 13937
rect 37105 13903 37139 13937
rect 37173 13903 37207 13937
rect 37241 13903 37275 13937
rect 37309 13903 37343 13937
rect 37377 13903 37411 13937
rect 37445 13903 37479 13937
rect 37513 13903 37547 13937
rect 37581 13903 37615 13937
rect 37649 13903 37683 13937
rect 37717 13903 37751 13937
rect 37785 13903 37819 13937
rect 37853 13903 37887 13937
rect 37921 13903 37955 13937
rect 37989 13903 38023 13937
rect 38057 13903 38091 13937
rect 38125 13903 38159 13937
rect 38193 13903 38227 13937
rect 38261 13903 38295 13937
rect 38329 13903 38363 13937
rect 38397 13903 38431 13937
rect 38465 13903 38499 13937
rect 36751 13759 36785 13793
rect 36751 13691 36785 13725
rect 36751 13623 36785 13657
rect 36751 13555 36785 13589
rect 36751 13487 36785 13521
rect 36751 13419 36785 13453
rect 36751 13351 36785 13385
rect 36751 13283 36785 13317
rect 36751 13215 36785 13249
rect 36751 13147 36785 13181
rect 36751 13079 36785 13113
rect 36751 13011 36785 13045
rect 36751 12943 36785 12977
rect 36751 12875 36785 12909
rect 36751 12807 36785 12841
rect 36751 12739 36785 12773
rect 36751 12671 36785 12705
rect 36751 12603 36785 12637
rect 38615 13759 38649 13793
rect 38615 13691 38649 13725
rect 38615 13623 38649 13657
rect 38615 13555 38649 13589
rect 38615 13487 38649 13521
rect 38615 13419 38649 13453
rect 38615 13351 38649 13385
rect 38615 13283 38649 13317
rect 38615 13215 38649 13249
rect 38615 13147 38649 13181
rect 38615 13079 38649 13113
rect 38615 13011 38649 13045
rect 38615 12943 38649 12977
rect 38615 12875 38649 12909
rect 38615 12807 38649 12841
rect 38615 12739 38649 12773
rect 38615 12671 38649 12705
rect 38615 12603 38649 12637
rect 36901 12459 36935 12493
rect 36969 12459 37003 12493
rect 37037 12459 37071 12493
rect 37105 12459 37139 12493
rect 37173 12459 37207 12493
rect 37241 12459 37275 12493
rect 37309 12459 37343 12493
rect 37377 12459 37411 12493
rect 37445 12459 37479 12493
rect 37513 12459 37547 12493
rect 37581 12459 37615 12493
rect 37649 12459 37683 12493
rect 37717 12459 37751 12493
rect 37785 12459 37819 12493
rect 37853 12459 37887 12493
rect 37921 12459 37955 12493
rect 37989 12459 38023 12493
rect 38057 12459 38091 12493
rect 38125 12459 38159 12493
rect 38193 12459 38227 12493
rect 38261 12459 38295 12493
rect 38329 12459 38363 12493
rect 38397 12459 38431 12493
rect 38465 12459 38499 12493
<< locali >>
rect 36718 13937 38682 13970
rect 36718 13903 36819 13937
rect 36853 13903 36891 13937
rect 36935 13903 36963 13937
rect 37003 13903 37035 13937
rect 37071 13903 37105 13937
rect 37141 13903 37173 13937
rect 37213 13903 37241 13937
rect 37285 13903 37309 13937
rect 37357 13903 37377 13937
rect 37429 13903 37445 13937
rect 37501 13903 37513 13937
rect 37573 13903 37581 13937
rect 37645 13903 37649 13937
rect 37751 13903 37755 13937
rect 37819 13903 37827 13937
rect 37887 13903 37899 13937
rect 37955 13903 37971 13937
rect 38023 13903 38043 13937
rect 38091 13903 38115 13937
rect 38159 13903 38187 13937
rect 38227 13903 38259 13937
rect 38295 13903 38329 13937
rect 38365 13903 38397 13937
rect 38437 13903 38465 13937
rect 38509 13903 38547 13937
rect 38581 13903 38682 13937
rect 36718 13870 38682 13903
rect 36718 13793 36818 13870
rect 36718 13757 36751 13793
rect 36785 13757 36818 13793
rect 36718 13725 36818 13757
rect 36718 13685 36751 13725
rect 36785 13685 36818 13725
rect 36718 13657 36818 13685
rect 36718 13613 36751 13657
rect 36785 13613 36818 13657
rect 36718 13589 36818 13613
rect 36718 13541 36751 13589
rect 36785 13541 36818 13589
rect 36718 13521 36818 13541
rect 36718 13469 36751 13521
rect 36785 13469 36818 13521
rect 36718 13453 36818 13469
rect 36718 13397 36751 13453
rect 36785 13397 36818 13453
rect 36718 13385 36818 13397
rect 36718 13325 36751 13385
rect 36785 13325 36818 13385
rect 36718 13317 36818 13325
rect 36718 13253 36751 13317
rect 36785 13253 36818 13317
rect 36718 13249 36818 13253
rect 36718 13147 36751 13249
rect 36785 13147 36818 13249
rect 36718 13143 36818 13147
rect 36718 13079 36751 13143
rect 36785 13079 36818 13143
rect 36718 13071 36818 13079
rect 36718 13011 36751 13071
rect 36785 13011 36818 13071
rect 36718 12999 36818 13011
rect 36718 12943 36751 12999
rect 36785 12943 36818 12999
rect 36718 12927 36818 12943
rect 36718 12875 36751 12927
rect 36785 12875 36818 12927
rect 36718 12855 36818 12875
rect 36718 12807 36751 12855
rect 36785 12807 36818 12855
rect 36718 12783 36818 12807
rect 36718 12739 36751 12783
rect 36785 12739 36818 12783
rect 36718 12711 36818 12739
rect 36718 12671 36751 12711
rect 36785 12671 36818 12711
rect 36718 12639 36818 12671
rect 36718 12603 36751 12639
rect 36785 12603 36818 12639
rect 36718 12526 36818 12603
rect 38582 13793 38682 13870
rect 38582 13757 38615 13793
rect 38649 13757 38682 13793
rect 38582 13725 38682 13757
rect 38582 13685 38615 13725
rect 38649 13685 38682 13725
rect 38582 13657 38682 13685
rect 38582 13613 38615 13657
rect 38649 13613 38682 13657
rect 38582 13589 38682 13613
rect 38582 13541 38615 13589
rect 38649 13541 38682 13589
rect 38582 13521 38682 13541
rect 38582 13469 38615 13521
rect 38649 13469 38682 13521
rect 38582 13453 38682 13469
rect 38582 13397 38615 13453
rect 38649 13397 38682 13453
rect 38582 13385 38682 13397
rect 38582 13325 38615 13385
rect 38649 13325 38682 13385
rect 38582 13317 38682 13325
rect 38582 13253 38615 13317
rect 38649 13253 38682 13317
rect 38582 13249 38682 13253
rect 38582 13147 38615 13249
rect 38649 13147 38682 13249
rect 38582 13143 38682 13147
rect 38582 13079 38615 13143
rect 38649 13079 38682 13143
rect 38582 13071 38682 13079
rect 38582 13011 38615 13071
rect 38649 13011 38682 13071
rect 38582 12999 38682 13011
rect 38582 12943 38615 12999
rect 38649 12943 38682 12999
rect 38582 12927 38682 12943
rect 38582 12875 38615 12927
rect 38649 12875 38682 12927
rect 38582 12855 38682 12875
rect 38582 12807 38615 12855
rect 38649 12807 38682 12855
rect 38582 12783 38682 12807
rect 38582 12739 38615 12783
rect 38649 12739 38682 12783
rect 38582 12711 38682 12739
rect 38582 12671 38615 12711
rect 38649 12671 38682 12711
rect 38582 12639 38682 12671
rect 38582 12603 38615 12639
rect 38649 12603 38682 12639
rect 38582 12526 38682 12603
rect 36718 12493 38682 12526
rect 36718 12459 36819 12493
rect 36853 12459 36891 12493
rect 36935 12459 36963 12493
rect 37003 12459 37035 12493
rect 37071 12459 37105 12493
rect 37141 12459 37173 12493
rect 37213 12459 37241 12493
rect 37285 12459 37309 12493
rect 37357 12459 37377 12493
rect 37429 12459 37445 12493
rect 37501 12459 37513 12493
rect 37573 12459 37581 12493
rect 37645 12459 37649 12493
rect 37751 12459 37755 12493
rect 37819 12459 37827 12493
rect 37887 12459 37899 12493
rect 37955 12459 37971 12493
rect 38023 12459 38043 12493
rect 38091 12459 38115 12493
rect 38159 12459 38187 12493
rect 38227 12459 38259 12493
rect 38295 12459 38329 12493
rect 38365 12459 38397 12493
rect 38437 12459 38465 12493
rect 38509 12459 38547 12493
rect 38581 12459 38682 12493
rect 36718 12426 38682 12459
rect -1114 362 -1103 396
rect -1069 362 -1031 396
rect -997 362 -959 396
rect -925 362 -914 396
rect -1188 327 -1154 360
rect -1188 255 -1154 293
rect -1188 183 -1154 221
rect -1188 111 -1154 149
rect -1188 39 -1154 77
rect -1188 -33 -1154 5
rect -1188 -100 -1154 -67
rect -872 328 -836 358
rect -872 294 -871 328
rect -837 294 -836 328
rect -872 256 -836 294
rect -872 222 -871 256
rect -837 222 -836 256
rect -872 184 -836 222
rect -872 150 -871 184
rect -837 150 -836 184
rect -872 112 -836 150
rect -872 78 -871 112
rect -837 78 -836 112
rect -872 40 -836 78
rect -872 6 -871 40
rect -837 6 -836 40
rect -872 -32 -836 6
rect -872 -66 -871 -32
rect -837 -66 -836 -32
rect -872 -96 -836 -66
rect -1116 -136 -1105 -102
rect -1071 -136 -1033 -102
rect -999 -136 -961 -102
rect -927 -136 -916 -102
<< viali >>
rect 36819 13903 36853 13937
rect 36891 13903 36901 13937
rect 36901 13903 36925 13937
rect 36963 13903 36969 13937
rect 36969 13903 36997 13937
rect 37035 13903 37037 13937
rect 37037 13903 37069 13937
rect 37107 13903 37139 13937
rect 37139 13903 37141 13937
rect 37179 13903 37207 13937
rect 37207 13903 37213 13937
rect 37251 13903 37275 13937
rect 37275 13903 37285 13937
rect 37323 13903 37343 13937
rect 37343 13903 37357 13937
rect 37395 13903 37411 13937
rect 37411 13903 37429 13937
rect 37467 13903 37479 13937
rect 37479 13903 37501 13937
rect 37539 13903 37547 13937
rect 37547 13903 37573 13937
rect 37611 13903 37615 13937
rect 37615 13903 37645 13937
rect 37683 13903 37717 13937
rect 37755 13903 37785 13937
rect 37785 13903 37789 13937
rect 37827 13903 37853 13937
rect 37853 13903 37861 13937
rect 37899 13903 37921 13937
rect 37921 13903 37933 13937
rect 37971 13903 37989 13937
rect 37989 13903 38005 13937
rect 38043 13903 38057 13937
rect 38057 13903 38077 13937
rect 38115 13903 38125 13937
rect 38125 13903 38149 13937
rect 38187 13903 38193 13937
rect 38193 13903 38221 13937
rect 38259 13903 38261 13937
rect 38261 13903 38293 13937
rect 38331 13903 38363 13937
rect 38363 13903 38365 13937
rect 38403 13903 38431 13937
rect 38431 13903 38437 13937
rect 38475 13903 38499 13937
rect 38499 13903 38509 13937
rect 38547 13903 38581 13937
rect 36751 13759 36785 13791
rect 36751 13757 36785 13759
rect 36751 13691 36785 13719
rect 36751 13685 36785 13691
rect 36751 13623 36785 13647
rect 36751 13613 36785 13623
rect 36751 13555 36785 13575
rect 36751 13541 36785 13555
rect 36751 13487 36785 13503
rect 36751 13469 36785 13487
rect 36751 13419 36785 13431
rect 36751 13397 36785 13419
rect 36751 13351 36785 13359
rect 36751 13325 36785 13351
rect 36751 13283 36785 13287
rect 36751 13253 36785 13283
rect 36751 13181 36785 13215
rect 36751 13113 36785 13143
rect 36751 13109 36785 13113
rect 36751 13045 36785 13071
rect 36751 13037 36785 13045
rect 36751 12977 36785 12999
rect 36751 12965 36785 12977
rect 36751 12909 36785 12927
rect 36751 12893 36785 12909
rect 36751 12841 36785 12855
rect 36751 12821 36785 12841
rect 36751 12773 36785 12783
rect 36751 12749 36785 12773
rect 36751 12705 36785 12711
rect 36751 12677 36785 12705
rect 36751 12637 36785 12639
rect 36751 12605 36785 12637
rect 38615 13759 38649 13791
rect 38615 13757 38649 13759
rect 38615 13691 38649 13719
rect 38615 13685 38649 13691
rect 38615 13623 38649 13647
rect 38615 13613 38649 13623
rect 38615 13555 38649 13575
rect 38615 13541 38649 13555
rect 38615 13487 38649 13503
rect 38615 13469 38649 13487
rect 38615 13419 38649 13431
rect 38615 13397 38649 13419
rect 38615 13351 38649 13359
rect 38615 13325 38649 13351
rect 38615 13283 38649 13287
rect 38615 13253 38649 13283
rect 38615 13181 38649 13215
rect 38615 13113 38649 13143
rect 38615 13109 38649 13113
rect 38615 13045 38649 13071
rect 38615 13037 38649 13045
rect 38615 12977 38649 12999
rect 38615 12965 38649 12977
rect 38615 12909 38649 12927
rect 38615 12893 38649 12909
rect 38615 12841 38649 12855
rect 38615 12821 38649 12841
rect 38615 12773 38649 12783
rect 38615 12749 38649 12773
rect 38615 12705 38649 12711
rect 38615 12677 38649 12705
rect 38615 12637 38649 12639
rect 38615 12605 38649 12637
rect 36819 12459 36853 12493
rect 36891 12459 36901 12493
rect 36901 12459 36925 12493
rect 36963 12459 36969 12493
rect 36969 12459 36997 12493
rect 37035 12459 37037 12493
rect 37037 12459 37069 12493
rect 37107 12459 37139 12493
rect 37139 12459 37141 12493
rect 37179 12459 37207 12493
rect 37207 12459 37213 12493
rect 37251 12459 37275 12493
rect 37275 12459 37285 12493
rect 37323 12459 37343 12493
rect 37343 12459 37357 12493
rect 37395 12459 37411 12493
rect 37411 12459 37429 12493
rect 37467 12459 37479 12493
rect 37479 12459 37501 12493
rect 37539 12459 37547 12493
rect 37547 12459 37573 12493
rect 37611 12459 37615 12493
rect 37615 12459 37645 12493
rect 37683 12459 37717 12493
rect 37755 12459 37785 12493
rect 37785 12459 37789 12493
rect 37827 12459 37853 12493
rect 37853 12459 37861 12493
rect 37899 12459 37921 12493
rect 37921 12459 37933 12493
rect 37971 12459 37989 12493
rect 37989 12459 38005 12493
rect 38043 12459 38057 12493
rect 38057 12459 38077 12493
rect 38115 12459 38125 12493
rect 38125 12459 38149 12493
rect 38187 12459 38193 12493
rect 38193 12459 38221 12493
rect 38259 12459 38261 12493
rect 38261 12459 38293 12493
rect 38331 12459 38363 12493
rect 38363 12459 38365 12493
rect 38403 12459 38431 12493
rect 38431 12459 38437 12493
rect 38475 12459 38499 12493
rect 38499 12459 38509 12493
rect 38547 12459 38581 12493
rect -1103 362 -1069 396
rect -1031 362 -997 396
rect -959 362 -925 396
rect -1188 293 -1154 327
rect -1188 221 -1154 255
rect -1188 149 -1154 183
rect -1188 77 -1154 111
rect -1188 5 -1154 39
rect -1188 -67 -1154 -33
rect -871 294 -837 328
rect -871 222 -837 256
rect -871 150 -837 184
rect -871 78 -837 112
rect -871 6 -837 40
rect -871 -66 -837 -32
rect -1105 -136 -1071 -102
rect -1033 -136 -999 -102
rect -961 -136 -927 -102
<< metal1 >>
rect 13280 17106 13352 17110
rect 13280 17054 13290 17106
rect 13342 17054 13352 17106
rect 13280 17050 13352 17054
rect 15638 17108 15698 17220
rect 15638 17056 15642 17108
rect 15694 17056 15698 17108
rect 15638 17046 15698 17056
rect 12484 16520 13584 16524
rect 12484 16468 12494 16520
rect 12546 16468 13584 16520
rect 12484 16464 13584 16468
rect 15632 16518 15704 16522
rect 15632 16466 15642 16518
rect 15694 16466 15704 16518
rect 15632 16462 15704 16466
rect -3432 14291 -1262 14548
rect -3432 13791 -2262 14291
rect -1762 13791 -1262 14291
rect -3432 13305 -1262 13791
rect -3432 1925 -3311 13305
rect -2939 1925 -1262 13305
rect 36712 13937 38688 13976
rect 36712 13903 36819 13937
rect 36853 13903 36891 13937
rect 36925 13903 36963 13937
rect 36997 13903 37035 13937
rect 37069 13903 37107 13937
rect 37141 13903 37179 13937
rect 37213 13903 37251 13937
rect 37285 13903 37323 13937
rect 37357 13903 37395 13937
rect 37429 13903 37467 13937
rect 37501 13903 37539 13937
rect 37573 13903 37611 13937
rect 37645 13903 37683 13937
rect 37717 13903 37755 13937
rect 37789 13903 37827 13937
rect 37861 13903 37899 13937
rect 37933 13903 37971 13937
rect 38005 13903 38043 13937
rect 38077 13903 38115 13937
rect 38149 13903 38187 13937
rect 38221 13903 38259 13937
rect 38293 13903 38331 13937
rect 38365 13903 38403 13937
rect 38437 13903 38475 13937
rect 38509 13903 38547 13937
rect 38581 13903 38688 13937
rect 36712 13864 38688 13903
rect 36712 13836 37434 13864
rect 36712 13791 36842 13836
rect 36712 13757 36751 13791
rect 36785 13757 36842 13791
rect 36712 13719 36842 13757
rect 36712 13685 36751 13719
rect 36785 13685 36842 13719
rect 36712 13647 36842 13685
rect 36712 13613 36751 13647
rect 36785 13613 36842 13647
rect 36712 13592 36842 13613
rect 37406 13592 37434 13836
rect 36712 13575 37434 13592
rect 36712 13541 36751 13575
rect 36785 13564 37434 13575
rect 37966 13836 38688 13864
rect 37966 13592 37994 13836
rect 38558 13791 38688 13836
rect 38558 13757 38615 13791
rect 38649 13757 38688 13791
rect 38558 13719 38688 13757
rect 38558 13685 38615 13719
rect 38649 13685 38688 13719
rect 38558 13647 38688 13685
rect 38558 13613 38615 13647
rect 38649 13613 38688 13647
rect 38558 13592 38688 13613
rect 37966 13575 38688 13592
rect 37966 13564 38615 13575
rect 36785 13541 36824 13564
rect 36712 13503 36824 13541
rect 36712 13469 36751 13503
rect 36785 13469 36824 13503
rect 36712 13431 36824 13469
rect 36712 13397 36751 13431
rect 36785 13397 36824 13431
rect 38576 13541 38615 13564
rect 38649 13541 38688 13575
rect 38576 13503 38688 13541
rect 38576 13469 38615 13503
rect 38649 13469 38688 13503
rect 38576 13431 38688 13469
rect 36712 13359 36824 13397
rect 36712 13325 36751 13359
rect 36785 13325 36824 13359
rect 36712 13287 36824 13325
rect 36712 13253 36751 13287
rect 36785 13253 36824 13287
rect 36890 13374 38514 13426
rect 36890 13322 36942 13374
rect 36994 13322 37006 13374
rect 37058 13322 37070 13374
rect 37122 13322 37134 13374
rect 37186 13322 37198 13374
rect 37250 13322 37262 13374
rect 37314 13322 37326 13374
rect 37378 13322 37390 13374
rect 37442 13322 37454 13374
rect 37506 13322 37518 13374
rect 37570 13322 37582 13374
rect 37634 13322 37646 13374
rect 37698 13322 37710 13374
rect 37762 13322 37774 13374
rect 37826 13322 37838 13374
rect 37890 13322 37902 13374
rect 37954 13322 37966 13374
rect 38018 13322 38030 13374
rect 38082 13322 38094 13374
rect 38146 13322 38158 13374
rect 38210 13322 38222 13374
rect 38274 13322 38286 13374
rect 38338 13322 38350 13374
rect 38402 13322 38414 13374
rect 38466 13322 38514 13374
rect 36890 13272 38514 13322
rect 38576 13397 38615 13431
rect 38649 13397 38688 13431
rect 38576 13359 38688 13397
rect 38576 13325 38615 13359
rect 38649 13325 38688 13359
rect 38576 13287 38688 13325
rect 36712 13215 36824 13253
rect 36712 13181 36751 13215
rect 36785 13181 36824 13215
rect 36712 13143 36824 13181
rect 36712 13109 36751 13143
rect 36785 13109 36824 13143
rect 36712 13071 36824 13109
rect 36712 13037 36751 13071
rect 36785 13037 36824 13071
rect 36712 12999 36824 13037
rect 36712 12965 36751 12999
rect 36785 12965 36824 12999
rect 36712 12927 36824 12965
rect 36712 12893 36751 12927
rect 36785 12893 36824 12927
rect 36712 12855 36824 12893
rect 36712 12821 36751 12855
rect 36785 12821 36824 12855
rect 36712 12783 36824 12821
rect 36712 12749 36751 12783
rect 36785 12749 36824 12783
rect 36712 12711 36824 12749
rect 36712 12677 36751 12711
rect 36785 12677 36824 12711
rect 36712 12639 36824 12677
rect 36712 12605 36751 12639
rect 36785 12605 36824 12639
rect 36712 12532 36824 12605
rect 36900 13130 37084 13272
rect 36900 12658 36960 13130
rect 37024 13044 37084 13130
rect 37414 12936 37474 13272
rect 37666 13190 37738 13194
rect 37666 13138 37676 13190
rect 37728 13138 37738 13190
rect 37666 13134 37738 13138
rect 37028 12658 37088 12753
rect 37156 12660 37216 12876
rect 37284 12662 37344 12748
rect 37540 12662 37600 12752
rect 37672 12662 37732 13134
rect 37930 12938 37990 13272
rect 38316 13135 38502 13272
rect 38316 13044 38376 13135
rect 37802 12662 37862 12750
rect 38058 12662 38118 12752
rect 36900 12598 37088 12658
rect 37150 12656 37222 12660
rect 37150 12604 37160 12656
rect 37212 12604 37222 12656
rect 37150 12600 37222 12604
rect 37284 12602 38118 12662
rect 38186 12660 38246 12844
rect 38314 12660 38374 12752
rect 38442 12660 38502 13135
rect 38180 12656 38252 12660
rect 38180 12604 38190 12656
rect 38242 12604 38252 12656
rect 38180 12600 38252 12604
rect 38314 12600 38502 12660
rect 38576 13253 38615 13287
rect 38649 13253 38688 13287
rect 38576 13215 38688 13253
rect 38576 13181 38615 13215
rect 38649 13181 38688 13215
rect 38576 13143 38688 13181
rect 38576 13109 38615 13143
rect 38649 13109 38688 13143
rect 38576 13071 38688 13109
rect 38576 13037 38615 13071
rect 38649 13037 38688 13071
rect 38576 12999 38688 13037
rect 38576 12965 38615 12999
rect 38649 12965 38688 12999
rect 38576 12927 38688 12965
rect 38576 12893 38615 12927
rect 38649 12893 38688 12927
rect 38576 12855 38688 12893
rect 38576 12821 38615 12855
rect 38649 12821 38688 12855
rect 38576 12783 38688 12821
rect 38576 12749 38615 12783
rect 38649 12749 38688 12783
rect 38576 12711 38688 12749
rect 38576 12677 38615 12711
rect 38649 12677 38688 12711
rect 38576 12639 38688 12677
rect 38576 12605 38615 12639
rect 38649 12605 38688 12639
rect 38576 12532 38688 12605
rect 36712 12493 38688 12532
rect 36712 12459 36819 12493
rect 36853 12459 36891 12493
rect 36925 12459 36963 12493
rect 36997 12459 37035 12493
rect 37069 12459 37107 12493
rect 37141 12459 37179 12493
rect 37213 12459 37251 12493
rect 37285 12459 37323 12493
rect 37357 12459 37395 12493
rect 37429 12459 37467 12493
rect 37501 12459 37539 12493
rect 37573 12459 37611 12493
rect 37645 12459 37683 12493
rect 37717 12459 37755 12493
rect 37789 12459 37827 12493
rect 37861 12459 37899 12493
rect 37933 12459 37971 12493
rect 38005 12459 38043 12493
rect 38077 12459 38115 12493
rect 38149 12459 38187 12493
rect 38221 12459 38259 12493
rect 38293 12459 38331 12493
rect 38365 12459 38403 12493
rect 38437 12459 38475 12493
rect 38509 12459 38547 12493
rect 38581 12459 38688 12493
rect 36712 12420 38688 12459
rect 12492 12062 12552 12072
rect 12492 12010 12496 12062
rect 12548 12010 12552 12062
rect 12492 12000 12552 12010
rect 13280 12062 13352 12066
rect 13280 12010 13290 12062
rect 13342 12010 13352 12062
rect 13280 12006 13352 12010
rect 12492 9970 12552 9980
rect 12492 9918 12496 9970
rect 12548 9918 12552 9970
rect 12492 9908 12552 9918
rect 12492 8728 12552 8738
rect 12492 8676 12496 8728
rect 12548 8676 12552 8728
rect 12492 8666 12552 8676
rect 12492 7492 12552 7502
rect 12492 7440 12496 7492
rect 12548 7440 12552 7492
rect 12492 7430 12552 7440
rect 12486 6966 12558 6970
rect 12486 6914 12496 6966
rect 12548 6914 12558 6966
rect 12486 6910 12558 6914
rect 13290 6966 13350 6976
rect 13290 6914 13294 6966
rect 13346 6914 13350 6966
rect 13290 6904 13350 6914
rect 13282 5382 13354 5386
rect 13282 5330 13292 5382
rect 13344 5330 13354 5382
rect 13282 5326 13354 5330
rect 41288 5248 41348 5402
rect 41288 5196 41292 5248
rect 41344 5196 41348 5248
rect 41288 5186 41348 5196
rect 11882 4726 11954 4730
rect 11882 4674 11892 4726
rect 11944 4674 11954 4726
rect 11882 4670 11954 4674
rect 13280 4726 13352 4730
rect 13280 4674 13290 4726
rect 13342 4674 13352 4726
rect 13280 4670 13352 4674
rect -3432 1842 -1262 1925
rect 8212 1394 8424 1454
rect 47814 1394 48076 1454
rect -1266 396 -810 414
rect -1266 394 -1103 396
rect -1364 362 -1103 394
rect -1069 362 -1031 396
rect -997 362 -959 396
rect -925 362 -810 396
rect -1364 344 -810 362
rect -1364 327 -1132 344
rect -1364 293 -1188 327
rect -1154 293 -1132 327
rect -1364 255 -1132 293
rect -894 328 -810 344
rect -894 294 -871 328
rect -837 294 -810 328
rect -1364 221 -1188 255
rect -1154 221 -1132 255
rect -1052 288 -980 292
rect -1052 236 -1042 288
rect -990 236 -980 288
rect -1052 232 -980 236
rect -894 256 -810 294
rect -1364 183 -1132 221
rect -1364 149 -1188 183
rect -1154 164 -1132 183
rect -894 222 -871 256
rect -837 222 -810 256
rect -894 184 -810 222
rect -998 166 -938 172
rect -1154 149 -1040 164
rect -1364 111 -1040 149
rect -1364 77 -1188 111
rect -1154 104 -1040 111
rect -1004 162 -932 166
rect -1004 110 -994 162
rect -942 110 -932 162
rect -1004 106 -932 110
rect -894 150 -871 184
rect -837 150 -810 184
rect -894 112 -810 150
rect -1154 77 -1132 104
rect -998 100 -938 106
rect -1364 39 -1132 77
rect -894 78 -871 112
rect -837 78 -810 112
rect -1364 5 -1188 39
rect -1154 5 -1132 39
rect -1364 -33 -1132 5
rect -1052 38 -980 42
rect -1052 -14 -1042 38
rect -990 -14 -980 38
rect -1052 -18 -980 -14
rect -894 40 -810 78
rect -894 6 -871 40
rect -837 6 -810 40
rect -1364 -67 -1188 -33
rect -1154 -67 -1132 -33
rect -1364 -68 -1132 -67
rect -894 -32 -810 6
rect -894 -66 -871 -32
rect -837 -66 -810 -32
rect -894 -68 -810 -66
rect -1364 -83 -808 -68
rect -1364 -120 -1192 -83
rect -1266 -135 -1192 -120
rect -1140 -135 -1128 -83
rect -1076 -102 -1064 -83
rect -1012 -102 -1000 -83
rect -948 -102 -936 -83
rect -1071 -135 -1064 -102
rect -884 -135 -872 -83
rect -820 -135 -808 -83
rect -1266 -136 -1105 -135
rect -1071 -136 -1033 -135
rect -999 -136 -961 -135
rect -927 -136 -808 -135
rect -1266 -152 -808 -136
rect -1266 -154 -1140 -152
rect -894 -154 -810 -152
<< via1 >>
rect 13290 17054 13342 17106
rect 15642 17056 15694 17108
rect 12494 16468 12546 16520
rect 15642 16466 15694 16518
rect -2262 13791 -1762 14291
rect -3311 1925 -2939 13305
rect 36842 13592 37406 13836
rect 37994 13592 38558 13836
rect 36942 13322 36994 13374
rect 37006 13322 37058 13374
rect 37070 13322 37122 13374
rect 37134 13322 37186 13374
rect 37198 13322 37250 13374
rect 37262 13322 37314 13374
rect 37326 13322 37378 13374
rect 37390 13322 37442 13374
rect 37454 13322 37506 13374
rect 37518 13322 37570 13374
rect 37582 13322 37634 13374
rect 37646 13322 37698 13374
rect 37710 13322 37762 13374
rect 37774 13322 37826 13374
rect 37838 13322 37890 13374
rect 37902 13322 37954 13374
rect 37966 13322 38018 13374
rect 38030 13322 38082 13374
rect 38094 13322 38146 13374
rect 38158 13322 38210 13374
rect 38222 13322 38274 13374
rect 38286 13322 38338 13374
rect 38350 13322 38402 13374
rect 38414 13322 38466 13374
rect 37676 13138 37728 13190
rect 37160 12604 37212 12656
rect 38190 12604 38242 12656
rect 12496 12010 12548 12062
rect 13290 12010 13342 12062
rect 12496 9918 12548 9970
rect 12496 8676 12548 8728
rect 12496 7440 12548 7492
rect 12496 6914 12548 6966
rect 13294 6914 13346 6966
rect 13292 5330 13344 5382
rect 41292 5196 41344 5248
rect 11892 4674 11944 4726
rect 13290 4674 13342 4726
rect -1042 236 -990 288
rect -994 110 -942 162
rect -1042 -14 -990 38
rect -1192 -135 -1140 -83
rect -1128 -102 -1076 -83
rect -1064 -102 -1012 -83
rect -1000 -102 -948 -83
rect -936 -102 -884 -83
rect -1128 -135 -1105 -102
rect -1105 -135 -1076 -102
rect -1064 -135 -1033 -102
rect -1033 -135 -1012 -102
rect -1000 -135 -999 -102
rect -999 -135 -961 -102
rect -961 -135 -948 -102
rect -936 -135 -927 -102
rect -927 -135 -884 -102
rect -872 -135 -820 -83
<< metal2 >>
rect 13286 17106 13346 17116
rect 13286 17054 13290 17106
rect 13342 17054 13346 17106
rect 12490 16520 12550 16530
rect 12490 16468 12494 16520
rect 12546 16468 12550 16520
rect 12490 16458 12550 16468
rect 13286 16400 13346 17054
rect 15632 17108 15704 17112
rect 15632 17056 15642 17108
rect 15694 17056 15704 17108
rect 15632 17052 15704 17056
rect 15638 16518 15698 17052
rect 15638 16466 15642 16518
rect 15694 16466 15698 16518
rect 15638 16456 15698 16466
rect 12492 15402 12552 15426
rect 12492 15346 12494 15402
rect 12550 15346 12552 15402
rect 12492 15236 12552 15346
rect -3432 14291 -1262 14548
rect -3432 13791 -2262 14291
rect -1762 13791 -1262 14291
rect -3432 13305 -1262 13791
rect 36824 13862 37424 13874
rect 36824 13836 36856 13862
rect 37392 13836 37424 13862
rect 36824 13592 36842 13836
rect 37406 13592 37424 13836
rect 36824 13566 36856 13592
rect 37392 13566 37424 13592
rect 36824 13554 37424 13566
rect 37976 13862 38576 13874
rect 37976 13836 38008 13862
rect 38544 13836 38576 13862
rect 37976 13592 37994 13836
rect 38558 13592 38576 13836
rect 37976 13566 38008 13592
rect 38544 13566 38576 13592
rect 37976 13554 38576 13566
rect -3432 13283 -3311 13305
rect -2939 13283 -1262 13305
rect -3432 1947 -3313 13283
rect -2937 1947 -1262 13283
rect 36890 13376 38514 13426
rect 36890 13374 36956 13376
rect 37012 13374 37036 13376
rect 37092 13374 37116 13376
rect 37172 13374 37196 13376
rect 37252 13374 37276 13376
rect 37332 13374 37356 13376
rect 37412 13374 37436 13376
rect 37492 13374 37516 13376
rect 37572 13374 37596 13376
rect 37652 13374 37676 13376
rect 37732 13374 37756 13376
rect 37812 13374 37836 13376
rect 37892 13374 37916 13376
rect 37972 13374 37996 13376
rect 38052 13374 38076 13376
rect 38132 13374 38156 13376
rect 38212 13374 38236 13376
rect 38292 13374 38316 13376
rect 38372 13374 38396 13376
rect 38452 13374 38514 13376
rect 36890 13322 36942 13374
rect 37186 13322 37196 13374
rect 37252 13322 37262 13374
rect 37506 13322 37516 13374
rect 37572 13322 37582 13374
rect 37826 13322 37836 13374
rect 37892 13322 37902 13374
rect 38146 13322 38156 13374
rect 38212 13322 38222 13374
rect 38466 13322 38514 13374
rect 36890 13320 36956 13322
rect 37012 13320 37036 13322
rect 37092 13320 37116 13322
rect 37172 13320 37196 13322
rect 37252 13320 37276 13322
rect 37332 13320 37356 13322
rect 37412 13320 37436 13322
rect 37492 13320 37516 13322
rect 37572 13320 37596 13322
rect 37652 13320 37676 13322
rect 37732 13320 37756 13322
rect 37812 13320 37836 13322
rect 37892 13320 37916 13322
rect 37972 13320 37996 13322
rect 38052 13320 38076 13322
rect 38132 13320 38156 13322
rect 38212 13320 38236 13322
rect 38292 13320 38316 13322
rect 38372 13320 38396 13322
rect 38452 13320 38514 13322
rect 36890 13272 38514 13320
rect 37672 13194 37732 13200
rect 39132 13194 39192 13203
rect 37672 13192 39192 13194
rect 37672 13190 39134 13192
rect 37672 13138 37676 13190
rect 37728 13138 39134 13190
rect 37672 13136 39134 13138
rect 39190 13136 39192 13192
rect 37672 13134 39192 13136
rect 37672 13128 37732 13134
rect 39132 13125 39192 13134
rect 37136 12660 37236 12678
rect 38186 12660 38246 12666
rect 37136 12656 38246 12660
rect 37136 12604 37160 12656
rect 37212 12604 38190 12656
rect 38242 12604 38246 12656
rect 37136 12600 38246 12604
rect 13286 12066 13346 12072
rect 12486 12062 13346 12066
rect 12486 12010 12496 12062
rect 12548 12010 13290 12062
rect 13342 12010 13346 12062
rect 12486 12006 13346 12010
rect 13286 12000 13346 12006
rect 12486 9970 13458 9974
rect 12486 9918 12496 9970
rect 12548 9918 13458 9970
rect 12486 9914 13458 9918
rect 34372 9972 34777 9974
rect 34372 9916 34710 9972
rect 34766 9916 34777 9972
rect 34372 9914 34777 9916
rect 12486 8728 13658 8732
rect 12486 8676 12496 8728
rect 12548 8676 13658 8728
rect 12486 8672 13658 8676
rect 12486 7492 13602 7496
rect 12486 7440 12496 7492
rect 12548 7440 13602 7492
rect 12486 7436 13602 7440
rect 12492 6970 12552 6976
rect 12492 6966 13356 6970
rect 12492 6914 12496 6966
rect 12548 6914 13294 6966
rect 13346 6914 13356 6966
rect 12492 6910 13356 6914
rect 12492 6904 12552 6910
rect 13288 5386 13348 5392
rect 12342 5382 13348 5386
rect 12342 5330 13292 5382
rect 13344 5330 13348 5382
rect 12342 5326 13348 5330
rect 13288 5320 13348 5326
rect 33930 5250 34179 5252
rect 33930 5194 34112 5250
rect 34168 5194 34179 5250
rect 33930 5192 34179 5194
rect 11888 4730 11948 4736
rect 13286 4730 13346 4736
rect 11888 4726 13346 4730
rect 11888 4674 11892 4726
rect 11944 4674 13290 4726
rect 13342 4674 13346 4726
rect 11888 4670 13346 4674
rect 11888 4664 11948 4670
rect 13286 4664 13346 4670
rect 11886 2776 11946 2954
rect 11886 2716 13454 2776
rect -3432 1925 -3311 1947
rect -2939 1925 -1262 1947
rect -3432 1842 -1262 1925
rect 264 1986 372 2003
rect 264 1930 290 1986
rect 346 1930 372 1986
rect 264 1913 372 1930
rect -1046 292 -986 298
rect -1046 288 -694 292
rect -1046 236 -1042 288
rect -990 236 -694 288
rect 37136 254 37236 12600
rect 38186 12594 38246 12600
rect 41279 6346 41444 6348
rect 41279 6290 41290 6346
rect 41346 6290 41444 6346
rect 41279 6288 41444 6290
rect 41288 5252 41348 5261
rect 41282 5250 41354 5252
rect 41282 5194 41290 5250
rect 41346 5194 41354 5250
rect 41282 5192 41354 5194
rect 41288 5183 41348 5192
rect 52714 2892 53274 2952
rect -1046 232 -694 236
rect 37127 232 37245 254
rect -1046 226 -986 232
rect -1012 164 -922 180
rect -1012 108 -995 164
rect -939 108 -922 164
rect -1012 94 -922 108
rect -1046 42 -986 48
rect -834 42 -774 232
rect 37127 176 37158 232
rect 37214 176 37245 232
rect 37127 154 37245 176
rect -1046 38 -774 42
rect -1046 -14 -1042 38
rect -990 -14 -774 38
rect -1046 -18 -774 -14
rect -1046 -24 -986 -18
rect -1212 -81 -806 -64
rect -1212 -137 -1194 -81
rect -1138 -83 -1114 -81
rect -1058 -83 -1034 -81
rect -978 -83 -954 -81
rect -898 -83 -874 -81
rect -1138 -135 -1128 -83
rect -884 -135 -874 -83
rect -1138 -137 -1114 -135
rect -1058 -137 -1034 -135
rect -978 -137 -954 -135
rect -898 -137 -874 -135
rect -818 -137 -806 -81
rect -1212 -154 -806 -137
<< via2 >>
rect 12494 15346 12550 15402
rect -2240 13813 -1784 14269
rect 36856 13836 37392 13862
rect 36856 13592 37392 13836
rect 36856 13566 37392 13592
rect 38008 13836 38544 13862
rect 38008 13592 38544 13836
rect 38008 13566 38544 13592
rect -3313 1947 -3311 13283
rect -3311 1947 -2939 13283
rect -2939 1947 -2937 13283
rect 36956 13374 37012 13376
rect 37036 13374 37092 13376
rect 37116 13374 37172 13376
rect 37196 13374 37252 13376
rect 37276 13374 37332 13376
rect 37356 13374 37412 13376
rect 37436 13374 37492 13376
rect 37516 13374 37572 13376
rect 37596 13374 37652 13376
rect 37676 13374 37732 13376
rect 37756 13374 37812 13376
rect 37836 13374 37892 13376
rect 37916 13374 37972 13376
rect 37996 13374 38052 13376
rect 38076 13374 38132 13376
rect 38156 13374 38212 13376
rect 38236 13374 38292 13376
rect 38316 13374 38372 13376
rect 38396 13374 38452 13376
rect 36956 13322 36994 13374
rect 36994 13322 37006 13374
rect 37006 13322 37012 13374
rect 37036 13322 37058 13374
rect 37058 13322 37070 13374
rect 37070 13322 37092 13374
rect 37116 13322 37122 13374
rect 37122 13322 37134 13374
rect 37134 13322 37172 13374
rect 37196 13322 37198 13374
rect 37198 13322 37250 13374
rect 37250 13322 37252 13374
rect 37276 13322 37314 13374
rect 37314 13322 37326 13374
rect 37326 13322 37332 13374
rect 37356 13322 37378 13374
rect 37378 13322 37390 13374
rect 37390 13322 37412 13374
rect 37436 13322 37442 13374
rect 37442 13322 37454 13374
rect 37454 13322 37492 13374
rect 37516 13322 37518 13374
rect 37518 13322 37570 13374
rect 37570 13322 37572 13374
rect 37596 13322 37634 13374
rect 37634 13322 37646 13374
rect 37646 13322 37652 13374
rect 37676 13322 37698 13374
rect 37698 13322 37710 13374
rect 37710 13322 37732 13374
rect 37756 13322 37762 13374
rect 37762 13322 37774 13374
rect 37774 13322 37812 13374
rect 37836 13322 37838 13374
rect 37838 13322 37890 13374
rect 37890 13322 37892 13374
rect 37916 13322 37954 13374
rect 37954 13322 37966 13374
rect 37966 13322 37972 13374
rect 37996 13322 38018 13374
rect 38018 13322 38030 13374
rect 38030 13322 38052 13374
rect 38076 13322 38082 13374
rect 38082 13322 38094 13374
rect 38094 13322 38132 13374
rect 38156 13322 38158 13374
rect 38158 13322 38210 13374
rect 38210 13322 38212 13374
rect 38236 13322 38274 13374
rect 38274 13322 38286 13374
rect 38286 13322 38292 13374
rect 38316 13322 38338 13374
rect 38338 13322 38350 13374
rect 38350 13322 38372 13374
rect 38396 13322 38402 13374
rect 38402 13322 38414 13374
rect 38414 13322 38452 13374
rect 36956 13320 37012 13322
rect 37036 13320 37092 13322
rect 37116 13320 37172 13322
rect 37196 13320 37252 13322
rect 37276 13320 37332 13322
rect 37356 13320 37412 13322
rect 37436 13320 37492 13322
rect 37516 13320 37572 13322
rect 37596 13320 37652 13322
rect 37676 13320 37732 13322
rect 37756 13320 37812 13322
rect 37836 13320 37892 13322
rect 37916 13320 37972 13322
rect 37996 13320 38052 13322
rect 38076 13320 38132 13322
rect 38156 13320 38212 13322
rect 38236 13320 38292 13322
rect 38316 13320 38372 13322
rect 38396 13320 38452 13322
rect 39134 13136 39190 13192
rect 34710 9916 34766 9972
rect 34112 5194 34168 5250
rect 290 1930 346 1986
rect 41290 6290 41346 6346
rect 41290 5248 41346 5250
rect 41290 5196 41292 5248
rect 41292 5196 41344 5248
rect 41344 5196 41346 5248
rect 41290 5194 41346 5196
rect -995 162 -939 164
rect -995 110 -994 162
rect -994 110 -942 162
rect -942 110 -939 162
rect -995 108 -939 110
rect 37158 176 37214 232
rect -1194 -83 -1138 -81
rect -1114 -83 -1058 -81
rect -1034 -83 -978 -81
rect -954 -83 -898 -81
rect -874 -83 -818 -81
rect -1194 -135 -1192 -83
rect -1192 -135 -1140 -83
rect -1140 -135 -1138 -83
rect -1114 -135 -1076 -83
rect -1076 -135 -1064 -83
rect -1064 -135 -1058 -83
rect -1034 -135 -1012 -83
rect -1012 -135 -1000 -83
rect -1000 -135 -978 -83
rect -954 -135 -948 -83
rect -948 -135 -936 -83
rect -936 -135 -898 -83
rect -874 -135 -872 -83
rect -872 -135 -820 -83
rect -820 -135 -818 -83
rect -1194 -137 -1138 -135
rect -1114 -137 -1058 -135
rect -1034 -137 -978 -135
rect -954 -137 -898 -135
rect -874 -137 -818 -135
<< metal3 >>
rect 12430 15424 12624 15426
rect 12430 15409 12636 15424
rect 12430 15345 12490 15409
rect 12554 15345 12636 15409
rect 12430 15328 12636 15345
rect 12430 15324 12624 15328
rect -3634 14544 -2794 14660
rect -16568 14361 -1528 14544
rect -16568 14355 -2341 14361
rect -16568 13731 -16380 14355
rect -15756 13737 -2341 14355
rect -1717 13737 -1528 14361
rect 52113 14346 52211 14351
rect 39110 14328 52212 14346
rect 39110 14264 52130 14328
rect 52194 14264 52212 14328
rect 39110 14246 52212 14264
rect -15756 13731 -1528 13737
rect -16568 13283 -1528 13731
rect 36814 13862 37434 13869
rect 36814 13826 36856 13862
rect 37392 13826 37434 13862
rect 36814 13602 36852 13826
rect 37396 13602 37434 13826
rect 36814 13566 36856 13602
rect 37392 13566 37434 13602
rect 36814 13559 37434 13566
rect 37966 13862 38586 13869
rect 37966 13826 38008 13862
rect 38544 13826 38586 13862
rect 37966 13602 38004 13826
rect 38548 13602 38586 13826
rect 37966 13566 38008 13602
rect 38544 13566 38586 13602
rect 37966 13559 38586 13566
rect -16568 1947 -3313 13283
rect -2937 1947 -1528 13283
rect 36890 13380 38514 13426
rect 36890 13316 36952 13380
rect 37016 13316 37032 13380
rect 37096 13316 37112 13380
rect 37176 13316 37192 13380
rect 37256 13316 37272 13380
rect 37336 13316 37352 13380
rect 37416 13316 37432 13380
rect 37496 13316 37512 13380
rect 37576 13316 37592 13380
rect 37656 13316 37672 13380
rect 37736 13316 37752 13380
rect 37816 13316 37832 13380
rect 37896 13316 37912 13380
rect 37976 13316 37992 13380
rect 38056 13316 38072 13380
rect 38136 13316 38152 13380
rect 38216 13316 38232 13380
rect 38296 13316 38312 13380
rect 38376 13316 38392 13380
rect 38456 13316 38514 13380
rect 36890 13272 38514 13316
rect 39110 13192 39210 14246
rect 52113 14241 52211 14246
rect 39110 13136 39134 13192
rect 39190 13136 39210 13192
rect 39110 13114 39210 13136
rect 34688 9972 41370 9992
rect 34688 9916 34710 9972
rect 34766 9916 41370 9972
rect 34688 9892 41370 9916
rect 41270 6346 41370 9892
rect 41270 6290 41290 6346
rect 41346 6290 41370 6346
rect 41270 6270 41370 6290
rect 34086 5250 41380 5270
rect 34086 5194 34112 5250
rect 34168 5194 41290 5250
rect 41346 5194 41380 5250
rect 34086 5170 41380 5194
rect -16568 360 -1528 1947
rect 268 1986 368 2008
rect 268 1930 290 1986
rect 346 1930 368 1986
rect 268 634 368 1930
rect -1016 496 -916 520
rect 268 513 370 634
rect -1016 432 -998 496
rect -934 432 -916 496
rect -16568 -458 -2656 360
rect -1016 164 -916 432
rect 263 496 373 513
rect 263 432 286 496
rect 350 432 373 496
rect 263 415 373 432
rect 268 414 370 415
rect -1016 108 -995 164
rect -939 108 -916 164
rect 270 254 370 414
rect 37131 254 37241 259
rect 270 232 37241 254
rect 270 176 37158 232
rect 37214 176 37241 232
rect 270 154 37241 176
rect 37131 149 37241 154
rect -1016 94 -916 108
rect -1212 -77 -806 -64
rect -1212 -141 -1198 -77
rect -1134 -141 -1118 -77
rect -1054 -141 -1038 -77
rect -974 -141 -958 -77
rect -894 -141 -878 -77
rect -814 -141 -806 -77
rect -1212 -154 -806 -141
<< via3 >>
rect 12490 15402 12554 15409
rect 12490 15346 12494 15402
rect 12494 15346 12550 15402
rect 12550 15346 12554 15402
rect 12490 15345 12554 15346
rect -16380 13731 -15756 14355
rect -2341 14269 -1717 14361
rect -2341 13813 -2240 14269
rect -2240 13813 -1784 14269
rect -1784 13813 -1717 14269
rect -2341 13737 -1717 13813
rect 52130 14264 52194 14328
rect 36852 13602 36856 13826
rect 36856 13602 37392 13826
rect 37392 13602 37396 13826
rect 38004 13602 38008 13826
rect 38008 13602 38544 13826
rect 38544 13602 38548 13826
rect 36952 13376 37016 13380
rect 36952 13320 36956 13376
rect 36956 13320 37012 13376
rect 37012 13320 37016 13376
rect 36952 13316 37016 13320
rect 37032 13376 37096 13380
rect 37032 13320 37036 13376
rect 37036 13320 37092 13376
rect 37092 13320 37096 13376
rect 37032 13316 37096 13320
rect 37112 13376 37176 13380
rect 37112 13320 37116 13376
rect 37116 13320 37172 13376
rect 37172 13320 37176 13376
rect 37112 13316 37176 13320
rect 37192 13376 37256 13380
rect 37192 13320 37196 13376
rect 37196 13320 37252 13376
rect 37252 13320 37256 13376
rect 37192 13316 37256 13320
rect 37272 13376 37336 13380
rect 37272 13320 37276 13376
rect 37276 13320 37332 13376
rect 37332 13320 37336 13376
rect 37272 13316 37336 13320
rect 37352 13376 37416 13380
rect 37352 13320 37356 13376
rect 37356 13320 37412 13376
rect 37412 13320 37416 13376
rect 37352 13316 37416 13320
rect 37432 13376 37496 13380
rect 37432 13320 37436 13376
rect 37436 13320 37492 13376
rect 37492 13320 37496 13376
rect 37432 13316 37496 13320
rect 37512 13376 37576 13380
rect 37512 13320 37516 13376
rect 37516 13320 37572 13376
rect 37572 13320 37576 13376
rect 37512 13316 37576 13320
rect 37592 13376 37656 13380
rect 37592 13320 37596 13376
rect 37596 13320 37652 13376
rect 37652 13320 37656 13376
rect 37592 13316 37656 13320
rect 37672 13376 37736 13380
rect 37672 13320 37676 13376
rect 37676 13320 37732 13376
rect 37732 13320 37736 13376
rect 37672 13316 37736 13320
rect 37752 13376 37816 13380
rect 37752 13320 37756 13376
rect 37756 13320 37812 13376
rect 37812 13320 37816 13376
rect 37752 13316 37816 13320
rect 37832 13376 37896 13380
rect 37832 13320 37836 13376
rect 37836 13320 37892 13376
rect 37892 13320 37896 13376
rect 37832 13316 37896 13320
rect 37912 13376 37976 13380
rect 37912 13320 37916 13376
rect 37916 13320 37972 13376
rect 37972 13320 37976 13376
rect 37912 13316 37976 13320
rect 37992 13376 38056 13380
rect 37992 13320 37996 13376
rect 37996 13320 38052 13376
rect 38052 13320 38056 13376
rect 37992 13316 38056 13320
rect 38072 13376 38136 13380
rect 38072 13320 38076 13376
rect 38076 13320 38132 13376
rect 38132 13320 38136 13376
rect 38072 13316 38136 13320
rect 38152 13376 38216 13380
rect 38152 13320 38156 13376
rect 38156 13320 38212 13376
rect 38212 13320 38216 13376
rect 38152 13316 38216 13320
rect 38232 13376 38296 13380
rect 38232 13320 38236 13376
rect 38236 13320 38292 13376
rect 38292 13320 38296 13376
rect 38232 13316 38296 13320
rect 38312 13376 38376 13380
rect 38312 13320 38316 13376
rect 38316 13320 38372 13376
rect 38372 13320 38376 13376
rect 38312 13316 38376 13320
rect 38392 13376 38456 13380
rect 38392 13320 38396 13376
rect 38396 13320 38452 13376
rect 38452 13320 38456 13376
rect 38392 13316 38456 13320
rect -998 432 -934 496
rect 286 432 350 496
rect -1198 -81 -1134 -77
rect -1198 -137 -1194 -81
rect -1194 -137 -1138 -81
rect -1138 -137 -1134 -81
rect -1198 -141 -1134 -137
rect -1118 -81 -1054 -77
rect -1118 -137 -1114 -81
rect -1114 -137 -1058 -81
rect -1058 -137 -1054 -81
rect -1118 -141 -1054 -137
rect -1038 -81 -974 -77
rect -1038 -137 -1034 -81
rect -1034 -137 -978 -81
rect -978 -137 -974 -81
rect -1038 -141 -974 -137
rect -958 -81 -894 -77
rect -958 -137 -954 -81
rect -954 -137 -898 -81
rect -898 -137 -894 -81
rect -958 -141 -894 -137
rect -878 -81 -814 -77
rect -878 -137 -874 -81
rect -874 -137 -818 -81
rect -818 -137 -814 -81
rect -878 -141 -814 -137
<< mimcap >>
rect -15382 14256 -9182 14344
rect -15382 14032 -9494 14256
rect -9270 14032 -9182 14256
rect -15382 13944 -9182 14032
rect -8982 14256 -2782 14344
rect -8982 14032 -3094 14256
rect -2870 14032 -2782 14256
rect -8982 13944 -2782 14032
rect -16468 13294 -15668 13362
rect -16468 7630 -15980 13294
rect -15756 7630 -15668 13294
rect -2424 13294 -1624 13362
rect -14528 12356 -9328 12444
rect -14528 7732 -9640 12356
rect -9416 7732 -9328 12356
rect -14528 7644 -9328 7732
rect -8928 12356 -3728 12444
rect -8928 7732 -4040 12356
rect -3816 7732 -3728 12356
rect -8928 7644 -3728 7732
rect -16468 7562 -15668 7630
rect -2424 7630 -1936 13294
rect -1712 7630 -1624 13294
rect -2424 7562 -1624 7630
rect -16468 6802 -15668 6870
rect -16468 1138 -15980 6802
rect -15756 1138 -15668 6802
rect -14528 6756 -9328 6844
rect -14528 2132 -9640 6756
rect -9416 2132 -9328 6756
rect -14528 2044 -9328 2132
rect -8928 6756 -3728 6844
rect -8928 2132 -4040 6756
rect -3816 2132 -3728 6756
rect -8928 2044 -3728 2132
rect -2424 6802 -1624 6870
rect -16468 1070 -15668 1138
rect -2424 1138 -1936 6802
rect -1712 1138 -1624 6802
rect -2424 1070 -1624 1138
rect -15882 356 -9682 444
rect -15882 132 -9994 356
rect -9770 132 -9682 356
rect -15882 44 -9682 132
rect -9482 356 -3282 444
rect -9482 132 -3594 356
rect -3370 132 -3282 356
rect -9482 44 -3282 132
<< mimcapcontact >>
rect -9494 14032 -9270 14256
rect -3094 14032 -2870 14256
rect -15980 7630 -15756 13294
rect -9640 7732 -9416 12356
rect -4040 7732 -3816 12356
rect -1936 7630 -1712 13294
rect -15980 1138 -15756 6802
rect -9640 2132 -9416 6756
rect -4040 2132 -3816 6756
rect -1936 1138 -1712 6802
rect -9994 132 -9770 356
rect -3594 132 -3370 356
<< metal4 >>
rect 34964 30648 37598 30770
rect 34964 30092 35354 30648
rect 35910 30092 37598 30648
rect 34964 29970 37598 30092
rect 12486 15409 12558 15410
rect 12486 15345 12490 15409
rect 12554 15345 12558 15409
rect 12486 15344 12558 15345
rect -4196 14544 -1528 14984
rect -16568 14361 -1528 14544
rect -16568 14355 -2341 14361
rect -16568 13731 -16380 14355
rect -15756 14256 -2341 14355
rect -15756 14032 -9494 14256
rect -9270 14032 -3094 14256
rect -2870 14032 -2341 14256
rect -15756 13737 -2341 14032
rect -1717 13737 -1528 14361
rect 52112 14328 52212 15426
rect 52112 14264 52130 14328
rect 52194 14264 52212 14328
rect 52112 14246 52212 14264
rect 35516 14048 36670 14050
rect -15756 13731 -1528 13737
rect -16568 13368 -1528 13731
rect -16568 13294 -15386 13368
rect -16568 7630 -15980 13294
rect -15756 7630 -15386 13294
rect -2828 13294 -1528 13368
rect -16568 6802 -15386 7630
rect -16568 1138 -15980 6802
rect -15756 1138 -15386 6802
rect -14628 12356 -3628 12544
rect -14628 7732 -9640 12356
rect -9416 7732 -4040 12356
rect -3816 7732 -3628 12356
rect -14628 6756 -3628 7732
rect -14628 2132 -9640 6756
rect -9416 2132 -4040 6756
rect -3816 2132 -3628 6756
rect -14628 1544 -3628 2132
rect -2828 7630 -1936 13294
rect -1712 7630 -1528 13294
rect 35232 13930 38760 14048
rect 35232 13374 35354 13930
rect 35910 13826 38760 13930
rect 35910 13602 36852 13826
rect 37396 13602 38004 13826
rect 38548 13602 38760 13826
rect 35910 13380 38760 13602
rect 35910 13374 36952 13380
rect 35232 13316 36952 13374
rect 37016 13316 37032 13380
rect 37096 13316 37112 13380
rect 37176 13316 37192 13380
rect 37256 13316 37272 13380
rect 37336 13316 37352 13380
rect 37416 13316 37432 13380
rect 37496 13316 37512 13380
rect 37576 13316 37592 13380
rect 37656 13316 37672 13380
rect 37736 13316 37752 13380
rect 37816 13316 37832 13380
rect 37896 13316 37912 13380
rect 37976 13316 37992 13380
rect 38056 13316 38072 13380
rect 38136 13316 38152 13380
rect 38216 13316 38232 13380
rect 38296 13316 38312 13380
rect 38376 13316 38392 13380
rect 38456 13316 38760 13380
rect 35232 13248 38760 13316
rect -2828 6802 -1528 7630
rect -2828 1760 -1936 6802
rect -3754 1496 -3628 1544
rect -3754 1396 -2814 1496
rect -16568 706 -15386 1138
rect -16568 620 -3244 706
rect -16566 356 -3244 620
rect -16566 132 -9994 356
rect -9770 132 -3594 356
rect -3370 132 -3244 356
rect -2914 340 -2814 1396
rect -2458 1138 -1936 1760
rect -1712 1138 -1528 6802
rect -2458 1002 -1528 1138
rect -2458 610 -1952 1002
rect -1017 514 -915 515
rect -1400 496 368 514
rect -1400 432 -998 496
rect -934 432 286 496
rect 350 432 368 496
rect -1400 414 368 432
rect -1400 340 -1300 414
rect -1017 413 -915 414
rect -2914 240 -1300 340
rect -16566 -32 -3244 132
rect -2652 -32 -1544 -30
rect -16566 -42 -1544 -32
rect -16566 -278 -16353 -42
rect -16117 -139 -1544 -42
rect -16117 -278 -1992 -139
rect -16566 -375 -1992 -278
rect -1756 -375 -1544 -139
rect -1198 -77 -814 -76
rect -1134 -141 -1118 -77
rect -1054 -141 -1038 -77
rect -974 -141 -958 -77
rect -894 -141 -878 -77
rect -1198 -142 -814 -141
rect -16566 -830 -1544 -375
rect 33872 -830 38596 -30
<< via4 >>
rect 35354 30092 35910 30648
rect -16346 13765 -15790 14321
rect -2307 13771 -1751 14327
rect 35354 13374 35910 13930
rect -16353 -278 -16117 -42
rect -1992 -375 -1756 -139
<< mimcap2 >>
rect -15382 13862 -9582 14344
rect -15382 13626 -15320 13862
rect -9644 13626 -9582 13862
rect -15382 13544 -9582 13626
rect -8982 13862 -3182 14344
rect -8982 13626 -8920 13862
rect -3244 13626 -3182 13862
rect -8982 13544 -3182 13626
rect -16468 7480 -16068 13362
rect -16468 7244 -16386 7480
rect -16150 7244 -16068 7480
rect -14528 7562 -9728 12444
rect -14528 7326 -14326 7562
rect -9930 7326 -9728 7562
rect -14528 7244 -9728 7326
rect -8928 7562 -4128 12444
rect -8928 7326 -8726 7562
rect -4330 7326 -4128 7562
rect -8928 7244 -4128 7326
rect -2424 7480 -2024 13362
rect -2424 7244 -2342 7480
rect -2106 7244 -2024 7480
rect -16468 7162 -16068 7244
rect -2424 7162 -2024 7244
rect -16468 988 -16068 6870
rect -14528 1962 -9728 6844
rect -14528 1726 -14326 1962
rect -9930 1726 -9728 1962
rect -14528 1644 -9728 1726
rect -8928 1962 -4128 6844
rect -8928 1726 -8726 1962
rect -4330 1726 -4128 1962
rect -8928 1644 -4128 1726
rect -16468 752 -16386 988
rect -16150 752 -16068 988
rect -16468 670 -16068 752
rect -2424 988 -2024 6870
rect -2424 752 -2342 988
rect -2106 752 -2024 988
rect -2424 670 -2024 752
rect -15882 -38 -10082 444
rect -15882 -274 -15820 -38
rect -10144 -274 -10082 -38
rect -15882 -356 -10082 -274
rect -9482 -38 -3682 444
rect -9482 -274 -9420 -38
rect -3744 -274 -3682 -38
rect -9482 -356 -3682 -274
<< mimcap2contact >>
rect -15320 13626 -9644 13862
rect -8920 13626 -3244 13862
rect -16386 7244 -16150 7480
rect -14326 7326 -9930 7562
rect -8726 7326 -4330 7562
rect -2342 7244 -2106 7480
rect -14326 1726 -9930 1962
rect -8726 1726 -4330 1962
rect -16386 752 -16150 988
rect -2342 752 -2106 988
rect -15820 -274 -10144 -38
rect -9420 -274 -3744 -38
<< metal5 >>
rect 35208 30648 36056 30794
rect 35208 30092 35354 30648
rect 35910 30092 36056 30648
rect 35208 29946 36056 30092
rect -16568 14327 -1528 14544
rect -16568 14321 -2307 14327
rect -16568 13765 -16346 14321
rect -15790 13862 -2307 14321
rect -15790 13765 -15320 13862
rect -16568 13626 -15320 13765
rect -9644 13626 -8920 13862
rect -3244 13771 -2307 13862
rect -1751 13771 -1528 14327
rect -3244 13626 -1528 13771
rect -16568 13368 -1528 13626
rect -16568 7562 -3364 13368
rect -16568 7480 -14326 7562
rect -16568 7244 -16386 7480
rect -16150 7326 -14326 7480
rect -9930 7326 -8726 7562
rect -4330 7326 -3364 7562
rect -16150 7244 -3364 7326
rect -16568 1962 -3364 7244
rect -16568 1726 -14326 1962
rect -9930 1726 -8726 1962
rect -4330 1844 -3364 1962
rect -2828 7480 -1528 13368
rect 35232 13930 36032 29946
rect 35232 13374 35354 13930
rect 35910 13374 36032 13930
rect 35232 13252 36032 13374
rect -2828 7244 -2342 7480
rect -2106 7244 -1528 7480
rect -2828 1844 -1528 7244
rect -4330 1726 -1528 1844
rect -16568 988 -1528 1726
rect -16568 752 -16386 988
rect -16150 752 -2342 988
rect -2106 752 -1528 988
rect -16568 360 -1528 752
rect -16568 -38 -1530 360
rect -16568 -42 -15820 -38
rect -16568 -278 -16353 -42
rect -16117 -274 -15820 -42
rect -10144 -274 -9420 -38
rect -3744 -139 -1530 -38
rect -3744 -274 -1992 -139
rect -16117 -278 -1992 -274
rect -16568 -375 -1992 -278
rect -1756 -375 -1530 -139
rect -16568 -458 -1530 -375
use se_fold_casc_wide_swing_ota  se_fold_casc_wide_swing_ota_1
timestamp 1626065694
transform 1 0 10950 0 1 26370
box -15168 -27248 25000 4400
use se_fold_casc_wide_swing_ota  se_fold_casc_wide_swing_ota_0
timestamp 1626065694
transform 1 0 51950 0 1 26370
box -15168 -27248 25000 4400
use sky130_fd_pr__nfet_01v8_HFLVLW  sky130_fd_pr__nfet_01v8_HFLVLW_0
timestamp 1626065694
transform 1 0 -1013 0 1 137
box -201 -299 201 285
use sky130_fd_pr__pfet_01v8_RC2RSP  sky130_fd_pr__pfet_01v8_RC2RSP_0
timestamp 1626065694
transform 1 0 37701 0 1 12898
box -839 -200 839 200
<< labels >>
flabel metal2 s 38146 12624 38158 12636 1 FreeSans 600 0 0 0 vpeakh
flabel metal1 s 37310 12672 37326 12682 1 FreeSans 600 0 0 0 verr
flabel metal4 s 37536 14028 37548 14038 1 FreeSans 600 0 0 0 VDD
flabel metal2 s -742 256 -736 264 1 FreeSans 600 0 0 0 rst
flabel metal2 s 53200 2918 53216 2930 1 FreeSans 600 0 0 0 vin
flabel metal2 s 12516 15272 12528 15284 1 FreeSans 600 0 0 0 vpeak_out
flabel metal4 s 36274 -344 36322 -292 1 FreeSans 600 0 0 0 VSS
flabel metal1 s 8324 1414 8342 1424 1 FreeSans 600 0 0 0 ibiasn2
flabel metal1 s 47952 1414 47972 1428 1 FreeSans 600 0 0 0 ibiasn1
flabel metal4 s -1544 284 -1530 294 1 FreeSans 600 0 0 0 vpeak
<< properties >>
string FIXED_BBOX 648 33828 2512 35272
<< end >>
