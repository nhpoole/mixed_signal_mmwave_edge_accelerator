magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -2605 -1448 2605 1448
<< pwell >>
rect -1345 -126 1345 126
<< nmoslvt >>
rect -1261 -100 -1061 100
rect -1003 -100 -803 100
rect -745 -100 -545 100
rect -487 -100 -287 100
rect -229 -100 -29 100
rect 29 -100 229 100
rect 287 -100 487 100
rect 545 -100 745 100
rect 803 -100 1003 100
rect 1061 -100 1261 100
<< ndiff >>
rect -1319 85 -1261 100
rect -1319 51 -1307 85
rect -1273 51 -1261 85
rect -1319 17 -1261 51
rect -1319 -17 -1307 17
rect -1273 -17 -1261 17
rect -1319 -51 -1261 -17
rect -1319 -85 -1307 -51
rect -1273 -85 -1261 -51
rect -1319 -100 -1261 -85
rect -1061 85 -1003 100
rect -1061 51 -1049 85
rect -1015 51 -1003 85
rect -1061 17 -1003 51
rect -1061 -17 -1049 17
rect -1015 -17 -1003 17
rect -1061 -51 -1003 -17
rect -1061 -85 -1049 -51
rect -1015 -85 -1003 -51
rect -1061 -100 -1003 -85
rect -803 85 -745 100
rect -803 51 -791 85
rect -757 51 -745 85
rect -803 17 -745 51
rect -803 -17 -791 17
rect -757 -17 -745 17
rect -803 -51 -745 -17
rect -803 -85 -791 -51
rect -757 -85 -745 -51
rect -803 -100 -745 -85
rect -545 85 -487 100
rect -545 51 -533 85
rect -499 51 -487 85
rect -545 17 -487 51
rect -545 -17 -533 17
rect -499 -17 -487 17
rect -545 -51 -487 -17
rect -545 -85 -533 -51
rect -499 -85 -487 -51
rect -545 -100 -487 -85
rect -287 85 -229 100
rect -287 51 -275 85
rect -241 51 -229 85
rect -287 17 -229 51
rect -287 -17 -275 17
rect -241 -17 -229 17
rect -287 -51 -229 -17
rect -287 -85 -275 -51
rect -241 -85 -229 -51
rect -287 -100 -229 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 229 85 287 100
rect 229 51 241 85
rect 275 51 287 85
rect 229 17 287 51
rect 229 -17 241 17
rect 275 -17 287 17
rect 229 -51 287 -17
rect 229 -85 241 -51
rect 275 -85 287 -51
rect 229 -100 287 -85
rect 487 85 545 100
rect 487 51 499 85
rect 533 51 545 85
rect 487 17 545 51
rect 487 -17 499 17
rect 533 -17 545 17
rect 487 -51 545 -17
rect 487 -85 499 -51
rect 533 -85 545 -51
rect 487 -100 545 -85
rect 745 85 803 100
rect 745 51 757 85
rect 791 51 803 85
rect 745 17 803 51
rect 745 -17 757 17
rect 791 -17 803 17
rect 745 -51 803 -17
rect 745 -85 757 -51
rect 791 -85 803 -51
rect 745 -100 803 -85
rect 1003 85 1061 100
rect 1003 51 1015 85
rect 1049 51 1061 85
rect 1003 17 1061 51
rect 1003 -17 1015 17
rect 1049 -17 1061 17
rect 1003 -51 1061 -17
rect 1003 -85 1015 -51
rect 1049 -85 1061 -51
rect 1003 -100 1061 -85
rect 1261 85 1319 100
rect 1261 51 1273 85
rect 1307 51 1319 85
rect 1261 17 1319 51
rect 1261 -17 1273 17
rect 1307 -17 1319 17
rect 1261 -51 1319 -17
rect 1261 -85 1273 -51
rect 1307 -85 1319 -51
rect 1261 -100 1319 -85
<< ndiffc >>
rect -1307 51 -1273 85
rect -1307 -17 -1273 17
rect -1307 -85 -1273 -51
rect -1049 51 -1015 85
rect -1049 -17 -1015 17
rect -1049 -85 -1015 -51
rect -791 51 -757 85
rect -791 -17 -757 17
rect -791 -85 -757 -51
rect -533 51 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -51
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
rect 499 51 533 85
rect 499 -17 533 17
rect 499 -85 533 -51
rect 757 51 791 85
rect 757 -17 791 17
rect 757 -85 791 -51
rect 1015 51 1049 85
rect 1015 -17 1049 17
rect 1015 -85 1049 -51
rect 1273 51 1307 85
rect 1273 -17 1307 17
rect 1273 -85 1307 -51
<< poly >>
rect -1227 172 -1095 188
rect -1227 155 -1178 172
rect -1261 138 -1178 155
rect -1144 155 -1095 172
rect -969 172 -837 188
rect -969 155 -920 172
rect -1144 138 -1061 155
rect -1261 100 -1061 138
rect -1003 138 -920 155
rect -886 155 -837 172
rect -711 172 -579 188
rect -711 155 -662 172
rect -886 138 -803 155
rect -1003 100 -803 138
rect -745 138 -662 155
rect -628 155 -579 172
rect -453 172 -321 188
rect -453 155 -404 172
rect -628 138 -545 155
rect -745 100 -545 138
rect -487 138 -404 155
rect -370 155 -321 172
rect -195 172 -63 188
rect -195 155 -146 172
rect -370 138 -287 155
rect -487 100 -287 138
rect -229 138 -146 155
rect -112 155 -63 172
rect 63 172 195 188
rect 63 155 112 172
rect -112 138 -29 155
rect -229 100 -29 138
rect 29 138 112 155
rect 146 155 195 172
rect 321 172 453 188
rect 321 155 370 172
rect 146 138 229 155
rect 29 100 229 138
rect 287 138 370 155
rect 404 155 453 172
rect 579 172 711 188
rect 579 155 628 172
rect 404 138 487 155
rect 287 100 487 138
rect 545 138 628 155
rect 662 155 711 172
rect 837 172 969 188
rect 837 155 886 172
rect 662 138 745 155
rect 545 100 745 138
rect 803 138 886 155
rect 920 155 969 172
rect 1095 172 1227 188
rect 1095 155 1144 172
rect 920 138 1003 155
rect 803 100 1003 138
rect 1061 138 1144 155
rect 1178 155 1227 172
rect 1178 138 1261 155
rect 1061 100 1261 138
rect -1261 -138 -1061 -100
rect -1261 -155 -1178 -138
rect -1227 -172 -1178 -155
rect -1144 -155 -1061 -138
rect -1003 -138 -803 -100
rect -1003 -155 -920 -138
rect -1144 -172 -1095 -155
rect -1227 -188 -1095 -172
rect -969 -172 -920 -155
rect -886 -155 -803 -138
rect -745 -138 -545 -100
rect -745 -155 -662 -138
rect -886 -172 -837 -155
rect -969 -188 -837 -172
rect -711 -172 -662 -155
rect -628 -155 -545 -138
rect -487 -138 -287 -100
rect -487 -155 -404 -138
rect -628 -172 -579 -155
rect -711 -188 -579 -172
rect -453 -172 -404 -155
rect -370 -155 -287 -138
rect -229 -138 -29 -100
rect -229 -155 -146 -138
rect -370 -172 -321 -155
rect -453 -188 -321 -172
rect -195 -172 -146 -155
rect -112 -155 -29 -138
rect 29 -138 229 -100
rect 29 -155 112 -138
rect -112 -172 -63 -155
rect -195 -188 -63 -172
rect 63 -172 112 -155
rect 146 -155 229 -138
rect 287 -138 487 -100
rect 287 -155 370 -138
rect 146 -172 195 -155
rect 63 -188 195 -172
rect 321 -172 370 -155
rect 404 -155 487 -138
rect 545 -138 745 -100
rect 545 -155 628 -138
rect 404 -172 453 -155
rect 321 -188 453 -172
rect 579 -172 628 -155
rect 662 -155 745 -138
rect 803 -138 1003 -100
rect 803 -155 886 -138
rect 662 -172 711 -155
rect 579 -188 711 -172
rect 837 -172 886 -155
rect 920 -155 1003 -138
rect 1061 -138 1261 -100
rect 1061 -155 1144 -138
rect 920 -172 969 -155
rect 837 -188 969 -172
rect 1095 -172 1144 -155
rect 1178 -155 1261 -138
rect 1178 -172 1227 -155
rect 1095 -188 1227 -172
<< polycont >>
rect -1178 138 -1144 172
rect -920 138 -886 172
rect -662 138 -628 172
rect -404 138 -370 172
rect -146 138 -112 172
rect 112 138 146 172
rect 370 138 404 172
rect 628 138 662 172
rect 886 138 920 172
rect 1144 138 1178 172
rect -1178 -172 -1144 -138
rect -920 -172 -886 -138
rect -662 -172 -628 -138
rect -404 -172 -370 -138
rect -146 -172 -112 -138
rect 112 -172 146 -138
rect 370 -172 404 -138
rect 628 -172 662 -138
rect 886 -172 920 -138
rect 1144 -172 1178 -138
<< locali >>
rect -1227 138 -1178 172
rect -1144 138 -1095 172
rect -969 138 -920 172
rect -886 138 -837 172
rect -711 138 -662 172
rect -628 138 -579 172
rect -453 138 -404 172
rect -370 138 -321 172
rect -195 138 -146 172
rect -112 138 -63 172
rect 63 138 112 172
rect 146 138 195 172
rect 321 138 370 172
rect 404 138 453 172
rect 579 138 628 172
rect 662 138 711 172
rect 837 138 886 172
rect 920 138 969 172
rect 1095 138 1144 172
rect 1178 138 1227 172
rect -1307 85 -1273 104
rect -1307 17 -1273 19
rect -1307 -19 -1273 -17
rect -1307 -104 -1273 -85
rect -1049 85 -1015 104
rect -1049 17 -1015 19
rect -1049 -19 -1015 -17
rect -1049 -104 -1015 -85
rect -791 85 -757 104
rect -791 17 -757 19
rect -791 -19 -757 -17
rect -791 -104 -757 -85
rect -533 85 -499 104
rect -533 17 -499 19
rect -533 -19 -499 -17
rect -533 -104 -499 -85
rect -275 85 -241 104
rect -275 17 -241 19
rect -275 -19 -241 -17
rect -275 -104 -241 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 241 85 275 104
rect 241 17 275 19
rect 241 -19 275 -17
rect 241 -104 275 -85
rect 499 85 533 104
rect 499 17 533 19
rect 499 -19 533 -17
rect 499 -104 533 -85
rect 757 85 791 104
rect 757 17 791 19
rect 757 -19 791 -17
rect 757 -104 791 -85
rect 1015 85 1049 104
rect 1015 17 1049 19
rect 1015 -19 1049 -17
rect 1015 -104 1049 -85
rect 1273 85 1307 104
rect 1273 17 1307 19
rect 1273 -19 1307 -17
rect 1273 -104 1307 -85
rect -1227 -172 -1178 -138
rect -1144 -172 -1095 -138
rect -969 -172 -920 -138
rect -886 -172 -837 -138
rect -711 -172 -662 -138
rect -628 -172 -579 -138
rect -453 -172 -404 -138
rect -370 -172 -321 -138
rect -195 -172 -146 -138
rect -112 -172 -63 -138
rect 63 -172 112 -138
rect 146 -172 195 -138
rect 321 -172 370 -138
rect 404 -172 453 -138
rect 579 -172 628 -138
rect 662 -172 711 -138
rect 837 -172 886 -138
rect 920 -172 969 -138
rect 1095 -172 1144 -138
rect 1178 -172 1227 -138
<< viali >>
rect -1178 138 -1144 172
rect -920 138 -886 172
rect -662 138 -628 172
rect -404 138 -370 172
rect -146 138 -112 172
rect 112 138 146 172
rect 370 138 404 172
rect 628 138 662 172
rect 886 138 920 172
rect 1144 138 1178 172
rect -1307 51 -1273 53
rect -1307 19 -1273 51
rect -1307 -51 -1273 -19
rect -1307 -53 -1273 -51
rect -1049 51 -1015 53
rect -1049 19 -1015 51
rect -1049 -51 -1015 -19
rect -1049 -53 -1015 -51
rect -791 51 -757 53
rect -791 19 -757 51
rect -791 -51 -757 -19
rect -791 -53 -757 -51
rect -533 51 -499 53
rect -533 19 -499 51
rect -533 -51 -499 -19
rect -533 -53 -499 -51
rect -275 51 -241 53
rect -275 19 -241 51
rect -275 -51 -241 -19
rect -275 -53 -241 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 241 51 275 53
rect 241 19 275 51
rect 241 -51 275 -19
rect 241 -53 275 -51
rect 499 51 533 53
rect 499 19 533 51
rect 499 -51 533 -19
rect 499 -53 533 -51
rect 757 51 791 53
rect 757 19 791 51
rect 757 -51 791 -19
rect 757 -53 791 -51
rect 1015 51 1049 53
rect 1015 19 1049 51
rect 1015 -51 1049 -19
rect 1015 -53 1049 -51
rect 1273 51 1307 53
rect 1273 19 1307 51
rect 1273 -51 1307 -19
rect 1273 -53 1307 -51
rect -1178 -172 -1144 -138
rect -920 -172 -886 -138
rect -662 -172 -628 -138
rect -404 -172 -370 -138
rect -146 -172 -112 -138
rect 112 -172 146 -138
rect 370 -172 404 -138
rect 628 -172 662 -138
rect 886 -172 920 -138
rect 1144 -172 1178 -138
<< metal1 >>
rect -1215 172 -1107 178
rect -1215 138 -1178 172
rect -1144 138 -1107 172
rect -1215 132 -1107 138
rect -957 172 -849 178
rect -957 138 -920 172
rect -886 138 -849 172
rect -957 132 -849 138
rect -699 172 -591 178
rect -699 138 -662 172
rect -628 138 -591 172
rect -699 132 -591 138
rect -441 172 -333 178
rect -441 138 -404 172
rect -370 138 -333 172
rect -441 132 -333 138
rect -183 172 -75 178
rect -183 138 -146 172
rect -112 138 -75 172
rect -183 132 -75 138
rect 75 172 183 178
rect 75 138 112 172
rect 146 138 183 172
rect 75 132 183 138
rect 333 172 441 178
rect 333 138 370 172
rect 404 138 441 172
rect 333 132 441 138
rect 591 172 699 178
rect 591 138 628 172
rect 662 138 699 172
rect 591 132 699 138
rect 849 172 957 178
rect 849 138 886 172
rect 920 138 957 172
rect 849 132 957 138
rect 1107 172 1215 178
rect 1107 138 1144 172
rect 1178 138 1215 172
rect 1107 132 1215 138
rect -1313 53 -1267 100
rect -1313 19 -1307 53
rect -1273 19 -1267 53
rect -1313 -19 -1267 19
rect -1313 -53 -1307 -19
rect -1273 -53 -1267 -19
rect -1313 -100 -1267 -53
rect -1055 53 -1009 100
rect -1055 19 -1049 53
rect -1015 19 -1009 53
rect -1055 -19 -1009 19
rect -1055 -53 -1049 -19
rect -1015 -53 -1009 -19
rect -1055 -100 -1009 -53
rect -797 53 -751 100
rect -797 19 -791 53
rect -757 19 -751 53
rect -797 -19 -751 19
rect -797 -53 -791 -19
rect -757 -53 -751 -19
rect -797 -100 -751 -53
rect -539 53 -493 100
rect -539 19 -533 53
rect -499 19 -493 53
rect -539 -19 -493 19
rect -539 -53 -533 -19
rect -499 -53 -493 -19
rect -539 -100 -493 -53
rect -281 53 -235 100
rect -281 19 -275 53
rect -241 19 -235 53
rect -281 -19 -235 19
rect -281 -53 -275 -19
rect -241 -53 -235 -19
rect -281 -100 -235 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 235 53 281 100
rect 235 19 241 53
rect 275 19 281 53
rect 235 -19 281 19
rect 235 -53 241 -19
rect 275 -53 281 -19
rect 235 -100 281 -53
rect 493 53 539 100
rect 493 19 499 53
rect 533 19 539 53
rect 493 -19 539 19
rect 493 -53 499 -19
rect 533 -53 539 -19
rect 493 -100 539 -53
rect 751 53 797 100
rect 751 19 757 53
rect 791 19 797 53
rect 751 -19 797 19
rect 751 -53 757 -19
rect 791 -53 797 -19
rect 751 -100 797 -53
rect 1009 53 1055 100
rect 1009 19 1015 53
rect 1049 19 1055 53
rect 1009 -19 1055 19
rect 1009 -53 1015 -19
rect 1049 -53 1055 -19
rect 1009 -100 1055 -53
rect 1267 53 1313 100
rect 1267 19 1273 53
rect 1307 19 1313 53
rect 1267 -19 1313 19
rect 1267 -53 1273 -19
rect 1307 -53 1313 -19
rect 1267 -100 1313 -53
rect -1215 -138 -1107 -132
rect -1215 -172 -1178 -138
rect -1144 -172 -1107 -138
rect -1215 -178 -1107 -172
rect -957 -138 -849 -132
rect -957 -172 -920 -138
rect -886 -172 -849 -138
rect -957 -178 -849 -172
rect -699 -138 -591 -132
rect -699 -172 -662 -138
rect -628 -172 -591 -138
rect -699 -178 -591 -172
rect -441 -138 -333 -132
rect -441 -172 -404 -138
rect -370 -172 -333 -138
rect -441 -178 -333 -172
rect -183 -138 -75 -132
rect -183 -172 -146 -138
rect -112 -172 -75 -138
rect -183 -178 -75 -172
rect 75 -138 183 -132
rect 75 -172 112 -138
rect 146 -172 183 -138
rect 75 -178 183 -172
rect 333 -138 441 -132
rect 333 -172 370 -138
rect 404 -172 441 -138
rect 333 -178 441 -172
rect 591 -138 699 -132
rect 591 -172 628 -138
rect 662 -172 699 -138
rect 591 -178 699 -172
rect 849 -138 957 -132
rect 849 -172 886 -138
rect 920 -172 957 -138
rect 849 -178 957 -172
rect 1107 -138 1215 -132
rect 1107 -172 1144 -138
rect 1178 -172 1215 -138
rect 1107 -178 1215 -172
<< end >>
