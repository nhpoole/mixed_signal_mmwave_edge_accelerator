magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -2689 -1548 2689 1548
<< pwell >>
rect -1429 -226 1429 226
<< nmos >>
rect -1345 -200 -945 200
rect -887 -200 -487 200
rect -429 -200 -29 200
rect 29 -200 429 200
rect 487 -200 887 200
rect 945 -200 1345 200
<< ndiff >>
rect -1403 187 -1345 200
rect -1403 153 -1391 187
rect -1357 153 -1345 187
rect -1403 119 -1345 153
rect -1403 85 -1391 119
rect -1357 85 -1345 119
rect -1403 51 -1345 85
rect -1403 17 -1391 51
rect -1357 17 -1345 51
rect -1403 -17 -1345 17
rect -1403 -51 -1391 -17
rect -1357 -51 -1345 -17
rect -1403 -85 -1345 -51
rect -1403 -119 -1391 -85
rect -1357 -119 -1345 -85
rect -1403 -153 -1345 -119
rect -1403 -187 -1391 -153
rect -1357 -187 -1345 -153
rect -1403 -200 -1345 -187
rect -945 187 -887 200
rect -945 153 -933 187
rect -899 153 -887 187
rect -945 119 -887 153
rect -945 85 -933 119
rect -899 85 -887 119
rect -945 51 -887 85
rect -945 17 -933 51
rect -899 17 -887 51
rect -945 -17 -887 17
rect -945 -51 -933 -17
rect -899 -51 -887 -17
rect -945 -85 -887 -51
rect -945 -119 -933 -85
rect -899 -119 -887 -85
rect -945 -153 -887 -119
rect -945 -187 -933 -153
rect -899 -187 -887 -153
rect -945 -200 -887 -187
rect -487 187 -429 200
rect -487 153 -475 187
rect -441 153 -429 187
rect -487 119 -429 153
rect -487 85 -475 119
rect -441 85 -429 119
rect -487 51 -429 85
rect -487 17 -475 51
rect -441 17 -429 51
rect -487 -17 -429 17
rect -487 -51 -475 -17
rect -441 -51 -429 -17
rect -487 -85 -429 -51
rect -487 -119 -475 -85
rect -441 -119 -429 -85
rect -487 -153 -429 -119
rect -487 -187 -475 -153
rect -441 -187 -429 -153
rect -487 -200 -429 -187
rect -29 187 29 200
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -200 29 -187
rect 429 187 487 200
rect 429 153 441 187
rect 475 153 487 187
rect 429 119 487 153
rect 429 85 441 119
rect 475 85 487 119
rect 429 51 487 85
rect 429 17 441 51
rect 475 17 487 51
rect 429 -17 487 17
rect 429 -51 441 -17
rect 475 -51 487 -17
rect 429 -85 487 -51
rect 429 -119 441 -85
rect 475 -119 487 -85
rect 429 -153 487 -119
rect 429 -187 441 -153
rect 475 -187 487 -153
rect 429 -200 487 -187
rect 887 187 945 200
rect 887 153 899 187
rect 933 153 945 187
rect 887 119 945 153
rect 887 85 899 119
rect 933 85 945 119
rect 887 51 945 85
rect 887 17 899 51
rect 933 17 945 51
rect 887 -17 945 17
rect 887 -51 899 -17
rect 933 -51 945 -17
rect 887 -85 945 -51
rect 887 -119 899 -85
rect 933 -119 945 -85
rect 887 -153 945 -119
rect 887 -187 899 -153
rect 933 -187 945 -153
rect 887 -200 945 -187
rect 1345 187 1403 200
rect 1345 153 1357 187
rect 1391 153 1403 187
rect 1345 119 1403 153
rect 1345 85 1357 119
rect 1391 85 1403 119
rect 1345 51 1403 85
rect 1345 17 1357 51
rect 1391 17 1403 51
rect 1345 -17 1403 17
rect 1345 -51 1357 -17
rect 1391 -51 1403 -17
rect 1345 -85 1403 -51
rect 1345 -119 1357 -85
rect 1391 -119 1403 -85
rect 1345 -153 1403 -119
rect 1345 -187 1357 -153
rect 1391 -187 1403 -153
rect 1345 -200 1403 -187
<< ndiffc >>
rect -1391 153 -1357 187
rect -1391 85 -1357 119
rect -1391 17 -1357 51
rect -1391 -51 -1357 -17
rect -1391 -119 -1357 -85
rect -1391 -187 -1357 -153
rect -933 153 -899 187
rect -933 85 -899 119
rect -933 17 -899 51
rect -933 -51 -899 -17
rect -933 -119 -899 -85
rect -933 -187 -899 -153
rect -475 153 -441 187
rect -475 85 -441 119
rect -475 17 -441 51
rect -475 -51 -441 -17
rect -475 -119 -441 -85
rect -475 -187 -441 -153
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect 441 153 475 187
rect 441 85 475 119
rect 441 17 475 51
rect 441 -51 475 -17
rect 441 -119 475 -85
rect 441 -187 475 -153
rect 899 153 933 187
rect 899 85 933 119
rect 899 17 933 51
rect 899 -51 933 -17
rect 899 -119 933 -85
rect 899 -187 933 -153
rect 1357 153 1391 187
rect 1357 85 1391 119
rect 1357 17 1391 51
rect 1357 -51 1391 -17
rect 1357 -119 1391 -85
rect 1357 -187 1391 -153
<< poly >>
rect -1271 272 -1019 288
rect -1271 255 -1230 272
rect -1345 238 -1230 255
rect -1196 238 -1162 272
rect -1128 238 -1094 272
rect -1060 255 -1019 272
rect -813 272 -561 288
rect -813 255 -772 272
rect -1060 238 -945 255
rect -1345 200 -945 238
rect -887 238 -772 255
rect -738 238 -704 272
rect -670 238 -636 272
rect -602 255 -561 272
rect -355 272 -103 288
rect -355 255 -314 272
rect -602 238 -487 255
rect -887 200 -487 238
rect -429 238 -314 255
rect -280 238 -246 272
rect -212 238 -178 272
rect -144 255 -103 272
rect 103 272 355 288
rect 103 255 144 272
rect -144 238 -29 255
rect -429 200 -29 238
rect 29 238 144 255
rect 178 238 212 272
rect 246 238 280 272
rect 314 255 355 272
rect 561 272 813 288
rect 561 255 602 272
rect 314 238 429 255
rect 29 200 429 238
rect 487 238 602 255
rect 636 238 670 272
rect 704 238 738 272
rect 772 255 813 272
rect 1019 272 1271 288
rect 1019 255 1060 272
rect 772 238 887 255
rect 487 200 887 238
rect 945 238 1060 255
rect 1094 238 1128 272
rect 1162 238 1196 272
rect 1230 255 1271 272
rect 1230 238 1345 255
rect 945 200 1345 238
rect -1345 -238 -945 -200
rect -1345 -255 -1230 -238
rect -1271 -272 -1230 -255
rect -1196 -272 -1162 -238
rect -1128 -272 -1094 -238
rect -1060 -255 -945 -238
rect -887 -238 -487 -200
rect -887 -255 -772 -238
rect -1060 -272 -1019 -255
rect -1271 -288 -1019 -272
rect -813 -272 -772 -255
rect -738 -272 -704 -238
rect -670 -272 -636 -238
rect -602 -255 -487 -238
rect -429 -238 -29 -200
rect -429 -255 -314 -238
rect -602 -272 -561 -255
rect -813 -288 -561 -272
rect -355 -272 -314 -255
rect -280 -272 -246 -238
rect -212 -272 -178 -238
rect -144 -255 -29 -238
rect 29 -238 429 -200
rect 29 -255 144 -238
rect -144 -272 -103 -255
rect -355 -288 -103 -272
rect 103 -272 144 -255
rect 178 -272 212 -238
rect 246 -272 280 -238
rect 314 -255 429 -238
rect 487 -238 887 -200
rect 487 -255 602 -238
rect 314 -272 355 -255
rect 103 -288 355 -272
rect 561 -272 602 -255
rect 636 -272 670 -238
rect 704 -272 738 -238
rect 772 -255 887 -238
rect 945 -238 1345 -200
rect 945 -255 1060 -238
rect 772 -272 813 -255
rect 561 -288 813 -272
rect 1019 -272 1060 -255
rect 1094 -272 1128 -238
rect 1162 -272 1196 -238
rect 1230 -255 1345 -238
rect 1230 -272 1271 -255
rect 1019 -288 1271 -272
<< polycont >>
rect -1230 238 -1196 272
rect -1162 238 -1128 272
rect -1094 238 -1060 272
rect -772 238 -738 272
rect -704 238 -670 272
rect -636 238 -602 272
rect -314 238 -280 272
rect -246 238 -212 272
rect -178 238 -144 272
rect 144 238 178 272
rect 212 238 246 272
rect 280 238 314 272
rect 602 238 636 272
rect 670 238 704 272
rect 738 238 772 272
rect 1060 238 1094 272
rect 1128 238 1162 272
rect 1196 238 1230 272
rect -1230 -272 -1196 -238
rect -1162 -272 -1128 -238
rect -1094 -272 -1060 -238
rect -772 -272 -738 -238
rect -704 -272 -670 -238
rect -636 -272 -602 -238
rect -314 -272 -280 -238
rect -246 -272 -212 -238
rect -178 -272 -144 -238
rect 144 -272 178 -238
rect 212 -272 246 -238
rect 280 -272 314 -238
rect 602 -272 636 -238
rect 670 -272 704 -238
rect 738 -272 772 -238
rect 1060 -272 1094 -238
rect 1128 -272 1162 -238
rect 1196 -272 1230 -238
<< locali >>
rect -1271 238 -1234 272
rect -1196 238 -1162 272
rect -1128 238 -1094 272
rect -1056 238 -1019 272
rect -813 238 -776 272
rect -738 238 -704 272
rect -670 238 -636 272
rect -598 238 -561 272
rect -355 238 -318 272
rect -280 238 -246 272
rect -212 238 -178 272
rect -140 238 -103 272
rect 103 238 140 272
rect 178 238 212 272
rect 246 238 280 272
rect 318 238 355 272
rect 561 238 598 272
rect 636 238 670 272
rect 704 238 738 272
rect 776 238 813 272
rect 1019 238 1056 272
rect 1094 238 1128 272
rect 1162 238 1196 272
rect 1234 238 1271 272
rect -1391 187 -1357 204
rect -1391 119 -1357 127
rect -1391 51 -1357 55
rect -1391 -55 -1357 -51
rect -1391 -127 -1357 -119
rect -1391 -204 -1357 -187
rect -933 187 -899 204
rect -933 119 -899 127
rect -933 51 -899 55
rect -933 -55 -899 -51
rect -933 -127 -899 -119
rect -933 -204 -899 -187
rect -475 187 -441 204
rect -475 119 -441 127
rect -475 51 -441 55
rect -475 -55 -441 -51
rect -475 -127 -441 -119
rect -475 -204 -441 -187
rect -17 187 17 204
rect -17 119 17 127
rect -17 51 17 55
rect -17 -55 17 -51
rect -17 -127 17 -119
rect -17 -204 17 -187
rect 441 187 475 204
rect 441 119 475 127
rect 441 51 475 55
rect 441 -55 475 -51
rect 441 -127 475 -119
rect 441 -204 475 -187
rect 899 187 933 204
rect 899 119 933 127
rect 899 51 933 55
rect 899 -55 933 -51
rect 899 -127 933 -119
rect 899 -204 933 -187
rect 1357 187 1391 204
rect 1357 119 1391 127
rect 1357 51 1391 55
rect 1357 -55 1391 -51
rect 1357 -127 1391 -119
rect 1357 -204 1391 -187
rect -1271 -272 -1234 -238
rect -1196 -272 -1162 -238
rect -1128 -272 -1094 -238
rect -1056 -272 -1019 -238
rect -813 -272 -776 -238
rect -738 -272 -704 -238
rect -670 -272 -636 -238
rect -598 -272 -561 -238
rect -355 -272 -318 -238
rect -280 -272 -246 -238
rect -212 -272 -178 -238
rect -140 -272 -103 -238
rect 103 -272 140 -238
rect 178 -272 212 -238
rect 246 -272 280 -238
rect 318 -272 355 -238
rect 561 -272 598 -238
rect 636 -272 670 -238
rect 704 -272 738 -238
rect 776 -272 813 -238
rect 1019 -272 1056 -238
rect 1094 -272 1128 -238
rect 1162 -272 1196 -238
rect 1234 -272 1271 -238
<< viali >>
rect -1234 238 -1230 272
rect -1230 238 -1200 272
rect -1162 238 -1128 272
rect -1090 238 -1060 272
rect -1060 238 -1056 272
rect -776 238 -772 272
rect -772 238 -742 272
rect -704 238 -670 272
rect -632 238 -602 272
rect -602 238 -598 272
rect -318 238 -314 272
rect -314 238 -284 272
rect -246 238 -212 272
rect -174 238 -144 272
rect -144 238 -140 272
rect 140 238 144 272
rect 144 238 174 272
rect 212 238 246 272
rect 284 238 314 272
rect 314 238 318 272
rect 598 238 602 272
rect 602 238 632 272
rect 670 238 704 272
rect 742 238 772 272
rect 772 238 776 272
rect 1056 238 1060 272
rect 1060 238 1090 272
rect 1128 238 1162 272
rect 1200 238 1230 272
rect 1230 238 1234 272
rect -1391 153 -1357 161
rect -1391 127 -1357 153
rect -1391 85 -1357 89
rect -1391 55 -1357 85
rect -1391 -17 -1357 17
rect -1391 -85 -1357 -55
rect -1391 -89 -1357 -85
rect -1391 -153 -1357 -127
rect -1391 -161 -1357 -153
rect -933 153 -899 161
rect -933 127 -899 153
rect -933 85 -899 89
rect -933 55 -899 85
rect -933 -17 -899 17
rect -933 -85 -899 -55
rect -933 -89 -899 -85
rect -933 -153 -899 -127
rect -933 -161 -899 -153
rect -475 153 -441 161
rect -475 127 -441 153
rect -475 85 -441 89
rect -475 55 -441 85
rect -475 -17 -441 17
rect -475 -85 -441 -55
rect -475 -89 -441 -85
rect -475 -153 -441 -127
rect -475 -161 -441 -153
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect 441 153 475 161
rect 441 127 475 153
rect 441 85 475 89
rect 441 55 475 85
rect 441 -17 475 17
rect 441 -85 475 -55
rect 441 -89 475 -85
rect 441 -153 475 -127
rect 441 -161 475 -153
rect 899 153 933 161
rect 899 127 933 153
rect 899 85 933 89
rect 899 55 933 85
rect 899 -17 933 17
rect 899 -85 933 -55
rect 899 -89 933 -85
rect 899 -153 933 -127
rect 899 -161 933 -153
rect 1357 153 1391 161
rect 1357 127 1391 153
rect 1357 85 1391 89
rect 1357 55 1391 85
rect 1357 -17 1391 17
rect 1357 -85 1391 -55
rect 1357 -89 1391 -85
rect 1357 -153 1391 -127
rect 1357 -161 1391 -153
rect -1234 -272 -1230 -238
rect -1230 -272 -1200 -238
rect -1162 -272 -1128 -238
rect -1090 -272 -1060 -238
rect -1060 -272 -1056 -238
rect -776 -272 -772 -238
rect -772 -272 -742 -238
rect -704 -272 -670 -238
rect -632 -272 -602 -238
rect -602 -272 -598 -238
rect -318 -272 -314 -238
rect -314 -272 -284 -238
rect -246 -272 -212 -238
rect -174 -272 -144 -238
rect -144 -272 -140 -238
rect 140 -272 144 -238
rect 144 -272 174 -238
rect 212 -272 246 -238
rect 284 -272 314 -238
rect 314 -272 318 -238
rect 598 -272 602 -238
rect 602 -272 632 -238
rect 670 -272 704 -238
rect 742 -272 772 -238
rect 772 -272 776 -238
rect 1056 -272 1060 -238
rect 1060 -272 1090 -238
rect 1128 -272 1162 -238
rect 1200 -272 1230 -238
rect 1230 -272 1234 -238
<< metal1 >>
rect -1249 272 -1041 278
rect -1249 238 -1234 272
rect -1200 238 -1162 272
rect -1128 238 -1090 272
rect -1056 238 -1041 272
rect -1249 232 -1041 238
rect -791 272 -583 278
rect -791 238 -776 272
rect -742 238 -704 272
rect -670 238 -632 272
rect -598 238 -583 272
rect -791 232 -583 238
rect -333 272 -125 278
rect -333 238 -318 272
rect -284 238 -246 272
rect -212 238 -174 272
rect -140 238 -125 272
rect -333 232 -125 238
rect 125 272 333 278
rect 125 238 140 272
rect 174 238 212 272
rect 246 238 284 272
rect 318 238 333 272
rect 125 232 333 238
rect 583 272 791 278
rect 583 238 598 272
rect 632 238 670 272
rect 704 238 742 272
rect 776 238 791 272
rect 583 232 791 238
rect 1041 272 1249 278
rect 1041 238 1056 272
rect 1090 238 1128 272
rect 1162 238 1200 272
rect 1234 238 1249 272
rect 1041 232 1249 238
rect -1397 161 -1351 200
rect -1397 127 -1391 161
rect -1357 127 -1351 161
rect -1397 89 -1351 127
rect -1397 55 -1391 89
rect -1357 55 -1351 89
rect -1397 17 -1351 55
rect -1397 -17 -1391 17
rect -1357 -17 -1351 17
rect -1397 -55 -1351 -17
rect -1397 -89 -1391 -55
rect -1357 -89 -1351 -55
rect -1397 -127 -1351 -89
rect -1397 -161 -1391 -127
rect -1357 -161 -1351 -127
rect -1397 -200 -1351 -161
rect -939 161 -893 200
rect -939 127 -933 161
rect -899 127 -893 161
rect -939 89 -893 127
rect -939 55 -933 89
rect -899 55 -893 89
rect -939 17 -893 55
rect -939 -17 -933 17
rect -899 -17 -893 17
rect -939 -55 -893 -17
rect -939 -89 -933 -55
rect -899 -89 -893 -55
rect -939 -127 -893 -89
rect -939 -161 -933 -127
rect -899 -161 -893 -127
rect -939 -200 -893 -161
rect -481 161 -435 200
rect -481 127 -475 161
rect -441 127 -435 161
rect -481 89 -435 127
rect -481 55 -475 89
rect -441 55 -435 89
rect -481 17 -435 55
rect -481 -17 -475 17
rect -441 -17 -435 17
rect -481 -55 -435 -17
rect -481 -89 -475 -55
rect -441 -89 -435 -55
rect -481 -127 -435 -89
rect -481 -161 -475 -127
rect -441 -161 -435 -127
rect -481 -200 -435 -161
rect -23 161 23 200
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -200 23 -161
rect 435 161 481 200
rect 435 127 441 161
rect 475 127 481 161
rect 435 89 481 127
rect 435 55 441 89
rect 475 55 481 89
rect 435 17 481 55
rect 435 -17 441 17
rect 475 -17 481 17
rect 435 -55 481 -17
rect 435 -89 441 -55
rect 475 -89 481 -55
rect 435 -127 481 -89
rect 435 -161 441 -127
rect 475 -161 481 -127
rect 435 -200 481 -161
rect 893 161 939 200
rect 893 127 899 161
rect 933 127 939 161
rect 893 89 939 127
rect 893 55 899 89
rect 933 55 939 89
rect 893 17 939 55
rect 893 -17 899 17
rect 933 -17 939 17
rect 893 -55 939 -17
rect 893 -89 899 -55
rect 933 -89 939 -55
rect 893 -127 939 -89
rect 893 -161 899 -127
rect 933 -161 939 -127
rect 893 -200 939 -161
rect 1351 161 1397 200
rect 1351 127 1357 161
rect 1391 127 1397 161
rect 1351 89 1397 127
rect 1351 55 1357 89
rect 1391 55 1397 89
rect 1351 17 1397 55
rect 1351 -17 1357 17
rect 1391 -17 1397 17
rect 1351 -55 1397 -17
rect 1351 -89 1357 -55
rect 1391 -89 1397 -55
rect 1351 -127 1397 -89
rect 1351 -161 1357 -127
rect 1391 -161 1397 -127
rect 1351 -200 1397 -161
rect -1249 -238 -1041 -232
rect -1249 -272 -1234 -238
rect -1200 -272 -1162 -238
rect -1128 -272 -1090 -238
rect -1056 -272 -1041 -238
rect -1249 -278 -1041 -272
rect -791 -238 -583 -232
rect -791 -272 -776 -238
rect -742 -272 -704 -238
rect -670 -272 -632 -238
rect -598 -272 -583 -238
rect -791 -278 -583 -272
rect -333 -238 -125 -232
rect -333 -272 -318 -238
rect -284 -272 -246 -238
rect -212 -272 -174 -238
rect -140 -272 -125 -238
rect -333 -278 -125 -272
rect 125 -238 333 -232
rect 125 -272 140 -238
rect 174 -272 212 -238
rect 246 -272 284 -238
rect 318 -272 333 -238
rect 125 -278 333 -272
rect 583 -238 791 -232
rect 583 -272 598 -238
rect 632 -272 670 -238
rect 704 -272 742 -238
rect 776 -272 791 -238
rect 583 -278 791 -272
rect 1041 -238 1249 -232
rect 1041 -272 1056 -238
rect 1090 -272 1128 -238
rect 1162 -272 1200 -238
rect 1234 -272 1249 -238
rect 1041 -278 1249 -272
<< end >>
