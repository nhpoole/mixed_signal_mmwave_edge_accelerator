magic
tech sky130A
magscale 1 2
timestamp 1625985445
<< nwell >>
rect -12082 15478 -10232 16318
rect -8617 15502 -7946 15800
rect -8617 15479 -8084 15502
rect -7962 15479 -7946 15502
<< pwell >>
rect -8558 15406 -8084 15421
rect -11841 14864 -10108 15384
rect -8558 15239 -7981 15406
rect -11841 14764 -10196 14864
<< viali >>
rect -8052 15430 -8004 15478
rect -7950 15434 -7902 15482
<< metal1 >>
rect 47792 27680 48000 27710
rect -1414 27642 -1354 27648
rect -8742 16408 -8682 16414
rect -1414 16408 -1354 27582
rect 47792 27564 47824 27680
rect 47022 25478 47376 25538
rect 47792 25514 48000 27564
rect 48306 27680 48488 27710
rect 48462 27564 48488 27680
rect 48306 25497 48488 27564
rect 47022 23538 47082 25478
rect 47244 23874 47250 23934
rect 47310 23874 47316 23934
rect 47022 23478 47802 23538
rect 48682 23478 50478 23538
rect 46972 21860 46978 21920
rect 47038 21860 47310 21920
rect -11462 16348 -10092 16408
rect -1420 16348 -1414 16408
rect -1354 16348 -1348 16408
rect -8742 16342 -8682 16348
rect -8340 15714 -8100 15810
rect -8299 15478 -7992 15484
rect -8299 15430 -8052 15478
rect -8004 15430 -7992 15478
rect -8299 15424 -7992 15430
rect -7962 15482 -7734 15488
rect -7962 15434 -7950 15482
rect -7902 15434 -7734 15482
rect -7962 15428 -7734 15434
rect -8340 15170 -8100 15266
rect -12478 14956 -12418 15054
rect -12484 14896 -12478 14956
rect -12418 14896 -12412 14956
rect -9878 14952 -9818 15078
rect -9884 14892 -9878 14952
rect -9818 14892 -9812 14952
rect -10006 14837 -9946 14843
rect -10006 14771 -9946 14777
rect -10508 14712 -10502 14730
rect -8750 14712 -8690 14718
rect -11460 14652 -9402 14712
rect -8750 14646 -8690 14652
rect -1792 14712 -1732 14718
rect -1732 14652 -1294 14712
rect -1792 14646 -1732 14652
rect 48494 8574 48554 8578
rect 48494 8514 49142 8574
rect 50076 8546 50476 23478
rect 50938 9048 50944 9108
rect 51004 9048 51010 9108
rect 48358 7491 48364 7551
rect 48424 7491 48430 7551
rect 48364 6176 48424 7491
rect 48494 6610 48554 8514
rect 50944 7650 51004 9048
rect 50812 7590 51004 7650
rect 49766 6818 52704 6878
rect 48494 6550 48854 6610
rect 48358 6116 48364 6176
rect 48424 6116 48430 6176
rect 8274 5144 8280 5204
rect 8340 5144 8346 5204
rect 3944 4926 4244 4986
rect 8280 4788 8340 5144
rect 48494 4610 48554 6550
rect 50810 5626 51006 5686
rect 57932 4926 58226 4986
rect 49930 4854 52710 4914
rect 48494 4550 48994 4610
rect 48494 2520 48554 4550
rect 49960 2854 52704 2914
rect 48494 2462 49148 2520
rect 48498 2460 49148 2462
rect 50008 764 52706 824
<< via1 >>
rect -1414 27582 -1354 27642
rect 47824 27564 48000 27680
rect 48306 27564 48462 27680
rect 47250 23874 47310 23934
rect 46978 21860 47038 21920
rect -8742 16348 -8682 16408
rect -1414 16348 -1354 16408
rect -12478 14896 -12418 14956
rect -9878 14892 -9818 14952
rect -10006 14777 -9946 14837
rect -8750 14652 -8690 14712
rect -1792 14652 -1732 14712
rect 50944 9048 51004 9108
rect 48364 7491 48424 7551
rect 48364 6116 48424 6176
rect 8280 5144 8340 5204
<< metal2 >>
rect 47796 27680 48490 27702
rect -1414 27642 -1354 27651
rect -1420 27582 -1414 27642
rect -1354 27582 -1348 27642
rect -1414 27573 -1354 27582
rect 47796 27564 47824 27680
rect 48462 27564 48490 27680
rect 47796 27536 48490 27564
rect 48230 24604 48398 24664
rect 48458 24604 48467 24664
rect 47615 24455 47624 24515
rect 47684 24455 47782 24515
rect 47250 23934 47310 23940
rect 42781 23874 42790 23934
rect 42850 23874 47250 23934
rect 47250 23868 47310 23874
rect 38874 23861 38964 23866
rect 38870 23781 38879 23861
rect 38959 23781 38968 23861
rect 38874 23705 38964 23781
rect 38874 23615 41091 23705
rect 41001 23527 41091 23615
rect 41001 23428 41091 23437
rect 47867 22604 47876 22664
rect 47936 22604 48046 22664
rect 48514 22455 48656 22515
rect 48716 22455 48725 22515
rect 49519 22328 49579 24074
rect 46978 21920 47038 21926
rect 42791 21860 42800 21920
rect 42860 21860 46978 21920
rect 46978 21854 47038 21860
rect 40228 21414 40328 21423
rect 36254 21314 40228 21414
rect 11206 18913 11306 18918
rect 11202 18823 11211 18913
rect 11301 18823 11310 18913
rect -1414 16408 -1354 16414
rect -8748 16348 -8742 16408
rect -8682 16348 -1414 16408
rect -1414 16342 -1354 16348
rect 10953 16318 10962 16418
rect 11062 16318 11071 16418
rect -13295 15325 -13286 15385
rect -13226 15325 -12580 15385
rect -10629 15325 -10620 15385
rect -10560 15325 -10006 15385
rect -1933 15092 -1924 15152
rect -1864 15092 -1855 15152
rect -12478 14956 -12418 14962
rect -13467 14610 -13377 14614
rect -12478 14610 -12418 14896
rect -9878 14952 -9818 14958
rect -10838 14777 -10006 14837
rect -9946 14777 -9940 14837
rect -13472 14605 -12418 14610
rect -13472 14515 -13467 14605
rect -13377 14515 -12418 14605
rect -13472 14510 -12418 14515
rect -13467 14506 -13377 14510
rect -9878 13120 -9818 14892
rect -1924 14838 -1864 15092
rect 10962 14983 11062 16318
rect 11206 15882 11306 18823
rect 36254 16193 36354 21314
rect 40228 21305 40328 21314
rect 65088 18913 65188 18918
rect 65084 18823 65093 18913
rect 65183 18823 65192 18913
rect 43134 17841 43262 17846
rect 38968 17829 39076 17834
rect 38964 17731 38973 17829
rect 39071 17731 39080 17829
rect 38968 17668 39076 17731
rect 43130 17723 43139 17841
rect 43257 17723 43266 17841
rect 47326 17831 47436 17836
rect 47322 17731 47331 17831
rect 47431 17731 47440 17831
rect 43134 17694 43262 17723
rect 38968 17560 41102 17668
rect 43134 17566 45316 17694
rect 40994 17516 41102 17560
rect 40994 17399 41102 17408
rect 45188 17526 45316 17566
rect 47326 17669 47436 17731
rect 47326 17559 49393 17669
rect 45188 17389 45316 17398
rect 49283 17507 49393 17559
rect 49283 17388 49393 17397
rect 36250 16103 36259 16193
rect 36349 16103 36358 16193
rect 36254 16098 36354 16103
rect 11197 15782 11206 15882
rect 11306 15782 11315 15882
rect 10958 14893 10967 14983
rect 11057 14893 11066 14983
rect 10962 14888 11062 14893
rect -8360 14778 -1864 14838
rect 11206 14812 11306 15782
rect 11197 14712 11206 14812
rect 11306 14712 11315 14812
rect 65088 14738 65188 18823
rect -8756 14652 -8750 14712
rect -8690 14652 -1792 14712
rect -1732 14652 -1726 14712
rect 65079 14638 65088 14738
rect 65188 14638 65197 14738
rect 36456 13814 36556 13823
rect 39253 13814 39343 13818
rect 36556 13809 39348 13814
rect 36556 13719 39253 13809
rect 39343 13719 39348 13809
rect 36556 13714 39348 13719
rect 36456 13705 36556 13714
rect 39253 13710 39343 13714
rect -9878 13051 -9818 13060
rect 42994 11727 43130 11732
rect 38844 11711 38950 11716
rect 38840 11615 38849 11711
rect 38945 11615 38954 11711
rect 38844 11553 38950 11615
rect 42990 11597 42999 11727
rect 43125 11597 43134 11727
rect 42994 11590 43134 11597
rect 38844 11447 40991 11553
rect 42994 11454 45158 11590
rect 40885 11381 40991 11447
rect 45050 11392 45158 11454
rect 45050 11275 45158 11284
rect 40885 11266 40991 11275
rect -9960 11043 -9846 11048
rect -9964 10939 -9955 11043
rect -9851 10939 -9842 11043
rect -5826 11027 -5720 11032
rect -9960 10871 -9846 10939
rect -5830 10931 -5821 11027
rect -5725 10931 -5716 11027
rect -5826 10891 -5720 10931
rect -9960 10757 -8667 10871
rect -5826 10785 -4683 10891
rect -8781 10725 -8667 10757
rect -8781 10602 -8667 10611
rect -4789 10715 -4683 10785
rect -4789 10600 -4683 10609
rect 36060 9306 36160 9315
rect 39009 9306 39099 9310
rect 36056 9206 36060 9306
rect 36160 9301 39104 9306
rect 36160 9211 39009 9301
rect 39099 9211 39104 9301
rect 36160 9206 39104 9211
rect 36060 9197 36160 9206
rect 39009 9202 39099 9206
rect 35833 9132 35935 9136
rect 35828 9127 51026 9132
rect 35828 9025 35833 9127
rect 35935 9108 51026 9127
rect 35935 9048 50944 9108
rect 51004 9048 51026 9108
rect 35935 9025 51026 9048
rect 35828 9020 51026 9025
rect 35833 9016 35935 9020
rect 49704 7640 49822 7700
rect 49882 7640 49891 7700
rect 48364 7551 48424 7557
rect 48424 7491 49184 7551
rect 48364 7485 48424 7491
rect 11382 7198 11442 7207
rect 9888 7138 11382 7198
rect 62341 7138 62350 7198
rect 62410 7138 62660 7198
rect 11382 7129 11442 7138
rect 50834 6944 51160 7004
rect 45907 6098 45916 6198
rect 46016 6176 48434 6198
rect 46016 6116 48364 6176
rect 48424 6116 48434 6176
rect 46016 6098 48434 6116
rect 49297 5676 49306 5736
rect 49366 5676 49510 5736
rect 49931 5527 49940 5587
rect 50000 5527 50009 5587
rect 8280 5204 8340 5210
rect 8271 5144 8280 5204
rect 8340 5144 8349 5204
rect 8280 5138 8340 5144
rect 38910 4099 39020 4104
rect 38906 3999 38915 4099
rect 39015 3999 39024 4099
rect 43082 4097 43192 4102
rect 38910 3971 39020 3999
rect 43078 3997 43087 4097
rect 43187 3997 43196 4097
rect 38910 3861 40895 3971
rect -10820 3835 -10716 3840
rect -10824 3741 -10815 3835
rect -10721 3741 -10712 3835
rect -6742 3827 -6642 3832
rect -10820 3688 -10716 3741
rect -6746 3737 -6737 3827
rect -6647 3737 -6638 3827
rect 40785 3799 40895 3861
rect 43082 3957 43192 3997
rect 43082 3847 45171 3957
rect -10820 3584 -8906 3688
rect -6742 3686 -6642 3737
rect -6742 3586 -4536 3686
rect 40785 3680 40895 3689
rect 45061 3787 45171 3847
rect 45061 3668 45171 3677
rect 49293 3676 49302 3736
rect 49362 3676 49472 3736
rect -9010 3514 -8906 3584
rect -9010 3401 -8906 3410
rect -4636 3510 -4536 3586
rect 49940 3527 50082 3587
rect 50142 3527 50151 3587
rect -4636 3401 -4536 3410
rect 50945 3400 51005 5146
rect 8042 1566 9100 1626
rect 46079 1610 46088 1670
rect 46148 1610 46157 1670
rect 8042 582 8102 1566
rect 46088 1497 46148 1610
rect 49734 1586 49828 1646
rect 49888 1586 49897 1646
rect 51100 1596 51160 6944
rect 66017 4876 66026 4936
rect 66086 4876 66095 4936
rect 66026 3818 66086 4876
rect 65964 3758 66086 3818
rect 62153 2933 62243 2942
rect 62243 2860 62414 2920
rect 62153 2834 62243 2843
rect 50940 1536 51160 1596
rect 46088 1437 49196 1497
rect 8033 522 8042 582
rect 8102 522 8111 582
<< via2 >>
rect -1414 27582 -1354 27642
rect 47824 27564 48000 27680
rect 48000 27564 48306 27680
rect 48306 27564 48462 27680
rect 48398 24604 48458 24664
rect 47624 24455 47684 24515
rect 42790 23874 42850 23934
rect 38879 23781 38959 23861
rect 41001 23437 41091 23527
rect 47876 22604 47936 22664
rect 48656 22455 48716 22515
rect 42800 21860 42860 21920
rect 40228 21314 40328 21414
rect 11211 18823 11301 18913
rect 10962 16318 11062 16418
rect -13286 15325 -13226 15385
rect -10620 15325 -10560 15385
rect -1924 15092 -1864 15152
rect -13467 14515 -13377 14605
rect 65093 18823 65183 18913
rect 38973 17731 39071 17829
rect 43139 17723 43257 17841
rect 47331 17731 47431 17831
rect 40994 17408 41102 17516
rect 45188 17398 45316 17526
rect 49283 17397 49393 17507
rect 36259 16103 36349 16193
rect 11206 15782 11306 15882
rect 10967 14893 11057 14983
rect 11206 14712 11306 14812
rect 65088 14638 65188 14738
rect 36456 13714 36556 13814
rect 39253 13719 39343 13809
rect -9878 13060 -9818 13120
rect 38849 11615 38945 11711
rect 42999 11597 43125 11727
rect 40885 11275 40991 11381
rect 45050 11284 45158 11392
rect -9955 10939 -9851 11043
rect -5821 10931 -5725 11027
rect -8781 10611 -8667 10725
rect -4789 10609 -4683 10715
rect 36060 9206 36160 9306
rect 39009 9211 39099 9301
rect 35833 9025 35935 9127
rect 49822 7640 49882 7700
rect 11382 7138 11442 7198
rect 62350 7138 62410 7198
rect 45916 6098 46016 6198
rect 49306 5676 49366 5736
rect 49940 5527 50000 5587
rect 8280 5144 8340 5204
rect 38915 3999 39015 4099
rect 43087 3997 43187 4097
rect -10815 3741 -10721 3835
rect -6737 3737 -6647 3827
rect 40785 3689 40895 3799
rect 45061 3677 45171 3787
rect 49302 3676 49362 3736
rect -9010 3410 -8906 3514
rect 50082 3527 50142 3587
rect -4636 3410 -4536 3510
rect 46088 1610 46148 1670
rect 49828 1586 49888 1646
rect 66026 4876 66086 4936
rect 62153 2843 62243 2933
rect 8042 522 8102 582
<< metal3 >>
rect 47796 27680 48490 27702
rect -1436 27647 -1330 27668
rect -1436 27583 -1419 27647
rect -1349 27583 -1330 27647
rect -1436 27582 -1414 27583
rect -1354 27582 -1330 27583
rect -1436 27562 -1330 27582
rect 47796 27564 47824 27680
rect 48462 27564 48490 27680
rect 47796 27536 48490 27564
rect 38430 26568 38578 26574
rect 37160 26420 38430 26494
rect 41348 26568 41506 26574
rect 38578 26420 41348 26494
rect 37160 26410 41348 26420
rect 41506 26410 42865 26494
rect 37160 25893 42865 26410
rect 37160 24776 37761 25893
rect 41522 25880 42865 25893
rect 37044 24644 37050 24776
rect 37182 24644 37761 24776
rect 36462 23470 36468 23570
rect 36568 23470 36574 23570
rect 36468 20168 36568 23470
rect 37160 22676 37761 24644
rect 42251 24768 42865 25880
rect 42251 24632 42912 24768
rect 43048 24632 43054 24768
rect 48378 24664 51894 24688
rect 38874 23861 38964 23912
rect 40401 23870 40503 24099
rect 42251 23934 42865 24632
rect 48378 24604 48398 24664
rect 48458 24604 51894 24664
rect 48378 24588 51894 24604
rect 46576 24534 46676 24540
rect 46676 24515 47704 24534
rect 46676 24455 47624 24515
rect 47684 24455 47704 24515
rect 46676 24434 47704 24455
rect 46576 24428 46676 24434
rect 42251 23874 42790 23934
rect 42850 23874 42865 23934
rect 38874 23781 38879 23861
rect 38959 23781 38964 23861
rect 38874 23776 38964 23781
rect 40396 23770 40402 23870
rect 40502 23770 40508 23870
rect 40401 23769 40503 23770
rect 41563 23712 41661 23717
rect 42030 23712 42130 23718
rect 41562 23711 42030 23712
rect 41562 23613 41563 23711
rect 41661 23613 42030 23711
rect 41562 23612 42030 23613
rect 41563 23607 41661 23612
rect 42030 23606 42130 23612
rect 39492 23567 39592 23568
rect 39487 23469 39493 23567
rect 39591 23469 39597 23567
rect 40996 23527 41096 23532
rect 39492 23348 39592 23469
rect 40996 23437 41001 23527
rect 41091 23437 41096 23527
rect 40996 23432 41096 23437
rect 41001 23229 41091 23432
rect 37070 22556 37076 22676
rect 37196 22556 37761 22676
rect 37160 21038 37761 22556
rect 42251 22658 42865 23874
rect 46404 22664 47952 22684
rect 42251 22518 42864 22658
rect 43004 22518 43010 22658
rect 46404 22604 47876 22664
rect 47936 22604 47952 22664
rect 46404 22584 47952 22604
rect 40228 21419 40328 22002
rect 42251 21920 42865 22518
rect 42251 21860 42800 21920
rect 42860 21860 42865 21920
rect 40223 21414 40333 21419
rect 40223 21314 40228 21414
rect 40328 21314 40333 21414
rect 40223 21309 40333 21314
rect 42251 21038 42865 21860
rect 46404 21381 46504 22584
rect 48640 22515 49860 22532
rect 48640 22455 48656 22515
rect 48716 22455 49860 22515
rect 48640 22432 49860 22455
rect 49760 21700 49860 22432
rect 49760 21594 49860 21600
rect 46399 21283 46405 21381
rect 46503 21283 46509 21381
rect 46404 21282 46504 21283
rect 51794 21066 51894 24588
rect 52138 23614 52144 23714
rect 52244 23614 52250 23714
rect 37160 20828 51393 21038
rect 51788 20966 51794 21066
rect 51894 20966 51900 21066
rect 37160 20490 40646 20828
rect 37160 20437 38494 20490
rect 37279 20420 38494 20437
rect 36468 19925 36572 20168
rect 36467 19827 36473 19925
rect 36571 19827 36577 19925
rect 11036 18913 11638 18918
rect 11036 18823 11211 18913
rect 11301 18823 11638 18913
rect 11036 18818 11638 18823
rect 36468 17152 36572 19827
rect 37279 19649 37879 20420
rect 38672 20456 40646 20490
rect 40846 20490 51393 20828
rect 40846 20456 40894 20490
rect 38672 20420 40894 20456
rect 38494 20306 38672 20312
rect 41072 20420 43294 20490
rect 40894 20306 41072 20312
rect 43472 20420 45420 20490
rect 43294 20306 43472 20312
rect 45598 20420 47594 20490
rect 45420 20306 45598 20312
rect 47772 20420 49994 20490
rect 47594 20306 47772 20312
rect 50172 20420 51393 20490
rect 49994 20306 50172 20312
rect 39072 19826 39078 19926
rect 39178 19826 46764 19926
rect 37279 18790 37881 19649
rect 39682 19460 39782 19826
rect 42460 19512 42560 19826
rect 46664 19432 46764 19826
rect 37144 18582 37150 18790
rect 37358 18582 37881 18790
rect 36468 17048 36852 17152
rect 10957 16418 11067 16423
rect 10957 16318 10962 16418
rect 11062 16318 11067 16418
rect 11464 16322 36558 16422
rect 10957 16313 11067 16318
rect 36254 16193 36354 16198
rect 36254 16103 36259 16193
rect 36349 16103 36354 16193
rect 11201 15882 11311 15887
rect 11201 15782 11206 15882
rect 11306 15782 36158 15882
rect 11201 15777 11311 15782
rect -13304 15385 -13204 15396
rect -13304 15325 -13286 15385
rect -13226 15325 -13204 15385
rect -13304 14732 -13204 15325
rect -10642 15385 -10542 15410
rect -10642 15325 -10620 15385
rect -10560 15325 -10542 15385
rect -10642 14732 -10542 15325
rect -1950 15152 35940 15182
rect -1950 15092 -1924 15152
rect -1864 15092 35940 15152
rect -1950 15070 35940 15092
rect -13304 14632 -10542 14732
rect -2396 14983 11062 14988
rect -2396 14893 10967 14983
rect 11057 14893 11062 14983
rect -2396 14888 11062 14893
rect -13472 14605 -13372 14610
rect -13472 14515 -13467 14605
rect -13377 14515 -13372 14605
rect -13472 10731 -13372 14515
rect -13477 10633 -13471 10731
rect -13373 10633 -13367 10731
rect -13472 10632 -13372 10633
rect -13304 3537 -13204 14632
rect -8836 14174 -8646 14180
rect -11154 14168 -11008 14174
rect -11154 14002 -11008 14022
rect -12476 13984 -8836 14002
rect -3940 14168 -3782 14174
rect -6346 14150 -6170 14156
rect -8646 13984 -6346 14002
rect -12476 13974 -6346 13984
rect -3940 14002 -3782 14010
rect -6170 13974 -2606 14002
rect -12476 13400 -2606 13974
rect -12476 13398 -7666 13400
rect -13108 13137 -13008 13138
rect -13113 13039 -13107 13137
rect -13009 13039 -13003 13137
rect -13108 12772 -13006 13039
rect -13106 9154 -13006 12772
rect -12476 11974 -11875 13398
rect -10580 13038 -10574 13138
rect -10474 13120 -7214 13138
rect -10474 13060 -9878 13120
rect -9818 13060 -7214 13120
rect -10474 13038 -7214 13060
rect -9994 12784 -9894 13038
rect -12630 11880 -12624 11974
rect -12530 11880 -11875 11974
rect -12476 10010 -11875 11880
rect -9960 11192 -9894 12784
rect -7314 12716 -7214 13038
rect -3207 12166 -2606 13400
rect -2396 12904 -2296 14888
rect 11201 14812 11311 14817
rect 10974 14810 11206 14812
rect -1756 14712 11206 14810
rect 11306 14712 11311 14812
rect -1756 14710 11311 14712
rect -2402 12804 -2396 12904
rect -2296 12804 -2290 12904
rect -3207 11856 -2604 12166
rect -3207 11764 -2524 11856
rect -2432 11764 -2426 11856
rect -3207 11566 -2604 11764
rect -9960 11043 -9846 11128
rect -9960 10939 -9955 11043
rect -9851 10939 -9846 11043
rect -9226 11029 -9126 11252
rect -9960 10934 -9846 10939
rect -9231 10931 -9225 11029
rect -9127 10931 -9121 11029
rect -5826 11027 -5720 11164
rect -5270 11029 -5170 11234
rect -5826 10931 -5821 11027
rect -5725 10931 -5720 11027
rect -5275 10931 -5269 11029
rect -5171 10931 -5165 11029
rect -9226 10930 -9126 10931
rect -5826 10926 -5720 10931
rect -5270 10930 -5170 10931
rect -8101 10882 -8003 10887
rect -7570 10882 -7470 10888
rect -8102 10881 -7570 10882
rect -8102 10783 -8101 10881
rect -8003 10783 -7570 10881
rect -8102 10782 -7570 10783
rect -3901 10880 -3803 10885
rect -3392 10880 -3292 10886
rect -8101 10777 -8003 10782
rect -7570 10776 -7470 10782
rect -3902 10879 -3392 10880
rect -3902 10781 -3901 10879
rect -3803 10781 -3392 10879
rect -3902 10780 -3392 10781
rect -3292 10780 -3288 10880
rect -3901 10775 -3803 10780
rect -3392 10774 -3292 10780
rect -6556 10733 -6456 10734
rect -10356 10731 -10256 10732
rect -10361 10633 -10355 10731
rect -10257 10633 -10251 10731
rect -8786 10725 -8662 10730
rect -10356 10588 -10256 10633
rect -8786 10611 -8781 10725
rect -8667 10611 -8662 10725
rect -8786 10606 -8662 10611
rect -10356 10476 -10202 10588
rect -10302 10450 -10202 10476
rect -12640 9930 -12634 10010
rect -12554 9930 -11875 10010
rect -13106 9054 -12632 9154
rect -13100 8619 -13000 8620
rect -13105 8521 -13099 8619
rect -13001 8521 -12995 8619
rect -13309 3439 -13303 3537
rect -13205 3439 -13199 3537
rect -13304 3438 -13204 3439
rect -13100 1627 -13000 8521
rect -12732 5665 -12632 9054
rect -12476 8260 -11875 9930
rect -10132 8620 -10032 10450
rect -8781 10315 -8667 10606
rect -7192 10492 -7190 10684
rect -6561 10635 -6555 10733
rect -6457 10635 -6451 10733
rect -4794 10715 -4678 10720
rect -6556 10476 -6456 10635
rect -4794 10609 -4789 10715
rect -4683 10609 -4678 10715
rect -4794 10604 -4678 10609
rect -4789 10433 -4683 10604
rect -3207 9848 -2606 11566
rect -1756 11018 -1656 14710
rect 11201 14707 11311 14710
rect -3207 9742 -2518 9848
rect -2412 9742 -2406 9848
rect -7192 8620 -7092 9154
rect -10540 8520 -10534 8620
rect -10434 8520 -7092 8620
rect -6953 8262 -6351 8264
rect -5974 8262 -4547 8264
rect -4183 8262 -3581 8264
rect -3207 8262 -2606 9742
rect -1758 8863 -1656 11018
rect 35828 9127 35940 15070
rect 36058 9716 36158 15782
rect 36254 15375 36354 16103
rect 36249 15277 36255 15375
rect 36353 15277 36359 15375
rect 35828 9025 35833 9127
rect 35935 9025 35940 9127
rect 35828 9020 35940 9025
rect 36054 9311 36158 9716
rect 36254 9541 36354 15277
rect 36458 13819 36558 16322
rect 36451 13814 36561 13819
rect 36451 13714 36456 13814
rect 36556 13714 36561 13814
rect 36451 13709 36561 13714
rect 36249 9443 36255 9541
rect 36353 9443 36359 9541
rect 36254 9442 36354 9443
rect 36054 9306 36165 9311
rect 36054 9206 36060 9306
rect 36160 9206 36165 9306
rect 36054 9201 36165 9206
rect -1761 8765 -1755 8863
rect -1657 8765 -1651 8863
rect -11351 8260 -2606 8262
rect -12476 7662 -2606 8260
rect 35229 7738 35327 7743
rect 11362 7737 35328 7738
rect -12476 7660 -6020 7662
rect -4183 7660 -3581 7662
rect -11204 7646 -10950 7660
rect -11204 7406 -11197 7646
rect -10957 7556 -10950 7646
rect -8792 7646 -8538 7660
rect -10957 7406 -10951 7556
rect -8792 7406 -8785 7646
rect -8545 7556 -8538 7646
rect -6380 7646 -6126 7660
rect -8545 7406 -8539 7556
rect -6380 7406 -6373 7646
rect -6133 7556 -6126 7646
rect -3968 7646 -3714 7660
rect -6133 7406 -6127 7556
rect -3968 7406 -3961 7646
rect -3721 7556 -3714 7646
rect 11362 7639 35229 7737
rect 35327 7639 35328 7737
rect 11362 7638 35328 7639
rect -3721 7406 -3715 7556
rect -11204 7056 -10954 7406
rect -11204 6814 -11198 7056
rect -10956 6814 -10954 7056
rect -11204 6812 -10954 6814
rect -8792 7056 -8542 7406
rect -8792 6814 -8786 7056
rect -8544 6814 -8542 7056
rect -8792 6812 -8542 6814
rect -6380 7056 -6130 7406
rect -6380 6814 -6374 7056
rect -6132 6814 -6130 7056
rect -6380 6812 -6130 6814
rect -3968 7056 -3718 7406
rect 11362 7198 11462 7638
rect 35229 7633 35327 7638
rect 11362 7138 11382 7198
rect 11442 7138 11462 7198
rect 11362 7102 11462 7138
rect -3968 6814 -3962 7056
rect -3720 6814 -3718 7056
rect -3968 6812 -3718 6814
rect -12474 6798 -2604 6812
rect -12475 6712 -2604 6798
rect -12475 6198 -2607 6712
rect -12737 5567 -12731 5665
rect -12633 5567 -12627 5665
rect -12732 5566 -12632 5567
rect -12475 4766 -11875 6198
rect -12592 4616 -12586 4766
rect -12436 4616 -11875 4766
rect -12475 2650 -11875 4616
rect -9948 5852 -7198 5952
rect -9948 4138 -9848 5852
rect -7298 5478 -7198 5852
rect -3207 4716 -2607 6198
rect -2426 5665 -2322 5666
rect -2427 5567 -2421 5665
rect -2323 5567 -2317 5665
rect -2426 5228 -2322 5567
rect -2426 5226 8314 5228
rect -2426 5204 8366 5226
rect -2426 5144 8280 5204
rect 8340 5144 8366 5204
rect -2426 5126 8366 5144
rect -2426 5124 8314 5126
rect -3207 4562 -2660 4716
rect -2506 4562 -2500 4716
rect -10820 3835 -10716 3856
rect -10820 3741 -10815 3835
rect -10721 3741 -10716 3835
rect -9366 3827 -9266 4098
rect -6742 3827 -6642 3888
rect -5144 3839 -5028 4060
rect -10820 3736 -10716 3741
rect -9371 3729 -9365 3827
rect -9267 3729 -9261 3827
rect -6742 3737 -6737 3827
rect -6647 3737 -6642 3827
rect -6742 3732 -6642 3737
rect -9366 3728 -9266 3729
rect -5149 3725 -5143 3839
rect -5029 3725 -5023 3839
rect -5144 3724 -5028 3725
rect -8085 3682 -7987 3687
rect -7554 3682 -7454 3688
rect -3885 3684 -3787 3689
rect -3382 3684 -3282 3690
rect -8086 3681 -7554 3682
rect -8086 3583 -8085 3681
rect -7987 3583 -7554 3681
rect -8086 3582 -7554 3583
rect -3886 3683 -3382 3684
rect -3886 3585 -3885 3683
rect -3787 3585 -3382 3683
rect -3886 3584 -3382 3585
rect -8085 3577 -7987 3582
rect -7554 3576 -7454 3582
rect -3885 3579 -3787 3584
rect -3382 3578 -3282 3584
rect -10168 3537 -10068 3538
rect -10173 3439 -10167 3537
rect -10069 3439 -10063 3537
rect -9015 3514 -8901 3519
rect -10168 3194 -10068 3439
rect -9015 3410 -9010 3514
rect -8906 3410 -8901 3514
rect -9015 3405 -8901 3410
rect -9010 3238 -8906 3405
rect -7176 3254 -7174 3446
rect -5914 3426 -5908 3542
rect -5792 3426 -5786 3542
rect -4641 3510 -4531 3515
rect -5908 3332 -5792 3426
rect -4641 3410 -4636 3510
rect -4536 3410 -4531 3510
rect -4641 3405 -4531 3410
rect -4636 3174 -4536 3405
rect -12586 2524 -12580 2650
rect -12454 2524 -11875 2650
rect -13103 1529 -13097 1627
rect -12999 1529 -12993 1627
rect -13100 1528 -13000 1529
rect -12475 1062 -11875 2524
rect -10086 1422 -9986 3082
rect -3207 3060 -2607 4562
rect -3207 2664 -2608 3060
rect -3207 2504 -2666 2664
rect -2506 2504 -2500 2664
rect -3207 2202 -2608 2504
rect 36054 2238 36158 9201
rect 36458 6197 36558 13709
rect 36748 13581 36852 17048
rect 37279 16650 37881 18582
rect 50792 18732 51393 20420
rect 50792 18570 51338 18732
rect 51500 18570 51506 18732
rect 38968 17829 39076 17892
rect 40416 17829 40516 18064
rect 43134 17841 43262 17960
rect 38968 17731 38973 17829
rect 39071 17731 39076 17829
rect 40411 17731 40417 17829
rect 40515 17731 40521 17829
rect 38968 17726 39076 17731
rect 40416 17730 40516 17731
rect 43134 17723 43139 17841
rect 43257 17723 43262 17841
rect 44642 17817 44742 18054
rect 47326 17831 47436 17902
rect 43134 17718 43262 17723
rect 44637 17719 44643 17817
rect 44741 17719 44747 17817
rect 47326 17731 47331 17831
rect 47431 17731 47436 17831
rect 48764 17827 48864 18046
rect 47326 17726 47436 17731
rect 48759 17729 48765 17827
rect 48863 17729 48869 17827
rect 48764 17728 48864 17729
rect 44642 17718 44742 17719
rect 41673 17678 41771 17683
rect 42204 17678 42304 17684
rect 45873 17678 45971 17683
rect 46404 17678 46504 17684
rect 50073 17678 50171 17683
rect 50604 17678 50704 17684
rect 41672 17677 42204 17678
rect 41672 17579 41673 17677
rect 41771 17579 42204 17677
rect 41672 17578 42204 17579
rect 45872 17677 46404 17678
rect 45872 17579 45873 17677
rect 45971 17579 46404 17677
rect 45872 17578 46404 17579
rect 50072 17677 50604 17678
rect 50072 17579 50073 17677
rect 50171 17579 50604 17677
rect 50072 17578 50604 17579
rect 41673 17573 41771 17578
rect 42204 17572 42304 17578
rect 45873 17573 45971 17578
rect 46404 17572 46504 17578
rect 50073 17573 50171 17578
rect 50604 17572 50704 17578
rect 45183 17526 45321 17531
rect 39618 17523 39718 17524
rect 43818 17523 43918 17524
rect 39613 17425 39619 17523
rect 39717 17425 39723 17523
rect 40989 17516 41107 17521
rect 39618 17384 39718 17425
rect 40989 17408 40994 17516
rect 41102 17408 41107 17516
rect 43813 17425 43819 17523
rect 43917 17425 43923 17523
rect 40989 17403 41107 17408
rect 39618 17272 39772 17384
rect 37073 16464 37079 16650
rect 37265 16464 37881 16650
rect 37279 14870 37881 16464
rect 39672 15376 39772 17272
rect 40994 17156 41102 17403
rect 43818 17272 43918 17425
rect 45183 17398 45188 17526
rect 45316 17398 45321 17526
rect 48018 17521 48118 17522
rect 48013 17423 48019 17521
rect 48117 17423 48123 17521
rect 49278 17507 49398 17512
rect 45183 17393 45321 17398
rect 45188 17194 45316 17393
rect 48018 17272 48118 17423
rect 49278 17397 49283 17507
rect 49393 17397 49398 17507
rect 49278 17392 49398 17397
rect 49283 17165 49393 17392
rect 50792 16638 51393 18570
rect 50792 16470 51364 16638
rect 51532 16470 51538 16638
rect 42582 15376 42682 15950
rect 46660 15376 46760 15844
rect 39292 15276 39298 15376
rect 39398 15276 46760 15376
rect 50792 14870 51393 16470
rect 37131 14316 51393 14870
rect 52144 14738 52244 23614
rect 65088 18913 65188 18918
rect 65088 18823 65093 18913
rect 65183 18823 65188 18913
rect 65088 18818 65188 18823
rect 52380 15100 52480 15106
rect 64976 15100 65076 16422
rect 52480 15000 65076 15100
rect 52380 14994 52480 15000
rect 65083 14738 65193 14743
rect 52144 14638 65088 14738
rect 65188 14638 65193 14738
rect 65083 14633 65193 14638
rect 37131 14260 38478 14316
rect 36743 13483 36749 13581
rect 36847 13483 36853 13581
rect 37131 13527 37731 14260
rect 38636 14260 40890 14316
rect 38478 14152 38636 14158
rect 41048 14260 43290 14316
rect 40890 14152 41048 14158
rect 43448 14260 45690 14316
rect 43290 14152 43448 14158
rect 45848 14268 47690 14316
rect 45848 14260 46992 14268
rect 45690 14152 45848 14158
rect 39248 13809 42430 13814
rect 39248 13719 39253 13809
rect 39343 13719 42430 13809
rect 39248 13714 42430 13719
rect 36748 13480 36852 13483
rect 37131 12668 37733 13527
rect 39568 13134 39668 13714
rect 42330 13394 42430 13714
rect 36996 12460 37002 12668
rect 37210 12460 37733 12668
rect 37131 10528 37733 12460
rect 46399 12734 46992 14260
rect 47848 14268 50090 14316
rect 47690 14152 47848 14158
rect 50248 14268 51393 14316
rect 50792 14264 51393 14268
rect 50090 14152 50248 14158
rect 46399 12610 46999 12734
rect 46399 12448 47030 12610
rect 47192 12448 47198 12610
rect 46399 12380 46999 12448
rect 38844 11711 38950 11868
rect 38844 11615 38849 11711
rect 38945 11615 38950 11711
rect 40292 11709 40392 11914
rect 42994 11727 43130 11854
rect 38844 11610 38950 11615
rect 40287 11611 40293 11709
rect 40391 11611 40397 11709
rect 40292 11610 40392 11611
rect 42994 11597 42999 11727
rect 43125 11597 43130 11727
rect 44512 11709 44612 11890
rect 44507 11611 44513 11709
rect 44611 11611 44617 11709
rect 44512 11610 44612 11611
rect 42994 11592 43130 11597
rect 41543 11560 41641 11565
rect 42074 11560 42174 11566
rect 45743 11560 45841 11565
rect 46218 11560 46318 11566
rect 41542 11559 42074 11560
rect 41542 11461 41543 11559
rect 41641 11461 42074 11559
rect 41542 11460 42074 11461
rect 45742 11559 46218 11560
rect 45742 11461 45743 11559
rect 45841 11461 46218 11559
rect 45742 11460 46218 11461
rect 41543 11455 41641 11460
rect 42074 11454 42174 11460
rect 45743 11455 45841 11460
rect 46218 11454 46318 11460
rect 39488 11411 39588 11412
rect 39483 11313 39489 11411
rect 39587 11313 39593 11411
rect 43688 11393 43788 11394
rect 40880 11381 40996 11386
rect 39488 11266 39588 11313
rect 40880 11275 40885 11381
rect 40991 11275 40996 11381
rect 43683 11295 43689 11393
rect 43787 11295 43793 11393
rect 45045 11392 45163 11397
rect 40880 11270 40996 11275
rect 39488 11154 39642 11266
rect 36925 10342 36931 10528
rect 37117 10342 37733 10528
rect 37131 8932 37733 10342
rect 39542 9306 39642 11154
rect 40885 10991 40991 11270
rect 43688 11154 43788 11295
rect 45045 11284 45050 11392
rect 45158 11284 45163 11392
rect 45045 11279 45163 11284
rect 45050 11168 45158 11279
rect 45008 11090 45158 11168
rect 45050 11088 45158 11090
rect 45010 11078 45158 11088
rect 45010 10952 45146 11078
rect 46399 10634 46992 12380
rect 46399 10510 46999 10634
rect 46399 10342 46992 10510
rect 47160 10342 47166 10510
rect 46399 9958 46999 10342
rect 42452 9306 42552 9832
rect 39004 9301 42552 9306
rect 39004 9211 39009 9301
rect 39099 9211 42552 9301
rect 39004 9206 42552 9211
rect 46399 9218 47037 9958
rect 46399 8932 46999 9218
rect 37131 8400 46999 8932
rect 37131 8330 38476 8400
rect 37131 8328 37731 8330
rect 38704 8398 46999 8400
rect 38704 8328 40888 8398
rect 40886 8312 40888 8328
rect 38476 8166 38704 8172
rect 41116 8328 43232 8398
rect 43230 8312 43232 8328
rect 40888 8164 41116 8170
rect 43460 8330 45620 8398
rect 43460 8328 44542 8330
rect 43232 8164 43460 8170
rect 45848 8348 46999 8398
rect 45848 8330 46992 8348
rect 45848 8310 45850 8330
rect 45620 8164 45848 8170
rect 36990 7638 36996 7738
rect 37096 7638 47596 7738
rect 53050 7722 53150 7728
rect 47496 7222 47596 7638
rect 49800 7700 53050 7722
rect 49800 7640 49822 7700
rect 49882 7640 53050 7700
rect 49800 7622 53050 7640
rect 53050 7616 53150 7622
rect 47494 7198 62432 7222
rect 38428 7174 38610 7180
rect 37150 7064 38428 7078
rect 37149 6992 38428 7064
rect 40828 7174 41010 7180
rect 38610 6992 40828 7078
rect 43240 7174 43422 7180
rect 41010 6992 43240 7078
rect 45640 7174 45822 7180
rect 43422 6992 45640 7078
rect 47494 7138 62350 7198
rect 62410 7138 62432 7198
rect 47494 7122 62432 7138
rect 45822 6992 47017 7078
rect 37149 6464 47017 6992
rect 36453 6099 36459 6197
rect 36557 6099 36563 6197
rect 36458 6098 36558 6099
rect 37149 5066 37749 6464
rect 45911 6198 46021 6203
rect 39048 6098 39054 6198
rect 39154 6098 45916 6198
rect 46016 6098 46021 6198
rect 39368 5682 39468 6098
rect 42330 5794 42430 6098
rect 45911 6093 46021 6098
rect 37014 4858 37020 5066
rect 37228 4858 37749 5066
rect 37149 2926 37749 4858
rect 46417 5008 47017 6464
rect 48476 5981 48576 5982
rect 48471 5883 48477 5981
rect 48575 5883 48581 5981
rect 48476 5758 48576 5883
rect 48476 5736 49388 5758
rect 48476 5676 49306 5736
rect 49366 5676 49388 5736
rect 48476 5658 49388 5676
rect 53048 5604 53148 5610
rect 49924 5587 53048 5604
rect 49924 5527 49940 5587
rect 50000 5527 53048 5587
rect 49924 5504 53048 5527
rect 53048 5498 53148 5504
rect 46417 4846 47048 5008
rect 47210 4846 47216 5008
rect 52183 4956 52281 4961
rect 52183 4955 66110 4956
rect 52281 4936 66110 4955
rect 52281 4876 66026 4936
rect 66086 4876 66110 4936
rect 52281 4857 66110 4876
rect 52183 4856 66110 4857
rect 52183 4851 52281 4856
rect 38910 4099 39020 4204
rect 40278 4105 40378 4356
rect 38910 3999 38915 4099
rect 39015 3999 39020 4099
rect 40273 4007 40279 4105
rect 40377 4007 40383 4105
rect 43082 4097 43192 4226
rect 40278 4006 40378 4007
rect 38910 3994 39020 3999
rect 43082 3997 43087 4097
rect 43187 3997 43192 4097
rect 44490 4089 44590 4350
rect 43082 3992 43192 3997
rect 44485 3991 44491 4089
rect 44589 3991 44595 4089
rect 44490 3990 44590 3991
rect 41543 3960 41641 3965
rect 42074 3960 42174 3966
rect 45743 3960 45841 3965
rect 46238 3960 46338 3966
rect 41542 3959 42074 3960
rect 41542 3861 41543 3959
rect 41641 3861 42074 3959
rect 41542 3860 42074 3861
rect 45742 3959 46238 3960
rect 45742 3861 45743 3959
rect 45841 3861 46238 3959
rect 45742 3860 46238 3861
rect 41543 3855 41641 3860
rect 42074 3854 42174 3860
rect 45743 3855 45841 3860
rect 46238 3854 46338 3860
rect 40780 3799 40900 3804
rect 43688 3799 43788 3800
rect 39488 3797 39588 3798
rect 39483 3699 39489 3797
rect 39587 3699 39593 3797
rect 39488 3666 39588 3699
rect 40780 3689 40785 3799
rect 40895 3689 40900 3799
rect 43683 3701 43689 3799
rect 43787 3701 43793 3799
rect 45056 3787 45176 3792
rect 40780 3684 40900 3689
rect 39488 3554 39642 3666
rect 36943 2740 36949 2926
rect 37135 2740 37749 2926
rect -7176 1422 -7076 1916
rect -10086 1322 -7076 1422
rect -3207 1064 -2607 2202
rect 36054 1691 36154 2238
rect -2334 1625 -2234 1626
rect -2339 1527 -2333 1625
rect -2235 1527 -2229 1625
rect 36049 1593 36055 1691
rect 36153 1593 36159 1691
rect 36054 1592 36154 1593
rect -7140 1062 -2607 1064
rect -12475 512 -2607 1062
rect -12475 460 -11156 512
rect -10918 460 -8744 512
rect -11156 268 -10918 274
rect -8506 460 -6332 512
rect -8744 268 -8506 274
rect -6094 462 -3920 512
rect -6094 460 -5990 462
rect -3978 460 -3920 462
rect -6332 268 -6094 274
rect -3682 462 -2607 512
rect -2334 602 -2230 1527
rect 37149 1330 37749 2740
rect 39542 1692 39642 3554
rect 40785 3463 40895 3684
rect 43688 3554 43788 3701
rect 45056 3677 45061 3787
rect 45171 3677 45176 3787
rect 45056 3672 45176 3677
rect 45061 3381 45171 3672
rect 46417 2908 47017 4846
rect 48482 3756 48582 3762
rect 48582 3736 49378 3756
rect 48582 3676 49302 3736
rect 49362 3676 49378 3736
rect 48582 3656 49378 3676
rect 48482 3650 48582 3656
rect 52181 3605 52283 3611
rect 50066 3587 52181 3604
rect 50066 3527 50082 3587
rect 50142 3527 52181 3587
rect 50066 3504 52181 3527
rect 52181 3497 52283 3503
rect 61918 2933 62248 2938
rect 46417 2740 47010 2908
rect 47178 2740 47184 2908
rect 61918 2843 62153 2933
rect 62243 2843 62248 2933
rect 53051 2834 53149 2839
rect 61918 2838 62248 2843
rect 61918 2834 62018 2838
rect 53051 2833 62018 2834
rect 42452 1692 42552 2232
rect 39160 1592 39166 1692
rect 39266 1670 46162 1692
rect 39266 1610 46088 1670
rect 46148 1610 46162 1670
rect 39266 1592 46162 1610
rect 46417 1330 47017 2740
rect 53149 2735 62018 2833
rect 53051 2734 62018 2735
rect 53051 2729 53149 2734
rect 52177 1672 52287 1678
rect 49806 1646 52177 1672
rect 49806 1586 49828 1646
rect 49888 1586 52177 1646
rect 49806 1562 52177 1586
rect 52177 1556 52287 1562
rect 37149 798 47017 1330
rect 37149 728 38494 798
rect 37149 726 37749 728
rect -2334 582 8126 602
rect -2334 522 8042 582
rect 8102 522 8126 582
rect 38722 796 47017 798
rect 38722 726 40906 796
rect 40904 710 40906 726
rect 38494 564 38722 570
rect 41134 726 43250 796
rect 43248 710 43250 726
rect 40906 562 41134 568
rect 43478 728 45638 796
rect 43478 726 44560 728
rect 43250 562 43478 568
rect 45866 746 47017 796
rect 45866 728 47016 746
rect 45866 708 45868 728
rect 45638 562 45866 568
rect -2334 502 8126 522
rect -2334 500 -2234 502
rect -3682 460 -3578 462
rect -3920 268 -3682 274
<< via3 >>
rect -1419 27642 -1349 27647
rect -1419 27583 -1414 27642
rect -1414 27583 -1354 27642
rect -1354 27583 -1349 27642
rect 47824 27564 48462 27680
rect 38430 26420 38578 26568
rect 41348 26410 41506 26568
rect 37050 24644 37182 24776
rect 36468 23470 36568 23570
rect 42912 24632 43048 24768
rect 46576 24434 46676 24534
rect 40402 23770 40502 23870
rect 41563 23613 41661 23711
rect 42030 23612 42130 23712
rect 39493 23469 39591 23567
rect 37076 22556 37196 22676
rect 42864 22518 43004 22658
rect 49760 21600 49860 21700
rect 46405 21283 46503 21381
rect 52144 23614 52244 23714
rect 51794 20966 51894 21066
rect 36473 19827 36571 19925
rect 38494 20312 38672 20490
rect 40894 20312 41072 20490
rect 43294 20312 43472 20490
rect 45420 20312 45598 20490
rect 47594 20312 47772 20490
rect 49994 20312 50172 20490
rect 39078 19826 39178 19926
rect 37150 18582 37358 18790
rect -13471 10633 -13373 10731
rect -11154 14022 -11008 14168
rect -8836 13984 -8646 14174
rect -6346 13974 -6170 14150
rect -3940 14010 -3782 14168
rect -13107 13039 -13009 13137
rect -10574 13038 -10474 13138
rect -12624 11880 -12530 11974
rect -2396 12804 -2296 12904
rect -2524 11764 -2432 11856
rect -9225 10931 -9127 11029
rect -5269 10931 -5171 11029
rect -8101 10783 -8003 10881
rect -7570 10782 -7470 10882
rect -3901 10781 -3803 10879
rect -3392 10780 -3292 10880
rect -10355 10633 -10257 10731
rect -12634 9930 -12554 10010
rect -13099 8521 -13001 8619
rect -13303 3439 -13205 3537
rect -6555 10635 -6457 10733
rect -2518 9742 -2412 9848
rect -10534 8520 -10434 8620
rect 36255 15277 36353 15375
rect 36255 9443 36353 9541
rect -1755 8765 -1657 8863
rect -11197 7406 -10957 7646
rect -8785 7406 -8545 7646
rect -6373 7406 -6133 7646
rect -3961 7406 -3721 7646
rect 35229 7639 35327 7737
rect -11198 6814 -10956 7056
rect -8786 6814 -8544 7056
rect -6374 6814 -6132 7056
rect -3962 6814 -3720 7056
rect -12731 5567 -12633 5665
rect -12586 4616 -12436 4766
rect -2421 5567 -2323 5665
rect -2660 4562 -2506 4716
rect -9365 3729 -9267 3827
rect -5143 3725 -5029 3839
rect -8085 3583 -7987 3681
rect -7554 3582 -7454 3682
rect -3885 3585 -3787 3683
rect -3382 3584 -3282 3684
rect -10167 3439 -10069 3537
rect -5908 3426 -5792 3542
rect -12580 2524 -12454 2650
rect -13097 1529 -12999 1627
rect -2666 2504 -2506 2664
rect 51338 18570 51500 18732
rect 40417 17731 40515 17829
rect 44643 17719 44741 17817
rect 48765 17729 48863 17827
rect 41673 17579 41771 17677
rect 42204 17578 42304 17678
rect 45873 17579 45971 17677
rect 46404 17578 46504 17678
rect 50073 17579 50171 17677
rect 50604 17578 50704 17678
rect 39619 17425 39717 17523
rect 43819 17425 43917 17523
rect 37079 16464 37265 16650
rect 48019 17423 48117 17521
rect 51364 16470 51532 16638
rect 39298 15276 39398 15376
rect 52380 15000 52480 15100
rect 36749 13483 36847 13581
rect 38478 14158 38636 14316
rect 40890 14158 41048 14316
rect 43290 14158 43448 14316
rect 45690 14158 45848 14316
rect 37002 12460 37210 12668
rect 47690 14158 47848 14316
rect 50090 14158 50248 14316
rect 47030 12448 47192 12610
rect 40293 11611 40391 11709
rect 44513 11611 44611 11709
rect 41543 11461 41641 11559
rect 42074 11460 42174 11560
rect 45743 11461 45841 11559
rect 46218 11460 46318 11560
rect 39489 11313 39587 11411
rect 43689 11295 43787 11393
rect 36931 10342 37117 10528
rect 46992 10342 47160 10510
rect 38476 8172 38704 8400
rect 40888 8170 41116 8398
rect 43232 8170 43460 8398
rect 45620 8170 45848 8398
rect 36996 7638 37096 7738
rect 53050 7622 53150 7722
rect 38428 6992 38610 7174
rect 40828 6992 41010 7174
rect 43240 6992 43422 7174
rect 45640 6992 45822 7174
rect 36459 6099 36557 6197
rect 39054 6098 39154 6198
rect 37020 4858 37228 5066
rect 48477 5883 48575 5981
rect 53048 5504 53148 5604
rect 47048 4846 47210 5008
rect 52183 4857 52281 4955
rect 40279 4007 40377 4105
rect 44491 3991 44589 4089
rect 41543 3861 41641 3959
rect 42074 3860 42174 3960
rect 45743 3861 45841 3959
rect 46238 3860 46338 3960
rect 39489 3699 39587 3797
rect 43689 3701 43787 3799
rect 36949 2740 37135 2926
rect -2333 1527 -2235 1625
rect 36055 1593 36153 1691
rect -11156 274 -10918 512
rect -8744 274 -8506 512
rect -6332 274 -6094 512
rect -3920 274 -3682 512
rect 48482 3656 48582 3756
rect 52181 3503 52283 3605
rect 47010 2740 47178 2908
rect 39166 1592 39266 1692
rect 53051 2735 53149 2833
rect 52177 1562 52287 1672
rect 38494 570 38722 798
rect 40906 568 41134 796
rect 43250 568 43478 796
rect 45638 568 45866 796
<< metal4 >>
rect 33530 27680 55572 28340
rect -1420 27647 -1348 27648
rect -1420 27583 -1419 27647
rect -1349 27583 -1348 27647
rect -1420 27582 -1348 27583
rect 33530 27564 47824 27680
rect 48462 27564 55572 27680
rect 33530 27540 55572 27564
rect 38429 26568 38579 26569
rect 38429 26420 38430 26568
rect 38578 26420 38579 26568
rect 38429 26419 38579 26420
rect 41347 26568 41507 26569
rect 38430 26166 38578 26419
rect 41347 26410 41348 26568
rect 41506 26410 41507 26568
rect 41347 26409 41507 26410
rect 41348 26105 41506 26409
rect 39530 25634 46676 25734
rect 39530 25280 39630 25634
rect 37049 24776 37183 24777
rect 37049 24644 37050 24776
rect 37182 24644 37586 24776
rect 37049 24643 37183 24644
rect 41418 24614 41928 24714
rect 40401 23870 40503 23871
rect 40401 23770 40402 23870
rect 40502 23770 40503 23870
rect 36467 23570 36569 23571
rect 36467 23568 36468 23570
rect 36462 23470 36468 23568
rect 36568 23568 36569 23570
rect 40401 23568 40503 23770
rect 36568 23567 40503 23568
rect 36568 23470 39493 23567
rect 36462 23469 39493 23470
rect 39591 23469 40503 23567
rect 36462 23468 40503 23469
rect 40401 23467 40503 23468
rect 41562 23711 41662 23712
rect 41562 23613 41563 23711
rect 41661 23613 41662 23711
rect 41562 23212 41662 23613
rect 37075 22676 37197 22677
rect 37075 22556 37076 22676
rect 37196 22556 37492 22676
rect 37075 22555 37197 22556
rect 39512 21694 39612 22074
rect 41828 21694 41928 24614
rect 42030 23714 42130 25634
rect 42911 24768 43049 24769
rect 42584 24632 42912 24768
rect 43048 24632 43049 24768
rect 42911 24631 43049 24632
rect 46576 24535 46676 25634
rect 46575 24534 46677 24535
rect 46575 24434 46576 24534
rect 46676 24434 46677 24534
rect 46575 24433 46677 24434
rect 52143 23714 52245 23715
rect 42030 23713 52144 23714
rect 42029 23712 52144 23713
rect 42029 23612 42030 23712
rect 42130 23614 52144 23712
rect 52244 23614 52245 23714
rect 42130 23612 42131 23614
rect 52143 23613 52245 23614
rect 42029 23611 42131 23612
rect 42863 22658 43005 22659
rect 42582 22518 42864 22658
rect 43004 22518 43005 22658
rect 42863 22517 43005 22518
rect 49759 21700 49861 21701
rect 49759 21694 49760 21700
rect 39512 21600 49760 21694
rect 49860 21694 49861 21700
rect 52380 21694 52480 21696
rect 49860 21600 52480 21694
rect 39512 21594 52480 21600
rect 46404 21381 46504 21382
rect 46404 21283 46405 21381
rect 46503 21283 46504 21381
rect 38494 20491 38672 20787
rect 40894 20491 41072 20787
rect 43294 20491 43472 20787
rect 45420 20491 45598 20787
rect 38493 20490 38673 20491
rect 38493 20312 38494 20490
rect 38672 20312 38673 20490
rect 38493 20311 38673 20312
rect 40893 20490 41073 20491
rect 40893 20312 40894 20490
rect 41072 20312 41073 20490
rect 40893 20311 41073 20312
rect 43293 20490 43473 20491
rect 43293 20312 43294 20490
rect 43472 20312 43473 20490
rect 43293 20311 43473 20312
rect 45419 20490 45599 20491
rect 45419 20312 45420 20490
rect 45598 20312 45599 20490
rect 45419 20311 45599 20312
rect 39077 19926 39179 19927
rect 36472 19925 39078 19926
rect 36472 19827 36473 19925
rect 36571 19827 39078 19925
rect 36472 19826 39078 19827
rect 39178 19826 39179 19926
rect 39077 19825 39179 19826
rect 46404 19700 46504 21283
rect 51793 21066 51895 21067
rect 51793 20966 51794 21066
rect 51894 20966 52248 21066
rect 51793 20965 51895 20966
rect 47594 20491 47772 20787
rect 49994 20491 50172 20787
rect 47593 20490 47773 20491
rect 47593 20312 47594 20490
rect 47772 20312 47773 20490
rect 47593 20311 47773 20312
rect 49993 20490 50173 20491
rect 49993 20312 49994 20490
rect 50172 20312 50173 20490
rect 49993 20311 50173 20312
rect 39640 19600 50704 19700
rect 39640 19246 39740 19600
rect 37149 18790 37359 18791
rect 37149 18582 37150 18790
rect 37358 18582 37676 18790
rect 37149 18581 37359 18582
rect 41528 18580 42068 18680
rect 40416 17829 40516 17830
rect 40416 17731 40417 17829
rect 40515 17731 40516 17829
rect 40416 17524 40516 17731
rect 39618 17523 40516 17524
rect 39618 17425 39619 17523
rect 39717 17425 40516 17523
rect 39618 17424 40516 17425
rect 41672 17677 41772 17678
rect 41672 17579 41673 17677
rect 41771 17579 41772 17677
rect 41672 17178 41772 17579
rect 37078 16650 37266 16651
rect 37078 16464 37079 16650
rect 37265 16464 37629 16650
rect 37078 16463 37266 16464
rect 39622 15660 39722 16040
rect 41968 15660 42068 18580
rect 42204 17679 42304 19600
rect 43840 19246 43940 19600
rect 45728 18580 46268 18680
rect 44642 17817 44742 17818
rect 44642 17719 44643 17817
rect 44741 17719 44742 17817
rect 42203 17678 42305 17679
rect 42203 17578 42204 17678
rect 42304 17578 42305 17678
rect 42203 17577 42305 17578
rect 44642 17524 44742 17719
rect 43818 17523 44742 17524
rect 43818 17425 43819 17523
rect 43917 17425 44742 17523
rect 43818 17424 44742 17425
rect 45872 17677 45972 17678
rect 45872 17579 45873 17677
rect 45971 17579 45972 17677
rect 45872 17178 45972 17579
rect 43822 15660 43922 16040
rect 46168 15660 46268 18580
rect 46404 17679 46504 19600
rect 48040 19246 48140 19600
rect 49928 18580 50468 18680
rect 48764 17827 48864 17828
rect 48764 17729 48765 17827
rect 48863 17729 48864 17827
rect 46403 17678 46505 17679
rect 46403 17578 46404 17678
rect 46504 17578 46505 17678
rect 46403 17577 46505 17578
rect 48764 17522 48864 17729
rect 48018 17521 48864 17522
rect 48018 17423 48019 17521
rect 48117 17423 48864 17521
rect 48018 17422 48864 17423
rect 50072 17677 50172 17678
rect 50072 17579 50073 17677
rect 50171 17579 50172 17677
rect 50072 17178 50172 17579
rect 48022 15660 48122 16040
rect 50368 15660 50468 18580
rect 50604 17679 50704 19600
rect 51337 18732 51501 18733
rect 51037 18570 51338 18732
rect 51500 18570 51501 18732
rect 51337 18569 51501 18570
rect 50603 17678 50705 17679
rect 50603 17578 50604 17678
rect 50704 17578 50705 17678
rect 50603 17577 50705 17578
rect 51363 16638 51533 16639
rect 51014 16470 51364 16638
rect 51532 16470 51533 16638
rect 51363 16469 51533 16470
rect 52148 15660 52248 20966
rect 39622 15560 52248 15660
rect 39297 15376 39399 15377
rect 36254 15375 39298 15376
rect 36254 15277 36255 15375
rect 36353 15277 39298 15375
rect 36254 15276 39298 15277
rect 39398 15276 39399 15376
rect 39297 15275 39399 15276
rect 52380 15101 52480 21594
rect 52379 15100 52481 15101
rect 52379 15000 52380 15100
rect 52480 15000 52481 15100
rect 52379 14999 52481 15000
rect 38478 14317 38636 14613
rect 40890 14317 41048 14613
rect 43290 14317 43448 14613
rect 45690 14317 45848 14613
rect 47690 14317 47848 14613
rect 50090 14317 50248 14613
rect 38477 14316 38637 14317
rect -8837 14174 -8645 14175
rect -11155 14168 -11007 14169
rect -11155 14022 -11154 14168
rect -11008 14022 -11007 14168
rect -11155 14021 -11007 14022
rect -11154 13679 -11008 14021
rect -8837 13984 -8836 14174
rect -8646 13984 -8645 14174
rect -3941 14168 -3781 14169
rect -8837 13983 -8645 13984
rect -6347 14150 -6169 14151
rect -8836 13619 -8646 13983
rect -6347 13974 -6346 14150
rect -6170 13974 -6169 14150
rect -3941 14010 -3940 14168
rect -3782 14010 -3781 14168
rect 38477 14158 38478 14316
rect 38636 14158 38637 14316
rect 38477 14157 38637 14158
rect 40889 14316 41049 14317
rect 40889 14158 40890 14316
rect 41048 14158 41049 14316
rect 40889 14157 41049 14158
rect 43289 14316 43449 14317
rect 43289 14158 43290 14316
rect 43448 14158 43449 14316
rect 43289 14157 43449 14158
rect 45689 14316 45849 14317
rect 45689 14158 45690 14316
rect 45848 14158 45849 14316
rect 45689 14157 45849 14158
rect 47689 14316 47849 14317
rect 47689 14158 47690 14316
rect 47848 14158 47849 14316
rect 47689 14157 47849 14158
rect 50089 14316 50249 14317
rect 50089 14158 50090 14316
rect 50248 14158 50249 14316
rect 50089 14157 50249 14158
rect -3941 14009 -3781 14010
rect -6347 13973 -6169 13974
rect -6346 13602 -6170 13973
rect -3940 13667 -3782 14009
rect 36748 13581 46318 13582
rect 36748 13483 36749 13581
rect 36847 13483 46318 13581
rect 36748 13482 46318 13483
rect -10575 13138 -10473 13139
rect -13108 13137 -10574 13138
rect -13108 13039 -13107 13137
rect -13009 13039 -10574 13137
rect -13108 13038 -10574 13039
rect -10474 13038 -10473 13138
rect 39510 13128 39610 13482
rect -10575 13037 -10473 13038
rect -2397 12904 -2295 12905
rect -10164 12804 -2396 12904
rect -2296 12804 -2295 12904
rect -10164 12450 -10064 12804
rect -12625 11974 -12529 11975
rect -12625 11880 -12624 11974
rect -12530 11880 -12207 11974
rect -12625 11879 -12529 11880
rect -8246 11784 -7706 11884
rect -9226 11029 -9126 11030
rect -9226 10931 -9225 11029
rect -9127 10931 -9126 11029
rect -9226 10732 -9126 10931
rect -13472 10731 -9126 10732
rect -13472 10633 -13471 10731
rect -13373 10633 -10355 10731
rect -10257 10633 -9126 10731
rect -13472 10632 -9126 10633
rect -8102 10881 -8002 10882
rect -8102 10783 -8101 10881
rect -8003 10783 -8002 10881
rect -8102 10382 -8002 10783
rect -12635 10010 -12553 10011
rect -12635 9930 -12634 10010
rect -12554 9930 -12204 10010
rect -12635 9929 -12553 9930
rect -10182 8864 -10082 9244
rect -7806 8864 -7706 11784
rect -7570 10883 -7470 12804
rect -5934 12450 -5834 12804
rect -4046 11784 -3506 11884
rect -5270 11029 -5170 11030
rect -5270 10931 -5269 11029
rect -5171 10931 -5170 11029
rect -7571 10882 -7469 10883
rect -7571 10782 -7570 10882
rect -7470 10782 -7469 10882
rect -7571 10781 -7469 10782
rect -5270 10734 -5170 10931
rect -6556 10733 -5170 10734
rect -6556 10635 -6555 10733
rect -6457 10635 -5170 10733
rect -6556 10634 -5170 10635
rect -3902 10879 -3802 10880
rect -3902 10781 -3901 10879
rect -3803 10781 -3802 10879
rect -3902 10382 -3802 10781
rect -5952 8864 -5852 9244
rect -3606 8864 -3506 11784
rect -3392 10881 -3292 12804
rect -2397 12803 -2295 12804
rect 37001 12668 37211 12669
rect 37001 12460 37002 12668
rect 37210 12460 37528 12668
rect 41398 12462 41938 12562
rect 37001 12459 37211 12460
rect -2525 11856 -2431 11857
rect -2892 11764 -2524 11856
rect -2432 11764 -2431 11856
rect -2525 11763 -2431 11764
rect 40292 11709 40392 11710
rect 40292 11611 40293 11709
rect 40391 11611 40392 11709
rect 40292 11412 40392 11611
rect 39488 11411 40392 11412
rect 39488 11313 39489 11411
rect 39587 11313 40392 11411
rect 39488 11312 40392 11313
rect 41542 11559 41642 11560
rect 41542 11461 41543 11559
rect 41641 11461 41642 11559
rect 41542 11060 41642 11461
rect -3393 10880 -3291 10881
rect -3393 10780 -3392 10880
rect -3292 10780 -3291 10880
rect -3393 10779 -3291 10780
rect -3392 10776 -3292 10779
rect 36930 10528 37118 10529
rect 36930 10342 36931 10528
rect 37117 10342 37481 10528
rect 36930 10341 37118 10342
rect -2519 9848 -2411 9849
rect -2891 9742 -2518 9848
rect -2412 9742 -2411 9848
rect -2519 9741 -2411 9742
rect 39492 9542 39592 9922
rect 41838 9542 41938 12462
rect 42074 11561 42174 13482
rect 43710 13128 43810 13482
rect 45598 12462 46138 12562
rect 44512 11709 44612 11710
rect 44512 11611 44513 11709
rect 44611 11611 44612 11709
rect 42073 11560 42175 11561
rect 42073 11460 42074 11560
rect 42174 11460 42175 11560
rect 42073 11459 42175 11460
rect 44512 11394 44612 11611
rect 43688 11393 44612 11394
rect 43688 11295 43689 11393
rect 43787 11295 44612 11393
rect 43688 11294 44612 11295
rect 45742 11559 45842 11560
rect 45742 11461 45743 11559
rect 45841 11461 45842 11559
rect 45742 11060 45842 11461
rect 43692 9542 43792 9922
rect 46038 9542 46138 12462
rect 46218 11561 46318 13482
rect 47029 12610 47193 12611
rect 46679 12448 47030 12610
rect 47192 12448 47193 12610
rect 47029 12447 47193 12448
rect 46217 11560 46319 11561
rect 46217 11460 46218 11560
rect 46318 11556 46319 11560
rect 46318 11460 53150 11556
rect 46217 11459 53150 11460
rect 46218 11456 53150 11459
rect 46991 10510 47161 10511
rect 46658 10342 46992 10510
rect 47160 10342 47161 10510
rect 46991 10341 47161 10342
rect 36254 9541 52282 9542
rect 36254 9443 36255 9541
rect 36353 9443 52282 9541
rect 36254 9442 52282 9443
rect -10182 8863 -1656 8864
rect -10182 8765 -1755 8863
rect -1657 8765 -1656 8863
rect -10182 8764 -1656 8765
rect 38476 8638 38704 8726
rect -10535 8620 -10433 8621
rect -13100 8619 -10534 8620
rect -13100 8521 -13099 8619
rect -13001 8521 -10534 8619
rect -13100 8520 -10534 8521
rect -10434 8520 -10433 8620
rect -10535 8519 -10433 8520
rect 38394 8400 38748 8638
rect 40888 8600 41116 8726
rect 38394 8172 38476 8400
rect 38704 8172 38748 8400
rect -11198 7646 -10956 8059
rect -11198 7406 -11197 7646
rect -10957 7406 -10956 7646
rect -11198 7057 -10956 7406
rect -8786 7646 -8544 8059
rect -8786 7406 -8785 7646
rect -8545 7406 -8544 7646
rect -8786 7057 -8544 7406
rect -6374 7646 -6132 8059
rect -6374 7406 -6373 7646
rect -6133 7406 -6132 7646
rect -6374 7057 -6132 7406
rect -3962 7646 -3720 8059
rect 36995 7738 37097 7739
rect -3962 7406 -3961 7646
rect -3721 7406 -3720 7646
rect 35228 7737 36996 7738
rect 35228 7639 35229 7737
rect 35327 7639 36996 7737
rect 35228 7638 36996 7639
rect 37096 7638 37097 7738
rect 36995 7637 37097 7638
rect -3962 7057 -3720 7406
rect 38394 7174 38748 8172
rect -11199 7056 -10955 7057
rect -11199 6814 -11198 7056
rect -10956 6814 -10955 7056
rect -11199 6813 -10955 6814
rect -8787 7056 -8543 7057
rect -8787 6814 -8786 7056
rect -8544 6814 -8543 7056
rect -8787 6813 -8543 6814
rect -6375 7056 -6131 7057
rect -6375 6814 -6374 7056
rect -6132 6814 -6131 7056
rect -6375 6813 -6131 6814
rect -3963 7056 -3719 7057
rect -3963 6814 -3962 7056
rect -3720 6814 -3719 7056
rect -3963 6813 -3719 6814
rect 38394 6992 38428 7174
rect 38610 6992 38748 7174
rect -11198 6413 -10956 6813
rect -9421 6658 -9070 6659
rect -9421 6338 -9420 6658
rect -8786 6413 -8544 6813
rect -6374 6413 -6132 6813
rect -3962 6413 -3720 6813
rect 38394 6640 38748 6992
rect 40796 8398 41150 8600
rect 40796 8170 40888 8398
rect 41116 8170 41150 8398
rect 40796 7174 41150 8170
rect 40796 6992 40828 7174
rect 41010 6992 41150 7174
rect 38428 6635 38610 6640
rect 40796 6630 41150 6992
rect 43168 8398 43504 8730
rect 43168 8170 43232 8398
rect 43460 8170 43504 8398
rect 43168 7174 43504 8170
rect 43168 6992 43240 7174
rect 43422 6992 43504 7174
rect 43168 6620 43504 6992
rect 45576 8398 45872 8746
rect 45576 8170 45620 8398
rect 45848 8170 45872 8398
rect 45576 7174 45872 8170
rect 45576 6992 45640 7174
rect 45822 6992 45872 7174
rect 45576 6630 45872 6992
rect -9421 6337 -9070 6338
rect 39053 6198 39155 6199
rect 36458 6197 39054 6198
rect 36458 6099 36459 6197
rect 36557 6099 39054 6197
rect 36458 6098 39054 6099
rect 39154 6098 39155 6198
rect 39053 6097 39155 6098
rect 39510 5981 48576 5982
rect 39510 5883 48477 5981
rect 48575 5883 48576 5981
rect 39510 5882 48576 5883
rect -12732 5665 -2322 5666
rect -12732 5567 -12731 5665
rect -12633 5567 -2421 5665
rect -2323 5567 -2322 5665
rect -12732 5566 -2322 5567
rect -10118 5212 -10018 5566
rect -12587 4766 -12435 4767
rect -12587 4616 -12586 4766
rect -12436 4616 -12157 4766
rect -12587 4615 -12435 4616
rect -8230 4546 -7690 4646
rect -9366 3827 -9266 3828
rect -9366 3729 -9365 3827
rect -9267 3729 -9266 3827
rect -9366 3538 -9266 3729
rect -13304 3537 -9266 3538
rect -13304 3439 -13303 3537
rect -13205 3439 -10167 3537
rect -10069 3439 -9266 3537
rect -13304 3438 -9266 3439
rect -8086 3681 -7986 3682
rect -8086 3583 -8085 3681
rect -7987 3583 -7986 3681
rect -8086 3144 -7986 3583
rect -12581 2650 -12453 2651
rect -12581 2524 -12580 2650
rect -12454 2524 -12079 2650
rect -12581 2523 -12453 2524
rect -10136 1628 -10036 2006
rect -13098 1627 -9512 1628
rect -13098 1529 -13097 1627
rect -12999 1626 -9512 1627
rect -7790 1626 -7690 4546
rect -7554 3683 -7454 5566
rect -5918 5212 -5818 5566
rect -4030 4546 -3490 4646
rect -5144 3839 -5028 3840
rect -5144 3725 -5143 3839
rect -5029 3725 -5028 3839
rect -7555 3682 -7453 3683
rect -7555 3582 -7554 3682
rect -7454 3582 -7453 3682
rect -7555 3581 -7453 3582
rect -5909 3542 -5791 3543
rect -5144 3542 -5028 3725
rect -5909 3426 -5908 3542
rect -5792 3426 -5028 3542
rect -3886 3683 -3786 3684
rect -3886 3585 -3885 3683
rect -3787 3585 -3786 3683
rect -5909 3425 -5791 3426
rect -3886 3144 -3786 3585
rect -5936 1626 -5836 2006
rect -3590 1626 -3490 4546
rect -3382 3685 -3282 5566
rect 39510 5528 39610 5882
rect 37019 5066 37229 5067
rect 37019 4858 37020 5066
rect 37228 4858 37546 5066
rect 41398 4862 41938 4962
rect 37019 4857 37229 4858
rect -2661 4716 -2505 4717
rect -2943 4562 -2660 4716
rect -2506 4562 -2505 4716
rect -2661 4561 -2505 4562
rect 40278 4105 40378 4106
rect 40278 4007 40279 4105
rect 40377 4007 40378 4105
rect 40278 3798 40378 4007
rect 39488 3797 40378 3798
rect 39488 3699 39489 3797
rect 39587 3699 40378 3797
rect 39488 3698 40378 3699
rect 41542 3959 41642 3960
rect 41542 3861 41543 3959
rect 41641 3861 41642 3959
rect -3383 3684 -3281 3685
rect -3383 3584 -3382 3684
rect -3282 3584 -3281 3684
rect -3383 3583 -3281 3584
rect 41542 3460 41642 3861
rect 36948 2926 37136 2927
rect 36948 2740 36949 2926
rect 37135 2740 37499 2926
rect 36948 2739 37136 2740
rect -2667 2664 -2505 2665
rect -2926 2504 -2666 2664
rect -2506 2504 -2505 2664
rect -2667 2503 -2505 2504
rect 39492 1942 39592 2322
rect 41838 1942 41938 4862
rect 42074 3961 42174 5882
rect 43710 5528 43810 5882
rect 45598 4862 46138 4962
rect 44490 4089 44590 4090
rect 44490 3991 44491 4089
rect 44589 3991 44590 4089
rect 42073 3960 42175 3961
rect 42073 3860 42074 3960
rect 42174 3860 42175 3960
rect 42073 3859 42175 3860
rect 44490 3800 44590 3991
rect 43688 3799 44590 3800
rect 43688 3701 43689 3799
rect 43787 3701 44590 3799
rect 43688 3700 44590 3701
rect 45742 3959 45842 3960
rect 45742 3861 45743 3959
rect 45841 3861 45842 3959
rect 45742 3460 45842 3861
rect 43692 1942 43792 2322
rect 46038 1942 46138 4862
rect 46238 3961 46338 5882
rect 47047 5008 47211 5009
rect 46697 4846 47048 5008
rect 47210 4846 47211 5008
rect 47047 4845 47211 4846
rect 52182 4955 52282 9442
rect 53050 7723 53150 11456
rect 53049 7722 53151 7723
rect 53049 7622 53050 7722
rect 53150 7622 53151 7722
rect 53049 7621 53151 7622
rect 53050 5605 53150 7621
rect 53047 5604 53150 5605
rect 53047 5504 53048 5604
rect 53148 5504 53150 5604
rect 53047 5503 53150 5504
rect 52182 4857 52183 4955
rect 52281 4857 52282 4955
rect 52182 4087 52282 4857
rect 46237 3960 46339 3961
rect 46237 3860 46238 3960
rect 46338 3860 46339 3960
rect 46237 3859 46339 3860
rect 48481 3756 48583 3757
rect 48481 3656 48482 3756
rect 48582 3656 48583 3756
rect 48481 3655 48583 3656
rect 47009 2908 47179 2909
rect 46676 2740 47010 2908
rect 47178 2740 47179 2908
rect 47009 2739 47179 2740
rect 48482 1942 48582 3655
rect 52181 3606 52283 4087
rect 52180 3605 52284 3606
rect 52180 3503 52181 3605
rect 52283 3503 52284 3605
rect 52180 3502 52284 3503
rect 39492 1842 48582 1942
rect 52181 1897 52283 3502
rect 53050 2833 53150 5503
rect 53050 2735 53051 2833
rect 53149 2735 53150 2833
rect 53050 2734 53150 2735
rect 39165 1692 39267 1693
rect 36054 1691 39166 1692
rect -12999 1625 -2234 1626
rect -12999 1529 -2333 1625
rect -13098 1528 -2333 1529
rect -10136 1527 -2333 1528
rect -2235 1527 -2234 1625
rect 36054 1593 36055 1691
rect 36153 1593 39166 1691
rect 36054 1592 39166 1593
rect 39266 1592 39267 1692
rect 52177 1673 52287 1897
rect 39165 1591 39267 1592
rect 52176 1672 52288 1673
rect 52176 1562 52177 1672
rect 52287 1562 52288 1672
rect 52176 1561 52288 1562
rect -10136 1526 -2234 1527
rect -11156 513 -10918 859
rect -8744 513 -8506 859
rect -6332 513 -6094 859
rect -3920 513 -3682 859
rect 38494 799 38722 1124
rect 38493 798 38723 799
rect 38493 570 38494 798
rect 38722 570 38723 798
rect 40906 797 41134 1124
rect 43250 797 43478 1124
rect 45638 797 45866 1124
rect 38493 569 38723 570
rect 40905 796 41135 797
rect -11157 512 -10917 513
rect -11157 274 -11156 512
rect -10918 274 -10917 512
rect -11157 273 -10917 274
rect -8745 512 -8505 513
rect -8745 274 -8744 512
rect -8506 274 -8505 512
rect -8745 273 -8505 274
rect -6333 512 -6093 513
rect -6333 274 -6332 512
rect -6094 274 -6093 512
rect -6333 273 -6093 274
rect -3921 512 -3681 513
rect -3921 274 -3920 512
rect -3682 274 -3681 512
rect -3921 273 -3681 274
rect -11156 140 -10918 273
rect -8744 140 -8506 273
rect -6332 140 -6094 273
rect -3920 140 -3682 273
rect 38494 140 38722 569
rect 40905 568 40906 796
rect 41134 568 41135 796
rect 40905 567 41135 568
rect 43249 796 43479 797
rect 43249 568 43250 796
rect 43478 568 43479 796
rect 43249 567 43479 568
rect 45637 796 45867 797
rect 45637 568 45638 796
rect 45866 568 45867 796
rect 45637 567 45867 568
rect 40906 140 41134 567
rect 43250 140 43478 567
rect 45638 140 45866 567
rect -13292 -660 378 140
rect 34882 -660 90192 140
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/diff_to_se_converter
timestamp 1624477805
transform 1 0 -8610 0 1 762
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_5 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/diff_to_se_converter
timestamp 1624477805
transform 1 0 -8648 0 1 2584
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_4 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/diff_to_se_converter
timestamp 1624477805
transform 1 0 -12124 0 1 2580
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_4 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/diff_to_se_converter
timestamp 1624477805
transform -1 0 -11093 0 1 762
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_4
timestamp 1624477805
transform 1 0 -10678 0 1 2584
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_1
timestamp 1624477805
transform -1 0 -6322 0 1 764
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_6
timestamp 1624477805
transform 1 0 -6488 0 1 2584
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_5
timestamp 1624477805
transform -1 0 -2958 0 1 2582
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_5
timestamp 1624477805
transform 1 0 -3839 0 1 764
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_7
timestamp 1624477805
transform 1 0 -4448 0 1 2584
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_2
timestamp 1624477805
transform 1 0 -8610 0 1 6498
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_6
timestamp 1624477805
transform -1 0 -11093 0 1 6498
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_10
timestamp 1624477805
transform 1 0 -8648 0 1 4684
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_6
timestamp 1624477805
transform 1 0 -12124 0 1 4684
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_8
timestamp 1624477805
transform 1 0 -10678 0 1 4684
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_3
timestamp 1624477805
transform -1 0 -6322 0 1 6500
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_9
timestamp 1624477805
transform 1 0 -6488 0 1 4684
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_7
timestamp 1624477805
transform 1 0 -3839 0 1 6500
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_7
timestamp 1624477805
transform -1 0 -2958 0 1 4686
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_11
timestamp 1624477805
transform 1 0 -4448 0 1 4684
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_22
timestamp 1624477805
transform 1 0 -12124 0 1 9780
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_46
timestamp 1624477805
transform 1 0 -10678 0 1 9784
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_22
timestamp 1624477805
transform 1 0 -8610 0 1 7962
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_23
timestamp 1624477805
transform -1 0 -11093 0 1 7962
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_42
timestamp 1624477805
transform 1 0 -8648 0 1 9784
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_43
timestamp 1624477805
transform 1 0 -6488 0 1 9784
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_23
timestamp 1624477805
transform -1 0 -6322 0 1 7964
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_22
timestamp 1624477805
transform 1 0 -3839 0 1 7964
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_40
timestamp 1624477805
transform 1 0 -4448 0 1 9784
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_20
timestamp 1624477805
transform -1 0 -2958 0 1 9782
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_23
timestamp 1624477805
transform 1 0 -12124 0 1 11884
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_47
timestamp 1624477805
transform 1 0 -10678 0 1 11884
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_21
timestamp 1624477805
transform -1 0 -11093 0 1 13698
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_20
timestamp 1624477805
transform 1 0 -8610 0 1 13698
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_44
timestamp 1624477805
transform 1 0 -8648 0 1 11884
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_45
timestamp 1624477805
transform 1 0 -6488 0 1 11884
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_21
timestamp 1624477805
transform -1 0 -6322 0 1 13700
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_20
timestamp 1624477805
transform 1 0 -3839 0 1 13700
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_41
timestamp 1624477805
transform 1 0 -4448 0 1 11884
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_21
timestamp 1624477805
transform -1 0 -2958 0 1 11886
box -350 -900 244 900
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform -1 0 -7834 0 1 15218
box -38 -48 314 592
use txgate  txgate_5 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/txgate
timestamp 1625985445
transform 1 0 -84715 0 1 -42708
box 74185 57360 76542 59116
use txgate  txgate_4
timestamp 1625985445
transform 1 0 -87315 0 1 -42708
box 74185 57360 76542 59116
use diff_fold_casc_ota  diff_fold_casc_ota_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/diff_fold_casc_ota
timestamp 1624477805
transform 1 0 10950 0 1 26540
box -12400 -27258 25000 1800
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_32
timestamp 1624477805
transform 1 0 38946 0 1 2850
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_17
timestamp 1624477805
transform 1 0 37500 0 1 2846
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_16
timestamp 1624477805
transform -1 0 38531 0 1 1028
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_37
timestamp 1624477805
transform 1 0 43136 0 1 2850
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_34
timestamp 1624477805
transform 1 0 40976 0 1 2850
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_17
timestamp 1624477805
transform 1 0 41014 0 1 1028
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_16
timestamp 1624477805
transform -1 0 43302 0 1 1030
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_39
timestamp 1624477805
transform 1 0 45176 0 1 2850
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_17
timestamp 1624477805
transform 1 0 45785 0 1 1030
box -1350 -300 1232 300
use txgate  txgate_6
timestamp 1625985445
transform 1 0 -25531 0 1 -56596
box 74185 57360 76542 59116
use txgate  txgate_1
timestamp 1625985445
transform 1 0 -25531 0 1 -54506
box 74185 57360 76542 59116
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_18
timestamp 1624477805
transform -1 0 46666 0 1 2848
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_18
timestamp 1624477805
transform -1 0 38531 0 1 6764
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_33
timestamp 1624477805
transform 1 0 38946 0 1 4950
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_16
timestamp 1624477805
transform 1 0 37500 0 1 4950
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_19
timestamp 1624477805
transform 1 0 41014 0 1 6764
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_18
timestamp 1624477805
transform -1 0 43302 0 1 6766
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_36
timestamp 1624477805
transform 1 0 43136 0 1 4950
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_35
timestamp 1624477805
transform 1 0 40976 0 1 4950
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_19
timestamp 1624477805
transform 1 0 45785 0 1 6766
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_38
timestamp 1624477805
transform 1 0 45176 0 1 4950
box -950 -900 838 900
use txgate  txgate_0
timestamp 1625985445
transform 1 0 -25531 0 1 -52506
box 74185 57360 76542 59116
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_19
timestamp 1624477805
transform -1 0 46666 0 1 4952
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_24
timestamp 1624477805
transform 1 0 38928 0 1 10452
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_13
timestamp 1624477805
transform 1 0 37482 0 1 10448
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_12
timestamp 1624477805
transform -1 0 38513 0 1 8630
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_26
timestamp 1624477805
transform 1 0 40958 0 1 10452
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_27
timestamp 1624477805
transform 1 0 43118 0 1 10452
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_13
timestamp 1624477805
transform -1 0 43284 0 1 8632
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_12
timestamp 1624477805
transform 1 0 40996 0 1 8630
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_30
timestamp 1624477805
transform 1 0 45158 0 1 10452
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_13
timestamp 1624477805
transform 1 0 45767 0 1 8632
box -1350 -300 1232 300
use txgate  txgate_7
timestamp 1625985445
transform 1 0 -25531 0 1 -50542
box 74185 57360 76542 59116
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_14
timestamp 1624477805
transform -1 0 46648 0 1 10450
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_25
timestamp 1624477805
transform 1 0 38928 0 1 12552
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_12
timestamp 1624477805
transform 1 0 37482 0 1 12552
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_28
timestamp 1624477805
transform 1 0 40958 0 1 12552
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_29
timestamp 1624477805
transform 1 0 43118 0 1 12552
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_31
timestamp 1624477805
transform 1 0 45158 0 1 12552
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_15
timestamp 1624477805
transform -1 0 46648 0 1 12554
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_14
timestamp 1624477805
transform -1 0 38513 0 1 14566
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_8
timestamp 1624477805
transform 1 0 37630 0 1 16570
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_13
timestamp 1624477805
transform 1 0 39076 0 1 16574
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_12
timestamp 1624477805
transform 1 0 41106 0 1 16574
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_15
timestamp 1624477805
transform 1 0 40996 0 1 14566
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_14
timestamp 1624477805
transform -1 0 43284 0 1 14568
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_14
timestamp 1624477805
transform 1 0 43266 0 1 16574
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_4
timestamp 1624477805
transform -1 0 45566 0 1 14568
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_15
timestamp 1624477805
transform 1 0 45306 0 1 16574
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_6
timestamp 1624477805
transform -1 0 47678 0 1 14568
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_23
timestamp 1624477805
transform 1 0 47462 0 1 16574
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_10
timestamp 1624477805
transform 1 0 50161 0 1 14568
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_22
timestamp 1624477805
transform 1 0 49502 0 1 16574
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_11
timestamp 1624477805
transform -1 0 51042 0 1 16570
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_3
timestamp 1624477805
transform -1 0 38513 0 1 20726
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_9
timestamp 1624477805
transform 1 0 37630 0 1 18674
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_17
timestamp 1624477805
transform 1 0 39076 0 1 18674
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_16
timestamp 1624477805
transform 1 0 41106 0 1 18674
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_9
timestamp 1624477805
transform 1 0 40996 0 1 20726
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_8
timestamp 1624477805
transform -1 0 43284 0 1 20728
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_18
timestamp 1624477805
transform 1 0 43266 0 1 18674
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_5
timestamp 1624477805
transform -1 0 45392 0 1 20728
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_19
timestamp 1624477805
transform 1 0 45306 0 1 18674
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_7
timestamp 1624477805
transform -1 0 47678 0 1 20728
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_20
timestamp 1624477805
transform 1 0 47462 0 1 18674
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_2
timestamp 1624477805
transform 1 0 50161 0 1 20728
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_21
timestamp 1624477805
transform 1 0 49502 0 1 18674
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_10
timestamp 1624477805
transform -1 0 51042 0 1 18674
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_1
timestamp 1624477805
transform 1 0 37516 0 1 22612
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_0
timestamp 1624477805
transform 1 0 37516 0 1 24716
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_3
timestamp 1624477805
transform 1 0 38968 0 1 24712
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_0
timestamp 1624477805
transform 1 0 38968 0 1 22612
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_2
timestamp 1624477805
transform 1 0 40998 0 1 24712
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_1
timestamp 1624477805
transform 1 0 40998 0 1 22612
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_3
timestamp 1624477805
transform 1 0 42616 0 1 22612
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_2
timestamp 1624477805
transform 1 0 42616 0 1 24716
box -350 -900 244 900
use txgate  txgate_2
timestamp 1625985445
transform 1 0 -26957 0 1 -35578
box 74185 57360 76542 59116
use txgate  txgate_3
timestamp 1625985445
transform 1 0 -26957 0 1 -33578
box 74185 57360 76542 59116
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_0
timestamp 1624477805
transform -1 0 38400 0 1 26180
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_1
timestamp 1624477805
transform -1 0 41400 0 1 26180
box -1350 -300 1232 300
use diff_fold_casc_ota  diff_fold_casc_ota_1
timestamp 1624477805
transform 1 0 64950 0 1 26540
box -12400 -27258 25000 1800
<< labels >>
flabel metal4 -9700 5602 -9690 5614 1 FreeSans 480 0 0 0 vip1
flabel metal4 -9752 1570 -9732 1586 1 FreeSans 480 0 0 0 vim1
flabel metal4 -5616 -342 -5562 -296 1 FreeSans 480 0 0 0 VSS
flabel metal4 39914 1890 39924 1898 1 FreeSans 480 0 0 0 venp1
flabel metal4 39912 5932 39922 5950 1 FreeSans 480 0 0 0 venm1
flabel metal4 39872 9472 39892 9486 1 FreeSans 480 0 0 0 vim2
flabel metal4 39942 13524 39962 13540 1 FreeSans 480 0 0 0 vip2
flabel metal4 40082 15590 40102 15606 1 FreeSans 480 0 0 0 venp2
flabel metal4 40024 19636 40048 19656 1 FreeSans 480 0 0 0 venm2
flabel metal4 40068 25698 40084 25712 1 FreeSans 480 0 0 0 vop
flabel metal4 49508 27900 49618 28008 1 FreeSans 480 0 0 0 VDD
flabel metal2 50956 4528 50982 4554 1 FreeSans 480 0 0 0 gain_ctrl_0
flabel metal2 49538 23440 49558 23458 1 FreeSans 480 0 0 0 gain_ctrl_1
flabel metal4 36296 7672 36328 7702 1 FreeSans 480 0 0 0 vocm
flabel metal1 3968 4954 3982 4962 1 FreeSans 480 0 0 0 ibiasn1
flabel metal1 57962 4966 57978 4972 1 FreeSans 480 0 0 0 ibiasn2
flabel metal1 -7768 15456 -7762 15460 1 FreeSans 480 0 0 0 rst_n
flabel metal1 -8136 15450 -8128 15458 1 FreeSans 480 0 0 0 rst
flabel metal3 -9694 13074 -9674 13090 1 FreeSans 480 0 0 0 vip1
flabel metal4 -9728 8802 -9684 8828 1 FreeSans 480 0 0 0 vop1
flabel metal4 -9734 12846 -9714 12872 1 FreeSans 480 0 0 0 vom1
flabel metal3 -9770 8556 -9744 8576 1 FreeSans 480 0 0 0 vim1
flabel metal3 -9338 5886 -9298 5918 1 FreeSans 480 0 0 0 vhpf
flabel metal3 -9718 1372 -9700 1386 1 FreeSans 480 0 0 0 vincm
flabel metal3 39912 1630 39926 1644 1 FreeSans 480 0 0 0 vop1
flabel metal3 39900 6144 39910 6156 1 FreeSans 480 0 0 0 vom1
flabel metal3 39848 9234 39866 9256 1 FreeSans 480 0 0 0 vop1
flabel metal3 39924 13774 39940 13786 1 FreeSans 480 0 0 0 vom1
flabel metal3 40106 19872 40122 19884 1 FreeSans 480 0 0 0 vip2
flabel metal3 40076 15316 40096 15328 1 FreeSans 480 0 0 0 vim2
flabel metal2 40896 23642 40916 23660 1 FreeSans 480 0 0 0 vim2
flabel metal4 39646 23514 39664 23536 1 FreeSans 480 0 0 0 vip2
flabel metal4 41878 23258 41900 23278 1 FreeSans 480 0 0 0 vom
<< end >>
