magic
tech sky130A
magscale 1 2
timestamp 1621035774
<< error_p >>
rect -1989 1950 -1929 3750
rect -1909 1950 -1849 3750
rect -70 1950 -10 3750
rect 10 1950 70 3750
rect 1849 1950 1909 3750
rect 1929 1950 1989 3750
rect -1989 50 -1929 1850
rect -1909 50 -1849 1850
rect -70 50 -10 1850
rect 10 50 70 1850
rect 1849 50 1909 1850
rect 1929 50 1989 1850
rect -1989 -1850 -1929 -50
rect -1909 -1850 -1849 -50
rect -70 -1850 -10 -50
rect 10 -1850 70 -50
rect 1849 -1850 1909 -50
rect 1929 -1850 1989 -50
rect -1989 -3750 -1929 -1950
rect -1909 -3750 -1849 -1950
rect -70 -3750 -10 -1950
rect 10 -3750 70 -1950
rect 1849 -3750 1909 -1950
rect 1929 -3750 1989 -1950
<< metal3 >>
rect -3828 3722 -1929 3750
rect -3828 1978 -2013 3722
rect -1949 1978 -1929 3722
rect -3828 1950 -1929 1978
rect -1909 3722 -10 3750
rect -1909 1978 -94 3722
rect -30 1978 -10 3722
rect -1909 1950 -10 1978
rect 10 3722 1909 3750
rect 10 1978 1825 3722
rect 1889 1978 1909 3722
rect 10 1950 1909 1978
rect 1929 3722 3828 3750
rect 1929 1978 3744 3722
rect 3808 1978 3828 3722
rect 1929 1950 3828 1978
rect -3828 1822 -1929 1850
rect -3828 78 -2013 1822
rect -1949 78 -1929 1822
rect -3828 50 -1929 78
rect -1909 1822 -10 1850
rect -1909 78 -94 1822
rect -30 78 -10 1822
rect -1909 50 -10 78
rect 10 1822 1909 1850
rect 10 78 1825 1822
rect 1889 78 1909 1822
rect 10 50 1909 78
rect 1929 1822 3828 1850
rect 1929 78 3744 1822
rect 3808 78 3828 1822
rect 1929 50 3828 78
rect -3828 -78 -1929 -50
rect -3828 -1822 -2013 -78
rect -1949 -1822 -1929 -78
rect -3828 -1850 -1929 -1822
rect -1909 -78 -10 -50
rect -1909 -1822 -94 -78
rect -30 -1822 -10 -78
rect -1909 -1850 -10 -1822
rect 10 -78 1909 -50
rect 10 -1822 1825 -78
rect 1889 -1822 1909 -78
rect 10 -1850 1909 -1822
rect 1929 -78 3828 -50
rect 1929 -1822 3744 -78
rect 3808 -1822 3828 -78
rect 1929 -1850 3828 -1822
rect -3828 -1978 -1929 -1950
rect -3828 -3722 -2013 -1978
rect -1949 -3722 -1929 -1978
rect -3828 -3750 -1929 -3722
rect -1909 -1978 -10 -1950
rect -1909 -3722 -94 -1978
rect -30 -3722 -10 -1978
rect -1909 -3750 -10 -3722
rect 10 -1978 1909 -1950
rect 10 -3722 1825 -1978
rect 1889 -3722 1909 -1978
rect 10 -3750 1909 -3722
rect 1929 -1978 3828 -1950
rect 1929 -3722 3744 -1978
rect 3808 -3722 3828 -1978
rect 1929 -3750 3828 -3722
<< via3 >>
rect -2013 1978 -1949 3722
rect -94 1978 -30 3722
rect 1825 1978 1889 3722
rect 3744 1978 3808 3722
rect -2013 78 -1949 1822
rect -94 78 -30 1822
rect 1825 78 1889 1822
rect 3744 78 3808 1822
rect -2013 -1822 -1949 -78
rect -94 -1822 -30 -78
rect 1825 -1822 1889 -78
rect 3744 -1822 3808 -78
rect -2013 -3722 -1949 -1978
rect -94 -3722 -30 -1978
rect 1825 -3722 1889 -1978
rect 3744 -3722 3808 -1978
<< mimcap >>
rect -3728 3610 -2128 3650
rect -3728 2090 -3688 3610
rect -2168 2090 -2128 3610
rect -3728 2050 -2128 2090
rect -1809 3610 -209 3650
rect -1809 2090 -1769 3610
rect -249 2090 -209 3610
rect -1809 2050 -209 2090
rect 110 3610 1710 3650
rect 110 2090 150 3610
rect 1670 2090 1710 3610
rect 110 2050 1710 2090
rect 2029 3610 3629 3650
rect 2029 2090 2069 3610
rect 3589 2090 3629 3610
rect 2029 2050 3629 2090
rect -3728 1710 -2128 1750
rect -3728 190 -3688 1710
rect -2168 190 -2128 1710
rect -3728 150 -2128 190
rect -1809 1710 -209 1750
rect -1809 190 -1769 1710
rect -249 190 -209 1710
rect -1809 150 -209 190
rect 110 1710 1710 1750
rect 110 190 150 1710
rect 1670 190 1710 1710
rect 110 150 1710 190
rect 2029 1710 3629 1750
rect 2029 190 2069 1710
rect 3589 190 3629 1710
rect 2029 150 3629 190
rect -3728 -190 -2128 -150
rect -3728 -1710 -3688 -190
rect -2168 -1710 -2128 -190
rect -3728 -1750 -2128 -1710
rect -1809 -190 -209 -150
rect -1809 -1710 -1769 -190
rect -249 -1710 -209 -190
rect -1809 -1750 -209 -1710
rect 110 -190 1710 -150
rect 110 -1710 150 -190
rect 1670 -1710 1710 -190
rect 110 -1750 1710 -1710
rect 2029 -190 3629 -150
rect 2029 -1710 2069 -190
rect 3589 -1710 3629 -190
rect 2029 -1750 3629 -1710
rect -3728 -2090 -2128 -2050
rect -3728 -3610 -3688 -2090
rect -2168 -3610 -2128 -2090
rect -3728 -3650 -2128 -3610
rect -1809 -2090 -209 -2050
rect -1809 -3610 -1769 -2090
rect -249 -3610 -209 -2090
rect -1809 -3650 -209 -3610
rect 110 -2090 1710 -2050
rect 110 -3610 150 -2090
rect 1670 -3610 1710 -2090
rect 110 -3650 1710 -3610
rect 2029 -2090 3629 -2050
rect 2029 -3610 2069 -2090
rect 3589 -3610 3629 -2090
rect 2029 -3650 3629 -3610
<< mimcapcontact >>
rect -3688 2090 -2168 3610
rect -1769 2090 -249 3610
rect 150 2090 1670 3610
rect 2069 2090 3589 3610
rect -3688 190 -2168 1710
rect -1769 190 -249 1710
rect 150 190 1670 1710
rect 2069 190 3589 1710
rect -3688 -1710 -2168 -190
rect -1769 -1710 -249 -190
rect 150 -1710 1670 -190
rect 2069 -1710 3589 -190
rect -3688 -3610 -2168 -2090
rect -1769 -3610 -249 -2090
rect 150 -3610 1670 -2090
rect 2069 -3610 3589 -2090
<< metal4 >>
rect -2980 3611 -2876 3800
rect -2060 3738 -1956 3800
rect -2060 3722 -1933 3738
rect -3689 3610 -2167 3611
rect -3689 2090 -3688 3610
rect -2168 2090 -2167 3610
rect -3689 2089 -2167 2090
rect -2980 1711 -2876 2089
rect -2060 1978 -2013 3722
rect -1949 1978 -1933 3722
rect -1061 3611 -957 3800
rect -141 3738 -37 3800
rect -141 3722 -14 3738
rect -1770 3610 -248 3611
rect -1770 2090 -1769 3610
rect -249 2090 -248 3610
rect -1770 2089 -248 2090
rect -2060 1962 -1933 1978
rect -2060 1838 -1956 1962
rect -2060 1822 -1933 1838
rect -3689 1710 -2167 1711
rect -3689 190 -3688 1710
rect -2168 190 -2167 1710
rect -3689 189 -2167 190
rect -2980 -189 -2876 189
rect -2060 78 -2013 1822
rect -1949 78 -1933 1822
rect -1061 1711 -957 2089
rect -141 1978 -94 3722
rect -30 1978 -14 3722
rect 858 3611 962 3800
rect 1778 3738 1882 3800
rect 1778 3722 1905 3738
rect 149 3610 1671 3611
rect 149 2090 150 3610
rect 1670 2090 1671 3610
rect 149 2089 1671 2090
rect -141 1962 -14 1978
rect -141 1838 -37 1962
rect -141 1822 -14 1838
rect -1770 1710 -248 1711
rect -1770 190 -1769 1710
rect -249 190 -248 1710
rect -1770 189 -248 190
rect -2060 62 -1933 78
rect -2060 -62 -1956 62
rect -2060 -78 -1933 -62
rect -3689 -190 -2167 -189
rect -3689 -1710 -3688 -190
rect -2168 -1710 -2167 -190
rect -3689 -1711 -2167 -1710
rect -2980 -2089 -2876 -1711
rect -2060 -1822 -2013 -78
rect -1949 -1822 -1933 -78
rect -1061 -189 -957 189
rect -141 78 -94 1822
rect -30 78 -14 1822
rect 858 1711 962 2089
rect 1778 1978 1825 3722
rect 1889 1978 1905 3722
rect 2777 3611 2881 3800
rect 3697 3738 3801 3800
rect 3697 3722 3824 3738
rect 2068 3610 3590 3611
rect 2068 2090 2069 3610
rect 3589 2090 3590 3610
rect 2068 2089 3590 2090
rect 1778 1962 1905 1978
rect 1778 1838 1882 1962
rect 1778 1822 1905 1838
rect 149 1710 1671 1711
rect 149 190 150 1710
rect 1670 190 1671 1710
rect 149 189 1671 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -1770 -190 -248 -189
rect -1770 -1710 -1769 -190
rect -249 -1710 -248 -190
rect -1770 -1711 -248 -1710
rect -2060 -1838 -1933 -1822
rect -2060 -1962 -1956 -1838
rect -2060 -1978 -1933 -1962
rect -3689 -2090 -2167 -2089
rect -3689 -3610 -3688 -2090
rect -2168 -3610 -2167 -2090
rect -3689 -3611 -2167 -3610
rect -2980 -3800 -2876 -3611
rect -2060 -3722 -2013 -1978
rect -1949 -3722 -1933 -1978
rect -1061 -2089 -957 -1711
rect -141 -1822 -94 -78
rect -30 -1822 -14 -78
rect 858 -189 962 189
rect 1778 78 1825 1822
rect 1889 78 1905 1822
rect 2777 1711 2881 2089
rect 3697 1978 3744 3722
rect 3808 1978 3824 3722
rect 3697 1962 3824 1978
rect 3697 1838 3801 1962
rect 3697 1822 3824 1838
rect 2068 1710 3590 1711
rect 2068 190 2069 1710
rect 3589 190 3590 1710
rect 2068 189 3590 190
rect 1778 62 1905 78
rect 1778 -62 1882 62
rect 1778 -78 1905 -62
rect 149 -190 1671 -189
rect 149 -1710 150 -190
rect 1670 -1710 1671 -190
rect 149 -1711 1671 -1710
rect -141 -1838 -14 -1822
rect -141 -1962 -37 -1838
rect -141 -1978 -14 -1962
rect -1770 -2090 -248 -2089
rect -1770 -3610 -1769 -2090
rect -249 -3610 -248 -2090
rect -1770 -3611 -248 -3610
rect -2060 -3738 -1933 -3722
rect -2060 -3800 -1956 -3738
rect -1061 -3800 -957 -3611
rect -141 -3722 -94 -1978
rect -30 -3722 -14 -1978
rect 858 -2089 962 -1711
rect 1778 -1822 1825 -78
rect 1889 -1822 1905 -78
rect 2777 -189 2881 189
rect 3697 78 3744 1822
rect 3808 78 3824 1822
rect 3697 62 3824 78
rect 3697 -62 3801 62
rect 3697 -78 3824 -62
rect 2068 -190 3590 -189
rect 2068 -1710 2069 -190
rect 3589 -1710 3590 -190
rect 2068 -1711 3590 -1710
rect 1778 -1838 1905 -1822
rect 1778 -1962 1882 -1838
rect 1778 -1978 1905 -1962
rect 149 -2090 1671 -2089
rect 149 -3610 150 -2090
rect 1670 -3610 1671 -2090
rect 149 -3611 1671 -3610
rect -141 -3738 -14 -3722
rect -141 -3800 -37 -3738
rect 858 -3800 962 -3611
rect 1778 -3722 1825 -1978
rect 1889 -3722 1905 -1978
rect 2777 -2089 2881 -1711
rect 3697 -1822 3744 -78
rect 3808 -1822 3824 -78
rect 3697 -1838 3824 -1822
rect 3697 -1962 3801 -1838
rect 3697 -1978 3824 -1962
rect 2068 -2090 3590 -2089
rect 2068 -3610 2069 -2090
rect 3589 -3610 3590 -2090
rect 2068 -3611 3590 -3610
rect 1778 -3738 1905 -3722
rect 1778 -3800 1882 -3738
rect 2777 -3800 2881 -3611
rect 3697 -3722 3744 -1978
rect 3808 -3722 3824 -1978
rect 3697 -3738 3824 -3722
rect 3697 -3800 3801 -3738
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 1929 1950 3729 3750
string parameters w 8.00 l 8.00 val 134.08 carea 2.00 cperi 0.19 nx 4 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
