magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -5447 -2160 5447 2160
<< nwell >>
rect -4187 -900 4187 900
<< pmoshvt >>
rect -4093 -800 -3693 800
rect -3635 -800 -3235 800
rect -3177 -800 -2777 800
rect -2719 -800 -2319 800
rect -2261 -800 -1861 800
rect -1803 -800 -1403 800
rect -1345 -800 -945 800
rect -887 -800 -487 800
rect -429 -800 -29 800
rect 29 -800 429 800
rect 487 -800 887 800
rect 945 -800 1345 800
rect 1403 -800 1803 800
rect 1861 -800 2261 800
rect 2319 -800 2719 800
rect 2777 -800 3177 800
rect 3235 -800 3635 800
rect 3693 -800 4093 800
<< pdiff >>
rect -4151 765 -4093 800
rect -4151 731 -4139 765
rect -4105 731 -4093 765
rect -4151 697 -4093 731
rect -4151 663 -4139 697
rect -4105 663 -4093 697
rect -4151 629 -4093 663
rect -4151 595 -4139 629
rect -4105 595 -4093 629
rect -4151 561 -4093 595
rect -4151 527 -4139 561
rect -4105 527 -4093 561
rect -4151 493 -4093 527
rect -4151 459 -4139 493
rect -4105 459 -4093 493
rect -4151 425 -4093 459
rect -4151 391 -4139 425
rect -4105 391 -4093 425
rect -4151 357 -4093 391
rect -4151 323 -4139 357
rect -4105 323 -4093 357
rect -4151 289 -4093 323
rect -4151 255 -4139 289
rect -4105 255 -4093 289
rect -4151 221 -4093 255
rect -4151 187 -4139 221
rect -4105 187 -4093 221
rect -4151 153 -4093 187
rect -4151 119 -4139 153
rect -4105 119 -4093 153
rect -4151 85 -4093 119
rect -4151 51 -4139 85
rect -4105 51 -4093 85
rect -4151 17 -4093 51
rect -4151 -17 -4139 17
rect -4105 -17 -4093 17
rect -4151 -51 -4093 -17
rect -4151 -85 -4139 -51
rect -4105 -85 -4093 -51
rect -4151 -119 -4093 -85
rect -4151 -153 -4139 -119
rect -4105 -153 -4093 -119
rect -4151 -187 -4093 -153
rect -4151 -221 -4139 -187
rect -4105 -221 -4093 -187
rect -4151 -255 -4093 -221
rect -4151 -289 -4139 -255
rect -4105 -289 -4093 -255
rect -4151 -323 -4093 -289
rect -4151 -357 -4139 -323
rect -4105 -357 -4093 -323
rect -4151 -391 -4093 -357
rect -4151 -425 -4139 -391
rect -4105 -425 -4093 -391
rect -4151 -459 -4093 -425
rect -4151 -493 -4139 -459
rect -4105 -493 -4093 -459
rect -4151 -527 -4093 -493
rect -4151 -561 -4139 -527
rect -4105 -561 -4093 -527
rect -4151 -595 -4093 -561
rect -4151 -629 -4139 -595
rect -4105 -629 -4093 -595
rect -4151 -663 -4093 -629
rect -4151 -697 -4139 -663
rect -4105 -697 -4093 -663
rect -4151 -731 -4093 -697
rect -4151 -765 -4139 -731
rect -4105 -765 -4093 -731
rect -4151 -800 -4093 -765
rect -3693 765 -3635 800
rect -3693 731 -3681 765
rect -3647 731 -3635 765
rect -3693 697 -3635 731
rect -3693 663 -3681 697
rect -3647 663 -3635 697
rect -3693 629 -3635 663
rect -3693 595 -3681 629
rect -3647 595 -3635 629
rect -3693 561 -3635 595
rect -3693 527 -3681 561
rect -3647 527 -3635 561
rect -3693 493 -3635 527
rect -3693 459 -3681 493
rect -3647 459 -3635 493
rect -3693 425 -3635 459
rect -3693 391 -3681 425
rect -3647 391 -3635 425
rect -3693 357 -3635 391
rect -3693 323 -3681 357
rect -3647 323 -3635 357
rect -3693 289 -3635 323
rect -3693 255 -3681 289
rect -3647 255 -3635 289
rect -3693 221 -3635 255
rect -3693 187 -3681 221
rect -3647 187 -3635 221
rect -3693 153 -3635 187
rect -3693 119 -3681 153
rect -3647 119 -3635 153
rect -3693 85 -3635 119
rect -3693 51 -3681 85
rect -3647 51 -3635 85
rect -3693 17 -3635 51
rect -3693 -17 -3681 17
rect -3647 -17 -3635 17
rect -3693 -51 -3635 -17
rect -3693 -85 -3681 -51
rect -3647 -85 -3635 -51
rect -3693 -119 -3635 -85
rect -3693 -153 -3681 -119
rect -3647 -153 -3635 -119
rect -3693 -187 -3635 -153
rect -3693 -221 -3681 -187
rect -3647 -221 -3635 -187
rect -3693 -255 -3635 -221
rect -3693 -289 -3681 -255
rect -3647 -289 -3635 -255
rect -3693 -323 -3635 -289
rect -3693 -357 -3681 -323
rect -3647 -357 -3635 -323
rect -3693 -391 -3635 -357
rect -3693 -425 -3681 -391
rect -3647 -425 -3635 -391
rect -3693 -459 -3635 -425
rect -3693 -493 -3681 -459
rect -3647 -493 -3635 -459
rect -3693 -527 -3635 -493
rect -3693 -561 -3681 -527
rect -3647 -561 -3635 -527
rect -3693 -595 -3635 -561
rect -3693 -629 -3681 -595
rect -3647 -629 -3635 -595
rect -3693 -663 -3635 -629
rect -3693 -697 -3681 -663
rect -3647 -697 -3635 -663
rect -3693 -731 -3635 -697
rect -3693 -765 -3681 -731
rect -3647 -765 -3635 -731
rect -3693 -800 -3635 -765
rect -3235 765 -3177 800
rect -3235 731 -3223 765
rect -3189 731 -3177 765
rect -3235 697 -3177 731
rect -3235 663 -3223 697
rect -3189 663 -3177 697
rect -3235 629 -3177 663
rect -3235 595 -3223 629
rect -3189 595 -3177 629
rect -3235 561 -3177 595
rect -3235 527 -3223 561
rect -3189 527 -3177 561
rect -3235 493 -3177 527
rect -3235 459 -3223 493
rect -3189 459 -3177 493
rect -3235 425 -3177 459
rect -3235 391 -3223 425
rect -3189 391 -3177 425
rect -3235 357 -3177 391
rect -3235 323 -3223 357
rect -3189 323 -3177 357
rect -3235 289 -3177 323
rect -3235 255 -3223 289
rect -3189 255 -3177 289
rect -3235 221 -3177 255
rect -3235 187 -3223 221
rect -3189 187 -3177 221
rect -3235 153 -3177 187
rect -3235 119 -3223 153
rect -3189 119 -3177 153
rect -3235 85 -3177 119
rect -3235 51 -3223 85
rect -3189 51 -3177 85
rect -3235 17 -3177 51
rect -3235 -17 -3223 17
rect -3189 -17 -3177 17
rect -3235 -51 -3177 -17
rect -3235 -85 -3223 -51
rect -3189 -85 -3177 -51
rect -3235 -119 -3177 -85
rect -3235 -153 -3223 -119
rect -3189 -153 -3177 -119
rect -3235 -187 -3177 -153
rect -3235 -221 -3223 -187
rect -3189 -221 -3177 -187
rect -3235 -255 -3177 -221
rect -3235 -289 -3223 -255
rect -3189 -289 -3177 -255
rect -3235 -323 -3177 -289
rect -3235 -357 -3223 -323
rect -3189 -357 -3177 -323
rect -3235 -391 -3177 -357
rect -3235 -425 -3223 -391
rect -3189 -425 -3177 -391
rect -3235 -459 -3177 -425
rect -3235 -493 -3223 -459
rect -3189 -493 -3177 -459
rect -3235 -527 -3177 -493
rect -3235 -561 -3223 -527
rect -3189 -561 -3177 -527
rect -3235 -595 -3177 -561
rect -3235 -629 -3223 -595
rect -3189 -629 -3177 -595
rect -3235 -663 -3177 -629
rect -3235 -697 -3223 -663
rect -3189 -697 -3177 -663
rect -3235 -731 -3177 -697
rect -3235 -765 -3223 -731
rect -3189 -765 -3177 -731
rect -3235 -800 -3177 -765
rect -2777 765 -2719 800
rect -2777 731 -2765 765
rect -2731 731 -2719 765
rect -2777 697 -2719 731
rect -2777 663 -2765 697
rect -2731 663 -2719 697
rect -2777 629 -2719 663
rect -2777 595 -2765 629
rect -2731 595 -2719 629
rect -2777 561 -2719 595
rect -2777 527 -2765 561
rect -2731 527 -2719 561
rect -2777 493 -2719 527
rect -2777 459 -2765 493
rect -2731 459 -2719 493
rect -2777 425 -2719 459
rect -2777 391 -2765 425
rect -2731 391 -2719 425
rect -2777 357 -2719 391
rect -2777 323 -2765 357
rect -2731 323 -2719 357
rect -2777 289 -2719 323
rect -2777 255 -2765 289
rect -2731 255 -2719 289
rect -2777 221 -2719 255
rect -2777 187 -2765 221
rect -2731 187 -2719 221
rect -2777 153 -2719 187
rect -2777 119 -2765 153
rect -2731 119 -2719 153
rect -2777 85 -2719 119
rect -2777 51 -2765 85
rect -2731 51 -2719 85
rect -2777 17 -2719 51
rect -2777 -17 -2765 17
rect -2731 -17 -2719 17
rect -2777 -51 -2719 -17
rect -2777 -85 -2765 -51
rect -2731 -85 -2719 -51
rect -2777 -119 -2719 -85
rect -2777 -153 -2765 -119
rect -2731 -153 -2719 -119
rect -2777 -187 -2719 -153
rect -2777 -221 -2765 -187
rect -2731 -221 -2719 -187
rect -2777 -255 -2719 -221
rect -2777 -289 -2765 -255
rect -2731 -289 -2719 -255
rect -2777 -323 -2719 -289
rect -2777 -357 -2765 -323
rect -2731 -357 -2719 -323
rect -2777 -391 -2719 -357
rect -2777 -425 -2765 -391
rect -2731 -425 -2719 -391
rect -2777 -459 -2719 -425
rect -2777 -493 -2765 -459
rect -2731 -493 -2719 -459
rect -2777 -527 -2719 -493
rect -2777 -561 -2765 -527
rect -2731 -561 -2719 -527
rect -2777 -595 -2719 -561
rect -2777 -629 -2765 -595
rect -2731 -629 -2719 -595
rect -2777 -663 -2719 -629
rect -2777 -697 -2765 -663
rect -2731 -697 -2719 -663
rect -2777 -731 -2719 -697
rect -2777 -765 -2765 -731
rect -2731 -765 -2719 -731
rect -2777 -800 -2719 -765
rect -2319 765 -2261 800
rect -2319 731 -2307 765
rect -2273 731 -2261 765
rect -2319 697 -2261 731
rect -2319 663 -2307 697
rect -2273 663 -2261 697
rect -2319 629 -2261 663
rect -2319 595 -2307 629
rect -2273 595 -2261 629
rect -2319 561 -2261 595
rect -2319 527 -2307 561
rect -2273 527 -2261 561
rect -2319 493 -2261 527
rect -2319 459 -2307 493
rect -2273 459 -2261 493
rect -2319 425 -2261 459
rect -2319 391 -2307 425
rect -2273 391 -2261 425
rect -2319 357 -2261 391
rect -2319 323 -2307 357
rect -2273 323 -2261 357
rect -2319 289 -2261 323
rect -2319 255 -2307 289
rect -2273 255 -2261 289
rect -2319 221 -2261 255
rect -2319 187 -2307 221
rect -2273 187 -2261 221
rect -2319 153 -2261 187
rect -2319 119 -2307 153
rect -2273 119 -2261 153
rect -2319 85 -2261 119
rect -2319 51 -2307 85
rect -2273 51 -2261 85
rect -2319 17 -2261 51
rect -2319 -17 -2307 17
rect -2273 -17 -2261 17
rect -2319 -51 -2261 -17
rect -2319 -85 -2307 -51
rect -2273 -85 -2261 -51
rect -2319 -119 -2261 -85
rect -2319 -153 -2307 -119
rect -2273 -153 -2261 -119
rect -2319 -187 -2261 -153
rect -2319 -221 -2307 -187
rect -2273 -221 -2261 -187
rect -2319 -255 -2261 -221
rect -2319 -289 -2307 -255
rect -2273 -289 -2261 -255
rect -2319 -323 -2261 -289
rect -2319 -357 -2307 -323
rect -2273 -357 -2261 -323
rect -2319 -391 -2261 -357
rect -2319 -425 -2307 -391
rect -2273 -425 -2261 -391
rect -2319 -459 -2261 -425
rect -2319 -493 -2307 -459
rect -2273 -493 -2261 -459
rect -2319 -527 -2261 -493
rect -2319 -561 -2307 -527
rect -2273 -561 -2261 -527
rect -2319 -595 -2261 -561
rect -2319 -629 -2307 -595
rect -2273 -629 -2261 -595
rect -2319 -663 -2261 -629
rect -2319 -697 -2307 -663
rect -2273 -697 -2261 -663
rect -2319 -731 -2261 -697
rect -2319 -765 -2307 -731
rect -2273 -765 -2261 -731
rect -2319 -800 -2261 -765
rect -1861 765 -1803 800
rect -1861 731 -1849 765
rect -1815 731 -1803 765
rect -1861 697 -1803 731
rect -1861 663 -1849 697
rect -1815 663 -1803 697
rect -1861 629 -1803 663
rect -1861 595 -1849 629
rect -1815 595 -1803 629
rect -1861 561 -1803 595
rect -1861 527 -1849 561
rect -1815 527 -1803 561
rect -1861 493 -1803 527
rect -1861 459 -1849 493
rect -1815 459 -1803 493
rect -1861 425 -1803 459
rect -1861 391 -1849 425
rect -1815 391 -1803 425
rect -1861 357 -1803 391
rect -1861 323 -1849 357
rect -1815 323 -1803 357
rect -1861 289 -1803 323
rect -1861 255 -1849 289
rect -1815 255 -1803 289
rect -1861 221 -1803 255
rect -1861 187 -1849 221
rect -1815 187 -1803 221
rect -1861 153 -1803 187
rect -1861 119 -1849 153
rect -1815 119 -1803 153
rect -1861 85 -1803 119
rect -1861 51 -1849 85
rect -1815 51 -1803 85
rect -1861 17 -1803 51
rect -1861 -17 -1849 17
rect -1815 -17 -1803 17
rect -1861 -51 -1803 -17
rect -1861 -85 -1849 -51
rect -1815 -85 -1803 -51
rect -1861 -119 -1803 -85
rect -1861 -153 -1849 -119
rect -1815 -153 -1803 -119
rect -1861 -187 -1803 -153
rect -1861 -221 -1849 -187
rect -1815 -221 -1803 -187
rect -1861 -255 -1803 -221
rect -1861 -289 -1849 -255
rect -1815 -289 -1803 -255
rect -1861 -323 -1803 -289
rect -1861 -357 -1849 -323
rect -1815 -357 -1803 -323
rect -1861 -391 -1803 -357
rect -1861 -425 -1849 -391
rect -1815 -425 -1803 -391
rect -1861 -459 -1803 -425
rect -1861 -493 -1849 -459
rect -1815 -493 -1803 -459
rect -1861 -527 -1803 -493
rect -1861 -561 -1849 -527
rect -1815 -561 -1803 -527
rect -1861 -595 -1803 -561
rect -1861 -629 -1849 -595
rect -1815 -629 -1803 -595
rect -1861 -663 -1803 -629
rect -1861 -697 -1849 -663
rect -1815 -697 -1803 -663
rect -1861 -731 -1803 -697
rect -1861 -765 -1849 -731
rect -1815 -765 -1803 -731
rect -1861 -800 -1803 -765
rect -1403 765 -1345 800
rect -1403 731 -1391 765
rect -1357 731 -1345 765
rect -1403 697 -1345 731
rect -1403 663 -1391 697
rect -1357 663 -1345 697
rect -1403 629 -1345 663
rect -1403 595 -1391 629
rect -1357 595 -1345 629
rect -1403 561 -1345 595
rect -1403 527 -1391 561
rect -1357 527 -1345 561
rect -1403 493 -1345 527
rect -1403 459 -1391 493
rect -1357 459 -1345 493
rect -1403 425 -1345 459
rect -1403 391 -1391 425
rect -1357 391 -1345 425
rect -1403 357 -1345 391
rect -1403 323 -1391 357
rect -1357 323 -1345 357
rect -1403 289 -1345 323
rect -1403 255 -1391 289
rect -1357 255 -1345 289
rect -1403 221 -1345 255
rect -1403 187 -1391 221
rect -1357 187 -1345 221
rect -1403 153 -1345 187
rect -1403 119 -1391 153
rect -1357 119 -1345 153
rect -1403 85 -1345 119
rect -1403 51 -1391 85
rect -1357 51 -1345 85
rect -1403 17 -1345 51
rect -1403 -17 -1391 17
rect -1357 -17 -1345 17
rect -1403 -51 -1345 -17
rect -1403 -85 -1391 -51
rect -1357 -85 -1345 -51
rect -1403 -119 -1345 -85
rect -1403 -153 -1391 -119
rect -1357 -153 -1345 -119
rect -1403 -187 -1345 -153
rect -1403 -221 -1391 -187
rect -1357 -221 -1345 -187
rect -1403 -255 -1345 -221
rect -1403 -289 -1391 -255
rect -1357 -289 -1345 -255
rect -1403 -323 -1345 -289
rect -1403 -357 -1391 -323
rect -1357 -357 -1345 -323
rect -1403 -391 -1345 -357
rect -1403 -425 -1391 -391
rect -1357 -425 -1345 -391
rect -1403 -459 -1345 -425
rect -1403 -493 -1391 -459
rect -1357 -493 -1345 -459
rect -1403 -527 -1345 -493
rect -1403 -561 -1391 -527
rect -1357 -561 -1345 -527
rect -1403 -595 -1345 -561
rect -1403 -629 -1391 -595
rect -1357 -629 -1345 -595
rect -1403 -663 -1345 -629
rect -1403 -697 -1391 -663
rect -1357 -697 -1345 -663
rect -1403 -731 -1345 -697
rect -1403 -765 -1391 -731
rect -1357 -765 -1345 -731
rect -1403 -800 -1345 -765
rect -945 765 -887 800
rect -945 731 -933 765
rect -899 731 -887 765
rect -945 697 -887 731
rect -945 663 -933 697
rect -899 663 -887 697
rect -945 629 -887 663
rect -945 595 -933 629
rect -899 595 -887 629
rect -945 561 -887 595
rect -945 527 -933 561
rect -899 527 -887 561
rect -945 493 -887 527
rect -945 459 -933 493
rect -899 459 -887 493
rect -945 425 -887 459
rect -945 391 -933 425
rect -899 391 -887 425
rect -945 357 -887 391
rect -945 323 -933 357
rect -899 323 -887 357
rect -945 289 -887 323
rect -945 255 -933 289
rect -899 255 -887 289
rect -945 221 -887 255
rect -945 187 -933 221
rect -899 187 -887 221
rect -945 153 -887 187
rect -945 119 -933 153
rect -899 119 -887 153
rect -945 85 -887 119
rect -945 51 -933 85
rect -899 51 -887 85
rect -945 17 -887 51
rect -945 -17 -933 17
rect -899 -17 -887 17
rect -945 -51 -887 -17
rect -945 -85 -933 -51
rect -899 -85 -887 -51
rect -945 -119 -887 -85
rect -945 -153 -933 -119
rect -899 -153 -887 -119
rect -945 -187 -887 -153
rect -945 -221 -933 -187
rect -899 -221 -887 -187
rect -945 -255 -887 -221
rect -945 -289 -933 -255
rect -899 -289 -887 -255
rect -945 -323 -887 -289
rect -945 -357 -933 -323
rect -899 -357 -887 -323
rect -945 -391 -887 -357
rect -945 -425 -933 -391
rect -899 -425 -887 -391
rect -945 -459 -887 -425
rect -945 -493 -933 -459
rect -899 -493 -887 -459
rect -945 -527 -887 -493
rect -945 -561 -933 -527
rect -899 -561 -887 -527
rect -945 -595 -887 -561
rect -945 -629 -933 -595
rect -899 -629 -887 -595
rect -945 -663 -887 -629
rect -945 -697 -933 -663
rect -899 -697 -887 -663
rect -945 -731 -887 -697
rect -945 -765 -933 -731
rect -899 -765 -887 -731
rect -945 -800 -887 -765
rect -487 765 -429 800
rect -487 731 -475 765
rect -441 731 -429 765
rect -487 697 -429 731
rect -487 663 -475 697
rect -441 663 -429 697
rect -487 629 -429 663
rect -487 595 -475 629
rect -441 595 -429 629
rect -487 561 -429 595
rect -487 527 -475 561
rect -441 527 -429 561
rect -487 493 -429 527
rect -487 459 -475 493
rect -441 459 -429 493
rect -487 425 -429 459
rect -487 391 -475 425
rect -441 391 -429 425
rect -487 357 -429 391
rect -487 323 -475 357
rect -441 323 -429 357
rect -487 289 -429 323
rect -487 255 -475 289
rect -441 255 -429 289
rect -487 221 -429 255
rect -487 187 -475 221
rect -441 187 -429 221
rect -487 153 -429 187
rect -487 119 -475 153
rect -441 119 -429 153
rect -487 85 -429 119
rect -487 51 -475 85
rect -441 51 -429 85
rect -487 17 -429 51
rect -487 -17 -475 17
rect -441 -17 -429 17
rect -487 -51 -429 -17
rect -487 -85 -475 -51
rect -441 -85 -429 -51
rect -487 -119 -429 -85
rect -487 -153 -475 -119
rect -441 -153 -429 -119
rect -487 -187 -429 -153
rect -487 -221 -475 -187
rect -441 -221 -429 -187
rect -487 -255 -429 -221
rect -487 -289 -475 -255
rect -441 -289 -429 -255
rect -487 -323 -429 -289
rect -487 -357 -475 -323
rect -441 -357 -429 -323
rect -487 -391 -429 -357
rect -487 -425 -475 -391
rect -441 -425 -429 -391
rect -487 -459 -429 -425
rect -487 -493 -475 -459
rect -441 -493 -429 -459
rect -487 -527 -429 -493
rect -487 -561 -475 -527
rect -441 -561 -429 -527
rect -487 -595 -429 -561
rect -487 -629 -475 -595
rect -441 -629 -429 -595
rect -487 -663 -429 -629
rect -487 -697 -475 -663
rect -441 -697 -429 -663
rect -487 -731 -429 -697
rect -487 -765 -475 -731
rect -441 -765 -429 -731
rect -487 -800 -429 -765
rect -29 765 29 800
rect -29 731 -17 765
rect 17 731 29 765
rect -29 697 29 731
rect -29 663 -17 697
rect 17 663 29 697
rect -29 629 29 663
rect -29 595 -17 629
rect 17 595 29 629
rect -29 561 29 595
rect -29 527 -17 561
rect 17 527 29 561
rect -29 493 29 527
rect -29 459 -17 493
rect 17 459 29 493
rect -29 425 29 459
rect -29 391 -17 425
rect 17 391 29 425
rect -29 357 29 391
rect -29 323 -17 357
rect 17 323 29 357
rect -29 289 29 323
rect -29 255 -17 289
rect 17 255 29 289
rect -29 221 29 255
rect -29 187 -17 221
rect 17 187 29 221
rect -29 153 29 187
rect -29 119 -17 153
rect 17 119 29 153
rect -29 85 29 119
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -119 29 -85
rect -29 -153 -17 -119
rect 17 -153 29 -119
rect -29 -187 29 -153
rect -29 -221 -17 -187
rect 17 -221 29 -187
rect -29 -255 29 -221
rect -29 -289 -17 -255
rect 17 -289 29 -255
rect -29 -323 29 -289
rect -29 -357 -17 -323
rect 17 -357 29 -323
rect -29 -391 29 -357
rect -29 -425 -17 -391
rect 17 -425 29 -391
rect -29 -459 29 -425
rect -29 -493 -17 -459
rect 17 -493 29 -459
rect -29 -527 29 -493
rect -29 -561 -17 -527
rect 17 -561 29 -527
rect -29 -595 29 -561
rect -29 -629 -17 -595
rect 17 -629 29 -595
rect -29 -663 29 -629
rect -29 -697 -17 -663
rect 17 -697 29 -663
rect -29 -731 29 -697
rect -29 -765 -17 -731
rect 17 -765 29 -731
rect -29 -800 29 -765
rect 429 765 487 800
rect 429 731 441 765
rect 475 731 487 765
rect 429 697 487 731
rect 429 663 441 697
rect 475 663 487 697
rect 429 629 487 663
rect 429 595 441 629
rect 475 595 487 629
rect 429 561 487 595
rect 429 527 441 561
rect 475 527 487 561
rect 429 493 487 527
rect 429 459 441 493
rect 475 459 487 493
rect 429 425 487 459
rect 429 391 441 425
rect 475 391 487 425
rect 429 357 487 391
rect 429 323 441 357
rect 475 323 487 357
rect 429 289 487 323
rect 429 255 441 289
rect 475 255 487 289
rect 429 221 487 255
rect 429 187 441 221
rect 475 187 487 221
rect 429 153 487 187
rect 429 119 441 153
rect 475 119 487 153
rect 429 85 487 119
rect 429 51 441 85
rect 475 51 487 85
rect 429 17 487 51
rect 429 -17 441 17
rect 475 -17 487 17
rect 429 -51 487 -17
rect 429 -85 441 -51
rect 475 -85 487 -51
rect 429 -119 487 -85
rect 429 -153 441 -119
rect 475 -153 487 -119
rect 429 -187 487 -153
rect 429 -221 441 -187
rect 475 -221 487 -187
rect 429 -255 487 -221
rect 429 -289 441 -255
rect 475 -289 487 -255
rect 429 -323 487 -289
rect 429 -357 441 -323
rect 475 -357 487 -323
rect 429 -391 487 -357
rect 429 -425 441 -391
rect 475 -425 487 -391
rect 429 -459 487 -425
rect 429 -493 441 -459
rect 475 -493 487 -459
rect 429 -527 487 -493
rect 429 -561 441 -527
rect 475 -561 487 -527
rect 429 -595 487 -561
rect 429 -629 441 -595
rect 475 -629 487 -595
rect 429 -663 487 -629
rect 429 -697 441 -663
rect 475 -697 487 -663
rect 429 -731 487 -697
rect 429 -765 441 -731
rect 475 -765 487 -731
rect 429 -800 487 -765
rect 887 765 945 800
rect 887 731 899 765
rect 933 731 945 765
rect 887 697 945 731
rect 887 663 899 697
rect 933 663 945 697
rect 887 629 945 663
rect 887 595 899 629
rect 933 595 945 629
rect 887 561 945 595
rect 887 527 899 561
rect 933 527 945 561
rect 887 493 945 527
rect 887 459 899 493
rect 933 459 945 493
rect 887 425 945 459
rect 887 391 899 425
rect 933 391 945 425
rect 887 357 945 391
rect 887 323 899 357
rect 933 323 945 357
rect 887 289 945 323
rect 887 255 899 289
rect 933 255 945 289
rect 887 221 945 255
rect 887 187 899 221
rect 933 187 945 221
rect 887 153 945 187
rect 887 119 899 153
rect 933 119 945 153
rect 887 85 945 119
rect 887 51 899 85
rect 933 51 945 85
rect 887 17 945 51
rect 887 -17 899 17
rect 933 -17 945 17
rect 887 -51 945 -17
rect 887 -85 899 -51
rect 933 -85 945 -51
rect 887 -119 945 -85
rect 887 -153 899 -119
rect 933 -153 945 -119
rect 887 -187 945 -153
rect 887 -221 899 -187
rect 933 -221 945 -187
rect 887 -255 945 -221
rect 887 -289 899 -255
rect 933 -289 945 -255
rect 887 -323 945 -289
rect 887 -357 899 -323
rect 933 -357 945 -323
rect 887 -391 945 -357
rect 887 -425 899 -391
rect 933 -425 945 -391
rect 887 -459 945 -425
rect 887 -493 899 -459
rect 933 -493 945 -459
rect 887 -527 945 -493
rect 887 -561 899 -527
rect 933 -561 945 -527
rect 887 -595 945 -561
rect 887 -629 899 -595
rect 933 -629 945 -595
rect 887 -663 945 -629
rect 887 -697 899 -663
rect 933 -697 945 -663
rect 887 -731 945 -697
rect 887 -765 899 -731
rect 933 -765 945 -731
rect 887 -800 945 -765
rect 1345 765 1403 800
rect 1345 731 1357 765
rect 1391 731 1403 765
rect 1345 697 1403 731
rect 1345 663 1357 697
rect 1391 663 1403 697
rect 1345 629 1403 663
rect 1345 595 1357 629
rect 1391 595 1403 629
rect 1345 561 1403 595
rect 1345 527 1357 561
rect 1391 527 1403 561
rect 1345 493 1403 527
rect 1345 459 1357 493
rect 1391 459 1403 493
rect 1345 425 1403 459
rect 1345 391 1357 425
rect 1391 391 1403 425
rect 1345 357 1403 391
rect 1345 323 1357 357
rect 1391 323 1403 357
rect 1345 289 1403 323
rect 1345 255 1357 289
rect 1391 255 1403 289
rect 1345 221 1403 255
rect 1345 187 1357 221
rect 1391 187 1403 221
rect 1345 153 1403 187
rect 1345 119 1357 153
rect 1391 119 1403 153
rect 1345 85 1403 119
rect 1345 51 1357 85
rect 1391 51 1403 85
rect 1345 17 1403 51
rect 1345 -17 1357 17
rect 1391 -17 1403 17
rect 1345 -51 1403 -17
rect 1345 -85 1357 -51
rect 1391 -85 1403 -51
rect 1345 -119 1403 -85
rect 1345 -153 1357 -119
rect 1391 -153 1403 -119
rect 1345 -187 1403 -153
rect 1345 -221 1357 -187
rect 1391 -221 1403 -187
rect 1345 -255 1403 -221
rect 1345 -289 1357 -255
rect 1391 -289 1403 -255
rect 1345 -323 1403 -289
rect 1345 -357 1357 -323
rect 1391 -357 1403 -323
rect 1345 -391 1403 -357
rect 1345 -425 1357 -391
rect 1391 -425 1403 -391
rect 1345 -459 1403 -425
rect 1345 -493 1357 -459
rect 1391 -493 1403 -459
rect 1345 -527 1403 -493
rect 1345 -561 1357 -527
rect 1391 -561 1403 -527
rect 1345 -595 1403 -561
rect 1345 -629 1357 -595
rect 1391 -629 1403 -595
rect 1345 -663 1403 -629
rect 1345 -697 1357 -663
rect 1391 -697 1403 -663
rect 1345 -731 1403 -697
rect 1345 -765 1357 -731
rect 1391 -765 1403 -731
rect 1345 -800 1403 -765
rect 1803 765 1861 800
rect 1803 731 1815 765
rect 1849 731 1861 765
rect 1803 697 1861 731
rect 1803 663 1815 697
rect 1849 663 1861 697
rect 1803 629 1861 663
rect 1803 595 1815 629
rect 1849 595 1861 629
rect 1803 561 1861 595
rect 1803 527 1815 561
rect 1849 527 1861 561
rect 1803 493 1861 527
rect 1803 459 1815 493
rect 1849 459 1861 493
rect 1803 425 1861 459
rect 1803 391 1815 425
rect 1849 391 1861 425
rect 1803 357 1861 391
rect 1803 323 1815 357
rect 1849 323 1861 357
rect 1803 289 1861 323
rect 1803 255 1815 289
rect 1849 255 1861 289
rect 1803 221 1861 255
rect 1803 187 1815 221
rect 1849 187 1861 221
rect 1803 153 1861 187
rect 1803 119 1815 153
rect 1849 119 1861 153
rect 1803 85 1861 119
rect 1803 51 1815 85
rect 1849 51 1861 85
rect 1803 17 1861 51
rect 1803 -17 1815 17
rect 1849 -17 1861 17
rect 1803 -51 1861 -17
rect 1803 -85 1815 -51
rect 1849 -85 1861 -51
rect 1803 -119 1861 -85
rect 1803 -153 1815 -119
rect 1849 -153 1861 -119
rect 1803 -187 1861 -153
rect 1803 -221 1815 -187
rect 1849 -221 1861 -187
rect 1803 -255 1861 -221
rect 1803 -289 1815 -255
rect 1849 -289 1861 -255
rect 1803 -323 1861 -289
rect 1803 -357 1815 -323
rect 1849 -357 1861 -323
rect 1803 -391 1861 -357
rect 1803 -425 1815 -391
rect 1849 -425 1861 -391
rect 1803 -459 1861 -425
rect 1803 -493 1815 -459
rect 1849 -493 1861 -459
rect 1803 -527 1861 -493
rect 1803 -561 1815 -527
rect 1849 -561 1861 -527
rect 1803 -595 1861 -561
rect 1803 -629 1815 -595
rect 1849 -629 1861 -595
rect 1803 -663 1861 -629
rect 1803 -697 1815 -663
rect 1849 -697 1861 -663
rect 1803 -731 1861 -697
rect 1803 -765 1815 -731
rect 1849 -765 1861 -731
rect 1803 -800 1861 -765
rect 2261 765 2319 800
rect 2261 731 2273 765
rect 2307 731 2319 765
rect 2261 697 2319 731
rect 2261 663 2273 697
rect 2307 663 2319 697
rect 2261 629 2319 663
rect 2261 595 2273 629
rect 2307 595 2319 629
rect 2261 561 2319 595
rect 2261 527 2273 561
rect 2307 527 2319 561
rect 2261 493 2319 527
rect 2261 459 2273 493
rect 2307 459 2319 493
rect 2261 425 2319 459
rect 2261 391 2273 425
rect 2307 391 2319 425
rect 2261 357 2319 391
rect 2261 323 2273 357
rect 2307 323 2319 357
rect 2261 289 2319 323
rect 2261 255 2273 289
rect 2307 255 2319 289
rect 2261 221 2319 255
rect 2261 187 2273 221
rect 2307 187 2319 221
rect 2261 153 2319 187
rect 2261 119 2273 153
rect 2307 119 2319 153
rect 2261 85 2319 119
rect 2261 51 2273 85
rect 2307 51 2319 85
rect 2261 17 2319 51
rect 2261 -17 2273 17
rect 2307 -17 2319 17
rect 2261 -51 2319 -17
rect 2261 -85 2273 -51
rect 2307 -85 2319 -51
rect 2261 -119 2319 -85
rect 2261 -153 2273 -119
rect 2307 -153 2319 -119
rect 2261 -187 2319 -153
rect 2261 -221 2273 -187
rect 2307 -221 2319 -187
rect 2261 -255 2319 -221
rect 2261 -289 2273 -255
rect 2307 -289 2319 -255
rect 2261 -323 2319 -289
rect 2261 -357 2273 -323
rect 2307 -357 2319 -323
rect 2261 -391 2319 -357
rect 2261 -425 2273 -391
rect 2307 -425 2319 -391
rect 2261 -459 2319 -425
rect 2261 -493 2273 -459
rect 2307 -493 2319 -459
rect 2261 -527 2319 -493
rect 2261 -561 2273 -527
rect 2307 -561 2319 -527
rect 2261 -595 2319 -561
rect 2261 -629 2273 -595
rect 2307 -629 2319 -595
rect 2261 -663 2319 -629
rect 2261 -697 2273 -663
rect 2307 -697 2319 -663
rect 2261 -731 2319 -697
rect 2261 -765 2273 -731
rect 2307 -765 2319 -731
rect 2261 -800 2319 -765
rect 2719 765 2777 800
rect 2719 731 2731 765
rect 2765 731 2777 765
rect 2719 697 2777 731
rect 2719 663 2731 697
rect 2765 663 2777 697
rect 2719 629 2777 663
rect 2719 595 2731 629
rect 2765 595 2777 629
rect 2719 561 2777 595
rect 2719 527 2731 561
rect 2765 527 2777 561
rect 2719 493 2777 527
rect 2719 459 2731 493
rect 2765 459 2777 493
rect 2719 425 2777 459
rect 2719 391 2731 425
rect 2765 391 2777 425
rect 2719 357 2777 391
rect 2719 323 2731 357
rect 2765 323 2777 357
rect 2719 289 2777 323
rect 2719 255 2731 289
rect 2765 255 2777 289
rect 2719 221 2777 255
rect 2719 187 2731 221
rect 2765 187 2777 221
rect 2719 153 2777 187
rect 2719 119 2731 153
rect 2765 119 2777 153
rect 2719 85 2777 119
rect 2719 51 2731 85
rect 2765 51 2777 85
rect 2719 17 2777 51
rect 2719 -17 2731 17
rect 2765 -17 2777 17
rect 2719 -51 2777 -17
rect 2719 -85 2731 -51
rect 2765 -85 2777 -51
rect 2719 -119 2777 -85
rect 2719 -153 2731 -119
rect 2765 -153 2777 -119
rect 2719 -187 2777 -153
rect 2719 -221 2731 -187
rect 2765 -221 2777 -187
rect 2719 -255 2777 -221
rect 2719 -289 2731 -255
rect 2765 -289 2777 -255
rect 2719 -323 2777 -289
rect 2719 -357 2731 -323
rect 2765 -357 2777 -323
rect 2719 -391 2777 -357
rect 2719 -425 2731 -391
rect 2765 -425 2777 -391
rect 2719 -459 2777 -425
rect 2719 -493 2731 -459
rect 2765 -493 2777 -459
rect 2719 -527 2777 -493
rect 2719 -561 2731 -527
rect 2765 -561 2777 -527
rect 2719 -595 2777 -561
rect 2719 -629 2731 -595
rect 2765 -629 2777 -595
rect 2719 -663 2777 -629
rect 2719 -697 2731 -663
rect 2765 -697 2777 -663
rect 2719 -731 2777 -697
rect 2719 -765 2731 -731
rect 2765 -765 2777 -731
rect 2719 -800 2777 -765
rect 3177 765 3235 800
rect 3177 731 3189 765
rect 3223 731 3235 765
rect 3177 697 3235 731
rect 3177 663 3189 697
rect 3223 663 3235 697
rect 3177 629 3235 663
rect 3177 595 3189 629
rect 3223 595 3235 629
rect 3177 561 3235 595
rect 3177 527 3189 561
rect 3223 527 3235 561
rect 3177 493 3235 527
rect 3177 459 3189 493
rect 3223 459 3235 493
rect 3177 425 3235 459
rect 3177 391 3189 425
rect 3223 391 3235 425
rect 3177 357 3235 391
rect 3177 323 3189 357
rect 3223 323 3235 357
rect 3177 289 3235 323
rect 3177 255 3189 289
rect 3223 255 3235 289
rect 3177 221 3235 255
rect 3177 187 3189 221
rect 3223 187 3235 221
rect 3177 153 3235 187
rect 3177 119 3189 153
rect 3223 119 3235 153
rect 3177 85 3235 119
rect 3177 51 3189 85
rect 3223 51 3235 85
rect 3177 17 3235 51
rect 3177 -17 3189 17
rect 3223 -17 3235 17
rect 3177 -51 3235 -17
rect 3177 -85 3189 -51
rect 3223 -85 3235 -51
rect 3177 -119 3235 -85
rect 3177 -153 3189 -119
rect 3223 -153 3235 -119
rect 3177 -187 3235 -153
rect 3177 -221 3189 -187
rect 3223 -221 3235 -187
rect 3177 -255 3235 -221
rect 3177 -289 3189 -255
rect 3223 -289 3235 -255
rect 3177 -323 3235 -289
rect 3177 -357 3189 -323
rect 3223 -357 3235 -323
rect 3177 -391 3235 -357
rect 3177 -425 3189 -391
rect 3223 -425 3235 -391
rect 3177 -459 3235 -425
rect 3177 -493 3189 -459
rect 3223 -493 3235 -459
rect 3177 -527 3235 -493
rect 3177 -561 3189 -527
rect 3223 -561 3235 -527
rect 3177 -595 3235 -561
rect 3177 -629 3189 -595
rect 3223 -629 3235 -595
rect 3177 -663 3235 -629
rect 3177 -697 3189 -663
rect 3223 -697 3235 -663
rect 3177 -731 3235 -697
rect 3177 -765 3189 -731
rect 3223 -765 3235 -731
rect 3177 -800 3235 -765
rect 3635 765 3693 800
rect 3635 731 3647 765
rect 3681 731 3693 765
rect 3635 697 3693 731
rect 3635 663 3647 697
rect 3681 663 3693 697
rect 3635 629 3693 663
rect 3635 595 3647 629
rect 3681 595 3693 629
rect 3635 561 3693 595
rect 3635 527 3647 561
rect 3681 527 3693 561
rect 3635 493 3693 527
rect 3635 459 3647 493
rect 3681 459 3693 493
rect 3635 425 3693 459
rect 3635 391 3647 425
rect 3681 391 3693 425
rect 3635 357 3693 391
rect 3635 323 3647 357
rect 3681 323 3693 357
rect 3635 289 3693 323
rect 3635 255 3647 289
rect 3681 255 3693 289
rect 3635 221 3693 255
rect 3635 187 3647 221
rect 3681 187 3693 221
rect 3635 153 3693 187
rect 3635 119 3647 153
rect 3681 119 3693 153
rect 3635 85 3693 119
rect 3635 51 3647 85
rect 3681 51 3693 85
rect 3635 17 3693 51
rect 3635 -17 3647 17
rect 3681 -17 3693 17
rect 3635 -51 3693 -17
rect 3635 -85 3647 -51
rect 3681 -85 3693 -51
rect 3635 -119 3693 -85
rect 3635 -153 3647 -119
rect 3681 -153 3693 -119
rect 3635 -187 3693 -153
rect 3635 -221 3647 -187
rect 3681 -221 3693 -187
rect 3635 -255 3693 -221
rect 3635 -289 3647 -255
rect 3681 -289 3693 -255
rect 3635 -323 3693 -289
rect 3635 -357 3647 -323
rect 3681 -357 3693 -323
rect 3635 -391 3693 -357
rect 3635 -425 3647 -391
rect 3681 -425 3693 -391
rect 3635 -459 3693 -425
rect 3635 -493 3647 -459
rect 3681 -493 3693 -459
rect 3635 -527 3693 -493
rect 3635 -561 3647 -527
rect 3681 -561 3693 -527
rect 3635 -595 3693 -561
rect 3635 -629 3647 -595
rect 3681 -629 3693 -595
rect 3635 -663 3693 -629
rect 3635 -697 3647 -663
rect 3681 -697 3693 -663
rect 3635 -731 3693 -697
rect 3635 -765 3647 -731
rect 3681 -765 3693 -731
rect 3635 -800 3693 -765
rect 4093 765 4151 800
rect 4093 731 4105 765
rect 4139 731 4151 765
rect 4093 697 4151 731
rect 4093 663 4105 697
rect 4139 663 4151 697
rect 4093 629 4151 663
rect 4093 595 4105 629
rect 4139 595 4151 629
rect 4093 561 4151 595
rect 4093 527 4105 561
rect 4139 527 4151 561
rect 4093 493 4151 527
rect 4093 459 4105 493
rect 4139 459 4151 493
rect 4093 425 4151 459
rect 4093 391 4105 425
rect 4139 391 4151 425
rect 4093 357 4151 391
rect 4093 323 4105 357
rect 4139 323 4151 357
rect 4093 289 4151 323
rect 4093 255 4105 289
rect 4139 255 4151 289
rect 4093 221 4151 255
rect 4093 187 4105 221
rect 4139 187 4151 221
rect 4093 153 4151 187
rect 4093 119 4105 153
rect 4139 119 4151 153
rect 4093 85 4151 119
rect 4093 51 4105 85
rect 4139 51 4151 85
rect 4093 17 4151 51
rect 4093 -17 4105 17
rect 4139 -17 4151 17
rect 4093 -51 4151 -17
rect 4093 -85 4105 -51
rect 4139 -85 4151 -51
rect 4093 -119 4151 -85
rect 4093 -153 4105 -119
rect 4139 -153 4151 -119
rect 4093 -187 4151 -153
rect 4093 -221 4105 -187
rect 4139 -221 4151 -187
rect 4093 -255 4151 -221
rect 4093 -289 4105 -255
rect 4139 -289 4151 -255
rect 4093 -323 4151 -289
rect 4093 -357 4105 -323
rect 4139 -357 4151 -323
rect 4093 -391 4151 -357
rect 4093 -425 4105 -391
rect 4139 -425 4151 -391
rect 4093 -459 4151 -425
rect 4093 -493 4105 -459
rect 4139 -493 4151 -459
rect 4093 -527 4151 -493
rect 4093 -561 4105 -527
rect 4139 -561 4151 -527
rect 4093 -595 4151 -561
rect 4093 -629 4105 -595
rect 4139 -629 4151 -595
rect 4093 -663 4151 -629
rect 4093 -697 4105 -663
rect 4139 -697 4151 -663
rect 4093 -731 4151 -697
rect 4093 -765 4105 -731
rect 4139 -765 4151 -731
rect 4093 -800 4151 -765
<< pdiffc >>
rect -4139 731 -4105 765
rect -4139 663 -4105 697
rect -4139 595 -4105 629
rect -4139 527 -4105 561
rect -4139 459 -4105 493
rect -4139 391 -4105 425
rect -4139 323 -4105 357
rect -4139 255 -4105 289
rect -4139 187 -4105 221
rect -4139 119 -4105 153
rect -4139 51 -4105 85
rect -4139 -17 -4105 17
rect -4139 -85 -4105 -51
rect -4139 -153 -4105 -119
rect -4139 -221 -4105 -187
rect -4139 -289 -4105 -255
rect -4139 -357 -4105 -323
rect -4139 -425 -4105 -391
rect -4139 -493 -4105 -459
rect -4139 -561 -4105 -527
rect -4139 -629 -4105 -595
rect -4139 -697 -4105 -663
rect -4139 -765 -4105 -731
rect -3681 731 -3647 765
rect -3681 663 -3647 697
rect -3681 595 -3647 629
rect -3681 527 -3647 561
rect -3681 459 -3647 493
rect -3681 391 -3647 425
rect -3681 323 -3647 357
rect -3681 255 -3647 289
rect -3681 187 -3647 221
rect -3681 119 -3647 153
rect -3681 51 -3647 85
rect -3681 -17 -3647 17
rect -3681 -85 -3647 -51
rect -3681 -153 -3647 -119
rect -3681 -221 -3647 -187
rect -3681 -289 -3647 -255
rect -3681 -357 -3647 -323
rect -3681 -425 -3647 -391
rect -3681 -493 -3647 -459
rect -3681 -561 -3647 -527
rect -3681 -629 -3647 -595
rect -3681 -697 -3647 -663
rect -3681 -765 -3647 -731
rect -3223 731 -3189 765
rect -3223 663 -3189 697
rect -3223 595 -3189 629
rect -3223 527 -3189 561
rect -3223 459 -3189 493
rect -3223 391 -3189 425
rect -3223 323 -3189 357
rect -3223 255 -3189 289
rect -3223 187 -3189 221
rect -3223 119 -3189 153
rect -3223 51 -3189 85
rect -3223 -17 -3189 17
rect -3223 -85 -3189 -51
rect -3223 -153 -3189 -119
rect -3223 -221 -3189 -187
rect -3223 -289 -3189 -255
rect -3223 -357 -3189 -323
rect -3223 -425 -3189 -391
rect -3223 -493 -3189 -459
rect -3223 -561 -3189 -527
rect -3223 -629 -3189 -595
rect -3223 -697 -3189 -663
rect -3223 -765 -3189 -731
rect -2765 731 -2731 765
rect -2765 663 -2731 697
rect -2765 595 -2731 629
rect -2765 527 -2731 561
rect -2765 459 -2731 493
rect -2765 391 -2731 425
rect -2765 323 -2731 357
rect -2765 255 -2731 289
rect -2765 187 -2731 221
rect -2765 119 -2731 153
rect -2765 51 -2731 85
rect -2765 -17 -2731 17
rect -2765 -85 -2731 -51
rect -2765 -153 -2731 -119
rect -2765 -221 -2731 -187
rect -2765 -289 -2731 -255
rect -2765 -357 -2731 -323
rect -2765 -425 -2731 -391
rect -2765 -493 -2731 -459
rect -2765 -561 -2731 -527
rect -2765 -629 -2731 -595
rect -2765 -697 -2731 -663
rect -2765 -765 -2731 -731
rect -2307 731 -2273 765
rect -2307 663 -2273 697
rect -2307 595 -2273 629
rect -2307 527 -2273 561
rect -2307 459 -2273 493
rect -2307 391 -2273 425
rect -2307 323 -2273 357
rect -2307 255 -2273 289
rect -2307 187 -2273 221
rect -2307 119 -2273 153
rect -2307 51 -2273 85
rect -2307 -17 -2273 17
rect -2307 -85 -2273 -51
rect -2307 -153 -2273 -119
rect -2307 -221 -2273 -187
rect -2307 -289 -2273 -255
rect -2307 -357 -2273 -323
rect -2307 -425 -2273 -391
rect -2307 -493 -2273 -459
rect -2307 -561 -2273 -527
rect -2307 -629 -2273 -595
rect -2307 -697 -2273 -663
rect -2307 -765 -2273 -731
rect -1849 731 -1815 765
rect -1849 663 -1815 697
rect -1849 595 -1815 629
rect -1849 527 -1815 561
rect -1849 459 -1815 493
rect -1849 391 -1815 425
rect -1849 323 -1815 357
rect -1849 255 -1815 289
rect -1849 187 -1815 221
rect -1849 119 -1815 153
rect -1849 51 -1815 85
rect -1849 -17 -1815 17
rect -1849 -85 -1815 -51
rect -1849 -153 -1815 -119
rect -1849 -221 -1815 -187
rect -1849 -289 -1815 -255
rect -1849 -357 -1815 -323
rect -1849 -425 -1815 -391
rect -1849 -493 -1815 -459
rect -1849 -561 -1815 -527
rect -1849 -629 -1815 -595
rect -1849 -697 -1815 -663
rect -1849 -765 -1815 -731
rect -1391 731 -1357 765
rect -1391 663 -1357 697
rect -1391 595 -1357 629
rect -1391 527 -1357 561
rect -1391 459 -1357 493
rect -1391 391 -1357 425
rect -1391 323 -1357 357
rect -1391 255 -1357 289
rect -1391 187 -1357 221
rect -1391 119 -1357 153
rect -1391 51 -1357 85
rect -1391 -17 -1357 17
rect -1391 -85 -1357 -51
rect -1391 -153 -1357 -119
rect -1391 -221 -1357 -187
rect -1391 -289 -1357 -255
rect -1391 -357 -1357 -323
rect -1391 -425 -1357 -391
rect -1391 -493 -1357 -459
rect -1391 -561 -1357 -527
rect -1391 -629 -1357 -595
rect -1391 -697 -1357 -663
rect -1391 -765 -1357 -731
rect -933 731 -899 765
rect -933 663 -899 697
rect -933 595 -899 629
rect -933 527 -899 561
rect -933 459 -899 493
rect -933 391 -899 425
rect -933 323 -899 357
rect -933 255 -899 289
rect -933 187 -899 221
rect -933 119 -899 153
rect -933 51 -899 85
rect -933 -17 -899 17
rect -933 -85 -899 -51
rect -933 -153 -899 -119
rect -933 -221 -899 -187
rect -933 -289 -899 -255
rect -933 -357 -899 -323
rect -933 -425 -899 -391
rect -933 -493 -899 -459
rect -933 -561 -899 -527
rect -933 -629 -899 -595
rect -933 -697 -899 -663
rect -933 -765 -899 -731
rect -475 731 -441 765
rect -475 663 -441 697
rect -475 595 -441 629
rect -475 527 -441 561
rect -475 459 -441 493
rect -475 391 -441 425
rect -475 323 -441 357
rect -475 255 -441 289
rect -475 187 -441 221
rect -475 119 -441 153
rect -475 51 -441 85
rect -475 -17 -441 17
rect -475 -85 -441 -51
rect -475 -153 -441 -119
rect -475 -221 -441 -187
rect -475 -289 -441 -255
rect -475 -357 -441 -323
rect -475 -425 -441 -391
rect -475 -493 -441 -459
rect -475 -561 -441 -527
rect -475 -629 -441 -595
rect -475 -697 -441 -663
rect -475 -765 -441 -731
rect -17 731 17 765
rect -17 663 17 697
rect -17 595 17 629
rect -17 527 17 561
rect -17 459 17 493
rect -17 391 17 425
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect -17 -425 17 -391
rect -17 -493 17 -459
rect -17 -561 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -663
rect -17 -765 17 -731
rect 441 731 475 765
rect 441 663 475 697
rect 441 595 475 629
rect 441 527 475 561
rect 441 459 475 493
rect 441 391 475 425
rect 441 323 475 357
rect 441 255 475 289
rect 441 187 475 221
rect 441 119 475 153
rect 441 51 475 85
rect 441 -17 475 17
rect 441 -85 475 -51
rect 441 -153 475 -119
rect 441 -221 475 -187
rect 441 -289 475 -255
rect 441 -357 475 -323
rect 441 -425 475 -391
rect 441 -493 475 -459
rect 441 -561 475 -527
rect 441 -629 475 -595
rect 441 -697 475 -663
rect 441 -765 475 -731
rect 899 731 933 765
rect 899 663 933 697
rect 899 595 933 629
rect 899 527 933 561
rect 899 459 933 493
rect 899 391 933 425
rect 899 323 933 357
rect 899 255 933 289
rect 899 187 933 221
rect 899 119 933 153
rect 899 51 933 85
rect 899 -17 933 17
rect 899 -85 933 -51
rect 899 -153 933 -119
rect 899 -221 933 -187
rect 899 -289 933 -255
rect 899 -357 933 -323
rect 899 -425 933 -391
rect 899 -493 933 -459
rect 899 -561 933 -527
rect 899 -629 933 -595
rect 899 -697 933 -663
rect 899 -765 933 -731
rect 1357 731 1391 765
rect 1357 663 1391 697
rect 1357 595 1391 629
rect 1357 527 1391 561
rect 1357 459 1391 493
rect 1357 391 1391 425
rect 1357 323 1391 357
rect 1357 255 1391 289
rect 1357 187 1391 221
rect 1357 119 1391 153
rect 1357 51 1391 85
rect 1357 -17 1391 17
rect 1357 -85 1391 -51
rect 1357 -153 1391 -119
rect 1357 -221 1391 -187
rect 1357 -289 1391 -255
rect 1357 -357 1391 -323
rect 1357 -425 1391 -391
rect 1357 -493 1391 -459
rect 1357 -561 1391 -527
rect 1357 -629 1391 -595
rect 1357 -697 1391 -663
rect 1357 -765 1391 -731
rect 1815 731 1849 765
rect 1815 663 1849 697
rect 1815 595 1849 629
rect 1815 527 1849 561
rect 1815 459 1849 493
rect 1815 391 1849 425
rect 1815 323 1849 357
rect 1815 255 1849 289
rect 1815 187 1849 221
rect 1815 119 1849 153
rect 1815 51 1849 85
rect 1815 -17 1849 17
rect 1815 -85 1849 -51
rect 1815 -153 1849 -119
rect 1815 -221 1849 -187
rect 1815 -289 1849 -255
rect 1815 -357 1849 -323
rect 1815 -425 1849 -391
rect 1815 -493 1849 -459
rect 1815 -561 1849 -527
rect 1815 -629 1849 -595
rect 1815 -697 1849 -663
rect 1815 -765 1849 -731
rect 2273 731 2307 765
rect 2273 663 2307 697
rect 2273 595 2307 629
rect 2273 527 2307 561
rect 2273 459 2307 493
rect 2273 391 2307 425
rect 2273 323 2307 357
rect 2273 255 2307 289
rect 2273 187 2307 221
rect 2273 119 2307 153
rect 2273 51 2307 85
rect 2273 -17 2307 17
rect 2273 -85 2307 -51
rect 2273 -153 2307 -119
rect 2273 -221 2307 -187
rect 2273 -289 2307 -255
rect 2273 -357 2307 -323
rect 2273 -425 2307 -391
rect 2273 -493 2307 -459
rect 2273 -561 2307 -527
rect 2273 -629 2307 -595
rect 2273 -697 2307 -663
rect 2273 -765 2307 -731
rect 2731 731 2765 765
rect 2731 663 2765 697
rect 2731 595 2765 629
rect 2731 527 2765 561
rect 2731 459 2765 493
rect 2731 391 2765 425
rect 2731 323 2765 357
rect 2731 255 2765 289
rect 2731 187 2765 221
rect 2731 119 2765 153
rect 2731 51 2765 85
rect 2731 -17 2765 17
rect 2731 -85 2765 -51
rect 2731 -153 2765 -119
rect 2731 -221 2765 -187
rect 2731 -289 2765 -255
rect 2731 -357 2765 -323
rect 2731 -425 2765 -391
rect 2731 -493 2765 -459
rect 2731 -561 2765 -527
rect 2731 -629 2765 -595
rect 2731 -697 2765 -663
rect 2731 -765 2765 -731
rect 3189 731 3223 765
rect 3189 663 3223 697
rect 3189 595 3223 629
rect 3189 527 3223 561
rect 3189 459 3223 493
rect 3189 391 3223 425
rect 3189 323 3223 357
rect 3189 255 3223 289
rect 3189 187 3223 221
rect 3189 119 3223 153
rect 3189 51 3223 85
rect 3189 -17 3223 17
rect 3189 -85 3223 -51
rect 3189 -153 3223 -119
rect 3189 -221 3223 -187
rect 3189 -289 3223 -255
rect 3189 -357 3223 -323
rect 3189 -425 3223 -391
rect 3189 -493 3223 -459
rect 3189 -561 3223 -527
rect 3189 -629 3223 -595
rect 3189 -697 3223 -663
rect 3189 -765 3223 -731
rect 3647 731 3681 765
rect 3647 663 3681 697
rect 3647 595 3681 629
rect 3647 527 3681 561
rect 3647 459 3681 493
rect 3647 391 3681 425
rect 3647 323 3681 357
rect 3647 255 3681 289
rect 3647 187 3681 221
rect 3647 119 3681 153
rect 3647 51 3681 85
rect 3647 -17 3681 17
rect 3647 -85 3681 -51
rect 3647 -153 3681 -119
rect 3647 -221 3681 -187
rect 3647 -289 3681 -255
rect 3647 -357 3681 -323
rect 3647 -425 3681 -391
rect 3647 -493 3681 -459
rect 3647 -561 3681 -527
rect 3647 -629 3681 -595
rect 3647 -697 3681 -663
rect 3647 -765 3681 -731
rect 4105 731 4139 765
rect 4105 663 4139 697
rect 4105 595 4139 629
rect 4105 527 4139 561
rect 4105 459 4139 493
rect 4105 391 4139 425
rect 4105 323 4139 357
rect 4105 255 4139 289
rect 4105 187 4139 221
rect 4105 119 4139 153
rect 4105 51 4139 85
rect 4105 -17 4139 17
rect 4105 -85 4139 -51
rect 4105 -153 4139 -119
rect 4105 -221 4139 -187
rect 4105 -289 4139 -255
rect 4105 -357 4139 -323
rect 4105 -425 4139 -391
rect 4105 -493 4139 -459
rect 4105 -561 4139 -527
rect 4105 -629 4139 -595
rect 4105 -697 4139 -663
rect 4105 -765 4139 -731
<< poly >>
rect -4019 881 -3767 897
rect -4019 864 -3978 881
rect -4093 847 -3978 864
rect -3944 847 -3910 881
rect -3876 847 -3842 881
rect -3808 864 -3767 881
rect -3561 881 -3309 897
rect -3561 864 -3520 881
rect -3808 847 -3693 864
rect -4093 800 -3693 847
rect -3635 847 -3520 864
rect -3486 847 -3452 881
rect -3418 847 -3384 881
rect -3350 864 -3309 881
rect -3103 881 -2851 897
rect -3103 864 -3062 881
rect -3350 847 -3235 864
rect -3635 800 -3235 847
rect -3177 847 -3062 864
rect -3028 847 -2994 881
rect -2960 847 -2926 881
rect -2892 864 -2851 881
rect -2645 881 -2393 897
rect -2645 864 -2604 881
rect -2892 847 -2777 864
rect -3177 800 -2777 847
rect -2719 847 -2604 864
rect -2570 847 -2536 881
rect -2502 847 -2468 881
rect -2434 864 -2393 881
rect -2187 881 -1935 897
rect -2187 864 -2146 881
rect -2434 847 -2319 864
rect -2719 800 -2319 847
rect -2261 847 -2146 864
rect -2112 847 -2078 881
rect -2044 847 -2010 881
rect -1976 864 -1935 881
rect -1729 881 -1477 897
rect -1729 864 -1688 881
rect -1976 847 -1861 864
rect -2261 800 -1861 847
rect -1803 847 -1688 864
rect -1654 847 -1620 881
rect -1586 847 -1552 881
rect -1518 864 -1477 881
rect -1271 881 -1019 897
rect -1271 864 -1230 881
rect -1518 847 -1403 864
rect -1803 800 -1403 847
rect -1345 847 -1230 864
rect -1196 847 -1162 881
rect -1128 847 -1094 881
rect -1060 864 -1019 881
rect -813 881 -561 897
rect -813 864 -772 881
rect -1060 847 -945 864
rect -1345 800 -945 847
rect -887 847 -772 864
rect -738 847 -704 881
rect -670 847 -636 881
rect -602 864 -561 881
rect -355 881 -103 897
rect -355 864 -314 881
rect -602 847 -487 864
rect -887 800 -487 847
rect -429 847 -314 864
rect -280 847 -246 881
rect -212 847 -178 881
rect -144 864 -103 881
rect 103 881 355 897
rect 103 864 144 881
rect -144 847 -29 864
rect -429 800 -29 847
rect 29 847 144 864
rect 178 847 212 881
rect 246 847 280 881
rect 314 864 355 881
rect 561 881 813 897
rect 561 864 602 881
rect 314 847 429 864
rect 29 800 429 847
rect 487 847 602 864
rect 636 847 670 881
rect 704 847 738 881
rect 772 864 813 881
rect 1019 881 1271 897
rect 1019 864 1060 881
rect 772 847 887 864
rect 487 800 887 847
rect 945 847 1060 864
rect 1094 847 1128 881
rect 1162 847 1196 881
rect 1230 864 1271 881
rect 1477 881 1729 897
rect 1477 864 1518 881
rect 1230 847 1345 864
rect 945 800 1345 847
rect 1403 847 1518 864
rect 1552 847 1586 881
rect 1620 847 1654 881
rect 1688 864 1729 881
rect 1935 881 2187 897
rect 1935 864 1976 881
rect 1688 847 1803 864
rect 1403 800 1803 847
rect 1861 847 1976 864
rect 2010 847 2044 881
rect 2078 847 2112 881
rect 2146 864 2187 881
rect 2393 881 2645 897
rect 2393 864 2434 881
rect 2146 847 2261 864
rect 1861 800 2261 847
rect 2319 847 2434 864
rect 2468 847 2502 881
rect 2536 847 2570 881
rect 2604 864 2645 881
rect 2851 881 3103 897
rect 2851 864 2892 881
rect 2604 847 2719 864
rect 2319 800 2719 847
rect 2777 847 2892 864
rect 2926 847 2960 881
rect 2994 847 3028 881
rect 3062 864 3103 881
rect 3309 881 3561 897
rect 3309 864 3350 881
rect 3062 847 3177 864
rect 2777 800 3177 847
rect 3235 847 3350 864
rect 3384 847 3418 881
rect 3452 847 3486 881
rect 3520 864 3561 881
rect 3767 881 4019 897
rect 3767 864 3808 881
rect 3520 847 3635 864
rect 3235 800 3635 847
rect 3693 847 3808 864
rect 3842 847 3876 881
rect 3910 847 3944 881
rect 3978 864 4019 881
rect 3978 847 4093 864
rect 3693 800 4093 847
rect -4093 -847 -3693 -800
rect -4093 -864 -3978 -847
rect -4019 -881 -3978 -864
rect -3944 -881 -3910 -847
rect -3876 -881 -3842 -847
rect -3808 -864 -3693 -847
rect -3635 -847 -3235 -800
rect -3635 -864 -3520 -847
rect -3808 -881 -3767 -864
rect -4019 -897 -3767 -881
rect -3561 -881 -3520 -864
rect -3486 -881 -3452 -847
rect -3418 -881 -3384 -847
rect -3350 -864 -3235 -847
rect -3177 -847 -2777 -800
rect -3177 -864 -3062 -847
rect -3350 -881 -3309 -864
rect -3561 -897 -3309 -881
rect -3103 -881 -3062 -864
rect -3028 -881 -2994 -847
rect -2960 -881 -2926 -847
rect -2892 -864 -2777 -847
rect -2719 -847 -2319 -800
rect -2719 -864 -2604 -847
rect -2892 -881 -2851 -864
rect -3103 -897 -2851 -881
rect -2645 -881 -2604 -864
rect -2570 -881 -2536 -847
rect -2502 -881 -2468 -847
rect -2434 -864 -2319 -847
rect -2261 -847 -1861 -800
rect -2261 -864 -2146 -847
rect -2434 -881 -2393 -864
rect -2645 -897 -2393 -881
rect -2187 -881 -2146 -864
rect -2112 -881 -2078 -847
rect -2044 -881 -2010 -847
rect -1976 -864 -1861 -847
rect -1803 -847 -1403 -800
rect -1803 -864 -1688 -847
rect -1976 -881 -1935 -864
rect -2187 -897 -1935 -881
rect -1729 -881 -1688 -864
rect -1654 -881 -1620 -847
rect -1586 -881 -1552 -847
rect -1518 -864 -1403 -847
rect -1345 -847 -945 -800
rect -1345 -864 -1230 -847
rect -1518 -881 -1477 -864
rect -1729 -897 -1477 -881
rect -1271 -881 -1230 -864
rect -1196 -881 -1162 -847
rect -1128 -881 -1094 -847
rect -1060 -864 -945 -847
rect -887 -847 -487 -800
rect -887 -864 -772 -847
rect -1060 -881 -1019 -864
rect -1271 -897 -1019 -881
rect -813 -881 -772 -864
rect -738 -881 -704 -847
rect -670 -881 -636 -847
rect -602 -864 -487 -847
rect -429 -847 -29 -800
rect -429 -864 -314 -847
rect -602 -881 -561 -864
rect -813 -897 -561 -881
rect -355 -881 -314 -864
rect -280 -881 -246 -847
rect -212 -881 -178 -847
rect -144 -864 -29 -847
rect 29 -847 429 -800
rect 29 -864 144 -847
rect -144 -881 -103 -864
rect -355 -897 -103 -881
rect 103 -881 144 -864
rect 178 -881 212 -847
rect 246 -881 280 -847
rect 314 -864 429 -847
rect 487 -847 887 -800
rect 487 -864 602 -847
rect 314 -881 355 -864
rect 103 -897 355 -881
rect 561 -881 602 -864
rect 636 -881 670 -847
rect 704 -881 738 -847
rect 772 -864 887 -847
rect 945 -847 1345 -800
rect 945 -864 1060 -847
rect 772 -881 813 -864
rect 561 -897 813 -881
rect 1019 -881 1060 -864
rect 1094 -881 1128 -847
rect 1162 -881 1196 -847
rect 1230 -864 1345 -847
rect 1403 -847 1803 -800
rect 1403 -864 1518 -847
rect 1230 -881 1271 -864
rect 1019 -897 1271 -881
rect 1477 -881 1518 -864
rect 1552 -881 1586 -847
rect 1620 -881 1654 -847
rect 1688 -864 1803 -847
rect 1861 -847 2261 -800
rect 1861 -864 1976 -847
rect 1688 -881 1729 -864
rect 1477 -897 1729 -881
rect 1935 -881 1976 -864
rect 2010 -881 2044 -847
rect 2078 -881 2112 -847
rect 2146 -864 2261 -847
rect 2319 -847 2719 -800
rect 2319 -864 2434 -847
rect 2146 -881 2187 -864
rect 1935 -897 2187 -881
rect 2393 -881 2434 -864
rect 2468 -881 2502 -847
rect 2536 -881 2570 -847
rect 2604 -864 2719 -847
rect 2777 -847 3177 -800
rect 2777 -864 2892 -847
rect 2604 -881 2645 -864
rect 2393 -897 2645 -881
rect 2851 -881 2892 -864
rect 2926 -881 2960 -847
rect 2994 -881 3028 -847
rect 3062 -864 3177 -847
rect 3235 -847 3635 -800
rect 3235 -864 3350 -847
rect 3062 -881 3103 -864
rect 2851 -897 3103 -881
rect 3309 -881 3350 -864
rect 3384 -881 3418 -847
rect 3452 -881 3486 -847
rect 3520 -864 3635 -847
rect 3693 -847 4093 -800
rect 3693 -864 3808 -847
rect 3520 -881 3561 -864
rect 3309 -897 3561 -881
rect 3767 -881 3808 -864
rect 3842 -881 3876 -847
rect 3910 -881 3944 -847
rect 3978 -864 4093 -847
rect 3978 -881 4019 -864
rect 3767 -897 4019 -881
<< polycont >>
rect -3978 847 -3944 881
rect -3910 847 -3876 881
rect -3842 847 -3808 881
rect -3520 847 -3486 881
rect -3452 847 -3418 881
rect -3384 847 -3350 881
rect -3062 847 -3028 881
rect -2994 847 -2960 881
rect -2926 847 -2892 881
rect -2604 847 -2570 881
rect -2536 847 -2502 881
rect -2468 847 -2434 881
rect -2146 847 -2112 881
rect -2078 847 -2044 881
rect -2010 847 -1976 881
rect -1688 847 -1654 881
rect -1620 847 -1586 881
rect -1552 847 -1518 881
rect -1230 847 -1196 881
rect -1162 847 -1128 881
rect -1094 847 -1060 881
rect -772 847 -738 881
rect -704 847 -670 881
rect -636 847 -602 881
rect -314 847 -280 881
rect -246 847 -212 881
rect -178 847 -144 881
rect 144 847 178 881
rect 212 847 246 881
rect 280 847 314 881
rect 602 847 636 881
rect 670 847 704 881
rect 738 847 772 881
rect 1060 847 1094 881
rect 1128 847 1162 881
rect 1196 847 1230 881
rect 1518 847 1552 881
rect 1586 847 1620 881
rect 1654 847 1688 881
rect 1976 847 2010 881
rect 2044 847 2078 881
rect 2112 847 2146 881
rect 2434 847 2468 881
rect 2502 847 2536 881
rect 2570 847 2604 881
rect 2892 847 2926 881
rect 2960 847 2994 881
rect 3028 847 3062 881
rect 3350 847 3384 881
rect 3418 847 3452 881
rect 3486 847 3520 881
rect 3808 847 3842 881
rect 3876 847 3910 881
rect 3944 847 3978 881
rect -3978 -881 -3944 -847
rect -3910 -881 -3876 -847
rect -3842 -881 -3808 -847
rect -3520 -881 -3486 -847
rect -3452 -881 -3418 -847
rect -3384 -881 -3350 -847
rect -3062 -881 -3028 -847
rect -2994 -881 -2960 -847
rect -2926 -881 -2892 -847
rect -2604 -881 -2570 -847
rect -2536 -881 -2502 -847
rect -2468 -881 -2434 -847
rect -2146 -881 -2112 -847
rect -2078 -881 -2044 -847
rect -2010 -881 -1976 -847
rect -1688 -881 -1654 -847
rect -1620 -881 -1586 -847
rect -1552 -881 -1518 -847
rect -1230 -881 -1196 -847
rect -1162 -881 -1128 -847
rect -1094 -881 -1060 -847
rect -772 -881 -738 -847
rect -704 -881 -670 -847
rect -636 -881 -602 -847
rect -314 -881 -280 -847
rect -246 -881 -212 -847
rect -178 -881 -144 -847
rect 144 -881 178 -847
rect 212 -881 246 -847
rect 280 -881 314 -847
rect 602 -881 636 -847
rect 670 -881 704 -847
rect 738 -881 772 -847
rect 1060 -881 1094 -847
rect 1128 -881 1162 -847
rect 1196 -881 1230 -847
rect 1518 -881 1552 -847
rect 1586 -881 1620 -847
rect 1654 -881 1688 -847
rect 1976 -881 2010 -847
rect 2044 -881 2078 -847
rect 2112 -881 2146 -847
rect 2434 -881 2468 -847
rect 2502 -881 2536 -847
rect 2570 -881 2604 -847
rect 2892 -881 2926 -847
rect 2960 -881 2994 -847
rect 3028 -881 3062 -847
rect 3350 -881 3384 -847
rect 3418 -881 3452 -847
rect 3486 -881 3520 -847
rect 3808 -881 3842 -847
rect 3876 -881 3910 -847
rect 3944 -881 3978 -847
<< locali >>
rect -4019 847 -3982 881
rect -3944 847 -3910 881
rect -3876 847 -3842 881
rect -3804 847 -3767 881
rect -3561 847 -3524 881
rect -3486 847 -3452 881
rect -3418 847 -3384 881
rect -3346 847 -3309 881
rect -3103 847 -3066 881
rect -3028 847 -2994 881
rect -2960 847 -2926 881
rect -2888 847 -2851 881
rect -2645 847 -2608 881
rect -2570 847 -2536 881
rect -2502 847 -2468 881
rect -2430 847 -2393 881
rect -2187 847 -2150 881
rect -2112 847 -2078 881
rect -2044 847 -2010 881
rect -1972 847 -1935 881
rect -1729 847 -1692 881
rect -1654 847 -1620 881
rect -1586 847 -1552 881
rect -1514 847 -1477 881
rect -1271 847 -1234 881
rect -1196 847 -1162 881
rect -1128 847 -1094 881
rect -1056 847 -1019 881
rect -813 847 -776 881
rect -738 847 -704 881
rect -670 847 -636 881
rect -598 847 -561 881
rect -355 847 -318 881
rect -280 847 -246 881
rect -212 847 -178 881
rect -140 847 -103 881
rect 103 847 140 881
rect 178 847 212 881
rect 246 847 280 881
rect 318 847 355 881
rect 561 847 598 881
rect 636 847 670 881
rect 704 847 738 881
rect 776 847 813 881
rect 1019 847 1056 881
rect 1094 847 1128 881
rect 1162 847 1196 881
rect 1234 847 1271 881
rect 1477 847 1514 881
rect 1552 847 1586 881
rect 1620 847 1654 881
rect 1692 847 1729 881
rect 1935 847 1972 881
rect 2010 847 2044 881
rect 2078 847 2112 881
rect 2150 847 2187 881
rect 2393 847 2430 881
rect 2468 847 2502 881
rect 2536 847 2570 881
rect 2608 847 2645 881
rect 2851 847 2888 881
rect 2926 847 2960 881
rect 2994 847 3028 881
rect 3066 847 3103 881
rect 3309 847 3346 881
rect 3384 847 3418 881
rect 3452 847 3486 881
rect 3524 847 3561 881
rect 3767 847 3804 881
rect 3842 847 3876 881
rect 3910 847 3944 881
rect 3982 847 4019 881
rect -4139 773 -4105 804
rect -4139 701 -4105 731
rect -4139 629 -4105 663
rect -4139 561 -4105 595
rect -4139 493 -4105 523
rect -4139 425 -4105 451
rect -4139 357 -4105 379
rect -4139 289 -4105 307
rect -4139 221 -4105 235
rect -4139 153 -4105 163
rect -4139 85 -4105 91
rect -4139 17 -4105 19
rect -4139 -19 -4105 -17
rect -4139 -91 -4105 -85
rect -4139 -163 -4105 -153
rect -4139 -235 -4105 -221
rect -4139 -307 -4105 -289
rect -4139 -379 -4105 -357
rect -4139 -451 -4105 -425
rect -4139 -523 -4105 -493
rect -4139 -595 -4105 -561
rect -4139 -663 -4105 -629
rect -4139 -731 -4105 -701
rect -4139 -804 -4105 -773
rect -3681 773 -3647 804
rect -3681 701 -3647 731
rect -3681 629 -3647 663
rect -3681 561 -3647 595
rect -3681 493 -3647 523
rect -3681 425 -3647 451
rect -3681 357 -3647 379
rect -3681 289 -3647 307
rect -3681 221 -3647 235
rect -3681 153 -3647 163
rect -3681 85 -3647 91
rect -3681 17 -3647 19
rect -3681 -19 -3647 -17
rect -3681 -91 -3647 -85
rect -3681 -163 -3647 -153
rect -3681 -235 -3647 -221
rect -3681 -307 -3647 -289
rect -3681 -379 -3647 -357
rect -3681 -451 -3647 -425
rect -3681 -523 -3647 -493
rect -3681 -595 -3647 -561
rect -3681 -663 -3647 -629
rect -3681 -731 -3647 -701
rect -3681 -804 -3647 -773
rect -3223 773 -3189 804
rect -3223 701 -3189 731
rect -3223 629 -3189 663
rect -3223 561 -3189 595
rect -3223 493 -3189 523
rect -3223 425 -3189 451
rect -3223 357 -3189 379
rect -3223 289 -3189 307
rect -3223 221 -3189 235
rect -3223 153 -3189 163
rect -3223 85 -3189 91
rect -3223 17 -3189 19
rect -3223 -19 -3189 -17
rect -3223 -91 -3189 -85
rect -3223 -163 -3189 -153
rect -3223 -235 -3189 -221
rect -3223 -307 -3189 -289
rect -3223 -379 -3189 -357
rect -3223 -451 -3189 -425
rect -3223 -523 -3189 -493
rect -3223 -595 -3189 -561
rect -3223 -663 -3189 -629
rect -3223 -731 -3189 -701
rect -3223 -804 -3189 -773
rect -2765 773 -2731 804
rect -2765 701 -2731 731
rect -2765 629 -2731 663
rect -2765 561 -2731 595
rect -2765 493 -2731 523
rect -2765 425 -2731 451
rect -2765 357 -2731 379
rect -2765 289 -2731 307
rect -2765 221 -2731 235
rect -2765 153 -2731 163
rect -2765 85 -2731 91
rect -2765 17 -2731 19
rect -2765 -19 -2731 -17
rect -2765 -91 -2731 -85
rect -2765 -163 -2731 -153
rect -2765 -235 -2731 -221
rect -2765 -307 -2731 -289
rect -2765 -379 -2731 -357
rect -2765 -451 -2731 -425
rect -2765 -523 -2731 -493
rect -2765 -595 -2731 -561
rect -2765 -663 -2731 -629
rect -2765 -731 -2731 -701
rect -2765 -804 -2731 -773
rect -2307 773 -2273 804
rect -2307 701 -2273 731
rect -2307 629 -2273 663
rect -2307 561 -2273 595
rect -2307 493 -2273 523
rect -2307 425 -2273 451
rect -2307 357 -2273 379
rect -2307 289 -2273 307
rect -2307 221 -2273 235
rect -2307 153 -2273 163
rect -2307 85 -2273 91
rect -2307 17 -2273 19
rect -2307 -19 -2273 -17
rect -2307 -91 -2273 -85
rect -2307 -163 -2273 -153
rect -2307 -235 -2273 -221
rect -2307 -307 -2273 -289
rect -2307 -379 -2273 -357
rect -2307 -451 -2273 -425
rect -2307 -523 -2273 -493
rect -2307 -595 -2273 -561
rect -2307 -663 -2273 -629
rect -2307 -731 -2273 -701
rect -2307 -804 -2273 -773
rect -1849 773 -1815 804
rect -1849 701 -1815 731
rect -1849 629 -1815 663
rect -1849 561 -1815 595
rect -1849 493 -1815 523
rect -1849 425 -1815 451
rect -1849 357 -1815 379
rect -1849 289 -1815 307
rect -1849 221 -1815 235
rect -1849 153 -1815 163
rect -1849 85 -1815 91
rect -1849 17 -1815 19
rect -1849 -19 -1815 -17
rect -1849 -91 -1815 -85
rect -1849 -163 -1815 -153
rect -1849 -235 -1815 -221
rect -1849 -307 -1815 -289
rect -1849 -379 -1815 -357
rect -1849 -451 -1815 -425
rect -1849 -523 -1815 -493
rect -1849 -595 -1815 -561
rect -1849 -663 -1815 -629
rect -1849 -731 -1815 -701
rect -1849 -804 -1815 -773
rect -1391 773 -1357 804
rect -1391 701 -1357 731
rect -1391 629 -1357 663
rect -1391 561 -1357 595
rect -1391 493 -1357 523
rect -1391 425 -1357 451
rect -1391 357 -1357 379
rect -1391 289 -1357 307
rect -1391 221 -1357 235
rect -1391 153 -1357 163
rect -1391 85 -1357 91
rect -1391 17 -1357 19
rect -1391 -19 -1357 -17
rect -1391 -91 -1357 -85
rect -1391 -163 -1357 -153
rect -1391 -235 -1357 -221
rect -1391 -307 -1357 -289
rect -1391 -379 -1357 -357
rect -1391 -451 -1357 -425
rect -1391 -523 -1357 -493
rect -1391 -595 -1357 -561
rect -1391 -663 -1357 -629
rect -1391 -731 -1357 -701
rect -1391 -804 -1357 -773
rect -933 773 -899 804
rect -933 701 -899 731
rect -933 629 -899 663
rect -933 561 -899 595
rect -933 493 -899 523
rect -933 425 -899 451
rect -933 357 -899 379
rect -933 289 -899 307
rect -933 221 -899 235
rect -933 153 -899 163
rect -933 85 -899 91
rect -933 17 -899 19
rect -933 -19 -899 -17
rect -933 -91 -899 -85
rect -933 -163 -899 -153
rect -933 -235 -899 -221
rect -933 -307 -899 -289
rect -933 -379 -899 -357
rect -933 -451 -899 -425
rect -933 -523 -899 -493
rect -933 -595 -899 -561
rect -933 -663 -899 -629
rect -933 -731 -899 -701
rect -933 -804 -899 -773
rect -475 773 -441 804
rect -475 701 -441 731
rect -475 629 -441 663
rect -475 561 -441 595
rect -475 493 -441 523
rect -475 425 -441 451
rect -475 357 -441 379
rect -475 289 -441 307
rect -475 221 -441 235
rect -475 153 -441 163
rect -475 85 -441 91
rect -475 17 -441 19
rect -475 -19 -441 -17
rect -475 -91 -441 -85
rect -475 -163 -441 -153
rect -475 -235 -441 -221
rect -475 -307 -441 -289
rect -475 -379 -441 -357
rect -475 -451 -441 -425
rect -475 -523 -441 -493
rect -475 -595 -441 -561
rect -475 -663 -441 -629
rect -475 -731 -441 -701
rect -475 -804 -441 -773
rect -17 773 17 804
rect -17 701 17 731
rect -17 629 17 663
rect -17 561 17 595
rect -17 493 17 523
rect -17 425 17 451
rect -17 357 17 379
rect -17 289 17 307
rect -17 221 17 235
rect -17 153 17 163
rect -17 85 17 91
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -91 17 -85
rect -17 -163 17 -153
rect -17 -235 17 -221
rect -17 -307 17 -289
rect -17 -379 17 -357
rect -17 -451 17 -425
rect -17 -523 17 -493
rect -17 -595 17 -561
rect -17 -663 17 -629
rect -17 -731 17 -701
rect -17 -804 17 -773
rect 441 773 475 804
rect 441 701 475 731
rect 441 629 475 663
rect 441 561 475 595
rect 441 493 475 523
rect 441 425 475 451
rect 441 357 475 379
rect 441 289 475 307
rect 441 221 475 235
rect 441 153 475 163
rect 441 85 475 91
rect 441 17 475 19
rect 441 -19 475 -17
rect 441 -91 475 -85
rect 441 -163 475 -153
rect 441 -235 475 -221
rect 441 -307 475 -289
rect 441 -379 475 -357
rect 441 -451 475 -425
rect 441 -523 475 -493
rect 441 -595 475 -561
rect 441 -663 475 -629
rect 441 -731 475 -701
rect 441 -804 475 -773
rect 899 773 933 804
rect 899 701 933 731
rect 899 629 933 663
rect 899 561 933 595
rect 899 493 933 523
rect 899 425 933 451
rect 899 357 933 379
rect 899 289 933 307
rect 899 221 933 235
rect 899 153 933 163
rect 899 85 933 91
rect 899 17 933 19
rect 899 -19 933 -17
rect 899 -91 933 -85
rect 899 -163 933 -153
rect 899 -235 933 -221
rect 899 -307 933 -289
rect 899 -379 933 -357
rect 899 -451 933 -425
rect 899 -523 933 -493
rect 899 -595 933 -561
rect 899 -663 933 -629
rect 899 -731 933 -701
rect 899 -804 933 -773
rect 1357 773 1391 804
rect 1357 701 1391 731
rect 1357 629 1391 663
rect 1357 561 1391 595
rect 1357 493 1391 523
rect 1357 425 1391 451
rect 1357 357 1391 379
rect 1357 289 1391 307
rect 1357 221 1391 235
rect 1357 153 1391 163
rect 1357 85 1391 91
rect 1357 17 1391 19
rect 1357 -19 1391 -17
rect 1357 -91 1391 -85
rect 1357 -163 1391 -153
rect 1357 -235 1391 -221
rect 1357 -307 1391 -289
rect 1357 -379 1391 -357
rect 1357 -451 1391 -425
rect 1357 -523 1391 -493
rect 1357 -595 1391 -561
rect 1357 -663 1391 -629
rect 1357 -731 1391 -701
rect 1357 -804 1391 -773
rect 1815 773 1849 804
rect 1815 701 1849 731
rect 1815 629 1849 663
rect 1815 561 1849 595
rect 1815 493 1849 523
rect 1815 425 1849 451
rect 1815 357 1849 379
rect 1815 289 1849 307
rect 1815 221 1849 235
rect 1815 153 1849 163
rect 1815 85 1849 91
rect 1815 17 1849 19
rect 1815 -19 1849 -17
rect 1815 -91 1849 -85
rect 1815 -163 1849 -153
rect 1815 -235 1849 -221
rect 1815 -307 1849 -289
rect 1815 -379 1849 -357
rect 1815 -451 1849 -425
rect 1815 -523 1849 -493
rect 1815 -595 1849 -561
rect 1815 -663 1849 -629
rect 1815 -731 1849 -701
rect 1815 -804 1849 -773
rect 2273 773 2307 804
rect 2273 701 2307 731
rect 2273 629 2307 663
rect 2273 561 2307 595
rect 2273 493 2307 523
rect 2273 425 2307 451
rect 2273 357 2307 379
rect 2273 289 2307 307
rect 2273 221 2307 235
rect 2273 153 2307 163
rect 2273 85 2307 91
rect 2273 17 2307 19
rect 2273 -19 2307 -17
rect 2273 -91 2307 -85
rect 2273 -163 2307 -153
rect 2273 -235 2307 -221
rect 2273 -307 2307 -289
rect 2273 -379 2307 -357
rect 2273 -451 2307 -425
rect 2273 -523 2307 -493
rect 2273 -595 2307 -561
rect 2273 -663 2307 -629
rect 2273 -731 2307 -701
rect 2273 -804 2307 -773
rect 2731 773 2765 804
rect 2731 701 2765 731
rect 2731 629 2765 663
rect 2731 561 2765 595
rect 2731 493 2765 523
rect 2731 425 2765 451
rect 2731 357 2765 379
rect 2731 289 2765 307
rect 2731 221 2765 235
rect 2731 153 2765 163
rect 2731 85 2765 91
rect 2731 17 2765 19
rect 2731 -19 2765 -17
rect 2731 -91 2765 -85
rect 2731 -163 2765 -153
rect 2731 -235 2765 -221
rect 2731 -307 2765 -289
rect 2731 -379 2765 -357
rect 2731 -451 2765 -425
rect 2731 -523 2765 -493
rect 2731 -595 2765 -561
rect 2731 -663 2765 -629
rect 2731 -731 2765 -701
rect 2731 -804 2765 -773
rect 3189 773 3223 804
rect 3189 701 3223 731
rect 3189 629 3223 663
rect 3189 561 3223 595
rect 3189 493 3223 523
rect 3189 425 3223 451
rect 3189 357 3223 379
rect 3189 289 3223 307
rect 3189 221 3223 235
rect 3189 153 3223 163
rect 3189 85 3223 91
rect 3189 17 3223 19
rect 3189 -19 3223 -17
rect 3189 -91 3223 -85
rect 3189 -163 3223 -153
rect 3189 -235 3223 -221
rect 3189 -307 3223 -289
rect 3189 -379 3223 -357
rect 3189 -451 3223 -425
rect 3189 -523 3223 -493
rect 3189 -595 3223 -561
rect 3189 -663 3223 -629
rect 3189 -731 3223 -701
rect 3189 -804 3223 -773
rect 3647 773 3681 804
rect 3647 701 3681 731
rect 3647 629 3681 663
rect 3647 561 3681 595
rect 3647 493 3681 523
rect 3647 425 3681 451
rect 3647 357 3681 379
rect 3647 289 3681 307
rect 3647 221 3681 235
rect 3647 153 3681 163
rect 3647 85 3681 91
rect 3647 17 3681 19
rect 3647 -19 3681 -17
rect 3647 -91 3681 -85
rect 3647 -163 3681 -153
rect 3647 -235 3681 -221
rect 3647 -307 3681 -289
rect 3647 -379 3681 -357
rect 3647 -451 3681 -425
rect 3647 -523 3681 -493
rect 3647 -595 3681 -561
rect 3647 -663 3681 -629
rect 3647 -731 3681 -701
rect 3647 -804 3681 -773
rect 4105 773 4139 804
rect 4105 701 4139 731
rect 4105 629 4139 663
rect 4105 561 4139 595
rect 4105 493 4139 523
rect 4105 425 4139 451
rect 4105 357 4139 379
rect 4105 289 4139 307
rect 4105 221 4139 235
rect 4105 153 4139 163
rect 4105 85 4139 91
rect 4105 17 4139 19
rect 4105 -19 4139 -17
rect 4105 -91 4139 -85
rect 4105 -163 4139 -153
rect 4105 -235 4139 -221
rect 4105 -307 4139 -289
rect 4105 -379 4139 -357
rect 4105 -451 4139 -425
rect 4105 -523 4139 -493
rect 4105 -595 4139 -561
rect 4105 -663 4139 -629
rect 4105 -731 4139 -701
rect 4105 -804 4139 -773
rect -4019 -881 -3982 -847
rect -3944 -881 -3910 -847
rect -3876 -881 -3842 -847
rect -3804 -881 -3767 -847
rect -3561 -881 -3524 -847
rect -3486 -881 -3452 -847
rect -3418 -881 -3384 -847
rect -3346 -881 -3309 -847
rect -3103 -881 -3066 -847
rect -3028 -881 -2994 -847
rect -2960 -881 -2926 -847
rect -2888 -881 -2851 -847
rect -2645 -881 -2608 -847
rect -2570 -881 -2536 -847
rect -2502 -881 -2468 -847
rect -2430 -881 -2393 -847
rect -2187 -881 -2150 -847
rect -2112 -881 -2078 -847
rect -2044 -881 -2010 -847
rect -1972 -881 -1935 -847
rect -1729 -881 -1692 -847
rect -1654 -881 -1620 -847
rect -1586 -881 -1552 -847
rect -1514 -881 -1477 -847
rect -1271 -881 -1234 -847
rect -1196 -881 -1162 -847
rect -1128 -881 -1094 -847
rect -1056 -881 -1019 -847
rect -813 -881 -776 -847
rect -738 -881 -704 -847
rect -670 -881 -636 -847
rect -598 -881 -561 -847
rect -355 -881 -318 -847
rect -280 -881 -246 -847
rect -212 -881 -178 -847
rect -140 -881 -103 -847
rect 103 -881 140 -847
rect 178 -881 212 -847
rect 246 -881 280 -847
rect 318 -881 355 -847
rect 561 -881 598 -847
rect 636 -881 670 -847
rect 704 -881 738 -847
rect 776 -881 813 -847
rect 1019 -881 1056 -847
rect 1094 -881 1128 -847
rect 1162 -881 1196 -847
rect 1234 -881 1271 -847
rect 1477 -881 1514 -847
rect 1552 -881 1586 -847
rect 1620 -881 1654 -847
rect 1692 -881 1729 -847
rect 1935 -881 1972 -847
rect 2010 -881 2044 -847
rect 2078 -881 2112 -847
rect 2150 -881 2187 -847
rect 2393 -881 2430 -847
rect 2468 -881 2502 -847
rect 2536 -881 2570 -847
rect 2608 -881 2645 -847
rect 2851 -881 2888 -847
rect 2926 -881 2960 -847
rect 2994 -881 3028 -847
rect 3066 -881 3103 -847
rect 3309 -881 3346 -847
rect 3384 -881 3418 -847
rect 3452 -881 3486 -847
rect 3524 -881 3561 -847
rect 3767 -881 3804 -847
rect 3842 -881 3876 -847
rect 3910 -881 3944 -847
rect 3982 -881 4019 -847
<< viali >>
rect -3982 847 -3978 881
rect -3978 847 -3948 881
rect -3910 847 -3876 881
rect -3838 847 -3808 881
rect -3808 847 -3804 881
rect -3524 847 -3520 881
rect -3520 847 -3490 881
rect -3452 847 -3418 881
rect -3380 847 -3350 881
rect -3350 847 -3346 881
rect -3066 847 -3062 881
rect -3062 847 -3032 881
rect -2994 847 -2960 881
rect -2922 847 -2892 881
rect -2892 847 -2888 881
rect -2608 847 -2604 881
rect -2604 847 -2574 881
rect -2536 847 -2502 881
rect -2464 847 -2434 881
rect -2434 847 -2430 881
rect -2150 847 -2146 881
rect -2146 847 -2116 881
rect -2078 847 -2044 881
rect -2006 847 -1976 881
rect -1976 847 -1972 881
rect -1692 847 -1688 881
rect -1688 847 -1658 881
rect -1620 847 -1586 881
rect -1548 847 -1518 881
rect -1518 847 -1514 881
rect -1234 847 -1230 881
rect -1230 847 -1200 881
rect -1162 847 -1128 881
rect -1090 847 -1060 881
rect -1060 847 -1056 881
rect -776 847 -772 881
rect -772 847 -742 881
rect -704 847 -670 881
rect -632 847 -602 881
rect -602 847 -598 881
rect -318 847 -314 881
rect -314 847 -284 881
rect -246 847 -212 881
rect -174 847 -144 881
rect -144 847 -140 881
rect 140 847 144 881
rect 144 847 174 881
rect 212 847 246 881
rect 284 847 314 881
rect 314 847 318 881
rect 598 847 602 881
rect 602 847 632 881
rect 670 847 704 881
rect 742 847 772 881
rect 772 847 776 881
rect 1056 847 1060 881
rect 1060 847 1090 881
rect 1128 847 1162 881
rect 1200 847 1230 881
rect 1230 847 1234 881
rect 1514 847 1518 881
rect 1518 847 1548 881
rect 1586 847 1620 881
rect 1658 847 1688 881
rect 1688 847 1692 881
rect 1972 847 1976 881
rect 1976 847 2006 881
rect 2044 847 2078 881
rect 2116 847 2146 881
rect 2146 847 2150 881
rect 2430 847 2434 881
rect 2434 847 2464 881
rect 2502 847 2536 881
rect 2574 847 2604 881
rect 2604 847 2608 881
rect 2888 847 2892 881
rect 2892 847 2922 881
rect 2960 847 2994 881
rect 3032 847 3062 881
rect 3062 847 3066 881
rect 3346 847 3350 881
rect 3350 847 3380 881
rect 3418 847 3452 881
rect 3490 847 3520 881
rect 3520 847 3524 881
rect 3804 847 3808 881
rect 3808 847 3838 881
rect 3876 847 3910 881
rect 3948 847 3978 881
rect 3978 847 3982 881
rect -4139 765 -4105 773
rect -4139 739 -4105 765
rect -4139 697 -4105 701
rect -4139 667 -4105 697
rect -4139 595 -4105 629
rect -4139 527 -4105 557
rect -4139 523 -4105 527
rect -4139 459 -4105 485
rect -4139 451 -4105 459
rect -4139 391 -4105 413
rect -4139 379 -4105 391
rect -4139 323 -4105 341
rect -4139 307 -4105 323
rect -4139 255 -4105 269
rect -4139 235 -4105 255
rect -4139 187 -4105 197
rect -4139 163 -4105 187
rect -4139 119 -4105 125
rect -4139 91 -4105 119
rect -4139 51 -4105 53
rect -4139 19 -4105 51
rect -4139 -51 -4105 -19
rect -4139 -53 -4105 -51
rect -4139 -119 -4105 -91
rect -4139 -125 -4105 -119
rect -4139 -187 -4105 -163
rect -4139 -197 -4105 -187
rect -4139 -255 -4105 -235
rect -4139 -269 -4105 -255
rect -4139 -323 -4105 -307
rect -4139 -341 -4105 -323
rect -4139 -391 -4105 -379
rect -4139 -413 -4105 -391
rect -4139 -459 -4105 -451
rect -4139 -485 -4105 -459
rect -4139 -527 -4105 -523
rect -4139 -557 -4105 -527
rect -4139 -629 -4105 -595
rect -4139 -697 -4105 -667
rect -4139 -701 -4105 -697
rect -4139 -765 -4105 -739
rect -4139 -773 -4105 -765
rect -3681 765 -3647 773
rect -3681 739 -3647 765
rect -3681 697 -3647 701
rect -3681 667 -3647 697
rect -3681 595 -3647 629
rect -3681 527 -3647 557
rect -3681 523 -3647 527
rect -3681 459 -3647 485
rect -3681 451 -3647 459
rect -3681 391 -3647 413
rect -3681 379 -3647 391
rect -3681 323 -3647 341
rect -3681 307 -3647 323
rect -3681 255 -3647 269
rect -3681 235 -3647 255
rect -3681 187 -3647 197
rect -3681 163 -3647 187
rect -3681 119 -3647 125
rect -3681 91 -3647 119
rect -3681 51 -3647 53
rect -3681 19 -3647 51
rect -3681 -51 -3647 -19
rect -3681 -53 -3647 -51
rect -3681 -119 -3647 -91
rect -3681 -125 -3647 -119
rect -3681 -187 -3647 -163
rect -3681 -197 -3647 -187
rect -3681 -255 -3647 -235
rect -3681 -269 -3647 -255
rect -3681 -323 -3647 -307
rect -3681 -341 -3647 -323
rect -3681 -391 -3647 -379
rect -3681 -413 -3647 -391
rect -3681 -459 -3647 -451
rect -3681 -485 -3647 -459
rect -3681 -527 -3647 -523
rect -3681 -557 -3647 -527
rect -3681 -629 -3647 -595
rect -3681 -697 -3647 -667
rect -3681 -701 -3647 -697
rect -3681 -765 -3647 -739
rect -3681 -773 -3647 -765
rect -3223 765 -3189 773
rect -3223 739 -3189 765
rect -3223 697 -3189 701
rect -3223 667 -3189 697
rect -3223 595 -3189 629
rect -3223 527 -3189 557
rect -3223 523 -3189 527
rect -3223 459 -3189 485
rect -3223 451 -3189 459
rect -3223 391 -3189 413
rect -3223 379 -3189 391
rect -3223 323 -3189 341
rect -3223 307 -3189 323
rect -3223 255 -3189 269
rect -3223 235 -3189 255
rect -3223 187 -3189 197
rect -3223 163 -3189 187
rect -3223 119 -3189 125
rect -3223 91 -3189 119
rect -3223 51 -3189 53
rect -3223 19 -3189 51
rect -3223 -51 -3189 -19
rect -3223 -53 -3189 -51
rect -3223 -119 -3189 -91
rect -3223 -125 -3189 -119
rect -3223 -187 -3189 -163
rect -3223 -197 -3189 -187
rect -3223 -255 -3189 -235
rect -3223 -269 -3189 -255
rect -3223 -323 -3189 -307
rect -3223 -341 -3189 -323
rect -3223 -391 -3189 -379
rect -3223 -413 -3189 -391
rect -3223 -459 -3189 -451
rect -3223 -485 -3189 -459
rect -3223 -527 -3189 -523
rect -3223 -557 -3189 -527
rect -3223 -629 -3189 -595
rect -3223 -697 -3189 -667
rect -3223 -701 -3189 -697
rect -3223 -765 -3189 -739
rect -3223 -773 -3189 -765
rect -2765 765 -2731 773
rect -2765 739 -2731 765
rect -2765 697 -2731 701
rect -2765 667 -2731 697
rect -2765 595 -2731 629
rect -2765 527 -2731 557
rect -2765 523 -2731 527
rect -2765 459 -2731 485
rect -2765 451 -2731 459
rect -2765 391 -2731 413
rect -2765 379 -2731 391
rect -2765 323 -2731 341
rect -2765 307 -2731 323
rect -2765 255 -2731 269
rect -2765 235 -2731 255
rect -2765 187 -2731 197
rect -2765 163 -2731 187
rect -2765 119 -2731 125
rect -2765 91 -2731 119
rect -2765 51 -2731 53
rect -2765 19 -2731 51
rect -2765 -51 -2731 -19
rect -2765 -53 -2731 -51
rect -2765 -119 -2731 -91
rect -2765 -125 -2731 -119
rect -2765 -187 -2731 -163
rect -2765 -197 -2731 -187
rect -2765 -255 -2731 -235
rect -2765 -269 -2731 -255
rect -2765 -323 -2731 -307
rect -2765 -341 -2731 -323
rect -2765 -391 -2731 -379
rect -2765 -413 -2731 -391
rect -2765 -459 -2731 -451
rect -2765 -485 -2731 -459
rect -2765 -527 -2731 -523
rect -2765 -557 -2731 -527
rect -2765 -629 -2731 -595
rect -2765 -697 -2731 -667
rect -2765 -701 -2731 -697
rect -2765 -765 -2731 -739
rect -2765 -773 -2731 -765
rect -2307 765 -2273 773
rect -2307 739 -2273 765
rect -2307 697 -2273 701
rect -2307 667 -2273 697
rect -2307 595 -2273 629
rect -2307 527 -2273 557
rect -2307 523 -2273 527
rect -2307 459 -2273 485
rect -2307 451 -2273 459
rect -2307 391 -2273 413
rect -2307 379 -2273 391
rect -2307 323 -2273 341
rect -2307 307 -2273 323
rect -2307 255 -2273 269
rect -2307 235 -2273 255
rect -2307 187 -2273 197
rect -2307 163 -2273 187
rect -2307 119 -2273 125
rect -2307 91 -2273 119
rect -2307 51 -2273 53
rect -2307 19 -2273 51
rect -2307 -51 -2273 -19
rect -2307 -53 -2273 -51
rect -2307 -119 -2273 -91
rect -2307 -125 -2273 -119
rect -2307 -187 -2273 -163
rect -2307 -197 -2273 -187
rect -2307 -255 -2273 -235
rect -2307 -269 -2273 -255
rect -2307 -323 -2273 -307
rect -2307 -341 -2273 -323
rect -2307 -391 -2273 -379
rect -2307 -413 -2273 -391
rect -2307 -459 -2273 -451
rect -2307 -485 -2273 -459
rect -2307 -527 -2273 -523
rect -2307 -557 -2273 -527
rect -2307 -629 -2273 -595
rect -2307 -697 -2273 -667
rect -2307 -701 -2273 -697
rect -2307 -765 -2273 -739
rect -2307 -773 -2273 -765
rect -1849 765 -1815 773
rect -1849 739 -1815 765
rect -1849 697 -1815 701
rect -1849 667 -1815 697
rect -1849 595 -1815 629
rect -1849 527 -1815 557
rect -1849 523 -1815 527
rect -1849 459 -1815 485
rect -1849 451 -1815 459
rect -1849 391 -1815 413
rect -1849 379 -1815 391
rect -1849 323 -1815 341
rect -1849 307 -1815 323
rect -1849 255 -1815 269
rect -1849 235 -1815 255
rect -1849 187 -1815 197
rect -1849 163 -1815 187
rect -1849 119 -1815 125
rect -1849 91 -1815 119
rect -1849 51 -1815 53
rect -1849 19 -1815 51
rect -1849 -51 -1815 -19
rect -1849 -53 -1815 -51
rect -1849 -119 -1815 -91
rect -1849 -125 -1815 -119
rect -1849 -187 -1815 -163
rect -1849 -197 -1815 -187
rect -1849 -255 -1815 -235
rect -1849 -269 -1815 -255
rect -1849 -323 -1815 -307
rect -1849 -341 -1815 -323
rect -1849 -391 -1815 -379
rect -1849 -413 -1815 -391
rect -1849 -459 -1815 -451
rect -1849 -485 -1815 -459
rect -1849 -527 -1815 -523
rect -1849 -557 -1815 -527
rect -1849 -629 -1815 -595
rect -1849 -697 -1815 -667
rect -1849 -701 -1815 -697
rect -1849 -765 -1815 -739
rect -1849 -773 -1815 -765
rect -1391 765 -1357 773
rect -1391 739 -1357 765
rect -1391 697 -1357 701
rect -1391 667 -1357 697
rect -1391 595 -1357 629
rect -1391 527 -1357 557
rect -1391 523 -1357 527
rect -1391 459 -1357 485
rect -1391 451 -1357 459
rect -1391 391 -1357 413
rect -1391 379 -1357 391
rect -1391 323 -1357 341
rect -1391 307 -1357 323
rect -1391 255 -1357 269
rect -1391 235 -1357 255
rect -1391 187 -1357 197
rect -1391 163 -1357 187
rect -1391 119 -1357 125
rect -1391 91 -1357 119
rect -1391 51 -1357 53
rect -1391 19 -1357 51
rect -1391 -51 -1357 -19
rect -1391 -53 -1357 -51
rect -1391 -119 -1357 -91
rect -1391 -125 -1357 -119
rect -1391 -187 -1357 -163
rect -1391 -197 -1357 -187
rect -1391 -255 -1357 -235
rect -1391 -269 -1357 -255
rect -1391 -323 -1357 -307
rect -1391 -341 -1357 -323
rect -1391 -391 -1357 -379
rect -1391 -413 -1357 -391
rect -1391 -459 -1357 -451
rect -1391 -485 -1357 -459
rect -1391 -527 -1357 -523
rect -1391 -557 -1357 -527
rect -1391 -629 -1357 -595
rect -1391 -697 -1357 -667
rect -1391 -701 -1357 -697
rect -1391 -765 -1357 -739
rect -1391 -773 -1357 -765
rect -933 765 -899 773
rect -933 739 -899 765
rect -933 697 -899 701
rect -933 667 -899 697
rect -933 595 -899 629
rect -933 527 -899 557
rect -933 523 -899 527
rect -933 459 -899 485
rect -933 451 -899 459
rect -933 391 -899 413
rect -933 379 -899 391
rect -933 323 -899 341
rect -933 307 -899 323
rect -933 255 -899 269
rect -933 235 -899 255
rect -933 187 -899 197
rect -933 163 -899 187
rect -933 119 -899 125
rect -933 91 -899 119
rect -933 51 -899 53
rect -933 19 -899 51
rect -933 -51 -899 -19
rect -933 -53 -899 -51
rect -933 -119 -899 -91
rect -933 -125 -899 -119
rect -933 -187 -899 -163
rect -933 -197 -899 -187
rect -933 -255 -899 -235
rect -933 -269 -899 -255
rect -933 -323 -899 -307
rect -933 -341 -899 -323
rect -933 -391 -899 -379
rect -933 -413 -899 -391
rect -933 -459 -899 -451
rect -933 -485 -899 -459
rect -933 -527 -899 -523
rect -933 -557 -899 -527
rect -933 -629 -899 -595
rect -933 -697 -899 -667
rect -933 -701 -899 -697
rect -933 -765 -899 -739
rect -933 -773 -899 -765
rect -475 765 -441 773
rect -475 739 -441 765
rect -475 697 -441 701
rect -475 667 -441 697
rect -475 595 -441 629
rect -475 527 -441 557
rect -475 523 -441 527
rect -475 459 -441 485
rect -475 451 -441 459
rect -475 391 -441 413
rect -475 379 -441 391
rect -475 323 -441 341
rect -475 307 -441 323
rect -475 255 -441 269
rect -475 235 -441 255
rect -475 187 -441 197
rect -475 163 -441 187
rect -475 119 -441 125
rect -475 91 -441 119
rect -475 51 -441 53
rect -475 19 -441 51
rect -475 -51 -441 -19
rect -475 -53 -441 -51
rect -475 -119 -441 -91
rect -475 -125 -441 -119
rect -475 -187 -441 -163
rect -475 -197 -441 -187
rect -475 -255 -441 -235
rect -475 -269 -441 -255
rect -475 -323 -441 -307
rect -475 -341 -441 -323
rect -475 -391 -441 -379
rect -475 -413 -441 -391
rect -475 -459 -441 -451
rect -475 -485 -441 -459
rect -475 -527 -441 -523
rect -475 -557 -441 -527
rect -475 -629 -441 -595
rect -475 -697 -441 -667
rect -475 -701 -441 -697
rect -475 -765 -441 -739
rect -475 -773 -441 -765
rect -17 765 17 773
rect -17 739 17 765
rect -17 697 17 701
rect -17 667 17 697
rect -17 595 17 629
rect -17 527 17 557
rect -17 523 17 527
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect -17 -527 17 -523
rect -17 -557 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -667
rect -17 -701 17 -697
rect -17 -765 17 -739
rect -17 -773 17 -765
rect 441 765 475 773
rect 441 739 475 765
rect 441 697 475 701
rect 441 667 475 697
rect 441 595 475 629
rect 441 527 475 557
rect 441 523 475 527
rect 441 459 475 485
rect 441 451 475 459
rect 441 391 475 413
rect 441 379 475 391
rect 441 323 475 341
rect 441 307 475 323
rect 441 255 475 269
rect 441 235 475 255
rect 441 187 475 197
rect 441 163 475 187
rect 441 119 475 125
rect 441 91 475 119
rect 441 51 475 53
rect 441 19 475 51
rect 441 -51 475 -19
rect 441 -53 475 -51
rect 441 -119 475 -91
rect 441 -125 475 -119
rect 441 -187 475 -163
rect 441 -197 475 -187
rect 441 -255 475 -235
rect 441 -269 475 -255
rect 441 -323 475 -307
rect 441 -341 475 -323
rect 441 -391 475 -379
rect 441 -413 475 -391
rect 441 -459 475 -451
rect 441 -485 475 -459
rect 441 -527 475 -523
rect 441 -557 475 -527
rect 441 -629 475 -595
rect 441 -697 475 -667
rect 441 -701 475 -697
rect 441 -765 475 -739
rect 441 -773 475 -765
rect 899 765 933 773
rect 899 739 933 765
rect 899 697 933 701
rect 899 667 933 697
rect 899 595 933 629
rect 899 527 933 557
rect 899 523 933 527
rect 899 459 933 485
rect 899 451 933 459
rect 899 391 933 413
rect 899 379 933 391
rect 899 323 933 341
rect 899 307 933 323
rect 899 255 933 269
rect 899 235 933 255
rect 899 187 933 197
rect 899 163 933 187
rect 899 119 933 125
rect 899 91 933 119
rect 899 51 933 53
rect 899 19 933 51
rect 899 -51 933 -19
rect 899 -53 933 -51
rect 899 -119 933 -91
rect 899 -125 933 -119
rect 899 -187 933 -163
rect 899 -197 933 -187
rect 899 -255 933 -235
rect 899 -269 933 -255
rect 899 -323 933 -307
rect 899 -341 933 -323
rect 899 -391 933 -379
rect 899 -413 933 -391
rect 899 -459 933 -451
rect 899 -485 933 -459
rect 899 -527 933 -523
rect 899 -557 933 -527
rect 899 -629 933 -595
rect 899 -697 933 -667
rect 899 -701 933 -697
rect 899 -765 933 -739
rect 899 -773 933 -765
rect 1357 765 1391 773
rect 1357 739 1391 765
rect 1357 697 1391 701
rect 1357 667 1391 697
rect 1357 595 1391 629
rect 1357 527 1391 557
rect 1357 523 1391 527
rect 1357 459 1391 485
rect 1357 451 1391 459
rect 1357 391 1391 413
rect 1357 379 1391 391
rect 1357 323 1391 341
rect 1357 307 1391 323
rect 1357 255 1391 269
rect 1357 235 1391 255
rect 1357 187 1391 197
rect 1357 163 1391 187
rect 1357 119 1391 125
rect 1357 91 1391 119
rect 1357 51 1391 53
rect 1357 19 1391 51
rect 1357 -51 1391 -19
rect 1357 -53 1391 -51
rect 1357 -119 1391 -91
rect 1357 -125 1391 -119
rect 1357 -187 1391 -163
rect 1357 -197 1391 -187
rect 1357 -255 1391 -235
rect 1357 -269 1391 -255
rect 1357 -323 1391 -307
rect 1357 -341 1391 -323
rect 1357 -391 1391 -379
rect 1357 -413 1391 -391
rect 1357 -459 1391 -451
rect 1357 -485 1391 -459
rect 1357 -527 1391 -523
rect 1357 -557 1391 -527
rect 1357 -629 1391 -595
rect 1357 -697 1391 -667
rect 1357 -701 1391 -697
rect 1357 -765 1391 -739
rect 1357 -773 1391 -765
rect 1815 765 1849 773
rect 1815 739 1849 765
rect 1815 697 1849 701
rect 1815 667 1849 697
rect 1815 595 1849 629
rect 1815 527 1849 557
rect 1815 523 1849 527
rect 1815 459 1849 485
rect 1815 451 1849 459
rect 1815 391 1849 413
rect 1815 379 1849 391
rect 1815 323 1849 341
rect 1815 307 1849 323
rect 1815 255 1849 269
rect 1815 235 1849 255
rect 1815 187 1849 197
rect 1815 163 1849 187
rect 1815 119 1849 125
rect 1815 91 1849 119
rect 1815 51 1849 53
rect 1815 19 1849 51
rect 1815 -51 1849 -19
rect 1815 -53 1849 -51
rect 1815 -119 1849 -91
rect 1815 -125 1849 -119
rect 1815 -187 1849 -163
rect 1815 -197 1849 -187
rect 1815 -255 1849 -235
rect 1815 -269 1849 -255
rect 1815 -323 1849 -307
rect 1815 -341 1849 -323
rect 1815 -391 1849 -379
rect 1815 -413 1849 -391
rect 1815 -459 1849 -451
rect 1815 -485 1849 -459
rect 1815 -527 1849 -523
rect 1815 -557 1849 -527
rect 1815 -629 1849 -595
rect 1815 -697 1849 -667
rect 1815 -701 1849 -697
rect 1815 -765 1849 -739
rect 1815 -773 1849 -765
rect 2273 765 2307 773
rect 2273 739 2307 765
rect 2273 697 2307 701
rect 2273 667 2307 697
rect 2273 595 2307 629
rect 2273 527 2307 557
rect 2273 523 2307 527
rect 2273 459 2307 485
rect 2273 451 2307 459
rect 2273 391 2307 413
rect 2273 379 2307 391
rect 2273 323 2307 341
rect 2273 307 2307 323
rect 2273 255 2307 269
rect 2273 235 2307 255
rect 2273 187 2307 197
rect 2273 163 2307 187
rect 2273 119 2307 125
rect 2273 91 2307 119
rect 2273 51 2307 53
rect 2273 19 2307 51
rect 2273 -51 2307 -19
rect 2273 -53 2307 -51
rect 2273 -119 2307 -91
rect 2273 -125 2307 -119
rect 2273 -187 2307 -163
rect 2273 -197 2307 -187
rect 2273 -255 2307 -235
rect 2273 -269 2307 -255
rect 2273 -323 2307 -307
rect 2273 -341 2307 -323
rect 2273 -391 2307 -379
rect 2273 -413 2307 -391
rect 2273 -459 2307 -451
rect 2273 -485 2307 -459
rect 2273 -527 2307 -523
rect 2273 -557 2307 -527
rect 2273 -629 2307 -595
rect 2273 -697 2307 -667
rect 2273 -701 2307 -697
rect 2273 -765 2307 -739
rect 2273 -773 2307 -765
rect 2731 765 2765 773
rect 2731 739 2765 765
rect 2731 697 2765 701
rect 2731 667 2765 697
rect 2731 595 2765 629
rect 2731 527 2765 557
rect 2731 523 2765 527
rect 2731 459 2765 485
rect 2731 451 2765 459
rect 2731 391 2765 413
rect 2731 379 2765 391
rect 2731 323 2765 341
rect 2731 307 2765 323
rect 2731 255 2765 269
rect 2731 235 2765 255
rect 2731 187 2765 197
rect 2731 163 2765 187
rect 2731 119 2765 125
rect 2731 91 2765 119
rect 2731 51 2765 53
rect 2731 19 2765 51
rect 2731 -51 2765 -19
rect 2731 -53 2765 -51
rect 2731 -119 2765 -91
rect 2731 -125 2765 -119
rect 2731 -187 2765 -163
rect 2731 -197 2765 -187
rect 2731 -255 2765 -235
rect 2731 -269 2765 -255
rect 2731 -323 2765 -307
rect 2731 -341 2765 -323
rect 2731 -391 2765 -379
rect 2731 -413 2765 -391
rect 2731 -459 2765 -451
rect 2731 -485 2765 -459
rect 2731 -527 2765 -523
rect 2731 -557 2765 -527
rect 2731 -629 2765 -595
rect 2731 -697 2765 -667
rect 2731 -701 2765 -697
rect 2731 -765 2765 -739
rect 2731 -773 2765 -765
rect 3189 765 3223 773
rect 3189 739 3223 765
rect 3189 697 3223 701
rect 3189 667 3223 697
rect 3189 595 3223 629
rect 3189 527 3223 557
rect 3189 523 3223 527
rect 3189 459 3223 485
rect 3189 451 3223 459
rect 3189 391 3223 413
rect 3189 379 3223 391
rect 3189 323 3223 341
rect 3189 307 3223 323
rect 3189 255 3223 269
rect 3189 235 3223 255
rect 3189 187 3223 197
rect 3189 163 3223 187
rect 3189 119 3223 125
rect 3189 91 3223 119
rect 3189 51 3223 53
rect 3189 19 3223 51
rect 3189 -51 3223 -19
rect 3189 -53 3223 -51
rect 3189 -119 3223 -91
rect 3189 -125 3223 -119
rect 3189 -187 3223 -163
rect 3189 -197 3223 -187
rect 3189 -255 3223 -235
rect 3189 -269 3223 -255
rect 3189 -323 3223 -307
rect 3189 -341 3223 -323
rect 3189 -391 3223 -379
rect 3189 -413 3223 -391
rect 3189 -459 3223 -451
rect 3189 -485 3223 -459
rect 3189 -527 3223 -523
rect 3189 -557 3223 -527
rect 3189 -629 3223 -595
rect 3189 -697 3223 -667
rect 3189 -701 3223 -697
rect 3189 -765 3223 -739
rect 3189 -773 3223 -765
rect 3647 765 3681 773
rect 3647 739 3681 765
rect 3647 697 3681 701
rect 3647 667 3681 697
rect 3647 595 3681 629
rect 3647 527 3681 557
rect 3647 523 3681 527
rect 3647 459 3681 485
rect 3647 451 3681 459
rect 3647 391 3681 413
rect 3647 379 3681 391
rect 3647 323 3681 341
rect 3647 307 3681 323
rect 3647 255 3681 269
rect 3647 235 3681 255
rect 3647 187 3681 197
rect 3647 163 3681 187
rect 3647 119 3681 125
rect 3647 91 3681 119
rect 3647 51 3681 53
rect 3647 19 3681 51
rect 3647 -51 3681 -19
rect 3647 -53 3681 -51
rect 3647 -119 3681 -91
rect 3647 -125 3681 -119
rect 3647 -187 3681 -163
rect 3647 -197 3681 -187
rect 3647 -255 3681 -235
rect 3647 -269 3681 -255
rect 3647 -323 3681 -307
rect 3647 -341 3681 -323
rect 3647 -391 3681 -379
rect 3647 -413 3681 -391
rect 3647 -459 3681 -451
rect 3647 -485 3681 -459
rect 3647 -527 3681 -523
rect 3647 -557 3681 -527
rect 3647 -629 3681 -595
rect 3647 -697 3681 -667
rect 3647 -701 3681 -697
rect 3647 -765 3681 -739
rect 3647 -773 3681 -765
rect 4105 765 4139 773
rect 4105 739 4139 765
rect 4105 697 4139 701
rect 4105 667 4139 697
rect 4105 595 4139 629
rect 4105 527 4139 557
rect 4105 523 4139 527
rect 4105 459 4139 485
rect 4105 451 4139 459
rect 4105 391 4139 413
rect 4105 379 4139 391
rect 4105 323 4139 341
rect 4105 307 4139 323
rect 4105 255 4139 269
rect 4105 235 4139 255
rect 4105 187 4139 197
rect 4105 163 4139 187
rect 4105 119 4139 125
rect 4105 91 4139 119
rect 4105 51 4139 53
rect 4105 19 4139 51
rect 4105 -51 4139 -19
rect 4105 -53 4139 -51
rect 4105 -119 4139 -91
rect 4105 -125 4139 -119
rect 4105 -187 4139 -163
rect 4105 -197 4139 -187
rect 4105 -255 4139 -235
rect 4105 -269 4139 -255
rect 4105 -323 4139 -307
rect 4105 -341 4139 -323
rect 4105 -391 4139 -379
rect 4105 -413 4139 -391
rect 4105 -459 4139 -451
rect 4105 -485 4139 -459
rect 4105 -527 4139 -523
rect 4105 -557 4139 -527
rect 4105 -629 4139 -595
rect 4105 -697 4139 -667
rect 4105 -701 4139 -697
rect 4105 -765 4139 -739
rect 4105 -773 4139 -765
rect -3982 -881 -3978 -847
rect -3978 -881 -3948 -847
rect -3910 -881 -3876 -847
rect -3838 -881 -3808 -847
rect -3808 -881 -3804 -847
rect -3524 -881 -3520 -847
rect -3520 -881 -3490 -847
rect -3452 -881 -3418 -847
rect -3380 -881 -3350 -847
rect -3350 -881 -3346 -847
rect -3066 -881 -3062 -847
rect -3062 -881 -3032 -847
rect -2994 -881 -2960 -847
rect -2922 -881 -2892 -847
rect -2892 -881 -2888 -847
rect -2608 -881 -2604 -847
rect -2604 -881 -2574 -847
rect -2536 -881 -2502 -847
rect -2464 -881 -2434 -847
rect -2434 -881 -2430 -847
rect -2150 -881 -2146 -847
rect -2146 -881 -2116 -847
rect -2078 -881 -2044 -847
rect -2006 -881 -1976 -847
rect -1976 -881 -1972 -847
rect -1692 -881 -1688 -847
rect -1688 -881 -1658 -847
rect -1620 -881 -1586 -847
rect -1548 -881 -1518 -847
rect -1518 -881 -1514 -847
rect -1234 -881 -1230 -847
rect -1230 -881 -1200 -847
rect -1162 -881 -1128 -847
rect -1090 -881 -1060 -847
rect -1060 -881 -1056 -847
rect -776 -881 -772 -847
rect -772 -881 -742 -847
rect -704 -881 -670 -847
rect -632 -881 -602 -847
rect -602 -881 -598 -847
rect -318 -881 -314 -847
rect -314 -881 -284 -847
rect -246 -881 -212 -847
rect -174 -881 -144 -847
rect -144 -881 -140 -847
rect 140 -881 144 -847
rect 144 -881 174 -847
rect 212 -881 246 -847
rect 284 -881 314 -847
rect 314 -881 318 -847
rect 598 -881 602 -847
rect 602 -881 632 -847
rect 670 -881 704 -847
rect 742 -881 772 -847
rect 772 -881 776 -847
rect 1056 -881 1060 -847
rect 1060 -881 1090 -847
rect 1128 -881 1162 -847
rect 1200 -881 1230 -847
rect 1230 -881 1234 -847
rect 1514 -881 1518 -847
rect 1518 -881 1548 -847
rect 1586 -881 1620 -847
rect 1658 -881 1688 -847
rect 1688 -881 1692 -847
rect 1972 -881 1976 -847
rect 1976 -881 2006 -847
rect 2044 -881 2078 -847
rect 2116 -881 2146 -847
rect 2146 -881 2150 -847
rect 2430 -881 2434 -847
rect 2434 -881 2464 -847
rect 2502 -881 2536 -847
rect 2574 -881 2604 -847
rect 2604 -881 2608 -847
rect 2888 -881 2892 -847
rect 2892 -881 2922 -847
rect 2960 -881 2994 -847
rect 3032 -881 3062 -847
rect 3062 -881 3066 -847
rect 3346 -881 3350 -847
rect 3350 -881 3380 -847
rect 3418 -881 3452 -847
rect 3490 -881 3520 -847
rect 3520 -881 3524 -847
rect 3804 -881 3808 -847
rect 3808 -881 3838 -847
rect 3876 -881 3910 -847
rect 3948 -881 3978 -847
rect 3978 -881 3982 -847
<< metal1 >>
rect -3997 881 -3789 887
rect -3997 847 -3982 881
rect -3948 847 -3910 881
rect -3876 847 -3838 881
rect -3804 847 -3789 881
rect -3997 841 -3789 847
rect -3539 881 -3331 887
rect -3539 847 -3524 881
rect -3490 847 -3452 881
rect -3418 847 -3380 881
rect -3346 847 -3331 881
rect -3539 841 -3331 847
rect -3081 881 -2873 887
rect -3081 847 -3066 881
rect -3032 847 -2994 881
rect -2960 847 -2922 881
rect -2888 847 -2873 881
rect -3081 841 -2873 847
rect -2623 881 -2415 887
rect -2623 847 -2608 881
rect -2574 847 -2536 881
rect -2502 847 -2464 881
rect -2430 847 -2415 881
rect -2623 841 -2415 847
rect -2165 881 -1957 887
rect -2165 847 -2150 881
rect -2116 847 -2078 881
rect -2044 847 -2006 881
rect -1972 847 -1957 881
rect -2165 841 -1957 847
rect -1707 881 -1499 887
rect -1707 847 -1692 881
rect -1658 847 -1620 881
rect -1586 847 -1548 881
rect -1514 847 -1499 881
rect -1707 841 -1499 847
rect -1249 881 -1041 887
rect -1249 847 -1234 881
rect -1200 847 -1162 881
rect -1128 847 -1090 881
rect -1056 847 -1041 881
rect -1249 841 -1041 847
rect -791 881 -583 887
rect -791 847 -776 881
rect -742 847 -704 881
rect -670 847 -632 881
rect -598 847 -583 881
rect -791 841 -583 847
rect -333 881 -125 887
rect -333 847 -318 881
rect -284 847 -246 881
rect -212 847 -174 881
rect -140 847 -125 881
rect -333 841 -125 847
rect 125 881 333 887
rect 125 847 140 881
rect 174 847 212 881
rect 246 847 284 881
rect 318 847 333 881
rect 125 841 333 847
rect 583 881 791 887
rect 583 847 598 881
rect 632 847 670 881
rect 704 847 742 881
rect 776 847 791 881
rect 583 841 791 847
rect 1041 881 1249 887
rect 1041 847 1056 881
rect 1090 847 1128 881
rect 1162 847 1200 881
rect 1234 847 1249 881
rect 1041 841 1249 847
rect 1499 881 1707 887
rect 1499 847 1514 881
rect 1548 847 1586 881
rect 1620 847 1658 881
rect 1692 847 1707 881
rect 1499 841 1707 847
rect 1957 881 2165 887
rect 1957 847 1972 881
rect 2006 847 2044 881
rect 2078 847 2116 881
rect 2150 847 2165 881
rect 1957 841 2165 847
rect 2415 881 2623 887
rect 2415 847 2430 881
rect 2464 847 2502 881
rect 2536 847 2574 881
rect 2608 847 2623 881
rect 2415 841 2623 847
rect 2873 881 3081 887
rect 2873 847 2888 881
rect 2922 847 2960 881
rect 2994 847 3032 881
rect 3066 847 3081 881
rect 2873 841 3081 847
rect 3331 881 3539 887
rect 3331 847 3346 881
rect 3380 847 3418 881
rect 3452 847 3490 881
rect 3524 847 3539 881
rect 3331 841 3539 847
rect 3789 881 3997 887
rect 3789 847 3804 881
rect 3838 847 3876 881
rect 3910 847 3948 881
rect 3982 847 3997 881
rect 3789 841 3997 847
rect -4145 773 -4099 800
rect -4145 739 -4139 773
rect -4105 739 -4099 773
rect -4145 701 -4099 739
rect -4145 667 -4139 701
rect -4105 667 -4099 701
rect -4145 629 -4099 667
rect -4145 595 -4139 629
rect -4105 595 -4099 629
rect -4145 557 -4099 595
rect -4145 523 -4139 557
rect -4105 523 -4099 557
rect -4145 485 -4099 523
rect -4145 451 -4139 485
rect -4105 451 -4099 485
rect -4145 413 -4099 451
rect -4145 379 -4139 413
rect -4105 379 -4099 413
rect -4145 341 -4099 379
rect -4145 307 -4139 341
rect -4105 307 -4099 341
rect -4145 269 -4099 307
rect -4145 235 -4139 269
rect -4105 235 -4099 269
rect -4145 197 -4099 235
rect -4145 163 -4139 197
rect -4105 163 -4099 197
rect -4145 125 -4099 163
rect -4145 91 -4139 125
rect -4105 91 -4099 125
rect -4145 53 -4099 91
rect -4145 19 -4139 53
rect -4105 19 -4099 53
rect -4145 -19 -4099 19
rect -4145 -53 -4139 -19
rect -4105 -53 -4099 -19
rect -4145 -91 -4099 -53
rect -4145 -125 -4139 -91
rect -4105 -125 -4099 -91
rect -4145 -163 -4099 -125
rect -4145 -197 -4139 -163
rect -4105 -197 -4099 -163
rect -4145 -235 -4099 -197
rect -4145 -269 -4139 -235
rect -4105 -269 -4099 -235
rect -4145 -307 -4099 -269
rect -4145 -341 -4139 -307
rect -4105 -341 -4099 -307
rect -4145 -379 -4099 -341
rect -4145 -413 -4139 -379
rect -4105 -413 -4099 -379
rect -4145 -451 -4099 -413
rect -4145 -485 -4139 -451
rect -4105 -485 -4099 -451
rect -4145 -523 -4099 -485
rect -4145 -557 -4139 -523
rect -4105 -557 -4099 -523
rect -4145 -595 -4099 -557
rect -4145 -629 -4139 -595
rect -4105 -629 -4099 -595
rect -4145 -667 -4099 -629
rect -4145 -701 -4139 -667
rect -4105 -701 -4099 -667
rect -4145 -739 -4099 -701
rect -4145 -773 -4139 -739
rect -4105 -773 -4099 -739
rect -4145 -800 -4099 -773
rect -3687 773 -3641 800
rect -3687 739 -3681 773
rect -3647 739 -3641 773
rect -3687 701 -3641 739
rect -3687 667 -3681 701
rect -3647 667 -3641 701
rect -3687 629 -3641 667
rect -3687 595 -3681 629
rect -3647 595 -3641 629
rect -3687 557 -3641 595
rect -3687 523 -3681 557
rect -3647 523 -3641 557
rect -3687 485 -3641 523
rect -3687 451 -3681 485
rect -3647 451 -3641 485
rect -3687 413 -3641 451
rect -3687 379 -3681 413
rect -3647 379 -3641 413
rect -3687 341 -3641 379
rect -3687 307 -3681 341
rect -3647 307 -3641 341
rect -3687 269 -3641 307
rect -3687 235 -3681 269
rect -3647 235 -3641 269
rect -3687 197 -3641 235
rect -3687 163 -3681 197
rect -3647 163 -3641 197
rect -3687 125 -3641 163
rect -3687 91 -3681 125
rect -3647 91 -3641 125
rect -3687 53 -3641 91
rect -3687 19 -3681 53
rect -3647 19 -3641 53
rect -3687 -19 -3641 19
rect -3687 -53 -3681 -19
rect -3647 -53 -3641 -19
rect -3687 -91 -3641 -53
rect -3687 -125 -3681 -91
rect -3647 -125 -3641 -91
rect -3687 -163 -3641 -125
rect -3687 -197 -3681 -163
rect -3647 -197 -3641 -163
rect -3687 -235 -3641 -197
rect -3687 -269 -3681 -235
rect -3647 -269 -3641 -235
rect -3687 -307 -3641 -269
rect -3687 -341 -3681 -307
rect -3647 -341 -3641 -307
rect -3687 -379 -3641 -341
rect -3687 -413 -3681 -379
rect -3647 -413 -3641 -379
rect -3687 -451 -3641 -413
rect -3687 -485 -3681 -451
rect -3647 -485 -3641 -451
rect -3687 -523 -3641 -485
rect -3687 -557 -3681 -523
rect -3647 -557 -3641 -523
rect -3687 -595 -3641 -557
rect -3687 -629 -3681 -595
rect -3647 -629 -3641 -595
rect -3687 -667 -3641 -629
rect -3687 -701 -3681 -667
rect -3647 -701 -3641 -667
rect -3687 -739 -3641 -701
rect -3687 -773 -3681 -739
rect -3647 -773 -3641 -739
rect -3687 -800 -3641 -773
rect -3229 773 -3183 800
rect -3229 739 -3223 773
rect -3189 739 -3183 773
rect -3229 701 -3183 739
rect -3229 667 -3223 701
rect -3189 667 -3183 701
rect -3229 629 -3183 667
rect -3229 595 -3223 629
rect -3189 595 -3183 629
rect -3229 557 -3183 595
rect -3229 523 -3223 557
rect -3189 523 -3183 557
rect -3229 485 -3183 523
rect -3229 451 -3223 485
rect -3189 451 -3183 485
rect -3229 413 -3183 451
rect -3229 379 -3223 413
rect -3189 379 -3183 413
rect -3229 341 -3183 379
rect -3229 307 -3223 341
rect -3189 307 -3183 341
rect -3229 269 -3183 307
rect -3229 235 -3223 269
rect -3189 235 -3183 269
rect -3229 197 -3183 235
rect -3229 163 -3223 197
rect -3189 163 -3183 197
rect -3229 125 -3183 163
rect -3229 91 -3223 125
rect -3189 91 -3183 125
rect -3229 53 -3183 91
rect -3229 19 -3223 53
rect -3189 19 -3183 53
rect -3229 -19 -3183 19
rect -3229 -53 -3223 -19
rect -3189 -53 -3183 -19
rect -3229 -91 -3183 -53
rect -3229 -125 -3223 -91
rect -3189 -125 -3183 -91
rect -3229 -163 -3183 -125
rect -3229 -197 -3223 -163
rect -3189 -197 -3183 -163
rect -3229 -235 -3183 -197
rect -3229 -269 -3223 -235
rect -3189 -269 -3183 -235
rect -3229 -307 -3183 -269
rect -3229 -341 -3223 -307
rect -3189 -341 -3183 -307
rect -3229 -379 -3183 -341
rect -3229 -413 -3223 -379
rect -3189 -413 -3183 -379
rect -3229 -451 -3183 -413
rect -3229 -485 -3223 -451
rect -3189 -485 -3183 -451
rect -3229 -523 -3183 -485
rect -3229 -557 -3223 -523
rect -3189 -557 -3183 -523
rect -3229 -595 -3183 -557
rect -3229 -629 -3223 -595
rect -3189 -629 -3183 -595
rect -3229 -667 -3183 -629
rect -3229 -701 -3223 -667
rect -3189 -701 -3183 -667
rect -3229 -739 -3183 -701
rect -3229 -773 -3223 -739
rect -3189 -773 -3183 -739
rect -3229 -800 -3183 -773
rect -2771 773 -2725 800
rect -2771 739 -2765 773
rect -2731 739 -2725 773
rect -2771 701 -2725 739
rect -2771 667 -2765 701
rect -2731 667 -2725 701
rect -2771 629 -2725 667
rect -2771 595 -2765 629
rect -2731 595 -2725 629
rect -2771 557 -2725 595
rect -2771 523 -2765 557
rect -2731 523 -2725 557
rect -2771 485 -2725 523
rect -2771 451 -2765 485
rect -2731 451 -2725 485
rect -2771 413 -2725 451
rect -2771 379 -2765 413
rect -2731 379 -2725 413
rect -2771 341 -2725 379
rect -2771 307 -2765 341
rect -2731 307 -2725 341
rect -2771 269 -2725 307
rect -2771 235 -2765 269
rect -2731 235 -2725 269
rect -2771 197 -2725 235
rect -2771 163 -2765 197
rect -2731 163 -2725 197
rect -2771 125 -2725 163
rect -2771 91 -2765 125
rect -2731 91 -2725 125
rect -2771 53 -2725 91
rect -2771 19 -2765 53
rect -2731 19 -2725 53
rect -2771 -19 -2725 19
rect -2771 -53 -2765 -19
rect -2731 -53 -2725 -19
rect -2771 -91 -2725 -53
rect -2771 -125 -2765 -91
rect -2731 -125 -2725 -91
rect -2771 -163 -2725 -125
rect -2771 -197 -2765 -163
rect -2731 -197 -2725 -163
rect -2771 -235 -2725 -197
rect -2771 -269 -2765 -235
rect -2731 -269 -2725 -235
rect -2771 -307 -2725 -269
rect -2771 -341 -2765 -307
rect -2731 -341 -2725 -307
rect -2771 -379 -2725 -341
rect -2771 -413 -2765 -379
rect -2731 -413 -2725 -379
rect -2771 -451 -2725 -413
rect -2771 -485 -2765 -451
rect -2731 -485 -2725 -451
rect -2771 -523 -2725 -485
rect -2771 -557 -2765 -523
rect -2731 -557 -2725 -523
rect -2771 -595 -2725 -557
rect -2771 -629 -2765 -595
rect -2731 -629 -2725 -595
rect -2771 -667 -2725 -629
rect -2771 -701 -2765 -667
rect -2731 -701 -2725 -667
rect -2771 -739 -2725 -701
rect -2771 -773 -2765 -739
rect -2731 -773 -2725 -739
rect -2771 -800 -2725 -773
rect -2313 773 -2267 800
rect -2313 739 -2307 773
rect -2273 739 -2267 773
rect -2313 701 -2267 739
rect -2313 667 -2307 701
rect -2273 667 -2267 701
rect -2313 629 -2267 667
rect -2313 595 -2307 629
rect -2273 595 -2267 629
rect -2313 557 -2267 595
rect -2313 523 -2307 557
rect -2273 523 -2267 557
rect -2313 485 -2267 523
rect -2313 451 -2307 485
rect -2273 451 -2267 485
rect -2313 413 -2267 451
rect -2313 379 -2307 413
rect -2273 379 -2267 413
rect -2313 341 -2267 379
rect -2313 307 -2307 341
rect -2273 307 -2267 341
rect -2313 269 -2267 307
rect -2313 235 -2307 269
rect -2273 235 -2267 269
rect -2313 197 -2267 235
rect -2313 163 -2307 197
rect -2273 163 -2267 197
rect -2313 125 -2267 163
rect -2313 91 -2307 125
rect -2273 91 -2267 125
rect -2313 53 -2267 91
rect -2313 19 -2307 53
rect -2273 19 -2267 53
rect -2313 -19 -2267 19
rect -2313 -53 -2307 -19
rect -2273 -53 -2267 -19
rect -2313 -91 -2267 -53
rect -2313 -125 -2307 -91
rect -2273 -125 -2267 -91
rect -2313 -163 -2267 -125
rect -2313 -197 -2307 -163
rect -2273 -197 -2267 -163
rect -2313 -235 -2267 -197
rect -2313 -269 -2307 -235
rect -2273 -269 -2267 -235
rect -2313 -307 -2267 -269
rect -2313 -341 -2307 -307
rect -2273 -341 -2267 -307
rect -2313 -379 -2267 -341
rect -2313 -413 -2307 -379
rect -2273 -413 -2267 -379
rect -2313 -451 -2267 -413
rect -2313 -485 -2307 -451
rect -2273 -485 -2267 -451
rect -2313 -523 -2267 -485
rect -2313 -557 -2307 -523
rect -2273 -557 -2267 -523
rect -2313 -595 -2267 -557
rect -2313 -629 -2307 -595
rect -2273 -629 -2267 -595
rect -2313 -667 -2267 -629
rect -2313 -701 -2307 -667
rect -2273 -701 -2267 -667
rect -2313 -739 -2267 -701
rect -2313 -773 -2307 -739
rect -2273 -773 -2267 -739
rect -2313 -800 -2267 -773
rect -1855 773 -1809 800
rect -1855 739 -1849 773
rect -1815 739 -1809 773
rect -1855 701 -1809 739
rect -1855 667 -1849 701
rect -1815 667 -1809 701
rect -1855 629 -1809 667
rect -1855 595 -1849 629
rect -1815 595 -1809 629
rect -1855 557 -1809 595
rect -1855 523 -1849 557
rect -1815 523 -1809 557
rect -1855 485 -1809 523
rect -1855 451 -1849 485
rect -1815 451 -1809 485
rect -1855 413 -1809 451
rect -1855 379 -1849 413
rect -1815 379 -1809 413
rect -1855 341 -1809 379
rect -1855 307 -1849 341
rect -1815 307 -1809 341
rect -1855 269 -1809 307
rect -1855 235 -1849 269
rect -1815 235 -1809 269
rect -1855 197 -1809 235
rect -1855 163 -1849 197
rect -1815 163 -1809 197
rect -1855 125 -1809 163
rect -1855 91 -1849 125
rect -1815 91 -1809 125
rect -1855 53 -1809 91
rect -1855 19 -1849 53
rect -1815 19 -1809 53
rect -1855 -19 -1809 19
rect -1855 -53 -1849 -19
rect -1815 -53 -1809 -19
rect -1855 -91 -1809 -53
rect -1855 -125 -1849 -91
rect -1815 -125 -1809 -91
rect -1855 -163 -1809 -125
rect -1855 -197 -1849 -163
rect -1815 -197 -1809 -163
rect -1855 -235 -1809 -197
rect -1855 -269 -1849 -235
rect -1815 -269 -1809 -235
rect -1855 -307 -1809 -269
rect -1855 -341 -1849 -307
rect -1815 -341 -1809 -307
rect -1855 -379 -1809 -341
rect -1855 -413 -1849 -379
rect -1815 -413 -1809 -379
rect -1855 -451 -1809 -413
rect -1855 -485 -1849 -451
rect -1815 -485 -1809 -451
rect -1855 -523 -1809 -485
rect -1855 -557 -1849 -523
rect -1815 -557 -1809 -523
rect -1855 -595 -1809 -557
rect -1855 -629 -1849 -595
rect -1815 -629 -1809 -595
rect -1855 -667 -1809 -629
rect -1855 -701 -1849 -667
rect -1815 -701 -1809 -667
rect -1855 -739 -1809 -701
rect -1855 -773 -1849 -739
rect -1815 -773 -1809 -739
rect -1855 -800 -1809 -773
rect -1397 773 -1351 800
rect -1397 739 -1391 773
rect -1357 739 -1351 773
rect -1397 701 -1351 739
rect -1397 667 -1391 701
rect -1357 667 -1351 701
rect -1397 629 -1351 667
rect -1397 595 -1391 629
rect -1357 595 -1351 629
rect -1397 557 -1351 595
rect -1397 523 -1391 557
rect -1357 523 -1351 557
rect -1397 485 -1351 523
rect -1397 451 -1391 485
rect -1357 451 -1351 485
rect -1397 413 -1351 451
rect -1397 379 -1391 413
rect -1357 379 -1351 413
rect -1397 341 -1351 379
rect -1397 307 -1391 341
rect -1357 307 -1351 341
rect -1397 269 -1351 307
rect -1397 235 -1391 269
rect -1357 235 -1351 269
rect -1397 197 -1351 235
rect -1397 163 -1391 197
rect -1357 163 -1351 197
rect -1397 125 -1351 163
rect -1397 91 -1391 125
rect -1357 91 -1351 125
rect -1397 53 -1351 91
rect -1397 19 -1391 53
rect -1357 19 -1351 53
rect -1397 -19 -1351 19
rect -1397 -53 -1391 -19
rect -1357 -53 -1351 -19
rect -1397 -91 -1351 -53
rect -1397 -125 -1391 -91
rect -1357 -125 -1351 -91
rect -1397 -163 -1351 -125
rect -1397 -197 -1391 -163
rect -1357 -197 -1351 -163
rect -1397 -235 -1351 -197
rect -1397 -269 -1391 -235
rect -1357 -269 -1351 -235
rect -1397 -307 -1351 -269
rect -1397 -341 -1391 -307
rect -1357 -341 -1351 -307
rect -1397 -379 -1351 -341
rect -1397 -413 -1391 -379
rect -1357 -413 -1351 -379
rect -1397 -451 -1351 -413
rect -1397 -485 -1391 -451
rect -1357 -485 -1351 -451
rect -1397 -523 -1351 -485
rect -1397 -557 -1391 -523
rect -1357 -557 -1351 -523
rect -1397 -595 -1351 -557
rect -1397 -629 -1391 -595
rect -1357 -629 -1351 -595
rect -1397 -667 -1351 -629
rect -1397 -701 -1391 -667
rect -1357 -701 -1351 -667
rect -1397 -739 -1351 -701
rect -1397 -773 -1391 -739
rect -1357 -773 -1351 -739
rect -1397 -800 -1351 -773
rect -939 773 -893 800
rect -939 739 -933 773
rect -899 739 -893 773
rect -939 701 -893 739
rect -939 667 -933 701
rect -899 667 -893 701
rect -939 629 -893 667
rect -939 595 -933 629
rect -899 595 -893 629
rect -939 557 -893 595
rect -939 523 -933 557
rect -899 523 -893 557
rect -939 485 -893 523
rect -939 451 -933 485
rect -899 451 -893 485
rect -939 413 -893 451
rect -939 379 -933 413
rect -899 379 -893 413
rect -939 341 -893 379
rect -939 307 -933 341
rect -899 307 -893 341
rect -939 269 -893 307
rect -939 235 -933 269
rect -899 235 -893 269
rect -939 197 -893 235
rect -939 163 -933 197
rect -899 163 -893 197
rect -939 125 -893 163
rect -939 91 -933 125
rect -899 91 -893 125
rect -939 53 -893 91
rect -939 19 -933 53
rect -899 19 -893 53
rect -939 -19 -893 19
rect -939 -53 -933 -19
rect -899 -53 -893 -19
rect -939 -91 -893 -53
rect -939 -125 -933 -91
rect -899 -125 -893 -91
rect -939 -163 -893 -125
rect -939 -197 -933 -163
rect -899 -197 -893 -163
rect -939 -235 -893 -197
rect -939 -269 -933 -235
rect -899 -269 -893 -235
rect -939 -307 -893 -269
rect -939 -341 -933 -307
rect -899 -341 -893 -307
rect -939 -379 -893 -341
rect -939 -413 -933 -379
rect -899 -413 -893 -379
rect -939 -451 -893 -413
rect -939 -485 -933 -451
rect -899 -485 -893 -451
rect -939 -523 -893 -485
rect -939 -557 -933 -523
rect -899 -557 -893 -523
rect -939 -595 -893 -557
rect -939 -629 -933 -595
rect -899 -629 -893 -595
rect -939 -667 -893 -629
rect -939 -701 -933 -667
rect -899 -701 -893 -667
rect -939 -739 -893 -701
rect -939 -773 -933 -739
rect -899 -773 -893 -739
rect -939 -800 -893 -773
rect -481 773 -435 800
rect -481 739 -475 773
rect -441 739 -435 773
rect -481 701 -435 739
rect -481 667 -475 701
rect -441 667 -435 701
rect -481 629 -435 667
rect -481 595 -475 629
rect -441 595 -435 629
rect -481 557 -435 595
rect -481 523 -475 557
rect -441 523 -435 557
rect -481 485 -435 523
rect -481 451 -475 485
rect -441 451 -435 485
rect -481 413 -435 451
rect -481 379 -475 413
rect -441 379 -435 413
rect -481 341 -435 379
rect -481 307 -475 341
rect -441 307 -435 341
rect -481 269 -435 307
rect -481 235 -475 269
rect -441 235 -435 269
rect -481 197 -435 235
rect -481 163 -475 197
rect -441 163 -435 197
rect -481 125 -435 163
rect -481 91 -475 125
rect -441 91 -435 125
rect -481 53 -435 91
rect -481 19 -475 53
rect -441 19 -435 53
rect -481 -19 -435 19
rect -481 -53 -475 -19
rect -441 -53 -435 -19
rect -481 -91 -435 -53
rect -481 -125 -475 -91
rect -441 -125 -435 -91
rect -481 -163 -435 -125
rect -481 -197 -475 -163
rect -441 -197 -435 -163
rect -481 -235 -435 -197
rect -481 -269 -475 -235
rect -441 -269 -435 -235
rect -481 -307 -435 -269
rect -481 -341 -475 -307
rect -441 -341 -435 -307
rect -481 -379 -435 -341
rect -481 -413 -475 -379
rect -441 -413 -435 -379
rect -481 -451 -435 -413
rect -481 -485 -475 -451
rect -441 -485 -435 -451
rect -481 -523 -435 -485
rect -481 -557 -475 -523
rect -441 -557 -435 -523
rect -481 -595 -435 -557
rect -481 -629 -475 -595
rect -441 -629 -435 -595
rect -481 -667 -435 -629
rect -481 -701 -475 -667
rect -441 -701 -435 -667
rect -481 -739 -435 -701
rect -481 -773 -475 -739
rect -441 -773 -435 -739
rect -481 -800 -435 -773
rect -23 773 23 800
rect -23 739 -17 773
rect 17 739 23 773
rect -23 701 23 739
rect -23 667 -17 701
rect 17 667 23 701
rect -23 629 23 667
rect -23 595 -17 629
rect 17 595 23 629
rect -23 557 23 595
rect -23 523 -17 557
rect 17 523 23 557
rect -23 485 23 523
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -523 23 -485
rect -23 -557 -17 -523
rect 17 -557 23 -523
rect -23 -595 23 -557
rect -23 -629 -17 -595
rect 17 -629 23 -595
rect -23 -667 23 -629
rect -23 -701 -17 -667
rect 17 -701 23 -667
rect -23 -739 23 -701
rect -23 -773 -17 -739
rect 17 -773 23 -739
rect -23 -800 23 -773
rect 435 773 481 800
rect 435 739 441 773
rect 475 739 481 773
rect 435 701 481 739
rect 435 667 441 701
rect 475 667 481 701
rect 435 629 481 667
rect 435 595 441 629
rect 475 595 481 629
rect 435 557 481 595
rect 435 523 441 557
rect 475 523 481 557
rect 435 485 481 523
rect 435 451 441 485
rect 475 451 481 485
rect 435 413 481 451
rect 435 379 441 413
rect 475 379 481 413
rect 435 341 481 379
rect 435 307 441 341
rect 475 307 481 341
rect 435 269 481 307
rect 435 235 441 269
rect 475 235 481 269
rect 435 197 481 235
rect 435 163 441 197
rect 475 163 481 197
rect 435 125 481 163
rect 435 91 441 125
rect 475 91 481 125
rect 435 53 481 91
rect 435 19 441 53
rect 475 19 481 53
rect 435 -19 481 19
rect 435 -53 441 -19
rect 475 -53 481 -19
rect 435 -91 481 -53
rect 435 -125 441 -91
rect 475 -125 481 -91
rect 435 -163 481 -125
rect 435 -197 441 -163
rect 475 -197 481 -163
rect 435 -235 481 -197
rect 435 -269 441 -235
rect 475 -269 481 -235
rect 435 -307 481 -269
rect 435 -341 441 -307
rect 475 -341 481 -307
rect 435 -379 481 -341
rect 435 -413 441 -379
rect 475 -413 481 -379
rect 435 -451 481 -413
rect 435 -485 441 -451
rect 475 -485 481 -451
rect 435 -523 481 -485
rect 435 -557 441 -523
rect 475 -557 481 -523
rect 435 -595 481 -557
rect 435 -629 441 -595
rect 475 -629 481 -595
rect 435 -667 481 -629
rect 435 -701 441 -667
rect 475 -701 481 -667
rect 435 -739 481 -701
rect 435 -773 441 -739
rect 475 -773 481 -739
rect 435 -800 481 -773
rect 893 773 939 800
rect 893 739 899 773
rect 933 739 939 773
rect 893 701 939 739
rect 893 667 899 701
rect 933 667 939 701
rect 893 629 939 667
rect 893 595 899 629
rect 933 595 939 629
rect 893 557 939 595
rect 893 523 899 557
rect 933 523 939 557
rect 893 485 939 523
rect 893 451 899 485
rect 933 451 939 485
rect 893 413 939 451
rect 893 379 899 413
rect 933 379 939 413
rect 893 341 939 379
rect 893 307 899 341
rect 933 307 939 341
rect 893 269 939 307
rect 893 235 899 269
rect 933 235 939 269
rect 893 197 939 235
rect 893 163 899 197
rect 933 163 939 197
rect 893 125 939 163
rect 893 91 899 125
rect 933 91 939 125
rect 893 53 939 91
rect 893 19 899 53
rect 933 19 939 53
rect 893 -19 939 19
rect 893 -53 899 -19
rect 933 -53 939 -19
rect 893 -91 939 -53
rect 893 -125 899 -91
rect 933 -125 939 -91
rect 893 -163 939 -125
rect 893 -197 899 -163
rect 933 -197 939 -163
rect 893 -235 939 -197
rect 893 -269 899 -235
rect 933 -269 939 -235
rect 893 -307 939 -269
rect 893 -341 899 -307
rect 933 -341 939 -307
rect 893 -379 939 -341
rect 893 -413 899 -379
rect 933 -413 939 -379
rect 893 -451 939 -413
rect 893 -485 899 -451
rect 933 -485 939 -451
rect 893 -523 939 -485
rect 893 -557 899 -523
rect 933 -557 939 -523
rect 893 -595 939 -557
rect 893 -629 899 -595
rect 933 -629 939 -595
rect 893 -667 939 -629
rect 893 -701 899 -667
rect 933 -701 939 -667
rect 893 -739 939 -701
rect 893 -773 899 -739
rect 933 -773 939 -739
rect 893 -800 939 -773
rect 1351 773 1397 800
rect 1351 739 1357 773
rect 1391 739 1397 773
rect 1351 701 1397 739
rect 1351 667 1357 701
rect 1391 667 1397 701
rect 1351 629 1397 667
rect 1351 595 1357 629
rect 1391 595 1397 629
rect 1351 557 1397 595
rect 1351 523 1357 557
rect 1391 523 1397 557
rect 1351 485 1397 523
rect 1351 451 1357 485
rect 1391 451 1397 485
rect 1351 413 1397 451
rect 1351 379 1357 413
rect 1391 379 1397 413
rect 1351 341 1397 379
rect 1351 307 1357 341
rect 1391 307 1397 341
rect 1351 269 1397 307
rect 1351 235 1357 269
rect 1391 235 1397 269
rect 1351 197 1397 235
rect 1351 163 1357 197
rect 1391 163 1397 197
rect 1351 125 1397 163
rect 1351 91 1357 125
rect 1391 91 1397 125
rect 1351 53 1397 91
rect 1351 19 1357 53
rect 1391 19 1397 53
rect 1351 -19 1397 19
rect 1351 -53 1357 -19
rect 1391 -53 1397 -19
rect 1351 -91 1397 -53
rect 1351 -125 1357 -91
rect 1391 -125 1397 -91
rect 1351 -163 1397 -125
rect 1351 -197 1357 -163
rect 1391 -197 1397 -163
rect 1351 -235 1397 -197
rect 1351 -269 1357 -235
rect 1391 -269 1397 -235
rect 1351 -307 1397 -269
rect 1351 -341 1357 -307
rect 1391 -341 1397 -307
rect 1351 -379 1397 -341
rect 1351 -413 1357 -379
rect 1391 -413 1397 -379
rect 1351 -451 1397 -413
rect 1351 -485 1357 -451
rect 1391 -485 1397 -451
rect 1351 -523 1397 -485
rect 1351 -557 1357 -523
rect 1391 -557 1397 -523
rect 1351 -595 1397 -557
rect 1351 -629 1357 -595
rect 1391 -629 1397 -595
rect 1351 -667 1397 -629
rect 1351 -701 1357 -667
rect 1391 -701 1397 -667
rect 1351 -739 1397 -701
rect 1351 -773 1357 -739
rect 1391 -773 1397 -739
rect 1351 -800 1397 -773
rect 1809 773 1855 800
rect 1809 739 1815 773
rect 1849 739 1855 773
rect 1809 701 1855 739
rect 1809 667 1815 701
rect 1849 667 1855 701
rect 1809 629 1855 667
rect 1809 595 1815 629
rect 1849 595 1855 629
rect 1809 557 1855 595
rect 1809 523 1815 557
rect 1849 523 1855 557
rect 1809 485 1855 523
rect 1809 451 1815 485
rect 1849 451 1855 485
rect 1809 413 1855 451
rect 1809 379 1815 413
rect 1849 379 1855 413
rect 1809 341 1855 379
rect 1809 307 1815 341
rect 1849 307 1855 341
rect 1809 269 1855 307
rect 1809 235 1815 269
rect 1849 235 1855 269
rect 1809 197 1855 235
rect 1809 163 1815 197
rect 1849 163 1855 197
rect 1809 125 1855 163
rect 1809 91 1815 125
rect 1849 91 1855 125
rect 1809 53 1855 91
rect 1809 19 1815 53
rect 1849 19 1855 53
rect 1809 -19 1855 19
rect 1809 -53 1815 -19
rect 1849 -53 1855 -19
rect 1809 -91 1855 -53
rect 1809 -125 1815 -91
rect 1849 -125 1855 -91
rect 1809 -163 1855 -125
rect 1809 -197 1815 -163
rect 1849 -197 1855 -163
rect 1809 -235 1855 -197
rect 1809 -269 1815 -235
rect 1849 -269 1855 -235
rect 1809 -307 1855 -269
rect 1809 -341 1815 -307
rect 1849 -341 1855 -307
rect 1809 -379 1855 -341
rect 1809 -413 1815 -379
rect 1849 -413 1855 -379
rect 1809 -451 1855 -413
rect 1809 -485 1815 -451
rect 1849 -485 1855 -451
rect 1809 -523 1855 -485
rect 1809 -557 1815 -523
rect 1849 -557 1855 -523
rect 1809 -595 1855 -557
rect 1809 -629 1815 -595
rect 1849 -629 1855 -595
rect 1809 -667 1855 -629
rect 1809 -701 1815 -667
rect 1849 -701 1855 -667
rect 1809 -739 1855 -701
rect 1809 -773 1815 -739
rect 1849 -773 1855 -739
rect 1809 -800 1855 -773
rect 2267 773 2313 800
rect 2267 739 2273 773
rect 2307 739 2313 773
rect 2267 701 2313 739
rect 2267 667 2273 701
rect 2307 667 2313 701
rect 2267 629 2313 667
rect 2267 595 2273 629
rect 2307 595 2313 629
rect 2267 557 2313 595
rect 2267 523 2273 557
rect 2307 523 2313 557
rect 2267 485 2313 523
rect 2267 451 2273 485
rect 2307 451 2313 485
rect 2267 413 2313 451
rect 2267 379 2273 413
rect 2307 379 2313 413
rect 2267 341 2313 379
rect 2267 307 2273 341
rect 2307 307 2313 341
rect 2267 269 2313 307
rect 2267 235 2273 269
rect 2307 235 2313 269
rect 2267 197 2313 235
rect 2267 163 2273 197
rect 2307 163 2313 197
rect 2267 125 2313 163
rect 2267 91 2273 125
rect 2307 91 2313 125
rect 2267 53 2313 91
rect 2267 19 2273 53
rect 2307 19 2313 53
rect 2267 -19 2313 19
rect 2267 -53 2273 -19
rect 2307 -53 2313 -19
rect 2267 -91 2313 -53
rect 2267 -125 2273 -91
rect 2307 -125 2313 -91
rect 2267 -163 2313 -125
rect 2267 -197 2273 -163
rect 2307 -197 2313 -163
rect 2267 -235 2313 -197
rect 2267 -269 2273 -235
rect 2307 -269 2313 -235
rect 2267 -307 2313 -269
rect 2267 -341 2273 -307
rect 2307 -341 2313 -307
rect 2267 -379 2313 -341
rect 2267 -413 2273 -379
rect 2307 -413 2313 -379
rect 2267 -451 2313 -413
rect 2267 -485 2273 -451
rect 2307 -485 2313 -451
rect 2267 -523 2313 -485
rect 2267 -557 2273 -523
rect 2307 -557 2313 -523
rect 2267 -595 2313 -557
rect 2267 -629 2273 -595
rect 2307 -629 2313 -595
rect 2267 -667 2313 -629
rect 2267 -701 2273 -667
rect 2307 -701 2313 -667
rect 2267 -739 2313 -701
rect 2267 -773 2273 -739
rect 2307 -773 2313 -739
rect 2267 -800 2313 -773
rect 2725 773 2771 800
rect 2725 739 2731 773
rect 2765 739 2771 773
rect 2725 701 2771 739
rect 2725 667 2731 701
rect 2765 667 2771 701
rect 2725 629 2771 667
rect 2725 595 2731 629
rect 2765 595 2771 629
rect 2725 557 2771 595
rect 2725 523 2731 557
rect 2765 523 2771 557
rect 2725 485 2771 523
rect 2725 451 2731 485
rect 2765 451 2771 485
rect 2725 413 2771 451
rect 2725 379 2731 413
rect 2765 379 2771 413
rect 2725 341 2771 379
rect 2725 307 2731 341
rect 2765 307 2771 341
rect 2725 269 2771 307
rect 2725 235 2731 269
rect 2765 235 2771 269
rect 2725 197 2771 235
rect 2725 163 2731 197
rect 2765 163 2771 197
rect 2725 125 2771 163
rect 2725 91 2731 125
rect 2765 91 2771 125
rect 2725 53 2771 91
rect 2725 19 2731 53
rect 2765 19 2771 53
rect 2725 -19 2771 19
rect 2725 -53 2731 -19
rect 2765 -53 2771 -19
rect 2725 -91 2771 -53
rect 2725 -125 2731 -91
rect 2765 -125 2771 -91
rect 2725 -163 2771 -125
rect 2725 -197 2731 -163
rect 2765 -197 2771 -163
rect 2725 -235 2771 -197
rect 2725 -269 2731 -235
rect 2765 -269 2771 -235
rect 2725 -307 2771 -269
rect 2725 -341 2731 -307
rect 2765 -341 2771 -307
rect 2725 -379 2771 -341
rect 2725 -413 2731 -379
rect 2765 -413 2771 -379
rect 2725 -451 2771 -413
rect 2725 -485 2731 -451
rect 2765 -485 2771 -451
rect 2725 -523 2771 -485
rect 2725 -557 2731 -523
rect 2765 -557 2771 -523
rect 2725 -595 2771 -557
rect 2725 -629 2731 -595
rect 2765 -629 2771 -595
rect 2725 -667 2771 -629
rect 2725 -701 2731 -667
rect 2765 -701 2771 -667
rect 2725 -739 2771 -701
rect 2725 -773 2731 -739
rect 2765 -773 2771 -739
rect 2725 -800 2771 -773
rect 3183 773 3229 800
rect 3183 739 3189 773
rect 3223 739 3229 773
rect 3183 701 3229 739
rect 3183 667 3189 701
rect 3223 667 3229 701
rect 3183 629 3229 667
rect 3183 595 3189 629
rect 3223 595 3229 629
rect 3183 557 3229 595
rect 3183 523 3189 557
rect 3223 523 3229 557
rect 3183 485 3229 523
rect 3183 451 3189 485
rect 3223 451 3229 485
rect 3183 413 3229 451
rect 3183 379 3189 413
rect 3223 379 3229 413
rect 3183 341 3229 379
rect 3183 307 3189 341
rect 3223 307 3229 341
rect 3183 269 3229 307
rect 3183 235 3189 269
rect 3223 235 3229 269
rect 3183 197 3229 235
rect 3183 163 3189 197
rect 3223 163 3229 197
rect 3183 125 3229 163
rect 3183 91 3189 125
rect 3223 91 3229 125
rect 3183 53 3229 91
rect 3183 19 3189 53
rect 3223 19 3229 53
rect 3183 -19 3229 19
rect 3183 -53 3189 -19
rect 3223 -53 3229 -19
rect 3183 -91 3229 -53
rect 3183 -125 3189 -91
rect 3223 -125 3229 -91
rect 3183 -163 3229 -125
rect 3183 -197 3189 -163
rect 3223 -197 3229 -163
rect 3183 -235 3229 -197
rect 3183 -269 3189 -235
rect 3223 -269 3229 -235
rect 3183 -307 3229 -269
rect 3183 -341 3189 -307
rect 3223 -341 3229 -307
rect 3183 -379 3229 -341
rect 3183 -413 3189 -379
rect 3223 -413 3229 -379
rect 3183 -451 3229 -413
rect 3183 -485 3189 -451
rect 3223 -485 3229 -451
rect 3183 -523 3229 -485
rect 3183 -557 3189 -523
rect 3223 -557 3229 -523
rect 3183 -595 3229 -557
rect 3183 -629 3189 -595
rect 3223 -629 3229 -595
rect 3183 -667 3229 -629
rect 3183 -701 3189 -667
rect 3223 -701 3229 -667
rect 3183 -739 3229 -701
rect 3183 -773 3189 -739
rect 3223 -773 3229 -739
rect 3183 -800 3229 -773
rect 3641 773 3687 800
rect 3641 739 3647 773
rect 3681 739 3687 773
rect 3641 701 3687 739
rect 3641 667 3647 701
rect 3681 667 3687 701
rect 3641 629 3687 667
rect 3641 595 3647 629
rect 3681 595 3687 629
rect 3641 557 3687 595
rect 3641 523 3647 557
rect 3681 523 3687 557
rect 3641 485 3687 523
rect 3641 451 3647 485
rect 3681 451 3687 485
rect 3641 413 3687 451
rect 3641 379 3647 413
rect 3681 379 3687 413
rect 3641 341 3687 379
rect 3641 307 3647 341
rect 3681 307 3687 341
rect 3641 269 3687 307
rect 3641 235 3647 269
rect 3681 235 3687 269
rect 3641 197 3687 235
rect 3641 163 3647 197
rect 3681 163 3687 197
rect 3641 125 3687 163
rect 3641 91 3647 125
rect 3681 91 3687 125
rect 3641 53 3687 91
rect 3641 19 3647 53
rect 3681 19 3687 53
rect 3641 -19 3687 19
rect 3641 -53 3647 -19
rect 3681 -53 3687 -19
rect 3641 -91 3687 -53
rect 3641 -125 3647 -91
rect 3681 -125 3687 -91
rect 3641 -163 3687 -125
rect 3641 -197 3647 -163
rect 3681 -197 3687 -163
rect 3641 -235 3687 -197
rect 3641 -269 3647 -235
rect 3681 -269 3687 -235
rect 3641 -307 3687 -269
rect 3641 -341 3647 -307
rect 3681 -341 3687 -307
rect 3641 -379 3687 -341
rect 3641 -413 3647 -379
rect 3681 -413 3687 -379
rect 3641 -451 3687 -413
rect 3641 -485 3647 -451
rect 3681 -485 3687 -451
rect 3641 -523 3687 -485
rect 3641 -557 3647 -523
rect 3681 -557 3687 -523
rect 3641 -595 3687 -557
rect 3641 -629 3647 -595
rect 3681 -629 3687 -595
rect 3641 -667 3687 -629
rect 3641 -701 3647 -667
rect 3681 -701 3687 -667
rect 3641 -739 3687 -701
rect 3641 -773 3647 -739
rect 3681 -773 3687 -739
rect 3641 -800 3687 -773
rect 4099 773 4145 800
rect 4099 739 4105 773
rect 4139 739 4145 773
rect 4099 701 4145 739
rect 4099 667 4105 701
rect 4139 667 4145 701
rect 4099 629 4145 667
rect 4099 595 4105 629
rect 4139 595 4145 629
rect 4099 557 4145 595
rect 4099 523 4105 557
rect 4139 523 4145 557
rect 4099 485 4145 523
rect 4099 451 4105 485
rect 4139 451 4145 485
rect 4099 413 4145 451
rect 4099 379 4105 413
rect 4139 379 4145 413
rect 4099 341 4145 379
rect 4099 307 4105 341
rect 4139 307 4145 341
rect 4099 269 4145 307
rect 4099 235 4105 269
rect 4139 235 4145 269
rect 4099 197 4145 235
rect 4099 163 4105 197
rect 4139 163 4145 197
rect 4099 125 4145 163
rect 4099 91 4105 125
rect 4139 91 4145 125
rect 4099 53 4145 91
rect 4099 19 4105 53
rect 4139 19 4145 53
rect 4099 -19 4145 19
rect 4099 -53 4105 -19
rect 4139 -53 4145 -19
rect 4099 -91 4145 -53
rect 4099 -125 4105 -91
rect 4139 -125 4145 -91
rect 4099 -163 4145 -125
rect 4099 -197 4105 -163
rect 4139 -197 4145 -163
rect 4099 -235 4145 -197
rect 4099 -269 4105 -235
rect 4139 -269 4145 -235
rect 4099 -307 4145 -269
rect 4099 -341 4105 -307
rect 4139 -341 4145 -307
rect 4099 -379 4145 -341
rect 4099 -413 4105 -379
rect 4139 -413 4145 -379
rect 4099 -451 4145 -413
rect 4099 -485 4105 -451
rect 4139 -485 4145 -451
rect 4099 -523 4145 -485
rect 4099 -557 4105 -523
rect 4139 -557 4145 -523
rect 4099 -595 4145 -557
rect 4099 -629 4105 -595
rect 4139 -629 4145 -595
rect 4099 -667 4145 -629
rect 4099 -701 4105 -667
rect 4139 -701 4145 -667
rect 4099 -739 4145 -701
rect 4099 -773 4105 -739
rect 4139 -773 4145 -739
rect 4099 -800 4145 -773
rect -3997 -847 -3789 -841
rect -3997 -881 -3982 -847
rect -3948 -881 -3910 -847
rect -3876 -881 -3838 -847
rect -3804 -881 -3789 -847
rect -3997 -887 -3789 -881
rect -3539 -847 -3331 -841
rect -3539 -881 -3524 -847
rect -3490 -881 -3452 -847
rect -3418 -881 -3380 -847
rect -3346 -881 -3331 -847
rect -3539 -887 -3331 -881
rect -3081 -847 -2873 -841
rect -3081 -881 -3066 -847
rect -3032 -881 -2994 -847
rect -2960 -881 -2922 -847
rect -2888 -881 -2873 -847
rect -3081 -887 -2873 -881
rect -2623 -847 -2415 -841
rect -2623 -881 -2608 -847
rect -2574 -881 -2536 -847
rect -2502 -881 -2464 -847
rect -2430 -881 -2415 -847
rect -2623 -887 -2415 -881
rect -2165 -847 -1957 -841
rect -2165 -881 -2150 -847
rect -2116 -881 -2078 -847
rect -2044 -881 -2006 -847
rect -1972 -881 -1957 -847
rect -2165 -887 -1957 -881
rect -1707 -847 -1499 -841
rect -1707 -881 -1692 -847
rect -1658 -881 -1620 -847
rect -1586 -881 -1548 -847
rect -1514 -881 -1499 -847
rect -1707 -887 -1499 -881
rect -1249 -847 -1041 -841
rect -1249 -881 -1234 -847
rect -1200 -881 -1162 -847
rect -1128 -881 -1090 -847
rect -1056 -881 -1041 -847
rect -1249 -887 -1041 -881
rect -791 -847 -583 -841
rect -791 -881 -776 -847
rect -742 -881 -704 -847
rect -670 -881 -632 -847
rect -598 -881 -583 -847
rect -791 -887 -583 -881
rect -333 -847 -125 -841
rect -333 -881 -318 -847
rect -284 -881 -246 -847
rect -212 -881 -174 -847
rect -140 -881 -125 -847
rect -333 -887 -125 -881
rect 125 -847 333 -841
rect 125 -881 140 -847
rect 174 -881 212 -847
rect 246 -881 284 -847
rect 318 -881 333 -847
rect 125 -887 333 -881
rect 583 -847 791 -841
rect 583 -881 598 -847
rect 632 -881 670 -847
rect 704 -881 742 -847
rect 776 -881 791 -847
rect 583 -887 791 -881
rect 1041 -847 1249 -841
rect 1041 -881 1056 -847
rect 1090 -881 1128 -847
rect 1162 -881 1200 -847
rect 1234 -881 1249 -847
rect 1041 -887 1249 -881
rect 1499 -847 1707 -841
rect 1499 -881 1514 -847
rect 1548 -881 1586 -847
rect 1620 -881 1658 -847
rect 1692 -881 1707 -847
rect 1499 -887 1707 -881
rect 1957 -847 2165 -841
rect 1957 -881 1972 -847
rect 2006 -881 2044 -847
rect 2078 -881 2116 -847
rect 2150 -881 2165 -847
rect 1957 -887 2165 -881
rect 2415 -847 2623 -841
rect 2415 -881 2430 -847
rect 2464 -881 2502 -847
rect 2536 -881 2574 -847
rect 2608 -881 2623 -847
rect 2415 -887 2623 -881
rect 2873 -847 3081 -841
rect 2873 -881 2888 -847
rect 2922 -881 2960 -847
rect 2994 -881 3032 -847
rect 3066 -881 3081 -847
rect 2873 -887 3081 -881
rect 3331 -847 3539 -841
rect 3331 -881 3346 -847
rect 3380 -881 3418 -847
rect 3452 -881 3490 -847
rect 3524 -881 3539 -847
rect 3331 -887 3539 -881
rect 3789 -847 3997 -841
rect 3789 -881 3804 -847
rect 3838 -881 3876 -847
rect 3910 -881 3948 -847
rect 3982 -881 3997 -847
rect 3789 -887 3997 -881
<< end >>
