magic
tech sky130A
timestamp 1621481787
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -589 -550 510 550
string parameters w 10.00 l 10.00 val 207.6 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 50
string library sky130
<< end >>
