magic
tech sky130A
magscale 1 2
timestamp 1625985445
<< locali >>
rect 121 14195 155 17901
rect 1409 119 1443 13141
rect 5365 12019 5399 14297
rect 5641 14195 5675 17017
rect 6745 14195 6779 14297
rect 8585 14195 8619 14297
rect 10241 14195 10275 14297
rect 5641 14161 6026 14195
rect 6670 14161 6779 14195
rect 8585 14161 8694 14195
rect 10166 14161 10275 14195
rect 8711 13141 8771 13175
rect 6302 13073 6411 13107
rect 6377 12903 6411 13073
rect 6653 13073 6762 13107
rect 6653 12971 6687 13073
rect 10609 12631 10643 14093
rect 10609 12597 10827 12631
rect 7866 12529 7958 12563
rect 7406 12461 7483 12495
rect 10166 12461 10459 12495
rect 10425 12359 10459 12461
rect 10425 12325 10551 12359
rect 5273 11985 5399 12019
rect 9982 11985 10091 12019
rect 5273 10931 5307 11985
rect 5549 11849 5934 11883
rect 5549 10999 5583 11849
rect 10057 11815 10091 11985
rect 10517 11543 10551 12325
rect 10425 11509 10551 11543
rect 5917 11441 6026 11475
rect 5917 11407 5951 11441
rect 10425 11407 10459 11509
rect 5641 11373 5951 11407
rect 10166 11373 10459 11407
rect 5641 11067 5675 11373
rect 7582 11330 7616 11339
rect 10793 11067 10827 12597
rect 5641 11033 5767 11067
rect 5549 10965 5675 10999
rect 5273 10897 5583 10931
rect 5549 10319 5583 10897
rect 5641 10727 5675 10965
rect 5733 10795 5767 11033
rect 10609 11033 10827 11067
rect 10609 10931 10643 11033
rect 10166 10897 10643 10931
rect 5733 10761 6026 10795
rect 10425 10591 10459 10761
rect 10425 10557 10551 10591
rect 6118 10421 6210 10455
rect 5549 10285 5934 10319
rect 5549 9639 5583 10285
rect 5641 9231 5675 10217
rect 10517 9911 10551 10557
rect 7466 9877 7500 9886
rect 10425 9877 10551 9911
rect 9321 9809 9430 9843
rect 9321 9707 9355 9809
rect 10425 9775 10459 9877
rect 10166 9741 10459 9775
rect 5641 9197 5934 9231
rect 8852 9154 8886 9163
rect 9137 8823 9171 8857
rect 9137 8789 9246 8823
rect 5549 8721 5934 8755
rect 5549 8619 5583 8721
rect 5457 8585 5583 8619
rect 10166 8585 10459 8619
rect 5457 8007 5491 8585
rect 10425 8483 10459 8585
rect 10425 8449 10551 8483
rect 5641 8109 5934 8143
rect 5457 7973 5583 8007
rect 5549 7803 5583 7973
rect 5549 7055 5583 7769
rect 5641 7667 5675 8109
rect 10517 7871 10551 8449
rect 10425 7837 10551 7871
rect 7466 7701 7500 7710
rect 10425 7667 10459 7837
rect 5641 7633 5934 7667
rect 9629 7633 9689 7667
rect 5825 7599 5859 7633
rect 6394 7157 6486 7191
rect 5549 7021 5934 7055
rect 7466 6613 7500 6622
rect 6118 6545 6486 6579
rect 8602 6545 9798 6579
rect 9999 6545 10459 6579
rect 6377 6443 6411 6545
rect 7481 5967 7515 6137
rect 7774 6069 7866 6103
rect 9062 6069 9154 6103
rect 8527 6001 8694 6035
rect 10425 5967 10459 6545
rect 7423 5933 7590 5967
rect 10166 5933 10459 5967
rect 6210 5865 6285 5899
<< viali >>
rect 121 17901 155 17935
rect 5641 17017 5675 17051
rect 121 14161 155 14195
rect 5365 14297 5399 14331
rect 1409 13141 1443 13175
rect 6193 14297 6227 14331
rect 6745 14297 6779 14331
rect 6561 14229 6595 14263
rect 8585 14297 8619 14331
rect 8125 14229 8159 14263
rect 10241 14297 10275 14331
rect 9229 14229 9263 14263
rect 6469 14161 6503 14195
rect 8033 14161 8067 14195
rect 8309 14161 8343 14195
rect 8861 14161 8895 14195
rect 9321 14161 9355 14195
rect 9965 14161 9999 14195
rect 7757 14093 7791 14127
rect 10609 14093 10643 14127
rect 7573 14025 7607 14059
rect 8769 14025 8803 14059
rect 7941 13957 7975 13991
rect 8033 13957 8067 13991
rect 9965 13957 9999 13991
rect 6561 13753 6595 13787
rect 6929 13753 6963 13787
rect 10149 13753 10183 13787
rect 8048 13549 8082 13583
rect 8309 13549 8343 13583
rect 8769 13549 8803 13583
rect 8677 13481 8711 13515
rect 9030 13481 9064 13515
rect 6653 13413 6687 13447
rect 8493 13413 8527 13447
rect 7205 13209 7239 13243
rect 9229 13209 9263 13243
rect 9965 13209 9999 13243
rect 8324 13141 8358 13175
rect 8677 13141 8711 13175
rect 6193 13005 6227 13039
rect 6929 13073 6963 13107
rect 9030 13073 9064 13107
rect 9137 13073 9171 13107
rect 9781 13073 9815 13107
rect 10057 13073 10091 13107
rect 8585 13005 8619 13039
rect 9413 13005 9447 13039
rect 9597 13005 9631 13039
rect 6653 12937 6687 12971
rect 6377 12869 6411 12903
rect 6745 12869 6779 12903
rect 9781 12869 9815 12903
rect 7389 12665 7423 12699
rect 6009 12529 6043 12563
rect 7665 12461 7699 12495
rect 8125 12461 8159 12495
rect 8769 12461 8803 12495
rect 6270 12393 6304 12427
rect 9030 12393 9064 12427
rect 8309 12325 8343 12359
rect 6285 12121 6319 12155
rect 9781 12121 9815 12155
rect 6837 11985 6871 12019
rect 7021 11985 7055 12019
rect 7205 11985 7239 12019
rect 7389 11985 7423 12019
rect 8478 11985 8512 12019
rect 9781 11985 9815 12019
rect 6101 11917 6135 11951
rect 6561 11917 6595 11951
rect 8217 11917 8251 11951
rect 6377 11849 6411 11883
rect 7021 11849 7055 11883
rect 9597 11849 9631 11883
rect 6745 11781 6779 11815
rect 7205 11781 7239 11815
rect 10057 11781 10091 11815
rect 6377 11577 6411 11611
rect 10057 11577 10091 11611
rect 7941 11509 7975 11543
rect 6193 11441 6227 11475
rect 7849 11373 7883 11407
rect 8125 11373 8159 11407
rect 8493 11373 8527 11407
rect 8754 11373 8788 11407
rect 7582 11296 7616 11330
rect 6469 11237 6503 11271
rect 8309 11237 8343 11271
rect 9873 11237 9907 11271
rect 7021 10965 7055 10999
rect 6009 10897 6043 10931
rect 6193 10897 6227 10931
rect 6561 10897 6595 10931
rect 6837 10905 6871 10939
rect 8769 10829 8803 10863
rect 9873 10829 9907 10863
rect 6561 10761 6595 10795
rect 7481 10761 7515 10795
rect 8585 10761 8619 10795
rect 9965 10761 9999 10795
rect 10425 10761 10459 10795
rect 5641 10693 5675 10727
rect 6653 10693 6687 10727
rect 10057 10693 10091 10727
rect 6653 10489 6687 10523
rect 10057 10489 10091 10523
rect 9873 10421 9907 10455
rect 6377 10353 6411 10387
rect 6101 10285 6135 10319
rect 6653 10285 6687 10319
rect 6837 10285 6871 10319
rect 6929 10285 6963 10319
rect 8493 10285 8527 10319
rect 8754 10285 8788 10319
rect 5549 9605 5583 9639
rect 5641 10217 5675 10251
rect 7190 10217 7224 10251
rect 6561 10149 6595 10183
rect 8309 10149 8343 10183
rect 9965 10149 9999 10183
rect 9781 9945 9815 9979
rect 7466 9886 7500 9920
rect 6561 9809 6595 9843
rect 7205 9809 7239 9843
rect 8953 9809 8987 9843
rect 9597 9809 9631 9843
rect 9965 9741 9999 9775
rect 6837 9673 6871 9707
rect 8585 9673 8619 9707
rect 9321 9673 9355 9707
rect 9597 9605 9631 9639
rect 7297 9265 7331 9299
rect 7573 9265 7607 9299
rect 7757 9265 7791 9299
rect 8033 9197 8067 9231
rect 8585 9197 8619 9231
rect 7030 9129 7064 9163
rect 7849 9129 7883 9163
rect 8217 9129 8251 9163
rect 8852 9120 8886 9154
rect 7389 9061 7423 9095
rect 9965 9061 9999 9095
rect 6009 8857 6043 8891
rect 6837 8857 6871 8891
rect 9137 8857 9171 8891
rect 9781 8857 9815 8891
rect 7466 8789 7500 8823
rect 9597 8789 9631 8823
rect 6193 8721 6227 8755
rect 6377 8721 6411 8755
rect 9413 8721 9447 8755
rect 6653 8653 6687 8687
rect 7205 8653 7239 8687
rect 9965 8653 9999 8687
rect 6469 8585 6503 8619
rect 8585 8517 8619 8551
rect 7849 8313 7883 8347
rect 7757 8245 7791 8279
rect 7297 8177 7331 8211
rect 7573 8109 7607 8143
rect 7849 8109 7883 8143
rect 8033 8109 8067 8143
rect 8493 8109 8527 8143
rect 9965 8109 9999 8143
rect 10149 8109 10183 8143
rect 5549 7769 5583 7803
rect 7052 8041 7086 8075
rect 8754 8041 8788 8075
rect 10057 8041 10091 8075
rect 7389 7973 7423 8007
rect 9873 7973 9907 8007
rect 6009 7769 6043 7803
rect 7021 7701 7055 7735
rect 7466 7710 7500 7744
rect 9229 7701 9263 7735
rect 6101 7633 6135 7667
rect 6193 7633 6227 7667
rect 6377 7633 6411 7667
rect 7205 7633 7239 7667
rect 9413 7633 9447 7667
rect 9689 7633 9723 7667
rect 10425 7633 10459 7667
rect 5825 7565 5859 7599
rect 6561 7565 6595 7599
rect 6837 7565 6871 7599
rect 9965 7565 9999 7599
rect 6653 7497 6687 7531
rect 9781 7497 9815 7531
rect 8585 7429 8619 7463
rect 10149 7429 10183 7463
rect 6101 7225 6135 7259
rect 8309 7225 8343 7259
rect 8493 7157 8527 7191
rect 6653 7089 6687 7123
rect 9873 7089 9907 7123
rect 6101 7021 6135 7055
rect 6193 7021 6227 7055
rect 6377 7021 6411 7055
rect 6929 7021 6963 7055
rect 6837 6953 6871 6987
rect 7190 6953 7224 6987
rect 9628 6953 9662 6987
rect 6009 6681 6043 6715
rect 7466 6622 7500 6656
rect 6653 6545 6687 6579
rect 7205 6545 7239 6579
rect 9965 6545 9999 6579
rect 6377 6409 6411 6443
rect 9781 6409 9815 6443
rect 6653 6341 6687 6375
rect 7021 6137 7055 6171
rect 7481 6137 7515 6171
rect 9597 6137 9631 6171
rect 9781 6137 9815 6171
rect 6653 6069 6687 6103
rect 6837 6001 6871 6035
rect 8217 6069 8251 6103
rect 8493 6001 8527 6035
rect 6377 5933 6411 5967
rect 7389 5933 7423 5967
rect 7757 5933 7791 5967
rect 8033 5933 8067 5967
rect 8861 5933 8895 5967
rect 9137 5933 9171 5967
rect 9321 5933 9355 5967
rect 9413 5933 9447 5967
rect 9597 5933 9631 5967
rect 9965 5933 9999 5967
rect 6285 5865 6319 5899
rect 6101 5797 6135 5831
rect 6561 5797 6595 5831
rect 1409 85 1443 119
<< metal1 >>
rect 14 17892 20 17944
rect 72 17932 78 17944
rect 109 17935 167 17941
rect 109 17932 121 17935
rect 72 17904 121 17932
rect 72 17892 78 17904
rect 109 17901 121 17904
rect 155 17901 167 17935
rect 109 17895 167 17901
rect 14 17008 20 17060
rect 72 17048 78 17060
rect 5629 17051 5687 17057
rect 5629 17048 5641 17051
rect 72 17020 5641 17048
rect 72 17008 78 17020
rect 5629 17017 5641 17020
rect 5675 17017 5687 17051
rect 5629 17011 5687 17017
rect 5796 14442 10304 14464
rect 5796 14390 5800 14442
rect 5852 14390 5864 14442
rect 5916 14390 5928 14442
rect 5980 14390 5992 14442
rect 6044 14390 6056 14442
rect 6108 14390 10304 14442
rect 5796 14368 10304 14390
rect 5353 14331 5411 14337
rect 5353 14297 5365 14331
rect 5399 14328 5411 14331
rect 6181 14331 6239 14337
rect 6181 14328 6193 14331
rect 5399 14300 6193 14328
rect 5399 14297 5411 14300
rect 5353 14291 5411 14297
rect 6181 14297 6193 14300
rect 6227 14297 6239 14331
rect 6181 14291 6239 14297
rect 6733 14331 6791 14337
rect 6733 14297 6745 14331
rect 6779 14328 6791 14331
rect 7190 14328 7196 14340
rect 6779 14300 7196 14328
rect 6779 14297 6791 14300
rect 6733 14291 6791 14297
rect 7190 14288 7196 14300
rect 7248 14328 7254 14340
rect 8573 14331 8631 14337
rect 8573 14328 8585 14331
rect 7248 14300 8585 14328
rect 7248 14288 7254 14300
rect 8573 14297 8585 14300
rect 8619 14328 8631 14331
rect 10229 14331 10287 14337
rect 10229 14328 10241 14331
rect 8619 14300 9444 14328
rect 8619 14297 8631 14300
rect 8573 14291 8631 14297
rect 9416 14294 9444 14300
rect 10060 14300 10241 14328
rect 10060 14294 10088 14300
rect 6549 14263 6607 14269
rect 6549 14229 6561 14263
rect 6595 14260 6607 14263
rect 6595 14232 6776 14260
rect 6595 14229 6607 14232
rect 6549 14223 6607 14229
rect 109 14195 167 14201
rect 109 14161 121 14195
rect 155 14192 167 14195
rect 6457 14195 6515 14201
rect 6457 14192 6469 14195
rect 155 14164 5304 14192
rect 155 14161 167 14164
rect 109 14155 167 14161
rect 5276 14124 5304 14164
rect 6288 14164 6469 14192
rect 6288 14124 6316 14164
rect 6457 14161 6469 14164
rect 6503 14161 6515 14195
rect 6457 14155 6515 14161
rect 5276 14096 6316 14124
rect 6748 14124 6776 14232
rect 7926 14220 7932 14272
rect 7984 14260 7990 14272
rect 8113 14263 8171 14269
rect 8113 14260 8125 14263
rect 7984 14232 8125 14260
rect 7984 14220 7990 14232
rect 8113 14229 8125 14232
rect 8159 14260 8171 14263
rect 9217 14263 9275 14269
rect 9416 14266 10088 14294
rect 10229 14297 10241 14300
rect 10275 14297 10287 14331
rect 10229 14291 10287 14297
rect 9217 14260 9229 14263
rect 8159 14232 9229 14260
rect 8159 14229 8171 14232
rect 8113 14223 8171 14229
rect 9217 14229 9229 14232
rect 9263 14229 9275 14263
rect 9217 14223 9275 14229
rect 8021 14195 8079 14201
rect 8021 14192 8033 14195
rect 7392 14164 8033 14192
rect 7392 14124 7420 14164
rect 8021 14161 8033 14164
rect 8067 14161 8079 14195
rect 8297 14195 8355 14201
rect 8297 14192 8309 14195
rect 8021 14155 8079 14161
rect 8220 14164 8309 14192
rect 6748 14096 7420 14124
rect 7742 14084 7748 14136
rect 7800 14124 7806 14136
rect 8110 14124 8116 14136
rect 7800 14096 8116 14124
rect 7800 14084 7806 14096
rect 8110 14084 8116 14096
rect 8168 14124 8174 14136
rect 8220 14124 8248 14164
rect 8297 14161 8309 14164
rect 8343 14161 8355 14195
rect 8297 14155 8355 14161
rect 8849 14195 8907 14201
rect 8849 14161 8861 14195
rect 8895 14192 8907 14195
rect 9309 14195 9367 14201
rect 9309 14192 9321 14195
rect 8895 14164 9321 14192
rect 8895 14161 8907 14164
rect 8849 14155 8907 14161
rect 9309 14161 9321 14164
rect 9355 14192 9367 14195
rect 9953 14195 10011 14201
rect 9953 14192 9965 14195
rect 9355 14164 9965 14192
rect 9355 14161 9367 14164
rect 9309 14155 9367 14161
rect 9953 14161 9965 14164
rect 9999 14192 10011 14195
rect 9999 14164 10088 14192
rect 9999 14161 10011 14164
rect 9953 14155 10011 14161
rect 8168 14096 8248 14124
rect 10060 14124 10088 14164
rect 10597 14127 10655 14133
rect 10597 14124 10609 14127
rect 10060 14096 10609 14124
rect 8168 14084 8174 14096
rect 10597 14093 10609 14096
rect 10643 14093 10655 14127
rect 10597 14087 10655 14093
rect 7561 14059 7619 14065
rect 7561 14025 7573 14059
rect 7607 14056 7619 14059
rect 8757 14059 8815 14065
rect 8757 14056 8769 14059
rect 7607 14028 8769 14056
rect 7607 14025 7619 14028
rect 7561 14019 7619 14025
rect 8757 14025 8769 14028
rect 8803 14056 8815 14059
rect 8846 14056 8852 14068
rect 8803 14028 8852 14056
rect 8803 14025 8815 14028
rect 8757 14019 8815 14025
rect 8846 14016 8852 14028
rect 8904 14016 8910 14068
rect 7650 13948 7656 14000
rect 7708 13988 7714 14000
rect 7929 13991 7987 13997
rect 7929 13988 7941 13991
rect 7708 13960 7941 13988
rect 7708 13948 7714 13960
rect 7929 13957 7941 13960
rect 7975 13957 7987 13991
rect 7929 13951 7987 13957
rect 8018 13948 8024 14000
rect 8076 13988 8082 14000
rect 8076 13960 8137 13988
rect 8076 13948 8082 13960
rect 9674 13948 9680 14000
rect 9732 13988 9738 14000
rect 9953 13991 10011 13997
rect 9953 13988 9965 13991
rect 9732 13960 9965 13988
rect 9732 13948 9738 13960
rect 9953 13957 9965 13960
rect 9999 13957 10011 13991
rect 9953 13951 10011 13957
rect 5796 13898 10304 13920
rect 5796 13846 8182 13898
rect 8234 13846 8246 13898
rect 8298 13846 8310 13898
rect 8362 13846 8374 13898
rect 8426 13846 8438 13898
rect 8490 13846 8502 13898
rect 8554 13846 8566 13898
rect 8618 13846 8630 13898
rect 8682 13846 8694 13898
rect 8746 13846 8758 13898
rect 8810 13846 10304 13898
rect 5796 13824 10304 13846
rect 14 13744 20 13796
rect 72 13784 78 13796
rect 6549 13787 6607 13793
rect 6549 13784 6561 13787
rect 72 13756 5764 13784
rect 72 13744 78 13756
rect 5736 13716 5764 13756
rect 6380 13756 6561 13784
rect 6380 13716 6408 13756
rect 6549 13753 6561 13756
rect 6595 13753 6607 13787
rect 6549 13747 6607 13753
rect 6917 13787 6975 13793
rect 6917 13753 6929 13787
rect 6963 13784 6975 13787
rect 7374 13784 7380 13796
rect 6963 13756 7380 13784
rect 6963 13753 6975 13756
rect 6917 13747 6975 13753
rect 7374 13744 7380 13756
rect 7432 13784 7438 13796
rect 7926 13784 7932 13796
rect 7432 13756 7932 13784
rect 7432 13744 7438 13756
rect 7926 13744 7932 13756
rect 7984 13744 7990 13796
rect 10137 13787 10195 13793
rect 10137 13753 10149 13787
rect 10183 13784 10195 13787
rect 15930 13784 15936 13796
rect 10183 13756 15936 13784
rect 10183 13753 10195 13756
rect 10137 13747 10195 13753
rect 15930 13744 15936 13756
rect 15988 13744 15994 13796
rect 5736 13688 6408 13716
rect 7650 13540 7656 13592
rect 7708 13580 7714 13592
rect 8036 13583 8094 13589
rect 8036 13580 8048 13583
rect 7708 13552 8048 13580
rect 7708 13540 7714 13552
rect 8036 13549 8048 13552
rect 8082 13549 8094 13583
rect 8036 13543 8094 13549
rect 8297 13583 8355 13589
rect 8297 13549 8309 13583
rect 8343 13580 8355 13583
rect 8757 13583 8815 13589
rect 8757 13580 8769 13583
rect 8343 13552 8769 13580
rect 8343 13549 8355 13552
rect 8297 13543 8355 13549
rect 8757 13549 8769 13552
rect 8803 13580 8815 13583
rect 8846 13580 8852 13592
rect 8803 13552 8852 13580
rect 8803 13549 8815 13552
rect 8757 13543 8815 13549
rect 8846 13540 8852 13552
rect 8904 13540 8910 13592
rect 8665 13515 8723 13521
rect 8665 13481 8677 13515
rect 8711 13512 8723 13515
rect 9018 13515 9076 13521
rect 8711 13484 8984 13512
rect 8711 13481 8723 13484
rect 8665 13475 8723 13481
rect 6641 13447 6699 13453
rect 6641 13413 6653 13447
rect 6687 13444 6699 13447
rect 6730 13444 6736 13456
rect 6687 13416 6736 13444
rect 6687 13413 6699 13416
rect 6641 13407 6699 13413
rect 6730 13404 6736 13416
rect 6788 13404 6794 13456
rect 8481 13447 8539 13453
rect 8481 13413 8493 13447
rect 8527 13444 8539 13447
rect 8754 13444 8760 13456
rect 8527 13416 8760 13444
rect 8527 13413 8539 13416
rect 8481 13407 8539 13413
rect 8754 13404 8760 13416
rect 8812 13404 8818 13456
rect 8956 13444 8984 13484
rect 9018 13481 9030 13515
rect 9064 13512 9076 13515
rect 9214 13512 9220 13524
rect 9064 13484 9220 13512
rect 9064 13481 9076 13484
rect 9018 13475 9076 13481
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 9416 13484 10364 13512
rect 9416 13444 9444 13484
rect 8956 13416 9444 13444
rect 5796 13354 10304 13376
rect 5796 13302 5800 13354
rect 5852 13302 5864 13354
rect 5916 13302 5928 13354
rect 5980 13302 5992 13354
rect 6044 13302 6056 13354
rect 6108 13302 10304 13354
rect 5796 13280 10304 13302
rect 7193 13243 7251 13249
rect 7193 13240 7205 13243
rect 1412 13212 5764 13240
rect 1412 13181 1440 13212
rect 1397 13175 1455 13181
rect 1397 13141 1409 13175
rect 1443 13141 1455 13175
rect 5736 13172 5764 13212
rect 6748 13212 7205 13240
rect 6748 13172 6776 13212
rect 7193 13209 7205 13212
rect 7239 13209 7251 13243
rect 9214 13240 9220 13252
rect 9159 13212 9220 13240
rect 7193 13203 7251 13209
rect 9214 13200 9220 13212
rect 9272 13200 9278 13252
rect 9953 13243 10011 13249
rect 9953 13240 9965 13243
rect 9508 13212 9965 13240
rect 5736 13144 6776 13172
rect 8312 13175 8370 13181
rect 1397 13135 1455 13141
rect 8312 13141 8324 13175
rect 8358 13172 8370 13175
rect 8665 13175 8723 13181
rect 8665 13172 8677 13175
rect 8358 13144 8677 13172
rect 8358 13141 8370 13144
rect 8312 13135 8370 13141
rect 8665 13141 8677 13144
rect 8711 13141 8723 13175
rect 8665 13135 8723 13141
rect 14 13064 20 13116
rect 72 13104 78 13116
rect 6917 13107 6975 13113
rect 72 13076 244 13104
rect 72 13064 78 13076
rect 216 13036 244 13076
rect 6917 13073 6929 13107
rect 6963 13104 6975 13107
rect 7006 13104 7012 13116
rect 6963 13076 7012 13104
rect 6963 13073 6975 13076
rect 6917 13067 6975 13073
rect 7006 13064 7012 13076
rect 7064 13064 7070 13116
rect 7742 13064 7748 13116
rect 7800 13104 7806 13116
rect 9018 13107 9076 13113
rect 9018 13104 9030 13107
rect 7800 13076 9030 13104
rect 7800 13064 7806 13076
rect 9018 13073 9030 13076
rect 9064 13073 9076 13107
rect 9018 13067 9076 13073
rect 9125 13107 9183 13113
rect 9125 13073 9137 13107
rect 9171 13104 9183 13107
rect 9508 13104 9536 13212
rect 9953 13209 9965 13212
rect 9999 13240 10011 13243
rect 10336 13240 10364 13484
rect 9999 13212 10364 13240
rect 9999 13209 10011 13212
rect 9953 13203 10011 13209
rect 9171 13076 9536 13104
rect 9171 13073 9183 13076
rect 9125 13067 9183 13073
rect 6181 13039 6239 13045
rect 6181 13036 6193 13039
rect 216 13008 6193 13036
rect 6181 13005 6193 13008
rect 6227 13005 6239 13039
rect 6181 12999 6239 13005
rect 8573 13039 8631 13045
rect 8573 13005 8585 13039
rect 8619 13036 8631 13039
rect 8846 13036 8852 13048
rect 8619 13008 8852 13036
rect 8619 13005 8631 13008
rect 8573 12999 8631 13005
rect 8846 12996 8852 13008
rect 8904 12996 8910 13048
rect 9033 13036 9061 13067
rect 9674 13064 9680 13116
rect 9732 13104 9738 13116
rect 9769 13107 9827 13113
rect 9769 13104 9781 13107
rect 9732 13076 9781 13104
rect 9732 13064 9738 13076
rect 9769 13073 9781 13076
rect 9815 13073 9827 13107
rect 9769 13067 9827 13073
rect 10045 13107 10103 13113
rect 10045 13073 10057 13107
rect 10091 13104 10103 13107
rect 15746 13104 15752 13116
rect 10091 13076 15752 13104
rect 10091 13073 10103 13076
rect 10045 13067 10103 13073
rect 9401 13039 9459 13045
rect 9401 13036 9413 13039
rect 9033 13008 9413 13036
rect 9401 13005 9413 13008
rect 9447 13005 9459 13039
rect 9401 12999 9459 13005
rect 9585 13039 9643 13045
rect 9585 13005 9597 13039
rect 9631 13036 9643 13039
rect 9784 13036 9812 13067
rect 15746 13064 15752 13076
rect 15804 13064 15810 13116
rect 9631 13008 9812 13036
rect 9631 13005 9643 13008
rect 9585 12999 9643 13005
rect 6641 12971 6699 12977
rect 6641 12937 6653 12971
rect 6687 12968 6699 12971
rect 6687 12940 7696 12968
rect 6687 12937 6699 12940
rect 6641 12931 6699 12937
rect 6362 12900 6368 12912
rect 6307 12872 6368 12900
rect 6362 12860 6368 12872
rect 6420 12860 6426 12912
rect 6730 12900 6736 12912
rect 6675 12872 6736 12900
rect 6730 12860 6736 12872
rect 6788 12860 6794 12912
rect 7668 12900 7696 12940
rect 9214 12900 9220 12912
rect 7668 12872 9220 12900
rect 9214 12860 9220 12872
rect 9272 12860 9278 12912
rect 9398 12860 9404 12912
rect 9456 12900 9462 12912
rect 9769 12903 9827 12909
rect 9769 12900 9781 12903
rect 9456 12872 9781 12900
rect 9456 12860 9462 12872
rect 9769 12869 9781 12872
rect 9815 12869 9827 12903
rect 9769 12863 9827 12869
rect 5796 12810 10304 12832
rect 5796 12758 8182 12810
rect 8234 12758 8246 12810
rect 8298 12758 8310 12810
rect 8362 12758 8374 12810
rect 8426 12758 8438 12810
rect 8490 12758 8502 12810
rect 8554 12758 8566 12810
rect 8618 12758 8630 12810
rect 8682 12758 8694 12810
rect 8746 12758 8758 12810
rect 8810 12758 10304 12810
rect 5796 12736 10304 12758
rect 7006 12656 7012 12708
rect 7064 12696 7070 12708
rect 7377 12699 7435 12705
rect 7377 12696 7389 12699
rect 7064 12668 7389 12696
rect 7064 12656 7070 12668
rect 7377 12665 7389 12668
rect 7423 12665 7435 12699
rect 7377 12659 7435 12665
rect 5994 12560 6000 12572
rect 5939 12532 6000 12560
rect 5994 12520 6000 12532
rect 6052 12520 6058 12572
rect 7653 12495 7711 12501
rect 7653 12492 7665 12495
rect 7024 12464 7665 12492
rect 6258 12427 6316 12433
rect 6258 12424 6270 12427
rect 5736 12396 6270 12424
rect 5736 12152 5764 12396
rect 6258 12393 6270 12396
rect 6304 12393 6316 12427
rect 6258 12387 6316 12393
rect 6914 12384 6920 12436
rect 6972 12424 6978 12436
rect 7024 12424 7052 12464
rect 7653 12461 7665 12464
rect 7699 12461 7711 12495
rect 7653 12455 7711 12461
rect 7742 12452 7748 12504
rect 7800 12492 7806 12504
rect 8113 12495 8171 12501
rect 8113 12492 8125 12495
rect 7800 12464 8125 12492
rect 7800 12452 7806 12464
rect 8113 12461 8125 12464
rect 8159 12461 8171 12495
rect 8113 12455 8171 12461
rect 8757 12495 8815 12501
rect 8757 12461 8769 12495
rect 8803 12492 8815 12495
rect 8846 12492 8852 12504
rect 8803 12464 8852 12492
rect 8803 12461 8815 12464
rect 8757 12455 8815 12461
rect 8846 12452 8852 12464
rect 8904 12452 8910 12504
rect 9030 12433 9036 12436
rect 6972 12396 7052 12424
rect 9018 12427 9036 12433
rect 6972 12384 6978 12396
rect 9018 12393 9030 12427
rect 9088 12424 9094 12436
rect 9088 12396 9137 12424
rect 9018 12387 9036 12393
rect 9030 12384 9036 12387
rect 9088 12384 9094 12396
rect 8297 12359 8355 12365
rect 8297 12325 8309 12359
rect 8343 12356 8355 12359
rect 8662 12356 8668 12368
rect 8343 12328 8668 12356
rect 8343 12325 8355 12328
rect 8297 12319 8355 12325
rect 8662 12316 8668 12328
rect 8720 12316 8726 12368
rect 5796 12266 10304 12288
rect 5796 12214 5800 12266
rect 5852 12214 5864 12266
rect 5916 12214 5928 12266
rect 5980 12214 5992 12266
rect 6044 12214 6056 12266
rect 6108 12214 10304 12266
rect 5796 12192 10304 12214
rect 6273 12155 6331 12161
rect 6273 12152 6285 12155
rect 5736 12124 6285 12152
rect 6273 12121 6285 12124
rect 6319 12121 6331 12155
rect 9769 12155 9827 12161
rect 9769 12152 9781 12155
rect 6273 12115 6331 12121
rect 7024 12124 9781 12152
rect 6362 11976 6368 12028
rect 6420 12016 6426 12028
rect 6825 12019 6883 12025
rect 6825 12016 6837 12019
rect 6420 11988 6837 12016
rect 6420 11976 6426 11988
rect 6825 11985 6837 11988
rect 6871 11985 6883 12019
rect 6825 11979 6883 11985
rect 6914 11976 6920 12028
rect 6972 12016 6978 12028
rect 7024 12025 7052 12124
rect 9769 12121 9781 12124
rect 9815 12121 9827 12155
rect 9769 12115 9827 12121
rect 7576 12056 8616 12084
rect 7009 12019 7067 12025
rect 7009 12016 7021 12019
rect 6972 11988 7021 12016
rect 6972 11976 6978 11988
rect 7009 11985 7021 11988
rect 7055 11985 7067 12019
rect 7009 11979 7067 11985
rect 7190 11976 7196 12028
rect 7248 11976 7254 12028
rect 7374 12016 7380 12028
rect 7319 11988 7380 12016
rect 7374 11976 7380 11988
rect 7432 12016 7438 12028
rect 7576 12016 7604 12056
rect 8588 12050 8616 12056
rect 7432 11988 7604 12016
rect 7432 11976 7438 11988
rect 7650 11976 7656 12028
rect 7708 12016 7714 12028
rect 8466 12019 8524 12025
rect 8588 12022 9260 12050
rect 8466 12016 8478 12019
rect 7708 11988 8478 12016
rect 7708 11976 7714 11988
rect 8466 11985 8478 11988
rect 8512 11985 8524 12019
rect 9232 12016 9260 12022
rect 9769 12019 9827 12025
rect 9769 12016 9781 12019
rect 9232 11988 9781 12016
rect 8466 11979 8524 11985
rect 9769 11985 9781 11988
rect 9815 11985 9827 12019
rect 9769 11979 9827 11985
rect 6086 11908 6092 11960
rect 6144 11948 6150 11960
rect 6549 11951 6607 11957
rect 6549 11948 6561 11951
rect 6144 11920 6561 11948
rect 6144 11908 6150 11920
rect 6549 11917 6561 11920
rect 6595 11917 6607 11951
rect 7208 11948 7236 11976
rect 7208 11920 7512 11948
rect 6549 11911 6607 11917
rect 6365 11883 6423 11889
rect 6365 11849 6377 11883
rect 6411 11880 6423 11883
rect 7009 11883 7067 11889
rect 7009 11880 7021 11883
rect 6411 11852 7021 11880
rect 6411 11849 6423 11852
rect 6365 11843 6423 11849
rect 7009 11849 7021 11852
rect 7055 11849 7067 11883
rect 7484 11880 7512 11920
rect 7558 11908 7564 11960
rect 7616 11948 7622 11960
rect 8205 11951 8263 11957
rect 8205 11948 8217 11951
rect 7616 11920 8217 11948
rect 7616 11908 7622 11920
rect 8205 11917 8217 11920
rect 8251 11917 8263 11951
rect 8205 11911 8263 11917
rect 7484 11852 8064 11880
rect 7009 11843 7067 11849
rect 6733 11815 6791 11821
rect 6733 11781 6745 11815
rect 6779 11812 6791 11815
rect 6822 11812 6828 11824
rect 6779 11784 6828 11812
rect 6779 11781 6791 11784
rect 6733 11775 6791 11781
rect 6822 11772 6828 11784
rect 6880 11772 6886 11824
rect 7193 11815 7251 11821
rect 7193 11781 7205 11815
rect 7239 11812 7251 11815
rect 7834 11812 7840 11824
rect 7239 11784 7840 11812
rect 7239 11781 7251 11784
rect 7193 11775 7251 11781
rect 7834 11772 7840 11784
rect 7892 11772 7898 11824
rect 8036 11812 8064 11852
rect 9214 11840 9220 11892
rect 9272 11880 9278 11892
rect 9585 11883 9643 11889
rect 9585 11880 9597 11883
rect 9272 11852 9597 11880
rect 9272 11840 9278 11852
rect 9585 11849 9597 11852
rect 9631 11849 9643 11883
rect 9585 11843 9643 11849
rect 10045 11815 10103 11821
rect 10045 11812 10057 11815
rect 8036 11784 10057 11812
rect 10045 11781 10057 11784
rect 10091 11812 10103 11815
rect 10091 11784 10364 11812
rect 10091 11781 10103 11784
rect 10045 11775 10103 11781
rect 5796 11722 10304 11744
rect 5796 11670 8182 11722
rect 8234 11670 8246 11722
rect 8298 11670 8310 11722
rect 8362 11670 8374 11722
rect 8426 11670 8438 11722
rect 8490 11670 8502 11722
rect 8554 11670 8566 11722
rect 8618 11670 8630 11722
rect 8682 11670 8694 11722
rect 8746 11670 8758 11722
rect 8810 11670 10304 11722
rect 5796 11648 10304 11670
rect 6365 11611 6423 11617
rect 6365 11577 6377 11611
rect 6411 11608 6423 11611
rect 7650 11608 7656 11620
rect 6411 11580 7656 11608
rect 6411 11577 6423 11580
rect 6365 11571 6423 11577
rect 7650 11568 7656 11580
rect 7708 11568 7714 11620
rect 10045 11611 10103 11617
rect 10045 11577 10057 11611
rect 10091 11608 10103 11611
rect 10336 11608 10364 11784
rect 10091 11580 10364 11608
rect 10091 11577 10103 11580
rect 10045 11571 10103 11577
rect 7834 11500 7840 11552
rect 7892 11540 7898 11552
rect 7929 11543 7987 11549
rect 7929 11540 7941 11543
rect 7892 11512 7941 11540
rect 7892 11500 7898 11512
rect 7929 11509 7941 11512
rect 7975 11509 7987 11543
rect 7929 11503 7987 11509
rect 6086 11432 6092 11484
rect 6144 11472 6150 11484
rect 6181 11475 6239 11481
rect 6181 11472 6193 11475
rect 6144 11444 6193 11472
rect 6144 11432 6150 11444
rect 6181 11441 6193 11444
rect 6227 11441 6239 11475
rect 6181 11435 6239 11441
rect 7558 11364 7564 11416
rect 7616 11404 7622 11416
rect 7837 11407 7895 11413
rect 7837 11404 7849 11407
rect 7616 11376 7849 11404
rect 7616 11364 7622 11376
rect 7837 11373 7849 11376
rect 7883 11373 7895 11407
rect 8113 11407 8171 11413
rect 8113 11404 8125 11407
rect 7837 11367 7895 11373
rect 7944 11376 8125 11404
rect 6822 11296 6828 11348
rect 6880 11336 6886 11348
rect 6880 11330 7628 11336
rect 6880 11308 7582 11330
rect 6880 11296 6886 11308
rect 7570 11296 7582 11308
rect 7616 11296 7628 11330
rect 7742 11296 7748 11348
rect 7800 11336 7806 11348
rect 7944 11336 7972 11376
rect 8113 11373 8125 11376
rect 8159 11373 8171 11407
rect 8478 11404 8484 11416
rect 8423 11376 8484 11404
rect 8113 11367 8171 11373
rect 8478 11364 8484 11376
rect 8536 11364 8542 11416
rect 8754 11413 8760 11416
rect 8742 11407 8760 11413
rect 8742 11404 8754 11407
rect 8699 11376 8754 11404
rect 8742 11373 8754 11376
rect 8742 11367 8760 11373
rect 8754 11364 8760 11367
rect 8812 11364 8818 11416
rect 7800 11308 7972 11336
rect 7800 11296 7806 11308
rect 7570 11290 7628 11296
rect 6362 11228 6368 11280
rect 6420 11268 6426 11280
rect 6457 11271 6515 11277
rect 6457 11268 6469 11271
rect 6420 11240 6469 11268
rect 6420 11228 6426 11240
rect 6457 11237 6469 11240
rect 6503 11237 6515 11271
rect 6457 11231 6515 11237
rect 8297 11271 8355 11277
rect 8297 11237 8309 11271
rect 8343 11268 8355 11271
rect 8846 11268 8852 11280
rect 8343 11240 8852 11268
rect 8343 11237 8355 11240
rect 8297 11231 8355 11237
rect 8846 11228 8852 11240
rect 8904 11228 8910 11280
rect 9582 11228 9588 11280
rect 9640 11268 9646 11280
rect 9861 11271 9919 11277
rect 9861 11268 9873 11271
rect 9640 11240 9873 11268
rect 9640 11228 9646 11240
rect 9861 11237 9873 11240
rect 9907 11237 9919 11271
rect 9861 11231 9919 11237
rect 5796 11178 10304 11200
rect 5796 11126 5800 11178
rect 5852 11126 5864 11178
rect 5916 11126 5928 11178
rect 5980 11126 5992 11178
rect 6044 11126 6056 11178
rect 6108 11126 10304 11178
rect 5796 11104 10304 11126
rect 6914 11064 6920 11076
rect 6012 11036 6920 11064
rect 6012 10940 6040 11036
rect 6840 10945 6868 11036
rect 6914 11024 6920 11036
rect 6972 11024 6978 11076
rect 7009 10999 7067 11005
rect 7009 10965 7021 10999
rect 7055 10996 7067 10999
rect 7098 10996 7104 11008
rect 7055 10968 7104 10996
rect 7055 10965 7067 10968
rect 7009 10959 7067 10965
rect 7098 10956 7104 10968
rect 7156 10956 7162 11008
rect 5994 10928 6000 10940
rect 5939 10900 6000 10928
rect 5994 10888 6000 10900
rect 6052 10888 6058 10940
rect 6178 10928 6184 10940
rect 6123 10900 6184 10928
rect 6178 10888 6184 10900
rect 6236 10888 6242 10940
rect 6546 10888 6552 10940
rect 6604 10888 6610 10940
rect 6825 10939 6883 10945
rect 6825 10905 6837 10939
rect 6871 10905 6883 10939
rect 6825 10899 6883 10905
rect 7650 10888 7656 10940
rect 7708 10888 7714 10940
rect 8757 10863 8815 10869
rect 8757 10829 8769 10863
rect 8803 10860 8815 10863
rect 8938 10860 8944 10872
rect 8803 10832 8944 10860
rect 8803 10829 8815 10832
rect 8757 10823 8815 10829
rect 8938 10820 8944 10832
rect 8996 10820 9002 10872
rect 9398 10820 9404 10872
rect 9456 10860 9462 10872
rect 9861 10863 9919 10869
rect 9861 10860 9873 10863
rect 9456 10832 9873 10860
rect 9456 10820 9462 10832
rect 9861 10829 9873 10832
rect 9907 10829 9919 10863
rect 9861 10823 9919 10829
rect 6546 10792 6552 10804
rect 5828 10764 6316 10792
rect 6491 10764 6552 10792
rect 5629 10727 5687 10733
rect 5629 10693 5641 10727
rect 5675 10724 5687 10727
rect 5828 10724 5856 10764
rect 5675 10696 5856 10724
rect 6288 10724 6316 10764
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 7466 10792 7472 10804
rect 7411 10764 7472 10792
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 8018 10752 8024 10804
rect 8076 10792 8082 10804
rect 8573 10795 8631 10801
rect 8573 10792 8585 10795
rect 8076 10764 8585 10792
rect 8076 10752 8082 10764
rect 8573 10761 8585 10764
rect 8619 10761 8631 10795
rect 8573 10755 8631 10761
rect 9953 10795 10011 10801
rect 9953 10761 9965 10795
rect 9999 10792 10011 10795
rect 10413 10795 10471 10801
rect 10413 10792 10425 10795
rect 9999 10764 10425 10792
rect 9999 10761 10011 10764
rect 9953 10755 10011 10761
rect 10413 10761 10425 10764
rect 10459 10761 10471 10795
rect 10413 10755 10471 10761
rect 6641 10727 6699 10733
rect 6641 10724 6653 10727
rect 6288 10696 6653 10724
rect 5675 10693 5687 10696
rect 5629 10687 5687 10693
rect 6641 10693 6653 10696
rect 6687 10693 6699 10727
rect 6641 10687 6699 10693
rect 10045 10727 10103 10733
rect 10045 10693 10057 10727
rect 10091 10724 10103 10727
rect 10091 10696 10364 10724
rect 10091 10693 10103 10696
rect 10045 10687 10103 10693
rect 5796 10634 10304 10656
rect 5796 10582 8182 10634
rect 8234 10582 8246 10634
rect 8298 10582 8310 10634
rect 8362 10582 8374 10634
rect 8426 10582 8438 10634
rect 8490 10582 8502 10634
rect 8554 10582 8566 10634
rect 8618 10582 8630 10634
rect 8682 10582 8694 10634
rect 8746 10582 8758 10634
rect 8810 10582 10304 10634
rect 5796 10560 10304 10582
rect 6270 10480 6276 10532
rect 6328 10520 6334 10532
rect 6641 10523 6699 10529
rect 6641 10520 6653 10523
rect 6328 10492 6653 10520
rect 6328 10480 6334 10492
rect 6641 10489 6653 10492
rect 6687 10489 6699 10523
rect 7098 10520 7104 10532
rect 6641 10483 6699 10489
rect 6840 10492 7104 10520
rect 5718 10344 5724 10396
rect 5776 10384 5782 10396
rect 6365 10387 6423 10393
rect 6365 10384 6377 10387
rect 5776 10356 6377 10384
rect 5776 10344 5782 10356
rect 6365 10353 6377 10356
rect 6411 10384 6423 10387
rect 6730 10384 6736 10396
rect 6411 10356 6736 10384
rect 6411 10353 6423 10356
rect 6365 10347 6423 10353
rect 6730 10344 6736 10356
rect 6788 10344 6794 10396
rect 5994 10276 6000 10328
rect 6052 10316 6058 10328
rect 6089 10319 6147 10325
rect 6089 10316 6101 10319
rect 6052 10288 6101 10316
rect 6052 10276 6058 10288
rect 6089 10285 6101 10288
rect 6135 10316 6147 10319
rect 6178 10316 6184 10328
rect 6135 10288 6184 10316
rect 6135 10285 6147 10288
rect 6089 10279 6147 10285
rect 6178 10276 6184 10288
rect 6236 10276 6242 10328
rect 6454 10276 6460 10328
rect 6512 10316 6518 10328
rect 6840 10325 6868 10492
rect 7098 10480 7104 10492
rect 7156 10480 7162 10532
rect 10045 10523 10103 10529
rect 10045 10489 10057 10523
rect 10091 10520 10103 10523
rect 10336 10520 10364 10696
rect 10091 10492 10364 10520
rect 10091 10489 10103 10492
rect 10045 10483 10103 10489
rect 9861 10455 9919 10461
rect 9861 10421 9873 10455
rect 9907 10452 9919 10455
rect 10226 10452 10232 10464
rect 9907 10424 10232 10452
rect 9907 10421 9919 10424
rect 9861 10415 9919 10421
rect 10226 10412 10232 10424
rect 10284 10412 10290 10464
rect 6641 10319 6699 10325
rect 6641 10316 6653 10319
rect 6512 10288 6653 10316
rect 6512 10276 6518 10288
rect 6641 10285 6653 10288
rect 6687 10285 6699 10319
rect 6825 10319 6883 10325
rect 6825 10316 6837 10319
rect 6641 10279 6699 10285
rect 6748 10288 6837 10316
rect 5629 10251 5687 10257
rect 5629 10217 5641 10251
rect 5675 10248 5687 10251
rect 6748 10248 6776 10288
rect 6825 10285 6837 10288
rect 6871 10285 6883 10319
rect 6825 10279 6883 10285
rect 6917 10319 6975 10325
rect 6917 10285 6929 10319
rect 6963 10316 6975 10319
rect 7466 10316 7472 10328
rect 6963 10288 7472 10316
rect 6963 10285 6975 10288
rect 6917 10279 6975 10285
rect 7466 10276 7472 10288
rect 7524 10276 7530 10328
rect 8478 10316 8484 10328
rect 8423 10288 8484 10316
rect 8478 10276 8484 10288
rect 8536 10276 8542 10328
rect 8754 10325 8760 10328
rect 8742 10319 8760 10325
rect 8742 10316 8754 10319
rect 8699 10288 8754 10316
rect 8742 10285 8754 10288
rect 8742 10279 8760 10285
rect 8754 10276 8760 10279
rect 8812 10276 8818 10328
rect 7190 10257 7196 10260
rect 7178 10251 7196 10257
rect 7178 10248 7190 10251
rect 5675 10220 6776 10248
rect 7135 10220 7190 10248
rect 5675 10217 5687 10220
rect 5629 10211 5687 10217
rect 7178 10217 7190 10220
rect 7178 10211 7196 10217
rect 7190 10208 7196 10211
rect 7248 10208 7254 10260
rect 9766 10248 9772 10260
rect 8956 10220 9772 10248
rect 6549 10183 6607 10189
rect 6549 10149 6561 10183
rect 6595 10180 6607 10183
rect 7006 10180 7012 10192
rect 6595 10152 7012 10180
rect 6595 10149 6607 10152
rect 6549 10143 6607 10149
rect 7006 10140 7012 10152
rect 7064 10140 7070 10192
rect 8297 10183 8355 10189
rect 8297 10149 8309 10183
rect 8343 10180 8355 10183
rect 8956 10180 8984 10220
rect 9766 10208 9772 10220
rect 9824 10208 9830 10260
rect 8343 10152 8984 10180
rect 8343 10149 8355 10152
rect 8297 10143 8355 10149
rect 9582 10140 9588 10192
rect 9640 10180 9646 10192
rect 9953 10183 10011 10189
rect 9953 10180 9965 10183
rect 9640 10152 9965 10180
rect 9640 10140 9646 10152
rect 9953 10149 9965 10152
rect 9999 10180 10011 10183
rect 9999 10152 10364 10180
rect 9999 10149 10011 10152
rect 9953 10143 10011 10149
rect 5796 10090 10304 10112
rect 5796 10038 5800 10090
rect 5852 10038 5864 10090
rect 5916 10038 5928 10090
rect 5980 10038 5992 10090
rect 6044 10038 6056 10090
rect 6108 10038 10304 10090
rect 5796 10016 10304 10038
rect 9122 9936 9128 9988
rect 9180 9976 9186 9988
rect 9769 9979 9827 9985
rect 9769 9976 9781 9979
rect 9180 9948 9781 9976
rect 9180 9936 9186 9948
rect 9769 9945 9781 9948
rect 9815 9945 9827 9979
rect 9769 9939 9827 9945
rect 7454 9920 7512 9926
rect 7006 9868 7012 9920
rect 7064 9908 7070 9920
rect 7454 9908 7466 9920
rect 7064 9886 7466 9908
rect 7500 9886 7512 9920
rect 7064 9880 7512 9886
rect 7064 9868 7070 9880
rect 7742 9868 7748 9920
rect 7800 9908 7806 9920
rect 7800 9880 9076 9908
rect 7800 9868 7806 9880
rect 6546 9840 6552 9852
rect 6491 9812 6552 9840
rect 6546 9800 6552 9812
rect 6604 9800 6610 9852
rect 7193 9843 7251 9849
rect 7193 9809 7205 9843
rect 7239 9840 7251 9843
rect 7466 9840 7472 9852
rect 7239 9812 7472 9840
rect 7239 9809 7251 9812
rect 7193 9803 7251 9809
rect 7466 9800 7472 9812
rect 7524 9800 7530 9852
rect 8938 9840 8944 9852
rect 8883 9812 8944 9840
rect 8938 9800 8944 9812
rect 8996 9800 9002 9852
rect 9048 9772 9076 9880
rect 10336 9874 10364 10152
rect 9585 9843 9643 9849
rect 9585 9809 9597 9843
rect 9631 9840 9643 9843
rect 9784 9846 10364 9874
rect 9784 9840 9812 9846
rect 9631 9812 9812 9840
rect 9631 9809 9643 9812
rect 9585 9803 9643 9809
rect 9953 9775 10011 9781
rect 9953 9772 9965 9775
rect 9048 9744 9965 9772
rect 9953 9741 9965 9744
rect 9999 9741 10011 9775
rect 9953 9735 10011 9741
rect 6822 9704 6828 9716
rect 5736 9676 6316 9704
rect 6767 9676 6828 9704
rect 5537 9639 5595 9645
rect 5537 9605 5549 9639
rect 5583 9636 5595 9639
rect 5736 9636 5764 9676
rect 5583 9608 5764 9636
rect 6288 9636 6316 9676
rect 6822 9664 6828 9676
rect 6880 9664 6886 9716
rect 8573 9707 8631 9713
rect 8573 9673 8585 9707
rect 8619 9704 8631 9707
rect 9309 9707 9367 9713
rect 9309 9704 9321 9707
rect 8619 9676 9321 9704
rect 8619 9673 8631 9676
rect 8573 9667 8631 9673
rect 9309 9673 9321 9676
rect 9355 9673 9367 9707
rect 9968 9704 9996 9735
rect 10502 9704 10508 9716
rect 9968 9676 10508 9704
rect 9309 9667 9367 9673
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 9585 9639 9643 9645
rect 9585 9636 9597 9639
rect 6288 9608 9597 9636
rect 5583 9605 5595 9608
rect 5537 9599 5595 9605
rect 9585 9605 9597 9608
rect 9631 9605 9643 9639
rect 9585 9599 9643 9605
rect 5796 9546 10304 9568
rect 5796 9494 8182 9546
rect 8234 9494 8246 9546
rect 8298 9494 8310 9546
rect 8362 9494 8374 9546
rect 8426 9494 8438 9546
rect 8490 9494 8502 9546
rect 8554 9494 8566 9546
rect 8618 9494 8630 9546
rect 8682 9494 8694 9546
rect 8746 9494 8758 9546
rect 8810 9494 10304 9546
rect 5796 9472 10304 9494
rect 7285 9299 7343 9305
rect 7285 9265 7297 9299
rect 7331 9296 7343 9299
rect 7374 9296 7380 9308
rect 7331 9268 7380 9296
rect 7331 9265 7343 9268
rect 7285 9259 7343 9265
rect 7374 9256 7380 9268
rect 7432 9256 7438 9308
rect 7558 9296 7564 9308
rect 7503 9268 7564 9296
rect 7558 9256 7564 9268
rect 7616 9256 7622 9308
rect 7745 9299 7803 9305
rect 7745 9265 7757 9299
rect 7791 9296 7803 9299
rect 8478 9296 8484 9308
rect 7791 9268 8484 9296
rect 7791 9265 7803 9268
rect 7745 9259 7803 9265
rect 8478 9256 8484 9268
rect 8536 9256 8542 9308
rect 8018 9228 8024 9240
rect 7963 9200 8024 9228
rect 8018 9188 8024 9200
rect 8076 9188 8082 9240
rect 8573 9231 8631 9237
rect 8573 9197 8585 9231
rect 8619 9228 8631 9231
rect 8846 9228 8852 9240
rect 8619 9200 8852 9228
rect 8619 9197 8631 9200
rect 8573 9191 8631 9197
rect 8846 9188 8852 9200
rect 8904 9188 8910 9240
rect 6822 9120 6828 9172
rect 6880 9160 6886 9172
rect 7018 9163 7076 9169
rect 7018 9160 7030 9163
rect 6880 9132 7030 9160
rect 6880 9120 6886 9132
rect 7018 9129 7030 9132
rect 7064 9129 7076 9163
rect 7018 9123 7076 9129
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 7837 9163 7895 9169
rect 7837 9160 7849 9163
rect 7800 9132 7849 9160
rect 7800 9120 7806 9132
rect 7837 9129 7849 9132
rect 7883 9129 7895 9163
rect 7837 9123 7895 9129
rect 8110 9120 8116 9172
rect 8168 9160 8174 9172
rect 8205 9163 8263 9169
rect 8205 9160 8217 9163
rect 8168 9132 8217 9160
rect 8168 9120 8174 9132
rect 8205 9129 8217 9132
rect 8251 9129 8263 9163
rect 9214 9160 9220 9172
rect 8205 9123 8263 9129
rect 8840 9154 9220 9160
rect 8840 9120 8852 9154
rect 8886 9132 9220 9154
rect 8886 9120 8898 9132
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 8840 9114 8898 9120
rect 7377 9095 7435 9101
rect 7377 9061 7389 9095
rect 7423 9092 7435 9095
rect 7558 9092 7564 9104
rect 7423 9064 7564 9092
rect 7423 9061 7435 9064
rect 7377 9055 7435 9061
rect 7558 9052 7564 9064
rect 7616 9052 7622 9104
rect 9950 9092 9956 9104
rect 9895 9064 9956 9092
rect 9950 9052 9956 9064
rect 10008 9052 10014 9104
rect 14 8984 20 9036
rect 72 8984 78 9036
rect 5796 9002 10304 9024
rect 32 8888 60 8984
rect 5796 8950 5800 9002
rect 5852 8950 5864 9002
rect 5916 8950 5928 9002
rect 5980 8950 5992 9002
rect 6044 8950 6056 9002
rect 6108 8950 10304 9002
rect 5796 8928 10304 8950
rect 5997 8891 6055 8897
rect 5997 8888 6009 8891
rect 32 8860 6009 8888
rect 5997 8857 6009 8860
rect 6043 8857 6055 8891
rect 6822 8888 6828 8900
rect 6767 8860 6828 8888
rect 5997 8851 6055 8857
rect 6822 8848 6828 8860
rect 6880 8848 6886 8900
rect 8478 8848 8484 8900
rect 8536 8888 8542 8900
rect 9125 8891 9183 8897
rect 9125 8888 9137 8891
rect 8536 8860 9137 8888
rect 8536 8848 8542 8860
rect 9125 8857 9137 8860
rect 9171 8857 9183 8891
rect 9125 8851 9183 8857
rect 9214 8848 9220 8900
rect 9272 8888 9278 8900
rect 9769 8891 9827 8897
rect 9769 8888 9781 8891
rect 9272 8860 9781 8888
rect 9272 8848 9278 8860
rect 9769 8857 9781 8860
rect 9815 8857 9827 8891
rect 9769 8851 9827 8857
rect 7454 8823 7512 8829
rect 7454 8789 7466 8823
rect 7500 8820 7512 8823
rect 7558 8820 7564 8832
rect 7500 8792 7564 8820
rect 7500 8789 7512 8792
rect 7454 8783 7512 8789
rect 7558 8780 7564 8792
rect 7616 8780 7622 8832
rect 9585 8823 9643 8829
rect 9585 8789 9597 8823
rect 9631 8820 9643 8823
rect 10226 8820 10232 8832
rect 9631 8792 10232 8820
rect 9631 8789 9643 8792
rect 9585 8783 9643 8789
rect 10226 8780 10232 8792
rect 10284 8780 10290 8832
rect 14 8712 20 8764
rect 72 8752 78 8764
rect 6181 8755 6239 8761
rect 6181 8752 6193 8755
rect 72 8724 244 8752
rect 72 8712 78 8724
rect 216 8684 244 8724
rect 6012 8724 6193 8752
rect 6012 8684 6040 8724
rect 6181 8721 6193 8724
rect 6227 8721 6239 8755
rect 6181 8715 6239 8721
rect 6365 8755 6423 8761
rect 6365 8721 6377 8755
rect 6411 8752 6423 8755
rect 6546 8752 6552 8764
rect 6411 8724 6552 8752
rect 6411 8721 6423 8724
rect 6365 8715 6423 8721
rect 6546 8712 6552 8724
rect 6604 8712 6610 8764
rect 8662 8712 8668 8764
rect 8720 8752 8726 8764
rect 9401 8755 9459 8761
rect 9401 8752 9413 8755
rect 8720 8724 9413 8752
rect 8720 8712 8726 8724
rect 9401 8721 9413 8724
rect 9447 8721 9459 8755
rect 9401 8715 9459 8721
rect 216 8656 6040 8684
rect 6641 8687 6699 8693
rect 6641 8653 6653 8687
rect 6687 8684 6699 8687
rect 6730 8684 6736 8696
rect 6687 8656 6736 8684
rect 6687 8653 6699 8656
rect 6641 8647 6699 8653
rect 6730 8644 6736 8656
rect 6788 8644 6794 8696
rect 6914 8644 6920 8696
rect 6972 8684 6978 8696
rect 7193 8687 7251 8693
rect 7193 8684 7205 8687
rect 6972 8656 7205 8684
rect 6972 8644 6978 8656
rect 7193 8653 7205 8656
rect 7239 8653 7251 8687
rect 7193 8647 7251 8653
rect 9953 8687 10011 8693
rect 9953 8653 9965 8687
rect 9999 8684 10011 8687
rect 10502 8684 10508 8696
rect 9999 8656 10508 8684
rect 9999 8653 10011 8656
rect 9953 8647 10011 8653
rect 10502 8644 10508 8656
rect 10560 8644 10566 8696
rect 6454 8616 6460 8628
rect 6399 8588 6460 8616
rect 6454 8576 6460 8588
rect 6512 8576 6518 8628
rect 8573 8551 8631 8557
rect 8573 8517 8585 8551
rect 8619 8548 8631 8551
rect 9030 8548 9036 8560
rect 8619 8520 9036 8548
rect 8619 8517 8631 8520
rect 8573 8511 8631 8517
rect 9030 8508 9036 8520
rect 9088 8508 9094 8560
rect 5796 8458 10304 8480
rect 5796 8406 8182 8458
rect 8234 8406 8246 8458
rect 8298 8406 8310 8458
rect 8362 8406 8374 8458
rect 8426 8406 8438 8458
rect 8490 8406 8502 8458
rect 8554 8406 8566 8458
rect 8618 8406 8630 8458
rect 8682 8406 8694 8458
rect 8746 8406 8758 8458
rect 8810 8406 10304 8458
rect 5796 8384 10304 8406
rect 6546 8304 6552 8356
rect 6604 8344 6610 8356
rect 7837 8347 7895 8353
rect 7837 8344 7849 8347
rect 6604 8316 7849 8344
rect 6604 8304 6610 8316
rect 7837 8313 7849 8316
rect 7883 8313 7895 8347
rect 7837 8307 7895 8313
rect 7742 8276 7748 8288
rect 7687 8248 7748 8276
rect 7742 8236 7748 8248
rect 7800 8236 7806 8288
rect 7285 8211 7343 8217
rect 7285 8177 7297 8211
rect 7331 8208 7343 8211
rect 7374 8208 7380 8220
rect 7331 8180 7380 8208
rect 7331 8177 7343 8180
rect 7285 8171 7343 8177
rect 7374 8168 7380 8180
rect 7432 8168 7438 8220
rect 7561 8143 7619 8149
rect 7561 8140 7573 8143
rect 7392 8112 7573 8140
rect 7040 8075 7098 8081
rect 7040 8041 7052 8075
rect 7086 8041 7098 8075
rect 7040 8035 7098 8041
rect 7055 8004 7083 8035
rect 7190 8032 7196 8084
rect 7248 8072 7254 8084
rect 7392 8072 7420 8112
rect 7561 8109 7573 8112
rect 7607 8109 7619 8143
rect 7561 8103 7619 8109
rect 7837 8143 7895 8149
rect 7837 8109 7849 8143
rect 7883 8140 7895 8143
rect 7926 8140 7932 8152
rect 7883 8112 7932 8140
rect 7883 8109 7895 8112
rect 7837 8103 7895 8109
rect 7926 8100 7932 8112
rect 7984 8100 7990 8152
rect 8018 8100 8024 8152
rect 8076 8140 8082 8152
rect 8478 8140 8484 8152
rect 8076 8112 8137 8140
rect 8423 8112 8484 8140
rect 8076 8100 8082 8112
rect 8478 8100 8484 8112
rect 8536 8100 8542 8152
rect 9766 8100 9772 8152
rect 9824 8140 9830 8152
rect 9953 8143 10011 8149
rect 9953 8140 9965 8143
rect 9824 8112 9965 8140
rect 9824 8100 9830 8112
rect 9953 8109 9965 8112
rect 9999 8109 10011 8143
rect 9953 8103 10011 8109
rect 10137 8143 10195 8149
rect 10137 8109 10149 8143
rect 10183 8140 10195 8143
rect 10226 8140 10232 8152
rect 10183 8112 10232 8140
rect 10183 8109 10195 8112
rect 10137 8103 10195 8109
rect 10226 8100 10232 8112
rect 10284 8100 10290 8152
rect 7248 8044 7420 8072
rect 8742 8075 8800 8081
rect 7248 8032 7254 8044
rect 8742 8041 8754 8075
rect 8788 8072 8800 8075
rect 8846 8072 8852 8084
rect 8788 8044 8852 8072
rect 8788 8041 8800 8044
rect 8742 8035 8800 8041
rect 8846 8032 8852 8044
rect 8904 8032 8910 8084
rect 10045 8075 10103 8081
rect 10045 8041 10057 8075
rect 10091 8072 10103 8075
rect 10318 8072 10324 8084
rect 10091 8044 10324 8072
rect 10091 8041 10103 8044
rect 10045 8035 10103 8041
rect 10318 8032 10324 8044
rect 10376 8032 10382 8084
rect 7377 8007 7435 8013
rect 7377 8004 7389 8007
rect 7055 7976 7389 8004
rect 7377 7973 7389 7976
rect 7423 7973 7435 8007
rect 7377 7967 7435 7973
rect 9861 8007 9919 8013
rect 9861 7973 9873 8007
rect 9907 8004 9919 8007
rect 10134 8004 10140 8016
rect 9907 7976 10140 8004
rect 9907 7973 9919 7976
rect 9861 7967 9919 7973
rect 10134 7964 10140 7976
rect 10192 7964 10198 8016
rect 5796 7914 10304 7936
rect 5796 7862 5800 7914
rect 5852 7862 5864 7914
rect 5916 7862 5928 7914
rect 5980 7862 5992 7914
rect 6044 7862 6056 7914
rect 6108 7862 10304 7914
rect 5796 7840 10304 7862
rect 5537 7803 5595 7809
rect 5537 7769 5549 7803
rect 5583 7800 5595 7803
rect 5997 7803 6055 7809
rect 5997 7800 6009 7803
rect 5583 7772 6009 7800
rect 5583 7769 5595 7772
rect 5537 7763 5595 7769
rect 5997 7769 6009 7772
rect 6043 7769 6055 7803
rect 5997 7763 6055 7769
rect 7454 7744 7512 7750
rect 7009 7735 7067 7741
rect 6104 7704 6960 7732
rect 6104 7673 6132 7704
rect 6089 7667 6147 7673
rect 6089 7633 6101 7667
rect 6135 7633 6147 7667
rect 6089 7627 6147 7633
rect 6181 7667 6239 7673
rect 6181 7633 6193 7667
rect 6227 7633 6239 7667
rect 6362 7664 6368 7676
rect 6307 7636 6368 7664
rect 6181 7627 6239 7633
rect 5813 7599 5871 7605
rect 5813 7565 5825 7599
rect 5859 7596 5871 7599
rect 6196 7596 6224 7627
rect 6362 7624 6368 7636
rect 6420 7624 6426 7676
rect 5859 7568 6224 7596
rect 5859 7565 5871 7568
rect 5813 7559 5871 7565
rect 6454 7556 6460 7608
rect 6512 7596 6518 7608
rect 6549 7599 6607 7605
rect 6549 7596 6561 7599
rect 6512 7568 6561 7596
rect 6512 7556 6518 7568
rect 6549 7565 6561 7568
rect 6595 7565 6607 7599
rect 6549 7559 6607 7565
rect 6730 7556 6736 7608
rect 6788 7596 6794 7608
rect 6825 7599 6883 7605
rect 6825 7596 6837 7599
rect 6788 7568 6837 7596
rect 6788 7556 6794 7568
rect 6825 7565 6837 7568
rect 6871 7565 6883 7599
rect 6825 7559 6883 7565
rect 6641 7531 6699 7537
rect 6641 7528 6653 7531
rect 6472 7500 6653 7528
rect 6472 7494 6500 7500
rect 5736 7466 6500 7494
rect 6641 7497 6653 7500
rect 6687 7497 6699 7531
rect 6641 7491 6699 7497
rect 5736 7256 5764 7466
rect 6932 7460 6960 7704
rect 7009 7701 7021 7735
rect 7055 7732 7067 7735
rect 7454 7732 7466 7744
rect 7055 7710 7466 7732
rect 7500 7710 7512 7744
rect 7055 7704 7512 7710
rect 7055 7701 7067 7704
rect 7009 7695 7067 7701
rect 9030 7692 9036 7744
rect 9088 7732 9094 7744
rect 9217 7735 9275 7741
rect 9217 7732 9229 7735
rect 9088 7704 9229 7732
rect 9088 7692 9094 7704
rect 9217 7701 9229 7704
rect 9263 7701 9275 7735
rect 9217 7695 9275 7701
rect 7193 7667 7251 7673
rect 7193 7633 7205 7667
rect 7239 7664 7251 7667
rect 7466 7664 7472 7676
rect 7239 7636 7472 7664
rect 7239 7633 7251 7636
rect 7193 7627 7251 7633
rect 7466 7624 7472 7636
rect 7524 7624 7530 7676
rect 9401 7667 9459 7673
rect 9401 7633 9413 7667
rect 9447 7633 9459 7667
rect 9401 7627 9459 7633
rect 9677 7667 9735 7673
rect 9677 7633 9689 7667
rect 9723 7664 9735 7667
rect 10413 7667 10471 7673
rect 10413 7664 10425 7667
rect 9723 7636 10425 7664
rect 9723 7633 9735 7636
rect 9677 7627 9735 7633
rect 10413 7633 10425 7636
rect 10459 7633 10471 7667
rect 10413 7627 10471 7633
rect 9122 7556 9128 7608
rect 9180 7596 9186 7608
rect 9416 7596 9444 7627
rect 9180 7568 9444 7596
rect 9953 7599 10011 7605
rect 9180 7556 9186 7568
rect 9953 7565 9965 7599
rect 9999 7596 10011 7599
rect 10502 7596 10508 7608
rect 9999 7568 10508 7596
rect 9999 7565 10011 7568
rect 9953 7559 10011 7565
rect 10502 7556 10508 7568
rect 10560 7556 10566 7608
rect 9766 7528 9772 7540
rect 9711 7500 9772 7528
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 8573 7463 8631 7469
rect 8573 7460 8585 7463
rect 6932 7432 8585 7460
rect 8573 7429 8585 7432
rect 8619 7429 8631 7463
rect 8573 7423 8631 7429
rect 9674 7420 9680 7472
rect 9732 7460 9738 7472
rect 10137 7463 10195 7469
rect 10137 7460 10149 7463
rect 9732 7432 10149 7460
rect 9732 7420 9738 7432
rect 10137 7429 10149 7432
rect 10183 7429 10195 7463
rect 10137 7423 10195 7429
rect 5796 7370 10304 7392
rect 5796 7318 8182 7370
rect 8234 7318 8246 7370
rect 8298 7318 8310 7370
rect 8362 7318 8374 7370
rect 8426 7318 8438 7370
rect 8490 7318 8502 7370
rect 8554 7318 8566 7370
rect 8618 7318 8630 7370
rect 8682 7318 8694 7370
rect 8746 7318 8758 7370
rect 8810 7318 10304 7370
rect 5796 7296 10304 7318
rect 6089 7259 6147 7265
rect 6089 7256 6101 7259
rect 5736 7228 6101 7256
rect 6089 7225 6101 7228
rect 6135 7225 6147 7259
rect 6089 7219 6147 7225
rect 7926 7216 7932 7268
rect 7984 7256 7990 7268
rect 8297 7259 8355 7265
rect 8297 7256 8309 7259
rect 7984 7228 8309 7256
rect 7984 7216 7990 7228
rect 8297 7225 8309 7228
rect 8343 7225 8355 7259
rect 8297 7219 8355 7225
rect 8018 7148 8024 7200
rect 8076 7188 8082 7200
rect 8481 7191 8539 7197
rect 8481 7188 8493 7191
rect 8076 7160 8493 7188
rect 8076 7148 8082 7160
rect 8481 7157 8493 7160
rect 8527 7157 8539 7191
rect 8481 7151 8539 7157
rect 6641 7123 6699 7129
rect 6104 7092 6408 7120
rect 6104 7061 6132 7092
rect 6380 7064 6408 7092
rect 6641 7089 6653 7123
rect 6687 7120 6699 7123
rect 6730 7120 6736 7132
rect 6687 7092 6736 7120
rect 6687 7089 6699 7092
rect 6641 7083 6699 7089
rect 6730 7080 6736 7092
rect 6788 7080 6794 7132
rect 9858 7120 9864 7132
rect 9803 7092 9864 7120
rect 9858 7080 9864 7092
rect 9916 7080 9922 7132
rect 6089 7055 6147 7061
rect 6089 7021 6101 7055
rect 6135 7021 6147 7055
rect 6089 7015 6147 7021
rect 6181 7055 6239 7061
rect 6181 7021 6193 7055
rect 6227 7021 6239 7055
rect 6181 7015 6239 7021
rect 6196 6984 6224 7015
rect 6362 7012 6368 7064
rect 6420 7012 6426 7064
rect 6917 7055 6975 7061
rect 6917 7021 6929 7055
rect 6963 7052 6975 7055
rect 7466 7052 7472 7064
rect 6963 7024 7472 7052
rect 6963 7021 6975 7024
rect 6917 7015 6975 7021
rect 7466 7012 7472 7024
rect 7524 7012 7530 7064
rect 6546 6984 6552 6996
rect 6196 6956 6552 6984
rect 6546 6944 6552 6956
rect 6604 6944 6610 6996
rect 9674 6993 9680 6996
rect 6825 6987 6883 6993
rect 6825 6953 6837 6987
rect 6871 6984 6883 6987
rect 7178 6987 7236 6993
rect 7178 6984 7190 6987
rect 6871 6956 7190 6984
rect 6871 6953 6883 6956
rect 6825 6947 6883 6953
rect 7178 6953 7190 6956
rect 7224 6953 7236 6987
rect 7178 6947 7236 6953
rect 9616 6987 9680 6993
rect 9616 6953 9628 6987
rect 9662 6953 9680 6987
rect 9616 6947 9680 6953
rect 9674 6944 9680 6947
rect 9732 6944 9738 6996
rect 5796 6826 10304 6848
rect 5796 6774 5800 6826
rect 5852 6774 5864 6826
rect 5916 6774 5928 6826
rect 5980 6774 5992 6826
rect 6044 6774 6056 6826
rect 6108 6774 10304 6826
rect 5796 6752 10304 6774
rect 106 6672 112 6724
rect 164 6712 170 6724
rect 5997 6715 6055 6721
rect 5997 6712 6009 6715
rect 164 6684 6009 6712
rect 164 6672 170 6684
rect 5997 6681 6009 6684
rect 6043 6681 6055 6715
rect 5997 6675 6055 6681
rect 7454 6656 7512 6662
rect 7098 6604 7104 6656
rect 7156 6644 7162 6656
rect 7454 6644 7466 6656
rect 7156 6622 7466 6644
rect 7500 6622 7512 6656
rect 7156 6616 7512 6622
rect 7156 6604 7162 6616
rect 6362 6536 6368 6588
rect 6420 6576 6426 6588
rect 6641 6579 6699 6585
rect 6641 6576 6653 6579
rect 6420 6548 6653 6576
rect 6420 6536 6426 6548
rect 6641 6545 6653 6548
rect 6687 6545 6699 6579
rect 6641 6539 6699 6545
rect 7193 6579 7251 6585
rect 7193 6545 7205 6579
rect 7239 6576 7251 6579
rect 7466 6576 7472 6588
rect 7239 6548 7472 6576
rect 7239 6545 7251 6548
rect 7193 6539 7251 6545
rect 7466 6536 7472 6548
rect 7524 6536 7530 6588
rect 9950 6576 9956 6588
rect 9895 6548 9956 6576
rect 9950 6536 9956 6548
rect 10008 6536 10014 6588
rect 8588 6480 9628 6508
rect 6365 6443 6423 6449
rect 6365 6409 6377 6443
rect 6411 6440 6423 6443
rect 6411 6412 7236 6440
rect 6411 6409 6423 6412
rect 6365 6403 6423 6409
rect 6638 6372 6644 6384
rect 6583 6344 6644 6372
rect 6638 6332 6644 6344
rect 6696 6332 6702 6384
rect 7208 6372 7236 6412
rect 8588 6372 8616 6480
rect 9600 6440 9628 6480
rect 9769 6443 9827 6449
rect 9769 6440 9781 6443
rect 9600 6412 9781 6440
rect 9769 6409 9781 6412
rect 9815 6409 9827 6443
rect 9769 6403 9827 6409
rect 7208 6344 8616 6372
rect 5796 6282 10304 6304
rect 5796 6230 8182 6282
rect 8234 6230 8246 6282
rect 8298 6230 8310 6282
rect 8362 6230 8374 6282
rect 8426 6230 8438 6282
rect 8490 6230 8502 6282
rect 8554 6230 8566 6282
rect 8618 6230 8630 6282
rect 8682 6230 8694 6282
rect 8746 6230 8758 6282
rect 8810 6230 10304 6282
rect 5796 6208 10304 6230
rect 7009 6171 7067 6177
rect 7009 6137 7021 6171
rect 7055 6168 7067 6171
rect 7098 6168 7104 6180
rect 7055 6140 7104 6168
rect 7055 6137 7067 6140
rect 7009 6131 7067 6137
rect 7098 6128 7104 6140
rect 7156 6128 7162 6180
rect 7469 6171 7527 6177
rect 7469 6137 7481 6171
rect 7515 6168 7527 6171
rect 9585 6171 9643 6177
rect 9585 6168 9597 6171
rect 7515 6140 9597 6168
rect 7515 6137 7527 6140
rect 7469 6131 7527 6137
rect 9585 6137 9597 6140
rect 9631 6137 9643 6171
rect 9766 6168 9772 6180
rect 9711 6140 9772 6168
rect 9585 6131 9643 6137
rect 9766 6128 9772 6140
rect 9824 6128 9830 6180
rect 6638 6100 6644 6112
rect 6583 6072 6644 6100
rect 6638 6060 6644 6072
rect 6696 6060 6702 6112
rect 8205 6103 8263 6109
rect 8205 6069 8217 6103
rect 8251 6100 8263 6103
rect 8846 6100 8852 6112
rect 8251 6072 8852 6100
rect 8251 6069 8263 6072
rect 6822 6032 6828 6044
rect 5552 6004 6224 6032
rect 6767 6004 6828 6032
rect 198 5924 204 5976
rect 256 5964 262 5976
rect 5552 5964 5580 6004
rect 256 5936 5580 5964
rect 6196 5964 6224 6004
rect 6822 5992 6828 6004
rect 6880 6032 6886 6044
rect 7024 6038 7880 6066
rect 8205 6063 8263 6069
rect 8846 6060 8852 6072
rect 8904 6060 8910 6112
rect 7024 6032 7052 6038
rect 6880 6004 7052 6032
rect 7852 6032 7880 6038
rect 7852 6004 8064 6032
rect 6880 5992 6886 6004
rect 6365 5967 6423 5973
rect 6365 5964 6377 5967
rect 6196 5936 6377 5964
rect 256 5924 262 5936
rect 6365 5933 6377 5936
rect 6411 5933 6423 5967
rect 7377 5967 7435 5973
rect 7377 5964 7389 5967
rect 6365 5927 6423 5933
rect 6932 5936 7389 5964
rect 6273 5899 6331 5905
rect 6273 5865 6285 5899
rect 6319 5896 6331 5899
rect 6932 5896 6960 5936
rect 7377 5933 7389 5936
rect 7423 5933 7435 5967
rect 7742 5964 7748 5976
rect 7687 5936 7748 5964
rect 7377 5927 7435 5933
rect 7742 5924 7748 5936
rect 7800 5924 7806 5976
rect 8036 5973 8064 6004
rect 8110 5992 8116 6044
rect 8168 6032 8174 6044
rect 8481 6035 8539 6041
rect 8481 6032 8493 6035
rect 8168 6004 8493 6032
rect 8168 5992 8174 6004
rect 8481 6001 8493 6004
rect 8527 6001 8539 6035
rect 10134 6032 10140 6044
rect 8481 5995 8539 6001
rect 9876 6004 10140 6032
rect 8021 5967 8079 5973
rect 8021 5933 8033 5967
rect 8067 5964 8079 5967
rect 8849 5967 8907 5973
rect 8849 5964 8861 5967
rect 8067 5936 8861 5964
rect 8067 5933 8079 5936
rect 8021 5927 8079 5933
rect 8849 5933 8861 5936
rect 8895 5933 8907 5967
rect 8849 5927 8907 5933
rect 8938 5924 8944 5976
rect 8996 5964 9002 5976
rect 9122 5964 9128 5976
rect 8996 5936 9128 5964
rect 8996 5924 9002 5936
rect 9122 5924 9128 5936
rect 9180 5924 9186 5976
rect 9309 5967 9367 5973
rect 9309 5964 9321 5967
rect 9232 5936 9321 5964
rect 9232 5896 9260 5936
rect 9309 5933 9321 5936
rect 9355 5933 9367 5967
rect 9309 5927 9367 5933
rect 9398 5924 9404 5976
rect 9456 5964 9462 5976
rect 9585 5967 9643 5973
rect 9456 5936 9517 5964
rect 9456 5924 9462 5936
rect 9585 5933 9597 5967
rect 9631 5964 9643 5967
rect 9876 5964 9904 6004
rect 10134 5992 10140 6004
rect 10192 5992 10198 6044
rect 9631 5936 9904 5964
rect 9631 5933 9643 5936
rect 9585 5927 9643 5933
rect 9950 5924 9956 5976
rect 10008 5964 10014 5976
rect 10008 5936 10069 5964
rect 10008 5924 10014 5936
rect 10318 5896 10324 5908
rect 6319 5868 6960 5896
rect 9048 5868 9444 5896
rect 6319 5865 6331 5868
rect 6273 5859 6331 5865
rect 9048 5862 9076 5868
rect 14 5788 20 5840
rect 72 5828 78 5840
rect 6089 5831 6147 5837
rect 6089 5828 6101 5831
rect 72 5800 244 5828
rect 72 5788 78 5800
rect 216 5760 244 5800
rect 5644 5800 6101 5828
rect 5644 5760 5672 5800
rect 6089 5797 6101 5800
rect 6135 5797 6147 5831
rect 6089 5791 6147 5797
rect 6549 5831 6607 5837
rect 6549 5797 6561 5831
rect 6595 5828 6607 5831
rect 7116 5834 9076 5862
rect 9416 5862 9444 5868
rect 10152 5868 10324 5896
rect 10152 5862 10180 5868
rect 9416 5834 10180 5862
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 7116 5828 7144 5834
rect 6595 5800 7144 5828
rect 6595 5797 6607 5800
rect 6549 5791 6607 5797
rect 216 5732 5672 5760
rect 5796 5738 10304 5760
rect 5796 5686 5800 5738
rect 5852 5686 5864 5738
rect 5916 5686 5928 5738
rect 5980 5686 5992 5738
rect 6044 5686 6056 5738
rect 6108 5686 10304 5738
rect 5796 5664 10304 5686
rect 6454 5584 6460 5636
rect 6512 5624 6518 5636
rect 7742 5624 7748 5636
rect 6512 5596 6684 5624
rect 6512 5584 6518 5596
rect 6656 5488 6684 5596
rect 7576 5596 7748 5624
rect 7576 5488 7604 5596
rect 7742 5584 7748 5596
rect 7800 5584 7806 5636
rect 6656 5460 7604 5488
rect 14 76 20 128
rect 72 116 78 128
rect 1397 119 1455 125
rect 1397 116 1409 119
rect 72 88 1409 116
rect 72 76 78 88
rect 1397 85 1409 88
rect 1443 85 1455 119
rect 1397 79 1455 85
<< via1 >>
rect 20 17892 72 17944
rect 20 17008 72 17060
rect 5800 14390 5852 14442
rect 5864 14390 5916 14442
rect 5928 14390 5980 14442
rect 5992 14390 6044 14442
rect 6056 14390 6108 14442
rect 7196 14288 7248 14340
rect 7932 14220 7984 14272
rect 7748 14127 7800 14136
rect 7748 14093 7757 14127
rect 7757 14093 7791 14127
rect 7791 14093 7800 14127
rect 7748 14084 7800 14093
rect 8116 14084 8168 14136
rect 8852 14016 8904 14068
rect 7656 13948 7708 14000
rect 8024 13991 8076 14000
rect 8024 13957 8033 13991
rect 8033 13957 8067 13991
rect 8067 13957 8076 13991
rect 8024 13948 8076 13957
rect 9680 13948 9732 14000
rect 8182 13846 8234 13898
rect 8246 13846 8298 13898
rect 8310 13846 8362 13898
rect 8374 13846 8426 13898
rect 8438 13846 8490 13898
rect 8502 13846 8554 13898
rect 8566 13846 8618 13898
rect 8630 13846 8682 13898
rect 8694 13846 8746 13898
rect 8758 13846 8810 13898
rect 20 13744 72 13796
rect 7380 13744 7432 13796
rect 7932 13744 7984 13796
rect 15936 13744 15988 13796
rect 7656 13540 7708 13592
rect 8852 13540 8904 13592
rect 6736 13404 6788 13456
rect 8760 13404 8812 13456
rect 9220 13472 9272 13524
rect 5800 13302 5852 13354
rect 5864 13302 5916 13354
rect 5928 13302 5980 13354
rect 5992 13302 6044 13354
rect 6056 13302 6108 13354
rect 9220 13243 9272 13252
rect 9220 13209 9229 13243
rect 9229 13209 9263 13243
rect 9263 13209 9272 13243
rect 9220 13200 9272 13209
rect 20 13064 72 13116
rect 7012 13064 7064 13116
rect 7748 13064 7800 13116
rect 8852 12996 8904 13048
rect 9680 13064 9732 13116
rect 15752 13064 15804 13116
rect 6368 12903 6420 12912
rect 6368 12869 6377 12903
rect 6377 12869 6411 12903
rect 6411 12869 6420 12903
rect 6368 12860 6420 12869
rect 6736 12903 6788 12912
rect 6736 12869 6745 12903
rect 6745 12869 6779 12903
rect 6779 12869 6788 12903
rect 6736 12860 6788 12869
rect 9220 12860 9272 12912
rect 9404 12860 9456 12912
rect 8182 12758 8234 12810
rect 8246 12758 8298 12810
rect 8310 12758 8362 12810
rect 8374 12758 8426 12810
rect 8438 12758 8490 12810
rect 8502 12758 8554 12810
rect 8566 12758 8618 12810
rect 8630 12758 8682 12810
rect 8694 12758 8746 12810
rect 8758 12758 8810 12810
rect 7012 12656 7064 12708
rect 6000 12563 6052 12572
rect 6000 12529 6009 12563
rect 6009 12529 6043 12563
rect 6043 12529 6052 12563
rect 6000 12520 6052 12529
rect 6920 12384 6972 12436
rect 7748 12452 7800 12504
rect 8852 12452 8904 12504
rect 9036 12427 9088 12436
rect 9036 12393 9064 12427
rect 9064 12393 9088 12427
rect 9036 12384 9088 12393
rect 8668 12316 8720 12368
rect 5800 12214 5852 12266
rect 5864 12214 5916 12266
rect 5928 12214 5980 12266
rect 5992 12214 6044 12266
rect 6056 12214 6108 12266
rect 6368 11976 6420 12028
rect 6920 11976 6972 12028
rect 7196 12019 7248 12028
rect 7196 11985 7205 12019
rect 7205 11985 7239 12019
rect 7239 11985 7248 12019
rect 7196 11976 7248 11985
rect 7380 12019 7432 12028
rect 7380 11985 7389 12019
rect 7389 11985 7423 12019
rect 7423 11985 7432 12019
rect 7380 11976 7432 11985
rect 7656 11976 7708 12028
rect 6092 11951 6144 11960
rect 6092 11917 6101 11951
rect 6101 11917 6135 11951
rect 6135 11917 6144 11951
rect 6092 11908 6144 11917
rect 7564 11908 7616 11960
rect 6828 11772 6880 11824
rect 7840 11772 7892 11824
rect 9220 11840 9272 11892
rect 8182 11670 8234 11722
rect 8246 11670 8298 11722
rect 8310 11670 8362 11722
rect 8374 11670 8426 11722
rect 8438 11670 8490 11722
rect 8502 11670 8554 11722
rect 8566 11670 8618 11722
rect 8630 11670 8682 11722
rect 8694 11670 8746 11722
rect 8758 11670 8810 11722
rect 7656 11568 7708 11620
rect 7840 11500 7892 11552
rect 6092 11432 6144 11484
rect 7564 11364 7616 11416
rect 6828 11296 6880 11348
rect 7748 11296 7800 11348
rect 8484 11407 8536 11416
rect 8484 11373 8493 11407
rect 8493 11373 8527 11407
rect 8527 11373 8536 11407
rect 8484 11364 8536 11373
rect 8760 11407 8812 11416
rect 8760 11373 8788 11407
rect 8788 11373 8812 11407
rect 8760 11364 8812 11373
rect 6368 11228 6420 11280
rect 8852 11228 8904 11280
rect 9588 11228 9640 11280
rect 5800 11126 5852 11178
rect 5864 11126 5916 11178
rect 5928 11126 5980 11178
rect 5992 11126 6044 11178
rect 6056 11126 6108 11178
rect 6920 11024 6972 11076
rect 7104 10956 7156 11008
rect 6000 10931 6052 10940
rect 6000 10897 6009 10931
rect 6009 10897 6043 10931
rect 6043 10897 6052 10931
rect 6000 10888 6052 10897
rect 6184 10931 6236 10940
rect 6184 10897 6193 10931
rect 6193 10897 6227 10931
rect 6227 10897 6236 10931
rect 6184 10888 6236 10897
rect 6552 10931 6604 10940
rect 6552 10897 6561 10931
rect 6561 10897 6595 10931
rect 6595 10897 6604 10931
rect 6552 10888 6604 10897
rect 7656 10888 7708 10940
rect 8944 10820 8996 10872
rect 9404 10820 9456 10872
rect 6552 10795 6604 10804
rect 6552 10761 6561 10795
rect 6561 10761 6595 10795
rect 6595 10761 6604 10795
rect 6552 10752 6604 10761
rect 7472 10795 7524 10804
rect 7472 10761 7481 10795
rect 7481 10761 7515 10795
rect 7515 10761 7524 10795
rect 7472 10752 7524 10761
rect 8024 10752 8076 10804
rect 8182 10582 8234 10634
rect 8246 10582 8298 10634
rect 8310 10582 8362 10634
rect 8374 10582 8426 10634
rect 8438 10582 8490 10634
rect 8502 10582 8554 10634
rect 8566 10582 8618 10634
rect 8630 10582 8682 10634
rect 8694 10582 8746 10634
rect 8758 10582 8810 10634
rect 6276 10480 6328 10532
rect 5724 10344 5776 10396
rect 6736 10344 6788 10396
rect 6000 10276 6052 10328
rect 6184 10276 6236 10328
rect 6460 10276 6512 10328
rect 7104 10480 7156 10532
rect 10232 10412 10284 10464
rect 7472 10276 7524 10328
rect 8484 10319 8536 10328
rect 8484 10285 8493 10319
rect 8493 10285 8527 10319
rect 8527 10285 8536 10319
rect 8484 10276 8536 10285
rect 8760 10319 8812 10328
rect 8760 10285 8788 10319
rect 8788 10285 8812 10319
rect 8760 10276 8812 10285
rect 7196 10251 7248 10260
rect 7196 10217 7224 10251
rect 7224 10217 7248 10251
rect 7196 10208 7248 10217
rect 7012 10140 7064 10192
rect 9772 10208 9824 10260
rect 9588 10140 9640 10192
rect 5800 10038 5852 10090
rect 5864 10038 5916 10090
rect 5928 10038 5980 10090
rect 5992 10038 6044 10090
rect 6056 10038 6108 10090
rect 9128 9936 9180 9988
rect 7012 9868 7064 9920
rect 7748 9868 7800 9920
rect 6552 9843 6604 9852
rect 6552 9809 6561 9843
rect 6561 9809 6595 9843
rect 6595 9809 6604 9843
rect 6552 9800 6604 9809
rect 7472 9800 7524 9852
rect 8944 9843 8996 9852
rect 8944 9809 8953 9843
rect 8953 9809 8987 9843
rect 8987 9809 8996 9843
rect 8944 9800 8996 9809
rect 6828 9707 6880 9716
rect 6828 9673 6837 9707
rect 6837 9673 6871 9707
rect 6871 9673 6880 9707
rect 6828 9664 6880 9673
rect 10508 9664 10560 9716
rect 8182 9494 8234 9546
rect 8246 9494 8298 9546
rect 8310 9494 8362 9546
rect 8374 9494 8426 9546
rect 8438 9494 8490 9546
rect 8502 9494 8554 9546
rect 8566 9494 8618 9546
rect 8630 9494 8682 9546
rect 8694 9494 8746 9546
rect 8758 9494 8810 9546
rect 7380 9256 7432 9308
rect 7564 9299 7616 9308
rect 7564 9265 7573 9299
rect 7573 9265 7607 9299
rect 7607 9265 7616 9299
rect 7564 9256 7616 9265
rect 8484 9256 8536 9308
rect 8024 9231 8076 9240
rect 8024 9197 8033 9231
rect 8033 9197 8067 9231
rect 8067 9197 8076 9231
rect 8024 9188 8076 9197
rect 8852 9188 8904 9240
rect 6828 9120 6880 9172
rect 7748 9120 7800 9172
rect 8116 9120 8168 9172
rect 9220 9120 9272 9172
rect 7564 9052 7616 9104
rect 9956 9095 10008 9104
rect 9956 9061 9965 9095
rect 9965 9061 9999 9095
rect 9999 9061 10008 9095
rect 9956 9052 10008 9061
rect 20 8984 72 9036
rect 5800 8950 5852 9002
rect 5864 8950 5916 9002
rect 5928 8950 5980 9002
rect 5992 8950 6044 9002
rect 6056 8950 6108 9002
rect 6828 8891 6880 8900
rect 6828 8857 6837 8891
rect 6837 8857 6871 8891
rect 6871 8857 6880 8891
rect 6828 8848 6880 8857
rect 8484 8848 8536 8900
rect 9220 8848 9272 8900
rect 7564 8780 7616 8832
rect 10232 8780 10284 8832
rect 20 8712 72 8764
rect 6552 8712 6604 8764
rect 8668 8712 8720 8764
rect 6736 8644 6788 8696
rect 6920 8644 6972 8696
rect 10508 8644 10560 8696
rect 6460 8619 6512 8628
rect 6460 8585 6469 8619
rect 6469 8585 6503 8619
rect 6503 8585 6512 8619
rect 6460 8576 6512 8585
rect 9036 8508 9088 8560
rect 8182 8406 8234 8458
rect 8246 8406 8298 8458
rect 8310 8406 8362 8458
rect 8374 8406 8426 8458
rect 8438 8406 8490 8458
rect 8502 8406 8554 8458
rect 8566 8406 8618 8458
rect 8630 8406 8682 8458
rect 8694 8406 8746 8458
rect 8758 8406 8810 8458
rect 6552 8304 6604 8356
rect 7748 8279 7800 8288
rect 7748 8245 7757 8279
rect 7757 8245 7791 8279
rect 7791 8245 7800 8279
rect 7748 8236 7800 8245
rect 7380 8168 7432 8220
rect 7196 8032 7248 8084
rect 7932 8100 7984 8152
rect 8024 8143 8076 8152
rect 8024 8109 8033 8143
rect 8033 8109 8067 8143
rect 8067 8109 8076 8143
rect 8484 8143 8536 8152
rect 8024 8100 8076 8109
rect 8484 8109 8493 8143
rect 8493 8109 8527 8143
rect 8527 8109 8536 8143
rect 8484 8100 8536 8109
rect 9772 8100 9824 8152
rect 10232 8100 10284 8152
rect 8852 8032 8904 8084
rect 10324 8032 10376 8084
rect 10140 7964 10192 8016
rect 5800 7862 5852 7914
rect 5864 7862 5916 7914
rect 5928 7862 5980 7914
rect 5992 7862 6044 7914
rect 6056 7862 6108 7914
rect 6368 7667 6420 7676
rect 6368 7633 6377 7667
rect 6377 7633 6411 7667
rect 6411 7633 6420 7667
rect 6368 7624 6420 7633
rect 6460 7556 6512 7608
rect 6736 7556 6788 7608
rect 9036 7692 9088 7744
rect 7472 7624 7524 7676
rect 9128 7556 9180 7608
rect 10508 7556 10560 7608
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 9680 7420 9732 7472
rect 8182 7318 8234 7370
rect 8246 7318 8298 7370
rect 8310 7318 8362 7370
rect 8374 7318 8426 7370
rect 8438 7318 8490 7370
rect 8502 7318 8554 7370
rect 8566 7318 8618 7370
rect 8630 7318 8682 7370
rect 8694 7318 8746 7370
rect 8758 7318 8810 7370
rect 7932 7216 7984 7268
rect 8024 7148 8076 7200
rect 6736 7080 6788 7132
rect 9864 7123 9916 7132
rect 9864 7089 9873 7123
rect 9873 7089 9907 7123
rect 9907 7089 9916 7123
rect 9864 7080 9916 7089
rect 6368 7055 6420 7064
rect 6368 7021 6377 7055
rect 6377 7021 6411 7055
rect 6411 7021 6420 7055
rect 6368 7012 6420 7021
rect 7472 7012 7524 7064
rect 6552 6944 6604 6996
rect 9680 6944 9732 6996
rect 5800 6774 5852 6826
rect 5864 6774 5916 6826
rect 5928 6774 5980 6826
rect 5992 6774 6044 6826
rect 6056 6774 6108 6826
rect 112 6672 164 6724
rect 7104 6604 7156 6656
rect 6368 6536 6420 6588
rect 7472 6536 7524 6588
rect 9956 6579 10008 6588
rect 9956 6545 9965 6579
rect 9965 6545 9999 6579
rect 9999 6545 10008 6579
rect 9956 6536 10008 6545
rect 6644 6375 6696 6384
rect 6644 6341 6653 6375
rect 6653 6341 6687 6375
rect 6687 6341 6696 6375
rect 6644 6332 6696 6341
rect 8182 6230 8234 6282
rect 8246 6230 8298 6282
rect 8310 6230 8362 6282
rect 8374 6230 8426 6282
rect 8438 6230 8490 6282
rect 8502 6230 8554 6282
rect 8566 6230 8618 6282
rect 8630 6230 8682 6282
rect 8694 6230 8746 6282
rect 8758 6230 8810 6282
rect 7104 6128 7156 6180
rect 9772 6171 9824 6180
rect 9772 6137 9781 6171
rect 9781 6137 9815 6171
rect 9815 6137 9824 6171
rect 9772 6128 9824 6137
rect 6644 6103 6696 6112
rect 6644 6069 6653 6103
rect 6653 6069 6687 6103
rect 6687 6069 6696 6103
rect 6644 6060 6696 6069
rect 6828 6035 6880 6044
rect 204 5924 256 5976
rect 6828 6001 6837 6035
rect 6837 6001 6871 6035
rect 6871 6001 6880 6035
rect 8852 6060 8904 6112
rect 6828 5992 6880 6001
rect 7748 5967 7800 5976
rect 7748 5933 7757 5967
rect 7757 5933 7791 5967
rect 7791 5933 7800 5967
rect 7748 5924 7800 5933
rect 8116 5992 8168 6044
rect 8944 5924 8996 5976
rect 9128 5967 9180 5976
rect 9128 5933 9137 5967
rect 9137 5933 9171 5967
rect 9171 5933 9180 5967
rect 9128 5924 9180 5933
rect 9404 5967 9456 5976
rect 9404 5933 9413 5967
rect 9413 5933 9447 5967
rect 9447 5933 9456 5967
rect 9404 5924 9456 5933
rect 10140 5992 10192 6044
rect 9956 5967 10008 5976
rect 9956 5933 9965 5967
rect 9965 5933 9999 5967
rect 9999 5933 10008 5967
rect 9956 5924 10008 5933
rect 20 5788 72 5840
rect 10324 5856 10376 5908
rect 5800 5686 5852 5738
rect 5864 5686 5916 5738
rect 5928 5686 5980 5738
rect 5992 5686 6044 5738
rect 6056 5686 6108 5738
rect 6460 5584 6512 5636
rect 7748 5584 7800 5636
rect 20 76 72 128
<< metal2 >>
rect 0 20080 97 20108
rect 32 17944 60 20080
rect 14 17892 20 17944
rect 72 17892 78 17944
rect 0 17836 97 17864
rect 32 17066 60 17836
rect 20 17060 72 17066
rect 20 17002 72 17008
rect 0 15592 97 15620
rect 32 13802 60 15592
rect 20 13796 72 13802
rect 20 13738 72 13744
rect 0 13348 97 13376
rect 32 13122 60 13348
rect 20 13116 72 13122
rect 20 13058 72 13064
rect 216 12493 244 20128
rect 5796 14444 6112 14464
rect 5796 14442 5806 14444
rect 5862 14442 5886 14444
rect 5942 14442 5966 14444
rect 6022 14442 6046 14444
rect 6102 14442 6112 14444
rect 5796 14390 5800 14442
rect 5862 14390 5864 14442
rect 6044 14390 6046 14442
rect 6108 14390 6112 14442
rect 5796 14388 5806 14390
rect 5862 14388 5886 14390
rect 5942 14388 5966 14390
rect 6022 14388 6046 14390
rect 6102 14388 6112 14390
rect 5796 14368 6112 14388
rect 7196 14340 7248 14346
rect 8036 14328 8064 20128
rect 15856 19904 15884 20128
rect 16003 20080 16100 20108
rect 15764 19876 15884 19904
rect 8036 14300 8156 14328
rect 7196 14282 7248 14288
rect 7208 13920 7236 14282
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 7748 14136 7800 14142
rect 7748 14078 7800 14084
rect 7656 14000 7708 14006
rect 7656 13942 7708 13948
rect 7116 13892 7236 13920
rect 6736 13456 6788 13462
rect 6736 13398 6788 13404
rect 5796 13356 6112 13376
rect 5796 13354 5806 13356
rect 5862 13354 5886 13356
rect 5942 13354 5966 13356
rect 6022 13354 6046 13356
rect 6102 13354 6112 13356
rect 5796 13302 5800 13354
rect 5862 13302 5864 13354
rect 6044 13302 6046 13354
rect 6108 13302 6112 13354
rect 5796 13300 5806 13302
rect 5862 13300 5886 13302
rect 5942 13300 5966 13302
rect 6022 13300 6046 13302
rect 6102 13300 6112 13302
rect 5796 13280 6112 13300
rect 6748 12918 6776 13398
rect 7116 13308 7144 13892
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7392 13376 7420 13738
rect 7668 13598 7696 13942
rect 7760 13920 7788 14078
rect 7760 13892 7834 13920
rect 7656 13592 7708 13598
rect 7656 13534 7708 13540
rect 7392 13348 7512 13376
rect 7116 13280 7236 13308
rect 7012 13116 7064 13122
rect 7012 13058 7064 13064
rect 6368 12912 6420 12918
rect 6368 12854 6420 12860
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6000 12572 6052 12578
rect 6052 12532 6224 12560
rect 6000 12514 6052 12520
rect 202 12484 258 12493
rect 202 12419 258 12428
rect 5796 12268 6112 12288
rect 5796 12266 5806 12268
rect 5862 12266 5886 12268
rect 5942 12266 5966 12268
rect 6022 12266 6046 12268
rect 6102 12266 6112 12268
rect 5796 12214 5800 12266
rect 5862 12214 5864 12266
rect 6044 12214 6046 12266
rect 6108 12214 6112 12266
rect 6196 12249 6224 12532
rect 5796 12212 5806 12214
rect 5862 12212 5886 12214
rect 5942 12212 5966 12214
rect 6022 12212 6046 12214
rect 6102 12212 6112 12214
rect 5796 12192 6112 12212
rect 6182 12240 6238 12249
rect 6182 12175 6238 12184
rect 6380 12034 6408 12854
rect 6550 12484 6606 12493
rect 6550 12419 6606 12428
rect 6368 12028 6420 12034
rect 6368 11970 6420 11976
rect 6092 11960 6144 11966
rect 6092 11902 6144 11908
rect 6104 11490 6132 11902
rect 6092 11484 6144 11490
rect 5736 11444 6092 11472
rect 0 11104 97 11132
rect 32 9036 60 11104
rect 5736 10402 5764 11444
rect 6380 11472 6408 11970
rect 6092 11426 6144 11432
rect 6288 11444 6408 11472
rect 5796 11180 6112 11200
rect 5796 11178 5806 11180
rect 5862 11178 5886 11180
rect 5942 11178 5966 11180
rect 6022 11178 6046 11180
rect 6102 11178 6112 11180
rect 5796 11126 5800 11178
rect 5862 11126 5864 11178
rect 6044 11126 6046 11178
rect 6108 11126 6112 11178
rect 5796 11124 5806 11126
rect 5862 11124 5886 11126
rect 5942 11124 5966 11126
rect 6022 11124 6046 11126
rect 6102 11124 6112 11126
rect 5796 11104 6112 11124
rect 6182 11020 6238 11029
rect 6000 10940 6052 10946
rect 6000 10882 6052 10888
rect 6182 10940 6238 10964
rect 6182 10888 6184 10940
rect 6236 10888 6238 10940
rect 6182 10882 6238 10888
rect 5724 10396 5776 10402
rect 5724 10338 5776 10344
rect 6012 10334 6040 10882
rect 6288 10538 6316 11444
rect 6368 11280 6420 11286
rect 6564 11273 6592 12419
rect 6368 11222 6420 11228
rect 6550 11264 6606 11273
rect 6276 10532 6328 10538
rect 6380 10520 6408 11222
rect 6550 11199 6606 11208
rect 6564 10946 6592 11199
rect 6748 11029 6776 12854
rect 7024 12714 7052 13058
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6932 12034 6960 12378
rect 7208 12034 7236 13280
rect 7484 12220 7512 13348
rect 7806 13308 7834 13892
rect 7944 13802 7972 14214
rect 8128 14142 8156 14300
rect 8116 14136 8168 14142
rect 8116 14078 8168 14084
rect 8852 14068 8904 14074
rect 8852 14010 8904 14016
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 7932 13796 7984 13802
rect 7932 13738 7984 13744
rect 8036 13716 8064 13942
rect 8160 13900 8832 13920
rect 8160 13898 8188 13900
rect 8244 13898 8268 13900
rect 8324 13898 8348 13900
rect 8404 13898 8428 13900
rect 8484 13898 8508 13900
rect 8564 13898 8588 13900
rect 8644 13898 8668 13900
rect 8724 13898 8748 13900
rect 8804 13898 8832 13900
rect 8160 13846 8182 13898
rect 8244 13846 8246 13898
rect 8426 13846 8428 13898
rect 8490 13846 8502 13898
rect 8564 13846 8566 13898
rect 8746 13846 8748 13898
rect 8810 13846 8832 13898
rect 8160 13844 8188 13846
rect 8244 13844 8268 13846
rect 8324 13844 8348 13846
rect 8404 13844 8428 13846
rect 8484 13844 8508 13846
rect 8564 13844 8588 13846
rect 8644 13844 8668 13846
rect 8724 13844 8748 13846
rect 8804 13844 8832 13846
rect 8160 13824 8832 13844
rect 8864 13784 8892 14010
rect 9680 14000 9732 14006
rect 9680 13942 9732 13948
rect 8772 13756 8892 13784
rect 8036 13688 8156 13716
rect 7760 13280 7834 13308
rect 7760 13122 7788 13280
rect 8128 13240 8156 13688
rect 8772 13462 8800 13756
rect 8852 13592 8904 13598
rect 8852 13534 8904 13540
rect 8760 13456 8812 13462
rect 8760 13398 8812 13404
rect 8036 13212 8156 13240
rect 7748 13116 7800 13122
rect 7748 13058 7800 13064
rect 7760 12510 7788 13058
rect 7748 12504 7800 12510
rect 7748 12446 7800 12452
rect 7392 12192 7512 12220
rect 7392 12034 7420 12192
rect 6920 12028 6972 12034
rect 6920 11970 6972 11976
rect 7196 12028 7248 12034
rect 7196 11970 7248 11976
rect 7380 12028 7432 12034
rect 7380 11970 7432 11976
rect 7656 12028 7708 12034
rect 7656 11970 7708 11976
rect 6828 11824 6880 11830
rect 6932 11812 6960 11970
rect 7564 11960 7616 11966
rect 7564 11902 7616 11908
rect 6932 11784 7052 11812
rect 6828 11766 6880 11772
rect 6840 11354 6868 11766
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 7024 11268 7052 11784
rect 7576 11422 7604 11902
rect 7668 11626 7696 11970
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7564 11416 7616 11422
rect 6932 11240 7052 11268
rect 7484 11376 7564 11404
rect 6932 11082 6960 11240
rect 6920 11076 6972 11082
rect 6734 11020 6790 11029
rect 6920 11018 6972 11024
rect 6734 10955 6790 10964
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 6552 10940 6604 10946
rect 6552 10882 6604 10888
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6380 10492 6500 10520
rect 6276 10474 6328 10480
rect 6472 10334 6500 10492
rect 6000 10328 6052 10334
rect 6000 10270 6052 10276
rect 6184 10328 6236 10334
rect 6184 10270 6236 10276
rect 6460 10328 6512 10334
rect 6460 10270 6512 10276
rect 5796 10092 6112 10112
rect 5796 10090 5806 10092
rect 5862 10090 5886 10092
rect 5942 10090 5966 10092
rect 6022 10090 6046 10092
rect 6102 10090 6112 10092
rect 5796 10038 5800 10090
rect 5862 10038 5864 10090
rect 6044 10038 6046 10090
rect 6108 10038 6112 10090
rect 5796 10036 5806 10038
rect 5862 10036 5886 10038
rect 5942 10036 5966 10038
rect 6022 10036 6046 10038
rect 6102 10036 6112 10038
rect 5796 10016 6112 10036
rect 6196 9199 6224 10270
rect 6564 9858 6592 10746
rect 7116 10538 7144 10950
rect 7484 10810 7512 11376
rect 7564 11358 7616 11364
rect 7760 11354 7788 12446
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 7852 11558 7880 11766
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7654 11264 7710 11273
rect 7654 11199 7710 11208
rect 7668 10946 7696 11199
rect 7656 10940 7708 10946
rect 7656 10882 7708 10888
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 6736 10396 6788 10402
rect 6736 10338 6788 10344
rect 6748 10175 6776 10338
rect 7484 10334 7512 10746
rect 7472 10328 7524 10334
rect 7472 10270 7524 10276
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7012 10192 7064 10198
rect 6734 10166 6790 10175
rect 7012 10134 7064 10140
rect 6734 10101 6790 10110
rect 6552 9852 6604 9858
rect 6552 9794 6604 9800
rect 6748 9636 6776 10101
rect 6918 9922 6974 9931
rect 7024 9926 7052 10134
rect 6918 9857 6974 9866
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 6828 9716 6880 9722
rect 6932 9704 6960 9857
rect 6880 9676 6960 9704
rect 7208 9704 7236 10202
rect 7484 9858 7512 10270
rect 7760 10175 7788 11290
rect 8036 10810 8064 13212
rect 8864 13054 8892 13534
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9232 13258 9260 13466
rect 9220 13252 9272 13258
rect 9220 13194 9272 13200
rect 9692 13122 9720 13942
rect 15764 13648 15792 19876
rect 15936 13796 15988 13802
rect 16037 13784 16065 20080
rect 15988 13756 16065 13784
rect 15936 13738 15988 13744
rect 15764 13620 15884 13648
rect 9680 13116 9732 13122
rect 9680 13058 9732 13064
rect 15752 13116 15804 13122
rect 15856 13104 15884 13620
rect 15804 13076 15884 13104
rect 15752 13058 15804 13064
rect 8852 13048 8904 13054
rect 8852 12990 8904 12996
rect 8160 12812 8832 12832
rect 8160 12810 8188 12812
rect 8244 12810 8268 12812
rect 8324 12810 8348 12812
rect 8404 12810 8428 12812
rect 8484 12810 8508 12812
rect 8564 12810 8588 12812
rect 8644 12810 8668 12812
rect 8724 12810 8748 12812
rect 8804 12810 8832 12812
rect 8160 12758 8182 12810
rect 8244 12758 8246 12810
rect 8426 12758 8428 12810
rect 8490 12758 8502 12810
rect 8564 12758 8566 12810
rect 8746 12758 8748 12810
rect 8810 12758 8832 12810
rect 8160 12756 8188 12758
rect 8244 12756 8268 12758
rect 8324 12756 8348 12758
rect 8404 12756 8428 12758
rect 8484 12756 8508 12758
rect 8564 12756 8588 12758
rect 8644 12756 8668 12758
rect 8724 12756 8748 12758
rect 8804 12756 8832 12758
rect 8160 12736 8832 12756
rect 8864 12510 8892 12990
rect 9220 12912 9272 12918
rect 9220 12854 9272 12860
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 8852 12504 8904 12510
rect 8852 12446 8904 12452
rect 8668 12368 8720 12374
rect 8668 12310 8720 12316
rect 8680 12016 8708 12310
rect 8864 12249 8892 12446
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 8850 12240 8906 12249
rect 8850 12175 8906 12184
rect 8680 11988 8892 12016
rect 8160 11724 8832 11744
rect 8160 11722 8188 11724
rect 8244 11722 8268 11724
rect 8324 11722 8348 11724
rect 8404 11722 8428 11724
rect 8484 11722 8508 11724
rect 8564 11722 8588 11724
rect 8644 11722 8668 11724
rect 8724 11722 8748 11724
rect 8804 11722 8832 11724
rect 8160 11670 8182 11722
rect 8244 11670 8246 11722
rect 8426 11670 8428 11722
rect 8490 11670 8502 11722
rect 8564 11670 8566 11722
rect 8746 11670 8748 11722
rect 8810 11670 8832 11722
rect 8160 11668 8188 11670
rect 8244 11668 8268 11670
rect 8324 11668 8348 11670
rect 8404 11668 8428 11670
rect 8484 11668 8508 11670
rect 8564 11668 8588 11670
rect 8644 11668 8668 11670
rect 8724 11668 8748 11670
rect 8804 11668 8832 11670
rect 8160 11648 8832 11668
rect 8864 11608 8892 11988
rect 9048 11676 9076 12378
rect 9232 11898 9260 12854
rect 9416 12696 9444 12854
rect 9416 12668 9536 12696
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9508 11744 9536 12668
rect 9416 11716 9536 11744
rect 9048 11648 9168 11676
rect 8772 11580 8892 11608
rect 8772 11422 8800 11580
rect 8484 11416 8536 11422
rect 8482 11386 8484 11395
rect 8760 11416 8812 11422
rect 8536 11386 8538 11395
rect 8760 11358 8812 11364
rect 8482 11321 8538 11330
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 8160 10636 8832 10656
rect 8160 10634 8188 10636
rect 8244 10634 8268 10636
rect 8324 10634 8348 10636
rect 8404 10634 8428 10636
rect 8484 10634 8508 10636
rect 8564 10634 8588 10636
rect 8644 10634 8668 10636
rect 8724 10634 8748 10636
rect 8804 10634 8832 10636
rect 8160 10582 8182 10634
rect 8244 10582 8246 10634
rect 8426 10582 8428 10634
rect 8490 10582 8502 10634
rect 8564 10582 8566 10634
rect 8746 10582 8748 10634
rect 8810 10582 8832 10634
rect 8160 10580 8188 10582
rect 8244 10580 8268 10582
rect 8324 10580 8348 10582
rect 8404 10580 8428 10582
rect 8484 10580 8508 10582
rect 8564 10580 8588 10582
rect 8644 10580 8668 10582
rect 8724 10580 8748 10582
rect 8804 10580 8832 10582
rect 8160 10560 8832 10580
rect 8864 10520 8892 11222
rect 8944 10872 8996 10878
rect 8944 10814 8996 10820
rect 8772 10492 8892 10520
rect 8772 10334 8800 10492
rect 8484 10328 8536 10334
rect 8482 10288 8484 10297
rect 8760 10328 8812 10334
rect 8536 10288 8538 10297
rect 8760 10270 8812 10276
rect 8482 10223 8538 10232
rect 7746 10166 7802 10175
rect 7746 10101 7802 10110
rect 7760 9926 7788 10101
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 8850 9922 8906 9931
rect 7472 9852 7524 9858
rect 7472 9794 7524 9800
rect 7208 9676 7328 9704
rect 6828 9658 6880 9664
rect 6564 9608 6776 9636
rect 6182 9190 6238 9199
rect 6182 9125 6238 9134
rect 14 8984 20 9036
rect 72 8984 78 9036
rect 5796 9004 6112 9024
rect 5796 9002 5806 9004
rect 5862 9002 5886 9004
rect 5942 9002 5966 9004
rect 6022 9002 6046 9004
rect 6102 9002 6112 9004
rect 0 8928 97 8956
rect 5796 8950 5800 9002
rect 5862 8950 5864 9002
rect 6044 8950 6046 9002
rect 6108 8950 6112 9002
rect 5796 8948 5806 8950
rect 5862 8948 5886 8950
rect 5942 8948 5966 8950
rect 6022 8948 6046 8950
rect 6102 8948 6112 8950
rect 5796 8928 6112 8948
rect 32 8770 60 8928
rect 20 8764 72 8770
rect 20 8706 72 8712
rect 5796 7916 6112 7936
rect 5796 7914 5806 7916
rect 5862 7914 5886 7916
rect 5942 7914 5966 7916
rect 6022 7914 6046 7916
rect 6102 7914 6112 7916
rect 5796 7862 5800 7914
rect 5862 7862 5864 7914
rect 6044 7862 6046 7914
rect 6108 7862 6112 7914
rect 5796 7860 5806 7862
rect 5862 7860 5886 7862
rect 5942 7860 5966 7862
rect 6022 7860 6046 7862
rect 6102 7860 6112 7862
rect 5796 7840 6112 7860
rect 6196 7664 6224 9125
rect 6564 8956 6592 9608
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6564 8928 6776 8956
rect 6552 8764 6604 8770
rect 6552 8706 6604 8712
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6472 8412 6500 8570
rect 6380 8384 6500 8412
rect 6380 7868 6408 8384
rect 6564 8362 6592 8706
rect 6748 8702 6776 8928
rect 6840 8906 6868 9114
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 6736 8696 6788 8702
rect 6932 8696 6960 9676
rect 6914 8644 6920 8696
rect 6972 8644 6978 8696
rect 6736 8638 6788 8644
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6564 8140 6592 8298
rect 6564 8112 6638 8140
rect 6380 7840 6500 7868
rect 6368 7676 6420 7682
rect 6196 7636 6368 7664
rect 6368 7618 6420 7624
rect 6380 7070 6408 7618
rect 6472 7614 6500 7840
rect 6460 7608 6512 7614
rect 6460 7550 6512 7556
rect 6610 7460 6638 8112
rect 6748 7936 6776 8638
rect 6932 8345 6960 8644
rect 6918 8336 6974 8345
rect 6918 8271 6974 8280
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7208 7936 7236 8026
rect 6748 7908 7236 7936
rect 6748 7614 6776 7908
rect 7300 7800 7328 9676
rect 7378 9434 7434 9443
rect 7378 9369 7434 9378
rect 7392 9314 7420 9369
rect 7380 9308 7432 9314
rect 7380 9250 7432 9256
rect 7378 8336 7434 8345
rect 7378 8271 7434 8280
rect 7392 8226 7420 8271
rect 7380 8220 7432 8226
rect 7380 8162 7432 8168
rect 7484 8101 7512 9794
rect 7564 9308 7616 9314
rect 7760 9296 7788 9862
rect 8850 9857 8906 9866
rect 8956 9858 8984 10814
rect 9140 10656 9168 11648
rect 9416 10878 9444 11716
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9404 10872 9456 10878
rect 9404 10814 9456 10820
rect 9140 10628 9260 10656
rect 9232 10180 9260 10628
rect 9600 10198 9628 11222
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9140 10152 9260 10180
rect 9588 10192 9640 10198
rect 9140 9994 9168 10152
rect 9588 10134 9640 10140
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 8160 9548 8832 9568
rect 8160 9546 8188 9548
rect 8244 9546 8268 9548
rect 8324 9546 8348 9548
rect 8404 9546 8428 9548
rect 8484 9546 8508 9548
rect 8564 9546 8588 9548
rect 8644 9546 8668 9548
rect 8724 9546 8748 9548
rect 8804 9546 8832 9548
rect 8160 9494 8182 9546
rect 8244 9494 8246 9546
rect 8426 9494 8428 9546
rect 8490 9494 8502 9546
rect 8564 9494 8566 9546
rect 8746 9494 8748 9546
rect 8810 9494 8832 9546
rect 8160 9492 8188 9494
rect 8244 9492 8268 9494
rect 8324 9492 8348 9494
rect 8404 9492 8428 9494
rect 8484 9492 8508 9494
rect 8564 9492 8588 9494
rect 8644 9492 8668 9494
rect 8724 9492 8748 9494
rect 8804 9492 8832 9494
rect 8160 9472 8832 9492
rect 7616 9268 7788 9296
rect 8484 9308 8536 9314
rect 7564 9250 7616 9256
rect 8484 9250 8536 9256
rect 8024 9240 8076 9246
rect 8022 9190 8024 9199
rect 8076 9190 8078 9199
rect 7748 9172 7800 9178
rect 8022 9125 8078 9134
rect 8116 9172 8168 9178
rect 7748 9114 7800 9120
rect 8116 9114 8168 9120
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7576 8838 7604 9046
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7760 8294 7788 9114
rect 8128 8616 8156 9114
rect 8496 8906 8524 9250
rect 8864 9246 8892 9857
rect 8944 9852 8996 9858
rect 8944 9794 8996 9800
rect 8852 9240 8904 9246
rect 8666 9190 8722 9199
rect 8852 9182 8904 9188
rect 9218 9190 9274 9199
rect 8666 9125 8722 9134
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 8680 8770 8708 9125
rect 8864 9024 8892 9182
rect 9218 9125 9220 9134
rect 9272 9125 9274 9134
rect 9220 9114 9272 9120
rect 9232 9102 9260 9114
rect 8864 8996 9628 9024
rect 9218 8946 9274 8955
rect 9218 8881 9220 8890
rect 9272 8881 9274 8890
rect 9220 8842 9272 8848
rect 8668 8764 8720 8770
rect 8668 8706 8720 8712
rect 8036 8588 8156 8616
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 8036 8158 8064 8588
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 8160 8460 8832 8480
rect 8160 8458 8188 8460
rect 8244 8458 8268 8460
rect 8324 8458 8348 8460
rect 8404 8458 8428 8460
rect 8484 8458 8508 8460
rect 8564 8458 8588 8460
rect 8644 8458 8668 8460
rect 8724 8458 8748 8460
rect 8804 8458 8832 8460
rect 8160 8406 8182 8458
rect 8244 8406 8246 8458
rect 8426 8406 8428 8458
rect 8490 8406 8502 8458
rect 8564 8406 8566 8458
rect 8746 8406 8748 8458
rect 8810 8406 8832 8458
rect 8160 8404 8188 8406
rect 8244 8404 8268 8406
rect 8324 8404 8348 8406
rect 8404 8404 8428 8406
rect 8484 8404 8508 8406
rect 8564 8404 8588 8406
rect 8644 8404 8668 8406
rect 8724 8404 8748 8406
rect 8804 8404 8832 8406
rect 8160 8384 8832 8404
rect 7932 8152 7984 8158
rect 7470 8092 7526 8101
rect 7932 8094 7984 8100
rect 8024 8152 8076 8158
rect 8484 8152 8536 8158
rect 8024 8094 8076 8100
rect 8482 8100 8484 8101
rect 8536 8100 8538 8101
rect 7470 8027 7526 8036
rect 7208 7772 7328 7800
rect 6736 7608 6788 7614
rect 6736 7550 6788 7556
rect 6564 7432 6638 7460
rect 6368 7064 6420 7070
rect 6368 7006 6420 7012
rect 5796 6828 6112 6848
rect 5796 6826 5806 6828
rect 5862 6826 5886 6828
rect 5942 6826 5966 6828
rect 6022 6826 6046 6828
rect 6102 6826 6112 6828
rect 5796 6774 5800 6826
rect 5862 6774 5864 6826
rect 6044 6774 6046 6826
rect 6108 6774 6112 6826
rect 5796 6772 5806 6774
rect 5862 6772 5886 6774
rect 5942 6772 5966 6774
rect 6022 6772 6046 6774
rect 6102 6772 6112 6774
rect 5796 6752 6112 6772
rect 112 6724 164 6730
rect 0 6684 112 6712
rect 112 6666 164 6672
rect 6380 6594 6408 7006
rect 6564 7002 6592 7432
rect 6748 7138 6776 7550
rect 6736 7132 6788 7138
rect 6736 7074 6788 7080
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6368 6588 6420 6594
rect 6368 6530 6420 6536
rect 204 5976 256 5982
rect 204 5918 256 5924
rect 20 5840 72 5846
rect 20 5782 72 5788
rect 32 4468 60 5782
rect 216 5760 244 5918
rect 6380 5896 6408 6530
rect 6748 6440 6776 7074
rect 7208 6848 7236 7772
rect 7484 7682 7512 8027
rect 7944 7936 7972 8094
rect 7852 7908 7972 7936
rect 7472 7676 7524 7682
rect 7472 7618 7524 7624
rect 7484 7070 7512 7618
rect 7852 7460 7880 7908
rect 7852 7432 7972 7460
rect 7944 7274 7972 7432
rect 7932 7268 7984 7274
rect 7932 7210 7984 7216
rect 8036 7206 8064 8094
rect 8482 8092 8538 8100
rect 8482 8027 8538 8036
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8160 7372 8832 7392
rect 8160 7370 8188 7372
rect 8244 7370 8268 7372
rect 8324 7370 8348 7372
rect 8404 7370 8428 7372
rect 8484 7370 8508 7372
rect 8564 7370 8588 7372
rect 8644 7370 8668 7372
rect 8724 7370 8748 7372
rect 8804 7370 8832 7372
rect 8160 7318 8182 7370
rect 8244 7318 8246 7370
rect 8426 7318 8428 7370
rect 8490 7318 8502 7370
rect 8564 7318 8566 7370
rect 8746 7318 8748 7370
rect 8810 7318 8832 7370
rect 8160 7316 8188 7318
rect 8244 7316 8268 7318
rect 8324 7316 8348 7318
rect 8404 7316 8428 7318
rect 8484 7316 8508 7318
rect 8564 7316 8588 7318
rect 8644 7316 8668 7318
rect 8724 7316 8748 7318
rect 8804 7316 8832 7318
rect 8160 7296 8832 7316
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 7472 7064 7524 7070
rect 7472 7006 7524 7012
rect 7208 6820 7328 6848
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 6748 6412 6868 6440
rect 6644 6384 6696 6390
rect 6644 6326 6696 6332
rect 6656 6118 6684 6326
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6840 6050 6868 6412
rect 7116 6186 7144 6598
rect 7104 6180 7156 6186
rect 7300 6168 7328 6820
rect 7484 6594 7512 7006
rect 7472 6588 7524 6594
rect 7472 6530 7524 6536
rect 8160 6284 8832 6304
rect 8160 6282 8188 6284
rect 8244 6282 8268 6284
rect 8324 6282 8348 6284
rect 8404 6282 8428 6284
rect 8484 6282 8508 6284
rect 8564 6282 8588 6284
rect 8644 6282 8668 6284
rect 8724 6282 8748 6284
rect 8804 6282 8832 6284
rect 8160 6230 8182 6282
rect 8244 6230 8246 6282
rect 8426 6230 8428 6282
rect 8490 6230 8502 6282
rect 8564 6230 8566 6282
rect 8746 6230 8748 6282
rect 8810 6230 8832 6282
rect 8160 6228 8188 6230
rect 8244 6228 8268 6230
rect 8324 6228 8348 6230
rect 8404 6228 8428 6230
rect 8484 6228 8508 6230
rect 8564 6228 8588 6230
rect 8644 6228 8668 6230
rect 8724 6228 8748 6230
rect 8804 6228 8832 6230
rect 8160 6208 8832 6228
rect 7300 6140 8156 6168
rect 7104 6122 7156 6128
rect 8128 6050 8156 6140
rect 8864 6118 8892 8026
rect 9048 7936 9076 8502
rect 9048 7908 9260 7936
rect 9048 7750 9076 7908
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9232 7664 9260 7908
rect 9232 7636 9444 7664
rect 9128 7608 9180 7614
rect 9128 7550 9180 7556
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 6828 6044 6880 6050
rect 8116 6044 8168 6050
rect 6828 5986 6880 5992
rect 7746 6018 7802 6027
rect 8116 5986 8168 5992
rect 8942 6018 8998 6027
rect 7746 5953 7748 5962
rect 7800 5953 7802 5962
rect 9140 5982 9168 7550
rect 9416 5982 9444 7636
rect 9600 7247 9628 8996
rect 9784 8158 9812 10202
rect 9956 9104 10008 9110
rect 9956 9046 10008 9052
rect 9772 8152 9824 8158
rect 9772 8094 9824 8100
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9586 7238 9642 7247
rect 9586 7173 9642 7182
rect 9692 7002 9720 7414
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9784 6186 9812 7482
rect 9862 7238 9918 7247
rect 9862 7173 9918 7182
rect 9876 7138 9904 7173
rect 9864 7132 9916 7138
rect 9864 7074 9916 7080
rect 9968 6594 9996 9046
rect 10244 8838 10272 10406
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10244 8158 10272 8774
rect 10520 8702 10548 9658
rect 10508 8696 10560 8702
rect 10508 8638 10560 8644
rect 10232 8152 10284 8158
rect 10232 8094 10284 8100
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 9956 6588 10008 6594
rect 9956 6530 10008 6536
rect 9772 6180 9824 6186
rect 9772 6122 9824 6128
rect 10152 6050 10180 7958
rect 10336 7392 10364 8026
rect 10520 7614 10548 8638
rect 10508 7608 10560 7614
rect 10508 7550 10560 7556
rect 10336 7364 10456 7392
rect 10428 6100 10456 7364
rect 10336 6072 10456 6100
rect 10140 6044 10192 6050
rect 9954 6018 10010 6027
rect 8942 5953 8944 5962
rect 7748 5918 7800 5924
rect 8996 5953 8998 5962
rect 9128 5976 9180 5982
rect 8944 5918 8996 5924
rect 9128 5918 9180 5924
rect 9404 5976 9456 5982
rect 10140 5986 10192 5992
rect 9954 5953 9956 5962
rect 9404 5918 9456 5924
rect 10008 5953 10010 5962
rect 9956 5918 10008 5924
rect 6380 5868 6500 5896
rect 216 5732 336 5760
rect 0 4440 97 4468
rect 308 4400 336 5732
rect 5796 5740 6112 5760
rect 5796 5738 5806 5740
rect 5862 5738 5886 5740
rect 5942 5738 5966 5740
rect 6022 5738 6046 5740
rect 6102 5738 6112 5740
rect 5796 5686 5800 5738
rect 5862 5686 5864 5738
rect 6044 5686 6046 5738
rect 6108 5686 6112 5738
rect 5796 5684 5806 5686
rect 5862 5684 5886 5686
rect 5942 5684 5966 5686
rect 6022 5684 6046 5686
rect 6102 5684 6112 5686
rect 5796 5664 6112 5684
rect 6472 5642 6500 5868
rect 7760 5642 7788 5918
rect 10336 5914 10364 6072
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 6460 5636 6512 5642
rect 6460 5578 6512 5584
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 216 4372 336 4400
rect 216 2224 244 4372
rect 0 2196 244 2224
rect 14 76 20 128
rect 72 76 78 128
rect 32 48 60 76
rect 0 20 97 48
<< via2 >>
rect 5806 14442 5862 14444
rect 5886 14442 5942 14444
rect 5966 14442 6022 14444
rect 6046 14442 6102 14444
rect 5806 14390 5852 14442
rect 5852 14390 5862 14442
rect 5886 14390 5916 14442
rect 5916 14390 5928 14442
rect 5928 14390 5942 14442
rect 5966 14390 5980 14442
rect 5980 14390 5992 14442
rect 5992 14390 6022 14442
rect 6046 14390 6056 14442
rect 6056 14390 6102 14442
rect 5806 14388 5862 14390
rect 5886 14388 5942 14390
rect 5966 14388 6022 14390
rect 6046 14388 6102 14390
rect 5806 13354 5862 13356
rect 5886 13354 5942 13356
rect 5966 13354 6022 13356
rect 6046 13354 6102 13356
rect 5806 13302 5852 13354
rect 5852 13302 5862 13354
rect 5886 13302 5916 13354
rect 5916 13302 5928 13354
rect 5928 13302 5942 13354
rect 5966 13302 5980 13354
rect 5980 13302 5992 13354
rect 5992 13302 6022 13354
rect 6046 13302 6056 13354
rect 6056 13302 6102 13354
rect 5806 13300 5862 13302
rect 5886 13300 5942 13302
rect 5966 13300 6022 13302
rect 6046 13300 6102 13302
rect 202 12428 258 12484
rect 5806 12266 5862 12268
rect 5886 12266 5942 12268
rect 5966 12266 6022 12268
rect 6046 12266 6102 12268
rect 5806 12214 5852 12266
rect 5852 12214 5862 12266
rect 5886 12214 5916 12266
rect 5916 12214 5928 12266
rect 5928 12214 5942 12266
rect 5966 12214 5980 12266
rect 5980 12214 5992 12266
rect 5992 12214 6022 12266
rect 6046 12214 6056 12266
rect 6056 12214 6102 12266
rect 5806 12212 5862 12214
rect 5886 12212 5942 12214
rect 5966 12212 6022 12214
rect 6046 12212 6102 12214
rect 6182 12184 6238 12240
rect 6550 12428 6606 12484
rect 5806 11178 5862 11180
rect 5886 11178 5942 11180
rect 5966 11178 6022 11180
rect 6046 11178 6102 11180
rect 5806 11126 5852 11178
rect 5852 11126 5862 11178
rect 5886 11126 5916 11178
rect 5916 11126 5928 11178
rect 5928 11126 5942 11178
rect 5966 11126 5980 11178
rect 5980 11126 5992 11178
rect 5992 11126 6022 11178
rect 6046 11126 6056 11178
rect 6056 11126 6102 11178
rect 5806 11124 5862 11126
rect 5886 11124 5942 11126
rect 5966 11124 6022 11126
rect 6046 11124 6102 11126
rect 6182 10964 6238 11020
rect 6550 11208 6606 11264
rect 8188 13898 8244 13900
rect 8268 13898 8324 13900
rect 8348 13898 8404 13900
rect 8428 13898 8484 13900
rect 8508 13898 8564 13900
rect 8588 13898 8644 13900
rect 8668 13898 8724 13900
rect 8748 13898 8804 13900
rect 8188 13846 8234 13898
rect 8234 13846 8244 13898
rect 8268 13846 8298 13898
rect 8298 13846 8310 13898
rect 8310 13846 8324 13898
rect 8348 13846 8362 13898
rect 8362 13846 8374 13898
rect 8374 13846 8404 13898
rect 8428 13846 8438 13898
rect 8438 13846 8484 13898
rect 8508 13846 8554 13898
rect 8554 13846 8564 13898
rect 8588 13846 8618 13898
rect 8618 13846 8630 13898
rect 8630 13846 8644 13898
rect 8668 13846 8682 13898
rect 8682 13846 8694 13898
rect 8694 13846 8724 13898
rect 8748 13846 8758 13898
rect 8758 13846 8804 13898
rect 8188 13844 8244 13846
rect 8268 13844 8324 13846
rect 8348 13844 8404 13846
rect 8428 13844 8484 13846
rect 8508 13844 8564 13846
rect 8588 13844 8644 13846
rect 8668 13844 8724 13846
rect 8748 13844 8804 13846
rect 6734 10964 6790 11020
rect 5806 10090 5862 10092
rect 5886 10090 5942 10092
rect 5966 10090 6022 10092
rect 6046 10090 6102 10092
rect 5806 10038 5852 10090
rect 5852 10038 5862 10090
rect 5886 10038 5916 10090
rect 5916 10038 5928 10090
rect 5928 10038 5942 10090
rect 5966 10038 5980 10090
rect 5980 10038 5992 10090
rect 5992 10038 6022 10090
rect 6046 10038 6056 10090
rect 6056 10038 6102 10090
rect 5806 10036 5862 10038
rect 5886 10036 5942 10038
rect 5966 10036 6022 10038
rect 6046 10036 6102 10038
rect 7654 11208 7710 11264
rect 6734 10110 6790 10166
rect 6918 9866 6974 9922
rect 8188 12810 8244 12812
rect 8268 12810 8324 12812
rect 8348 12810 8404 12812
rect 8428 12810 8484 12812
rect 8508 12810 8564 12812
rect 8588 12810 8644 12812
rect 8668 12810 8724 12812
rect 8748 12810 8804 12812
rect 8188 12758 8234 12810
rect 8234 12758 8244 12810
rect 8268 12758 8298 12810
rect 8298 12758 8310 12810
rect 8310 12758 8324 12810
rect 8348 12758 8362 12810
rect 8362 12758 8374 12810
rect 8374 12758 8404 12810
rect 8428 12758 8438 12810
rect 8438 12758 8484 12810
rect 8508 12758 8554 12810
rect 8554 12758 8564 12810
rect 8588 12758 8618 12810
rect 8618 12758 8630 12810
rect 8630 12758 8644 12810
rect 8668 12758 8682 12810
rect 8682 12758 8694 12810
rect 8694 12758 8724 12810
rect 8748 12758 8758 12810
rect 8758 12758 8804 12810
rect 8188 12756 8244 12758
rect 8268 12756 8324 12758
rect 8348 12756 8404 12758
rect 8428 12756 8484 12758
rect 8508 12756 8564 12758
rect 8588 12756 8644 12758
rect 8668 12756 8724 12758
rect 8748 12756 8804 12758
rect 8850 12184 8906 12240
rect 8188 11722 8244 11724
rect 8268 11722 8324 11724
rect 8348 11722 8404 11724
rect 8428 11722 8484 11724
rect 8508 11722 8564 11724
rect 8588 11722 8644 11724
rect 8668 11722 8724 11724
rect 8748 11722 8804 11724
rect 8188 11670 8234 11722
rect 8234 11670 8244 11722
rect 8268 11670 8298 11722
rect 8298 11670 8310 11722
rect 8310 11670 8324 11722
rect 8348 11670 8362 11722
rect 8362 11670 8374 11722
rect 8374 11670 8404 11722
rect 8428 11670 8438 11722
rect 8438 11670 8484 11722
rect 8508 11670 8554 11722
rect 8554 11670 8564 11722
rect 8588 11670 8618 11722
rect 8618 11670 8630 11722
rect 8630 11670 8644 11722
rect 8668 11670 8682 11722
rect 8682 11670 8694 11722
rect 8694 11670 8724 11722
rect 8748 11670 8758 11722
rect 8758 11670 8804 11722
rect 8188 11668 8244 11670
rect 8268 11668 8324 11670
rect 8348 11668 8404 11670
rect 8428 11668 8484 11670
rect 8508 11668 8564 11670
rect 8588 11668 8644 11670
rect 8668 11668 8724 11670
rect 8748 11668 8804 11670
rect 8482 11364 8484 11386
rect 8484 11364 8536 11386
rect 8536 11364 8538 11386
rect 8482 11330 8538 11364
rect 8188 10634 8244 10636
rect 8268 10634 8324 10636
rect 8348 10634 8404 10636
rect 8428 10634 8484 10636
rect 8508 10634 8564 10636
rect 8588 10634 8644 10636
rect 8668 10634 8724 10636
rect 8748 10634 8804 10636
rect 8188 10582 8234 10634
rect 8234 10582 8244 10634
rect 8268 10582 8298 10634
rect 8298 10582 8310 10634
rect 8310 10582 8324 10634
rect 8348 10582 8362 10634
rect 8362 10582 8374 10634
rect 8374 10582 8404 10634
rect 8428 10582 8438 10634
rect 8438 10582 8484 10634
rect 8508 10582 8554 10634
rect 8554 10582 8564 10634
rect 8588 10582 8618 10634
rect 8618 10582 8630 10634
rect 8630 10582 8644 10634
rect 8668 10582 8682 10634
rect 8682 10582 8694 10634
rect 8694 10582 8724 10634
rect 8748 10582 8758 10634
rect 8758 10582 8804 10634
rect 8188 10580 8244 10582
rect 8268 10580 8324 10582
rect 8348 10580 8404 10582
rect 8428 10580 8484 10582
rect 8508 10580 8564 10582
rect 8588 10580 8644 10582
rect 8668 10580 8724 10582
rect 8748 10580 8804 10582
rect 8482 10276 8484 10288
rect 8484 10276 8536 10288
rect 8536 10276 8538 10288
rect 8482 10232 8538 10276
rect 7746 10110 7802 10166
rect 8850 9866 8906 9922
rect 6182 9134 6238 9190
rect 5806 9002 5862 9004
rect 5886 9002 5942 9004
rect 5966 9002 6022 9004
rect 6046 9002 6102 9004
rect 5806 8950 5852 9002
rect 5852 8950 5862 9002
rect 5886 8950 5916 9002
rect 5916 8950 5928 9002
rect 5928 8950 5942 9002
rect 5966 8950 5980 9002
rect 5980 8950 5992 9002
rect 5992 8950 6022 9002
rect 6046 8950 6056 9002
rect 6056 8950 6102 9002
rect 5806 8948 5862 8950
rect 5886 8948 5942 8950
rect 5966 8948 6022 8950
rect 6046 8948 6102 8950
rect 5806 7914 5862 7916
rect 5886 7914 5942 7916
rect 5966 7914 6022 7916
rect 6046 7914 6102 7916
rect 5806 7862 5852 7914
rect 5852 7862 5862 7914
rect 5886 7862 5916 7914
rect 5916 7862 5928 7914
rect 5928 7862 5942 7914
rect 5966 7862 5980 7914
rect 5980 7862 5992 7914
rect 5992 7862 6022 7914
rect 6046 7862 6056 7914
rect 6056 7862 6102 7914
rect 5806 7860 5862 7862
rect 5886 7860 5942 7862
rect 5966 7860 6022 7862
rect 6046 7860 6102 7862
rect 6918 8280 6974 8336
rect 7378 9378 7434 9434
rect 7378 8280 7434 8336
rect 8188 9546 8244 9548
rect 8268 9546 8324 9548
rect 8348 9546 8404 9548
rect 8428 9546 8484 9548
rect 8508 9546 8564 9548
rect 8588 9546 8644 9548
rect 8668 9546 8724 9548
rect 8748 9546 8804 9548
rect 8188 9494 8234 9546
rect 8234 9494 8244 9546
rect 8268 9494 8298 9546
rect 8298 9494 8310 9546
rect 8310 9494 8324 9546
rect 8348 9494 8362 9546
rect 8362 9494 8374 9546
rect 8374 9494 8404 9546
rect 8428 9494 8438 9546
rect 8438 9494 8484 9546
rect 8508 9494 8554 9546
rect 8554 9494 8564 9546
rect 8588 9494 8618 9546
rect 8618 9494 8630 9546
rect 8630 9494 8644 9546
rect 8668 9494 8682 9546
rect 8682 9494 8694 9546
rect 8694 9494 8724 9546
rect 8748 9494 8758 9546
rect 8758 9494 8804 9546
rect 8188 9492 8244 9494
rect 8268 9492 8324 9494
rect 8348 9492 8404 9494
rect 8428 9492 8484 9494
rect 8508 9492 8564 9494
rect 8588 9492 8644 9494
rect 8668 9492 8724 9494
rect 8748 9492 8804 9494
rect 8022 9188 8024 9190
rect 8024 9188 8076 9190
rect 8076 9188 8078 9190
rect 8022 9134 8078 9188
rect 8666 9134 8722 9190
rect 9218 9172 9274 9190
rect 9218 9134 9220 9172
rect 9220 9134 9272 9172
rect 9272 9134 9274 9172
rect 9218 8900 9274 8946
rect 9218 8890 9220 8900
rect 9220 8890 9272 8900
rect 9272 8890 9274 8900
rect 8188 8458 8244 8460
rect 8268 8458 8324 8460
rect 8348 8458 8404 8460
rect 8428 8458 8484 8460
rect 8508 8458 8564 8460
rect 8588 8458 8644 8460
rect 8668 8458 8724 8460
rect 8748 8458 8804 8460
rect 8188 8406 8234 8458
rect 8234 8406 8244 8458
rect 8268 8406 8298 8458
rect 8298 8406 8310 8458
rect 8310 8406 8324 8458
rect 8348 8406 8362 8458
rect 8362 8406 8374 8458
rect 8374 8406 8404 8458
rect 8428 8406 8438 8458
rect 8438 8406 8484 8458
rect 8508 8406 8554 8458
rect 8554 8406 8564 8458
rect 8588 8406 8618 8458
rect 8618 8406 8630 8458
rect 8630 8406 8644 8458
rect 8668 8406 8682 8458
rect 8682 8406 8694 8458
rect 8694 8406 8724 8458
rect 8748 8406 8758 8458
rect 8758 8406 8804 8458
rect 8188 8404 8244 8406
rect 8268 8404 8324 8406
rect 8348 8404 8404 8406
rect 8428 8404 8484 8406
rect 8508 8404 8564 8406
rect 8588 8404 8644 8406
rect 8668 8404 8724 8406
rect 8748 8404 8804 8406
rect 7470 8036 7526 8092
rect 5806 6826 5862 6828
rect 5886 6826 5942 6828
rect 5966 6826 6022 6828
rect 6046 6826 6102 6828
rect 5806 6774 5852 6826
rect 5852 6774 5862 6826
rect 5886 6774 5916 6826
rect 5916 6774 5928 6826
rect 5928 6774 5942 6826
rect 5966 6774 5980 6826
rect 5980 6774 5992 6826
rect 5992 6774 6022 6826
rect 6046 6774 6056 6826
rect 6056 6774 6102 6826
rect 5806 6772 5862 6774
rect 5886 6772 5942 6774
rect 5966 6772 6022 6774
rect 6046 6772 6102 6774
rect 8482 8036 8538 8092
rect 8188 7370 8244 7372
rect 8268 7370 8324 7372
rect 8348 7370 8404 7372
rect 8428 7370 8484 7372
rect 8508 7370 8564 7372
rect 8588 7370 8644 7372
rect 8668 7370 8724 7372
rect 8748 7370 8804 7372
rect 8188 7318 8234 7370
rect 8234 7318 8244 7370
rect 8268 7318 8298 7370
rect 8298 7318 8310 7370
rect 8310 7318 8324 7370
rect 8348 7318 8362 7370
rect 8362 7318 8374 7370
rect 8374 7318 8404 7370
rect 8428 7318 8438 7370
rect 8438 7318 8484 7370
rect 8508 7318 8554 7370
rect 8554 7318 8564 7370
rect 8588 7318 8618 7370
rect 8618 7318 8630 7370
rect 8630 7318 8644 7370
rect 8668 7318 8682 7370
rect 8682 7318 8694 7370
rect 8694 7318 8724 7370
rect 8748 7318 8758 7370
rect 8758 7318 8804 7370
rect 8188 7316 8244 7318
rect 8268 7316 8324 7318
rect 8348 7316 8404 7318
rect 8428 7316 8484 7318
rect 8508 7316 8564 7318
rect 8588 7316 8644 7318
rect 8668 7316 8724 7318
rect 8748 7316 8804 7318
rect 8188 6282 8244 6284
rect 8268 6282 8324 6284
rect 8348 6282 8404 6284
rect 8428 6282 8484 6284
rect 8508 6282 8564 6284
rect 8588 6282 8644 6284
rect 8668 6282 8724 6284
rect 8748 6282 8804 6284
rect 8188 6230 8234 6282
rect 8234 6230 8244 6282
rect 8268 6230 8298 6282
rect 8298 6230 8310 6282
rect 8310 6230 8324 6282
rect 8348 6230 8362 6282
rect 8362 6230 8374 6282
rect 8374 6230 8404 6282
rect 8428 6230 8438 6282
rect 8438 6230 8484 6282
rect 8508 6230 8554 6282
rect 8554 6230 8564 6282
rect 8588 6230 8618 6282
rect 8618 6230 8630 6282
rect 8630 6230 8644 6282
rect 8668 6230 8682 6282
rect 8682 6230 8694 6282
rect 8694 6230 8724 6282
rect 8748 6230 8758 6282
rect 8758 6230 8804 6282
rect 8188 6228 8244 6230
rect 8268 6228 8324 6230
rect 8348 6228 8404 6230
rect 8428 6228 8484 6230
rect 8508 6228 8564 6230
rect 8588 6228 8644 6230
rect 8668 6228 8724 6230
rect 8748 6228 8804 6230
rect 7746 5976 7802 6018
rect 7746 5962 7748 5976
rect 7748 5962 7800 5976
rect 7800 5962 7802 5976
rect 8942 5976 8998 6018
rect 9586 7182 9642 7238
rect 9862 7182 9918 7238
rect 8942 5962 8944 5976
rect 8944 5962 8996 5976
rect 8996 5962 8998 5976
rect 9954 5976 10010 6018
rect 9954 5962 9956 5976
rect 9956 5962 10008 5976
rect 10008 5962 10010 5976
rect 5806 5738 5862 5740
rect 5886 5738 5942 5740
rect 5966 5738 6022 5740
rect 6046 5738 6102 5740
rect 5806 5686 5852 5738
rect 5852 5686 5862 5738
rect 5886 5686 5916 5738
rect 5916 5686 5928 5738
rect 5928 5686 5942 5738
rect 5966 5686 5980 5738
rect 5980 5686 5992 5738
rect 5992 5686 6022 5738
rect 6046 5686 6056 5738
rect 6056 5686 6102 5738
rect 5806 5684 5862 5686
rect 5886 5684 5942 5686
rect 5966 5684 6022 5686
rect 6046 5684 6102 5686
<< metal3 >>
rect 5796 14448 6112 14464
rect 5796 14384 5802 14448
rect 5866 14384 5882 14448
rect 5946 14384 5962 14448
rect 6026 14384 6042 14448
rect 6106 14384 6112 14448
rect 5796 14368 6112 14384
rect 8160 13904 8832 13920
rect 8160 13840 8184 13904
rect 8248 13840 8264 13904
rect 8328 13840 8344 13904
rect 8408 13840 8424 13904
rect 8488 13840 8504 13904
rect 8568 13840 8584 13904
rect 8648 13840 8664 13904
rect 8728 13840 8744 13904
rect 8808 13840 8832 13904
rect 8160 13824 8832 13840
rect 5796 13360 6112 13376
rect 5796 13296 5802 13360
rect 5866 13296 5882 13360
rect 5946 13296 5962 13360
rect 6026 13296 6042 13360
rect 6106 13296 6112 13360
rect 5796 13280 6112 13296
rect 8160 12816 8832 12832
rect 8160 12752 8184 12816
rect 8248 12752 8264 12816
rect 8328 12752 8344 12816
rect 8408 12752 8424 12816
rect 8488 12752 8504 12816
rect 8568 12752 8584 12816
rect 8648 12752 8664 12816
rect 8728 12752 8744 12816
rect 8808 12752 8832 12816
rect 8160 12736 8832 12752
rect 197 12486 263 12489
rect 6545 12486 6611 12489
rect 197 12484 6611 12486
rect 197 12428 202 12484
rect 258 12428 6550 12484
rect 6606 12428 6611 12484
rect 197 12426 6611 12428
rect 197 12423 263 12426
rect 6545 12423 6611 12426
rect 5796 12272 6112 12288
rect 5796 12208 5802 12272
rect 5866 12208 5882 12272
rect 5946 12208 5962 12272
rect 6026 12208 6042 12272
rect 6106 12208 6112 12272
rect 5796 12192 6112 12208
rect 6177 12242 6243 12245
rect 7874 12242 7880 12244
rect 6177 12240 7880 12242
rect 6177 12184 6182 12240
rect 6238 12184 7880 12240
rect 6177 12182 7880 12184
rect 6177 12179 6243 12182
rect 7874 12180 7880 12182
rect 7944 12242 7950 12244
rect 8845 12242 8911 12245
rect 7944 12240 8911 12242
rect 7944 12184 8850 12240
rect 8906 12184 8911 12240
rect 7944 12182 8911 12184
rect 7944 12180 7950 12182
rect 8845 12179 8911 12182
rect 8160 11728 8832 11744
rect 8160 11664 8184 11728
rect 8248 11664 8264 11728
rect 8328 11664 8344 11728
rect 8408 11664 8424 11728
rect 8488 11664 8504 11728
rect 8568 11664 8584 11728
rect 8648 11664 8664 11728
rect 8728 11664 8744 11728
rect 8808 11664 8832 11728
rect 8160 11648 8832 11664
rect 7874 11326 7880 11390
rect 7944 11388 7950 11390
rect 8477 11388 8543 11391
rect 7944 11386 8543 11388
rect 7944 11330 8482 11386
rect 8538 11330 8543 11386
rect 7944 11328 8543 11330
rect 7944 11326 7950 11328
rect 8477 11325 8543 11328
rect 6545 11266 6611 11269
rect 7649 11266 7715 11269
rect 6545 11264 7715 11266
rect 6545 11208 6550 11264
rect 6606 11208 7654 11264
rect 7710 11208 7715 11264
rect 6545 11206 7715 11208
rect 6545 11203 6611 11206
rect 7649 11203 7715 11206
rect 5796 11184 6112 11200
rect 5796 11120 5802 11184
rect 5866 11120 5882 11184
rect 5946 11120 5962 11184
rect 6026 11120 6042 11184
rect 6106 11120 6112 11184
rect 5796 11104 6112 11120
rect 6177 11022 6243 11025
rect 6729 11022 6795 11025
rect 6177 11020 6795 11022
rect 6177 10964 6182 11020
rect 6238 10964 6734 11020
rect 6790 10964 6795 11020
rect 6177 10962 6795 10964
rect 6177 10959 6243 10962
rect 6729 10959 6795 10962
rect 8160 10640 8832 10656
rect 8160 10576 8184 10640
rect 8248 10576 8264 10640
rect 8328 10576 8344 10640
rect 8408 10576 8424 10640
rect 8488 10576 8504 10640
rect 8568 10576 8584 10640
rect 8648 10576 8664 10640
rect 8728 10576 8744 10640
rect 8808 10576 8832 10640
rect 8160 10560 8832 10576
rect 7874 10228 7880 10292
rect 7944 10290 7950 10292
rect 8477 10290 8543 10293
rect 7944 10288 8543 10290
rect 7944 10232 8482 10288
rect 8538 10232 8543 10288
rect 7944 10230 8543 10232
rect 7944 10228 7950 10230
rect 8477 10227 8543 10230
rect 6729 10168 6795 10171
rect 7741 10168 7807 10171
rect 6729 10166 7807 10168
rect 5796 10096 6112 10112
rect 6729 10110 6734 10166
rect 6790 10110 7746 10166
rect 7802 10110 7807 10166
rect 6729 10108 7807 10110
rect 6729 10105 6795 10108
rect 7741 10105 7807 10108
rect 5796 10032 5802 10096
rect 5866 10032 5882 10096
rect 5946 10032 5962 10096
rect 6026 10032 6042 10096
rect 6106 10032 6112 10096
rect 5796 10016 6112 10032
rect 6913 9924 6979 9927
rect 7874 9924 7880 9926
rect 6913 9922 7880 9924
rect 6913 9866 6918 9922
rect 6974 9866 7880 9922
rect 6913 9864 7880 9866
rect 6913 9861 6979 9864
rect 7376 9439 7436 9864
rect 7874 9862 7880 9864
rect 7944 9924 7950 9926
rect 8845 9924 8911 9927
rect 7944 9922 8911 9924
rect 7944 9866 8850 9922
rect 8906 9866 8911 9922
rect 7944 9864 8911 9866
rect 7944 9862 7950 9864
rect 8845 9861 8911 9864
rect 8160 9552 8832 9568
rect 8160 9488 8184 9552
rect 8248 9488 8264 9552
rect 8328 9488 8344 9552
rect 8408 9488 8424 9552
rect 8488 9488 8504 9552
rect 8568 9488 8584 9552
rect 8648 9488 8664 9552
rect 8728 9488 8744 9552
rect 8808 9488 8832 9552
rect 8160 9472 8832 9488
rect 7373 9434 7439 9439
rect 7373 9378 7378 9434
rect 7434 9378 7439 9434
rect 7373 9373 7439 9378
rect 6177 9192 6243 9195
rect 8017 9192 8083 9195
rect 8661 9192 8727 9195
rect 6177 9190 8727 9192
rect 6177 9134 6182 9190
rect 6238 9134 8022 9190
rect 8078 9134 8666 9190
rect 8722 9134 8727 9190
rect 6177 9132 8727 9134
rect 6177 9129 6243 9132
rect 8017 9129 8083 9132
rect 8661 9129 8727 9132
rect 9213 9190 9279 9195
rect 9213 9134 9218 9190
rect 9274 9134 9279 9190
rect 9213 9129 9279 9134
rect 5796 9008 6112 9024
rect 5796 8944 5802 9008
rect 5866 8944 5882 9008
rect 5946 8944 5962 9008
rect 6026 8944 6042 9008
rect 6106 8944 6112 9008
rect 9216 8951 9276 9129
rect 5796 8928 6112 8944
rect 9213 8946 9279 8951
rect 9213 8890 9218 8946
rect 9274 8890 9279 8946
rect 9213 8885 9279 8890
rect 8160 8464 8832 8480
rect 8160 8400 8184 8464
rect 8248 8400 8264 8464
rect 8328 8400 8344 8464
rect 8408 8400 8424 8464
rect 8488 8400 8504 8464
rect 8568 8400 8584 8464
rect 8648 8400 8664 8464
rect 8728 8400 8744 8464
rect 8808 8400 8832 8464
rect 8160 8384 8832 8400
rect 6913 8338 6979 8341
rect 7373 8338 7439 8341
rect 6913 8336 7439 8338
rect 6913 8280 6918 8336
rect 6974 8280 7378 8336
rect 7434 8280 7439 8336
rect 6913 8278 7439 8280
rect 6913 8275 6979 8278
rect 7373 8275 7439 8278
rect 7465 8094 7531 8097
rect 8477 8094 8543 8097
rect 7465 8092 8543 8094
rect 7465 8036 7470 8092
rect 7526 8036 8482 8092
rect 8538 8036 8543 8092
rect 7465 8034 8543 8036
rect 7465 8031 7531 8034
rect 8477 8031 8543 8034
rect 5796 7920 6112 7936
rect 5796 7856 5802 7920
rect 5866 7856 5882 7920
rect 5946 7856 5962 7920
rect 6026 7856 6042 7920
rect 6106 7856 6112 7920
rect 5796 7840 6112 7856
rect 8160 7376 8832 7392
rect 8160 7312 8184 7376
rect 8248 7312 8264 7376
rect 8328 7312 8344 7376
rect 8408 7312 8424 7376
rect 8488 7312 8504 7376
rect 8568 7312 8584 7376
rect 8648 7312 8664 7376
rect 8728 7312 8744 7376
rect 8808 7312 8832 7376
rect 8160 7296 8832 7312
rect 9581 7240 9647 7243
rect 9857 7240 9923 7243
rect 9581 7238 9923 7240
rect 9581 7182 9586 7238
rect 9642 7182 9862 7238
rect 9918 7182 9923 7238
rect 9581 7180 9923 7182
rect 9581 7177 9647 7180
rect 9857 7177 9923 7180
rect 5796 6832 6112 6848
rect 5796 6768 5802 6832
rect 5866 6768 5882 6832
rect 5946 6768 5962 6832
rect 6026 6768 6042 6832
rect 6106 6768 6112 6832
rect 5796 6752 6112 6768
rect 8160 6288 8832 6304
rect 8160 6224 8184 6288
rect 8248 6224 8264 6288
rect 8328 6224 8344 6288
rect 8408 6224 8424 6288
rect 8488 6224 8504 6288
rect 8568 6224 8584 6288
rect 8648 6224 8664 6288
rect 8728 6224 8744 6288
rect 8808 6224 8832 6288
rect 8160 6208 8832 6224
rect 7741 6020 7807 6023
rect 8937 6020 9003 6023
rect 9949 6020 10015 6023
rect 7741 6018 10015 6020
rect 7741 5962 7746 6018
rect 7802 5962 8942 6018
rect 8998 5962 9954 6018
rect 10010 5962 10015 6018
rect 7741 5960 10015 5962
rect 7741 5957 7807 5960
rect 8937 5957 9003 5960
rect 9949 5957 10015 5960
rect 5796 5744 6112 5760
rect 5796 5680 5802 5744
rect 5866 5680 5882 5744
rect 5946 5680 5962 5744
rect 6026 5680 6042 5744
rect 6106 5680 6112 5744
rect 5796 5664 6112 5680
<< via3 >>
rect 5802 14444 5866 14448
rect 5802 14388 5806 14444
rect 5806 14388 5862 14444
rect 5862 14388 5866 14444
rect 5802 14384 5866 14388
rect 5882 14444 5946 14448
rect 5882 14388 5886 14444
rect 5886 14388 5942 14444
rect 5942 14388 5946 14444
rect 5882 14384 5946 14388
rect 5962 14444 6026 14448
rect 5962 14388 5966 14444
rect 5966 14388 6022 14444
rect 6022 14388 6026 14444
rect 5962 14384 6026 14388
rect 6042 14444 6106 14448
rect 6042 14388 6046 14444
rect 6046 14388 6102 14444
rect 6102 14388 6106 14444
rect 6042 14384 6106 14388
rect 8184 13900 8248 13904
rect 8184 13844 8188 13900
rect 8188 13844 8244 13900
rect 8244 13844 8248 13900
rect 8184 13840 8248 13844
rect 8264 13900 8328 13904
rect 8264 13844 8268 13900
rect 8268 13844 8324 13900
rect 8324 13844 8328 13900
rect 8264 13840 8328 13844
rect 8344 13900 8408 13904
rect 8344 13844 8348 13900
rect 8348 13844 8404 13900
rect 8404 13844 8408 13900
rect 8344 13840 8408 13844
rect 8424 13900 8488 13904
rect 8424 13844 8428 13900
rect 8428 13844 8484 13900
rect 8484 13844 8488 13900
rect 8424 13840 8488 13844
rect 8504 13900 8568 13904
rect 8504 13844 8508 13900
rect 8508 13844 8564 13900
rect 8564 13844 8568 13900
rect 8504 13840 8568 13844
rect 8584 13900 8648 13904
rect 8584 13844 8588 13900
rect 8588 13844 8644 13900
rect 8644 13844 8648 13900
rect 8584 13840 8648 13844
rect 8664 13900 8728 13904
rect 8664 13844 8668 13900
rect 8668 13844 8724 13900
rect 8724 13844 8728 13900
rect 8664 13840 8728 13844
rect 8744 13900 8808 13904
rect 8744 13844 8748 13900
rect 8748 13844 8804 13900
rect 8804 13844 8808 13900
rect 8744 13840 8808 13844
rect 5802 13356 5866 13360
rect 5802 13300 5806 13356
rect 5806 13300 5862 13356
rect 5862 13300 5866 13356
rect 5802 13296 5866 13300
rect 5882 13356 5946 13360
rect 5882 13300 5886 13356
rect 5886 13300 5942 13356
rect 5942 13300 5946 13356
rect 5882 13296 5946 13300
rect 5962 13356 6026 13360
rect 5962 13300 5966 13356
rect 5966 13300 6022 13356
rect 6022 13300 6026 13356
rect 5962 13296 6026 13300
rect 6042 13356 6106 13360
rect 6042 13300 6046 13356
rect 6046 13300 6102 13356
rect 6102 13300 6106 13356
rect 6042 13296 6106 13300
rect 8184 12812 8248 12816
rect 8184 12756 8188 12812
rect 8188 12756 8244 12812
rect 8244 12756 8248 12812
rect 8184 12752 8248 12756
rect 8264 12812 8328 12816
rect 8264 12756 8268 12812
rect 8268 12756 8324 12812
rect 8324 12756 8328 12812
rect 8264 12752 8328 12756
rect 8344 12812 8408 12816
rect 8344 12756 8348 12812
rect 8348 12756 8404 12812
rect 8404 12756 8408 12812
rect 8344 12752 8408 12756
rect 8424 12812 8488 12816
rect 8424 12756 8428 12812
rect 8428 12756 8484 12812
rect 8484 12756 8488 12812
rect 8424 12752 8488 12756
rect 8504 12812 8568 12816
rect 8504 12756 8508 12812
rect 8508 12756 8564 12812
rect 8564 12756 8568 12812
rect 8504 12752 8568 12756
rect 8584 12812 8648 12816
rect 8584 12756 8588 12812
rect 8588 12756 8644 12812
rect 8644 12756 8648 12812
rect 8584 12752 8648 12756
rect 8664 12812 8728 12816
rect 8664 12756 8668 12812
rect 8668 12756 8724 12812
rect 8724 12756 8728 12812
rect 8664 12752 8728 12756
rect 8744 12812 8808 12816
rect 8744 12756 8748 12812
rect 8748 12756 8804 12812
rect 8804 12756 8808 12812
rect 8744 12752 8808 12756
rect 5802 12268 5866 12272
rect 5802 12212 5806 12268
rect 5806 12212 5862 12268
rect 5862 12212 5866 12268
rect 5802 12208 5866 12212
rect 5882 12268 5946 12272
rect 5882 12212 5886 12268
rect 5886 12212 5942 12268
rect 5942 12212 5946 12268
rect 5882 12208 5946 12212
rect 5962 12268 6026 12272
rect 5962 12212 5966 12268
rect 5966 12212 6022 12268
rect 6022 12212 6026 12268
rect 5962 12208 6026 12212
rect 6042 12268 6106 12272
rect 6042 12212 6046 12268
rect 6046 12212 6102 12268
rect 6102 12212 6106 12268
rect 6042 12208 6106 12212
rect 7880 12180 7944 12244
rect 8184 11724 8248 11728
rect 8184 11668 8188 11724
rect 8188 11668 8244 11724
rect 8244 11668 8248 11724
rect 8184 11664 8248 11668
rect 8264 11724 8328 11728
rect 8264 11668 8268 11724
rect 8268 11668 8324 11724
rect 8324 11668 8328 11724
rect 8264 11664 8328 11668
rect 8344 11724 8408 11728
rect 8344 11668 8348 11724
rect 8348 11668 8404 11724
rect 8404 11668 8408 11724
rect 8344 11664 8408 11668
rect 8424 11724 8488 11728
rect 8424 11668 8428 11724
rect 8428 11668 8484 11724
rect 8484 11668 8488 11724
rect 8424 11664 8488 11668
rect 8504 11724 8568 11728
rect 8504 11668 8508 11724
rect 8508 11668 8564 11724
rect 8564 11668 8568 11724
rect 8504 11664 8568 11668
rect 8584 11724 8648 11728
rect 8584 11668 8588 11724
rect 8588 11668 8644 11724
rect 8644 11668 8648 11724
rect 8584 11664 8648 11668
rect 8664 11724 8728 11728
rect 8664 11668 8668 11724
rect 8668 11668 8724 11724
rect 8724 11668 8728 11724
rect 8664 11664 8728 11668
rect 8744 11724 8808 11728
rect 8744 11668 8748 11724
rect 8748 11668 8804 11724
rect 8804 11668 8808 11724
rect 8744 11664 8808 11668
rect 7880 11326 7944 11390
rect 5802 11180 5866 11184
rect 5802 11124 5806 11180
rect 5806 11124 5862 11180
rect 5862 11124 5866 11180
rect 5802 11120 5866 11124
rect 5882 11180 5946 11184
rect 5882 11124 5886 11180
rect 5886 11124 5942 11180
rect 5942 11124 5946 11180
rect 5882 11120 5946 11124
rect 5962 11180 6026 11184
rect 5962 11124 5966 11180
rect 5966 11124 6022 11180
rect 6022 11124 6026 11180
rect 5962 11120 6026 11124
rect 6042 11180 6106 11184
rect 6042 11124 6046 11180
rect 6046 11124 6102 11180
rect 6102 11124 6106 11180
rect 6042 11120 6106 11124
rect 8184 10636 8248 10640
rect 8184 10580 8188 10636
rect 8188 10580 8244 10636
rect 8244 10580 8248 10636
rect 8184 10576 8248 10580
rect 8264 10636 8328 10640
rect 8264 10580 8268 10636
rect 8268 10580 8324 10636
rect 8324 10580 8328 10636
rect 8264 10576 8328 10580
rect 8344 10636 8408 10640
rect 8344 10580 8348 10636
rect 8348 10580 8404 10636
rect 8404 10580 8408 10636
rect 8344 10576 8408 10580
rect 8424 10636 8488 10640
rect 8424 10580 8428 10636
rect 8428 10580 8484 10636
rect 8484 10580 8488 10636
rect 8424 10576 8488 10580
rect 8504 10636 8568 10640
rect 8504 10580 8508 10636
rect 8508 10580 8564 10636
rect 8564 10580 8568 10636
rect 8504 10576 8568 10580
rect 8584 10636 8648 10640
rect 8584 10580 8588 10636
rect 8588 10580 8644 10636
rect 8644 10580 8648 10636
rect 8584 10576 8648 10580
rect 8664 10636 8728 10640
rect 8664 10580 8668 10636
rect 8668 10580 8724 10636
rect 8724 10580 8728 10636
rect 8664 10576 8728 10580
rect 8744 10636 8808 10640
rect 8744 10580 8748 10636
rect 8748 10580 8804 10636
rect 8804 10580 8808 10636
rect 8744 10576 8808 10580
rect 7880 10228 7944 10292
rect 5802 10092 5866 10096
rect 5802 10036 5806 10092
rect 5806 10036 5862 10092
rect 5862 10036 5866 10092
rect 5802 10032 5866 10036
rect 5882 10092 5946 10096
rect 5882 10036 5886 10092
rect 5886 10036 5942 10092
rect 5942 10036 5946 10092
rect 5882 10032 5946 10036
rect 5962 10092 6026 10096
rect 5962 10036 5966 10092
rect 5966 10036 6022 10092
rect 6022 10036 6026 10092
rect 5962 10032 6026 10036
rect 6042 10092 6106 10096
rect 6042 10036 6046 10092
rect 6046 10036 6102 10092
rect 6102 10036 6106 10092
rect 6042 10032 6106 10036
rect 7880 9862 7944 9926
rect 8184 9548 8248 9552
rect 8184 9492 8188 9548
rect 8188 9492 8244 9548
rect 8244 9492 8248 9548
rect 8184 9488 8248 9492
rect 8264 9548 8328 9552
rect 8264 9492 8268 9548
rect 8268 9492 8324 9548
rect 8324 9492 8328 9548
rect 8264 9488 8328 9492
rect 8344 9548 8408 9552
rect 8344 9492 8348 9548
rect 8348 9492 8404 9548
rect 8404 9492 8408 9548
rect 8344 9488 8408 9492
rect 8424 9548 8488 9552
rect 8424 9492 8428 9548
rect 8428 9492 8484 9548
rect 8484 9492 8488 9548
rect 8424 9488 8488 9492
rect 8504 9548 8568 9552
rect 8504 9492 8508 9548
rect 8508 9492 8564 9548
rect 8564 9492 8568 9548
rect 8504 9488 8568 9492
rect 8584 9548 8648 9552
rect 8584 9492 8588 9548
rect 8588 9492 8644 9548
rect 8644 9492 8648 9548
rect 8584 9488 8648 9492
rect 8664 9548 8728 9552
rect 8664 9492 8668 9548
rect 8668 9492 8724 9548
rect 8724 9492 8728 9548
rect 8664 9488 8728 9492
rect 8744 9548 8808 9552
rect 8744 9492 8748 9548
rect 8748 9492 8804 9548
rect 8804 9492 8808 9548
rect 8744 9488 8808 9492
rect 5802 9004 5866 9008
rect 5802 8948 5806 9004
rect 5806 8948 5862 9004
rect 5862 8948 5866 9004
rect 5802 8944 5866 8948
rect 5882 9004 5946 9008
rect 5882 8948 5886 9004
rect 5886 8948 5942 9004
rect 5942 8948 5946 9004
rect 5882 8944 5946 8948
rect 5962 9004 6026 9008
rect 5962 8948 5966 9004
rect 5966 8948 6022 9004
rect 6022 8948 6026 9004
rect 5962 8944 6026 8948
rect 6042 9004 6106 9008
rect 6042 8948 6046 9004
rect 6046 8948 6102 9004
rect 6102 8948 6106 9004
rect 6042 8944 6106 8948
rect 8184 8460 8248 8464
rect 8184 8404 8188 8460
rect 8188 8404 8244 8460
rect 8244 8404 8248 8460
rect 8184 8400 8248 8404
rect 8264 8460 8328 8464
rect 8264 8404 8268 8460
rect 8268 8404 8324 8460
rect 8324 8404 8328 8460
rect 8264 8400 8328 8404
rect 8344 8460 8408 8464
rect 8344 8404 8348 8460
rect 8348 8404 8404 8460
rect 8404 8404 8408 8460
rect 8344 8400 8408 8404
rect 8424 8460 8488 8464
rect 8424 8404 8428 8460
rect 8428 8404 8484 8460
rect 8484 8404 8488 8460
rect 8424 8400 8488 8404
rect 8504 8460 8568 8464
rect 8504 8404 8508 8460
rect 8508 8404 8564 8460
rect 8564 8404 8568 8460
rect 8504 8400 8568 8404
rect 8584 8460 8648 8464
rect 8584 8404 8588 8460
rect 8588 8404 8644 8460
rect 8644 8404 8648 8460
rect 8584 8400 8648 8404
rect 8664 8460 8728 8464
rect 8664 8404 8668 8460
rect 8668 8404 8724 8460
rect 8724 8404 8728 8460
rect 8664 8400 8728 8404
rect 8744 8460 8808 8464
rect 8744 8404 8748 8460
rect 8748 8404 8804 8460
rect 8804 8404 8808 8460
rect 8744 8400 8808 8404
rect 5802 7916 5866 7920
rect 5802 7860 5806 7916
rect 5806 7860 5862 7916
rect 5862 7860 5866 7916
rect 5802 7856 5866 7860
rect 5882 7916 5946 7920
rect 5882 7860 5886 7916
rect 5886 7860 5942 7916
rect 5942 7860 5946 7916
rect 5882 7856 5946 7860
rect 5962 7916 6026 7920
rect 5962 7860 5966 7916
rect 5966 7860 6022 7916
rect 6022 7860 6026 7916
rect 5962 7856 6026 7860
rect 6042 7916 6106 7920
rect 6042 7860 6046 7916
rect 6046 7860 6102 7916
rect 6102 7860 6106 7916
rect 6042 7856 6106 7860
rect 8184 7372 8248 7376
rect 8184 7316 8188 7372
rect 8188 7316 8244 7372
rect 8244 7316 8248 7372
rect 8184 7312 8248 7316
rect 8264 7372 8328 7376
rect 8264 7316 8268 7372
rect 8268 7316 8324 7372
rect 8324 7316 8328 7372
rect 8264 7312 8328 7316
rect 8344 7372 8408 7376
rect 8344 7316 8348 7372
rect 8348 7316 8404 7372
rect 8404 7316 8408 7372
rect 8344 7312 8408 7316
rect 8424 7372 8488 7376
rect 8424 7316 8428 7372
rect 8428 7316 8484 7372
rect 8484 7316 8488 7372
rect 8424 7312 8488 7316
rect 8504 7372 8568 7376
rect 8504 7316 8508 7372
rect 8508 7316 8564 7372
rect 8564 7316 8568 7372
rect 8504 7312 8568 7316
rect 8584 7372 8648 7376
rect 8584 7316 8588 7372
rect 8588 7316 8644 7372
rect 8644 7316 8648 7372
rect 8584 7312 8648 7316
rect 8664 7372 8728 7376
rect 8664 7316 8668 7372
rect 8668 7316 8724 7372
rect 8724 7316 8728 7372
rect 8664 7312 8728 7316
rect 8744 7372 8808 7376
rect 8744 7316 8748 7372
rect 8748 7316 8804 7372
rect 8804 7316 8808 7372
rect 8744 7312 8808 7316
rect 5802 6828 5866 6832
rect 5802 6772 5806 6828
rect 5806 6772 5862 6828
rect 5862 6772 5866 6828
rect 5802 6768 5866 6772
rect 5882 6828 5946 6832
rect 5882 6772 5886 6828
rect 5886 6772 5942 6828
rect 5942 6772 5946 6828
rect 5882 6768 5946 6772
rect 5962 6828 6026 6832
rect 5962 6772 5966 6828
rect 5966 6772 6022 6828
rect 6022 6772 6026 6828
rect 5962 6768 6026 6772
rect 6042 6828 6106 6832
rect 6042 6772 6046 6828
rect 6046 6772 6102 6828
rect 6102 6772 6106 6828
rect 6042 6768 6106 6772
rect 8184 6284 8248 6288
rect 8184 6228 8188 6284
rect 8188 6228 8244 6284
rect 8244 6228 8248 6284
rect 8184 6224 8248 6228
rect 8264 6284 8328 6288
rect 8264 6228 8268 6284
rect 8268 6228 8324 6284
rect 8324 6228 8328 6284
rect 8264 6224 8328 6228
rect 8344 6284 8408 6288
rect 8344 6228 8348 6284
rect 8348 6228 8404 6284
rect 8404 6228 8408 6284
rect 8344 6224 8408 6228
rect 8424 6284 8488 6288
rect 8424 6228 8428 6284
rect 8428 6228 8484 6284
rect 8484 6228 8488 6284
rect 8424 6224 8488 6228
rect 8504 6284 8568 6288
rect 8504 6228 8508 6284
rect 8508 6228 8564 6284
rect 8564 6228 8568 6284
rect 8504 6224 8568 6228
rect 8584 6284 8648 6288
rect 8584 6228 8588 6284
rect 8588 6228 8644 6284
rect 8644 6228 8648 6284
rect 8584 6224 8648 6228
rect 8664 6284 8728 6288
rect 8664 6228 8668 6284
rect 8668 6228 8724 6284
rect 8724 6228 8728 6284
rect 8664 6224 8728 6228
rect 8744 6284 8808 6288
rect 8744 6228 8748 6284
rect 8748 6228 8804 6284
rect 8804 6228 8808 6284
rect 8744 6224 8808 6228
rect 5802 5740 5866 5744
rect 5802 5684 5806 5740
rect 5806 5684 5862 5740
rect 5862 5684 5866 5740
rect 5802 5680 5866 5684
rect 5882 5740 5946 5744
rect 5882 5684 5886 5740
rect 5886 5684 5942 5740
rect 5942 5684 5946 5740
rect 5882 5680 5946 5684
rect 5962 5740 6026 5744
rect 5962 5684 5966 5740
rect 5966 5684 6022 5740
rect 6022 5684 6026 5740
rect 5962 5680 6026 5684
rect 6042 5740 6106 5744
rect 6042 5684 6046 5740
rect 6046 5684 6102 5740
rect 6102 5684 6106 5740
rect 6042 5680 6106 5684
<< metal4 >>
rect 900 19254 2532 20128
rect 900 19018 958 19254
rect 1194 19018 1278 19254
rect 1514 19018 1598 19254
rect 1834 19018 1918 19254
rect 2154 19018 2238 19254
rect 2474 19018 2532 19254
rect 900 18934 2532 19018
rect 900 18698 958 18934
rect 1194 18698 1278 18934
rect 1514 18698 1598 18934
rect 1834 18698 1918 18934
rect 2154 18698 2238 18934
rect 2474 18698 2532 18934
rect 900 18614 2532 18698
rect 900 18378 958 18614
rect 1194 18378 1278 18614
rect 1514 18378 1598 18614
rect 1834 18378 1918 18614
rect 2154 18378 2238 18614
rect 2474 18378 2532 18614
rect 900 18294 2532 18378
rect 900 18058 958 18294
rect 1194 18058 1278 18294
rect 1514 18058 1598 18294
rect 1834 18058 1918 18294
rect 2154 18058 2238 18294
rect 2474 18058 2532 18294
rect 900 17974 2532 18058
rect 900 17738 958 17974
rect 1194 17738 1278 17974
rect 1514 17738 1598 17974
rect 1834 17738 1918 17974
rect 2154 17738 2238 17974
rect 2474 17738 2532 17974
rect 900 14214 2532 17738
rect 900 13978 958 14214
rect 1194 13978 1278 14214
rect 1514 13978 1598 14214
rect 1834 13978 1918 14214
rect 2154 13978 2238 14214
rect 2474 13978 2532 14214
rect 900 13894 2532 13978
rect 900 13658 958 13894
rect 1194 13658 1278 13894
rect 1514 13658 1598 13894
rect 1834 13658 1918 13894
rect 2154 13658 2238 13894
rect 2474 13658 2532 13894
rect 900 8774 2532 13658
rect 900 8538 958 8774
rect 1194 8538 1278 8774
rect 1514 8538 1598 8774
rect 1834 8538 1918 8774
rect 2154 8538 2238 8774
rect 2474 8538 2532 8774
rect 900 8454 2532 8538
rect 900 8218 958 8454
rect 1194 8218 1278 8454
rect 1514 8218 1598 8454
rect 1834 8218 1918 8454
rect 2154 8218 2238 8454
rect 2474 8218 2532 8454
rect 900 2390 2532 8218
rect 900 2154 958 2390
rect 1194 2154 1278 2390
rect 1514 2154 1598 2390
rect 1834 2154 1918 2390
rect 2154 2154 2238 2390
rect 2474 2154 2532 2390
rect 900 2070 2532 2154
rect 900 1834 958 2070
rect 1194 1834 1278 2070
rect 1514 1834 1598 2070
rect 1834 1834 1918 2070
rect 2154 1834 2238 2070
rect 2474 1834 2532 2070
rect 900 1750 2532 1834
rect 900 1514 958 1750
rect 1194 1514 1278 1750
rect 1514 1514 1598 1750
rect 1834 1514 1918 1750
rect 2154 1514 2238 1750
rect 2474 1514 2532 1750
rect 900 1430 2532 1514
rect 900 1194 958 1430
rect 1194 1194 1278 1430
rect 1514 1194 1598 1430
rect 1834 1194 1918 1430
rect 2154 1194 2238 1430
rect 2474 1194 2532 1430
rect 900 1110 2532 1194
rect 900 874 958 1110
rect 1194 874 1278 1110
rect 1514 874 1598 1110
rect 1834 874 1918 1110
rect 2154 874 2238 1110
rect 2474 874 2532 1110
rect 900 0 2532 874
rect 3348 16806 4980 20128
rect 3348 16570 3406 16806
rect 3642 16570 3726 16806
rect 3962 16570 4046 16806
rect 4282 16570 4366 16806
rect 4602 16570 4686 16806
rect 4922 16570 4980 16806
rect 3348 16486 4980 16570
rect 3348 16250 3406 16486
rect 3642 16250 3726 16486
rect 3962 16250 4046 16486
rect 4282 16250 4366 16486
rect 4602 16250 4686 16486
rect 4922 16250 4980 16486
rect 3348 16166 4980 16250
rect 3348 15930 3406 16166
rect 3642 15930 3726 16166
rect 3962 15930 4046 16166
rect 4282 15930 4366 16166
rect 4602 15930 4686 16166
rect 4922 15930 4980 16166
rect 3348 15846 4980 15930
rect 3348 15610 3406 15846
rect 3642 15610 3726 15846
rect 3962 15610 4046 15846
rect 4282 15610 4366 15846
rect 4602 15610 4686 15846
rect 4922 15610 4980 15846
rect 3348 15526 4980 15610
rect 3348 15290 3406 15526
rect 3642 15290 3726 15526
rect 3962 15290 4046 15526
rect 4282 15290 4366 15526
rect 4602 15290 4686 15526
rect 4922 15290 4980 15526
rect 3348 11494 4980 15290
rect 3348 11258 3406 11494
rect 3642 11258 3726 11494
rect 3962 11258 4046 11494
rect 4282 11258 4366 11494
rect 4602 11258 4686 11494
rect 4922 11258 4980 11494
rect 3348 11174 4980 11258
rect 3348 10938 3406 11174
rect 3642 10938 3726 11174
rect 3962 10938 4046 11174
rect 4282 10938 4366 11174
rect 4602 10938 4686 11174
rect 4922 10938 4980 11174
rect 3348 6054 4980 10938
rect 3348 5818 3406 6054
rect 3642 5818 3726 6054
rect 3962 5818 4046 6054
rect 4282 5818 4366 6054
rect 4602 5818 4686 6054
rect 4922 5818 4980 6054
rect 3348 5734 4980 5818
rect 3348 5498 3406 5734
rect 3642 5498 3726 5734
rect 3962 5498 4046 5734
rect 4282 5498 4366 5734
rect 4602 5498 4686 5734
rect 4922 5498 4980 5734
rect 3348 4838 4980 5498
rect 3348 4602 3406 4838
rect 3642 4602 3726 4838
rect 3962 4602 4046 4838
rect 4282 4602 4366 4838
rect 4602 4602 4686 4838
rect 4922 4602 4980 4838
rect 3348 4518 4980 4602
rect 3348 4282 3406 4518
rect 3642 4282 3726 4518
rect 3962 4282 4046 4518
rect 4282 4282 4366 4518
rect 4602 4282 4686 4518
rect 4922 4282 4980 4518
rect 3348 4198 4980 4282
rect 3348 3962 3406 4198
rect 3642 3962 3726 4198
rect 3962 3962 4046 4198
rect 4282 3962 4366 4198
rect 4602 3962 4686 4198
rect 4922 3962 4980 4198
rect 3348 3878 4980 3962
rect 3348 3642 3406 3878
rect 3642 3642 3726 3878
rect 3962 3642 4046 3878
rect 4282 3642 4366 3878
rect 4602 3642 4686 3878
rect 4922 3642 4980 3878
rect 3348 3558 4980 3642
rect 3348 3322 3406 3558
rect 3642 3322 3726 3558
rect 3962 3322 4046 3558
rect 4282 3322 4366 3558
rect 4602 3322 4686 3558
rect 4922 3322 4980 3558
rect 3348 0 4980 3322
rect 5440 19254 6112 19312
rect 5440 19018 5498 19254
rect 5734 19018 5818 19254
rect 6054 19018 6112 19254
rect 5440 18934 6112 19018
rect 5440 18698 5498 18934
rect 5734 18698 5818 18934
rect 6054 18698 6112 18934
rect 5440 18614 6112 18698
rect 5440 18378 5498 18614
rect 5734 18378 5818 18614
rect 6054 18378 6112 18614
rect 5440 18294 6112 18378
rect 5440 18058 5498 18294
rect 5734 18058 5818 18294
rect 6054 18058 6112 18294
rect 5440 17974 6112 18058
rect 5440 17738 5498 17974
rect 5734 17738 5818 17974
rect 6054 17738 6112 17974
rect 5440 14448 6112 17738
rect 5440 14384 5802 14448
rect 5866 14384 5882 14448
rect 5946 14384 5962 14448
rect 6026 14384 6042 14448
rect 6106 14384 6112 14448
rect 5440 14214 6112 14384
rect 5440 13978 5498 14214
rect 5734 13978 5818 14214
rect 6054 13978 6112 14214
rect 5440 13894 6112 13978
rect 5440 13658 5498 13894
rect 5734 13658 5818 13894
rect 6054 13658 6112 13894
rect 5440 13360 6112 13658
rect 5440 13296 5802 13360
rect 5866 13296 5882 13360
rect 5946 13296 5962 13360
rect 6026 13296 6042 13360
rect 6106 13296 6112 13360
rect 5440 12272 6112 13296
rect 5440 12208 5802 12272
rect 5866 12208 5882 12272
rect 5946 12208 5962 12272
rect 6026 12208 6042 12272
rect 6106 12208 6112 12272
rect 8160 16806 8832 16864
rect 8160 16570 8218 16806
rect 8454 16570 8538 16806
rect 8774 16570 8832 16806
rect 8160 16486 8832 16570
rect 8160 16250 8218 16486
rect 8454 16250 8538 16486
rect 8774 16250 8832 16486
rect 8160 16166 8832 16250
rect 8160 15930 8218 16166
rect 8454 15930 8538 16166
rect 8774 15930 8832 16166
rect 8160 15846 8832 15930
rect 8160 15610 8218 15846
rect 8454 15610 8538 15846
rect 8774 15610 8832 15846
rect 8160 15526 8832 15610
rect 8160 15290 8218 15526
rect 8454 15290 8538 15526
rect 8774 15290 8832 15526
rect 8160 13904 8832 15290
rect 8160 13840 8184 13904
rect 8248 13840 8264 13904
rect 8328 13840 8344 13904
rect 8408 13840 8424 13904
rect 8488 13840 8504 13904
rect 8568 13840 8584 13904
rect 8648 13840 8664 13904
rect 8728 13840 8744 13904
rect 8808 13840 8832 13904
rect 8160 12816 8832 13840
rect 8160 12752 8184 12816
rect 8248 12752 8264 12816
rect 8328 12752 8344 12816
rect 8408 12752 8424 12816
rect 8488 12752 8504 12816
rect 8568 12752 8584 12816
rect 8648 12752 8664 12816
rect 8728 12752 8744 12816
rect 8808 12752 8832 12816
rect 5440 11184 6112 12208
rect 7879 12244 7945 12245
rect 7879 12180 7880 12244
rect 7944 12180 7945 12244
rect 7879 12179 7945 12180
rect 7882 11391 7942 12179
rect 8160 11728 8832 12752
rect 8160 11664 8184 11728
rect 8248 11664 8264 11728
rect 8328 11664 8344 11728
rect 8408 11664 8424 11728
rect 8488 11664 8504 11728
rect 8568 11664 8584 11728
rect 8648 11664 8664 11728
rect 8728 11664 8744 11728
rect 8808 11664 8832 11728
rect 8160 11494 8832 11664
rect 7879 11390 7945 11391
rect 7879 11326 7880 11390
rect 7944 11326 7945 11390
rect 7879 11325 7945 11326
rect 5440 11120 5802 11184
rect 5866 11120 5882 11184
rect 5946 11120 5962 11184
rect 6026 11120 6042 11184
rect 6106 11120 6112 11184
rect 5440 10096 6112 11120
rect 7882 10293 7942 11325
rect 8160 11258 8218 11494
rect 8454 11258 8538 11494
rect 8774 11258 8832 11494
rect 8160 11174 8832 11258
rect 8160 10938 8218 11174
rect 8454 10938 8538 11174
rect 8774 10938 8832 11174
rect 8160 10640 8832 10938
rect 8160 10576 8184 10640
rect 8248 10576 8264 10640
rect 8328 10576 8344 10640
rect 8408 10576 8424 10640
rect 8488 10576 8504 10640
rect 8568 10576 8584 10640
rect 8648 10576 8664 10640
rect 8728 10576 8744 10640
rect 8808 10576 8832 10640
rect 7879 10292 7945 10293
rect 7879 10228 7880 10292
rect 7944 10228 7945 10292
rect 7879 10227 7945 10228
rect 5440 10032 5802 10096
rect 5866 10032 5882 10096
rect 5946 10032 5962 10096
rect 6026 10032 6042 10096
rect 6106 10032 6112 10096
rect 5440 9008 6112 10032
rect 7882 9927 7942 10227
rect 7879 9926 7945 9927
rect 7879 9862 7880 9926
rect 7944 9862 7945 9926
rect 7879 9861 7945 9862
rect 5440 8944 5802 9008
rect 5866 8944 5882 9008
rect 5946 8944 5962 9008
rect 6026 8944 6042 9008
rect 6106 8944 6112 9008
rect 5440 8774 6112 8944
rect 5440 8538 5498 8774
rect 5734 8538 5818 8774
rect 6054 8538 6112 8774
rect 5440 8454 6112 8538
rect 5440 8218 5498 8454
rect 5734 8218 5818 8454
rect 6054 8218 6112 8454
rect 5440 7920 6112 8218
rect 5440 7856 5802 7920
rect 5866 7856 5882 7920
rect 5946 7856 5962 7920
rect 6026 7856 6042 7920
rect 6106 7856 6112 7920
rect 5440 6832 6112 7856
rect 5440 6768 5802 6832
rect 5866 6768 5882 6832
rect 5946 6768 5962 6832
rect 6026 6768 6042 6832
rect 6106 6768 6112 6832
rect 5440 5744 6112 6768
rect 5440 5680 5802 5744
rect 5866 5680 5882 5744
rect 5946 5680 5962 5744
rect 6026 5680 6042 5744
rect 6106 5680 6112 5744
rect 5440 2390 6112 5680
rect 8160 9552 8832 10576
rect 8160 9488 8184 9552
rect 8248 9488 8264 9552
rect 8328 9488 8344 9552
rect 8408 9488 8424 9552
rect 8488 9488 8504 9552
rect 8568 9488 8584 9552
rect 8648 9488 8664 9552
rect 8728 9488 8744 9552
rect 8808 9488 8832 9552
rect 8160 8464 8832 9488
rect 8160 8400 8184 8464
rect 8248 8400 8264 8464
rect 8328 8400 8344 8464
rect 8408 8400 8424 8464
rect 8488 8400 8504 8464
rect 8568 8400 8584 8464
rect 8648 8400 8664 8464
rect 8728 8400 8744 8464
rect 8808 8400 8832 8464
rect 8160 7376 8832 8400
rect 8160 7312 8184 7376
rect 8248 7312 8264 7376
rect 8328 7312 8344 7376
rect 8408 7312 8424 7376
rect 8488 7312 8504 7376
rect 8568 7312 8584 7376
rect 8648 7312 8664 7376
rect 8728 7312 8744 7376
rect 8808 7312 8832 7376
rect 8160 6288 8832 7312
rect 8160 6224 8184 6288
rect 8248 6224 8264 6288
rect 8328 6224 8344 6288
rect 8408 6224 8424 6288
rect 8488 6224 8504 6288
rect 8568 6224 8584 6288
rect 8648 6224 8664 6288
rect 8728 6224 8744 6288
rect 8808 6224 8832 6288
rect 8160 6054 8832 6224
rect 8160 5818 8218 6054
rect 8454 5818 8538 6054
rect 8774 5818 8832 6054
rect 8160 5734 8832 5818
rect 8160 5498 8218 5734
rect 8454 5498 8538 5734
rect 8774 5498 8832 5734
rect 8160 4838 8832 5498
rect 8160 4602 8218 4838
rect 8454 4602 8538 4838
rect 8774 4602 8832 4838
rect 8160 4518 8832 4602
rect 8160 4282 8218 4518
rect 8454 4282 8538 4518
rect 8774 4282 8832 4518
rect 8160 4198 8832 4282
rect 8160 3962 8218 4198
rect 8454 3962 8538 4198
rect 8774 3962 8832 4198
rect 8160 3878 8832 3962
rect 8160 3642 8218 3878
rect 8454 3642 8538 3878
rect 8774 3642 8832 3878
rect 8160 3558 8832 3642
rect 8160 3322 8218 3558
rect 8454 3322 8538 3558
rect 8774 3322 8832 3558
rect 8160 3264 8832 3322
rect 11120 16806 12752 20128
rect 11120 16570 11178 16806
rect 11414 16570 11498 16806
rect 11734 16570 11818 16806
rect 12054 16570 12138 16806
rect 12374 16570 12458 16806
rect 12694 16570 12752 16806
rect 11120 16486 12752 16570
rect 11120 16250 11178 16486
rect 11414 16250 11498 16486
rect 11734 16250 11818 16486
rect 12054 16250 12138 16486
rect 12374 16250 12458 16486
rect 12694 16250 12752 16486
rect 11120 16166 12752 16250
rect 11120 15930 11178 16166
rect 11414 15930 11498 16166
rect 11734 15930 11818 16166
rect 12054 15930 12138 16166
rect 12374 15930 12458 16166
rect 12694 15930 12752 16166
rect 11120 15846 12752 15930
rect 11120 15610 11178 15846
rect 11414 15610 11498 15846
rect 11734 15610 11818 15846
rect 12054 15610 12138 15846
rect 12374 15610 12458 15846
rect 12694 15610 12752 15846
rect 11120 15526 12752 15610
rect 11120 15290 11178 15526
rect 11414 15290 11498 15526
rect 11734 15290 11818 15526
rect 12054 15290 12138 15526
rect 12374 15290 12458 15526
rect 12694 15290 12752 15526
rect 11120 11494 12752 15290
rect 11120 11258 11178 11494
rect 11414 11258 11498 11494
rect 11734 11258 11818 11494
rect 12054 11258 12138 11494
rect 12374 11258 12458 11494
rect 12694 11258 12752 11494
rect 11120 11174 12752 11258
rect 11120 10938 11178 11174
rect 11414 10938 11498 11174
rect 11734 10938 11818 11174
rect 12054 10938 12138 11174
rect 12374 10938 12458 11174
rect 12694 10938 12752 11174
rect 11120 6054 12752 10938
rect 11120 5818 11178 6054
rect 11414 5818 11498 6054
rect 11734 5818 11818 6054
rect 12054 5818 12138 6054
rect 12374 5818 12458 6054
rect 12694 5818 12752 6054
rect 11120 5734 12752 5818
rect 11120 5498 11178 5734
rect 11414 5498 11498 5734
rect 11734 5498 11818 5734
rect 12054 5498 12138 5734
rect 12374 5498 12458 5734
rect 12694 5498 12752 5734
rect 11120 4838 12752 5498
rect 11120 4602 11178 4838
rect 11414 4602 11498 4838
rect 11734 4602 11818 4838
rect 12054 4602 12138 4838
rect 12374 4602 12458 4838
rect 12694 4602 12752 4838
rect 11120 4518 12752 4602
rect 11120 4282 11178 4518
rect 11414 4282 11498 4518
rect 11734 4282 11818 4518
rect 12054 4282 12138 4518
rect 12374 4282 12458 4518
rect 12694 4282 12752 4518
rect 11120 4198 12752 4282
rect 11120 3962 11178 4198
rect 11414 3962 11498 4198
rect 11734 3962 11818 4198
rect 12054 3962 12138 4198
rect 12374 3962 12458 4198
rect 12694 3962 12752 4198
rect 11120 3878 12752 3962
rect 11120 3642 11178 3878
rect 11414 3642 11498 3878
rect 11734 3642 11818 3878
rect 12054 3642 12138 3878
rect 12374 3642 12458 3878
rect 12694 3642 12752 3878
rect 11120 3558 12752 3642
rect 11120 3322 11178 3558
rect 11414 3322 11498 3558
rect 11734 3322 11818 3558
rect 12054 3322 12138 3558
rect 12374 3322 12458 3558
rect 12694 3322 12752 3558
rect 5440 2154 5498 2390
rect 5734 2154 5818 2390
rect 6054 2154 6112 2390
rect 5440 2070 6112 2154
rect 5440 1834 5498 2070
rect 5734 1834 5818 2070
rect 6054 1834 6112 2070
rect 5440 1750 6112 1834
rect 5440 1514 5498 1750
rect 5734 1514 5818 1750
rect 6054 1514 6112 1750
rect 5440 1430 6112 1514
rect 5440 1194 5498 1430
rect 5734 1194 5818 1430
rect 6054 1194 6112 1430
rect 5440 1110 6112 1194
rect 5440 874 5498 1110
rect 5734 874 5818 1110
rect 6054 874 6112 1110
rect 5440 816 6112 874
rect 11120 0 12752 3322
rect 13568 19254 15200 20128
rect 13568 19018 13626 19254
rect 13862 19018 13946 19254
rect 14182 19018 14266 19254
rect 14502 19018 14586 19254
rect 14822 19018 14906 19254
rect 15142 19018 15200 19254
rect 13568 18934 15200 19018
rect 13568 18698 13626 18934
rect 13862 18698 13946 18934
rect 14182 18698 14266 18934
rect 14502 18698 14586 18934
rect 14822 18698 14906 18934
rect 15142 18698 15200 18934
rect 13568 18614 15200 18698
rect 13568 18378 13626 18614
rect 13862 18378 13946 18614
rect 14182 18378 14266 18614
rect 14502 18378 14586 18614
rect 14822 18378 14906 18614
rect 15142 18378 15200 18614
rect 13568 18294 15200 18378
rect 13568 18058 13626 18294
rect 13862 18058 13946 18294
rect 14182 18058 14266 18294
rect 14502 18058 14586 18294
rect 14822 18058 14906 18294
rect 15142 18058 15200 18294
rect 13568 17974 15200 18058
rect 13568 17738 13626 17974
rect 13862 17738 13946 17974
rect 14182 17738 14266 17974
rect 14502 17738 14586 17974
rect 14822 17738 14906 17974
rect 15142 17738 15200 17974
rect 13568 14214 15200 17738
rect 13568 13978 13626 14214
rect 13862 13978 13946 14214
rect 14182 13978 14266 14214
rect 14502 13978 14586 14214
rect 14822 13978 14906 14214
rect 15142 13978 15200 14214
rect 13568 13894 15200 13978
rect 13568 13658 13626 13894
rect 13862 13658 13946 13894
rect 14182 13658 14266 13894
rect 14502 13658 14586 13894
rect 14822 13658 14906 13894
rect 15142 13658 15200 13894
rect 13568 8774 15200 13658
rect 13568 8538 13626 8774
rect 13862 8538 13946 8774
rect 14182 8538 14266 8774
rect 14502 8538 14586 8774
rect 14822 8538 14906 8774
rect 15142 8538 15200 8774
rect 13568 8454 15200 8538
rect 13568 8218 13626 8454
rect 13862 8218 13946 8454
rect 14182 8218 14266 8454
rect 14502 8218 14586 8454
rect 14822 8218 14906 8454
rect 15142 8218 15200 8454
rect 13568 2390 15200 8218
rect 13568 2154 13626 2390
rect 13862 2154 13946 2390
rect 14182 2154 14266 2390
rect 14502 2154 14586 2390
rect 14822 2154 14906 2390
rect 15142 2154 15200 2390
rect 13568 2070 15200 2154
rect 13568 1834 13626 2070
rect 13862 1834 13946 2070
rect 14182 1834 14266 2070
rect 14502 1834 14586 2070
rect 14822 1834 14906 2070
rect 15142 1834 15200 2070
rect 13568 1750 15200 1834
rect 13568 1514 13626 1750
rect 13862 1514 13946 1750
rect 14182 1514 14266 1750
rect 14502 1514 14586 1750
rect 14822 1514 14906 1750
rect 15142 1514 15200 1750
rect 13568 1430 15200 1514
rect 13568 1194 13626 1430
rect 13862 1194 13946 1430
rect 14182 1194 14266 1430
rect 14502 1194 14586 1430
rect 14822 1194 14906 1430
rect 15142 1194 15200 1430
rect 13568 1110 15200 1194
rect 13568 874 13626 1110
rect 13862 874 13946 1110
rect 14182 874 14266 1110
rect 14502 874 14586 1110
rect 14822 874 14906 1110
rect 15142 874 15200 1110
rect 13568 0 15200 874
<< via4 >>
rect 958 19018 1194 19254
rect 1278 19018 1514 19254
rect 1598 19018 1834 19254
rect 1918 19018 2154 19254
rect 2238 19018 2474 19254
rect 958 18698 1194 18934
rect 1278 18698 1514 18934
rect 1598 18698 1834 18934
rect 1918 18698 2154 18934
rect 2238 18698 2474 18934
rect 958 18378 1194 18614
rect 1278 18378 1514 18614
rect 1598 18378 1834 18614
rect 1918 18378 2154 18614
rect 2238 18378 2474 18614
rect 958 18058 1194 18294
rect 1278 18058 1514 18294
rect 1598 18058 1834 18294
rect 1918 18058 2154 18294
rect 2238 18058 2474 18294
rect 958 17738 1194 17974
rect 1278 17738 1514 17974
rect 1598 17738 1834 17974
rect 1918 17738 2154 17974
rect 2238 17738 2474 17974
rect 958 13978 1194 14214
rect 1278 13978 1514 14214
rect 1598 13978 1834 14214
rect 1918 13978 2154 14214
rect 2238 13978 2474 14214
rect 958 13658 1194 13894
rect 1278 13658 1514 13894
rect 1598 13658 1834 13894
rect 1918 13658 2154 13894
rect 2238 13658 2474 13894
rect 958 8538 1194 8774
rect 1278 8538 1514 8774
rect 1598 8538 1834 8774
rect 1918 8538 2154 8774
rect 2238 8538 2474 8774
rect 958 8218 1194 8454
rect 1278 8218 1514 8454
rect 1598 8218 1834 8454
rect 1918 8218 2154 8454
rect 2238 8218 2474 8454
rect 958 2154 1194 2390
rect 1278 2154 1514 2390
rect 1598 2154 1834 2390
rect 1918 2154 2154 2390
rect 2238 2154 2474 2390
rect 958 1834 1194 2070
rect 1278 1834 1514 2070
rect 1598 1834 1834 2070
rect 1918 1834 2154 2070
rect 2238 1834 2474 2070
rect 958 1514 1194 1750
rect 1278 1514 1514 1750
rect 1598 1514 1834 1750
rect 1918 1514 2154 1750
rect 2238 1514 2474 1750
rect 958 1194 1194 1430
rect 1278 1194 1514 1430
rect 1598 1194 1834 1430
rect 1918 1194 2154 1430
rect 2238 1194 2474 1430
rect 958 874 1194 1110
rect 1278 874 1514 1110
rect 1598 874 1834 1110
rect 1918 874 2154 1110
rect 2238 874 2474 1110
rect 3406 16570 3642 16806
rect 3726 16570 3962 16806
rect 4046 16570 4282 16806
rect 4366 16570 4602 16806
rect 4686 16570 4922 16806
rect 3406 16250 3642 16486
rect 3726 16250 3962 16486
rect 4046 16250 4282 16486
rect 4366 16250 4602 16486
rect 4686 16250 4922 16486
rect 3406 15930 3642 16166
rect 3726 15930 3962 16166
rect 4046 15930 4282 16166
rect 4366 15930 4602 16166
rect 4686 15930 4922 16166
rect 3406 15610 3642 15846
rect 3726 15610 3962 15846
rect 4046 15610 4282 15846
rect 4366 15610 4602 15846
rect 4686 15610 4922 15846
rect 3406 15290 3642 15526
rect 3726 15290 3962 15526
rect 4046 15290 4282 15526
rect 4366 15290 4602 15526
rect 4686 15290 4922 15526
rect 3406 11258 3642 11494
rect 3726 11258 3962 11494
rect 4046 11258 4282 11494
rect 4366 11258 4602 11494
rect 4686 11258 4922 11494
rect 3406 10938 3642 11174
rect 3726 10938 3962 11174
rect 4046 10938 4282 11174
rect 4366 10938 4602 11174
rect 4686 10938 4922 11174
rect 3406 5818 3642 6054
rect 3726 5818 3962 6054
rect 4046 5818 4282 6054
rect 4366 5818 4602 6054
rect 4686 5818 4922 6054
rect 3406 5498 3642 5734
rect 3726 5498 3962 5734
rect 4046 5498 4282 5734
rect 4366 5498 4602 5734
rect 4686 5498 4922 5734
rect 3406 4602 3642 4838
rect 3726 4602 3962 4838
rect 4046 4602 4282 4838
rect 4366 4602 4602 4838
rect 4686 4602 4922 4838
rect 3406 4282 3642 4518
rect 3726 4282 3962 4518
rect 4046 4282 4282 4518
rect 4366 4282 4602 4518
rect 4686 4282 4922 4518
rect 3406 3962 3642 4198
rect 3726 3962 3962 4198
rect 4046 3962 4282 4198
rect 4366 3962 4602 4198
rect 4686 3962 4922 4198
rect 3406 3642 3642 3878
rect 3726 3642 3962 3878
rect 4046 3642 4282 3878
rect 4366 3642 4602 3878
rect 4686 3642 4922 3878
rect 3406 3322 3642 3558
rect 3726 3322 3962 3558
rect 4046 3322 4282 3558
rect 4366 3322 4602 3558
rect 4686 3322 4922 3558
rect 5498 19018 5734 19254
rect 5818 19018 6054 19254
rect 5498 18698 5734 18934
rect 5818 18698 6054 18934
rect 5498 18378 5734 18614
rect 5818 18378 6054 18614
rect 5498 18058 5734 18294
rect 5818 18058 6054 18294
rect 5498 17738 5734 17974
rect 5818 17738 6054 17974
rect 5498 13978 5734 14214
rect 5818 13978 6054 14214
rect 5498 13658 5734 13894
rect 5818 13658 6054 13894
rect 8218 16570 8454 16806
rect 8538 16570 8774 16806
rect 8218 16250 8454 16486
rect 8538 16250 8774 16486
rect 8218 15930 8454 16166
rect 8538 15930 8774 16166
rect 8218 15610 8454 15846
rect 8538 15610 8774 15846
rect 8218 15290 8454 15526
rect 8538 15290 8774 15526
rect 8218 11258 8454 11494
rect 8538 11258 8774 11494
rect 8218 10938 8454 11174
rect 8538 10938 8774 11174
rect 5498 8538 5734 8774
rect 5818 8538 6054 8774
rect 5498 8218 5734 8454
rect 5818 8218 6054 8454
rect 8218 5818 8454 6054
rect 8538 5818 8774 6054
rect 8218 5498 8454 5734
rect 8538 5498 8774 5734
rect 8218 4602 8454 4838
rect 8538 4602 8774 4838
rect 8218 4282 8454 4518
rect 8538 4282 8774 4518
rect 8218 3962 8454 4198
rect 8538 3962 8774 4198
rect 8218 3642 8454 3878
rect 8538 3642 8774 3878
rect 8218 3322 8454 3558
rect 8538 3322 8774 3558
rect 11178 16570 11414 16806
rect 11498 16570 11734 16806
rect 11818 16570 12054 16806
rect 12138 16570 12374 16806
rect 12458 16570 12694 16806
rect 11178 16250 11414 16486
rect 11498 16250 11734 16486
rect 11818 16250 12054 16486
rect 12138 16250 12374 16486
rect 12458 16250 12694 16486
rect 11178 15930 11414 16166
rect 11498 15930 11734 16166
rect 11818 15930 12054 16166
rect 12138 15930 12374 16166
rect 12458 15930 12694 16166
rect 11178 15610 11414 15846
rect 11498 15610 11734 15846
rect 11818 15610 12054 15846
rect 12138 15610 12374 15846
rect 12458 15610 12694 15846
rect 11178 15290 11414 15526
rect 11498 15290 11734 15526
rect 11818 15290 12054 15526
rect 12138 15290 12374 15526
rect 12458 15290 12694 15526
rect 11178 11258 11414 11494
rect 11498 11258 11734 11494
rect 11818 11258 12054 11494
rect 12138 11258 12374 11494
rect 12458 11258 12694 11494
rect 11178 10938 11414 11174
rect 11498 10938 11734 11174
rect 11818 10938 12054 11174
rect 12138 10938 12374 11174
rect 12458 10938 12694 11174
rect 11178 5818 11414 6054
rect 11498 5818 11734 6054
rect 11818 5818 12054 6054
rect 12138 5818 12374 6054
rect 12458 5818 12694 6054
rect 11178 5498 11414 5734
rect 11498 5498 11734 5734
rect 11818 5498 12054 5734
rect 12138 5498 12374 5734
rect 12458 5498 12694 5734
rect 11178 4602 11414 4838
rect 11498 4602 11734 4838
rect 11818 4602 12054 4838
rect 12138 4602 12374 4838
rect 12458 4602 12694 4838
rect 11178 4282 11414 4518
rect 11498 4282 11734 4518
rect 11818 4282 12054 4518
rect 12138 4282 12374 4518
rect 12458 4282 12694 4518
rect 11178 3962 11414 4198
rect 11498 3962 11734 4198
rect 11818 3962 12054 4198
rect 12138 3962 12374 4198
rect 12458 3962 12694 4198
rect 11178 3642 11414 3878
rect 11498 3642 11734 3878
rect 11818 3642 12054 3878
rect 12138 3642 12374 3878
rect 12458 3642 12694 3878
rect 11178 3322 11414 3558
rect 11498 3322 11734 3558
rect 11818 3322 12054 3558
rect 12138 3322 12374 3558
rect 12458 3322 12694 3558
rect 5498 2154 5734 2390
rect 5818 2154 6054 2390
rect 5498 1834 5734 2070
rect 5818 1834 6054 2070
rect 5498 1514 5734 1750
rect 5818 1514 6054 1750
rect 5498 1194 5734 1430
rect 5818 1194 6054 1430
rect 5498 874 5734 1110
rect 5818 874 6054 1110
rect 13626 19018 13862 19254
rect 13946 19018 14182 19254
rect 14266 19018 14502 19254
rect 14586 19018 14822 19254
rect 14906 19018 15142 19254
rect 13626 18698 13862 18934
rect 13946 18698 14182 18934
rect 14266 18698 14502 18934
rect 14586 18698 14822 18934
rect 14906 18698 15142 18934
rect 13626 18378 13862 18614
rect 13946 18378 14182 18614
rect 14266 18378 14502 18614
rect 14586 18378 14822 18614
rect 14906 18378 15142 18614
rect 13626 18058 13862 18294
rect 13946 18058 14182 18294
rect 14266 18058 14502 18294
rect 14586 18058 14822 18294
rect 14906 18058 15142 18294
rect 13626 17738 13862 17974
rect 13946 17738 14182 17974
rect 14266 17738 14502 17974
rect 14586 17738 14822 17974
rect 14906 17738 15142 17974
rect 13626 13978 13862 14214
rect 13946 13978 14182 14214
rect 14266 13978 14502 14214
rect 14586 13978 14822 14214
rect 14906 13978 15142 14214
rect 13626 13658 13862 13894
rect 13946 13658 14182 13894
rect 14266 13658 14502 13894
rect 14586 13658 14822 13894
rect 14906 13658 15142 13894
rect 13626 8538 13862 8774
rect 13946 8538 14182 8774
rect 14266 8538 14502 8774
rect 14586 8538 14822 8774
rect 14906 8538 15142 8774
rect 13626 8218 13862 8454
rect 13946 8218 14182 8454
rect 14266 8218 14502 8454
rect 14586 8218 14822 8454
rect 14906 8218 15142 8454
rect 13626 2154 13862 2390
rect 13946 2154 14182 2390
rect 14266 2154 14502 2390
rect 14586 2154 14822 2390
rect 14906 2154 15142 2390
rect 13626 1834 13862 2070
rect 13946 1834 14182 2070
rect 14266 1834 14502 2070
rect 14586 1834 14822 2070
rect 14906 1834 15142 2070
rect 13626 1514 13862 1750
rect 13946 1514 14182 1750
rect 14266 1514 14502 1750
rect 14586 1514 14822 1750
rect 14906 1514 15142 1750
rect 13626 1194 13862 1430
rect 13946 1194 14182 1430
rect 14266 1194 14502 1430
rect 14586 1194 14822 1430
rect 14906 1194 15142 1430
rect 13626 874 13862 1110
rect 13946 874 14182 1110
rect 14266 874 14502 1110
rect 14586 874 14822 1110
rect 14906 874 15142 1110
<< metal5 >>
rect 0 19254 16100 19312
rect 0 19018 958 19254
rect 1194 19018 1278 19254
rect 1514 19018 1598 19254
rect 1834 19018 1918 19254
rect 2154 19018 2238 19254
rect 2474 19018 5498 19254
rect 5734 19018 5818 19254
rect 6054 19018 13626 19254
rect 13862 19018 13946 19254
rect 14182 19018 14266 19254
rect 14502 19018 14586 19254
rect 14822 19018 14906 19254
rect 15142 19018 16100 19254
rect 0 18934 16100 19018
rect 0 18698 958 18934
rect 1194 18698 1278 18934
rect 1514 18698 1598 18934
rect 1834 18698 1918 18934
rect 2154 18698 2238 18934
rect 2474 18698 5498 18934
rect 5734 18698 5818 18934
rect 6054 18698 13626 18934
rect 13862 18698 13946 18934
rect 14182 18698 14266 18934
rect 14502 18698 14586 18934
rect 14822 18698 14906 18934
rect 15142 18698 16100 18934
rect 0 18614 16100 18698
rect 0 18378 958 18614
rect 1194 18378 1278 18614
rect 1514 18378 1598 18614
rect 1834 18378 1918 18614
rect 2154 18378 2238 18614
rect 2474 18378 5498 18614
rect 5734 18378 5818 18614
rect 6054 18378 13626 18614
rect 13862 18378 13946 18614
rect 14182 18378 14266 18614
rect 14502 18378 14586 18614
rect 14822 18378 14906 18614
rect 15142 18378 16100 18614
rect 0 18294 16100 18378
rect 0 18058 958 18294
rect 1194 18058 1278 18294
rect 1514 18058 1598 18294
rect 1834 18058 1918 18294
rect 2154 18058 2238 18294
rect 2474 18058 5498 18294
rect 5734 18058 5818 18294
rect 6054 18058 13626 18294
rect 13862 18058 13946 18294
rect 14182 18058 14266 18294
rect 14502 18058 14586 18294
rect 14822 18058 14906 18294
rect 15142 18058 16100 18294
rect 0 17974 16100 18058
rect 0 17738 958 17974
rect 1194 17738 1278 17974
rect 1514 17738 1598 17974
rect 1834 17738 1918 17974
rect 2154 17738 2238 17974
rect 2474 17738 5498 17974
rect 5734 17738 5818 17974
rect 6054 17738 13626 17974
rect 13862 17738 13946 17974
rect 14182 17738 14266 17974
rect 14502 17738 14586 17974
rect 14822 17738 14906 17974
rect 15142 17738 16100 17974
rect 0 17680 16100 17738
rect 0 16806 16100 16864
rect 0 16570 3406 16806
rect 3642 16570 3726 16806
rect 3962 16570 4046 16806
rect 4282 16570 4366 16806
rect 4602 16570 4686 16806
rect 4922 16570 8218 16806
rect 8454 16570 8538 16806
rect 8774 16570 11178 16806
rect 11414 16570 11498 16806
rect 11734 16570 11818 16806
rect 12054 16570 12138 16806
rect 12374 16570 12458 16806
rect 12694 16570 16100 16806
rect 0 16486 16100 16570
rect 0 16250 3406 16486
rect 3642 16250 3726 16486
rect 3962 16250 4046 16486
rect 4282 16250 4366 16486
rect 4602 16250 4686 16486
rect 4922 16250 8218 16486
rect 8454 16250 8538 16486
rect 8774 16250 11178 16486
rect 11414 16250 11498 16486
rect 11734 16250 11818 16486
rect 12054 16250 12138 16486
rect 12374 16250 12458 16486
rect 12694 16250 16100 16486
rect 0 16166 16100 16250
rect 0 15930 3406 16166
rect 3642 15930 3726 16166
rect 3962 15930 4046 16166
rect 4282 15930 4366 16166
rect 4602 15930 4686 16166
rect 4922 15930 8218 16166
rect 8454 15930 8538 16166
rect 8774 15930 11178 16166
rect 11414 15930 11498 16166
rect 11734 15930 11818 16166
rect 12054 15930 12138 16166
rect 12374 15930 12458 16166
rect 12694 15930 16100 16166
rect 0 15846 16100 15930
rect 0 15610 3406 15846
rect 3642 15610 3726 15846
rect 3962 15610 4046 15846
rect 4282 15610 4366 15846
rect 4602 15610 4686 15846
rect 4922 15610 8218 15846
rect 8454 15610 8538 15846
rect 8774 15610 11178 15846
rect 11414 15610 11498 15846
rect 11734 15610 11818 15846
rect 12054 15610 12138 15846
rect 12374 15610 12458 15846
rect 12694 15610 16100 15846
rect 0 15526 16100 15610
rect 0 15290 3406 15526
rect 3642 15290 3726 15526
rect 3962 15290 4046 15526
rect 4282 15290 4366 15526
rect 4602 15290 4686 15526
rect 4922 15290 8218 15526
rect 8454 15290 8538 15526
rect 8774 15290 11178 15526
rect 11414 15290 11498 15526
rect 11734 15290 11818 15526
rect 12054 15290 12138 15526
rect 12374 15290 12458 15526
rect 12694 15290 16100 15526
rect 0 15232 16100 15290
rect 900 14214 15200 14272
rect 900 13978 958 14214
rect 1194 13978 1278 14214
rect 1514 13978 1598 14214
rect 1834 13978 1918 14214
rect 2154 13978 2238 14214
rect 2474 13978 5498 14214
rect 5734 13978 5818 14214
rect 6054 13978 13626 14214
rect 13862 13978 13946 14214
rect 14182 13978 14266 14214
rect 14502 13978 14586 14214
rect 14822 13978 14906 14214
rect 15142 13978 15200 14214
rect 900 13894 15200 13978
rect 900 13658 958 13894
rect 1194 13658 1278 13894
rect 1514 13658 1598 13894
rect 1834 13658 1918 13894
rect 2154 13658 2238 13894
rect 2474 13658 5498 13894
rect 5734 13658 5818 13894
rect 6054 13658 13626 13894
rect 13862 13658 13946 13894
rect 14182 13658 14266 13894
rect 14502 13658 14586 13894
rect 14822 13658 14906 13894
rect 15142 13658 15200 13894
rect 900 13600 15200 13658
rect 3348 11494 12752 11552
rect 3348 11258 3406 11494
rect 3642 11258 3726 11494
rect 3962 11258 4046 11494
rect 4282 11258 4366 11494
rect 4602 11258 4686 11494
rect 4922 11258 8218 11494
rect 8454 11258 8538 11494
rect 8774 11258 11178 11494
rect 11414 11258 11498 11494
rect 11734 11258 11818 11494
rect 12054 11258 12138 11494
rect 12374 11258 12458 11494
rect 12694 11258 12752 11494
rect 3348 11174 12752 11258
rect 3348 10938 3406 11174
rect 3642 10938 3726 11174
rect 3962 10938 4046 11174
rect 4282 10938 4366 11174
rect 4602 10938 4686 11174
rect 4922 10938 8218 11174
rect 8454 10938 8538 11174
rect 8774 10938 11178 11174
rect 11414 10938 11498 11174
rect 11734 10938 11818 11174
rect 12054 10938 12138 11174
rect 12374 10938 12458 11174
rect 12694 10938 12752 11174
rect 3348 10880 12752 10938
rect 900 8774 15200 8832
rect 900 8538 958 8774
rect 1194 8538 1278 8774
rect 1514 8538 1598 8774
rect 1834 8538 1918 8774
rect 2154 8538 2238 8774
rect 2474 8538 5498 8774
rect 5734 8538 5818 8774
rect 6054 8538 13626 8774
rect 13862 8538 13946 8774
rect 14182 8538 14266 8774
rect 14502 8538 14586 8774
rect 14822 8538 14906 8774
rect 15142 8538 15200 8774
rect 900 8454 15200 8538
rect 900 8218 958 8454
rect 1194 8218 1278 8454
rect 1514 8218 1598 8454
rect 1834 8218 1918 8454
rect 2154 8218 2238 8454
rect 2474 8218 5498 8454
rect 5734 8218 5818 8454
rect 6054 8218 13626 8454
rect 13862 8218 13946 8454
rect 14182 8218 14266 8454
rect 14502 8218 14586 8454
rect 14822 8218 14906 8454
rect 15142 8218 15200 8454
rect 900 8160 15200 8218
rect 3348 6054 12752 6112
rect 3348 5818 3406 6054
rect 3642 5818 3726 6054
rect 3962 5818 4046 6054
rect 4282 5818 4366 6054
rect 4602 5818 4686 6054
rect 4922 5818 8218 6054
rect 8454 5818 8538 6054
rect 8774 5818 11178 6054
rect 11414 5818 11498 6054
rect 11734 5818 11818 6054
rect 12054 5818 12138 6054
rect 12374 5818 12458 6054
rect 12694 5818 12752 6054
rect 3348 5734 12752 5818
rect 3348 5498 3406 5734
rect 3642 5498 3726 5734
rect 3962 5498 4046 5734
rect 4282 5498 4366 5734
rect 4602 5498 4686 5734
rect 4922 5498 8218 5734
rect 8454 5498 8538 5734
rect 8774 5498 11178 5734
rect 11414 5498 11498 5734
rect 11734 5498 11818 5734
rect 12054 5498 12138 5734
rect 12374 5498 12458 5734
rect 12694 5498 12752 5734
rect 3348 5440 12752 5498
rect 0 4838 16100 4896
rect 0 4602 3406 4838
rect 3642 4602 3726 4838
rect 3962 4602 4046 4838
rect 4282 4602 4366 4838
rect 4602 4602 4686 4838
rect 4922 4602 8218 4838
rect 8454 4602 8538 4838
rect 8774 4602 11178 4838
rect 11414 4602 11498 4838
rect 11734 4602 11818 4838
rect 12054 4602 12138 4838
rect 12374 4602 12458 4838
rect 12694 4602 16100 4838
rect 0 4518 16100 4602
rect 0 4282 3406 4518
rect 3642 4282 3726 4518
rect 3962 4282 4046 4518
rect 4282 4282 4366 4518
rect 4602 4282 4686 4518
rect 4922 4282 8218 4518
rect 8454 4282 8538 4518
rect 8774 4282 11178 4518
rect 11414 4282 11498 4518
rect 11734 4282 11818 4518
rect 12054 4282 12138 4518
rect 12374 4282 12458 4518
rect 12694 4282 16100 4518
rect 0 4198 16100 4282
rect 0 3962 3406 4198
rect 3642 3962 3726 4198
rect 3962 3962 4046 4198
rect 4282 3962 4366 4198
rect 4602 3962 4686 4198
rect 4922 3962 8218 4198
rect 8454 3962 8538 4198
rect 8774 3962 11178 4198
rect 11414 3962 11498 4198
rect 11734 3962 11818 4198
rect 12054 3962 12138 4198
rect 12374 3962 12458 4198
rect 12694 3962 16100 4198
rect 0 3878 16100 3962
rect 0 3642 3406 3878
rect 3642 3642 3726 3878
rect 3962 3642 4046 3878
rect 4282 3642 4366 3878
rect 4602 3642 4686 3878
rect 4922 3642 8218 3878
rect 8454 3642 8538 3878
rect 8774 3642 11178 3878
rect 11414 3642 11498 3878
rect 11734 3642 11818 3878
rect 12054 3642 12138 3878
rect 12374 3642 12458 3878
rect 12694 3642 16100 3878
rect 0 3558 16100 3642
rect 0 3322 3406 3558
rect 3642 3322 3726 3558
rect 3962 3322 4046 3558
rect 4282 3322 4366 3558
rect 4602 3322 4686 3558
rect 4922 3322 8218 3558
rect 8454 3322 8538 3558
rect 8774 3322 11178 3558
rect 11414 3322 11498 3558
rect 11734 3322 11818 3558
rect 12054 3322 12138 3558
rect 12374 3322 12458 3558
rect 12694 3322 16100 3558
rect 0 3264 16100 3322
rect 0 2390 16100 2448
rect 0 2154 958 2390
rect 1194 2154 1278 2390
rect 1514 2154 1598 2390
rect 1834 2154 1918 2390
rect 2154 2154 2238 2390
rect 2474 2154 5498 2390
rect 5734 2154 5818 2390
rect 6054 2154 13626 2390
rect 13862 2154 13946 2390
rect 14182 2154 14266 2390
rect 14502 2154 14586 2390
rect 14822 2154 14906 2390
rect 15142 2154 16100 2390
rect 0 2070 16100 2154
rect 0 1834 958 2070
rect 1194 1834 1278 2070
rect 1514 1834 1598 2070
rect 1834 1834 1918 2070
rect 2154 1834 2238 2070
rect 2474 1834 5498 2070
rect 5734 1834 5818 2070
rect 6054 1834 13626 2070
rect 13862 1834 13946 2070
rect 14182 1834 14266 2070
rect 14502 1834 14586 2070
rect 14822 1834 14906 2070
rect 15142 1834 16100 2070
rect 0 1750 16100 1834
rect 0 1514 958 1750
rect 1194 1514 1278 1750
rect 1514 1514 1598 1750
rect 1834 1514 1918 1750
rect 2154 1514 2238 1750
rect 2474 1514 5498 1750
rect 5734 1514 5818 1750
rect 6054 1514 13626 1750
rect 13862 1514 13946 1750
rect 14182 1514 14266 1750
rect 14502 1514 14586 1750
rect 14822 1514 14906 1750
rect 15142 1514 16100 1750
rect 0 1430 16100 1514
rect 0 1194 958 1430
rect 1194 1194 1278 1430
rect 1514 1194 1598 1430
rect 1834 1194 1918 1430
rect 2154 1194 2238 1430
rect 2474 1194 5498 1430
rect 5734 1194 5818 1430
rect 6054 1194 13626 1430
rect 13862 1194 13946 1430
rect 14182 1194 14266 1430
rect 14502 1194 14586 1430
rect 14822 1194 14906 1430
rect 15142 1194 16100 1430
rect 0 1110 16100 1194
rect 0 874 958 1110
rect 1194 874 1278 1110
rect 1514 874 1598 1110
rect 1834 874 1918 1110
rect 2154 874 2238 1110
rect 2474 874 5498 1110
rect 5734 874 5818 1110
rect 6054 874 13626 1110
rect 13862 874 13946 1110
rect 14182 874 14266 1110
rect 14502 874 14586 1110
rect 14822 874 14906 1110
rect 15142 874 16100 1110
rect 0 816 16100 874
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform 1 0 5796 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  U72 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform -1 0 6256 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  U70
timestamp 1625971452
transform -1 0 6164 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILL_36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform 1 0 6164 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_70 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform 1 0 5888 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_66
timestamp 1625971452
transform 1 0 5796 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  U80
timestamp 1625971452
transform -1 0 6624 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U96 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform -1 0 6716 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILL_69
timestamp 1625971452
transform 1 0 6256 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_65
timestamp 1625971452
transform 1 0 6348 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__and2_0  U11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform 1 0 6624 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__fill_4  FILL_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform 1 0 7176 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILL_11
timestamp 1625971452
transform 1 0 6716 0 -1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_2
timestamp 1625971452
transform 1 0 7084 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_5
timestamp 1625971452
transform 1 0 7084 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  dac_select_bits_reg_5_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform 1 0 7176 0 -1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_3
timestamp 1625971452
transform 1 0 8372 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform 1 0 8648 0 -1 6800
box -38 -48 774 592
use sky130_fd_sc_hd__and2_0  U15
timestamp 1625971452
transform -1 0 9108 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  U13
timestamp 1625971452
transform 1 0 7820 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  U98
timestamp 1625971452
transform 1 0 9108 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U97
timestamp 1625971452
transform -1 0 7820 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILL_37
timestamp 1625971452
transform 1 0 8464 0 1 5712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_68
timestamp 1625971452
transform 1 0 8280 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_64
timestamp 1625971452
transform 1 0 9568 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_35
timestamp 1625971452
transform 1 0 9384 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  U71
timestamp 1625971452
transform -1 0 9660 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U69
timestamp 1625971452
transform 1 0 9752 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_1  U106 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform -1 0 10212 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_4
timestamp 1625971452
transform 1 0 9660 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_6
timestamp 1625971452
transform 1 0 9660 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_67
timestamp 1625971452
transform 1 0 10212 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_63
timestamp 1625971452
transform 1 0 10212 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_34
timestamp 1625971452
transform 1 0 10028 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_7
timestamp 1625971452
transform 1 0 5796 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  dac_select_bits_reg_4_
timestamp 1625971452
transform 1 0 6900 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_0  U9
timestamp 1625971452
transform 1 0 6440 0 1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  U95
timestamp 1625971452
transform -1 0 6440 0 1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U94
timestamp 1625971452
transform -1 0 6164 0 1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_8
timestamp 1625971452
transform 1 0 8372 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  dac_mask_reg_4_
timestamp 1625971452
transform -1 0 9936 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_9
timestamp 1625971452
transform 1 0 10212 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_33
timestamp 1625971452
transform 1 0 9936 0 1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_62
timestamp 1625971452
transform 1 0 10120 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_10
timestamp 1625971452
transform 1 0 7084 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__nor2b_1  U108
timestamp 1625971452
transform 1 0 6164 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  dac_select_bits_reg_3_
timestamp 1625971452
transform 1 0 7176 0 -1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_0  U7
timestamp 1625971452
transform 1 0 6624 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  U73
timestamp 1625971452
transform -1 0 6164 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILL_61
timestamp 1625971452
transform 1 0 5796 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__nor2b_1  U105
timestamp 1625971452
transform 1 0 9200 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__fill_4  FILL_10
timestamp 1625971452
transform 1 0 8648 0 -1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_32
timestamp 1625971452
transform 1 0 9016 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_11
timestamp 1625971452
transform 1 0 9660 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__and2_0  U10
timestamp 1625971452
transform 1 0 9752 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILL_60
timestamp 1625971452
transform 1 0 10212 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_12
timestamp 1625971452
transform 1 0 5796 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  dac_mask_reg_3_
timestamp 1625971452
transform -1 0 7360 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_0  U8
timestamp 1625971452
transform -1 0 7820 0 1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_13
timestamp 1625971452
transform 1 0 8372 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  dac_select_bits_reg_6_
timestamp 1625971452
transform 1 0 8464 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_1  U81
timestamp 1625971452
transform 1 0 7820 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILL_31
timestamp 1625971452
transform 1 0 8096 0 1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_59
timestamp 1625971452
transform 1 0 8280 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_14
timestamp 1625971452
transform 1 0 10212 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  U79
timestamp 1625971452
transform 1 0 9936 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_15
timestamp 1625971452
transform 1 0 7084 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  dac_mask_reg_6_
timestamp 1625971452
transform 1 0 7176 0 -1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_0  U6
timestamp 1625971452
transform 1 0 6440 0 -1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  U82
timestamp 1625971452
transform -1 0 6440 0 -1 8976
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  U74
timestamp 1625971452
transform 1 0 5888 0 -1 8976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILL_30
timestamp 1625971452
transform 1 0 6900 0 -1 8976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_58
timestamp 1625971452
transform 1 0 5796 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__nor2b_1  U104
timestamp 1625971452
transform -1 0 9660 0 -1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__fill_4  FILL_9
timestamp 1625971452
transform 1 0 8648 0 -1 8976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_29
timestamp 1625971452
transform 1 0 9016 0 -1 8976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_16
timestamp 1625971452
transform 1 0 9660 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__and2_0  U12
timestamp 1625971452
transform -1 0 10212 0 -1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILL_57
timestamp 1625971452
transform 1 0 10212 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_17
timestamp 1625971452
transform 1 0 5796 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_20
timestamp 1625971452
transform 1 0 7084 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_4  CTS_ccl_a_inv_00003 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform -1 0 6992 0 -1 10064
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  dac_mask_reg_2_
timestamp 1625971452
transform -1 0 7360 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  dac_select_bits_reg_0_
timestamp 1625971452
transform 1 0 7176 0 -1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_4  FILL_8
timestamp 1625971452
transform 1 0 5796 0 -1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__and2_0  U14
timestamp 1625971452
transform -1 0 7820 0 1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILL_27
timestamp 1625971452
transform 1 0 6164 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_54
timestamp 1625971452
transform 1 0 6992 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_18
timestamp 1625971452
transform 1 0 8372 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  clk_gate_dac_select_bits_reg_LTIE $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform -1 0 9200 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_1  U107
timestamp 1625971452
transform -1 0 8280 0 1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  dac_mask_reg_5_
timestamp 1625971452
transform 1 0 8556 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILL_26
timestamp 1625971452
transform 1 0 8648 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILL_25
timestamp 1625971452
transform 1 0 9200 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_56
timestamp 1625971452
transform 1 0 8280 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_55
timestamp 1625971452
transform 1 0 8464 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_53
timestamp 1625971452
transform 1 0 8832 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_19
timestamp 1625971452
transform 1 0 10212 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_21
timestamp 1625971452
transform 1 0 9660 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__and2_0  U21
timestamp 1625971452
transform -1 0 10212 0 -1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  U67
timestamp 1625971452
transform -1 0 9660 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILL_28
timestamp 1625971452
transform 1 0 10028 0 1 8976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_52
timestamp 1625971452
transform 1 0 10212 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_22
timestamp 1625971452
transform 1 0 5796 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  dac_select_bits_reg_7_
timestamp 1625971452
transform 1 0 6900 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_0  U16
timestamp 1625971452
transform 1 0 6164 0 1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  U91
timestamp 1625971452
transform -1 0 6164 0 1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U75
timestamp 1625971452
transform 1 0 6624 0 1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_23
timestamp 1625971452
transform 1 0 8372 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  dac_mask_reg_7_
timestamp 1625971452
transform 1 0 8464 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_24
timestamp 1625971452
transform 1 0 10212 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  U100
timestamp 1625971452
transform 1 0 9936 0 1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_25
timestamp 1625971452
transform 1 0 7084 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  CTS_ccl_a_inv_00006 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform -1 0 6624 0 -1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__sdlclkp_4  clk_gate_dac_select_bits_reg_latch $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform -1 0 8832 0 -1 11152
box -38 -48 1694 592
use sky130_fd_sc_hd__nor2b_1  U109
timestamp 1625971452
transform -1 0 7084 0 -1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  U92
timestamp 1625971452
transform 1 0 5980 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILL_24
timestamp 1625971452
transform 1 0 5796 0 -1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILL_2
timestamp 1625971452
transform 1 0 8832 0 -1 11152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_26
timestamp 1625971452
transform 1 0 9660 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  U102 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform -1 0 10212 0 -1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILL_51
timestamp 1625971452
transform 1 0 9568 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_50
timestamp 1625971452
transform 1 0 9752 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_49
timestamp 1625971452
transform 1 0 10212 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_27
timestamp 1625971452
transform 1 0 5796 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  dac_select_bits_reg_2_
timestamp 1625971452
transform -1 0 7912 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_0  U3
timestamp 1625971452
transform 1 0 5980 0 1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILL_48
timestamp 1625971452
transform 1 0 5888 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_28
timestamp 1625971452
transform 1 0 8372 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  dac_mask_reg_0_
timestamp 1625971452
transform 1 0 8464 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_0  U17
timestamp 1625971452
transform 1 0 7912 0 1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_29
timestamp 1625971452
transform 1 0 10212 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  U83
timestamp 1625971452
transform -1 0 10212 0 1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_30
timestamp 1625971452
transform 1 0 7084 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_1
timestamp 1625971452
transform 1 0 7452 0 -1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__and2_0  U5
timestamp 1625971452
transform 1 0 6348 0 -1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  U4
timestamp 1625971452
transform 1 0 5888 0 -1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  U103
timestamp 1625971452
transform 1 0 7176 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U93
timestamp 1625971452
transform -1 0 7084 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILL_47
timestamp 1625971452
transform 1 0 5796 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  dac_select_bits_reg_1_
timestamp 1625971452
transform 1 0 8188 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  U90 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform -1 0 10028 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_31
timestamp 1625971452
transform 1 0 9660 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_23
timestamp 1625971452
transform 1 0 10028 0 -1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_46
timestamp 1625971452
transform 1 0 10212 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_32
timestamp 1625971452
transform 1 0 5796 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__nor2b_1  U110
timestamp 1625971452
transform 1 0 7452 0 1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  dac_mask_reg_1_
timestamp 1625971452
transform 1 0 5980 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILL_45
timestamp 1625971452
transform 1 0 5888 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_33
timestamp 1625971452
transform 1 0 8372 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  state_r_reg_0_
timestamp 1625971452
transform 1 0 8740 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_0  U22
timestamp 1625971452
transform 1 0 7912 0 1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILL_22
timestamp 1625971452
transform 1 0 8464 0 1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_44
timestamp 1625971452
transform 1 0 8648 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_34
timestamp 1625971452
transform 1 0 10212 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_43
timestamp 1625971452
transform 1 0 5980 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_21
timestamp 1625971452
transform 1 0 5796 0 -1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILL_19
timestamp 1625971452
transform 1 0 6256 0 1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_1  U78
timestamp 1625971452
transform -1 0 6716 0 1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  U76
timestamp 1625971452
transform -1 0 6348 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__fill_4  FILL_7
timestamp 1625971452
transform 1 0 6348 0 -1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILL_6
timestamp 1625971452
transform 1 0 5888 0 1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_37
timestamp 1625971452
transform 1 0 5796 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_42
timestamp 1625971452
transform 1 0 6992 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_18
timestamp 1625971452
transform 1 0 6716 0 1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  U77
timestamp 1625971452
transform 1 0 6716 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_35
timestamp 1625971452
transform 1 0 7084 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  run_adc_n_reg
timestamp 1625971452
transform -1 0 8648 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  state_r_reg_1_
timestamp 1625971452
transform -1 0 8372 0 1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_38
timestamp 1625971452
transform 1 0 8372 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  out_valid_reg
timestamp 1625971452
transform 1 0 8740 0 1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2b_1  U18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform -1 0 9200 0 -1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  U19
timestamp 1625971452
transform -1 0 9660 0 -1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  U86
timestamp 1625971452
transform 1 0 8464 0 1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILL_41
timestamp 1625971452
transform 1 0 8648 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_36
timestamp 1625971452
transform 1 0 9660 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_39
timestamp 1625971452
transform 1 0 10212 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_1  U101 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform 1 0 9752 0 -1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_20
timestamp 1625971452
transform 1 0 10120 0 -1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  U88
timestamp 1625971452
transform -1 0 6716 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_40
timestamp 1625971452
transform 1 0 5796 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_41
timestamp 1625971452
transform 1 0 7084 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILL_5
timestamp 1625971452
transform 1 0 6716 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILL_4
timestamp 1625971452
transform 1 0 7176 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  U68
timestamp 1625971452
transform -1 0 6256 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILL_17
timestamp 1625971452
transform 1 0 6256 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_40
timestamp 1625971452
transform 1 0 5888 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  U85
timestamp 1625971452
transform -1 0 8924 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_42
timestamp 1625971452
transform 1 0 8372 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__and2_0  U20
timestamp 1625971452
transform 1 0 7544 0 -1 14416
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  U84
timestamp 1625971452
transform 1 0 9200 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  U89 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1625971452
transform -1 0 8372 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_16
timestamp 1625971452
transform 1 0 8464 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILL_15
timestamp 1625971452
transform 1 0 8924 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_39
timestamp 1625971452
transform 1 0 9108 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_43
timestamp 1625971452
transform 1 0 9660 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  U99
timestamp 1625971452
transform 1 0 9936 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILL_14
timestamp 1625971452
transform 1 0 9476 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILL_13
timestamp 1625971452
transform 1 0 9752 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_38
timestamp 1625971452
transform 1 0 10212 0 -1 14416
box -38 -48 130 592
<< labels >>
rlabel metal2 s 216 20031 244 20128 6 clk
port 0 nsew signal input
rlabel metal2 s 8036 20031 8064 20128 6 rst_n
port 1 nsew signal input
rlabel metal2 s 15856 20031 15884 20128 6 adc_start
port 2 nsew signal input
rlabel metal2 s 0 20080 97 20108 6 comparator_val
port 3 nsew signal input
rlabel metal2 s 0 20 97 48 6 run_adc_n
port 4 nsew signal tristate
rlabel metal2 s 0 2196 97 2224 6 adc_val[7]
port 5 nsew signal tristate
rlabel metal2 s 0 4440 97 4468 6 adc_val[6]
port 6 nsew signal tristate
rlabel metal2 s 0 6684 97 6712 6 adc_val[5]
port 7 nsew signal tristate
rlabel metal2 s 0 8928 97 8956 6 adc_val[4]
port 8 nsew signal tristate
rlabel metal2 s 0 11104 97 11132 6 adc_val[3]
port 9 nsew signal tristate
rlabel metal2 s 0 13348 97 13376 6 adc_val[2]
port 10 nsew signal tristate
rlabel metal2 s 0 15592 97 15620 6 adc_val[1]
port 11 nsew signal tristate
rlabel metal2 s 0 17836 97 17864 6 adc_val[0]
port 12 nsew signal tristate
rlabel metal2 s 16003 20080 16100 20108 6 out_valid
port 13 nsew signal tristate
rlabel metal5 s 14468 17680 16100 19312 6 VSS
port 14 nsew ground bidirectional
rlabel metal5 s 0 17680 1632 19312 6 VSS
port 15 nsew ground bidirectional
rlabel metal5 s 14468 816 16100 2448 6 VSS
port 16 nsew ground bidirectional
rlabel metal5 s 0 816 1632 2448 6 VSS
port 17 nsew ground bidirectional
rlabel metal4 s 13568 18496 15200 20128 6 VSS
port 18 nsew ground bidirectional
rlabel metal4 s 13568 0 15200 1632 6 VSS
port 19 nsew ground bidirectional
rlabel metal4 s 900 18496 2532 20128 6 VSS
port 20 nsew ground bidirectional
rlabel metal4 s 900 0 2532 1632 6 VSS
port 21 nsew ground bidirectional
rlabel metal5 s 14468 15232 16100 16864 6 VDD
port 22 nsew power bidirectional
rlabel metal5 s 0 15232 1632 16864 6 VDD
port 23 nsew power bidirectional
rlabel metal5 s 14468 3264 16100 4896 6 VDD
port 24 nsew power bidirectional
rlabel metal5 s 0 3264 1632 4896 6 VDD
port 25 nsew power bidirectional
rlabel metal4 s 11120 18496 12752 20128 6 VDD
port 26 nsew power bidirectional
rlabel metal4 s 11120 0 12752 1632 6 VDD
port 27 nsew power bidirectional
rlabel metal4 s 3348 18496 4980 20128 6 VDD
port 28 nsew power bidirectional
rlabel metal4 s 3348 0 4980 1632 6 VDD
port 29 nsew power bidirectional
<< end >>
