magic
tech sky130A
timestamp 1626486988
<< checkpaint >>
rect -798 -654 798 654
<< metal2 >>
rect -168 14 168 24
rect -168 -14 -154 14
rect -126 -14 -114 14
rect -86 -14 -74 14
rect -46 -14 -34 14
rect -6 -14 6 14
rect 34 -14 46 14
rect 74 -14 86 14
rect 114 -14 126 14
rect 154 -14 168 14
rect -168 -24 168 -14
<< via2 >>
rect -154 -14 -126 14
rect -114 -14 -86 14
rect -74 -14 -46 14
rect -34 -14 -6 14
rect 6 -14 34 14
rect 46 -14 74 14
rect 86 -14 114 14
rect 126 -14 154 14
<< metal3 >>
rect -168 14 168 24
rect -168 -14 -154 14
rect -126 -14 -114 14
rect -86 -14 -74 14
rect -46 -14 -34 14
rect -6 -14 6 14
rect 34 -14 46 14
rect 74 -14 86 14
rect 114 -14 126 14
rect 154 -14 168 14
rect -168 -24 168 -14
<< end >>
