magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< nwell >>
rect 342 -8918 24858 1758
<< pwell >>
rect -12358 -27258 24958 -11142
<< nmos >>
rect 2628 -12318 3588 -11718
rect 3646 -12318 4606 -11718
rect 4664 -12318 5624 -11718
rect 5682 -12318 6642 -11718
rect 6700 -12318 7660 -11718
rect 7718 -12318 8678 -11718
rect 8736 -12318 9696 -11718
rect 9754 -12318 10714 -11718
rect 10772 -12318 11732 -11718
rect 11790 -12318 12750 -11718
rect 12808 -12318 13768 -11718
rect 13826 -12318 14786 -11718
rect 14844 -12318 15804 -11718
rect 15862 -12318 16822 -11718
rect 16880 -12318 17840 -11718
rect 17898 -12318 18858 -11718
rect 18916 -12318 19876 -11718
rect 19934 -12318 20894 -11718
rect 20952 -12318 21912 -11718
rect 21970 -12318 22930 -11718
rect 2628 -13552 3588 -12952
rect 3646 -13552 4606 -12952
rect 4664 -13552 5624 -12952
rect 5682 -13552 6642 -12952
rect 6700 -13552 7660 -12952
rect 7718 -13552 8678 -12952
rect 8736 -13552 9696 -12952
rect 9754 -13552 10714 -12952
rect 10772 -13552 11732 -12952
rect 11790 -13552 12750 -12952
rect 12808 -13552 13768 -12952
rect 13826 -13552 14786 -12952
rect 14844 -13552 15804 -12952
rect 15862 -13552 16822 -12952
rect 16880 -13552 17840 -12952
rect 17898 -13552 18858 -12952
rect 18916 -13552 19876 -12952
rect 19934 -13552 20894 -12952
rect 20952 -13552 21912 -12952
rect 21970 -13552 22930 -12952
rect 2628 -14784 3588 -14184
rect 3646 -14784 4606 -14184
rect 4664 -14784 5624 -14184
rect 5682 -14784 6642 -14184
rect 6700 -14784 7660 -14184
rect 7718 -14784 8678 -14184
rect 8736 -14784 9696 -14184
rect 9754 -14784 10714 -14184
rect 10772 -14784 11732 -14184
rect 11790 -14784 12750 -14184
rect 12808 -14784 13768 -14184
rect 13826 -14784 14786 -14184
rect 14844 -14784 15804 -14184
rect 15862 -14784 16822 -14184
rect 16880 -14784 17840 -14184
rect 17898 -14784 18858 -14184
rect 18916 -14784 19876 -14184
rect 19934 -14784 20894 -14184
rect 20952 -14784 21912 -14184
rect 21970 -14784 22930 -14184
rect 2626 -16018 3586 -15418
rect 3644 -16018 4604 -15418
rect 4662 -16018 5622 -15418
rect 5680 -16018 6640 -15418
rect 6698 -16018 7658 -15418
rect 7716 -16018 8676 -15418
rect 8734 -16018 9694 -15418
rect 9752 -16018 10712 -15418
rect 10770 -16018 11730 -15418
rect 11788 -16018 12748 -15418
rect 12806 -16018 13766 -15418
rect 13824 -16018 14784 -15418
rect 14842 -16018 15802 -15418
rect 15860 -16018 16820 -15418
rect 16878 -16018 17838 -15418
rect 17896 -16018 18856 -15418
rect 18914 -16018 19874 -15418
rect 19932 -16018 20892 -15418
rect 20950 -16018 21910 -15418
rect 21968 -16018 22928 -15418
rect 2626 -17252 3586 -16652
rect 3644 -17252 4604 -16652
rect 4662 -17252 5622 -16652
rect 5680 -17252 6640 -16652
rect 6698 -17252 7658 -16652
rect 7716 -17252 8676 -16652
rect 8734 -17252 9694 -16652
rect 9752 -17252 10712 -16652
rect 10770 -17252 11730 -16652
rect 11788 -17252 12748 -16652
rect 12806 -17252 13766 -16652
rect 13824 -17252 14784 -16652
rect 14842 -17252 15802 -16652
rect 15860 -17252 16820 -16652
rect 16878 -17252 17838 -16652
rect 17896 -17252 18856 -16652
rect 18914 -17252 19874 -16652
rect 19932 -17252 20892 -16652
rect 20950 -17252 21910 -16652
rect 21968 -17252 22928 -16652
rect 2626 -18484 3586 -17884
rect 3644 -18484 4604 -17884
rect 4662 -18484 5622 -17884
rect 5680 -18484 6640 -17884
rect 6698 -18484 7658 -17884
rect 7716 -18484 8676 -17884
rect 8734 -18484 9694 -17884
rect 9752 -18484 10712 -17884
rect 10770 -18484 11730 -17884
rect 11788 -18484 12748 -17884
rect 12806 -18484 13766 -17884
rect 13824 -18484 14784 -17884
rect 14842 -18484 15802 -17884
rect 15860 -18484 16820 -17884
rect 16878 -18484 17838 -17884
rect 17896 -18484 18856 -17884
rect 18914 -18484 19874 -17884
rect 19932 -18484 20892 -17884
rect 20950 -18484 21910 -17884
rect 21968 -18484 22928 -17884
rect 2626 -19718 3586 -19118
rect 3644 -19718 4604 -19118
rect 4662 -19718 5622 -19118
rect 5680 -19718 6640 -19118
rect 6698 -19718 7658 -19118
rect 7716 -19718 8676 -19118
rect 8734 -19718 9694 -19118
rect 9752 -19718 10712 -19118
rect 10770 -19718 11730 -19118
rect 11788 -19718 12748 -19118
rect 12806 -19718 13766 -19118
rect 13824 -19718 14784 -19118
rect 14842 -19718 15802 -19118
rect 15860 -19718 16820 -19118
rect 16878 -19718 17838 -19118
rect 17896 -19718 18856 -19118
rect 18914 -19718 19874 -19118
rect 19932 -19718 20892 -19118
rect 20950 -19718 21910 -19118
rect 21968 -19718 22928 -19118
rect 2626 -20952 3586 -20352
rect 3644 -20952 4604 -20352
rect 4662 -20952 5622 -20352
rect 5680 -20952 6640 -20352
rect 6698 -20952 7658 -20352
rect 7716 -20952 8676 -20352
rect 8734 -20952 9694 -20352
rect 9752 -20952 10712 -20352
rect 10770 -20952 11730 -20352
rect 11788 -20952 12748 -20352
rect 12806 -20952 13766 -20352
rect 13824 -20952 14784 -20352
rect 14842 -20952 15802 -20352
rect 15860 -20952 16820 -20352
rect 16878 -20952 17838 -20352
rect 17896 -20952 18856 -20352
rect 18914 -20952 19874 -20352
rect 19932 -20952 20892 -20352
rect 20950 -20952 21910 -20352
rect 21968 -20952 22928 -20352
rect -9359 -22381 -8399 -21781
rect -8341 -22381 -7381 -21781
rect -7323 -22381 -6363 -21781
rect -6305 -22381 -5345 -21781
rect -5287 -22381 -4327 -21781
rect -4269 -22381 -3309 -21781
rect 2626 -22184 3586 -21584
rect 3644 -22184 4604 -21584
rect 4662 -22184 5622 -21584
rect 5680 -22184 6640 -21584
rect 6698 -22184 7658 -21584
rect 7716 -22184 8676 -21584
rect 8734 -22184 9694 -21584
rect 9752 -22184 10712 -21584
rect 10770 -22184 11730 -21584
rect 11788 -22184 12748 -21584
rect 12806 -22184 13766 -21584
rect 13824 -22184 14784 -21584
rect 14842 -22184 15802 -21584
rect 15860 -22184 16820 -21584
rect 16878 -22184 17838 -21584
rect 17896 -22184 18856 -21584
rect 18914 -22184 19874 -21584
rect 19932 -22184 20892 -21584
rect 20950 -22184 21910 -21584
rect 21968 -22184 22928 -21584
rect -9360 -23494 -8400 -22894
rect -8342 -23494 -7382 -22894
rect -7324 -23494 -6364 -22894
rect -6306 -23494 -5346 -22894
rect -5288 -23494 -4328 -22894
rect -4270 -23494 -3310 -22894
rect 2626 -23418 3586 -22818
rect 3644 -23418 4604 -22818
rect 4662 -23418 5622 -22818
rect 5680 -23418 6640 -22818
rect 6698 -23418 7658 -22818
rect 7716 -23418 8676 -22818
rect 8734 -23418 9694 -22818
rect 9752 -23418 10712 -22818
rect 10770 -23418 11730 -22818
rect 11788 -23418 12748 -22818
rect 12806 -23418 13766 -22818
rect 13824 -23418 14784 -22818
rect 14842 -23418 15802 -22818
rect 15860 -23418 16820 -22818
rect 16878 -23418 17838 -22818
rect 17896 -23418 18856 -22818
rect 18914 -23418 19874 -22818
rect 19932 -23418 20892 -22818
rect 20950 -23418 21910 -22818
rect 21968 -23418 22928 -22818
rect -9359 -24605 -8399 -24005
rect -8341 -24605 -7381 -24005
rect -7323 -24605 -6363 -24005
rect -6305 -24605 -5345 -24005
rect -5287 -24605 -4327 -24005
rect -4269 -24605 -3309 -24005
rect 2626 -24652 3586 -24052
rect 3644 -24652 4604 -24052
rect 4662 -24652 5622 -24052
rect 5680 -24652 6640 -24052
rect 6698 -24652 7658 -24052
rect 7716 -24652 8676 -24052
rect 8734 -24652 9694 -24052
rect 9752 -24652 10712 -24052
rect 10770 -24652 11730 -24052
rect 11788 -24652 12748 -24052
rect 12806 -24652 13766 -24052
rect 13824 -24652 14784 -24052
rect 14842 -24652 15802 -24052
rect 15860 -24652 16820 -24052
rect 16878 -24652 17838 -24052
rect 17896 -24652 18856 -24052
rect 18914 -24652 19874 -24052
rect 19932 -24652 20892 -24052
rect 20950 -24652 21910 -24052
rect 21968 -24652 22928 -24052
rect -9360 -25718 -8400 -25118
rect -8342 -25718 -7382 -25118
rect -7324 -25718 -6364 -25118
rect -6306 -25718 -5346 -25118
rect -5288 -25718 -4328 -25118
rect -4270 -25718 -3310 -25118
rect 2626 -25884 3586 -25284
rect 3644 -25884 4604 -25284
rect 4662 -25884 5622 -25284
rect 5680 -25884 6640 -25284
rect 6698 -25884 7658 -25284
rect 7716 -25884 8676 -25284
rect 8734 -25884 9694 -25284
rect 9752 -25884 10712 -25284
rect 10770 -25884 11730 -25284
rect 11788 -25884 12748 -25284
rect 12806 -25884 13766 -25284
rect 13824 -25884 14784 -25284
rect 14842 -25884 15802 -25284
rect 15860 -25884 16820 -25284
rect 16878 -25884 17838 -25284
rect 17896 -25884 18856 -25284
rect 18914 -25884 19874 -25284
rect 19932 -25884 20892 -25284
rect 20950 -25884 21910 -25284
rect 21968 -25884 22928 -25284
<< pmos >>
rect 3672 -5090 3832 -4690
rect 3890 -5090 4050 -4690
rect 4108 -5090 4268 -4690
rect 4326 -5090 4486 -4690
rect 4544 -5090 4704 -4690
rect 4762 -5090 4922 -4690
rect 4980 -5090 5140 -4690
rect 5198 -5090 5358 -4690
rect 5416 -5090 5576 -4690
rect 5634 -5090 5794 -4690
rect 3672 -6028 3832 -5628
rect 3890 -6028 4050 -5628
rect 4108 -6028 4268 -5628
rect 4326 -6028 4486 -5628
rect 4544 -6028 4704 -5628
rect 4762 -6028 4922 -5628
rect 4980 -6028 5140 -5628
rect 5198 -6028 5358 -5628
rect 5416 -6028 5576 -5628
rect 5634 -6028 5794 -5628
rect 3672 -6966 3832 -6566
rect 3890 -6966 4050 -6566
rect 4108 -6966 4268 -6566
rect 4326 -6966 4486 -6566
rect 4544 -6966 4704 -6566
rect 4762 -6966 4922 -6566
rect 4980 -6966 5140 -6566
rect 5198 -6966 5358 -6566
rect 5416 -6966 5576 -6566
rect 5634 -6966 5794 -6566
rect 3672 -7904 3832 -7504
rect 3890 -7904 4050 -7504
rect 4108 -7904 4268 -7504
rect 4326 -7904 4486 -7504
rect 4544 -7904 4704 -7504
rect 4762 -7904 4922 -7504
rect 4980 -7904 5140 -7504
rect 5198 -7904 5358 -7504
rect 5416 -7904 5576 -7504
rect 5634 -7904 5794 -7504
<< nmoslvt >>
rect -9138 -13112 -8178 -12512
rect -8120 -13112 -7160 -12512
rect -7102 -13112 -6142 -12512
rect -6084 -13112 -5124 -12512
rect -5066 -13112 -4106 -12512
rect -4048 -13112 -3088 -12512
rect -3030 -13112 -2070 -12512
rect -2012 -13112 -1052 -12512
rect -994 -13112 -34 -12512
rect -9138 -13930 -8178 -13330
rect -8120 -13930 -7160 -13330
rect -7102 -13930 -6142 -13330
rect -6084 -13930 -5124 -13330
rect -5066 -13930 -4106 -13330
rect -4048 -13930 -3088 -13330
rect -3030 -13930 -2070 -13330
rect -2012 -13930 -1052 -13330
rect -994 -13930 -34 -13330
rect -9138 -14748 -8178 -14148
rect -8120 -14748 -7160 -14148
rect -7102 -14748 -6142 -14148
rect -6084 -14748 -5124 -14148
rect -5066 -14748 -4106 -14148
rect -4048 -14748 -3088 -14148
rect -3030 -14748 -2070 -14148
rect -2012 -14748 -1052 -14148
rect -994 -14748 -34 -14148
rect -9138 -15566 -8178 -14966
rect -8120 -15566 -7160 -14966
rect -7102 -15566 -6142 -14966
rect -6084 -15566 -5124 -14966
rect -5066 -15566 -4106 -14966
rect -4048 -15566 -3088 -14966
rect -3030 -15566 -2070 -14966
rect -2012 -15566 -1052 -14966
rect -994 -15566 -34 -14966
rect -9138 -16384 -8178 -15784
rect -8120 -16384 -7160 -15784
rect -7102 -16384 -6142 -15784
rect -6084 -16384 -5124 -15784
rect -5066 -16384 -4106 -15784
rect -4048 -16384 -3088 -15784
rect -3030 -16384 -2070 -15784
rect -2012 -16384 -1052 -15784
rect -994 -16384 -34 -15784
rect -9138 -17202 -8178 -16602
rect -8120 -17202 -7160 -16602
rect -7102 -17202 -6142 -16602
rect -6084 -17202 -5124 -16602
rect -5066 -17202 -4106 -16602
rect -4048 -17202 -3088 -16602
rect -3030 -17202 -2070 -16602
rect -2012 -17202 -1052 -16602
rect -994 -17202 -34 -16602
rect -9138 -18020 -8178 -17420
rect -8120 -18020 -7160 -17420
rect -7102 -18020 -6142 -17420
rect -6084 -18020 -5124 -17420
rect -5066 -18020 -4106 -17420
rect -4048 -18020 -3088 -17420
rect -3030 -18020 -2070 -17420
rect -2012 -18020 -1052 -17420
rect -994 -18020 -34 -17420
rect -9138 -18838 -8178 -18238
rect -8120 -18838 -7160 -18238
rect -7102 -18838 -6142 -18238
rect -6084 -18838 -5124 -18238
rect -5066 -18838 -4106 -18238
rect -4048 -18838 -3088 -18238
rect -3030 -18838 -2070 -18238
rect -2012 -18838 -1052 -18238
rect -994 -18838 -34 -18238
rect -2278 -19822 -2118 -19622
rect -2060 -19822 -1900 -19622
rect -1842 -19822 -1682 -19622
rect -1624 -19822 -1464 -19622
rect -1406 -19822 -1246 -19622
rect -1188 -19822 -1028 -19622
rect -970 -19822 -810 -19622
rect -752 -19822 -592 -19622
rect -534 -19822 -374 -19622
rect -316 -19822 -156 -19622
rect -2278 -20654 -2118 -20454
rect -2060 -20654 -1900 -20454
rect -1842 -20654 -1682 -20454
rect -1624 -20654 -1464 -20454
rect -1406 -20654 -1246 -20454
rect -1188 -20654 -1028 -20454
rect -970 -20654 -810 -20454
rect -752 -20654 -592 -20454
rect -534 -20654 -374 -20454
rect -316 -20654 -156 -20454
rect -2364 -22380 -2124 -21780
rect -2066 -22380 -1826 -21780
rect -1768 -22380 -1528 -21780
rect -1470 -22380 -1230 -21780
rect -1172 -22380 -932 -21780
rect -874 -22380 -634 -21780
rect -576 -22380 -336 -21780
rect -278 -22380 -38 -21780
rect 20 -22380 260 -21780
rect 318 -22380 558 -21780
rect 616 -22380 856 -21780
rect -2364 -23492 -2124 -22892
rect -2066 -23492 -1826 -22892
rect -1768 -23492 -1528 -22892
rect -1470 -23492 -1230 -22892
rect -1172 -23492 -932 -22892
rect -874 -23492 -634 -22892
rect -576 -23492 -336 -22892
rect -278 -23492 -38 -22892
rect 20 -23492 260 -22892
rect 318 -23492 558 -22892
rect 616 -23492 856 -22892
rect -2366 -24604 -2126 -24004
rect -2068 -24604 -1828 -24004
rect -1770 -24604 -1530 -24004
rect -1472 -24604 -1232 -24004
rect -1174 -24604 -934 -24004
rect -876 -24604 -636 -24004
rect -578 -24604 -338 -24004
rect -280 -24604 -40 -24004
rect 18 -24604 258 -24004
rect 316 -24604 556 -24004
rect 614 -24604 854 -24004
rect -2366 -25714 -2126 -25114
rect -2068 -25714 -1828 -25114
rect -1770 -25714 -1530 -25114
rect -1472 -25714 -1232 -25114
rect -1174 -25714 -934 -25114
rect -876 -25714 -636 -25114
rect -578 -25714 -338 -25114
rect -280 -25714 -40 -25114
rect 18 -25714 258 -25114
rect 316 -25714 556 -25114
rect 614 -25714 854 -25114
<< ndiff >>
rect 2570 -11730 2628 -11718
rect 2570 -12306 2582 -11730
rect 2616 -12306 2628 -11730
rect 2570 -12318 2628 -12306
rect 3588 -11730 3646 -11718
rect 3588 -12306 3600 -11730
rect 3634 -12306 3646 -11730
rect 3588 -12318 3646 -12306
rect 4606 -11730 4664 -11718
rect 4606 -12306 4618 -11730
rect 4652 -12306 4664 -11730
rect 4606 -12318 4664 -12306
rect 5624 -11730 5682 -11718
rect 5624 -12306 5636 -11730
rect 5670 -12306 5682 -11730
rect 5624 -12318 5682 -12306
rect 6642 -11730 6700 -11718
rect 6642 -12306 6654 -11730
rect 6688 -12306 6700 -11730
rect 6642 -12318 6700 -12306
rect 7660 -11730 7718 -11718
rect 7660 -12306 7672 -11730
rect 7706 -12306 7718 -11730
rect 7660 -12318 7718 -12306
rect 8678 -11730 8736 -11718
rect 8678 -12306 8690 -11730
rect 8724 -12306 8736 -11730
rect 8678 -12318 8736 -12306
rect 9696 -11730 9754 -11718
rect 9696 -12306 9708 -11730
rect 9742 -12306 9754 -11730
rect 9696 -12318 9754 -12306
rect 10714 -11730 10772 -11718
rect 10714 -12306 10726 -11730
rect 10760 -12306 10772 -11730
rect 10714 -12318 10772 -12306
rect 11732 -11730 11790 -11718
rect 11732 -12306 11744 -11730
rect 11778 -12306 11790 -11730
rect 11732 -12318 11790 -12306
rect 12750 -11730 12808 -11718
rect 12750 -12306 12762 -11730
rect 12796 -12306 12808 -11730
rect 12750 -12318 12808 -12306
rect 13768 -11730 13826 -11718
rect 13768 -12306 13780 -11730
rect 13814 -12306 13826 -11730
rect 13768 -12318 13826 -12306
rect 14786 -11730 14844 -11718
rect 14786 -12306 14798 -11730
rect 14832 -12306 14844 -11730
rect 14786 -12318 14844 -12306
rect 15804 -11730 15862 -11718
rect 15804 -12306 15816 -11730
rect 15850 -12306 15862 -11730
rect 15804 -12318 15862 -12306
rect 16822 -11730 16880 -11718
rect 16822 -12306 16834 -11730
rect 16868 -12306 16880 -11730
rect 16822 -12318 16880 -12306
rect 17840 -11730 17898 -11718
rect 17840 -12306 17852 -11730
rect 17886 -12306 17898 -11730
rect 17840 -12318 17898 -12306
rect 18858 -11730 18916 -11718
rect 18858 -12306 18870 -11730
rect 18904 -12306 18916 -11730
rect 18858 -12318 18916 -12306
rect 19876 -11730 19934 -11718
rect 19876 -12306 19888 -11730
rect 19922 -12306 19934 -11730
rect 19876 -12318 19934 -12306
rect 20894 -11730 20952 -11718
rect 20894 -12306 20906 -11730
rect 20940 -12306 20952 -11730
rect 20894 -12318 20952 -12306
rect 21912 -11730 21970 -11718
rect 21912 -12306 21924 -11730
rect 21958 -12306 21970 -11730
rect 21912 -12318 21970 -12306
rect 22930 -11730 22988 -11718
rect 22930 -12306 22942 -11730
rect 22976 -12306 22988 -11730
rect 22930 -12318 22988 -12306
rect -9196 -12524 -9138 -12512
rect -9196 -13100 -9184 -12524
rect -9150 -13100 -9138 -12524
rect -9196 -13112 -9138 -13100
rect -8178 -12524 -8120 -12512
rect -8178 -13100 -8166 -12524
rect -8132 -13100 -8120 -12524
rect -8178 -13112 -8120 -13100
rect -7160 -12524 -7102 -12512
rect -7160 -13100 -7148 -12524
rect -7114 -13100 -7102 -12524
rect -7160 -13112 -7102 -13100
rect -6142 -12524 -6084 -12512
rect -6142 -13100 -6130 -12524
rect -6096 -13100 -6084 -12524
rect -6142 -13112 -6084 -13100
rect -5124 -12524 -5066 -12512
rect -5124 -13100 -5112 -12524
rect -5078 -13100 -5066 -12524
rect -5124 -13112 -5066 -13100
rect -4106 -12524 -4048 -12512
rect -4106 -13100 -4094 -12524
rect -4060 -13100 -4048 -12524
rect -4106 -13112 -4048 -13100
rect -3088 -12524 -3030 -12512
rect -3088 -13100 -3076 -12524
rect -3042 -13100 -3030 -12524
rect -3088 -13112 -3030 -13100
rect -2070 -12524 -2012 -12512
rect -2070 -13100 -2058 -12524
rect -2024 -13100 -2012 -12524
rect -2070 -13112 -2012 -13100
rect -1052 -12524 -994 -12512
rect -1052 -13100 -1040 -12524
rect -1006 -13100 -994 -12524
rect -1052 -13112 -994 -13100
rect -34 -12524 24 -12512
rect -34 -13100 -22 -12524
rect 12 -13100 24 -12524
rect -34 -13112 24 -13100
rect 2570 -12964 2628 -12952
rect -9196 -13342 -9138 -13330
rect -9196 -13918 -9184 -13342
rect -9150 -13918 -9138 -13342
rect -9196 -13930 -9138 -13918
rect -8178 -13342 -8120 -13330
rect -8178 -13918 -8166 -13342
rect -8132 -13918 -8120 -13342
rect -8178 -13930 -8120 -13918
rect -7160 -13342 -7102 -13330
rect -7160 -13918 -7148 -13342
rect -7114 -13918 -7102 -13342
rect -7160 -13930 -7102 -13918
rect -6142 -13342 -6084 -13330
rect -6142 -13918 -6130 -13342
rect -6096 -13918 -6084 -13342
rect -6142 -13930 -6084 -13918
rect -5124 -13342 -5066 -13330
rect -5124 -13918 -5112 -13342
rect -5078 -13918 -5066 -13342
rect -5124 -13930 -5066 -13918
rect -4106 -13342 -4048 -13330
rect -4106 -13918 -4094 -13342
rect -4060 -13918 -4048 -13342
rect -4106 -13930 -4048 -13918
rect -3088 -13342 -3030 -13330
rect -3088 -13918 -3076 -13342
rect -3042 -13918 -3030 -13342
rect -3088 -13930 -3030 -13918
rect -2070 -13342 -2012 -13330
rect -2070 -13918 -2058 -13342
rect -2024 -13918 -2012 -13342
rect -2070 -13930 -2012 -13918
rect -1052 -13342 -994 -13330
rect -1052 -13918 -1040 -13342
rect -1006 -13918 -994 -13342
rect -1052 -13930 -994 -13918
rect -34 -13342 24 -13330
rect -34 -13918 -22 -13342
rect 12 -13918 24 -13342
rect 2570 -13540 2582 -12964
rect 2616 -13540 2628 -12964
rect 2570 -13552 2628 -13540
rect 3588 -12964 3646 -12952
rect 3588 -13540 3600 -12964
rect 3634 -13540 3646 -12964
rect 3588 -13552 3646 -13540
rect 4606 -12964 4664 -12952
rect 4606 -13540 4618 -12964
rect 4652 -13540 4664 -12964
rect 4606 -13552 4664 -13540
rect 5624 -12964 5682 -12952
rect 5624 -13540 5636 -12964
rect 5670 -13540 5682 -12964
rect 5624 -13552 5682 -13540
rect 6642 -12964 6700 -12952
rect 6642 -13540 6654 -12964
rect 6688 -13540 6700 -12964
rect 6642 -13552 6700 -13540
rect 7660 -12964 7718 -12952
rect 7660 -13540 7672 -12964
rect 7706 -13540 7718 -12964
rect 7660 -13552 7718 -13540
rect 8678 -12964 8736 -12952
rect 8678 -13540 8690 -12964
rect 8724 -13540 8736 -12964
rect 8678 -13552 8736 -13540
rect 9696 -12964 9754 -12952
rect 9696 -13540 9708 -12964
rect 9742 -13540 9754 -12964
rect 9696 -13552 9754 -13540
rect 10714 -12964 10772 -12952
rect 10714 -13540 10726 -12964
rect 10760 -13540 10772 -12964
rect 10714 -13552 10772 -13540
rect 11732 -12964 11790 -12952
rect 11732 -13540 11744 -12964
rect 11778 -13540 11790 -12964
rect 11732 -13552 11790 -13540
rect 12750 -12964 12808 -12952
rect 12750 -13540 12762 -12964
rect 12796 -13540 12808 -12964
rect 12750 -13552 12808 -13540
rect 13768 -12964 13826 -12952
rect 13768 -13540 13780 -12964
rect 13814 -13540 13826 -12964
rect 13768 -13552 13826 -13540
rect 14786 -12964 14844 -12952
rect 14786 -13540 14798 -12964
rect 14832 -13540 14844 -12964
rect 14786 -13552 14844 -13540
rect 15804 -12964 15862 -12952
rect 15804 -13540 15816 -12964
rect 15850 -13540 15862 -12964
rect 15804 -13552 15862 -13540
rect 16822 -12964 16880 -12952
rect 16822 -13540 16834 -12964
rect 16868 -13540 16880 -12964
rect 16822 -13552 16880 -13540
rect 17840 -12964 17898 -12952
rect 17840 -13540 17852 -12964
rect 17886 -13540 17898 -12964
rect 17840 -13552 17898 -13540
rect 18858 -12964 18916 -12952
rect 18858 -13540 18870 -12964
rect 18904 -13540 18916 -12964
rect 18858 -13552 18916 -13540
rect 19876 -12964 19934 -12952
rect 19876 -13540 19888 -12964
rect 19922 -13540 19934 -12964
rect 19876 -13552 19934 -13540
rect 20894 -12964 20952 -12952
rect 20894 -13540 20906 -12964
rect 20940 -13540 20952 -12964
rect 20894 -13552 20952 -13540
rect 21912 -12964 21970 -12952
rect 21912 -13540 21924 -12964
rect 21958 -13540 21970 -12964
rect 21912 -13552 21970 -13540
rect 22930 -12964 22988 -12952
rect 22930 -13540 22942 -12964
rect 22976 -13540 22988 -12964
rect 22930 -13552 22988 -13540
rect -34 -13930 24 -13918
rect -9196 -14160 -9138 -14148
rect -9196 -14736 -9184 -14160
rect -9150 -14736 -9138 -14160
rect -9196 -14748 -9138 -14736
rect -8178 -14160 -8120 -14148
rect -8178 -14736 -8166 -14160
rect -8132 -14736 -8120 -14160
rect -8178 -14748 -8120 -14736
rect -7160 -14160 -7102 -14148
rect -7160 -14736 -7148 -14160
rect -7114 -14736 -7102 -14160
rect -7160 -14748 -7102 -14736
rect -6142 -14160 -6084 -14148
rect -6142 -14736 -6130 -14160
rect -6096 -14736 -6084 -14160
rect -6142 -14748 -6084 -14736
rect -5124 -14160 -5066 -14148
rect -5124 -14736 -5112 -14160
rect -5078 -14736 -5066 -14160
rect -5124 -14748 -5066 -14736
rect -4106 -14160 -4048 -14148
rect -4106 -14736 -4094 -14160
rect -4060 -14736 -4048 -14160
rect -4106 -14748 -4048 -14736
rect -3088 -14160 -3030 -14148
rect -3088 -14736 -3076 -14160
rect -3042 -14736 -3030 -14160
rect -3088 -14748 -3030 -14736
rect -2070 -14160 -2012 -14148
rect -2070 -14736 -2058 -14160
rect -2024 -14736 -2012 -14160
rect -2070 -14748 -2012 -14736
rect -1052 -14160 -994 -14148
rect -1052 -14736 -1040 -14160
rect -1006 -14736 -994 -14160
rect -1052 -14748 -994 -14736
rect -34 -14160 24 -14148
rect -34 -14736 -22 -14160
rect 12 -14736 24 -14160
rect -34 -14748 24 -14736
rect 2570 -14196 2628 -14184
rect 2570 -14772 2582 -14196
rect 2616 -14772 2628 -14196
rect 2570 -14784 2628 -14772
rect 3588 -14196 3646 -14184
rect 3588 -14772 3600 -14196
rect 3634 -14772 3646 -14196
rect 3588 -14784 3646 -14772
rect 4606 -14196 4664 -14184
rect 4606 -14772 4618 -14196
rect 4652 -14772 4664 -14196
rect 4606 -14784 4664 -14772
rect 5624 -14196 5682 -14184
rect 5624 -14772 5636 -14196
rect 5670 -14772 5682 -14196
rect 5624 -14784 5682 -14772
rect 6642 -14196 6700 -14184
rect 6642 -14772 6654 -14196
rect 6688 -14772 6700 -14196
rect 6642 -14784 6700 -14772
rect 7660 -14196 7718 -14184
rect 7660 -14772 7672 -14196
rect 7706 -14772 7718 -14196
rect 7660 -14784 7718 -14772
rect 8678 -14196 8736 -14184
rect 8678 -14772 8690 -14196
rect 8724 -14772 8736 -14196
rect 8678 -14784 8736 -14772
rect 9696 -14196 9754 -14184
rect 9696 -14772 9708 -14196
rect 9742 -14772 9754 -14196
rect 9696 -14784 9754 -14772
rect 10714 -14196 10772 -14184
rect 10714 -14772 10726 -14196
rect 10760 -14772 10772 -14196
rect 10714 -14784 10772 -14772
rect 11732 -14196 11790 -14184
rect 11732 -14772 11744 -14196
rect 11778 -14772 11790 -14196
rect 11732 -14784 11790 -14772
rect 12750 -14196 12808 -14184
rect 12750 -14772 12762 -14196
rect 12796 -14772 12808 -14196
rect 12750 -14784 12808 -14772
rect 13768 -14196 13826 -14184
rect 13768 -14772 13780 -14196
rect 13814 -14772 13826 -14196
rect 13768 -14784 13826 -14772
rect 14786 -14196 14844 -14184
rect 14786 -14772 14798 -14196
rect 14832 -14772 14844 -14196
rect 14786 -14784 14844 -14772
rect 15804 -14196 15862 -14184
rect 15804 -14772 15816 -14196
rect 15850 -14772 15862 -14196
rect 15804 -14784 15862 -14772
rect 16822 -14196 16880 -14184
rect 16822 -14772 16834 -14196
rect 16868 -14772 16880 -14196
rect 16822 -14784 16880 -14772
rect 17840 -14196 17898 -14184
rect 17840 -14772 17852 -14196
rect 17886 -14772 17898 -14196
rect 17840 -14784 17898 -14772
rect 18858 -14196 18916 -14184
rect 18858 -14772 18870 -14196
rect 18904 -14772 18916 -14196
rect 18858 -14784 18916 -14772
rect 19876 -14196 19934 -14184
rect 19876 -14772 19888 -14196
rect 19922 -14772 19934 -14196
rect 19876 -14784 19934 -14772
rect 20894 -14196 20952 -14184
rect 20894 -14772 20906 -14196
rect 20940 -14772 20952 -14196
rect 20894 -14784 20952 -14772
rect 21912 -14196 21970 -14184
rect 21912 -14772 21924 -14196
rect 21958 -14772 21970 -14196
rect 21912 -14784 21970 -14772
rect 22930 -14196 22988 -14184
rect 22930 -14772 22942 -14196
rect 22976 -14772 22988 -14196
rect 22930 -14784 22988 -14772
rect -9196 -14978 -9138 -14966
rect -9196 -15554 -9184 -14978
rect -9150 -15554 -9138 -14978
rect -9196 -15566 -9138 -15554
rect -8178 -14978 -8120 -14966
rect -8178 -15554 -8166 -14978
rect -8132 -15554 -8120 -14978
rect -8178 -15566 -8120 -15554
rect -7160 -14978 -7102 -14966
rect -7160 -15554 -7148 -14978
rect -7114 -15554 -7102 -14978
rect -7160 -15566 -7102 -15554
rect -6142 -14978 -6084 -14966
rect -6142 -15554 -6130 -14978
rect -6096 -15554 -6084 -14978
rect -6142 -15566 -6084 -15554
rect -5124 -14978 -5066 -14966
rect -5124 -15554 -5112 -14978
rect -5078 -15554 -5066 -14978
rect -5124 -15566 -5066 -15554
rect -4106 -14978 -4048 -14966
rect -4106 -15554 -4094 -14978
rect -4060 -15554 -4048 -14978
rect -4106 -15566 -4048 -15554
rect -3088 -14978 -3030 -14966
rect -3088 -15554 -3076 -14978
rect -3042 -15554 -3030 -14978
rect -3088 -15566 -3030 -15554
rect -2070 -14978 -2012 -14966
rect -2070 -15554 -2058 -14978
rect -2024 -15554 -2012 -14978
rect -2070 -15566 -2012 -15554
rect -1052 -14978 -994 -14966
rect -1052 -15554 -1040 -14978
rect -1006 -15554 -994 -14978
rect -1052 -15566 -994 -15554
rect -34 -14978 24 -14966
rect -34 -15554 -22 -14978
rect 12 -15554 24 -14978
rect -34 -15566 24 -15554
rect 2568 -15430 2626 -15418
rect -9196 -15796 -9138 -15784
rect -9196 -16372 -9184 -15796
rect -9150 -16372 -9138 -15796
rect -9196 -16384 -9138 -16372
rect -8178 -15796 -8120 -15784
rect -8178 -16372 -8166 -15796
rect -8132 -16372 -8120 -15796
rect -8178 -16384 -8120 -16372
rect -7160 -15796 -7102 -15784
rect -7160 -16372 -7148 -15796
rect -7114 -16372 -7102 -15796
rect -7160 -16384 -7102 -16372
rect -6142 -15796 -6084 -15784
rect -6142 -16372 -6130 -15796
rect -6096 -16372 -6084 -15796
rect -6142 -16384 -6084 -16372
rect -5124 -15796 -5066 -15784
rect -5124 -16372 -5112 -15796
rect -5078 -16372 -5066 -15796
rect -5124 -16384 -5066 -16372
rect -4106 -15796 -4048 -15784
rect -4106 -16372 -4094 -15796
rect -4060 -16372 -4048 -15796
rect -4106 -16384 -4048 -16372
rect -3088 -15796 -3030 -15784
rect -3088 -16372 -3076 -15796
rect -3042 -16372 -3030 -15796
rect -3088 -16384 -3030 -16372
rect -2070 -15796 -2012 -15784
rect -2070 -16372 -2058 -15796
rect -2024 -16372 -2012 -15796
rect -2070 -16384 -2012 -16372
rect -1052 -15796 -994 -15784
rect -1052 -16372 -1040 -15796
rect -1006 -16372 -994 -15796
rect -1052 -16384 -994 -16372
rect -34 -15796 24 -15784
rect -34 -16372 -22 -15796
rect 12 -16372 24 -15796
rect 2568 -16006 2580 -15430
rect 2614 -16006 2626 -15430
rect 2568 -16018 2626 -16006
rect 3586 -15430 3644 -15418
rect 3586 -16006 3598 -15430
rect 3632 -16006 3644 -15430
rect 3586 -16018 3644 -16006
rect 4604 -15430 4662 -15418
rect 4604 -16006 4616 -15430
rect 4650 -16006 4662 -15430
rect 4604 -16018 4662 -16006
rect 5622 -15430 5680 -15418
rect 5622 -16006 5634 -15430
rect 5668 -16006 5680 -15430
rect 5622 -16018 5680 -16006
rect 6640 -15430 6698 -15418
rect 6640 -16006 6652 -15430
rect 6686 -16006 6698 -15430
rect 6640 -16018 6698 -16006
rect 7658 -15430 7716 -15418
rect 7658 -16006 7670 -15430
rect 7704 -16006 7716 -15430
rect 7658 -16018 7716 -16006
rect 8676 -15430 8734 -15418
rect 8676 -16006 8688 -15430
rect 8722 -16006 8734 -15430
rect 8676 -16018 8734 -16006
rect 9694 -15430 9752 -15418
rect 9694 -16006 9706 -15430
rect 9740 -16006 9752 -15430
rect 9694 -16018 9752 -16006
rect 10712 -15430 10770 -15418
rect 10712 -16006 10724 -15430
rect 10758 -16006 10770 -15430
rect 10712 -16018 10770 -16006
rect 11730 -15430 11788 -15418
rect 11730 -16006 11742 -15430
rect 11776 -16006 11788 -15430
rect 11730 -16018 11788 -16006
rect 12748 -15430 12806 -15418
rect 12748 -16006 12760 -15430
rect 12794 -16006 12806 -15430
rect 12748 -16018 12806 -16006
rect 13766 -15430 13824 -15418
rect 13766 -16006 13778 -15430
rect 13812 -16006 13824 -15430
rect 13766 -16018 13824 -16006
rect 14784 -15430 14842 -15418
rect 14784 -16006 14796 -15430
rect 14830 -16006 14842 -15430
rect 14784 -16018 14842 -16006
rect 15802 -15430 15860 -15418
rect 15802 -16006 15814 -15430
rect 15848 -16006 15860 -15430
rect 15802 -16018 15860 -16006
rect 16820 -15430 16878 -15418
rect 16820 -16006 16832 -15430
rect 16866 -16006 16878 -15430
rect 16820 -16018 16878 -16006
rect 17838 -15430 17896 -15418
rect 17838 -16006 17850 -15430
rect 17884 -16006 17896 -15430
rect 17838 -16018 17896 -16006
rect 18856 -15430 18914 -15418
rect 18856 -16006 18868 -15430
rect 18902 -16006 18914 -15430
rect 18856 -16018 18914 -16006
rect 19874 -15430 19932 -15418
rect 19874 -16006 19886 -15430
rect 19920 -16006 19932 -15430
rect 19874 -16018 19932 -16006
rect 20892 -15430 20950 -15418
rect 20892 -16006 20904 -15430
rect 20938 -16006 20950 -15430
rect 20892 -16018 20950 -16006
rect 21910 -15430 21968 -15418
rect 21910 -16006 21922 -15430
rect 21956 -16006 21968 -15430
rect 21910 -16018 21968 -16006
rect 22928 -15430 22986 -15418
rect 22928 -16006 22940 -15430
rect 22974 -16006 22986 -15430
rect 22928 -16018 22986 -16006
rect -34 -16384 24 -16372
rect -9196 -16614 -9138 -16602
rect -9196 -17190 -9184 -16614
rect -9150 -17190 -9138 -16614
rect -9196 -17202 -9138 -17190
rect -8178 -16614 -8120 -16602
rect -8178 -17190 -8166 -16614
rect -8132 -17190 -8120 -16614
rect -8178 -17202 -8120 -17190
rect -7160 -16614 -7102 -16602
rect -7160 -17190 -7148 -16614
rect -7114 -17190 -7102 -16614
rect -7160 -17202 -7102 -17190
rect -6142 -16614 -6084 -16602
rect -6142 -17190 -6130 -16614
rect -6096 -17190 -6084 -16614
rect -6142 -17202 -6084 -17190
rect -5124 -16614 -5066 -16602
rect -5124 -17190 -5112 -16614
rect -5078 -17190 -5066 -16614
rect -5124 -17202 -5066 -17190
rect -4106 -16614 -4048 -16602
rect -4106 -17190 -4094 -16614
rect -4060 -17190 -4048 -16614
rect -4106 -17202 -4048 -17190
rect -3088 -16614 -3030 -16602
rect -3088 -17190 -3076 -16614
rect -3042 -17190 -3030 -16614
rect -3088 -17202 -3030 -17190
rect -2070 -16614 -2012 -16602
rect -2070 -17190 -2058 -16614
rect -2024 -17190 -2012 -16614
rect -2070 -17202 -2012 -17190
rect -1052 -16614 -994 -16602
rect -1052 -17190 -1040 -16614
rect -1006 -17190 -994 -16614
rect -1052 -17202 -994 -17190
rect -34 -16614 24 -16602
rect -34 -17190 -22 -16614
rect 12 -17190 24 -16614
rect -34 -17202 24 -17190
rect 2568 -16664 2626 -16652
rect 2568 -17240 2580 -16664
rect 2614 -17240 2626 -16664
rect 2568 -17252 2626 -17240
rect 3586 -16664 3644 -16652
rect 3586 -17240 3598 -16664
rect 3632 -17240 3644 -16664
rect 3586 -17252 3644 -17240
rect 4604 -16664 4662 -16652
rect 4604 -17240 4616 -16664
rect 4650 -17240 4662 -16664
rect 4604 -17252 4662 -17240
rect 5622 -16664 5680 -16652
rect 5622 -17240 5634 -16664
rect 5668 -17240 5680 -16664
rect 5622 -17252 5680 -17240
rect 6640 -16664 6698 -16652
rect 6640 -17240 6652 -16664
rect 6686 -17240 6698 -16664
rect 6640 -17252 6698 -17240
rect 7658 -16664 7716 -16652
rect 7658 -17240 7670 -16664
rect 7704 -17240 7716 -16664
rect 7658 -17252 7716 -17240
rect 8676 -16664 8734 -16652
rect 8676 -17240 8688 -16664
rect 8722 -17240 8734 -16664
rect 8676 -17252 8734 -17240
rect 9694 -16664 9752 -16652
rect 9694 -17240 9706 -16664
rect 9740 -17240 9752 -16664
rect 9694 -17252 9752 -17240
rect 10712 -16664 10770 -16652
rect 10712 -17240 10724 -16664
rect 10758 -17240 10770 -16664
rect 10712 -17252 10770 -17240
rect 11730 -16664 11788 -16652
rect 11730 -17240 11742 -16664
rect 11776 -17240 11788 -16664
rect 11730 -17252 11788 -17240
rect 12748 -16664 12806 -16652
rect 12748 -17240 12760 -16664
rect 12794 -17240 12806 -16664
rect 12748 -17252 12806 -17240
rect 13766 -16664 13824 -16652
rect 13766 -17240 13778 -16664
rect 13812 -17240 13824 -16664
rect 13766 -17252 13824 -17240
rect 14784 -16664 14842 -16652
rect 14784 -17240 14796 -16664
rect 14830 -17240 14842 -16664
rect 14784 -17252 14842 -17240
rect 15802 -16664 15860 -16652
rect 15802 -17240 15814 -16664
rect 15848 -17240 15860 -16664
rect 15802 -17252 15860 -17240
rect 16820 -16664 16878 -16652
rect 16820 -17240 16832 -16664
rect 16866 -17240 16878 -16664
rect 16820 -17252 16878 -17240
rect 17838 -16664 17896 -16652
rect 17838 -17240 17850 -16664
rect 17884 -17240 17896 -16664
rect 17838 -17252 17896 -17240
rect 18856 -16664 18914 -16652
rect 18856 -17240 18868 -16664
rect 18902 -17240 18914 -16664
rect 18856 -17252 18914 -17240
rect 19874 -16664 19932 -16652
rect 19874 -17240 19886 -16664
rect 19920 -17240 19932 -16664
rect 19874 -17252 19932 -17240
rect 20892 -16664 20950 -16652
rect 20892 -17240 20904 -16664
rect 20938 -17240 20950 -16664
rect 20892 -17252 20950 -17240
rect 21910 -16664 21968 -16652
rect 21910 -17240 21922 -16664
rect 21956 -17240 21968 -16664
rect 21910 -17252 21968 -17240
rect 22928 -16664 22986 -16652
rect 22928 -17240 22940 -16664
rect 22974 -17240 22986 -16664
rect 22928 -17252 22986 -17240
rect -9196 -17432 -9138 -17420
rect -9196 -18008 -9184 -17432
rect -9150 -18008 -9138 -17432
rect -9196 -18020 -9138 -18008
rect -8178 -17432 -8120 -17420
rect -8178 -18008 -8166 -17432
rect -8132 -18008 -8120 -17432
rect -8178 -18020 -8120 -18008
rect -7160 -17432 -7102 -17420
rect -7160 -18008 -7148 -17432
rect -7114 -18008 -7102 -17432
rect -7160 -18020 -7102 -18008
rect -6142 -17432 -6084 -17420
rect -6142 -18008 -6130 -17432
rect -6096 -18008 -6084 -17432
rect -6142 -18020 -6084 -18008
rect -5124 -17432 -5066 -17420
rect -5124 -18008 -5112 -17432
rect -5078 -18008 -5066 -17432
rect -5124 -18020 -5066 -18008
rect -4106 -17432 -4048 -17420
rect -4106 -18008 -4094 -17432
rect -4060 -18008 -4048 -17432
rect -4106 -18020 -4048 -18008
rect -3088 -17432 -3030 -17420
rect -3088 -18008 -3076 -17432
rect -3042 -18008 -3030 -17432
rect -3088 -18020 -3030 -18008
rect -2070 -17432 -2012 -17420
rect -2070 -18008 -2058 -17432
rect -2024 -18008 -2012 -17432
rect -2070 -18020 -2012 -18008
rect -1052 -17432 -994 -17420
rect -1052 -18008 -1040 -17432
rect -1006 -18008 -994 -17432
rect -1052 -18020 -994 -18008
rect -34 -17432 24 -17420
rect -34 -18008 -22 -17432
rect 12 -18008 24 -17432
rect -34 -18020 24 -18008
rect 2568 -17896 2626 -17884
rect -9196 -18250 -9138 -18238
rect -9196 -18826 -9184 -18250
rect -9150 -18826 -9138 -18250
rect -9196 -18838 -9138 -18826
rect -8178 -18250 -8120 -18238
rect -8178 -18826 -8166 -18250
rect -8132 -18826 -8120 -18250
rect -8178 -18838 -8120 -18826
rect -7160 -18250 -7102 -18238
rect -7160 -18826 -7148 -18250
rect -7114 -18826 -7102 -18250
rect -7160 -18838 -7102 -18826
rect -6142 -18250 -6084 -18238
rect -6142 -18826 -6130 -18250
rect -6096 -18826 -6084 -18250
rect -6142 -18838 -6084 -18826
rect -5124 -18250 -5066 -18238
rect -5124 -18826 -5112 -18250
rect -5078 -18826 -5066 -18250
rect -5124 -18838 -5066 -18826
rect -4106 -18250 -4048 -18238
rect -4106 -18826 -4094 -18250
rect -4060 -18826 -4048 -18250
rect -4106 -18838 -4048 -18826
rect -3088 -18250 -3030 -18238
rect -3088 -18826 -3076 -18250
rect -3042 -18826 -3030 -18250
rect -3088 -18838 -3030 -18826
rect -2070 -18250 -2012 -18238
rect -2070 -18826 -2058 -18250
rect -2024 -18826 -2012 -18250
rect -2070 -18838 -2012 -18826
rect -1052 -18250 -994 -18238
rect -1052 -18826 -1040 -18250
rect -1006 -18826 -994 -18250
rect -1052 -18838 -994 -18826
rect -34 -18250 24 -18238
rect -34 -18826 -22 -18250
rect 12 -18826 24 -18250
rect 2568 -18472 2580 -17896
rect 2614 -18472 2626 -17896
rect 2568 -18484 2626 -18472
rect 3586 -17896 3644 -17884
rect 3586 -18472 3598 -17896
rect 3632 -18472 3644 -17896
rect 3586 -18484 3644 -18472
rect 4604 -17896 4662 -17884
rect 4604 -18472 4616 -17896
rect 4650 -18472 4662 -17896
rect 4604 -18484 4662 -18472
rect 5622 -17896 5680 -17884
rect 5622 -18472 5634 -17896
rect 5668 -18472 5680 -17896
rect 5622 -18484 5680 -18472
rect 6640 -17896 6698 -17884
rect 6640 -18472 6652 -17896
rect 6686 -18472 6698 -17896
rect 6640 -18484 6698 -18472
rect 7658 -17896 7716 -17884
rect 7658 -18472 7670 -17896
rect 7704 -18472 7716 -17896
rect 7658 -18484 7716 -18472
rect 8676 -17896 8734 -17884
rect 8676 -18472 8688 -17896
rect 8722 -18472 8734 -17896
rect 8676 -18484 8734 -18472
rect 9694 -17896 9752 -17884
rect 9694 -18472 9706 -17896
rect 9740 -18472 9752 -17896
rect 9694 -18484 9752 -18472
rect 10712 -17896 10770 -17884
rect 10712 -18472 10724 -17896
rect 10758 -18472 10770 -17896
rect 10712 -18484 10770 -18472
rect 11730 -17896 11788 -17884
rect 11730 -18472 11742 -17896
rect 11776 -18472 11788 -17896
rect 11730 -18484 11788 -18472
rect 12748 -17896 12806 -17884
rect 12748 -18472 12760 -17896
rect 12794 -18472 12806 -17896
rect 12748 -18484 12806 -18472
rect 13766 -17896 13824 -17884
rect 13766 -18472 13778 -17896
rect 13812 -18472 13824 -17896
rect 13766 -18484 13824 -18472
rect 14784 -17896 14842 -17884
rect 14784 -18472 14796 -17896
rect 14830 -18472 14842 -17896
rect 14784 -18484 14842 -18472
rect 15802 -17896 15860 -17884
rect 15802 -18472 15814 -17896
rect 15848 -18472 15860 -17896
rect 15802 -18484 15860 -18472
rect 16820 -17896 16878 -17884
rect 16820 -18472 16832 -17896
rect 16866 -18472 16878 -17896
rect 16820 -18484 16878 -18472
rect 17838 -17896 17896 -17884
rect 17838 -18472 17850 -17896
rect 17884 -18472 17896 -17896
rect 17838 -18484 17896 -18472
rect 18856 -17896 18914 -17884
rect 18856 -18472 18868 -17896
rect 18902 -18472 18914 -17896
rect 18856 -18484 18914 -18472
rect 19874 -17896 19932 -17884
rect 19874 -18472 19886 -17896
rect 19920 -18472 19932 -17896
rect 19874 -18484 19932 -18472
rect 20892 -17896 20950 -17884
rect 20892 -18472 20904 -17896
rect 20938 -18472 20950 -17896
rect 20892 -18484 20950 -18472
rect 21910 -17896 21968 -17884
rect 21910 -18472 21922 -17896
rect 21956 -18472 21968 -17896
rect 21910 -18484 21968 -18472
rect 22928 -17896 22986 -17884
rect 22928 -18472 22940 -17896
rect 22974 -18472 22986 -17896
rect 22928 -18484 22986 -18472
rect -34 -18838 24 -18826
rect 2568 -19130 2626 -19118
rect -2336 -19634 -2278 -19622
rect -2336 -19810 -2324 -19634
rect -2290 -19810 -2278 -19634
rect -2336 -19822 -2278 -19810
rect -2118 -19634 -2060 -19622
rect -2118 -19810 -2106 -19634
rect -2072 -19810 -2060 -19634
rect -2118 -19822 -2060 -19810
rect -1900 -19634 -1842 -19622
rect -1900 -19810 -1888 -19634
rect -1854 -19810 -1842 -19634
rect -1900 -19822 -1842 -19810
rect -1682 -19634 -1624 -19622
rect -1682 -19810 -1670 -19634
rect -1636 -19810 -1624 -19634
rect -1682 -19822 -1624 -19810
rect -1464 -19634 -1406 -19622
rect -1464 -19810 -1452 -19634
rect -1418 -19810 -1406 -19634
rect -1464 -19822 -1406 -19810
rect -1246 -19634 -1188 -19622
rect -1246 -19810 -1234 -19634
rect -1200 -19810 -1188 -19634
rect -1246 -19822 -1188 -19810
rect -1028 -19634 -970 -19622
rect -1028 -19810 -1016 -19634
rect -982 -19810 -970 -19634
rect -1028 -19822 -970 -19810
rect -810 -19634 -752 -19622
rect -810 -19810 -798 -19634
rect -764 -19810 -752 -19634
rect -810 -19822 -752 -19810
rect -592 -19634 -534 -19622
rect -592 -19810 -580 -19634
rect -546 -19810 -534 -19634
rect -592 -19822 -534 -19810
rect -374 -19634 -316 -19622
rect -374 -19810 -362 -19634
rect -328 -19810 -316 -19634
rect -374 -19822 -316 -19810
rect -156 -19634 -98 -19622
rect -156 -19810 -144 -19634
rect -110 -19810 -98 -19634
rect 2568 -19706 2580 -19130
rect 2614 -19706 2626 -19130
rect 2568 -19718 2626 -19706
rect 3586 -19130 3644 -19118
rect 3586 -19706 3598 -19130
rect 3632 -19706 3644 -19130
rect 3586 -19718 3644 -19706
rect 4604 -19130 4662 -19118
rect 4604 -19706 4616 -19130
rect 4650 -19706 4662 -19130
rect 4604 -19718 4662 -19706
rect 5622 -19130 5680 -19118
rect 5622 -19706 5634 -19130
rect 5668 -19706 5680 -19130
rect 5622 -19718 5680 -19706
rect 6640 -19130 6698 -19118
rect 6640 -19706 6652 -19130
rect 6686 -19706 6698 -19130
rect 6640 -19718 6698 -19706
rect 7658 -19130 7716 -19118
rect 7658 -19706 7670 -19130
rect 7704 -19706 7716 -19130
rect 7658 -19718 7716 -19706
rect 8676 -19130 8734 -19118
rect 8676 -19706 8688 -19130
rect 8722 -19706 8734 -19130
rect 8676 -19718 8734 -19706
rect 9694 -19130 9752 -19118
rect 9694 -19706 9706 -19130
rect 9740 -19706 9752 -19130
rect 9694 -19718 9752 -19706
rect 10712 -19130 10770 -19118
rect 10712 -19706 10724 -19130
rect 10758 -19706 10770 -19130
rect 10712 -19718 10770 -19706
rect 11730 -19130 11788 -19118
rect 11730 -19706 11742 -19130
rect 11776 -19706 11788 -19130
rect 11730 -19718 11788 -19706
rect 12748 -19130 12806 -19118
rect 12748 -19706 12760 -19130
rect 12794 -19706 12806 -19130
rect 12748 -19718 12806 -19706
rect 13766 -19130 13824 -19118
rect 13766 -19706 13778 -19130
rect 13812 -19706 13824 -19130
rect 13766 -19718 13824 -19706
rect 14784 -19130 14842 -19118
rect 14784 -19706 14796 -19130
rect 14830 -19706 14842 -19130
rect 14784 -19718 14842 -19706
rect 15802 -19130 15860 -19118
rect 15802 -19706 15814 -19130
rect 15848 -19706 15860 -19130
rect 15802 -19718 15860 -19706
rect 16820 -19130 16878 -19118
rect 16820 -19706 16832 -19130
rect 16866 -19706 16878 -19130
rect 16820 -19718 16878 -19706
rect 17838 -19130 17896 -19118
rect 17838 -19706 17850 -19130
rect 17884 -19706 17896 -19130
rect 17838 -19718 17896 -19706
rect 18856 -19130 18914 -19118
rect 18856 -19706 18868 -19130
rect 18902 -19706 18914 -19130
rect 18856 -19718 18914 -19706
rect 19874 -19130 19932 -19118
rect 19874 -19706 19886 -19130
rect 19920 -19706 19932 -19130
rect 19874 -19718 19932 -19706
rect 20892 -19130 20950 -19118
rect 20892 -19706 20904 -19130
rect 20938 -19706 20950 -19130
rect 20892 -19718 20950 -19706
rect 21910 -19130 21968 -19118
rect 21910 -19706 21922 -19130
rect 21956 -19706 21968 -19130
rect 21910 -19718 21968 -19706
rect 22928 -19130 22986 -19118
rect 22928 -19706 22940 -19130
rect 22974 -19706 22986 -19130
rect 22928 -19718 22986 -19706
rect -156 -19822 -98 -19810
rect 2568 -20364 2626 -20352
rect -2336 -20466 -2278 -20454
rect -2336 -20642 -2324 -20466
rect -2290 -20642 -2278 -20466
rect -2336 -20654 -2278 -20642
rect -2118 -20466 -2060 -20454
rect -2118 -20642 -2106 -20466
rect -2072 -20642 -2060 -20466
rect -2118 -20654 -2060 -20642
rect -1900 -20466 -1842 -20454
rect -1900 -20642 -1888 -20466
rect -1854 -20642 -1842 -20466
rect -1900 -20654 -1842 -20642
rect -1682 -20466 -1624 -20454
rect -1682 -20642 -1670 -20466
rect -1636 -20642 -1624 -20466
rect -1682 -20654 -1624 -20642
rect -1464 -20466 -1406 -20454
rect -1464 -20642 -1452 -20466
rect -1418 -20642 -1406 -20466
rect -1464 -20654 -1406 -20642
rect -1246 -20466 -1188 -20454
rect -1246 -20642 -1234 -20466
rect -1200 -20642 -1188 -20466
rect -1246 -20654 -1188 -20642
rect -1028 -20466 -970 -20454
rect -1028 -20642 -1016 -20466
rect -982 -20642 -970 -20466
rect -1028 -20654 -970 -20642
rect -810 -20466 -752 -20454
rect -810 -20642 -798 -20466
rect -764 -20642 -752 -20466
rect -810 -20654 -752 -20642
rect -592 -20466 -534 -20454
rect -592 -20642 -580 -20466
rect -546 -20642 -534 -20466
rect -592 -20654 -534 -20642
rect -374 -20466 -316 -20454
rect -374 -20642 -362 -20466
rect -328 -20642 -316 -20466
rect -374 -20654 -316 -20642
rect -156 -20466 -98 -20454
rect -156 -20642 -144 -20466
rect -110 -20642 -98 -20466
rect -156 -20654 -98 -20642
rect 2568 -20940 2580 -20364
rect 2614 -20940 2626 -20364
rect 2568 -20952 2626 -20940
rect 3586 -20364 3644 -20352
rect 3586 -20940 3598 -20364
rect 3632 -20940 3644 -20364
rect 3586 -20952 3644 -20940
rect 4604 -20364 4662 -20352
rect 4604 -20940 4616 -20364
rect 4650 -20940 4662 -20364
rect 4604 -20952 4662 -20940
rect 5622 -20364 5680 -20352
rect 5622 -20940 5634 -20364
rect 5668 -20940 5680 -20364
rect 5622 -20952 5680 -20940
rect 6640 -20364 6698 -20352
rect 6640 -20940 6652 -20364
rect 6686 -20940 6698 -20364
rect 6640 -20952 6698 -20940
rect 7658 -20364 7716 -20352
rect 7658 -20940 7670 -20364
rect 7704 -20940 7716 -20364
rect 7658 -20952 7716 -20940
rect 8676 -20364 8734 -20352
rect 8676 -20940 8688 -20364
rect 8722 -20940 8734 -20364
rect 8676 -20952 8734 -20940
rect 9694 -20364 9752 -20352
rect 9694 -20940 9706 -20364
rect 9740 -20940 9752 -20364
rect 9694 -20952 9752 -20940
rect 10712 -20364 10770 -20352
rect 10712 -20940 10724 -20364
rect 10758 -20940 10770 -20364
rect 10712 -20952 10770 -20940
rect 11730 -20364 11788 -20352
rect 11730 -20940 11742 -20364
rect 11776 -20940 11788 -20364
rect 11730 -20952 11788 -20940
rect 12748 -20364 12806 -20352
rect 12748 -20940 12760 -20364
rect 12794 -20940 12806 -20364
rect 12748 -20952 12806 -20940
rect 13766 -20364 13824 -20352
rect 13766 -20940 13778 -20364
rect 13812 -20940 13824 -20364
rect 13766 -20952 13824 -20940
rect 14784 -20364 14842 -20352
rect 14784 -20940 14796 -20364
rect 14830 -20940 14842 -20364
rect 14784 -20952 14842 -20940
rect 15802 -20364 15860 -20352
rect 15802 -20940 15814 -20364
rect 15848 -20940 15860 -20364
rect 15802 -20952 15860 -20940
rect 16820 -20364 16878 -20352
rect 16820 -20940 16832 -20364
rect 16866 -20940 16878 -20364
rect 16820 -20952 16878 -20940
rect 17838 -20364 17896 -20352
rect 17838 -20940 17850 -20364
rect 17884 -20940 17896 -20364
rect 17838 -20952 17896 -20940
rect 18856 -20364 18914 -20352
rect 18856 -20940 18868 -20364
rect 18902 -20940 18914 -20364
rect 18856 -20952 18914 -20940
rect 19874 -20364 19932 -20352
rect 19874 -20940 19886 -20364
rect 19920 -20940 19932 -20364
rect 19874 -20952 19932 -20940
rect 20892 -20364 20950 -20352
rect 20892 -20940 20904 -20364
rect 20938 -20940 20950 -20364
rect 20892 -20952 20950 -20940
rect 21910 -20364 21968 -20352
rect 21910 -20940 21922 -20364
rect 21956 -20940 21968 -20364
rect 21910 -20952 21968 -20940
rect 22928 -20364 22986 -20352
rect 22928 -20940 22940 -20364
rect 22974 -20940 22986 -20364
rect 22928 -20952 22986 -20940
rect 2568 -21596 2626 -21584
rect -9417 -21793 -9359 -21781
rect -9417 -22369 -9405 -21793
rect -9371 -22369 -9359 -21793
rect -9417 -22381 -9359 -22369
rect -8399 -21793 -8341 -21781
rect -8399 -22369 -8387 -21793
rect -8353 -22369 -8341 -21793
rect -8399 -22381 -8341 -22369
rect -7381 -21793 -7323 -21781
rect -7381 -22369 -7369 -21793
rect -7335 -22369 -7323 -21793
rect -7381 -22381 -7323 -22369
rect -6363 -21793 -6305 -21781
rect -6363 -22369 -6351 -21793
rect -6317 -22369 -6305 -21793
rect -6363 -22381 -6305 -22369
rect -5345 -21793 -5287 -21781
rect -5345 -22369 -5333 -21793
rect -5299 -22369 -5287 -21793
rect -5345 -22381 -5287 -22369
rect -4327 -21793 -4269 -21781
rect -4327 -22369 -4315 -21793
rect -4281 -22369 -4269 -21793
rect -4327 -22381 -4269 -22369
rect -3309 -21793 -3251 -21781
rect -3309 -22369 -3297 -21793
rect -3263 -22369 -3251 -21793
rect -3309 -22381 -3251 -22369
rect -2422 -21792 -2364 -21780
rect -2422 -22368 -2410 -21792
rect -2376 -22368 -2364 -21792
rect -2422 -22380 -2364 -22368
rect -2124 -21792 -2066 -21780
rect -2124 -22368 -2112 -21792
rect -2078 -22368 -2066 -21792
rect -2124 -22380 -2066 -22368
rect -1826 -21792 -1768 -21780
rect -1826 -22368 -1814 -21792
rect -1780 -22368 -1768 -21792
rect -1826 -22380 -1768 -22368
rect -1528 -21792 -1470 -21780
rect -1528 -22368 -1516 -21792
rect -1482 -22368 -1470 -21792
rect -1528 -22380 -1470 -22368
rect -1230 -21792 -1172 -21780
rect -1230 -22368 -1218 -21792
rect -1184 -22368 -1172 -21792
rect -1230 -22380 -1172 -22368
rect -932 -21792 -874 -21780
rect -932 -22368 -920 -21792
rect -886 -22368 -874 -21792
rect -932 -22380 -874 -22368
rect -634 -21792 -576 -21780
rect -634 -22368 -622 -21792
rect -588 -22368 -576 -21792
rect -634 -22380 -576 -22368
rect -336 -21792 -278 -21780
rect -336 -22368 -324 -21792
rect -290 -22368 -278 -21792
rect -336 -22380 -278 -22368
rect -38 -21792 20 -21780
rect -38 -22368 -26 -21792
rect 8 -22368 20 -21792
rect -38 -22380 20 -22368
rect 260 -21792 318 -21780
rect 260 -22368 272 -21792
rect 306 -22368 318 -21792
rect 260 -22380 318 -22368
rect 558 -21792 616 -21780
rect 558 -22368 570 -21792
rect 604 -22368 616 -21792
rect 558 -22380 616 -22368
rect 856 -21792 914 -21780
rect 856 -22368 868 -21792
rect 902 -22368 914 -21792
rect 2568 -22172 2580 -21596
rect 2614 -22172 2626 -21596
rect 2568 -22184 2626 -22172
rect 3586 -21596 3644 -21584
rect 3586 -22172 3598 -21596
rect 3632 -22172 3644 -21596
rect 3586 -22184 3644 -22172
rect 4604 -21596 4662 -21584
rect 4604 -22172 4616 -21596
rect 4650 -22172 4662 -21596
rect 4604 -22184 4662 -22172
rect 5622 -21596 5680 -21584
rect 5622 -22172 5634 -21596
rect 5668 -22172 5680 -21596
rect 5622 -22184 5680 -22172
rect 6640 -21596 6698 -21584
rect 6640 -22172 6652 -21596
rect 6686 -22172 6698 -21596
rect 6640 -22184 6698 -22172
rect 7658 -21596 7716 -21584
rect 7658 -22172 7670 -21596
rect 7704 -22172 7716 -21596
rect 7658 -22184 7716 -22172
rect 8676 -21596 8734 -21584
rect 8676 -22172 8688 -21596
rect 8722 -22172 8734 -21596
rect 8676 -22184 8734 -22172
rect 9694 -21596 9752 -21584
rect 9694 -22172 9706 -21596
rect 9740 -22172 9752 -21596
rect 9694 -22184 9752 -22172
rect 10712 -21596 10770 -21584
rect 10712 -22172 10724 -21596
rect 10758 -22172 10770 -21596
rect 10712 -22184 10770 -22172
rect 11730 -21596 11788 -21584
rect 11730 -22172 11742 -21596
rect 11776 -22172 11788 -21596
rect 11730 -22184 11788 -22172
rect 12748 -21596 12806 -21584
rect 12748 -22172 12760 -21596
rect 12794 -22172 12806 -21596
rect 12748 -22184 12806 -22172
rect 13766 -21596 13824 -21584
rect 13766 -22172 13778 -21596
rect 13812 -22172 13824 -21596
rect 13766 -22184 13824 -22172
rect 14784 -21596 14842 -21584
rect 14784 -22172 14796 -21596
rect 14830 -22172 14842 -21596
rect 14784 -22184 14842 -22172
rect 15802 -21596 15860 -21584
rect 15802 -22172 15814 -21596
rect 15848 -22172 15860 -21596
rect 15802 -22184 15860 -22172
rect 16820 -21596 16878 -21584
rect 16820 -22172 16832 -21596
rect 16866 -22172 16878 -21596
rect 16820 -22184 16878 -22172
rect 17838 -21596 17896 -21584
rect 17838 -22172 17850 -21596
rect 17884 -22172 17896 -21596
rect 17838 -22184 17896 -22172
rect 18856 -21596 18914 -21584
rect 18856 -22172 18868 -21596
rect 18902 -22172 18914 -21596
rect 18856 -22184 18914 -22172
rect 19874 -21596 19932 -21584
rect 19874 -22172 19886 -21596
rect 19920 -22172 19932 -21596
rect 19874 -22184 19932 -22172
rect 20892 -21596 20950 -21584
rect 20892 -22172 20904 -21596
rect 20938 -22172 20950 -21596
rect 20892 -22184 20950 -22172
rect 21910 -21596 21968 -21584
rect 21910 -22172 21922 -21596
rect 21956 -22172 21968 -21596
rect 21910 -22184 21968 -22172
rect 22928 -21596 22986 -21584
rect 22928 -22172 22940 -21596
rect 22974 -22172 22986 -21596
rect 22928 -22184 22986 -22172
rect 856 -22380 914 -22368
rect 2568 -22830 2626 -22818
rect -9418 -22906 -9360 -22894
rect -9418 -23482 -9406 -22906
rect -9372 -23482 -9360 -22906
rect -9418 -23494 -9360 -23482
rect -8400 -22906 -8342 -22894
rect -8400 -23482 -8388 -22906
rect -8354 -23482 -8342 -22906
rect -8400 -23494 -8342 -23482
rect -7382 -22906 -7324 -22894
rect -7382 -23482 -7370 -22906
rect -7336 -23482 -7324 -22906
rect -7382 -23494 -7324 -23482
rect -6364 -22906 -6306 -22894
rect -6364 -23482 -6352 -22906
rect -6318 -23482 -6306 -22906
rect -6364 -23494 -6306 -23482
rect -5346 -22906 -5288 -22894
rect -5346 -23482 -5334 -22906
rect -5300 -23482 -5288 -22906
rect -5346 -23494 -5288 -23482
rect -4328 -22906 -4270 -22894
rect -4328 -23482 -4316 -22906
rect -4282 -23482 -4270 -22906
rect -4328 -23494 -4270 -23482
rect -3310 -22906 -3252 -22894
rect -3310 -23482 -3298 -22906
rect -3264 -23482 -3252 -22906
rect -3310 -23494 -3252 -23482
rect -2422 -22904 -2364 -22892
rect -2422 -23480 -2410 -22904
rect -2376 -23480 -2364 -22904
rect -2422 -23492 -2364 -23480
rect -2124 -22904 -2066 -22892
rect -2124 -23480 -2112 -22904
rect -2078 -23480 -2066 -22904
rect -2124 -23492 -2066 -23480
rect -1826 -22904 -1768 -22892
rect -1826 -23480 -1814 -22904
rect -1780 -23480 -1768 -22904
rect -1826 -23492 -1768 -23480
rect -1528 -22904 -1470 -22892
rect -1528 -23480 -1516 -22904
rect -1482 -23480 -1470 -22904
rect -1528 -23492 -1470 -23480
rect -1230 -22904 -1172 -22892
rect -1230 -23480 -1218 -22904
rect -1184 -23480 -1172 -22904
rect -1230 -23492 -1172 -23480
rect -932 -22904 -874 -22892
rect -932 -23480 -920 -22904
rect -886 -23480 -874 -22904
rect -932 -23492 -874 -23480
rect -634 -22904 -576 -22892
rect -634 -23480 -622 -22904
rect -588 -23480 -576 -22904
rect -634 -23492 -576 -23480
rect -336 -22904 -278 -22892
rect -336 -23480 -324 -22904
rect -290 -23480 -278 -22904
rect -336 -23492 -278 -23480
rect -38 -22904 20 -22892
rect -38 -23480 -26 -22904
rect 8 -23480 20 -22904
rect -38 -23492 20 -23480
rect 260 -22904 318 -22892
rect 260 -23480 272 -22904
rect 306 -23480 318 -22904
rect 260 -23492 318 -23480
rect 558 -22904 616 -22892
rect 558 -23480 570 -22904
rect 604 -23480 616 -22904
rect 558 -23492 616 -23480
rect 856 -22904 914 -22892
rect 856 -23480 868 -22904
rect 902 -23480 914 -22904
rect 2568 -23406 2580 -22830
rect 2614 -23406 2626 -22830
rect 2568 -23418 2626 -23406
rect 3586 -22830 3644 -22818
rect 3586 -23406 3598 -22830
rect 3632 -23406 3644 -22830
rect 3586 -23418 3644 -23406
rect 4604 -22830 4662 -22818
rect 4604 -23406 4616 -22830
rect 4650 -23406 4662 -22830
rect 4604 -23418 4662 -23406
rect 5622 -22830 5680 -22818
rect 5622 -23406 5634 -22830
rect 5668 -23406 5680 -22830
rect 5622 -23418 5680 -23406
rect 6640 -22830 6698 -22818
rect 6640 -23406 6652 -22830
rect 6686 -23406 6698 -22830
rect 6640 -23418 6698 -23406
rect 7658 -22830 7716 -22818
rect 7658 -23406 7670 -22830
rect 7704 -23406 7716 -22830
rect 7658 -23418 7716 -23406
rect 8676 -22830 8734 -22818
rect 8676 -23406 8688 -22830
rect 8722 -23406 8734 -22830
rect 8676 -23418 8734 -23406
rect 9694 -22830 9752 -22818
rect 9694 -23406 9706 -22830
rect 9740 -23406 9752 -22830
rect 9694 -23418 9752 -23406
rect 10712 -22830 10770 -22818
rect 10712 -23406 10724 -22830
rect 10758 -23406 10770 -22830
rect 10712 -23418 10770 -23406
rect 11730 -22830 11788 -22818
rect 11730 -23406 11742 -22830
rect 11776 -23406 11788 -22830
rect 11730 -23418 11788 -23406
rect 12748 -22830 12806 -22818
rect 12748 -23406 12760 -22830
rect 12794 -23406 12806 -22830
rect 12748 -23418 12806 -23406
rect 13766 -22830 13824 -22818
rect 13766 -23406 13778 -22830
rect 13812 -23406 13824 -22830
rect 13766 -23418 13824 -23406
rect 14784 -22830 14842 -22818
rect 14784 -23406 14796 -22830
rect 14830 -23406 14842 -22830
rect 14784 -23418 14842 -23406
rect 15802 -22830 15860 -22818
rect 15802 -23406 15814 -22830
rect 15848 -23406 15860 -22830
rect 15802 -23418 15860 -23406
rect 16820 -22830 16878 -22818
rect 16820 -23406 16832 -22830
rect 16866 -23406 16878 -22830
rect 16820 -23418 16878 -23406
rect 17838 -22830 17896 -22818
rect 17838 -23406 17850 -22830
rect 17884 -23406 17896 -22830
rect 17838 -23418 17896 -23406
rect 18856 -22830 18914 -22818
rect 18856 -23406 18868 -22830
rect 18902 -23406 18914 -22830
rect 18856 -23418 18914 -23406
rect 19874 -22830 19932 -22818
rect 19874 -23406 19886 -22830
rect 19920 -23406 19932 -22830
rect 19874 -23418 19932 -23406
rect 20892 -22830 20950 -22818
rect 20892 -23406 20904 -22830
rect 20938 -23406 20950 -22830
rect 20892 -23418 20950 -23406
rect 21910 -22830 21968 -22818
rect 21910 -23406 21922 -22830
rect 21956 -23406 21968 -22830
rect 21910 -23418 21968 -23406
rect 22928 -22830 22986 -22818
rect 22928 -23406 22940 -22830
rect 22974 -23406 22986 -22830
rect 22928 -23418 22986 -23406
rect 856 -23492 914 -23480
rect -9417 -24017 -9359 -24005
rect -9417 -24593 -9405 -24017
rect -9371 -24593 -9359 -24017
rect -9417 -24605 -9359 -24593
rect -8399 -24017 -8341 -24005
rect -8399 -24593 -8387 -24017
rect -8353 -24593 -8341 -24017
rect -8399 -24605 -8341 -24593
rect -7381 -24017 -7323 -24005
rect -7381 -24593 -7369 -24017
rect -7335 -24593 -7323 -24017
rect -7381 -24605 -7323 -24593
rect -6363 -24017 -6305 -24005
rect -6363 -24593 -6351 -24017
rect -6317 -24593 -6305 -24017
rect -6363 -24605 -6305 -24593
rect -5345 -24017 -5287 -24005
rect -5345 -24593 -5333 -24017
rect -5299 -24593 -5287 -24017
rect -5345 -24605 -5287 -24593
rect -4327 -24017 -4269 -24005
rect -4327 -24593 -4315 -24017
rect -4281 -24593 -4269 -24017
rect -4327 -24605 -4269 -24593
rect -3309 -24017 -3251 -24005
rect -3309 -24593 -3297 -24017
rect -3263 -24593 -3251 -24017
rect -3309 -24605 -3251 -24593
rect -2424 -24016 -2366 -24004
rect -2424 -24592 -2412 -24016
rect -2378 -24592 -2366 -24016
rect -2424 -24604 -2366 -24592
rect -2126 -24016 -2068 -24004
rect -2126 -24592 -2114 -24016
rect -2080 -24592 -2068 -24016
rect -2126 -24604 -2068 -24592
rect -1828 -24016 -1770 -24004
rect -1828 -24592 -1816 -24016
rect -1782 -24592 -1770 -24016
rect -1828 -24604 -1770 -24592
rect -1530 -24016 -1472 -24004
rect -1530 -24592 -1518 -24016
rect -1484 -24592 -1472 -24016
rect -1530 -24604 -1472 -24592
rect -1232 -24016 -1174 -24004
rect -1232 -24592 -1220 -24016
rect -1186 -24592 -1174 -24016
rect -1232 -24604 -1174 -24592
rect -934 -24016 -876 -24004
rect -934 -24592 -922 -24016
rect -888 -24592 -876 -24016
rect -934 -24604 -876 -24592
rect -636 -24016 -578 -24004
rect -636 -24592 -624 -24016
rect -590 -24592 -578 -24016
rect -636 -24604 -578 -24592
rect -338 -24016 -280 -24004
rect -338 -24592 -326 -24016
rect -292 -24592 -280 -24016
rect -338 -24604 -280 -24592
rect -40 -24016 18 -24004
rect -40 -24592 -28 -24016
rect 6 -24592 18 -24016
rect -40 -24604 18 -24592
rect 258 -24016 316 -24004
rect 258 -24592 270 -24016
rect 304 -24592 316 -24016
rect 258 -24604 316 -24592
rect 556 -24016 614 -24004
rect 556 -24592 568 -24016
rect 602 -24592 614 -24016
rect 556 -24604 614 -24592
rect 854 -24016 912 -24004
rect 854 -24592 866 -24016
rect 900 -24592 912 -24016
rect 854 -24604 912 -24592
rect 2568 -24064 2626 -24052
rect 2568 -24640 2580 -24064
rect 2614 -24640 2626 -24064
rect 2568 -24652 2626 -24640
rect 3586 -24064 3644 -24052
rect 3586 -24640 3598 -24064
rect 3632 -24640 3644 -24064
rect 3586 -24652 3644 -24640
rect 4604 -24064 4662 -24052
rect 4604 -24640 4616 -24064
rect 4650 -24640 4662 -24064
rect 4604 -24652 4662 -24640
rect 5622 -24064 5680 -24052
rect 5622 -24640 5634 -24064
rect 5668 -24640 5680 -24064
rect 5622 -24652 5680 -24640
rect 6640 -24064 6698 -24052
rect 6640 -24640 6652 -24064
rect 6686 -24640 6698 -24064
rect 6640 -24652 6698 -24640
rect 7658 -24064 7716 -24052
rect 7658 -24640 7670 -24064
rect 7704 -24640 7716 -24064
rect 7658 -24652 7716 -24640
rect 8676 -24064 8734 -24052
rect 8676 -24640 8688 -24064
rect 8722 -24640 8734 -24064
rect 8676 -24652 8734 -24640
rect 9694 -24064 9752 -24052
rect 9694 -24640 9706 -24064
rect 9740 -24640 9752 -24064
rect 9694 -24652 9752 -24640
rect 10712 -24064 10770 -24052
rect 10712 -24640 10724 -24064
rect 10758 -24640 10770 -24064
rect 10712 -24652 10770 -24640
rect 11730 -24064 11788 -24052
rect 11730 -24640 11742 -24064
rect 11776 -24640 11788 -24064
rect 11730 -24652 11788 -24640
rect 12748 -24064 12806 -24052
rect 12748 -24640 12760 -24064
rect 12794 -24640 12806 -24064
rect 12748 -24652 12806 -24640
rect 13766 -24064 13824 -24052
rect 13766 -24640 13778 -24064
rect 13812 -24640 13824 -24064
rect 13766 -24652 13824 -24640
rect 14784 -24064 14842 -24052
rect 14784 -24640 14796 -24064
rect 14830 -24640 14842 -24064
rect 14784 -24652 14842 -24640
rect 15802 -24064 15860 -24052
rect 15802 -24640 15814 -24064
rect 15848 -24640 15860 -24064
rect 15802 -24652 15860 -24640
rect 16820 -24064 16878 -24052
rect 16820 -24640 16832 -24064
rect 16866 -24640 16878 -24064
rect 16820 -24652 16878 -24640
rect 17838 -24064 17896 -24052
rect 17838 -24640 17850 -24064
rect 17884 -24640 17896 -24064
rect 17838 -24652 17896 -24640
rect 18856 -24064 18914 -24052
rect 18856 -24640 18868 -24064
rect 18902 -24640 18914 -24064
rect 18856 -24652 18914 -24640
rect 19874 -24064 19932 -24052
rect 19874 -24640 19886 -24064
rect 19920 -24640 19932 -24064
rect 19874 -24652 19932 -24640
rect 20892 -24064 20950 -24052
rect 20892 -24640 20904 -24064
rect 20938 -24640 20950 -24064
rect 20892 -24652 20950 -24640
rect 21910 -24064 21968 -24052
rect 21910 -24640 21922 -24064
rect 21956 -24640 21968 -24064
rect 21910 -24652 21968 -24640
rect 22928 -24064 22986 -24052
rect 22928 -24640 22940 -24064
rect 22974 -24640 22986 -24064
rect 22928 -24652 22986 -24640
rect -9418 -25130 -9360 -25118
rect -9418 -25706 -9406 -25130
rect -9372 -25706 -9360 -25130
rect -9418 -25718 -9360 -25706
rect -8400 -25130 -8342 -25118
rect -8400 -25706 -8388 -25130
rect -8354 -25706 -8342 -25130
rect -8400 -25718 -8342 -25706
rect -7382 -25130 -7324 -25118
rect -7382 -25706 -7370 -25130
rect -7336 -25706 -7324 -25130
rect -7382 -25718 -7324 -25706
rect -6364 -25130 -6306 -25118
rect -6364 -25706 -6352 -25130
rect -6318 -25706 -6306 -25130
rect -6364 -25718 -6306 -25706
rect -5346 -25130 -5288 -25118
rect -5346 -25706 -5334 -25130
rect -5300 -25706 -5288 -25130
rect -5346 -25718 -5288 -25706
rect -4328 -25130 -4270 -25118
rect -4328 -25706 -4316 -25130
rect -4282 -25706 -4270 -25130
rect -4328 -25718 -4270 -25706
rect -3310 -25130 -3252 -25118
rect -3310 -25706 -3298 -25130
rect -3264 -25706 -3252 -25130
rect -3310 -25718 -3252 -25706
rect -2424 -25126 -2366 -25114
rect -2424 -25702 -2412 -25126
rect -2378 -25702 -2366 -25126
rect -2424 -25714 -2366 -25702
rect -2126 -25126 -2068 -25114
rect -2126 -25702 -2114 -25126
rect -2080 -25702 -2068 -25126
rect -2126 -25714 -2068 -25702
rect -1828 -25126 -1770 -25114
rect -1828 -25702 -1816 -25126
rect -1782 -25702 -1770 -25126
rect -1828 -25714 -1770 -25702
rect -1530 -25126 -1472 -25114
rect -1530 -25702 -1518 -25126
rect -1484 -25702 -1472 -25126
rect -1530 -25714 -1472 -25702
rect -1232 -25126 -1174 -25114
rect -1232 -25702 -1220 -25126
rect -1186 -25702 -1174 -25126
rect -1232 -25714 -1174 -25702
rect -934 -25126 -876 -25114
rect -934 -25702 -922 -25126
rect -888 -25702 -876 -25126
rect -934 -25714 -876 -25702
rect -636 -25126 -578 -25114
rect -636 -25702 -624 -25126
rect -590 -25702 -578 -25126
rect -636 -25714 -578 -25702
rect -338 -25126 -280 -25114
rect -338 -25702 -326 -25126
rect -292 -25702 -280 -25126
rect -338 -25714 -280 -25702
rect -40 -25126 18 -25114
rect -40 -25702 -28 -25126
rect 6 -25702 18 -25126
rect -40 -25714 18 -25702
rect 258 -25126 316 -25114
rect 258 -25702 270 -25126
rect 304 -25702 316 -25126
rect 258 -25714 316 -25702
rect 556 -25126 614 -25114
rect 556 -25702 568 -25126
rect 602 -25702 614 -25126
rect 556 -25714 614 -25702
rect 854 -25126 912 -25114
rect 854 -25702 866 -25126
rect 900 -25702 912 -25126
rect 854 -25714 912 -25702
rect 2568 -25296 2626 -25284
rect 2568 -25872 2580 -25296
rect 2614 -25872 2626 -25296
rect 2568 -25884 2626 -25872
rect 3586 -25296 3644 -25284
rect 3586 -25872 3598 -25296
rect 3632 -25872 3644 -25296
rect 3586 -25884 3644 -25872
rect 4604 -25296 4662 -25284
rect 4604 -25872 4616 -25296
rect 4650 -25872 4662 -25296
rect 4604 -25884 4662 -25872
rect 5622 -25296 5680 -25284
rect 5622 -25872 5634 -25296
rect 5668 -25872 5680 -25296
rect 5622 -25884 5680 -25872
rect 6640 -25296 6698 -25284
rect 6640 -25872 6652 -25296
rect 6686 -25872 6698 -25296
rect 6640 -25884 6698 -25872
rect 7658 -25296 7716 -25284
rect 7658 -25872 7670 -25296
rect 7704 -25872 7716 -25296
rect 7658 -25884 7716 -25872
rect 8676 -25296 8734 -25284
rect 8676 -25872 8688 -25296
rect 8722 -25872 8734 -25296
rect 8676 -25884 8734 -25872
rect 9694 -25296 9752 -25284
rect 9694 -25872 9706 -25296
rect 9740 -25872 9752 -25296
rect 9694 -25884 9752 -25872
rect 10712 -25296 10770 -25284
rect 10712 -25872 10724 -25296
rect 10758 -25872 10770 -25296
rect 10712 -25884 10770 -25872
rect 11730 -25296 11788 -25284
rect 11730 -25872 11742 -25296
rect 11776 -25872 11788 -25296
rect 11730 -25884 11788 -25872
rect 12748 -25296 12806 -25284
rect 12748 -25872 12760 -25296
rect 12794 -25872 12806 -25296
rect 12748 -25884 12806 -25872
rect 13766 -25296 13824 -25284
rect 13766 -25872 13778 -25296
rect 13812 -25872 13824 -25296
rect 13766 -25884 13824 -25872
rect 14784 -25296 14842 -25284
rect 14784 -25872 14796 -25296
rect 14830 -25872 14842 -25296
rect 14784 -25884 14842 -25872
rect 15802 -25296 15860 -25284
rect 15802 -25872 15814 -25296
rect 15848 -25872 15860 -25296
rect 15802 -25884 15860 -25872
rect 16820 -25296 16878 -25284
rect 16820 -25872 16832 -25296
rect 16866 -25872 16878 -25296
rect 16820 -25884 16878 -25872
rect 17838 -25296 17896 -25284
rect 17838 -25872 17850 -25296
rect 17884 -25872 17896 -25296
rect 17838 -25884 17896 -25872
rect 18856 -25296 18914 -25284
rect 18856 -25872 18868 -25296
rect 18902 -25872 18914 -25296
rect 18856 -25884 18914 -25872
rect 19874 -25296 19932 -25284
rect 19874 -25872 19886 -25296
rect 19920 -25872 19932 -25296
rect 19874 -25884 19932 -25872
rect 20892 -25296 20950 -25284
rect 20892 -25872 20904 -25296
rect 20938 -25872 20950 -25296
rect 20892 -25884 20950 -25872
rect 21910 -25296 21968 -25284
rect 21910 -25872 21922 -25296
rect 21956 -25872 21968 -25296
rect 21910 -25884 21968 -25872
rect 22928 -25296 22986 -25284
rect 22928 -25872 22940 -25296
rect 22974 -25872 22986 -25296
rect 22928 -25884 22986 -25872
<< pdiff >>
rect 3614 -4702 3672 -4690
rect 3614 -5078 3626 -4702
rect 3660 -5078 3672 -4702
rect 3614 -5090 3672 -5078
rect 3832 -4702 3890 -4690
rect 3832 -5078 3844 -4702
rect 3878 -5078 3890 -4702
rect 3832 -5090 3890 -5078
rect 4050 -4702 4108 -4690
rect 4050 -5078 4062 -4702
rect 4096 -5078 4108 -4702
rect 4050 -5090 4108 -5078
rect 4268 -4702 4326 -4690
rect 4268 -5078 4280 -4702
rect 4314 -5078 4326 -4702
rect 4268 -5090 4326 -5078
rect 4486 -4702 4544 -4690
rect 4486 -5078 4498 -4702
rect 4532 -5078 4544 -4702
rect 4486 -5090 4544 -5078
rect 4704 -4702 4762 -4690
rect 4704 -5078 4716 -4702
rect 4750 -5078 4762 -4702
rect 4704 -5090 4762 -5078
rect 4922 -4702 4980 -4690
rect 4922 -5078 4934 -4702
rect 4968 -5078 4980 -4702
rect 4922 -5090 4980 -5078
rect 5140 -4702 5198 -4690
rect 5140 -5078 5152 -4702
rect 5186 -5078 5198 -4702
rect 5140 -5090 5198 -5078
rect 5358 -4702 5416 -4690
rect 5358 -5078 5370 -4702
rect 5404 -5078 5416 -4702
rect 5358 -5090 5416 -5078
rect 5576 -4702 5634 -4690
rect 5576 -5078 5588 -4702
rect 5622 -5078 5634 -4702
rect 5576 -5090 5634 -5078
rect 5794 -4702 5852 -4690
rect 5794 -5078 5806 -4702
rect 5840 -5078 5852 -4702
rect 5794 -5090 5852 -5078
rect 3614 -5640 3672 -5628
rect 3614 -6016 3626 -5640
rect 3660 -6016 3672 -5640
rect 3614 -6028 3672 -6016
rect 3832 -5640 3890 -5628
rect 3832 -6016 3844 -5640
rect 3878 -6016 3890 -5640
rect 3832 -6028 3890 -6016
rect 4050 -5640 4108 -5628
rect 4050 -6016 4062 -5640
rect 4096 -6016 4108 -5640
rect 4050 -6028 4108 -6016
rect 4268 -5640 4326 -5628
rect 4268 -6016 4280 -5640
rect 4314 -6016 4326 -5640
rect 4268 -6028 4326 -6016
rect 4486 -5640 4544 -5628
rect 4486 -6016 4498 -5640
rect 4532 -6016 4544 -5640
rect 4486 -6028 4544 -6016
rect 4704 -5640 4762 -5628
rect 4704 -6016 4716 -5640
rect 4750 -6016 4762 -5640
rect 4704 -6028 4762 -6016
rect 4922 -5640 4980 -5628
rect 4922 -6016 4934 -5640
rect 4968 -6016 4980 -5640
rect 4922 -6028 4980 -6016
rect 5140 -5640 5198 -5628
rect 5140 -6016 5152 -5640
rect 5186 -6016 5198 -5640
rect 5140 -6028 5198 -6016
rect 5358 -5640 5416 -5628
rect 5358 -6016 5370 -5640
rect 5404 -6016 5416 -5640
rect 5358 -6028 5416 -6016
rect 5576 -5640 5634 -5628
rect 5576 -6016 5588 -5640
rect 5622 -6016 5634 -5640
rect 5576 -6028 5634 -6016
rect 5794 -5640 5852 -5628
rect 5794 -6016 5806 -5640
rect 5840 -6016 5852 -5640
rect 5794 -6028 5852 -6016
rect 3614 -6578 3672 -6566
rect 3614 -6954 3626 -6578
rect 3660 -6954 3672 -6578
rect 3614 -6966 3672 -6954
rect 3832 -6578 3890 -6566
rect 3832 -6954 3844 -6578
rect 3878 -6954 3890 -6578
rect 3832 -6966 3890 -6954
rect 4050 -6578 4108 -6566
rect 4050 -6954 4062 -6578
rect 4096 -6954 4108 -6578
rect 4050 -6966 4108 -6954
rect 4268 -6578 4326 -6566
rect 4268 -6954 4280 -6578
rect 4314 -6954 4326 -6578
rect 4268 -6966 4326 -6954
rect 4486 -6578 4544 -6566
rect 4486 -6954 4498 -6578
rect 4532 -6954 4544 -6578
rect 4486 -6966 4544 -6954
rect 4704 -6578 4762 -6566
rect 4704 -6954 4716 -6578
rect 4750 -6954 4762 -6578
rect 4704 -6966 4762 -6954
rect 4922 -6578 4980 -6566
rect 4922 -6954 4934 -6578
rect 4968 -6954 4980 -6578
rect 4922 -6966 4980 -6954
rect 5140 -6578 5198 -6566
rect 5140 -6954 5152 -6578
rect 5186 -6954 5198 -6578
rect 5140 -6966 5198 -6954
rect 5358 -6578 5416 -6566
rect 5358 -6954 5370 -6578
rect 5404 -6954 5416 -6578
rect 5358 -6966 5416 -6954
rect 5576 -6578 5634 -6566
rect 5576 -6954 5588 -6578
rect 5622 -6954 5634 -6578
rect 5576 -6966 5634 -6954
rect 5794 -6578 5852 -6566
rect 5794 -6954 5806 -6578
rect 5840 -6954 5852 -6578
rect 5794 -6966 5852 -6954
rect 3614 -7516 3672 -7504
rect 3614 -7892 3626 -7516
rect 3660 -7892 3672 -7516
rect 3614 -7904 3672 -7892
rect 3832 -7516 3890 -7504
rect 3832 -7892 3844 -7516
rect 3878 -7892 3890 -7516
rect 3832 -7904 3890 -7892
rect 4050 -7516 4108 -7504
rect 4050 -7892 4062 -7516
rect 4096 -7892 4108 -7516
rect 4050 -7904 4108 -7892
rect 4268 -7516 4326 -7504
rect 4268 -7892 4280 -7516
rect 4314 -7892 4326 -7516
rect 4268 -7904 4326 -7892
rect 4486 -7516 4544 -7504
rect 4486 -7892 4498 -7516
rect 4532 -7892 4544 -7516
rect 4486 -7904 4544 -7892
rect 4704 -7516 4762 -7504
rect 4704 -7892 4716 -7516
rect 4750 -7892 4762 -7516
rect 4704 -7904 4762 -7892
rect 4922 -7516 4980 -7504
rect 4922 -7892 4934 -7516
rect 4968 -7892 4980 -7516
rect 4922 -7904 4980 -7892
rect 5140 -7516 5198 -7504
rect 5140 -7892 5152 -7516
rect 5186 -7892 5198 -7516
rect 5140 -7904 5198 -7892
rect 5358 -7516 5416 -7504
rect 5358 -7892 5370 -7516
rect 5404 -7892 5416 -7516
rect 5358 -7904 5416 -7892
rect 5576 -7516 5634 -7504
rect 5576 -7892 5588 -7516
rect 5622 -7892 5634 -7516
rect 5576 -7904 5634 -7892
rect 5794 -7516 5852 -7504
rect 5794 -7892 5806 -7516
rect 5840 -7892 5852 -7516
rect 5794 -7904 5852 -7892
<< ndiffc >>
rect 2582 -12306 2616 -11730
rect 3600 -12306 3634 -11730
rect 4618 -12306 4652 -11730
rect 5636 -12306 5670 -11730
rect 6654 -12306 6688 -11730
rect 7672 -12306 7706 -11730
rect 8690 -12306 8724 -11730
rect 9708 -12306 9742 -11730
rect 10726 -12306 10760 -11730
rect 11744 -12306 11778 -11730
rect 12762 -12306 12796 -11730
rect 13780 -12306 13814 -11730
rect 14798 -12306 14832 -11730
rect 15816 -12306 15850 -11730
rect 16834 -12306 16868 -11730
rect 17852 -12306 17886 -11730
rect 18870 -12306 18904 -11730
rect 19888 -12306 19922 -11730
rect 20906 -12306 20940 -11730
rect 21924 -12306 21958 -11730
rect 22942 -12306 22976 -11730
rect -9184 -13100 -9150 -12524
rect -8166 -13100 -8132 -12524
rect -7148 -13100 -7114 -12524
rect -6130 -13100 -6096 -12524
rect -5112 -13100 -5078 -12524
rect -4094 -13100 -4060 -12524
rect -3076 -13100 -3042 -12524
rect -2058 -13100 -2024 -12524
rect -1040 -13100 -1006 -12524
rect -22 -13100 12 -12524
rect -9184 -13918 -9150 -13342
rect -8166 -13918 -8132 -13342
rect -7148 -13918 -7114 -13342
rect -6130 -13918 -6096 -13342
rect -5112 -13918 -5078 -13342
rect -4094 -13918 -4060 -13342
rect -3076 -13918 -3042 -13342
rect -2058 -13918 -2024 -13342
rect -1040 -13918 -1006 -13342
rect -22 -13918 12 -13342
rect 2582 -13540 2616 -12964
rect 3600 -13540 3634 -12964
rect 4618 -13540 4652 -12964
rect 5636 -13540 5670 -12964
rect 6654 -13540 6688 -12964
rect 7672 -13540 7706 -12964
rect 8690 -13540 8724 -12964
rect 9708 -13540 9742 -12964
rect 10726 -13540 10760 -12964
rect 11744 -13540 11778 -12964
rect 12762 -13540 12796 -12964
rect 13780 -13540 13814 -12964
rect 14798 -13540 14832 -12964
rect 15816 -13540 15850 -12964
rect 16834 -13540 16868 -12964
rect 17852 -13540 17886 -12964
rect 18870 -13540 18904 -12964
rect 19888 -13540 19922 -12964
rect 20906 -13540 20940 -12964
rect 21924 -13540 21958 -12964
rect 22942 -13540 22976 -12964
rect -9184 -14736 -9150 -14160
rect -8166 -14736 -8132 -14160
rect -7148 -14736 -7114 -14160
rect -6130 -14736 -6096 -14160
rect -5112 -14736 -5078 -14160
rect -4094 -14736 -4060 -14160
rect -3076 -14736 -3042 -14160
rect -2058 -14736 -2024 -14160
rect -1040 -14736 -1006 -14160
rect -22 -14736 12 -14160
rect 2582 -14772 2616 -14196
rect 3600 -14772 3634 -14196
rect 4618 -14772 4652 -14196
rect 5636 -14772 5670 -14196
rect 6654 -14772 6688 -14196
rect 7672 -14772 7706 -14196
rect 8690 -14772 8724 -14196
rect 9708 -14772 9742 -14196
rect 10726 -14772 10760 -14196
rect 11744 -14772 11778 -14196
rect 12762 -14772 12796 -14196
rect 13780 -14772 13814 -14196
rect 14798 -14772 14832 -14196
rect 15816 -14772 15850 -14196
rect 16834 -14772 16868 -14196
rect 17852 -14772 17886 -14196
rect 18870 -14772 18904 -14196
rect 19888 -14772 19922 -14196
rect 20906 -14772 20940 -14196
rect 21924 -14772 21958 -14196
rect 22942 -14772 22976 -14196
rect -9184 -15554 -9150 -14978
rect -8166 -15554 -8132 -14978
rect -7148 -15554 -7114 -14978
rect -6130 -15554 -6096 -14978
rect -5112 -15554 -5078 -14978
rect -4094 -15554 -4060 -14978
rect -3076 -15554 -3042 -14978
rect -2058 -15554 -2024 -14978
rect -1040 -15554 -1006 -14978
rect -22 -15554 12 -14978
rect -9184 -16372 -9150 -15796
rect -8166 -16372 -8132 -15796
rect -7148 -16372 -7114 -15796
rect -6130 -16372 -6096 -15796
rect -5112 -16372 -5078 -15796
rect -4094 -16372 -4060 -15796
rect -3076 -16372 -3042 -15796
rect -2058 -16372 -2024 -15796
rect -1040 -16372 -1006 -15796
rect -22 -16372 12 -15796
rect 2580 -16006 2614 -15430
rect 3598 -16006 3632 -15430
rect 4616 -16006 4650 -15430
rect 5634 -16006 5668 -15430
rect 6652 -16006 6686 -15430
rect 7670 -16006 7704 -15430
rect 8688 -16006 8722 -15430
rect 9706 -16006 9740 -15430
rect 10724 -16006 10758 -15430
rect 11742 -16006 11776 -15430
rect 12760 -16006 12794 -15430
rect 13778 -16006 13812 -15430
rect 14796 -16006 14830 -15430
rect 15814 -16006 15848 -15430
rect 16832 -16006 16866 -15430
rect 17850 -16006 17884 -15430
rect 18868 -16006 18902 -15430
rect 19886 -16006 19920 -15430
rect 20904 -16006 20938 -15430
rect 21922 -16006 21956 -15430
rect 22940 -16006 22974 -15430
rect -9184 -17190 -9150 -16614
rect -8166 -17190 -8132 -16614
rect -7148 -17190 -7114 -16614
rect -6130 -17190 -6096 -16614
rect -5112 -17190 -5078 -16614
rect -4094 -17190 -4060 -16614
rect -3076 -17190 -3042 -16614
rect -2058 -17190 -2024 -16614
rect -1040 -17190 -1006 -16614
rect -22 -17190 12 -16614
rect 2580 -17240 2614 -16664
rect 3598 -17240 3632 -16664
rect 4616 -17240 4650 -16664
rect 5634 -17240 5668 -16664
rect 6652 -17240 6686 -16664
rect 7670 -17240 7704 -16664
rect 8688 -17240 8722 -16664
rect 9706 -17240 9740 -16664
rect 10724 -17240 10758 -16664
rect 11742 -17240 11776 -16664
rect 12760 -17240 12794 -16664
rect 13778 -17240 13812 -16664
rect 14796 -17240 14830 -16664
rect 15814 -17240 15848 -16664
rect 16832 -17240 16866 -16664
rect 17850 -17240 17884 -16664
rect 18868 -17240 18902 -16664
rect 19886 -17240 19920 -16664
rect 20904 -17240 20938 -16664
rect 21922 -17240 21956 -16664
rect 22940 -17240 22974 -16664
rect -9184 -18008 -9150 -17432
rect -8166 -18008 -8132 -17432
rect -7148 -18008 -7114 -17432
rect -6130 -18008 -6096 -17432
rect -5112 -18008 -5078 -17432
rect -4094 -18008 -4060 -17432
rect -3076 -18008 -3042 -17432
rect -2058 -18008 -2024 -17432
rect -1040 -18008 -1006 -17432
rect -22 -18008 12 -17432
rect -9184 -18826 -9150 -18250
rect -8166 -18826 -8132 -18250
rect -7148 -18826 -7114 -18250
rect -6130 -18826 -6096 -18250
rect -5112 -18826 -5078 -18250
rect -4094 -18826 -4060 -18250
rect -3076 -18826 -3042 -18250
rect -2058 -18826 -2024 -18250
rect -1040 -18826 -1006 -18250
rect -22 -18826 12 -18250
rect 2580 -18472 2614 -17896
rect 3598 -18472 3632 -17896
rect 4616 -18472 4650 -17896
rect 5634 -18472 5668 -17896
rect 6652 -18472 6686 -17896
rect 7670 -18472 7704 -17896
rect 8688 -18472 8722 -17896
rect 9706 -18472 9740 -17896
rect 10724 -18472 10758 -17896
rect 11742 -18472 11776 -17896
rect 12760 -18472 12794 -17896
rect 13778 -18472 13812 -17896
rect 14796 -18472 14830 -17896
rect 15814 -18472 15848 -17896
rect 16832 -18472 16866 -17896
rect 17850 -18472 17884 -17896
rect 18868 -18472 18902 -17896
rect 19886 -18472 19920 -17896
rect 20904 -18472 20938 -17896
rect 21922 -18472 21956 -17896
rect 22940 -18472 22974 -17896
rect -2324 -19810 -2290 -19634
rect -2106 -19810 -2072 -19634
rect -1888 -19810 -1854 -19634
rect -1670 -19810 -1636 -19634
rect -1452 -19810 -1418 -19634
rect -1234 -19810 -1200 -19634
rect -1016 -19810 -982 -19634
rect -798 -19810 -764 -19634
rect -580 -19810 -546 -19634
rect -362 -19810 -328 -19634
rect -144 -19810 -110 -19634
rect 2580 -19706 2614 -19130
rect 3598 -19706 3632 -19130
rect 4616 -19706 4650 -19130
rect 5634 -19706 5668 -19130
rect 6652 -19706 6686 -19130
rect 7670 -19706 7704 -19130
rect 8688 -19706 8722 -19130
rect 9706 -19706 9740 -19130
rect 10724 -19706 10758 -19130
rect 11742 -19706 11776 -19130
rect 12760 -19706 12794 -19130
rect 13778 -19706 13812 -19130
rect 14796 -19706 14830 -19130
rect 15814 -19706 15848 -19130
rect 16832 -19706 16866 -19130
rect 17850 -19706 17884 -19130
rect 18868 -19706 18902 -19130
rect 19886 -19706 19920 -19130
rect 20904 -19706 20938 -19130
rect 21922 -19706 21956 -19130
rect 22940 -19706 22974 -19130
rect -2324 -20642 -2290 -20466
rect -2106 -20642 -2072 -20466
rect -1888 -20642 -1854 -20466
rect -1670 -20642 -1636 -20466
rect -1452 -20642 -1418 -20466
rect -1234 -20642 -1200 -20466
rect -1016 -20642 -982 -20466
rect -798 -20642 -764 -20466
rect -580 -20642 -546 -20466
rect -362 -20642 -328 -20466
rect -144 -20642 -110 -20466
rect 2580 -20940 2614 -20364
rect 3598 -20940 3632 -20364
rect 4616 -20940 4650 -20364
rect 5634 -20940 5668 -20364
rect 6652 -20940 6686 -20364
rect 7670 -20940 7704 -20364
rect 8688 -20940 8722 -20364
rect 9706 -20940 9740 -20364
rect 10724 -20940 10758 -20364
rect 11742 -20940 11776 -20364
rect 12760 -20940 12794 -20364
rect 13778 -20940 13812 -20364
rect 14796 -20940 14830 -20364
rect 15814 -20940 15848 -20364
rect 16832 -20940 16866 -20364
rect 17850 -20940 17884 -20364
rect 18868 -20940 18902 -20364
rect 19886 -20940 19920 -20364
rect 20904 -20940 20938 -20364
rect 21922 -20940 21956 -20364
rect 22940 -20940 22974 -20364
rect -9405 -22369 -9371 -21793
rect -8387 -22369 -8353 -21793
rect -7369 -22369 -7335 -21793
rect -6351 -22369 -6317 -21793
rect -5333 -22369 -5299 -21793
rect -4315 -22369 -4281 -21793
rect -3297 -22369 -3263 -21793
rect -2410 -22368 -2376 -21792
rect -2112 -22368 -2078 -21792
rect -1814 -22368 -1780 -21792
rect -1516 -22368 -1482 -21792
rect -1218 -22368 -1184 -21792
rect -920 -22368 -886 -21792
rect -622 -22368 -588 -21792
rect -324 -22368 -290 -21792
rect -26 -22368 8 -21792
rect 272 -22368 306 -21792
rect 570 -22368 604 -21792
rect 868 -22368 902 -21792
rect 2580 -22172 2614 -21596
rect 3598 -22172 3632 -21596
rect 4616 -22172 4650 -21596
rect 5634 -22172 5668 -21596
rect 6652 -22172 6686 -21596
rect 7670 -22172 7704 -21596
rect 8688 -22172 8722 -21596
rect 9706 -22172 9740 -21596
rect 10724 -22172 10758 -21596
rect 11742 -22172 11776 -21596
rect 12760 -22172 12794 -21596
rect 13778 -22172 13812 -21596
rect 14796 -22172 14830 -21596
rect 15814 -22172 15848 -21596
rect 16832 -22172 16866 -21596
rect 17850 -22172 17884 -21596
rect 18868 -22172 18902 -21596
rect 19886 -22172 19920 -21596
rect 20904 -22172 20938 -21596
rect 21922 -22172 21956 -21596
rect 22940 -22172 22974 -21596
rect -9406 -23482 -9372 -22906
rect -8388 -23482 -8354 -22906
rect -7370 -23482 -7336 -22906
rect -6352 -23482 -6318 -22906
rect -5334 -23482 -5300 -22906
rect -4316 -23482 -4282 -22906
rect -3298 -23482 -3264 -22906
rect -2410 -23480 -2376 -22904
rect -2112 -23480 -2078 -22904
rect -1814 -23480 -1780 -22904
rect -1516 -23480 -1482 -22904
rect -1218 -23480 -1184 -22904
rect -920 -23480 -886 -22904
rect -622 -23480 -588 -22904
rect -324 -23480 -290 -22904
rect -26 -23480 8 -22904
rect 272 -23480 306 -22904
rect 570 -23480 604 -22904
rect 868 -23480 902 -22904
rect 2580 -23406 2614 -22830
rect 3598 -23406 3632 -22830
rect 4616 -23406 4650 -22830
rect 5634 -23406 5668 -22830
rect 6652 -23406 6686 -22830
rect 7670 -23406 7704 -22830
rect 8688 -23406 8722 -22830
rect 9706 -23406 9740 -22830
rect 10724 -23406 10758 -22830
rect 11742 -23406 11776 -22830
rect 12760 -23406 12794 -22830
rect 13778 -23406 13812 -22830
rect 14796 -23406 14830 -22830
rect 15814 -23406 15848 -22830
rect 16832 -23406 16866 -22830
rect 17850 -23406 17884 -22830
rect 18868 -23406 18902 -22830
rect 19886 -23406 19920 -22830
rect 20904 -23406 20938 -22830
rect 21922 -23406 21956 -22830
rect 22940 -23406 22974 -22830
rect -9405 -24593 -9371 -24017
rect -8387 -24593 -8353 -24017
rect -7369 -24593 -7335 -24017
rect -6351 -24593 -6317 -24017
rect -5333 -24593 -5299 -24017
rect -4315 -24593 -4281 -24017
rect -3297 -24593 -3263 -24017
rect -2412 -24592 -2378 -24016
rect -2114 -24592 -2080 -24016
rect -1816 -24592 -1782 -24016
rect -1518 -24592 -1484 -24016
rect -1220 -24592 -1186 -24016
rect -922 -24592 -888 -24016
rect -624 -24592 -590 -24016
rect -326 -24592 -292 -24016
rect -28 -24592 6 -24016
rect 270 -24592 304 -24016
rect 568 -24592 602 -24016
rect 866 -24592 900 -24016
rect 2580 -24640 2614 -24064
rect 3598 -24640 3632 -24064
rect 4616 -24640 4650 -24064
rect 5634 -24640 5668 -24064
rect 6652 -24640 6686 -24064
rect 7670 -24640 7704 -24064
rect 8688 -24640 8722 -24064
rect 9706 -24640 9740 -24064
rect 10724 -24640 10758 -24064
rect 11742 -24640 11776 -24064
rect 12760 -24640 12794 -24064
rect 13778 -24640 13812 -24064
rect 14796 -24640 14830 -24064
rect 15814 -24640 15848 -24064
rect 16832 -24640 16866 -24064
rect 17850 -24640 17884 -24064
rect 18868 -24640 18902 -24064
rect 19886 -24640 19920 -24064
rect 20904 -24640 20938 -24064
rect 21922 -24640 21956 -24064
rect 22940 -24640 22974 -24064
rect -9406 -25706 -9372 -25130
rect -8388 -25706 -8354 -25130
rect -7370 -25706 -7336 -25130
rect -6352 -25706 -6318 -25130
rect -5334 -25706 -5300 -25130
rect -4316 -25706 -4282 -25130
rect -3298 -25706 -3264 -25130
rect -2412 -25702 -2378 -25126
rect -2114 -25702 -2080 -25126
rect -1816 -25702 -1782 -25126
rect -1518 -25702 -1484 -25126
rect -1220 -25702 -1186 -25126
rect -922 -25702 -888 -25126
rect -624 -25702 -590 -25126
rect -326 -25702 -292 -25126
rect -28 -25702 6 -25126
rect 270 -25702 304 -25126
rect 568 -25702 602 -25126
rect 866 -25702 900 -25126
rect 2580 -25872 2614 -25296
rect 3598 -25872 3632 -25296
rect 4616 -25872 4650 -25296
rect 5634 -25872 5668 -25296
rect 6652 -25872 6686 -25296
rect 7670 -25872 7704 -25296
rect 8688 -25872 8722 -25296
rect 9706 -25872 9740 -25296
rect 10724 -25872 10758 -25296
rect 11742 -25872 11776 -25296
rect 12760 -25872 12794 -25296
rect 13778 -25872 13812 -25296
rect 14796 -25872 14830 -25296
rect 15814 -25872 15848 -25296
rect 16832 -25872 16866 -25296
rect 17850 -25872 17884 -25296
rect 18868 -25872 18902 -25296
rect 19886 -25872 19920 -25296
rect 20904 -25872 20938 -25296
rect 21922 -25872 21956 -25296
rect 22940 -25872 22974 -25296
<< pdiffc >>
rect 3626 -5078 3660 -4702
rect 3844 -5078 3878 -4702
rect 4062 -5078 4096 -4702
rect 4280 -5078 4314 -4702
rect 4498 -5078 4532 -4702
rect 4716 -5078 4750 -4702
rect 4934 -5078 4968 -4702
rect 5152 -5078 5186 -4702
rect 5370 -5078 5404 -4702
rect 5588 -5078 5622 -4702
rect 5806 -5078 5840 -4702
rect 3626 -6016 3660 -5640
rect 3844 -6016 3878 -5640
rect 4062 -6016 4096 -5640
rect 4280 -6016 4314 -5640
rect 4498 -6016 4532 -5640
rect 4716 -6016 4750 -5640
rect 4934 -6016 4968 -5640
rect 5152 -6016 5186 -5640
rect 5370 -6016 5404 -5640
rect 5588 -6016 5622 -5640
rect 5806 -6016 5840 -5640
rect 3626 -6954 3660 -6578
rect 3844 -6954 3878 -6578
rect 4062 -6954 4096 -6578
rect 4280 -6954 4314 -6578
rect 4498 -6954 4532 -6578
rect 4716 -6954 4750 -6578
rect 4934 -6954 4968 -6578
rect 5152 -6954 5186 -6578
rect 5370 -6954 5404 -6578
rect 5588 -6954 5622 -6578
rect 5806 -6954 5840 -6578
rect 3626 -7892 3660 -7516
rect 3844 -7892 3878 -7516
rect 4062 -7892 4096 -7516
rect 4280 -7892 4314 -7516
rect 4498 -7892 4532 -7516
rect 4716 -7892 4750 -7516
rect 4934 -7892 4968 -7516
rect 5152 -7892 5186 -7516
rect 5370 -7892 5404 -7516
rect 5588 -7892 5622 -7516
rect 5806 -7892 5840 -7516
<< psubdiff >>
rect -12322 -11278 -12160 -11178
rect 24760 -11278 24922 -11178
rect -12322 -11340 -12222 -11278
rect 24822 -11340 24922 -11278
rect -12322 -27122 -12222 -27060
rect 24822 -27122 24922 -27060
rect -12322 -27222 -12160 -27122
rect 24760 -27222 24922 -27122
<< nsubdiff >>
rect 378 1622 540 1722
rect 24660 1622 24822 1722
rect 378 1560 478 1622
rect 24722 1560 24822 1622
rect 378 -8782 478 -8720
rect 24722 -8782 24822 -8720
rect 378 -8882 540 -8782
rect 24660 -8882 24822 -8782
<< psubdiffcont >>
rect -12160 -11278 24760 -11178
rect -12322 -27060 -12222 -11340
rect 24822 -27060 24922 -11340
rect -12160 -27222 24760 -27122
<< nsubdiffcont >>
rect 540 1622 24660 1722
rect 378 -8720 478 1560
rect 24722 -8720 24822 1560
rect 540 -8882 24660 -8782
<< poly >>
rect 3698 -4609 3806 -4593
rect 3698 -4626 3714 -4609
rect 3672 -4643 3714 -4626
rect 3790 -4626 3806 -4609
rect 3916 -4609 4024 -4593
rect 3916 -4626 3932 -4609
rect 3790 -4643 3832 -4626
rect 3672 -4690 3832 -4643
rect 3890 -4643 3932 -4626
rect 4008 -4626 4024 -4609
rect 4134 -4609 4242 -4593
rect 4134 -4626 4150 -4609
rect 4008 -4643 4050 -4626
rect 3890 -4690 4050 -4643
rect 4108 -4643 4150 -4626
rect 4226 -4626 4242 -4609
rect 4352 -4609 4460 -4593
rect 4352 -4626 4368 -4609
rect 4226 -4643 4268 -4626
rect 4108 -4690 4268 -4643
rect 4326 -4643 4368 -4626
rect 4444 -4626 4460 -4609
rect 4570 -4609 4678 -4593
rect 4570 -4626 4586 -4609
rect 4444 -4643 4486 -4626
rect 4326 -4690 4486 -4643
rect 4544 -4643 4586 -4626
rect 4662 -4626 4678 -4609
rect 4788 -4609 4896 -4593
rect 4788 -4626 4804 -4609
rect 4662 -4643 4704 -4626
rect 4544 -4690 4704 -4643
rect 4762 -4643 4804 -4626
rect 4880 -4626 4896 -4609
rect 5006 -4609 5114 -4593
rect 5006 -4626 5022 -4609
rect 4880 -4643 4922 -4626
rect 4762 -4690 4922 -4643
rect 4980 -4643 5022 -4626
rect 5098 -4626 5114 -4609
rect 5224 -4609 5332 -4593
rect 5224 -4626 5240 -4609
rect 5098 -4643 5140 -4626
rect 4980 -4690 5140 -4643
rect 5198 -4643 5240 -4626
rect 5316 -4626 5332 -4609
rect 5442 -4609 5550 -4593
rect 5442 -4626 5458 -4609
rect 5316 -4643 5358 -4626
rect 5198 -4690 5358 -4643
rect 5416 -4643 5458 -4626
rect 5534 -4626 5550 -4609
rect 5660 -4609 5768 -4593
rect 5660 -4626 5676 -4609
rect 5534 -4643 5576 -4626
rect 5416 -4690 5576 -4643
rect 5634 -4643 5676 -4626
rect 5752 -4626 5768 -4609
rect 5752 -4643 5794 -4626
rect 5634 -4690 5794 -4643
rect 3672 -5137 3832 -5090
rect 3672 -5154 3714 -5137
rect 3698 -5171 3714 -5154
rect 3790 -5154 3832 -5137
rect 3890 -5137 4050 -5090
rect 3890 -5154 3932 -5137
rect 3790 -5171 3806 -5154
rect 3698 -5187 3806 -5171
rect 3916 -5171 3932 -5154
rect 4008 -5154 4050 -5137
rect 4108 -5137 4268 -5090
rect 4108 -5154 4150 -5137
rect 4008 -5171 4024 -5154
rect 3916 -5187 4024 -5171
rect 4134 -5171 4150 -5154
rect 4226 -5154 4268 -5137
rect 4326 -5137 4486 -5090
rect 4326 -5154 4368 -5137
rect 4226 -5171 4242 -5154
rect 4134 -5187 4242 -5171
rect 4352 -5171 4368 -5154
rect 4444 -5154 4486 -5137
rect 4544 -5137 4704 -5090
rect 4544 -5154 4586 -5137
rect 4444 -5171 4460 -5154
rect 4352 -5187 4460 -5171
rect 4570 -5171 4586 -5154
rect 4662 -5154 4704 -5137
rect 4762 -5137 4922 -5090
rect 4762 -5154 4804 -5137
rect 4662 -5171 4678 -5154
rect 4570 -5187 4678 -5171
rect 4788 -5171 4804 -5154
rect 4880 -5154 4922 -5137
rect 4980 -5137 5140 -5090
rect 4980 -5154 5022 -5137
rect 4880 -5171 4896 -5154
rect 4788 -5187 4896 -5171
rect 5006 -5171 5022 -5154
rect 5098 -5154 5140 -5137
rect 5198 -5137 5358 -5090
rect 5198 -5154 5240 -5137
rect 5098 -5171 5114 -5154
rect 5006 -5187 5114 -5171
rect 5224 -5171 5240 -5154
rect 5316 -5154 5358 -5137
rect 5416 -5137 5576 -5090
rect 5416 -5154 5458 -5137
rect 5316 -5171 5332 -5154
rect 5224 -5187 5332 -5171
rect 5442 -5171 5458 -5154
rect 5534 -5154 5576 -5137
rect 5634 -5137 5794 -5090
rect 5634 -5154 5676 -5137
rect 5534 -5171 5550 -5154
rect 5442 -5187 5550 -5171
rect 5660 -5171 5676 -5154
rect 5752 -5154 5794 -5137
rect 5752 -5171 5768 -5154
rect 5660 -5187 5768 -5171
rect 3698 -5547 3806 -5531
rect 3698 -5564 3714 -5547
rect 3672 -5581 3714 -5564
rect 3790 -5564 3806 -5547
rect 3916 -5547 4024 -5531
rect 3916 -5564 3932 -5547
rect 3790 -5581 3832 -5564
rect 3672 -5628 3832 -5581
rect 3890 -5581 3932 -5564
rect 4008 -5564 4024 -5547
rect 4134 -5547 4242 -5531
rect 4134 -5564 4150 -5547
rect 4008 -5581 4050 -5564
rect 3890 -5628 4050 -5581
rect 4108 -5581 4150 -5564
rect 4226 -5564 4242 -5547
rect 4352 -5547 4460 -5531
rect 4352 -5564 4368 -5547
rect 4226 -5581 4268 -5564
rect 4108 -5628 4268 -5581
rect 4326 -5581 4368 -5564
rect 4444 -5564 4460 -5547
rect 4570 -5547 4678 -5531
rect 4570 -5564 4586 -5547
rect 4444 -5581 4486 -5564
rect 4326 -5628 4486 -5581
rect 4544 -5581 4586 -5564
rect 4662 -5564 4678 -5547
rect 4788 -5547 4896 -5531
rect 4788 -5564 4804 -5547
rect 4662 -5581 4704 -5564
rect 4544 -5628 4704 -5581
rect 4762 -5581 4804 -5564
rect 4880 -5564 4896 -5547
rect 5006 -5547 5114 -5531
rect 5006 -5564 5022 -5547
rect 4880 -5581 4922 -5564
rect 4762 -5628 4922 -5581
rect 4980 -5581 5022 -5564
rect 5098 -5564 5114 -5547
rect 5224 -5547 5332 -5531
rect 5224 -5564 5240 -5547
rect 5098 -5581 5140 -5564
rect 4980 -5628 5140 -5581
rect 5198 -5581 5240 -5564
rect 5316 -5564 5332 -5547
rect 5442 -5547 5550 -5531
rect 5442 -5564 5458 -5547
rect 5316 -5581 5358 -5564
rect 5198 -5628 5358 -5581
rect 5416 -5581 5458 -5564
rect 5534 -5564 5550 -5547
rect 5660 -5547 5768 -5531
rect 5660 -5564 5676 -5547
rect 5534 -5581 5576 -5564
rect 5416 -5628 5576 -5581
rect 5634 -5581 5676 -5564
rect 5752 -5564 5768 -5547
rect 5752 -5581 5794 -5564
rect 5634 -5628 5794 -5581
rect 3672 -6075 3832 -6028
rect 3672 -6092 3714 -6075
rect 3698 -6109 3714 -6092
rect 3790 -6092 3832 -6075
rect 3890 -6075 4050 -6028
rect 3890 -6092 3932 -6075
rect 3790 -6109 3806 -6092
rect 3698 -6125 3806 -6109
rect 3916 -6109 3932 -6092
rect 4008 -6092 4050 -6075
rect 4108 -6075 4268 -6028
rect 4108 -6092 4150 -6075
rect 4008 -6109 4024 -6092
rect 3916 -6125 4024 -6109
rect 4134 -6109 4150 -6092
rect 4226 -6092 4268 -6075
rect 4326 -6075 4486 -6028
rect 4326 -6092 4368 -6075
rect 4226 -6109 4242 -6092
rect 4134 -6125 4242 -6109
rect 4352 -6109 4368 -6092
rect 4444 -6092 4486 -6075
rect 4544 -6075 4704 -6028
rect 4544 -6092 4586 -6075
rect 4444 -6109 4460 -6092
rect 4352 -6125 4460 -6109
rect 4570 -6109 4586 -6092
rect 4662 -6092 4704 -6075
rect 4762 -6075 4922 -6028
rect 4762 -6092 4804 -6075
rect 4662 -6109 4678 -6092
rect 4570 -6125 4678 -6109
rect 4788 -6109 4804 -6092
rect 4880 -6092 4922 -6075
rect 4980 -6075 5140 -6028
rect 4980 -6092 5022 -6075
rect 4880 -6109 4896 -6092
rect 4788 -6125 4896 -6109
rect 5006 -6109 5022 -6092
rect 5098 -6092 5140 -6075
rect 5198 -6075 5358 -6028
rect 5198 -6092 5240 -6075
rect 5098 -6109 5114 -6092
rect 5006 -6125 5114 -6109
rect 5224 -6109 5240 -6092
rect 5316 -6092 5358 -6075
rect 5416 -6075 5576 -6028
rect 5416 -6092 5458 -6075
rect 5316 -6109 5332 -6092
rect 5224 -6125 5332 -6109
rect 5442 -6109 5458 -6092
rect 5534 -6092 5576 -6075
rect 5634 -6075 5794 -6028
rect 5634 -6092 5676 -6075
rect 5534 -6109 5550 -6092
rect 5442 -6125 5550 -6109
rect 5660 -6109 5676 -6092
rect 5752 -6092 5794 -6075
rect 5752 -6109 5768 -6092
rect 5660 -6125 5768 -6109
rect 3698 -6485 3806 -6469
rect 3698 -6502 3714 -6485
rect 3672 -6519 3714 -6502
rect 3790 -6502 3806 -6485
rect 3916 -6485 4024 -6469
rect 3916 -6502 3932 -6485
rect 3790 -6519 3832 -6502
rect 3672 -6566 3832 -6519
rect 3890 -6519 3932 -6502
rect 4008 -6502 4024 -6485
rect 4134 -6485 4242 -6469
rect 4134 -6502 4150 -6485
rect 4008 -6519 4050 -6502
rect 3890 -6566 4050 -6519
rect 4108 -6519 4150 -6502
rect 4226 -6502 4242 -6485
rect 4352 -6485 4460 -6469
rect 4352 -6502 4368 -6485
rect 4226 -6519 4268 -6502
rect 4108 -6566 4268 -6519
rect 4326 -6519 4368 -6502
rect 4444 -6502 4460 -6485
rect 4570 -6485 4678 -6469
rect 4570 -6502 4586 -6485
rect 4444 -6519 4486 -6502
rect 4326 -6566 4486 -6519
rect 4544 -6519 4586 -6502
rect 4662 -6502 4678 -6485
rect 4788 -6485 4896 -6469
rect 4788 -6502 4804 -6485
rect 4662 -6519 4704 -6502
rect 4544 -6566 4704 -6519
rect 4762 -6519 4804 -6502
rect 4880 -6502 4896 -6485
rect 5006 -6485 5114 -6469
rect 5006 -6502 5022 -6485
rect 4880 -6519 4922 -6502
rect 4762 -6566 4922 -6519
rect 4980 -6519 5022 -6502
rect 5098 -6502 5114 -6485
rect 5224 -6485 5332 -6469
rect 5224 -6502 5240 -6485
rect 5098 -6519 5140 -6502
rect 4980 -6566 5140 -6519
rect 5198 -6519 5240 -6502
rect 5316 -6502 5332 -6485
rect 5442 -6485 5550 -6469
rect 5442 -6502 5458 -6485
rect 5316 -6519 5358 -6502
rect 5198 -6566 5358 -6519
rect 5416 -6519 5458 -6502
rect 5534 -6502 5550 -6485
rect 5660 -6485 5768 -6469
rect 5660 -6502 5676 -6485
rect 5534 -6519 5576 -6502
rect 5416 -6566 5576 -6519
rect 5634 -6519 5676 -6502
rect 5752 -6502 5768 -6485
rect 5752 -6519 5794 -6502
rect 5634 -6566 5794 -6519
rect 3672 -7013 3832 -6966
rect 3672 -7030 3714 -7013
rect 3698 -7047 3714 -7030
rect 3790 -7030 3832 -7013
rect 3890 -7013 4050 -6966
rect 3890 -7030 3932 -7013
rect 3790 -7047 3806 -7030
rect 3698 -7063 3806 -7047
rect 3916 -7047 3932 -7030
rect 4008 -7030 4050 -7013
rect 4108 -7013 4268 -6966
rect 4108 -7030 4150 -7013
rect 4008 -7047 4024 -7030
rect 3916 -7063 4024 -7047
rect 4134 -7047 4150 -7030
rect 4226 -7030 4268 -7013
rect 4326 -7013 4486 -6966
rect 4326 -7030 4368 -7013
rect 4226 -7047 4242 -7030
rect 4134 -7063 4242 -7047
rect 4352 -7047 4368 -7030
rect 4444 -7030 4486 -7013
rect 4544 -7013 4704 -6966
rect 4544 -7030 4586 -7013
rect 4444 -7047 4460 -7030
rect 4352 -7063 4460 -7047
rect 4570 -7047 4586 -7030
rect 4662 -7030 4704 -7013
rect 4762 -7013 4922 -6966
rect 4762 -7030 4804 -7013
rect 4662 -7047 4678 -7030
rect 4570 -7063 4678 -7047
rect 4788 -7047 4804 -7030
rect 4880 -7030 4922 -7013
rect 4980 -7013 5140 -6966
rect 4980 -7030 5022 -7013
rect 4880 -7047 4896 -7030
rect 4788 -7063 4896 -7047
rect 5006 -7047 5022 -7030
rect 5098 -7030 5140 -7013
rect 5198 -7013 5358 -6966
rect 5198 -7030 5240 -7013
rect 5098 -7047 5114 -7030
rect 5006 -7063 5114 -7047
rect 5224 -7047 5240 -7030
rect 5316 -7030 5358 -7013
rect 5416 -7013 5576 -6966
rect 5416 -7030 5458 -7013
rect 5316 -7047 5332 -7030
rect 5224 -7063 5332 -7047
rect 5442 -7047 5458 -7030
rect 5534 -7030 5576 -7013
rect 5634 -7013 5794 -6966
rect 5634 -7030 5676 -7013
rect 5534 -7047 5550 -7030
rect 5442 -7063 5550 -7047
rect 5660 -7047 5676 -7030
rect 5752 -7030 5794 -7013
rect 5752 -7047 5768 -7030
rect 5660 -7063 5768 -7047
rect 3698 -7423 3806 -7407
rect 3698 -7440 3714 -7423
rect 3672 -7457 3714 -7440
rect 3790 -7440 3806 -7423
rect 3916 -7423 4024 -7407
rect 3916 -7440 3932 -7423
rect 3790 -7457 3832 -7440
rect 3672 -7504 3832 -7457
rect 3890 -7457 3932 -7440
rect 4008 -7440 4024 -7423
rect 4134 -7423 4242 -7407
rect 4134 -7440 4150 -7423
rect 4008 -7457 4050 -7440
rect 3890 -7504 4050 -7457
rect 4108 -7457 4150 -7440
rect 4226 -7440 4242 -7423
rect 4352 -7423 4460 -7407
rect 4352 -7440 4368 -7423
rect 4226 -7457 4268 -7440
rect 4108 -7504 4268 -7457
rect 4326 -7457 4368 -7440
rect 4444 -7440 4460 -7423
rect 4570 -7423 4678 -7407
rect 4570 -7440 4586 -7423
rect 4444 -7457 4486 -7440
rect 4326 -7504 4486 -7457
rect 4544 -7457 4586 -7440
rect 4662 -7440 4678 -7423
rect 4788 -7423 4896 -7407
rect 4788 -7440 4804 -7423
rect 4662 -7457 4704 -7440
rect 4544 -7504 4704 -7457
rect 4762 -7457 4804 -7440
rect 4880 -7440 4896 -7423
rect 5006 -7423 5114 -7407
rect 5006 -7440 5022 -7423
rect 4880 -7457 4922 -7440
rect 4762 -7504 4922 -7457
rect 4980 -7457 5022 -7440
rect 5098 -7440 5114 -7423
rect 5224 -7423 5332 -7407
rect 5224 -7440 5240 -7423
rect 5098 -7457 5140 -7440
rect 4980 -7504 5140 -7457
rect 5198 -7457 5240 -7440
rect 5316 -7440 5332 -7423
rect 5442 -7423 5550 -7407
rect 5442 -7440 5458 -7423
rect 5316 -7457 5358 -7440
rect 5198 -7504 5358 -7457
rect 5416 -7457 5458 -7440
rect 5534 -7440 5550 -7423
rect 5660 -7423 5768 -7407
rect 5660 -7440 5676 -7423
rect 5534 -7457 5576 -7440
rect 5416 -7504 5576 -7457
rect 5634 -7457 5676 -7440
rect 5752 -7440 5768 -7423
rect 5752 -7457 5794 -7440
rect 5634 -7504 5794 -7457
rect 3672 -7951 3832 -7904
rect 3672 -7968 3714 -7951
rect 3698 -7985 3714 -7968
rect 3790 -7968 3832 -7951
rect 3890 -7951 4050 -7904
rect 3890 -7968 3932 -7951
rect 3790 -7985 3806 -7968
rect 3698 -8001 3806 -7985
rect 3916 -7985 3932 -7968
rect 4008 -7968 4050 -7951
rect 4108 -7951 4268 -7904
rect 4108 -7968 4150 -7951
rect 4008 -7985 4024 -7968
rect 3916 -8001 4024 -7985
rect 4134 -7985 4150 -7968
rect 4226 -7968 4268 -7951
rect 4326 -7951 4486 -7904
rect 4326 -7968 4368 -7951
rect 4226 -7985 4242 -7968
rect 4134 -8001 4242 -7985
rect 4352 -7985 4368 -7968
rect 4444 -7968 4486 -7951
rect 4544 -7951 4704 -7904
rect 4544 -7968 4586 -7951
rect 4444 -7985 4460 -7968
rect 4352 -8001 4460 -7985
rect 4570 -7985 4586 -7968
rect 4662 -7968 4704 -7951
rect 4762 -7951 4922 -7904
rect 4762 -7968 4804 -7951
rect 4662 -7985 4678 -7968
rect 4570 -8001 4678 -7985
rect 4788 -7985 4804 -7968
rect 4880 -7968 4922 -7951
rect 4980 -7951 5140 -7904
rect 4980 -7968 5022 -7951
rect 4880 -7985 4896 -7968
rect 4788 -8001 4896 -7985
rect 5006 -7985 5022 -7968
rect 5098 -7968 5140 -7951
rect 5198 -7951 5358 -7904
rect 5198 -7968 5240 -7951
rect 5098 -7985 5114 -7968
rect 5006 -8001 5114 -7985
rect 5224 -7985 5240 -7968
rect 5316 -7968 5358 -7951
rect 5416 -7951 5576 -7904
rect 5416 -7968 5458 -7951
rect 5316 -7985 5332 -7968
rect 5224 -8001 5332 -7985
rect 5442 -7985 5458 -7968
rect 5534 -7968 5576 -7951
rect 5634 -7951 5794 -7904
rect 5634 -7968 5676 -7951
rect 5534 -7985 5550 -7968
rect 5442 -8001 5550 -7985
rect 5660 -7985 5676 -7968
rect 5752 -7968 5794 -7951
rect 5752 -7985 5768 -7968
rect 5660 -8001 5768 -7985
rect 2814 -11646 3402 -11630
rect 2814 -11663 2830 -11646
rect 2628 -11680 2830 -11663
rect 3386 -11663 3402 -11646
rect 3832 -11646 4420 -11630
rect 3832 -11663 3848 -11646
rect 3386 -11680 3588 -11663
rect 2628 -11718 3588 -11680
rect 3646 -11680 3848 -11663
rect 4404 -11663 4420 -11646
rect 4850 -11646 5438 -11630
rect 4850 -11663 4866 -11646
rect 4404 -11680 4606 -11663
rect 3646 -11718 4606 -11680
rect 4664 -11680 4866 -11663
rect 5422 -11663 5438 -11646
rect 5868 -11646 6456 -11630
rect 5868 -11663 5884 -11646
rect 5422 -11680 5624 -11663
rect 4664 -11718 5624 -11680
rect 5682 -11680 5884 -11663
rect 6440 -11663 6456 -11646
rect 6886 -11646 7474 -11630
rect 6886 -11663 6902 -11646
rect 6440 -11680 6642 -11663
rect 5682 -11718 6642 -11680
rect 6700 -11680 6902 -11663
rect 7458 -11663 7474 -11646
rect 7904 -11646 8492 -11630
rect 7904 -11663 7920 -11646
rect 7458 -11680 7660 -11663
rect 6700 -11718 7660 -11680
rect 7718 -11680 7920 -11663
rect 8476 -11663 8492 -11646
rect 8922 -11646 9510 -11630
rect 8922 -11663 8938 -11646
rect 8476 -11680 8678 -11663
rect 7718 -11718 8678 -11680
rect 8736 -11680 8938 -11663
rect 9494 -11663 9510 -11646
rect 9940 -11646 10528 -11630
rect 9940 -11663 9956 -11646
rect 9494 -11680 9696 -11663
rect 8736 -11718 9696 -11680
rect 9754 -11680 9956 -11663
rect 10512 -11663 10528 -11646
rect 10958 -11646 11546 -11630
rect 10958 -11663 10974 -11646
rect 10512 -11680 10714 -11663
rect 9754 -11718 10714 -11680
rect 10772 -11680 10974 -11663
rect 11530 -11663 11546 -11646
rect 11976 -11646 12564 -11630
rect 11976 -11663 11992 -11646
rect 11530 -11680 11732 -11663
rect 10772 -11718 11732 -11680
rect 11790 -11680 11992 -11663
rect 12548 -11663 12564 -11646
rect 12994 -11646 13582 -11630
rect 12994 -11663 13010 -11646
rect 12548 -11680 12750 -11663
rect 11790 -11718 12750 -11680
rect 12808 -11680 13010 -11663
rect 13566 -11663 13582 -11646
rect 14012 -11646 14600 -11630
rect 14012 -11663 14028 -11646
rect 13566 -11680 13768 -11663
rect 12808 -11718 13768 -11680
rect 13826 -11680 14028 -11663
rect 14584 -11663 14600 -11646
rect 15030 -11646 15618 -11630
rect 15030 -11663 15046 -11646
rect 14584 -11680 14786 -11663
rect 13826 -11718 14786 -11680
rect 14844 -11680 15046 -11663
rect 15602 -11663 15618 -11646
rect 16048 -11646 16636 -11630
rect 16048 -11663 16064 -11646
rect 15602 -11680 15804 -11663
rect 14844 -11718 15804 -11680
rect 15862 -11680 16064 -11663
rect 16620 -11663 16636 -11646
rect 17066 -11646 17654 -11630
rect 17066 -11663 17082 -11646
rect 16620 -11680 16822 -11663
rect 15862 -11718 16822 -11680
rect 16880 -11680 17082 -11663
rect 17638 -11663 17654 -11646
rect 18084 -11646 18672 -11630
rect 18084 -11663 18100 -11646
rect 17638 -11680 17840 -11663
rect 16880 -11718 17840 -11680
rect 17898 -11680 18100 -11663
rect 18656 -11663 18672 -11646
rect 19102 -11646 19690 -11630
rect 19102 -11663 19118 -11646
rect 18656 -11680 18858 -11663
rect 17898 -11718 18858 -11680
rect 18916 -11680 19118 -11663
rect 19674 -11663 19690 -11646
rect 20120 -11646 20708 -11630
rect 20120 -11663 20136 -11646
rect 19674 -11680 19876 -11663
rect 18916 -11718 19876 -11680
rect 19934 -11680 20136 -11663
rect 20692 -11663 20708 -11646
rect 21138 -11646 21726 -11630
rect 21138 -11663 21154 -11646
rect 20692 -11680 20894 -11663
rect 19934 -11718 20894 -11680
rect 20952 -11680 21154 -11663
rect 21710 -11663 21726 -11646
rect 22156 -11646 22744 -11630
rect 22156 -11663 22172 -11646
rect 21710 -11680 21912 -11663
rect 20952 -11718 21912 -11680
rect 21970 -11680 22172 -11663
rect 22728 -11663 22744 -11646
rect 22728 -11680 22930 -11663
rect 21970 -11718 22930 -11680
rect 2628 -12356 3588 -12318
rect 2628 -12373 2830 -12356
rect 2814 -12390 2830 -12373
rect 3386 -12373 3588 -12356
rect 3646 -12356 4606 -12318
rect 3646 -12373 3848 -12356
rect 3386 -12390 3402 -12373
rect 2814 -12406 3402 -12390
rect 3832 -12390 3848 -12373
rect 4404 -12373 4606 -12356
rect 4664 -12356 5624 -12318
rect 4664 -12373 4866 -12356
rect 4404 -12390 4420 -12373
rect 3832 -12406 4420 -12390
rect 4850 -12390 4866 -12373
rect 5422 -12373 5624 -12356
rect 5682 -12356 6642 -12318
rect 5682 -12373 5884 -12356
rect 5422 -12390 5438 -12373
rect 4850 -12406 5438 -12390
rect 5868 -12390 5884 -12373
rect 6440 -12373 6642 -12356
rect 6700 -12356 7660 -12318
rect 6700 -12373 6902 -12356
rect 6440 -12390 6456 -12373
rect 5868 -12406 6456 -12390
rect 6886 -12390 6902 -12373
rect 7458 -12373 7660 -12356
rect 7718 -12356 8678 -12318
rect 7718 -12373 7920 -12356
rect 7458 -12390 7474 -12373
rect 6886 -12406 7474 -12390
rect 7904 -12390 7920 -12373
rect 8476 -12373 8678 -12356
rect 8736 -12356 9696 -12318
rect 8736 -12373 8938 -12356
rect 8476 -12390 8492 -12373
rect 7904 -12406 8492 -12390
rect 8922 -12390 8938 -12373
rect 9494 -12373 9696 -12356
rect 9754 -12356 10714 -12318
rect 9754 -12373 9956 -12356
rect 9494 -12390 9510 -12373
rect 8922 -12406 9510 -12390
rect 9940 -12390 9956 -12373
rect 10512 -12373 10714 -12356
rect 10772 -12356 11732 -12318
rect 10772 -12373 10974 -12356
rect 10512 -12390 10528 -12373
rect 9940 -12406 10528 -12390
rect 10958 -12390 10974 -12373
rect 11530 -12373 11732 -12356
rect 11790 -12356 12750 -12318
rect 11790 -12373 11992 -12356
rect 11530 -12390 11546 -12373
rect 10958 -12406 11546 -12390
rect 11976 -12390 11992 -12373
rect 12548 -12373 12750 -12356
rect 12808 -12356 13768 -12318
rect 12808 -12373 13010 -12356
rect 12548 -12390 12564 -12373
rect 11976 -12406 12564 -12390
rect 12994 -12390 13010 -12373
rect 13566 -12373 13768 -12356
rect 13826 -12356 14786 -12318
rect 13826 -12373 14028 -12356
rect 13566 -12390 13582 -12373
rect 12994 -12406 13582 -12390
rect 14012 -12390 14028 -12373
rect 14584 -12373 14786 -12356
rect 14844 -12356 15804 -12318
rect 14844 -12373 15046 -12356
rect 14584 -12390 14600 -12373
rect 14012 -12406 14600 -12390
rect 15030 -12390 15046 -12373
rect 15602 -12373 15804 -12356
rect 15862 -12356 16822 -12318
rect 15862 -12373 16064 -12356
rect 15602 -12390 15618 -12373
rect 15030 -12406 15618 -12390
rect 16048 -12390 16064 -12373
rect 16620 -12373 16822 -12356
rect 16880 -12356 17840 -12318
rect 16880 -12373 17082 -12356
rect 16620 -12390 16636 -12373
rect 16048 -12406 16636 -12390
rect 17066 -12390 17082 -12373
rect 17638 -12373 17840 -12356
rect 17898 -12356 18858 -12318
rect 17898 -12373 18100 -12356
rect 17638 -12390 17654 -12373
rect 17066 -12406 17654 -12390
rect 18084 -12390 18100 -12373
rect 18656 -12373 18858 -12356
rect 18916 -12356 19876 -12318
rect 18916 -12373 19118 -12356
rect 18656 -12390 18672 -12373
rect 18084 -12406 18672 -12390
rect 19102 -12390 19118 -12373
rect 19674 -12373 19876 -12356
rect 19934 -12356 20894 -12318
rect 19934 -12373 20136 -12356
rect 19674 -12390 19690 -12373
rect 19102 -12406 19690 -12390
rect 20120 -12390 20136 -12373
rect 20692 -12373 20894 -12356
rect 20952 -12356 21912 -12318
rect 20952 -12373 21154 -12356
rect 20692 -12390 20708 -12373
rect 20120 -12406 20708 -12390
rect 21138 -12390 21154 -12373
rect 21710 -12373 21912 -12356
rect 21970 -12356 22930 -12318
rect 21970 -12373 22172 -12356
rect 21710 -12390 21726 -12373
rect 21138 -12406 21726 -12390
rect 22156 -12390 22172 -12373
rect 22728 -12373 22930 -12356
rect 22728 -12390 22744 -12373
rect 22156 -12406 22744 -12390
rect -8952 -12440 -8364 -12424
rect -8952 -12457 -8936 -12440
rect -9138 -12474 -8936 -12457
rect -8380 -12457 -8364 -12440
rect -7934 -12440 -7346 -12424
rect -7934 -12457 -7918 -12440
rect -8380 -12474 -8178 -12457
rect -9138 -12512 -8178 -12474
rect -8120 -12474 -7918 -12457
rect -7362 -12457 -7346 -12440
rect -6916 -12440 -6328 -12424
rect -6916 -12457 -6900 -12440
rect -7362 -12474 -7160 -12457
rect -8120 -12512 -7160 -12474
rect -7102 -12474 -6900 -12457
rect -6344 -12457 -6328 -12440
rect -5898 -12440 -5310 -12424
rect -5898 -12457 -5882 -12440
rect -6344 -12474 -6142 -12457
rect -7102 -12512 -6142 -12474
rect -6084 -12474 -5882 -12457
rect -5326 -12457 -5310 -12440
rect -4880 -12440 -4292 -12424
rect -4880 -12457 -4864 -12440
rect -5326 -12474 -5124 -12457
rect -6084 -12512 -5124 -12474
rect -5066 -12474 -4864 -12457
rect -4308 -12457 -4292 -12440
rect -3862 -12440 -3274 -12424
rect -3862 -12457 -3846 -12440
rect -4308 -12474 -4106 -12457
rect -5066 -12512 -4106 -12474
rect -4048 -12474 -3846 -12457
rect -3290 -12457 -3274 -12440
rect -2844 -12440 -2256 -12424
rect -2844 -12457 -2828 -12440
rect -3290 -12474 -3088 -12457
rect -4048 -12512 -3088 -12474
rect -3030 -12474 -2828 -12457
rect -2272 -12457 -2256 -12440
rect -1826 -12440 -1238 -12424
rect -1826 -12457 -1810 -12440
rect -2272 -12474 -2070 -12457
rect -3030 -12512 -2070 -12474
rect -2012 -12474 -1810 -12457
rect -1254 -12457 -1238 -12440
rect -808 -12440 -220 -12424
rect -808 -12457 -792 -12440
rect -1254 -12474 -1052 -12457
rect -2012 -12512 -1052 -12474
rect -994 -12474 -792 -12457
rect -236 -12457 -220 -12440
rect -236 -12474 -34 -12457
rect -994 -12512 -34 -12474
rect 2814 -12880 3402 -12864
rect 2814 -12897 2830 -12880
rect 2628 -12914 2830 -12897
rect 3386 -12897 3402 -12880
rect 3832 -12880 4420 -12864
rect 3832 -12897 3848 -12880
rect 3386 -12914 3588 -12897
rect 2628 -12952 3588 -12914
rect 3646 -12914 3848 -12897
rect 4404 -12897 4420 -12880
rect 4850 -12880 5438 -12864
rect 4850 -12897 4866 -12880
rect 4404 -12914 4606 -12897
rect 3646 -12952 4606 -12914
rect 4664 -12914 4866 -12897
rect 5422 -12897 5438 -12880
rect 5868 -12880 6456 -12864
rect 5868 -12897 5884 -12880
rect 5422 -12914 5624 -12897
rect 4664 -12952 5624 -12914
rect 5682 -12914 5884 -12897
rect 6440 -12897 6456 -12880
rect 6886 -12880 7474 -12864
rect 6886 -12897 6902 -12880
rect 6440 -12914 6642 -12897
rect 5682 -12952 6642 -12914
rect 6700 -12914 6902 -12897
rect 7458 -12897 7474 -12880
rect 7904 -12880 8492 -12864
rect 7904 -12897 7920 -12880
rect 7458 -12914 7660 -12897
rect 6700 -12952 7660 -12914
rect 7718 -12914 7920 -12897
rect 8476 -12897 8492 -12880
rect 8922 -12880 9510 -12864
rect 8922 -12897 8938 -12880
rect 8476 -12914 8678 -12897
rect 7718 -12952 8678 -12914
rect 8736 -12914 8938 -12897
rect 9494 -12897 9510 -12880
rect 9940 -12880 10528 -12864
rect 9940 -12897 9956 -12880
rect 9494 -12914 9696 -12897
rect 8736 -12952 9696 -12914
rect 9754 -12914 9956 -12897
rect 10512 -12897 10528 -12880
rect 10958 -12880 11546 -12864
rect 10958 -12897 10974 -12880
rect 10512 -12914 10714 -12897
rect 9754 -12952 10714 -12914
rect 10772 -12914 10974 -12897
rect 11530 -12897 11546 -12880
rect 11976 -12880 12564 -12864
rect 11976 -12897 11992 -12880
rect 11530 -12914 11732 -12897
rect 10772 -12952 11732 -12914
rect 11790 -12914 11992 -12897
rect 12548 -12897 12564 -12880
rect 12994 -12880 13582 -12864
rect 12994 -12897 13010 -12880
rect 12548 -12914 12750 -12897
rect 11790 -12952 12750 -12914
rect 12808 -12914 13010 -12897
rect 13566 -12897 13582 -12880
rect 14012 -12880 14600 -12864
rect 14012 -12897 14028 -12880
rect 13566 -12914 13768 -12897
rect 12808 -12952 13768 -12914
rect 13826 -12914 14028 -12897
rect 14584 -12897 14600 -12880
rect 15030 -12880 15618 -12864
rect 15030 -12897 15046 -12880
rect 14584 -12914 14786 -12897
rect 13826 -12952 14786 -12914
rect 14844 -12914 15046 -12897
rect 15602 -12897 15618 -12880
rect 16048 -12880 16636 -12864
rect 16048 -12897 16064 -12880
rect 15602 -12914 15804 -12897
rect 14844 -12952 15804 -12914
rect 15862 -12914 16064 -12897
rect 16620 -12897 16636 -12880
rect 17066 -12880 17654 -12864
rect 17066 -12897 17082 -12880
rect 16620 -12914 16822 -12897
rect 15862 -12952 16822 -12914
rect 16880 -12914 17082 -12897
rect 17638 -12897 17654 -12880
rect 18084 -12880 18672 -12864
rect 18084 -12897 18100 -12880
rect 17638 -12914 17840 -12897
rect 16880 -12952 17840 -12914
rect 17898 -12914 18100 -12897
rect 18656 -12897 18672 -12880
rect 19102 -12880 19690 -12864
rect 19102 -12897 19118 -12880
rect 18656 -12914 18858 -12897
rect 17898 -12952 18858 -12914
rect 18916 -12914 19118 -12897
rect 19674 -12897 19690 -12880
rect 20120 -12880 20708 -12864
rect 20120 -12897 20136 -12880
rect 19674 -12914 19876 -12897
rect 18916 -12952 19876 -12914
rect 19934 -12914 20136 -12897
rect 20692 -12897 20708 -12880
rect 21138 -12880 21726 -12864
rect 21138 -12897 21154 -12880
rect 20692 -12914 20894 -12897
rect 19934 -12952 20894 -12914
rect 20952 -12914 21154 -12897
rect 21710 -12897 21726 -12880
rect 22156 -12880 22744 -12864
rect 22156 -12897 22172 -12880
rect 21710 -12914 21912 -12897
rect 20952 -12952 21912 -12914
rect 21970 -12914 22172 -12897
rect 22728 -12897 22744 -12880
rect 22728 -12914 22930 -12897
rect 21970 -12952 22930 -12914
rect -9138 -13150 -8178 -13112
rect -9138 -13167 -8936 -13150
rect -8952 -13184 -8936 -13167
rect -8380 -13167 -8178 -13150
rect -8120 -13150 -7160 -13112
rect -8120 -13167 -7918 -13150
rect -8380 -13184 -8364 -13167
rect -8952 -13200 -8364 -13184
rect -7934 -13184 -7918 -13167
rect -7362 -13167 -7160 -13150
rect -7102 -13150 -6142 -13112
rect -7102 -13167 -6900 -13150
rect -7362 -13184 -7346 -13167
rect -7934 -13200 -7346 -13184
rect -6916 -13184 -6900 -13167
rect -6344 -13167 -6142 -13150
rect -6084 -13150 -5124 -13112
rect -6084 -13167 -5882 -13150
rect -6344 -13184 -6328 -13167
rect -6916 -13200 -6328 -13184
rect -5898 -13184 -5882 -13167
rect -5326 -13167 -5124 -13150
rect -5066 -13150 -4106 -13112
rect -5066 -13167 -4864 -13150
rect -5326 -13184 -5310 -13167
rect -5898 -13200 -5310 -13184
rect -4880 -13184 -4864 -13167
rect -4308 -13167 -4106 -13150
rect -4048 -13150 -3088 -13112
rect -4048 -13167 -3846 -13150
rect -4308 -13184 -4292 -13167
rect -4880 -13200 -4292 -13184
rect -3862 -13184 -3846 -13167
rect -3290 -13167 -3088 -13150
rect -3030 -13150 -2070 -13112
rect -3030 -13167 -2828 -13150
rect -3290 -13184 -3274 -13167
rect -3862 -13200 -3274 -13184
rect -2844 -13184 -2828 -13167
rect -2272 -13167 -2070 -13150
rect -2012 -13150 -1052 -13112
rect -2012 -13167 -1810 -13150
rect -2272 -13184 -2256 -13167
rect -2844 -13200 -2256 -13184
rect -1826 -13184 -1810 -13167
rect -1254 -13167 -1052 -13150
rect -994 -13150 -34 -13112
rect -994 -13167 -792 -13150
rect -1254 -13184 -1238 -13167
rect -1826 -13200 -1238 -13184
rect -808 -13184 -792 -13167
rect -236 -13167 -34 -13150
rect -236 -13184 -220 -13167
rect -808 -13200 -220 -13184
rect -8952 -13258 -8364 -13242
rect -8952 -13275 -8936 -13258
rect -9138 -13292 -8936 -13275
rect -8380 -13275 -8364 -13258
rect -7934 -13258 -7346 -13242
rect -7934 -13275 -7918 -13258
rect -8380 -13292 -8178 -13275
rect -9138 -13330 -8178 -13292
rect -8120 -13292 -7918 -13275
rect -7362 -13275 -7346 -13258
rect -6916 -13258 -6328 -13242
rect -6916 -13275 -6900 -13258
rect -7362 -13292 -7160 -13275
rect -8120 -13330 -7160 -13292
rect -7102 -13292 -6900 -13275
rect -6344 -13275 -6328 -13258
rect -5898 -13258 -5310 -13242
rect -5898 -13275 -5882 -13258
rect -6344 -13292 -6142 -13275
rect -7102 -13330 -6142 -13292
rect -6084 -13292 -5882 -13275
rect -5326 -13275 -5310 -13258
rect -4880 -13258 -4292 -13242
rect -4880 -13275 -4864 -13258
rect -5326 -13292 -5124 -13275
rect -6084 -13330 -5124 -13292
rect -5066 -13292 -4864 -13275
rect -4308 -13275 -4292 -13258
rect -3862 -13258 -3274 -13242
rect -3862 -13275 -3846 -13258
rect -4308 -13292 -4106 -13275
rect -5066 -13330 -4106 -13292
rect -4048 -13292 -3846 -13275
rect -3290 -13275 -3274 -13258
rect -2844 -13258 -2256 -13242
rect -2844 -13275 -2828 -13258
rect -3290 -13292 -3088 -13275
rect -4048 -13330 -3088 -13292
rect -3030 -13292 -2828 -13275
rect -2272 -13275 -2256 -13258
rect -1826 -13258 -1238 -13242
rect -1826 -13275 -1810 -13258
rect -2272 -13292 -2070 -13275
rect -3030 -13330 -2070 -13292
rect -2012 -13292 -1810 -13275
rect -1254 -13275 -1238 -13258
rect -808 -13258 -220 -13242
rect -808 -13275 -792 -13258
rect -1254 -13292 -1052 -13275
rect -2012 -13330 -1052 -13292
rect -994 -13292 -792 -13275
rect -236 -13275 -220 -13258
rect -236 -13292 -34 -13275
rect -994 -13330 -34 -13292
rect 2628 -13590 3588 -13552
rect 2628 -13607 2830 -13590
rect 2814 -13624 2830 -13607
rect 3386 -13607 3588 -13590
rect 3646 -13590 4606 -13552
rect 3646 -13607 3848 -13590
rect 3386 -13624 3402 -13607
rect 2814 -13640 3402 -13624
rect 3832 -13624 3848 -13607
rect 4404 -13607 4606 -13590
rect 4664 -13590 5624 -13552
rect 4664 -13607 4866 -13590
rect 4404 -13624 4420 -13607
rect 3832 -13640 4420 -13624
rect 4850 -13624 4866 -13607
rect 5422 -13607 5624 -13590
rect 5682 -13590 6642 -13552
rect 5682 -13607 5884 -13590
rect 5422 -13624 5438 -13607
rect 4850 -13640 5438 -13624
rect 5868 -13624 5884 -13607
rect 6440 -13607 6642 -13590
rect 6700 -13590 7660 -13552
rect 6700 -13607 6902 -13590
rect 6440 -13624 6456 -13607
rect 5868 -13640 6456 -13624
rect 6886 -13624 6902 -13607
rect 7458 -13607 7660 -13590
rect 7718 -13590 8678 -13552
rect 7718 -13607 7920 -13590
rect 7458 -13624 7474 -13607
rect 6886 -13640 7474 -13624
rect 7904 -13624 7920 -13607
rect 8476 -13607 8678 -13590
rect 8736 -13590 9696 -13552
rect 8736 -13607 8938 -13590
rect 8476 -13624 8492 -13607
rect 7904 -13640 8492 -13624
rect 8922 -13624 8938 -13607
rect 9494 -13607 9696 -13590
rect 9754 -13590 10714 -13552
rect 9754 -13607 9956 -13590
rect 9494 -13624 9510 -13607
rect 8922 -13640 9510 -13624
rect 9940 -13624 9956 -13607
rect 10512 -13607 10714 -13590
rect 10772 -13590 11732 -13552
rect 10772 -13607 10974 -13590
rect 10512 -13624 10528 -13607
rect 9940 -13640 10528 -13624
rect 10958 -13624 10974 -13607
rect 11530 -13607 11732 -13590
rect 11790 -13590 12750 -13552
rect 11790 -13607 11992 -13590
rect 11530 -13624 11546 -13607
rect 10958 -13640 11546 -13624
rect 11976 -13624 11992 -13607
rect 12548 -13607 12750 -13590
rect 12808 -13590 13768 -13552
rect 12808 -13607 13010 -13590
rect 12548 -13624 12564 -13607
rect 11976 -13640 12564 -13624
rect 12994 -13624 13010 -13607
rect 13566 -13607 13768 -13590
rect 13826 -13590 14786 -13552
rect 13826 -13607 14028 -13590
rect 13566 -13624 13582 -13607
rect 12994 -13640 13582 -13624
rect 14012 -13624 14028 -13607
rect 14584 -13607 14786 -13590
rect 14844 -13590 15804 -13552
rect 14844 -13607 15046 -13590
rect 14584 -13624 14600 -13607
rect 14012 -13640 14600 -13624
rect 15030 -13624 15046 -13607
rect 15602 -13607 15804 -13590
rect 15862 -13590 16822 -13552
rect 15862 -13607 16064 -13590
rect 15602 -13624 15618 -13607
rect 15030 -13640 15618 -13624
rect 16048 -13624 16064 -13607
rect 16620 -13607 16822 -13590
rect 16880 -13590 17840 -13552
rect 16880 -13607 17082 -13590
rect 16620 -13624 16636 -13607
rect 16048 -13640 16636 -13624
rect 17066 -13624 17082 -13607
rect 17638 -13607 17840 -13590
rect 17898 -13590 18858 -13552
rect 17898 -13607 18100 -13590
rect 17638 -13624 17654 -13607
rect 17066 -13640 17654 -13624
rect 18084 -13624 18100 -13607
rect 18656 -13607 18858 -13590
rect 18916 -13590 19876 -13552
rect 18916 -13607 19118 -13590
rect 18656 -13624 18672 -13607
rect 18084 -13640 18672 -13624
rect 19102 -13624 19118 -13607
rect 19674 -13607 19876 -13590
rect 19934 -13590 20894 -13552
rect 19934 -13607 20136 -13590
rect 19674 -13624 19690 -13607
rect 19102 -13640 19690 -13624
rect 20120 -13624 20136 -13607
rect 20692 -13607 20894 -13590
rect 20952 -13590 21912 -13552
rect 20952 -13607 21154 -13590
rect 20692 -13624 20708 -13607
rect 20120 -13640 20708 -13624
rect 21138 -13624 21154 -13607
rect 21710 -13607 21912 -13590
rect 21970 -13590 22930 -13552
rect 21970 -13607 22172 -13590
rect 21710 -13624 21726 -13607
rect 21138 -13640 21726 -13624
rect 22156 -13624 22172 -13607
rect 22728 -13607 22930 -13590
rect 22728 -13624 22744 -13607
rect 22156 -13640 22744 -13624
rect -9138 -13968 -8178 -13930
rect -9138 -13985 -8936 -13968
rect -8952 -14002 -8936 -13985
rect -8380 -13985 -8178 -13968
rect -8120 -13968 -7160 -13930
rect -8120 -13985 -7918 -13968
rect -8380 -14002 -8364 -13985
rect -8952 -14018 -8364 -14002
rect -7934 -14002 -7918 -13985
rect -7362 -13985 -7160 -13968
rect -7102 -13968 -6142 -13930
rect -7102 -13985 -6900 -13968
rect -7362 -14002 -7346 -13985
rect -7934 -14018 -7346 -14002
rect -6916 -14002 -6900 -13985
rect -6344 -13985 -6142 -13968
rect -6084 -13968 -5124 -13930
rect -6084 -13985 -5882 -13968
rect -6344 -14002 -6328 -13985
rect -6916 -14018 -6328 -14002
rect -5898 -14002 -5882 -13985
rect -5326 -13985 -5124 -13968
rect -5066 -13968 -4106 -13930
rect -5066 -13985 -4864 -13968
rect -5326 -14002 -5310 -13985
rect -5898 -14018 -5310 -14002
rect -4880 -14002 -4864 -13985
rect -4308 -13985 -4106 -13968
rect -4048 -13968 -3088 -13930
rect -4048 -13985 -3846 -13968
rect -4308 -14002 -4292 -13985
rect -4880 -14018 -4292 -14002
rect -3862 -14002 -3846 -13985
rect -3290 -13985 -3088 -13968
rect -3030 -13968 -2070 -13930
rect -3030 -13985 -2828 -13968
rect -3290 -14002 -3274 -13985
rect -3862 -14018 -3274 -14002
rect -2844 -14002 -2828 -13985
rect -2272 -13985 -2070 -13968
rect -2012 -13968 -1052 -13930
rect -2012 -13985 -1810 -13968
rect -2272 -14002 -2256 -13985
rect -2844 -14018 -2256 -14002
rect -1826 -14002 -1810 -13985
rect -1254 -13985 -1052 -13968
rect -994 -13968 -34 -13930
rect -994 -13985 -792 -13968
rect -1254 -14002 -1238 -13985
rect -1826 -14018 -1238 -14002
rect -808 -14002 -792 -13985
rect -236 -13985 -34 -13968
rect -236 -14002 -220 -13985
rect -808 -14018 -220 -14002
rect -8952 -14076 -8364 -14060
rect -8952 -14093 -8936 -14076
rect -9138 -14110 -8936 -14093
rect -8380 -14093 -8364 -14076
rect -7934 -14076 -7346 -14060
rect -7934 -14093 -7918 -14076
rect -8380 -14110 -8178 -14093
rect -9138 -14148 -8178 -14110
rect -8120 -14110 -7918 -14093
rect -7362 -14093 -7346 -14076
rect -6916 -14076 -6328 -14060
rect -6916 -14093 -6900 -14076
rect -7362 -14110 -7160 -14093
rect -8120 -14148 -7160 -14110
rect -7102 -14110 -6900 -14093
rect -6344 -14093 -6328 -14076
rect -5898 -14076 -5310 -14060
rect -5898 -14093 -5882 -14076
rect -6344 -14110 -6142 -14093
rect -7102 -14148 -6142 -14110
rect -6084 -14110 -5882 -14093
rect -5326 -14093 -5310 -14076
rect -4880 -14076 -4292 -14060
rect -4880 -14093 -4864 -14076
rect -5326 -14110 -5124 -14093
rect -6084 -14148 -5124 -14110
rect -5066 -14110 -4864 -14093
rect -4308 -14093 -4292 -14076
rect -3862 -14076 -3274 -14060
rect -3862 -14093 -3846 -14076
rect -4308 -14110 -4106 -14093
rect -5066 -14148 -4106 -14110
rect -4048 -14110 -3846 -14093
rect -3290 -14093 -3274 -14076
rect -2844 -14076 -2256 -14060
rect -2844 -14093 -2828 -14076
rect -3290 -14110 -3088 -14093
rect -4048 -14148 -3088 -14110
rect -3030 -14110 -2828 -14093
rect -2272 -14093 -2256 -14076
rect -1826 -14076 -1238 -14060
rect -1826 -14093 -1810 -14076
rect -2272 -14110 -2070 -14093
rect -3030 -14148 -2070 -14110
rect -2012 -14110 -1810 -14093
rect -1254 -14093 -1238 -14076
rect -808 -14076 -220 -14060
rect -808 -14093 -792 -14076
rect -1254 -14110 -1052 -14093
rect -2012 -14148 -1052 -14110
rect -994 -14110 -792 -14093
rect -236 -14093 -220 -14076
rect -236 -14110 -34 -14093
rect -994 -14148 -34 -14110
rect 2814 -14112 3402 -14096
rect 2814 -14129 2830 -14112
rect 2628 -14146 2830 -14129
rect 3386 -14129 3402 -14112
rect 3832 -14112 4420 -14096
rect 3832 -14129 3848 -14112
rect 3386 -14146 3588 -14129
rect 2628 -14184 3588 -14146
rect 3646 -14146 3848 -14129
rect 4404 -14129 4420 -14112
rect 4850 -14112 5438 -14096
rect 4850 -14129 4866 -14112
rect 4404 -14146 4606 -14129
rect 3646 -14184 4606 -14146
rect 4664 -14146 4866 -14129
rect 5422 -14129 5438 -14112
rect 5868 -14112 6456 -14096
rect 5868 -14129 5884 -14112
rect 5422 -14146 5624 -14129
rect 4664 -14184 5624 -14146
rect 5682 -14146 5884 -14129
rect 6440 -14129 6456 -14112
rect 6886 -14112 7474 -14096
rect 6886 -14129 6902 -14112
rect 6440 -14146 6642 -14129
rect 5682 -14184 6642 -14146
rect 6700 -14146 6902 -14129
rect 7458 -14129 7474 -14112
rect 7904 -14112 8492 -14096
rect 7904 -14129 7920 -14112
rect 7458 -14146 7660 -14129
rect 6700 -14184 7660 -14146
rect 7718 -14146 7920 -14129
rect 8476 -14129 8492 -14112
rect 8922 -14112 9510 -14096
rect 8922 -14129 8938 -14112
rect 8476 -14146 8678 -14129
rect 7718 -14184 8678 -14146
rect 8736 -14146 8938 -14129
rect 9494 -14129 9510 -14112
rect 9940 -14112 10528 -14096
rect 9940 -14129 9956 -14112
rect 9494 -14146 9696 -14129
rect 8736 -14184 9696 -14146
rect 9754 -14146 9956 -14129
rect 10512 -14129 10528 -14112
rect 10958 -14112 11546 -14096
rect 10958 -14129 10974 -14112
rect 10512 -14146 10714 -14129
rect 9754 -14184 10714 -14146
rect 10772 -14146 10974 -14129
rect 11530 -14129 11546 -14112
rect 11976 -14112 12564 -14096
rect 11976 -14129 11992 -14112
rect 11530 -14146 11732 -14129
rect 10772 -14184 11732 -14146
rect 11790 -14146 11992 -14129
rect 12548 -14129 12564 -14112
rect 12994 -14112 13582 -14096
rect 12994 -14129 13010 -14112
rect 12548 -14146 12750 -14129
rect 11790 -14184 12750 -14146
rect 12808 -14146 13010 -14129
rect 13566 -14129 13582 -14112
rect 14012 -14112 14600 -14096
rect 14012 -14129 14028 -14112
rect 13566 -14146 13768 -14129
rect 12808 -14184 13768 -14146
rect 13826 -14146 14028 -14129
rect 14584 -14129 14600 -14112
rect 15030 -14112 15618 -14096
rect 15030 -14129 15046 -14112
rect 14584 -14146 14786 -14129
rect 13826 -14184 14786 -14146
rect 14844 -14146 15046 -14129
rect 15602 -14129 15618 -14112
rect 16048 -14112 16636 -14096
rect 16048 -14129 16064 -14112
rect 15602 -14146 15804 -14129
rect 14844 -14184 15804 -14146
rect 15862 -14146 16064 -14129
rect 16620 -14129 16636 -14112
rect 17066 -14112 17654 -14096
rect 17066 -14129 17082 -14112
rect 16620 -14146 16822 -14129
rect 15862 -14184 16822 -14146
rect 16880 -14146 17082 -14129
rect 17638 -14129 17654 -14112
rect 18084 -14112 18672 -14096
rect 18084 -14129 18100 -14112
rect 17638 -14146 17840 -14129
rect 16880 -14184 17840 -14146
rect 17898 -14146 18100 -14129
rect 18656 -14129 18672 -14112
rect 19102 -14112 19690 -14096
rect 19102 -14129 19118 -14112
rect 18656 -14146 18858 -14129
rect 17898 -14184 18858 -14146
rect 18916 -14146 19118 -14129
rect 19674 -14129 19690 -14112
rect 20120 -14112 20708 -14096
rect 20120 -14129 20136 -14112
rect 19674 -14146 19876 -14129
rect 18916 -14184 19876 -14146
rect 19934 -14146 20136 -14129
rect 20692 -14129 20708 -14112
rect 21138 -14112 21726 -14096
rect 21138 -14129 21154 -14112
rect 20692 -14146 20894 -14129
rect 19934 -14184 20894 -14146
rect 20952 -14146 21154 -14129
rect 21710 -14129 21726 -14112
rect 22156 -14112 22744 -14096
rect 22156 -14129 22172 -14112
rect 21710 -14146 21912 -14129
rect 20952 -14184 21912 -14146
rect 21970 -14146 22172 -14129
rect 22728 -14129 22744 -14112
rect 22728 -14146 22930 -14129
rect 21970 -14184 22930 -14146
rect -9138 -14786 -8178 -14748
rect -9138 -14803 -8936 -14786
rect -8952 -14820 -8936 -14803
rect -8380 -14803 -8178 -14786
rect -8120 -14786 -7160 -14748
rect -8120 -14803 -7918 -14786
rect -8380 -14820 -8364 -14803
rect -8952 -14836 -8364 -14820
rect -7934 -14820 -7918 -14803
rect -7362 -14803 -7160 -14786
rect -7102 -14786 -6142 -14748
rect -7102 -14803 -6900 -14786
rect -7362 -14820 -7346 -14803
rect -7934 -14836 -7346 -14820
rect -6916 -14820 -6900 -14803
rect -6344 -14803 -6142 -14786
rect -6084 -14786 -5124 -14748
rect -6084 -14803 -5882 -14786
rect -6344 -14820 -6328 -14803
rect -6916 -14836 -6328 -14820
rect -5898 -14820 -5882 -14803
rect -5326 -14803 -5124 -14786
rect -5066 -14786 -4106 -14748
rect -5066 -14803 -4864 -14786
rect -5326 -14820 -5310 -14803
rect -5898 -14836 -5310 -14820
rect -4880 -14820 -4864 -14803
rect -4308 -14803 -4106 -14786
rect -4048 -14786 -3088 -14748
rect -4048 -14803 -3846 -14786
rect -4308 -14820 -4292 -14803
rect -4880 -14836 -4292 -14820
rect -3862 -14820 -3846 -14803
rect -3290 -14803 -3088 -14786
rect -3030 -14786 -2070 -14748
rect -3030 -14803 -2828 -14786
rect -3290 -14820 -3274 -14803
rect -3862 -14836 -3274 -14820
rect -2844 -14820 -2828 -14803
rect -2272 -14803 -2070 -14786
rect -2012 -14786 -1052 -14748
rect -2012 -14803 -1810 -14786
rect -2272 -14820 -2256 -14803
rect -2844 -14836 -2256 -14820
rect -1826 -14820 -1810 -14803
rect -1254 -14803 -1052 -14786
rect -994 -14786 -34 -14748
rect -994 -14803 -792 -14786
rect -1254 -14820 -1238 -14803
rect -1826 -14836 -1238 -14820
rect -808 -14820 -792 -14803
rect -236 -14803 -34 -14786
rect -236 -14820 -220 -14803
rect -808 -14836 -220 -14820
rect 2628 -14822 3588 -14784
rect 2628 -14839 2830 -14822
rect 2814 -14856 2830 -14839
rect 3386 -14839 3588 -14822
rect 3646 -14822 4606 -14784
rect 3646 -14839 3848 -14822
rect 3386 -14856 3402 -14839
rect 2814 -14872 3402 -14856
rect 3832 -14856 3848 -14839
rect 4404 -14839 4606 -14822
rect 4664 -14822 5624 -14784
rect 4664 -14839 4866 -14822
rect 4404 -14856 4420 -14839
rect 3832 -14872 4420 -14856
rect 4850 -14856 4866 -14839
rect 5422 -14839 5624 -14822
rect 5682 -14822 6642 -14784
rect 5682 -14839 5884 -14822
rect 5422 -14856 5438 -14839
rect 4850 -14872 5438 -14856
rect 5868 -14856 5884 -14839
rect 6440 -14839 6642 -14822
rect 6700 -14822 7660 -14784
rect 6700 -14839 6902 -14822
rect 6440 -14856 6456 -14839
rect 5868 -14872 6456 -14856
rect 6886 -14856 6902 -14839
rect 7458 -14839 7660 -14822
rect 7718 -14822 8678 -14784
rect 7718 -14839 7920 -14822
rect 7458 -14856 7474 -14839
rect 6886 -14872 7474 -14856
rect 7904 -14856 7920 -14839
rect 8476 -14839 8678 -14822
rect 8736 -14822 9696 -14784
rect 8736 -14839 8938 -14822
rect 8476 -14856 8492 -14839
rect 7904 -14872 8492 -14856
rect 8922 -14856 8938 -14839
rect 9494 -14839 9696 -14822
rect 9754 -14822 10714 -14784
rect 9754 -14839 9956 -14822
rect 9494 -14856 9510 -14839
rect 8922 -14872 9510 -14856
rect 9940 -14856 9956 -14839
rect 10512 -14839 10714 -14822
rect 10772 -14822 11732 -14784
rect 10772 -14839 10974 -14822
rect 10512 -14856 10528 -14839
rect 9940 -14872 10528 -14856
rect 10958 -14856 10974 -14839
rect 11530 -14839 11732 -14822
rect 11790 -14822 12750 -14784
rect 11790 -14839 11992 -14822
rect 11530 -14856 11546 -14839
rect 10958 -14872 11546 -14856
rect 11976 -14856 11992 -14839
rect 12548 -14839 12750 -14822
rect 12808 -14822 13768 -14784
rect 12808 -14839 13010 -14822
rect 12548 -14856 12564 -14839
rect 11976 -14872 12564 -14856
rect 12994 -14856 13010 -14839
rect 13566 -14839 13768 -14822
rect 13826 -14822 14786 -14784
rect 13826 -14839 14028 -14822
rect 13566 -14856 13582 -14839
rect 12994 -14872 13582 -14856
rect 14012 -14856 14028 -14839
rect 14584 -14839 14786 -14822
rect 14844 -14822 15804 -14784
rect 14844 -14839 15046 -14822
rect 14584 -14856 14600 -14839
rect 14012 -14872 14600 -14856
rect 15030 -14856 15046 -14839
rect 15602 -14839 15804 -14822
rect 15862 -14822 16822 -14784
rect 15862 -14839 16064 -14822
rect 15602 -14856 15618 -14839
rect 15030 -14872 15618 -14856
rect 16048 -14856 16064 -14839
rect 16620 -14839 16822 -14822
rect 16880 -14822 17840 -14784
rect 16880 -14839 17082 -14822
rect 16620 -14856 16636 -14839
rect 16048 -14872 16636 -14856
rect 17066 -14856 17082 -14839
rect 17638 -14839 17840 -14822
rect 17898 -14822 18858 -14784
rect 17898 -14839 18100 -14822
rect 17638 -14856 17654 -14839
rect 17066 -14872 17654 -14856
rect 18084 -14856 18100 -14839
rect 18656 -14839 18858 -14822
rect 18916 -14822 19876 -14784
rect 18916 -14839 19118 -14822
rect 18656 -14856 18672 -14839
rect 18084 -14872 18672 -14856
rect 19102 -14856 19118 -14839
rect 19674 -14839 19876 -14822
rect 19934 -14822 20894 -14784
rect 19934 -14839 20136 -14822
rect 19674 -14856 19690 -14839
rect 19102 -14872 19690 -14856
rect 20120 -14856 20136 -14839
rect 20692 -14839 20894 -14822
rect 20952 -14822 21912 -14784
rect 20952 -14839 21154 -14822
rect 20692 -14856 20708 -14839
rect 20120 -14872 20708 -14856
rect 21138 -14856 21154 -14839
rect 21710 -14839 21912 -14822
rect 21970 -14822 22930 -14784
rect 21970 -14839 22172 -14822
rect 21710 -14856 21726 -14839
rect 21138 -14872 21726 -14856
rect 22156 -14856 22172 -14839
rect 22728 -14839 22930 -14822
rect 22728 -14856 22744 -14839
rect 22156 -14872 22744 -14856
rect -8952 -14894 -8364 -14878
rect -8952 -14911 -8936 -14894
rect -9138 -14928 -8936 -14911
rect -8380 -14911 -8364 -14894
rect -7934 -14894 -7346 -14878
rect -7934 -14911 -7918 -14894
rect -8380 -14928 -8178 -14911
rect -9138 -14966 -8178 -14928
rect -8120 -14928 -7918 -14911
rect -7362 -14911 -7346 -14894
rect -6916 -14894 -6328 -14878
rect -6916 -14911 -6900 -14894
rect -7362 -14928 -7160 -14911
rect -8120 -14966 -7160 -14928
rect -7102 -14928 -6900 -14911
rect -6344 -14911 -6328 -14894
rect -5898 -14894 -5310 -14878
rect -5898 -14911 -5882 -14894
rect -6344 -14928 -6142 -14911
rect -7102 -14966 -6142 -14928
rect -6084 -14928 -5882 -14911
rect -5326 -14911 -5310 -14894
rect -4880 -14894 -4292 -14878
rect -4880 -14911 -4864 -14894
rect -5326 -14928 -5124 -14911
rect -6084 -14966 -5124 -14928
rect -5066 -14928 -4864 -14911
rect -4308 -14911 -4292 -14894
rect -3862 -14894 -3274 -14878
rect -3862 -14911 -3846 -14894
rect -4308 -14928 -4106 -14911
rect -5066 -14966 -4106 -14928
rect -4048 -14928 -3846 -14911
rect -3290 -14911 -3274 -14894
rect -2844 -14894 -2256 -14878
rect -2844 -14911 -2828 -14894
rect -3290 -14928 -3088 -14911
rect -4048 -14966 -3088 -14928
rect -3030 -14928 -2828 -14911
rect -2272 -14911 -2256 -14894
rect -1826 -14894 -1238 -14878
rect -1826 -14911 -1810 -14894
rect -2272 -14928 -2070 -14911
rect -3030 -14966 -2070 -14928
rect -2012 -14928 -1810 -14911
rect -1254 -14911 -1238 -14894
rect -808 -14894 -220 -14878
rect -808 -14911 -792 -14894
rect -1254 -14928 -1052 -14911
rect -2012 -14966 -1052 -14928
rect -994 -14928 -792 -14911
rect -236 -14911 -220 -14894
rect -236 -14928 -34 -14911
rect -994 -14966 -34 -14928
rect 2812 -15346 3400 -15330
rect 2812 -15363 2828 -15346
rect 2626 -15380 2828 -15363
rect 3384 -15363 3400 -15346
rect 3830 -15346 4418 -15330
rect 3830 -15363 3846 -15346
rect 3384 -15380 3586 -15363
rect 2626 -15418 3586 -15380
rect 3644 -15380 3846 -15363
rect 4402 -15363 4418 -15346
rect 4848 -15346 5436 -15330
rect 4848 -15363 4864 -15346
rect 4402 -15380 4604 -15363
rect 3644 -15418 4604 -15380
rect 4662 -15380 4864 -15363
rect 5420 -15363 5436 -15346
rect 5866 -15346 6454 -15330
rect 5866 -15363 5882 -15346
rect 5420 -15380 5622 -15363
rect 4662 -15418 5622 -15380
rect 5680 -15380 5882 -15363
rect 6438 -15363 6454 -15346
rect 6884 -15346 7472 -15330
rect 6884 -15363 6900 -15346
rect 6438 -15380 6640 -15363
rect 5680 -15418 6640 -15380
rect 6698 -15380 6900 -15363
rect 7456 -15363 7472 -15346
rect 7902 -15346 8490 -15330
rect 7902 -15363 7918 -15346
rect 7456 -15380 7658 -15363
rect 6698 -15418 7658 -15380
rect 7716 -15380 7918 -15363
rect 8474 -15363 8490 -15346
rect 8920 -15346 9508 -15330
rect 8920 -15363 8936 -15346
rect 8474 -15380 8676 -15363
rect 7716 -15418 8676 -15380
rect 8734 -15380 8936 -15363
rect 9492 -15363 9508 -15346
rect 9938 -15346 10526 -15330
rect 9938 -15363 9954 -15346
rect 9492 -15380 9694 -15363
rect 8734 -15418 9694 -15380
rect 9752 -15380 9954 -15363
rect 10510 -15363 10526 -15346
rect 10956 -15346 11544 -15330
rect 10956 -15363 10972 -15346
rect 10510 -15380 10712 -15363
rect 9752 -15418 10712 -15380
rect 10770 -15380 10972 -15363
rect 11528 -15363 11544 -15346
rect 11974 -15346 12562 -15330
rect 11974 -15363 11990 -15346
rect 11528 -15380 11730 -15363
rect 10770 -15418 11730 -15380
rect 11788 -15380 11990 -15363
rect 12546 -15363 12562 -15346
rect 12992 -15346 13580 -15330
rect 12992 -15363 13008 -15346
rect 12546 -15380 12748 -15363
rect 11788 -15418 12748 -15380
rect 12806 -15380 13008 -15363
rect 13564 -15363 13580 -15346
rect 14010 -15346 14598 -15330
rect 14010 -15363 14026 -15346
rect 13564 -15380 13766 -15363
rect 12806 -15418 13766 -15380
rect 13824 -15380 14026 -15363
rect 14582 -15363 14598 -15346
rect 15028 -15346 15616 -15330
rect 15028 -15363 15044 -15346
rect 14582 -15380 14784 -15363
rect 13824 -15418 14784 -15380
rect 14842 -15380 15044 -15363
rect 15600 -15363 15616 -15346
rect 16046 -15346 16634 -15330
rect 16046 -15363 16062 -15346
rect 15600 -15380 15802 -15363
rect 14842 -15418 15802 -15380
rect 15860 -15380 16062 -15363
rect 16618 -15363 16634 -15346
rect 17064 -15346 17652 -15330
rect 17064 -15363 17080 -15346
rect 16618 -15380 16820 -15363
rect 15860 -15418 16820 -15380
rect 16878 -15380 17080 -15363
rect 17636 -15363 17652 -15346
rect 18082 -15346 18670 -15330
rect 18082 -15363 18098 -15346
rect 17636 -15380 17838 -15363
rect 16878 -15418 17838 -15380
rect 17896 -15380 18098 -15363
rect 18654 -15363 18670 -15346
rect 19100 -15346 19688 -15330
rect 19100 -15363 19116 -15346
rect 18654 -15380 18856 -15363
rect 17896 -15418 18856 -15380
rect 18914 -15380 19116 -15363
rect 19672 -15363 19688 -15346
rect 20118 -15346 20706 -15330
rect 20118 -15363 20134 -15346
rect 19672 -15380 19874 -15363
rect 18914 -15418 19874 -15380
rect 19932 -15380 20134 -15363
rect 20690 -15363 20706 -15346
rect 21136 -15346 21724 -15330
rect 21136 -15363 21152 -15346
rect 20690 -15380 20892 -15363
rect 19932 -15418 20892 -15380
rect 20950 -15380 21152 -15363
rect 21708 -15363 21724 -15346
rect 22154 -15346 22742 -15330
rect 22154 -15363 22170 -15346
rect 21708 -15380 21910 -15363
rect 20950 -15418 21910 -15380
rect 21968 -15380 22170 -15363
rect 22726 -15363 22742 -15346
rect 22726 -15380 22928 -15363
rect 21968 -15418 22928 -15380
rect -9138 -15604 -8178 -15566
rect -9138 -15621 -8936 -15604
rect -8952 -15638 -8936 -15621
rect -8380 -15621 -8178 -15604
rect -8120 -15604 -7160 -15566
rect -8120 -15621 -7918 -15604
rect -8380 -15638 -8364 -15621
rect -8952 -15654 -8364 -15638
rect -7934 -15638 -7918 -15621
rect -7362 -15621 -7160 -15604
rect -7102 -15604 -6142 -15566
rect -7102 -15621 -6900 -15604
rect -7362 -15638 -7346 -15621
rect -7934 -15654 -7346 -15638
rect -6916 -15638 -6900 -15621
rect -6344 -15621 -6142 -15604
rect -6084 -15604 -5124 -15566
rect -6084 -15621 -5882 -15604
rect -6344 -15638 -6328 -15621
rect -6916 -15654 -6328 -15638
rect -5898 -15638 -5882 -15621
rect -5326 -15621 -5124 -15604
rect -5066 -15604 -4106 -15566
rect -5066 -15621 -4864 -15604
rect -5326 -15638 -5310 -15621
rect -5898 -15654 -5310 -15638
rect -4880 -15638 -4864 -15621
rect -4308 -15621 -4106 -15604
rect -4048 -15604 -3088 -15566
rect -4048 -15621 -3846 -15604
rect -4308 -15638 -4292 -15621
rect -4880 -15654 -4292 -15638
rect -3862 -15638 -3846 -15621
rect -3290 -15621 -3088 -15604
rect -3030 -15604 -2070 -15566
rect -3030 -15621 -2828 -15604
rect -3290 -15638 -3274 -15621
rect -3862 -15654 -3274 -15638
rect -2844 -15638 -2828 -15621
rect -2272 -15621 -2070 -15604
rect -2012 -15604 -1052 -15566
rect -2012 -15621 -1810 -15604
rect -2272 -15638 -2256 -15621
rect -2844 -15654 -2256 -15638
rect -1826 -15638 -1810 -15621
rect -1254 -15621 -1052 -15604
rect -994 -15604 -34 -15566
rect -994 -15621 -792 -15604
rect -1254 -15638 -1238 -15621
rect -1826 -15654 -1238 -15638
rect -808 -15638 -792 -15621
rect -236 -15621 -34 -15604
rect -236 -15638 -220 -15621
rect -808 -15654 -220 -15638
rect -8952 -15712 -8364 -15696
rect -8952 -15729 -8936 -15712
rect -9138 -15746 -8936 -15729
rect -8380 -15729 -8364 -15712
rect -7934 -15712 -7346 -15696
rect -7934 -15729 -7918 -15712
rect -8380 -15746 -8178 -15729
rect -9138 -15784 -8178 -15746
rect -8120 -15746 -7918 -15729
rect -7362 -15729 -7346 -15712
rect -6916 -15712 -6328 -15696
rect -6916 -15729 -6900 -15712
rect -7362 -15746 -7160 -15729
rect -8120 -15784 -7160 -15746
rect -7102 -15746 -6900 -15729
rect -6344 -15729 -6328 -15712
rect -5898 -15712 -5310 -15696
rect -5898 -15729 -5882 -15712
rect -6344 -15746 -6142 -15729
rect -7102 -15784 -6142 -15746
rect -6084 -15746 -5882 -15729
rect -5326 -15729 -5310 -15712
rect -4880 -15712 -4292 -15696
rect -4880 -15729 -4864 -15712
rect -5326 -15746 -5124 -15729
rect -6084 -15784 -5124 -15746
rect -5066 -15746 -4864 -15729
rect -4308 -15729 -4292 -15712
rect -3862 -15712 -3274 -15696
rect -3862 -15729 -3846 -15712
rect -4308 -15746 -4106 -15729
rect -5066 -15784 -4106 -15746
rect -4048 -15746 -3846 -15729
rect -3290 -15729 -3274 -15712
rect -2844 -15712 -2256 -15696
rect -2844 -15729 -2828 -15712
rect -3290 -15746 -3088 -15729
rect -4048 -15784 -3088 -15746
rect -3030 -15746 -2828 -15729
rect -2272 -15729 -2256 -15712
rect -1826 -15712 -1238 -15696
rect -1826 -15729 -1810 -15712
rect -2272 -15746 -2070 -15729
rect -3030 -15784 -2070 -15746
rect -2012 -15746 -1810 -15729
rect -1254 -15729 -1238 -15712
rect -808 -15712 -220 -15696
rect -808 -15729 -792 -15712
rect -1254 -15746 -1052 -15729
rect -2012 -15784 -1052 -15746
rect -994 -15746 -792 -15729
rect -236 -15729 -220 -15712
rect -236 -15746 -34 -15729
rect -994 -15784 -34 -15746
rect 2626 -16056 3586 -16018
rect 2626 -16073 2828 -16056
rect 2812 -16090 2828 -16073
rect 3384 -16073 3586 -16056
rect 3644 -16056 4604 -16018
rect 3644 -16073 3846 -16056
rect 3384 -16090 3400 -16073
rect 2812 -16106 3400 -16090
rect 3830 -16090 3846 -16073
rect 4402 -16073 4604 -16056
rect 4662 -16056 5622 -16018
rect 4662 -16073 4864 -16056
rect 4402 -16090 4418 -16073
rect 3830 -16106 4418 -16090
rect 4848 -16090 4864 -16073
rect 5420 -16073 5622 -16056
rect 5680 -16056 6640 -16018
rect 5680 -16073 5882 -16056
rect 5420 -16090 5436 -16073
rect 4848 -16106 5436 -16090
rect 5866 -16090 5882 -16073
rect 6438 -16073 6640 -16056
rect 6698 -16056 7658 -16018
rect 6698 -16073 6900 -16056
rect 6438 -16090 6454 -16073
rect 5866 -16106 6454 -16090
rect 6884 -16090 6900 -16073
rect 7456 -16073 7658 -16056
rect 7716 -16056 8676 -16018
rect 7716 -16073 7918 -16056
rect 7456 -16090 7472 -16073
rect 6884 -16106 7472 -16090
rect 7902 -16090 7918 -16073
rect 8474 -16073 8676 -16056
rect 8734 -16056 9694 -16018
rect 8734 -16073 8936 -16056
rect 8474 -16090 8490 -16073
rect 7902 -16106 8490 -16090
rect 8920 -16090 8936 -16073
rect 9492 -16073 9694 -16056
rect 9752 -16056 10712 -16018
rect 9752 -16073 9954 -16056
rect 9492 -16090 9508 -16073
rect 8920 -16106 9508 -16090
rect 9938 -16090 9954 -16073
rect 10510 -16073 10712 -16056
rect 10770 -16056 11730 -16018
rect 10770 -16073 10972 -16056
rect 10510 -16090 10526 -16073
rect 9938 -16106 10526 -16090
rect 10956 -16090 10972 -16073
rect 11528 -16073 11730 -16056
rect 11788 -16056 12748 -16018
rect 11788 -16073 11990 -16056
rect 11528 -16090 11544 -16073
rect 10956 -16106 11544 -16090
rect 11974 -16090 11990 -16073
rect 12546 -16073 12748 -16056
rect 12806 -16056 13766 -16018
rect 12806 -16073 13008 -16056
rect 12546 -16090 12562 -16073
rect 11974 -16106 12562 -16090
rect 12992 -16090 13008 -16073
rect 13564 -16073 13766 -16056
rect 13824 -16056 14784 -16018
rect 13824 -16073 14026 -16056
rect 13564 -16090 13580 -16073
rect 12992 -16106 13580 -16090
rect 14010 -16090 14026 -16073
rect 14582 -16073 14784 -16056
rect 14842 -16056 15802 -16018
rect 14842 -16073 15044 -16056
rect 14582 -16090 14598 -16073
rect 14010 -16106 14598 -16090
rect 15028 -16090 15044 -16073
rect 15600 -16073 15802 -16056
rect 15860 -16056 16820 -16018
rect 15860 -16073 16062 -16056
rect 15600 -16090 15616 -16073
rect 15028 -16106 15616 -16090
rect 16046 -16090 16062 -16073
rect 16618 -16073 16820 -16056
rect 16878 -16056 17838 -16018
rect 16878 -16073 17080 -16056
rect 16618 -16090 16634 -16073
rect 16046 -16106 16634 -16090
rect 17064 -16090 17080 -16073
rect 17636 -16073 17838 -16056
rect 17896 -16056 18856 -16018
rect 17896 -16073 18098 -16056
rect 17636 -16090 17652 -16073
rect 17064 -16106 17652 -16090
rect 18082 -16090 18098 -16073
rect 18654 -16073 18856 -16056
rect 18914 -16056 19874 -16018
rect 18914 -16073 19116 -16056
rect 18654 -16090 18670 -16073
rect 18082 -16106 18670 -16090
rect 19100 -16090 19116 -16073
rect 19672 -16073 19874 -16056
rect 19932 -16056 20892 -16018
rect 19932 -16073 20134 -16056
rect 19672 -16090 19688 -16073
rect 19100 -16106 19688 -16090
rect 20118 -16090 20134 -16073
rect 20690 -16073 20892 -16056
rect 20950 -16056 21910 -16018
rect 20950 -16073 21152 -16056
rect 20690 -16090 20706 -16073
rect 20118 -16106 20706 -16090
rect 21136 -16090 21152 -16073
rect 21708 -16073 21910 -16056
rect 21968 -16056 22928 -16018
rect 21968 -16073 22170 -16056
rect 21708 -16090 21724 -16073
rect 21136 -16106 21724 -16090
rect 22154 -16090 22170 -16073
rect 22726 -16073 22928 -16056
rect 22726 -16090 22742 -16073
rect 22154 -16106 22742 -16090
rect -9138 -16422 -8178 -16384
rect -9138 -16439 -8936 -16422
rect -8952 -16456 -8936 -16439
rect -8380 -16439 -8178 -16422
rect -8120 -16422 -7160 -16384
rect -8120 -16439 -7918 -16422
rect -8380 -16456 -8364 -16439
rect -8952 -16472 -8364 -16456
rect -7934 -16456 -7918 -16439
rect -7362 -16439 -7160 -16422
rect -7102 -16422 -6142 -16384
rect -7102 -16439 -6900 -16422
rect -7362 -16456 -7346 -16439
rect -7934 -16472 -7346 -16456
rect -6916 -16456 -6900 -16439
rect -6344 -16439 -6142 -16422
rect -6084 -16422 -5124 -16384
rect -6084 -16439 -5882 -16422
rect -6344 -16456 -6328 -16439
rect -6916 -16472 -6328 -16456
rect -5898 -16456 -5882 -16439
rect -5326 -16439 -5124 -16422
rect -5066 -16422 -4106 -16384
rect -5066 -16439 -4864 -16422
rect -5326 -16456 -5310 -16439
rect -5898 -16472 -5310 -16456
rect -4880 -16456 -4864 -16439
rect -4308 -16439 -4106 -16422
rect -4048 -16422 -3088 -16384
rect -4048 -16439 -3846 -16422
rect -4308 -16456 -4292 -16439
rect -4880 -16472 -4292 -16456
rect -3862 -16456 -3846 -16439
rect -3290 -16439 -3088 -16422
rect -3030 -16422 -2070 -16384
rect -3030 -16439 -2828 -16422
rect -3290 -16456 -3274 -16439
rect -3862 -16472 -3274 -16456
rect -2844 -16456 -2828 -16439
rect -2272 -16439 -2070 -16422
rect -2012 -16422 -1052 -16384
rect -2012 -16439 -1810 -16422
rect -2272 -16456 -2256 -16439
rect -2844 -16472 -2256 -16456
rect -1826 -16456 -1810 -16439
rect -1254 -16439 -1052 -16422
rect -994 -16422 -34 -16384
rect -994 -16439 -792 -16422
rect -1254 -16456 -1238 -16439
rect -1826 -16472 -1238 -16456
rect -808 -16456 -792 -16439
rect -236 -16439 -34 -16422
rect -236 -16456 -220 -16439
rect -808 -16472 -220 -16456
rect -8952 -16530 -8364 -16514
rect -8952 -16547 -8936 -16530
rect -9138 -16564 -8936 -16547
rect -8380 -16547 -8364 -16530
rect -7934 -16530 -7346 -16514
rect -7934 -16547 -7918 -16530
rect -8380 -16564 -8178 -16547
rect -9138 -16602 -8178 -16564
rect -8120 -16564 -7918 -16547
rect -7362 -16547 -7346 -16530
rect -6916 -16530 -6328 -16514
rect -6916 -16547 -6900 -16530
rect -7362 -16564 -7160 -16547
rect -8120 -16602 -7160 -16564
rect -7102 -16564 -6900 -16547
rect -6344 -16547 -6328 -16530
rect -5898 -16530 -5310 -16514
rect -5898 -16547 -5882 -16530
rect -6344 -16564 -6142 -16547
rect -7102 -16602 -6142 -16564
rect -6084 -16564 -5882 -16547
rect -5326 -16547 -5310 -16530
rect -4880 -16530 -4292 -16514
rect -4880 -16547 -4864 -16530
rect -5326 -16564 -5124 -16547
rect -6084 -16602 -5124 -16564
rect -5066 -16564 -4864 -16547
rect -4308 -16547 -4292 -16530
rect -3862 -16530 -3274 -16514
rect -3862 -16547 -3846 -16530
rect -4308 -16564 -4106 -16547
rect -5066 -16602 -4106 -16564
rect -4048 -16564 -3846 -16547
rect -3290 -16547 -3274 -16530
rect -2844 -16530 -2256 -16514
rect -2844 -16547 -2828 -16530
rect -3290 -16564 -3088 -16547
rect -4048 -16602 -3088 -16564
rect -3030 -16564 -2828 -16547
rect -2272 -16547 -2256 -16530
rect -1826 -16530 -1238 -16514
rect -1826 -16547 -1810 -16530
rect -2272 -16564 -2070 -16547
rect -3030 -16602 -2070 -16564
rect -2012 -16564 -1810 -16547
rect -1254 -16547 -1238 -16530
rect -808 -16530 -220 -16514
rect -808 -16547 -792 -16530
rect -1254 -16564 -1052 -16547
rect -2012 -16602 -1052 -16564
rect -994 -16564 -792 -16547
rect -236 -16547 -220 -16530
rect -236 -16564 -34 -16547
rect -994 -16602 -34 -16564
rect 2812 -16580 3400 -16564
rect 2812 -16597 2828 -16580
rect 2626 -16614 2828 -16597
rect 3384 -16597 3400 -16580
rect 3830 -16580 4418 -16564
rect 3830 -16597 3846 -16580
rect 3384 -16614 3586 -16597
rect 2626 -16652 3586 -16614
rect 3644 -16614 3846 -16597
rect 4402 -16597 4418 -16580
rect 4848 -16580 5436 -16564
rect 4848 -16597 4864 -16580
rect 4402 -16614 4604 -16597
rect 3644 -16652 4604 -16614
rect 4662 -16614 4864 -16597
rect 5420 -16597 5436 -16580
rect 5866 -16580 6454 -16564
rect 5866 -16597 5882 -16580
rect 5420 -16614 5622 -16597
rect 4662 -16652 5622 -16614
rect 5680 -16614 5882 -16597
rect 6438 -16597 6454 -16580
rect 6884 -16580 7472 -16564
rect 6884 -16597 6900 -16580
rect 6438 -16614 6640 -16597
rect 5680 -16652 6640 -16614
rect 6698 -16614 6900 -16597
rect 7456 -16597 7472 -16580
rect 7902 -16580 8490 -16564
rect 7902 -16597 7918 -16580
rect 7456 -16614 7658 -16597
rect 6698 -16652 7658 -16614
rect 7716 -16614 7918 -16597
rect 8474 -16597 8490 -16580
rect 8920 -16580 9508 -16564
rect 8920 -16597 8936 -16580
rect 8474 -16614 8676 -16597
rect 7716 -16652 8676 -16614
rect 8734 -16614 8936 -16597
rect 9492 -16597 9508 -16580
rect 9938 -16580 10526 -16564
rect 9938 -16597 9954 -16580
rect 9492 -16614 9694 -16597
rect 8734 -16652 9694 -16614
rect 9752 -16614 9954 -16597
rect 10510 -16597 10526 -16580
rect 10956 -16580 11544 -16564
rect 10956 -16597 10972 -16580
rect 10510 -16614 10712 -16597
rect 9752 -16652 10712 -16614
rect 10770 -16614 10972 -16597
rect 11528 -16597 11544 -16580
rect 11974 -16580 12562 -16564
rect 11974 -16597 11990 -16580
rect 11528 -16614 11730 -16597
rect 10770 -16652 11730 -16614
rect 11788 -16614 11990 -16597
rect 12546 -16597 12562 -16580
rect 12992 -16580 13580 -16564
rect 12992 -16597 13008 -16580
rect 12546 -16614 12748 -16597
rect 11788 -16652 12748 -16614
rect 12806 -16614 13008 -16597
rect 13564 -16597 13580 -16580
rect 14010 -16580 14598 -16564
rect 14010 -16597 14026 -16580
rect 13564 -16614 13766 -16597
rect 12806 -16652 13766 -16614
rect 13824 -16614 14026 -16597
rect 14582 -16597 14598 -16580
rect 15028 -16580 15616 -16564
rect 15028 -16597 15044 -16580
rect 14582 -16614 14784 -16597
rect 13824 -16652 14784 -16614
rect 14842 -16614 15044 -16597
rect 15600 -16597 15616 -16580
rect 16046 -16580 16634 -16564
rect 16046 -16597 16062 -16580
rect 15600 -16614 15802 -16597
rect 14842 -16652 15802 -16614
rect 15860 -16614 16062 -16597
rect 16618 -16597 16634 -16580
rect 17064 -16580 17652 -16564
rect 17064 -16597 17080 -16580
rect 16618 -16614 16820 -16597
rect 15860 -16652 16820 -16614
rect 16878 -16614 17080 -16597
rect 17636 -16597 17652 -16580
rect 18082 -16580 18670 -16564
rect 18082 -16597 18098 -16580
rect 17636 -16614 17838 -16597
rect 16878 -16652 17838 -16614
rect 17896 -16614 18098 -16597
rect 18654 -16597 18670 -16580
rect 19100 -16580 19688 -16564
rect 19100 -16597 19116 -16580
rect 18654 -16614 18856 -16597
rect 17896 -16652 18856 -16614
rect 18914 -16614 19116 -16597
rect 19672 -16597 19688 -16580
rect 20118 -16580 20706 -16564
rect 20118 -16597 20134 -16580
rect 19672 -16614 19874 -16597
rect 18914 -16652 19874 -16614
rect 19932 -16614 20134 -16597
rect 20690 -16597 20706 -16580
rect 21136 -16580 21724 -16564
rect 21136 -16597 21152 -16580
rect 20690 -16614 20892 -16597
rect 19932 -16652 20892 -16614
rect 20950 -16614 21152 -16597
rect 21708 -16597 21724 -16580
rect 22154 -16580 22742 -16564
rect 22154 -16597 22170 -16580
rect 21708 -16614 21910 -16597
rect 20950 -16652 21910 -16614
rect 21968 -16614 22170 -16597
rect 22726 -16597 22742 -16580
rect 22726 -16614 22928 -16597
rect 21968 -16652 22928 -16614
rect -9138 -17240 -8178 -17202
rect -9138 -17257 -8936 -17240
rect -8952 -17274 -8936 -17257
rect -8380 -17257 -8178 -17240
rect -8120 -17240 -7160 -17202
rect -8120 -17257 -7918 -17240
rect -8380 -17274 -8364 -17257
rect -8952 -17290 -8364 -17274
rect -7934 -17274 -7918 -17257
rect -7362 -17257 -7160 -17240
rect -7102 -17240 -6142 -17202
rect -7102 -17257 -6900 -17240
rect -7362 -17274 -7346 -17257
rect -7934 -17290 -7346 -17274
rect -6916 -17274 -6900 -17257
rect -6344 -17257 -6142 -17240
rect -6084 -17240 -5124 -17202
rect -6084 -17257 -5882 -17240
rect -6344 -17274 -6328 -17257
rect -6916 -17290 -6328 -17274
rect -5898 -17274 -5882 -17257
rect -5326 -17257 -5124 -17240
rect -5066 -17240 -4106 -17202
rect -5066 -17257 -4864 -17240
rect -5326 -17274 -5310 -17257
rect -5898 -17290 -5310 -17274
rect -4880 -17274 -4864 -17257
rect -4308 -17257 -4106 -17240
rect -4048 -17240 -3088 -17202
rect -4048 -17257 -3846 -17240
rect -4308 -17274 -4292 -17257
rect -4880 -17290 -4292 -17274
rect -3862 -17274 -3846 -17257
rect -3290 -17257 -3088 -17240
rect -3030 -17240 -2070 -17202
rect -3030 -17257 -2828 -17240
rect -3290 -17274 -3274 -17257
rect -3862 -17290 -3274 -17274
rect -2844 -17274 -2828 -17257
rect -2272 -17257 -2070 -17240
rect -2012 -17240 -1052 -17202
rect -2012 -17257 -1810 -17240
rect -2272 -17274 -2256 -17257
rect -2844 -17290 -2256 -17274
rect -1826 -17274 -1810 -17257
rect -1254 -17257 -1052 -17240
rect -994 -17240 -34 -17202
rect -994 -17257 -792 -17240
rect -1254 -17274 -1238 -17257
rect -1826 -17290 -1238 -17274
rect -808 -17274 -792 -17257
rect -236 -17257 -34 -17240
rect -236 -17274 -220 -17257
rect -808 -17290 -220 -17274
rect 2626 -17290 3586 -17252
rect 2626 -17307 2828 -17290
rect 2812 -17324 2828 -17307
rect 3384 -17307 3586 -17290
rect 3644 -17290 4604 -17252
rect 3644 -17307 3846 -17290
rect 3384 -17324 3400 -17307
rect -8952 -17348 -8364 -17332
rect -8952 -17365 -8936 -17348
rect -9138 -17382 -8936 -17365
rect -8380 -17365 -8364 -17348
rect -7934 -17348 -7346 -17332
rect -7934 -17365 -7918 -17348
rect -8380 -17382 -8178 -17365
rect -9138 -17420 -8178 -17382
rect -8120 -17382 -7918 -17365
rect -7362 -17365 -7346 -17348
rect -6916 -17348 -6328 -17332
rect -6916 -17365 -6900 -17348
rect -7362 -17382 -7160 -17365
rect -8120 -17420 -7160 -17382
rect -7102 -17382 -6900 -17365
rect -6344 -17365 -6328 -17348
rect -5898 -17348 -5310 -17332
rect -5898 -17365 -5882 -17348
rect -6344 -17382 -6142 -17365
rect -7102 -17420 -6142 -17382
rect -6084 -17382 -5882 -17365
rect -5326 -17365 -5310 -17348
rect -4880 -17348 -4292 -17332
rect -4880 -17365 -4864 -17348
rect -5326 -17382 -5124 -17365
rect -6084 -17420 -5124 -17382
rect -5066 -17382 -4864 -17365
rect -4308 -17365 -4292 -17348
rect -3862 -17348 -3274 -17332
rect -3862 -17365 -3846 -17348
rect -4308 -17382 -4106 -17365
rect -5066 -17420 -4106 -17382
rect -4048 -17382 -3846 -17365
rect -3290 -17365 -3274 -17348
rect -2844 -17348 -2256 -17332
rect -2844 -17365 -2828 -17348
rect -3290 -17382 -3088 -17365
rect -4048 -17420 -3088 -17382
rect -3030 -17382 -2828 -17365
rect -2272 -17365 -2256 -17348
rect -1826 -17348 -1238 -17332
rect -1826 -17365 -1810 -17348
rect -2272 -17382 -2070 -17365
rect -3030 -17420 -2070 -17382
rect -2012 -17382 -1810 -17365
rect -1254 -17365 -1238 -17348
rect -808 -17348 -220 -17332
rect 2812 -17340 3400 -17324
rect 3830 -17324 3846 -17307
rect 4402 -17307 4604 -17290
rect 4662 -17290 5622 -17252
rect 4662 -17307 4864 -17290
rect 4402 -17324 4418 -17307
rect 3830 -17340 4418 -17324
rect 4848 -17324 4864 -17307
rect 5420 -17307 5622 -17290
rect 5680 -17290 6640 -17252
rect 5680 -17307 5882 -17290
rect 5420 -17324 5436 -17307
rect 4848 -17340 5436 -17324
rect 5866 -17324 5882 -17307
rect 6438 -17307 6640 -17290
rect 6698 -17290 7658 -17252
rect 6698 -17307 6900 -17290
rect 6438 -17324 6454 -17307
rect 5866 -17340 6454 -17324
rect 6884 -17324 6900 -17307
rect 7456 -17307 7658 -17290
rect 7716 -17290 8676 -17252
rect 7716 -17307 7918 -17290
rect 7456 -17324 7472 -17307
rect 6884 -17340 7472 -17324
rect 7902 -17324 7918 -17307
rect 8474 -17307 8676 -17290
rect 8734 -17290 9694 -17252
rect 8734 -17307 8936 -17290
rect 8474 -17324 8490 -17307
rect 7902 -17340 8490 -17324
rect 8920 -17324 8936 -17307
rect 9492 -17307 9694 -17290
rect 9752 -17290 10712 -17252
rect 9752 -17307 9954 -17290
rect 9492 -17324 9508 -17307
rect 8920 -17340 9508 -17324
rect 9938 -17324 9954 -17307
rect 10510 -17307 10712 -17290
rect 10770 -17290 11730 -17252
rect 10770 -17307 10972 -17290
rect 10510 -17324 10526 -17307
rect 9938 -17340 10526 -17324
rect 10956 -17324 10972 -17307
rect 11528 -17307 11730 -17290
rect 11788 -17290 12748 -17252
rect 11788 -17307 11990 -17290
rect 11528 -17324 11544 -17307
rect 10956 -17340 11544 -17324
rect 11974 -17324 11990 -17307
rect 12546 -17307 12748 -17290
rect 12806 -17290 13766 -17252
rect 12806 -17307 13008 -17290
rect 12546 -17324 12562 -17307
rect 11974 -17340 12562 -17324
rect 12992 -17324 13008 -17307
rect 13564 -17307 13766 -17290
rect 13824 -17290 14784 -17252
rect 13824 -17307 14026 -17290
rect 13564 -17324 13580 -17307
rect 12992 -17340 13580 -17324
rect 14010 -17324 14026 -17307
rect 14582 -17307 14784 -17290
rect 14842 -17290 15802 -17252
rect 14842 -17307 15044 -17290
rect 14582 -17324 14598 -17307
rect 14010 -17340 14598 -17324
rect 15028 -17324 15044 -17307
rect 15600 -17307 15802 -17290
rect 15860 -17290 16820 -17252
rect 15860 -17307 16062 -17290
rect 15600 -17324 15616 -17307
rect 15028 -17340 15616 -17324
rect 16046 -17324 16062 -17307
rect 16618 -17307 16820 -17290
rect 16878 -17290 17838 -17252
rect 16878 -17307 17080 -17290
rect 16618 -17324 16634 -17307
rect 16046 -17340 16634 -17324
rect 17064 -17324 17080 -17307
rect 17636 -17307 17838 -17290
rect 17896 -17290 18856 -17252
rect 17896 -17307 18098 -17290
rect 17636 -17324 17652 -17307
rect 17064 -17340 17652 -17324
rect 18082 -17324 18098 -17307
rect 18654 -17307 18856 -17290
rect 18914 -17290 19874 -17252
rect 18914 -17307 19116 -17290
rect 18654 -17324 18670 -17307
rect 18082 -17340 18670 -17324
rect 19100 -17324 19116 -17307
rect 19672 -17307 19874 -17290
rect 19932 -17290 20892 -17252
rect 19932 -17307 20134 -17290
rect 19672 -17324 19688 -17307
rect 19100 -17340 19688 -17324
rect 20118 -17324 20134 -17307
rect 20690 -17307 20892 -17290
rect 20950 -17290 21910 -17252
rect 20950 -17307 21152 -17290
rect 20690 -17324 20706 -17307
rect 20118 -17340 20706 -17324
rect 21136 -17324 21152 -17307
rect 21708 -17307 21910 -17290
rect 21968 -17290 22928 -17252
rect 21968 -17307 22170 -17290
rect 21708 -17324 21724 -17307
rect 21136 -17340 21724 -17324
rect 22154 -17324 22170 -17307
rect 22726 -17307 22928 -17290
rect 22726 -17324 22742 -17307
rect 22154 -17340 22742 -17324
rect -808 -17365 -792 -17348
rect -1254 -17382 -1052 -17365
rect -2012 -17420 -1052 -17382
rect -994 -17382 -792 -17365
rect -236 -17365 -220 -17348
rect -236 -17382 -34 -17365
rect -994 -17420 -34 -17382
rect 2812 -17812 3400 -17796
rect 2812 -17829 2828 -17812
rect 2626 -17846 2828 -17829
rect 3384 -17829 3400 -17812
rect 3830 -17812 4418 -17796
rect 3830 -17829 3846 -17812
rect 3384 -17846 3586 -17829
rect 2626 -17884 3586 -17846
rect 3644 -17846 3846 -17829
rect 4402 -17829 4418 -17812
rect 4848 -17812 5436 -17796
rect 4848 -17829 4864 -17812
rect 4402 -17846 4604 -17829
rect 3644 -17884 4604 -17846
rect 4662 -17846 4864 -17829
rect 5420 -17829 5436 -17812
rect 5866 -17812 6454 -17796
rect 5866 -17829 5882 -17812
rect 5420 -17846 5622 -17829
rect 4662 -17884 5622 -17846
rect 5680 -17846 5882 -17829
rect 6438 -17829 6454 -17812
rect 6884 -17812 7472 -17796
rect 6884 -17829 6900 -17812
rect 6438 -17846 6640 -17829
rect 5680 -17884 6640 -17846
rect 6698 -17846 6900 -17829
rect 7456 -17829 7472 -17812
rect 7902 -17812 8490 -17796
rect 7902 -17829 7918 -17812
rect 7456 -17846 7658 -17829
rect 6698 -17884 7658 -17846
rect 7716 -17846 7918 -17829
rect 8474 -17829 8490 -17812
rect 8920 -17812 9508 -17796
rect 8920 -17829 8936 -17812
rect 8474 -17846 8676 -17829
rect 7716 -17884 8676 -17846
rect 8734 -17846 8936 -17829
rect 9492 -17829 9508 -17812
rect 9938 -17812 10526 -17796
rect 9938 -17829 9954 -17812
rect 9492 -17846 9694 -17829
rect 8734 -17884 9694 -17846
rect 9752 -17846 9954 -17829
rect 10510 -17829 10526 -17812
rect 10956 -17812 11544 -17796
rect 10956 -17829 10972 -17812
rect 10510 -17846 10712 -17829
rect 9752 -17884 10712 -17846
rect 10770 -17846 10972 -17829
rect 11528 -17829 11544 -17812
rect 11974 -17812 12562 -17796
rect 11974 -17829 11990 -17812
rect 11528 -17846 11730 -17829
rect 10770 -17884 11730 -17846
rect 11788 -17846 11990 -17829
rect 12546 -17829 12562 -17812
rect 12992 -17812 13580 -17796
rect 12992 -17829 13008 -17812
rect 12546 -17846 12748 -17829
rect 11788 -17884 12748 -17846
rect 12806 -17846 13008 -17829
rect 13564 -17829 13580 -17812
rect 14010 -17812 14598 -17796
rect 14010 -17829 14026 -17812
rect 13564 -17846 13766 -17829
rect 12806 -17884 13766 -17846
rect 13824 -17846 14026 -17829
rect 14582 -17829 14598 -17812
rect 15028 -17812 15616 -17796
rect 15028 -17829 15044 -17812
rect 14582 -17846 14784 -17829
rect 13824 -17884 14784 -17846
rect 14842 -17846 15044 -17829
rect 15600 -17829 15616 -17812
rect 16046 -17812 16634 -17796
rect 16046 -17829 16062 -17812
rect 15600 -17846 15802 -17829
rect 14842 -17884 15802 -17846
rect 15860 -17846 16062 -17829
rect 16618 -17829 16634 -17812
rect 17064 -17812 17652 -17796
rect 17064 -17829 17080 -17812
rect 16618 -17846 16820 -17829
rect 15860 -17884 16820 -17846
rect 16878 -17846 17080 -17829
rect 17636 -17829 17652 -17812
rect 18082 -17812 18670 -17796
rect 18082 -17829 18098 -17812
rect 17636 -17846 17838 -17829
rect 16878 -17884 17838 -17846
rect 17896 -17846 18098 -17829
rect 18654 -17829 18670 -17812
rect 19100 -17812 19688 -17796
rect 19100 -17829 19116 -17812
rect 18654 -17846 18856 -17829
rect 17896 -17884 18856 -17846
rect 18914 -17846 19116 -17829
rect 19672 -17829 19688 -17812
rect 20118 -17812 20706 -17796
rect 20118 -17829 20134 -17812
rect 19672 -17846 19874 -17829
rect 18914 -17884 19874 -17846
rect 19932 -17846 20134 -17829
rect 20690 -17829 20706 -17812
rect 21136 -17812 21724 -17796
rect 21136 -17829 21152 -17812
rect 20690 -17846 20892 -17829
rect 19932 -17884 20892 -17846
rect 20950 -17846 21152 -17829
rect 21708 -17829 21724 -17812
rect 22154 -17812 22742 -17796
rect 22154 -17829 22170 -17812
rect 21708 -17846 21910 -17829
rect 20950 -17884 21910 -17846
rect 21968 -17846 22170 -17829
rect 22726 -17829 22742 -17812
rect 22726 -17846 22928 -17829
rect 21968 -17884 22928 -17846
rect -9138 -18058 -8178 -18020
rect -9138 -18075 -8936 -18058
rect -8952 -18092 -8936 -18075
rect -8380 -18075 -8178 -18058
rect -8120 -18058 -7160 -18020
rect -8120 -18075 -7918 -18058
rect -8380 -18092 -8364 -18075
rect -8952 -18108 -8364 -18092
rect -7934 -18092 -7918 -18075
rect -7362 -18075 -7160 -18058
rect -7102 -18058 -6142 -18020
rect -7102 -18075 -6900 -18058
rect -7362 -18092 -7346 -18075
rect -7934 -18108 -7346 -18092
rect -6916 -18092 -6900 -18075
rect -6344 -18075 -6142 -18058
rect -6084 -18058 -5124 -18020
rect -6084 -18075 -5882 -18058
rect -6344 -18092 -6328 -18075
rect -6916 -18108 -6328 -18092
rect -5898 -18092 -5882 -18075
rect -5326 -18075 -5124 -18058
rect -5066 -18058 -4106 -18020
rect -5066 -18075 -4864 -18058
rect -5326 -18092 -5310 -18075
rect -5898 -18108 -5310 -18092
rect -4880 -18092 -4864 -18075
rect -4308 -18075 -4106 -18058
rect -4048 -18058 -3088 -18020
rect -4048 -18075 -3846 -18058
rect -4308 -18092 -4292 -18075
rect -4880 -18108 -4292 -18092
rect -3862 -18092 -3846 -18075
rect -3290 -18075 -3088 -18058
rect -3030 -18058 -2070 -18020
rect -3030 -18075 -2828 -18058
rect -3290 -18092 -3274 -18075
rect -3862 -18108 -3274 -18092
rect -2844 -18092 -2828 -18075
rect -2272 -18075 -2070 -18058
rect -2012 -18058 -1052 -18020
rect -2012 -18075 -1810 -18058
rect -2272 -18092 -2256 -18075
rect -2844 -18108 -2256 -18092
rect -1826 -18092 -1810 -18075
rect -1254 -18075 -1052 -18058
rect -994 -18058 -34 -18020
rect -994 -18075 -792 -18058
rect -1254 -18092 -1238 -18075
rect -1826 -18108 -1238 -18092
rect -808 -18092 -792 -18075
rect -236 -18075 -34 -18058
rect -236 -18092 -220 -18075
rect -808 -18108 -220 -18092
rect -8952 -18166 -8364 -18150
rect -8952 -18183 -8936 -18166
rect -9138 -18200 -8936 -18183
rect -8380 -18183 -8364 -18166
rect -7934 -18166 -7346 -18150
rect -7934 -18183 -7918 -18166
rect -8380 -18200 -8178 -18183
rect -9138 -18238 -8178 -18200
rect -8120 -18200 -7918 -18183
rect -7362 -18183 -7346 -18166
rect -6916 -18166 -6328 -18150
rect -6916 -18183 -6900 -18166
rect -7362 -18200 -7160 -18183
rect -8120 -18238 -7160 -18200
rect -7102 -18200 -6900 -18183
rect -6344 -18183 -6328 -18166
rect -5898 -18166 -5310 -18150
rect -5898 -18183 -5882 -18166
rect -6344 -18200 -6142 -18183
rect -7102 -18238 -6142 -18200
rect -6084 -18200 -5882 -18183
rect -5326 -18183 -5310 -18166
rect -4880 -18166 -4292 -18150
rect -4880 -18183 -4864 -18166
rect -5326 -18200 -5124 -18183
rect -6084 -18238 -5124 -18200
rect -5066 -18200 -4864 -18183
rect -4308 -18183 -4292 -18166
rect -3862 -18166 -3274 -18150
rect -3862 -18183 -3846 -18166
rect -4308 -18200 -4106 -18183
rect -5066 -18238 -4106 -18200
rect -4048 -18200 -3846 -18183
rect -3290 -18183 -3274 -18166
rect -2844 -18166 -2256 -18150
rect -2844 -18183 -2828 -18166
rect -3290 -18200 -3088 -18183
rect -4048 -18238 -3088 -18200
rect -3030 -18200 -2828 -18183
rect -2272 -18183 -2256 -18166
rect -1826 -18166 -1238 -18150
rect -1826 -18183 -1810 -18166
rect -2272 -18200 -2070 -18183
rect -3030 -18238 -2070 -18200
rect -2012 -18200 -1810 -18183
rect -1254 -18183 -1238 -18166
rect -808 -18166 -220 -18150
rect -808 -18183 -792 -18166
rect -1254 -18200 -1052 -18183
rect -2012 -18238 -1052 -18200
rect -994 -18200 -792 -18183
rect -236 -18183 -220 -18166
rect -236 -18200 -34 -18183
rect -994 -18238 -34 -18200
rect 2626 -18522 3586 -18484
rect 2626 -18539 2828 -18522
rect 2812 -18556 2828 -18539
rect 3384 -18539 3586 -18522
rect 3644 -18522 4604 -18484
rect 3644 -18539 3846 -18522
rect 3384 -18556 3400 -18539
rect 2812 -18572 3400 -18556
rect 3830 -18556 3846 -18539
rect 4402 -18539 4604 -18522
rect 4662 -18522 5622 -18484
rect 4662 -18539 4864 -18522
rect 4402 -18556 4418 -18539
rect 3830 -18572 4418 -18556
rect 4848 -18556 4864 -18539
rect 5420 -18539 5622 -18522
rect 5680 -18522 6640 -18484
rect 5680 -18539 5882 -18522
rect 5420 -18556 5436 -18539
rect 4848 -18572 5436 -18556
rect 5866 -18556 5882 -18539
rect 6438 -18539 6640 -18522
rect 6698 -18522 7658 -18484
rect 6698 -18539 6900 -18522
rect 6438 -18556 6454 -18539
rect 5866 -18572 6454 -18556
rect 6884 -18556 6900 -18539
rect 7456 -18539 7658 -18522
rect 7716 -18522 8676 -18484
rect 7716 -18539 7918 -18522
rect 7456 -18556 7472 -18539
rect 6884 -18572 7472 -18556
rect 7902 -18556 7918 -18539
rect 8474 -18539 8676 -18522
rect 8734 -18522 9694 -18484
rect 8734 -18539 8936 -18522
rect 8474 -18556 8490 -18539
rect 7902 -18572 8490 -18556
rect 8920 -18556 8936 -18539
rect 9492 -18539 9694 -18522
rect 9752 -18522 10712 -18484
rect 9752 -18539 9954 -18522
rect 9492 -18556 9508 -18539
rect 8920 -18572 9508 -18556
rect 9938 -18556 9954 -18539
rect 10510 -18539 10712 -18522
rect 10770 -18522 11730 -18484
rect 10770 -18539 10972 -18522
rect 10510 -18556 10526 -18539
rect 9938 -18572 10526 -18556
rect 10956 -18556 10972 -18539
rect 11528 -18539 11730 -18522
rect 11788 -18522 12748 -18484
rect 11788 -18539 11990 -18522
rect 11528 -18556 11544 -18539
rect 10956 -18572 11544 -18556
rect 11974 -18556 11990 -18539
rect 12546 -18539 12748 -18522
rect 12806 -18522 13766 -18484
rect 12806 -18539 13008 -18522
rect 12546 -18556 12562 -18539
rect 11974 -18572 12562 -18556
rect 12992 -18556 13008 -18539
rect 13564 -18539 13766 -18522
rect 13824 -18522 14784 -18484
rect 13824 -18539 14026 -18522
rect 13564 -18556 13580 -18539
rect 12992 -18572 13580 -18556
rect 14010 -18556 14026 -18539
rect 14582 -18539 14784 -18522
rect 14842 -18522 15802 -18484
rect 14842 -18539 15044 -18522
rect 14582 -18556 14598 -18539
rect 14010 -18572 14598 -18556
rect 15028 -18556 15044 -18539
rect 15600 -18539 15802 -18522
rect 15860 -18522 16820 -18484
rect 15860 -18539 16062 -18522
rect 15600 -18556 15616 -18539
rect 15028 -18572 15616 -18556
rect 16046 -18556 16062 -18539
rect 16618 -18539 16820 -18522
rect 16878 -18522 17838 -18484
rect 16878 -18539 17080 -18522
rect 16618 -18556 16634 -18539
rect 16046 -18572 16634 -18556
rect 17064 -18556 17080 -18539
rect 17636 -18539 17838 -18522
rect 17896 -18522 18856 -18484
rect 17896 -18539 18098 -18522
rect 17636 -18556 17652 -18539
rect 17064 -18572 17652 -18556
rect 18082 -18556 18098 -18539
rect 18654 -18539 18856 -18522
rect 18914 -18522 19874 -18484
rect 18914 -18539 19116 -18522
rect 18654 -18556 18670 -18539
rect 18082 -18572 18670 -18556
rect 19100 -18556 19116 -18539
rect 19672 -18539 19874 -18522
rect 19932 -18522 20892 -18484
rect 19932 -18539 20134 -18522
rect 19672 -18556 19688 -18539
rect 19100 -18572 19688 -18556
rect 20118 -18556 20134 -18539
rect 20690 -18539 20892 -18522
rect 20950 -18522 21910 -18484
rect 20950 -18539 21152 -18522
rect 20690 -18556 20706 -18539
rect 20118 -18572 20706 -18556
rect 21136 -18556 21152 -18539
rect 21708 -18539 21910 -18522
rect 21968 -18522 22928 -18484
rect 21968 -18539 22170 -18522
rect 21708 -18556 21724 -18539
rect 21136 -18572 21724 -18556
rect 22154 -18556 22170 -18539
rect 22726 -18539 22928 -18522
rect 22726 -18556 22742 -18539
rect 22154 -18572 22742 -18556
rect -9138 -18876 -8178 -18838
rect -9138 -18893 -8936 -18876
rect -8952 -18910 -8936 -18893
rect -8380 -18893 -8178 -18876
rect -8120 -18876 -7160 -18838
rect -8120 -18893 -7918 -18876
rect -8380 -18910 -8364 -18893
rect -8952 -18926 -8364 -18910
rect -7934 -18910 -7918 -18893
rect -7362 -18893 -7160 -18876
rect -7102 -18876 -6142 -18838
rect -7102 -18893 -6900 -18876
rect -7362 -18910 -7346 -18893
rect -7934 -18926 -7346 -18910
rect -6916 -18910 -6900 -18893
rect -6344 -18893 -6142 -18876
rect -6084 -18876 -5124 -18838
rect -6084 -18893 -5882 -18876
rect -6344 -18910 -6328 -18893
rect -6916 -18926 -6328 -18910
rect -5898 -18910 -5882 -18893
rect -5326 -18893 -5124 -18876
rect -5066 -18876 -4106 -18838
rect -5066 -18893 -4864 -18876
rect -5326 -18910 -5310 -18893
rect -5898 -18926 -5310 -18910
rect -4880 -18910 -4864 -18893
rect -4308 -18893 -4106 -18876
rect -4048 -18876 -3088 -18838
rect -4048 -18893 -3846 -18876
rect -4308 -18910 -4292 -18893
rect -4880 -18926 -4292 -18910
rect -3862 -18910 -3846 -18893
rect -3290 -18893 -3088 -18876
rect -3030 -18876 -2070 -18838
rect -3030 -18893 -2828 -18876
rect -3290 -18910 -3274 -18893
rect -3862 -18926 -3274 -18910
rect -2844 -18910 -2828 -18893
rect -2272 -18893 -2070 -18876
rect -2012 -18876 -1052 -18838
rect -2012 -18893 -1810 -18876
rect -2272 -18910 -2256 -18893
rect -2844 -18926 -2256 -18910
rect -1826 -18910 -1810 -18893
rect -1254 -18893 -1052 -18876
rect -994 -18876 -34 -18838
rect -994 -18893 -792 -18876
rect -1254 -18910 -1238 -18893
rect -1826 -18926 -1238 -18910
rect -808 -18910 -792 -18893
rect -236 -18893 -34 -18876
rect -236 -18910 -220 -18893
rect -808 -18926 -220 -18910
rect 2812 -19046 3400 -19030
rect 2812 -19063 2828 -19046
rect 2626 -19080 2828 -19063
rect 3384 -19063 3400 -19046
rect 3830 -19046 4418 -19030
rect 3830 -19063 3846 -19046
rect 3384 -19080 3586 -19063
rect 2626 -19118 3586 -19080
rect 3644 -19080 3846 -19063
rect 4402 -19063 4418 -19046
rect 4848 -19046 5436 -19030
rect 4848 -19063 4864 -19046
rect 4402 -19080 4604 -19063
rect 3644 -19118 4604 -19080
rect 4662 -19080 4864 -19063
rect 5420 -19063 5436 -19046
rect 5866 -19046 6454 -19030
rect 5866 -19063 5882 -19046
rect 5420 -19080 5622 -19063
rect 4662 -19118 5622 -19080
rect 5680 -19080 5882 -19063
rect 6438 -19063 6454 -19046
rect 6884 -19046 7472 -19030
rect 6884 -19063 6900 -19046
rect 6438 -19080 6640 -19063
rect 5680 -19118 6640 -19080
rect 6698 -19080 6900 -19063
rect 7456 -19063 7472 -19046
rect 7902 -19046 8490 -19030
rect 7902 -19063 7918 -19046
rect 7456 -19080 7658 -19063
rect 6698 -19118 7658 -19080
rect 7716 -19080 7918 -19063
rect 8474 -19063 8490 -19046
rect 8920 -19046 9508 -19030
rect 8920 -19063 8936 -19046
rect 8474 -19080 8676 -19063
rect 7716 -19118 8676 -19080
rect 8734 -19080 8936 -19063
rect 9492 -19063 9508 -19046
rect 9938 -19046 10526 -19030
rect 9938 -19063 9954 -19046
rect 9492 -19080 9694 -19063
rect 8734 -19118 9694 -19080
rect 9752 -19080 9954 -19063
rect 10510 -19063 10526 -19046
rect 10956 -19046 11544 -19030
rect 10956 -19063 10972 -19046
rect 10510 -19080 10712 -19063
rect 9752 -19118 10712 -19080
rect 10770 -19080 10972 -19063
rect 11528 -19063 11544 -19046
rect 11974 -19046 12562 -19030
rect 11974 -19063 11990 -19046
rect 11528 -19080 11730 -19063
rect 10770 -19118 11730 -19080
rect 11788 -19080 11990 -19063
rect 12546 -19063 12562 -19046
rect 12992 -19046 13580 -19030
rect 12992 -19063 13008 -19046
rect 12546 -19080 12748 -19063
rect 11788 -19118 12748 -19080
rect 12806 -19080 13008 -19063
rect 13564 -19063 13580 -19046
rect 14010 -19046 14598 -19030
rect 14010 -19063 14026 -19046
rect 13564 -19080 13766 -19063
rect 12806 -19118 13766 -19080
rect 13824 -19080 14026 -19063
rect 14582 -19063 14598 -19046
rect 15028 -19046 15616 -19030
rect 15028 -19063 15044 -19046
rect 14582 -19080 14784 -19063
rect 13824 -19118 14784 -19080
rect 14842 -19080 15044 -19063
rect 15600 -19063 15616 -19046
rect 16046 -19046 16634 -19030
rect 16046 -19063 16062 -19046
rect 15600 -19080 15802 -19063
rect 14842 -19118 15802 -19080
rect 15860 -19080 16062 -19063
rect 16618 -19063 16634 -19046
rect 17064 -19046 17652 -19030
rect 17064 -19063 17080 -19046
rect 16618 -19080 16820 -19063
rect 15860 -19118 16820 -19080
rect 16878 -19080 17080 -19063
rect 17636 -19063 17652 -19046
rect 18082 -19046 18670 -19030
rect 18082 -19063 18098 -19046
rect 17636 -19080 17838 -19063
rect 16878 -19118 17838 -19080
rect 17896 -19080 18098 -19063
rect 18654 -19063 18670 -19046
rect 19100 -19046 19688 -19030
rect 19100 -19063 19116 -19046
rect 18654 -19080 18856 -19063
rect 17896 -19118 18856 -19080
rect 18914 -19080 19116 -19063
rect 19672 -19063 19688 -19046
rect 20118 -19046 20706 -19030
rect 20118 -19063 20134 -19046
rect 19672 -19080 19874 -19063
rect 18914 -19118 19874 -19080
rect 19932 -19080 20134 -19063
rect 20690 -19063 20706 -19046
rect 21136 -19046 21724 -19030
rect 21136 -19063 21152 -19046
rect 20690 -19080 20892 -19063
rect 19932 -19118 20892 -19080
rect 20950 -19080 21152 -19063
rect 21708 -19063 21724 -19046
rect 22154 -19046 22742 -19030
rect 22154 -19063 22170 -19046
rect 21708 -19080 21910 -19063
rect 20950 -19118 21910 -19080
rect 21968 -19080 22170 -19063
rect 22726 -19063 22742 -19046
rect 22726 -19080 22928 -19063
rect 21968 -19118 22928 -19080
rect -2252 -19550 -2144 -19534
rect -2252 -19567 -2236 -19550
rect -2278 -19584 -2236 -19567
rect -2160 -19567 -2144 -19550
rect -2034 -19550 -1926 -19534
rect -2034 -19567 -2018 -19550
rect -2160 -19584 -2118 -19567
rect -2278 -19622 -2118 -19584
rect -2060 -19584 -2018 -19567
rect -1942 -19567 -1926 -19550
rect -1816 -19550 -1708 -19534
rect -1816 -19567 -1800 -19550
rect -1942 -19584 -1900 -19567
rect -2060 -19622 -1900 -19584
rect -1842 -19584 -1800 -19567
rect -1724 -19567 -1708 -19550
rect -1598 -19550 -1490 -19534
rect -1598 -19567 -1582 -19550
rect -1724 -19584 -1682 -19567
rect -1842 -19622 -1682 -19584
rect -1624 -19584 -1582 -19567
rect -1506 -19567 -1490 -19550
rect -1380 -19550 -1272 -19534
rect -1380 -19567 -1364 -19550
rect -1506 -19584 -1464 -19567
rect -1624 -19622 -1464 -19584
rect -1406 -19584 -1364 -19567
rect -1288 -19567 -1272 -19550
rect -1162 -19550 -1054 -19534
rect -1162 -19567 -1146 -19550
rect -1288 -19584 -1246 -19567
rect -1406 -19622 -1246 -19584
rect -1188 -19584 -1146 -19567
rect -1070 -19567 -1054 -19550
rect -944 -19550 -836 -19534
rect -944 -19567 -928 -19550
rect -1070 -19584 -1028 -19567
rect -1188 -19622 -1028 -19584
rect -970 -19584 -928 -19567
rect -852 -19567 -836 -19550
rect -726 -19550 -618 -19534
rect -726 -19567 -710 -19550
rect -852 -19584 -810 -19567
rect -970 -19622 -810 -19584
rect -752 -19584 -710 -19567
rect -634 -19567 -618 -19550
rect -508 -19550 -400 -19534
rect -508 -19567 -492 -19550
rect -634 -19584 -592 -19567
rect -752 -19622 -592 -19584
rect -534 -19584 -492 -19567
rect -416 -19567 -400 -19550
rect -290 -19550 -182 -19534
rect -290 -19567 -274 -19550
rect -416 -19584 -374 -19567
rect -534 -19622 -374 -19584
rect -316 -19584 -274 -19567
rect -198 -19567 -182 -19550
rect -198 -19584 -156 -19567
rect -316 -19622 -156 -19584
rect 2626 -19756 3586 -19718
rect 2626 -19773 2828 -19756
rect 2812 -19790 2828 -19773
rect 3384 -19773 3586 -19756
rect 3644 -19756 4604 -19718
rect 3644 -19773 3846 -19756
rect 3384 -19790 3400 -19773
rect 2812 -19806 3400 -19790
rect 3830 -19790 3846 -19773
rect 4402 -19773 4604 -19756
rect 4662 -19756 5622 -19718
rect 4662 -19773 4864 -19756
rect 4402 -19790 4418 -19773
rect 3830 -19806 4418 -19790
rect 4848 -19790 4864 -19773
rect 5420 -19773 5622 -19756
rect 5680 -19756 6640 -19718
rect 5680 -19773 5882 -19756
rect 5420 -19790 5436 -19773
rect 4848 -19806 5436 -19790
rect 5866 -19790 5882 -19773
rect 6438 -19773 6640 -19756
rect 6698 -19756 7658 -19718
rect 6698 -19773 6900 -19756
rect 6438 -19790 6454 -19773
rect 5866 -19806 6454 -19790
rect 6884 -19790 6900 -19773
rect 7456 -19773 7658 -19756
rect 7716 -19756 8676 -19718
rect 7716 -19773 7918 -19756
rect 7456 -19790 7472 -19773
rect 6884 -19806 7472 -19790
rect 7902 -19790 7918 -19773
rect 8474 -19773 8676 -19756
rect 8734 -19756 9694 -19718
rect 8734 -19773 8936 -19756
rect 8474 -19790 8490 -19773
rect 7902 -19806 8490 -19790
rect 8920 -19790 8936 -19773
rect 9492 -19773 9694 -19756
rect 9752 -19756 10712 -19718
rect 9752 -19773 9954 -19756
rect 9492 -19790 9508 -19773
rect 8920 -19806 9508 -19790
rect 9938 -19790 9954 -19773
rect 10510 -19773 10712 -19756
rect 10770 -19756 11730 -19718
rect 10770 -19773 10972 -19756
rect 10510 -19790 10526 -19773
rect 9938 -19806 10526 -19790
rect 10956 -19790 10972 -19773
rect 11528 -19773 11730 -19756
rect 11788 -19756 12748 -19718
rect 11788 -19773 11990 -19756
rect 11528 -19790 11544 -19773
rect 10956 -19806 11544 -19790
rect 11974 -19790 11990 -19773
rect 12546 -19773 12748 -19756
rect 12806 -19756 13766 -19718
rect 12806 -19773 13008 -19756
rect 12546 -19790 12562 -19773
rect 11974 -19806 12562 -19790
rect 12992 -19790 13008 -19773
rect 13564 -19773 13766 -19756
rect 13824 -19756 14784 -19718
rect 13824 -19773 14026 -19756
rect 13564 -19790 13580 -19773
rect 12992 -19806 13580 -19790
rect 14010 -19790 14026 -19773
rect 14582 -19773 14784 -19756
rect 14842 -19756 15802 -19718
rect 14842 -19773 15044 -19756
rect 14582 -19790 14598 -19773
rect 14010 -19806 14598 -19790
rect 15028 -19790 15044 -19773
rect 15600 -19773 15802 -19756
rect 15860 -19756 16820 -19718
rect 15860 -19773 16062 -19756
rect 15600 -19790 15616 -19773
rect 15028 -19806 15616 -19790
rect 16046 -19790 16062 -19773
rect 16618 -19773 16820 -19756
rect 16878 -19756 17838 -19718
rect 16878 -19773 17080 -19756
rect 16618 -19790 16634 -19773
rect 16046 -19806 16634 -19790
rect 17064 -19790 17080 -19773
rect 17636 -19773 17838 -19756
rect 17896 -19756 18856 -19718
rect 17896 -19773 18098 -19756
rect 17636 -19790 17652 -19773
rect 17064 -19806 17652 -19790
rect 18082 -19790 18098 -19773
rect 18654 -19773 18856 -19756
rect 18914 -19756 19874 -19718
rect 18914 -19773 19116 -19756
rect 18654 -19790 18670 -19773
rect 18082 -19806 18670 -19790
rect 19100 -19790 19116 -19773
rect 19672 -19773 19874 -19756
rect 19932 -19756 20892 -19718
rect 19932 -19773 20134 -19756
rect 19672 -19790 19688 -19773
rect 19100 -19806 19688 -19790
rect 20118 -19790 20134 -19773
rect 20690 -19773 20892 -19756
rect 20950 -19756 21910 -19718
rect 20950 -19773 21152 -19756
rect 20690 -19790 20706 -19773
rect 20118 -19806 20706 -19790
rect 21136 -19790 21152 -19773
rect 21708 -19773 21910 -19756
rect 21968 -19756 22928 -19718
rect 21968 -19773 22170 -19756
rect 21708 -19790 21724 -19773
rect 21136 -19806 21724 -19790
rect 22154 -19790 22170 -19773
rect 22726 -19773 22928 -19756
rect 22726 -19790 22742 -19773
rect 22154 -19806 22742 -19790
rect -2278 -19860 -2118 -19822
rect -2278 -19877 -2236 -19860
rect -2252 -19894 -2236 -19877
rect -2160 -19877 -2118 -19860
rect -2060 -19860 -1900 -19822
rect -2060 -19877 -2018 -19860
rect -2160 -19894 -2144 -19877
rect -2252 -19910 -2144 -19894
rect -2034 -19894 -2018 -19877
rect -1942 -19877 -1900 -19860
rect -1842 -19860 -1682 -19822
rect -1842 -19877 -1800 -19860
rect -1942 -19894 -1926 -19877
rect -2034 -19910 -1926 -19894
rect -1816 -19894 -1800 -19877
rect -1724 -19877 -1682 -19860
rect -1624 -19860 -1464 -19822
rect -1624 -19877 -1582 -19860
rect -1724 -19894 -1708 -19877
rect -1816 -19910 -1708 -19894
rect -1598 -19894 -1582 -19877
rect -1506 -19877 -1464 -19860
rect -1406 -19860 -1246 -19822
rect -1406 -19877 -1364 -19860
rect -1506 -19894 -1490 -19877
rect -1598 -19910 -1490 -19894
rect -1380 -19894 -1364 -19877
rect -1288 -19877 -1246 -19860
rect -1188 -19860 -1028 -19822
rect -1188 -19877 -1146 -19860
rect -1288 -19894 -1272 -19877
rect -1380 -19910 -1272 -19894
rect -1162 -19894 -1146 -19877
rect -1070 -19877 -1028 -19860
rect -970 -19860 -810 -19822
rect -970 -19877 -928 -19860
rect -1070 -19894 -1054 -19877
rect -1162 -19910 -1054 -19894
rect -944 -19894 -928 -19877
rect -852 -19877 -810 -19860
rect -752 -19860 -592 -19822
rect -752 -19877 -710 -19860
rect -852 -19894 -836 -19877
rect -944 -19910 -836 -19894
rect -726 -19894 -710 -19877
rect -634 -19877 -592 -19860
rect -534 -19860 -374 -19822
rect -534 -19877 -492 -19860
rect -634 -19894 -618 -19877
rect -726 -19910 -618 -19894
rect -508 -19894 -492 -19877
rect -416 -19877 -374 -19860
rect -316 -19860 -156 -19822
rect -316 -19877 -274 -19860
rect -416 -19894 -400 -19877
rect -508 -19910 -400 -19894
rect -290 -19894 -274 -19877
rect -198 -19877 -156 -19860
rect -198 -19894 -182 -19877
rect -290 -19910 -182 -19894
rect 2812 -20280 3400 -20264
rect 2812 -20297 2828 -20280
rect 2626 -20314 2828 -20297
rect 3384 -20297 3400 -20280
rect 3830 -20280 4418 -20264
rect 3830 -20297 3846 -20280
rect 3384 -20314 3586 -20297
rect 2626 -20352 3586 -20314
rect 3644 -20314 3846 -20297
rect 4402 -20297 4418 -20280
rect 4848 -20280 5436 -20264
rect 4848 -20297 4864 -20280
rect 4402 -20314 4604 -20297
rect 3644 -20352 4604 -20314
rect 4662 -20314 4864 -20297
rect 5420 -20297 5436 -20280
rect 5866 -20280 6454 -20264
rect 5866 -20297 5882 -20280
rect 5420 -20314 5622 -20297
rect 4662 -20352 5622 -20314
rect 5680 -20314 5882 -20297
rect 6438 -20297 6454 -20280
rect 6884 -20280 7472 -20264
rect 6884 -20297 6900 -20280
rect 6438 -20314 6640 -20297
rect 5680 -20352 6640 -20314
rect 6698 -20314 6900 -20297
rect 7456 -20297 7472 -20280
rect 7902 -20280 8490 -20264
rect 7902 -20297 7918 -20280
rect 7456 -20314 7658 -20297
rect 6698 -20352 7658 -20314
rect 7716 -20314 7918 -20297
rect 8474 -20297 8490 -20280
rect 8920 -20280 9508 -20264
rect 8920 -20297 8936 -20280
rect 8474 -20314 8676 -20297
rect 7716 -20352 8676 -20314
rect 8734 -20314 8936 -20297
rect 9492 -20297 9508 -20280
rect 9938 -20280 10526 -20264
rect 9938 -20297 9954 -20280
rect 9492 -20314 9694 -20297
rect 8734 -20352 9694 -20314
rect 9752 -20314 9954 -20297
rect 10510 -20297 10526 -20280
rect 10956 -20280 11544 -20264
rect 10956 -20297 10972 -20280
rect 10510 -20314 10712 -20297
rect 9752 -20352 10712 -20314
rect 10770 -20314 10972 -20297
rect 11528 -20297 11544 -20280
rect 11974 -20280 12562 -20264
rect 11974 -20297 11990 -20280
rect 11528 -20314 11730 -20297
rect 10770 -20352 11730 -20314
rect 11788 -20314 11990 -20297
rect 12546 -20297 12562 -20280
rect 12992 -20280 13580 -20264
rect 12992 -20297 13008 -20280
rect 12546 -20314 12748 -20297
rect 11788 -20352 12748 -20314
rect 12806 -20314 13008 -20297
rect 13564 -20297 13580 -20280
rect 14010 -20280 14598 -20264
rect 14010 -20297 14026 -20280
rect 13564 -20314 13766 -20297
rect 12806 -20352 13766 -20314
rect 13824 -20314 14026 -20297
rect 14582 -20297 14598 -20280
rect 15028 -20280 15616 -20264
rect 15028 -20297 15044 -20280
rect 14582 -20314 14784 -20297
rect 13824 -20352 14784 -20314
rect 14842 -20314 15044 -20297
rect 15600 -20297 15616 -20280
rect 16046 -20280 16634 -20264
rect 16046 -20297 16062 -20280
rect 15600 -20314 15802 -20297
rect 14842 -20352 15802 -20314
rect 15860 -20314 16062 -20297
rect 16618 -20297 16634 -20280
rect 17064 -20280 17652 -20264
rect 17064 -20297 17080 -20280
rect 16618 -20314 16820 -20297
rect 15860 -20352 16820 -20314
rect 16878 -20314 17080 -20297
rect 17636 -20297 17652 -20280
rect 18082 -20280 18670 -20264
rect 18082 -20297 18098 -20280
rect 17636 -20314 17838 -20297
rect 16878 -20352 17838 -20314
rect 17896 -20314 18098 -20297
rect 18654 -20297 18670 -20280
rect 19100 -20280 19688 -20264
rect 19100 -20297 19116 -20280
rect 18654 -20314 18856 -20297
rect 17896 -20352 18856 -20314
rect 18914 -20314 19116 -20297
rect 19672 -20297 19688 -20280
rect 20118 -20280 20706 -20264
rect 20118 -20297 20134 -20280
rect 19672 -20314 19874 -20297
rect 18914 -20352 19874 -20314
rect 19932 -20314 20134 -20297
rect 20690 -20297 20706 -20280
rect 21136 -20280 21724 -20264
rect 21136 -20297 21152 -20280
rect 20690 -20314 20892 -20297
rect 19932 -20352 20892 -20314
rect 20950 -20314 21152 -20297
rect 21708 -20297 21724 -20280
rect 22154 -20280 22742 -20264
rect 22154 -20297 22170 -20280
rect 21708 -20314 21910 -20297
rect 20950 -20352 21910 -20314
rect 21968 -20314 22170 -20297
rect 22726 -20297 22742 -20280
rect 22726 -20314 22928 -20297
rect 21968 -20352 22928 -20314
rect -2252 -20382 -2144 -20366
rect -2252 -20399 -2236 -20382
rect -2278 -20416 -2236 -20399
rect -2160 -20399 -2144 -20382
rect -2034 -20382 -1926 -20366
rect -2034 -20399 -2018 -20382
rect -2160 -20416 -2118 -20399
rect -2278 -20454 -2118 -20416
rect -2060 -20416 -2018 -20399
rect -1942 -20399 -1926 -20382
rect -1816 -20382 -1708 -20366
rect -1816 -20399 -1800 -20382
rect -1942 -20416 -1900 -20399
rect -2060 -20454 -1900 -20416
rect -1842 -20416 -1800 -20399
rect -1724 -20399 -1708 -20382
rect -1598 -20382 -1490 -20366
rect -1598 -20399 -1582 -20382
rect -1724 -20416 -1682 -20399
rect -1842 -20454 -1682 -20416
rect -1624 -20416 -1582 -20399
rect -1506 -20399 -1490 -20382
rect -1380 -20382 -1272 -20366
rect -1380 -20399 -1364 -20382
rect -1506 -20416 -1464 -20399
rect -1624 -20454 -1464 -20416
rect -1406 -20416 -1364 -20399
rect -1288 -20399 -1272 -20382
rect -1162 -20382 -1054 -20366
rect -1162 -20399 -1146 -20382
rect -1288 -20416 -1246 -20399
rect -1406 -20454 -1246 -20416
rect -1188 -20416 -1146 -20399
rect -1070 -20399 -1054 -20382
rect -944 -20382 -836 -20366
rect -944 -20399 -928 -20382
rect -1070 -20416 -1028 -20399
rect -1188 -20454 -1028 -20416
rect -970 -20416 -928 -20399
rect -852 -20399 -836 -20382
rect -726 -20382 -618 -20366
rect -726 -20399 -710 -20382
rect -852 -20416 -810 -20399
rect -970 -20454 -810 -20416
rect -752 -20416 -710 -20399
rect -634 -20399 -618 -20382
rect -508 -20382 -400 -20366
rect -508 -20399 -492 -20382
rect -634 -20416 -592 -20399
rect -752 -20454 -592 -20416
rect -534 -20416 -492 -20399
rect -416 -20399 -400 -20382
rect -290 -20382 -182 -20366
rect -290 -20399 -274 -20382
rect -416 -20416 -374 -20399
rect -534 -20454 -374 -20416
rect -316 -20416 -274 -20399
rect -198 -20399 -182 -20382
rect -198 -20416 -156 -20399
rect -316 -20454 -156 -20416
rect -2278 -20692 -2118 -20654
rect -2278 -20709 -2236 -20692
rect -2252 -20726 -2236 -20709
rect -2160 -20709 -2118 -20692
rect -2060 -20692 -1900 -20654
rect -2060 -20709 -2018 -20692
rect -2160 -20726 -2144 -20709
rect -2252 -20742 -2144 -20726
rect -2034 -20726 -2018 -20709
rect -1942 -20709 -1900 -20692
rect -1842 -20692 -1682 -20654
rect -1842 -20709 -1800 -20692
rect -1942 -20726 -1926 -20709
rect -2034 -20742 -1926 -20726
rect -1816 -20726 -1800 -20709
rect -1724 -20709 -1682 -20692
rect -1624 -20692 -1464 -20654
rect -1624 -20709 -1582 -20692
rect -1724 -20726 -1708 -20709
rect -1816 -20742 -1708 -20726
rect -1598 -20726 -1582 -20709
rect -1506 -20709 -1464 -20692
rect -1406 -20692 -1246 -20654
rect -1406 -20709 -1364 -20692
rect -1506 -20726 -1490 -20709
rect -1598 -20742 -1490 -20726
rect -1380 -20726 -1364 -20709
rect -1288 -20709 -1246 -20692
rect -1188 -20692 -1028 -20654
rect -1188 -20709 -1146 -20692
rect -1288 -20726 -1272 -20709
rect -1380 -20742 -1272 -20726
rect -1162 -20726 -1146 -20709
rect -1070 -20709 -1028 -20692
rect -970 -20692 -810 -20654
rect -970 -20709 -928 -20692
rect -1070 -20726 -1054 -20709
rect -1162 -20742 -1054 -20726
rect -944 -20726 -928 -20709
rect -852 -20709 -810 -20692
rect -752 -20692 -592 -20654
rect -752 -20709 -710 -20692
rect -852 -20726 -836 -20709
rect -944 -20742 -836 -20726
rect -726 -20726 -710 -20709
rect -634 -20709 -592 -20692
rect -534 -20692 -374 -20654
rect -534 -20709 -492 -20692
rect -634 -20726 -618 -20709
rect -726 -20742 -618 -20726
rect -508 -20726 -492 -20709
rect -416 -20709 -374 -20692
rect -316 -20692 -156 -20654
rect -316 -20709 -274 -20692
rect -416 -20726 -400 -20709
rect -508 -20742 -400 -20726
rect -290 -20726 -274 -20709
rect -198 -20709 -156 -20692
rect -198 -20726 -182 -20709
rect -290 -20742 -182 -20726
rect 2626 -20990 3586 -20952
rect 2626 -21007 2828 -20990
rect 2812 -21024 2828 -21007
rect 3384 -21007 3586 -20990
rect 3644 -20990 4604 -20952
rect 3644 -21007 3846 -20990
rect 3384 -21024 3400 -21007
rect 2812 -21040 3400 -21024
rect 3830 -21024 3846 -21007
rect 4402 -21007 4604 -20990
rect 4662 -20990 5622 -20952
rect 4662 -21007 4864 -20990
rect 4402 -21024 4418 -21007
rect 3830 -21040 4418 -21024
rect 4848 -21024 4864 -21007
rect 5420 -21007 5622 -20990
rect 5680 -20990 6640 -20952
rect 5680 -21007 5882 -20990
rect 5420 -21024 5436 -21007
rect 4848 -21040 5436 -21024
rect 5866 -21024 5882 -21007
rect 6438 -21007 6640 -20990
rect 6698 -20990 7658 -20952
rect 6698 -21007 6900 -20990
rect 6438 -21024 6454 -21007
rect 5866 -21040 6454 -21024
rect 6884 -21024 6900 -21007
rect 7456 -21007 7658 -20990
rect 7716 -20990 8676 -20952
rect 7716 -21007 7918 -20990
rect 7456 -21024 7472 -21007
rect 6884 -21040 7472 -21024
rect 7902 -21024 7918 -21007
rect 8474 -21007 8676 -20990
rect 8734 -20990 9694 -20952
rect 8734 -21007 8936 -20990
rect 8474 -21024 8490 -21007
rect 7902 -21040 8490 -21024
rect 8920 -21024 8936 -21007
rect 9492 -21007 9694 -20990
rect 9752 -20990 10712 -20952
rect 9752 -21007 9954 -20990
rect 9492 -21024 9508 -21007
rect 8920 -21040 9508 -21024
rect 9938 -21024 9954 -21007
rect 10510 -21007 10712 -20990
rect 10770 -20990 11730 -20952
rect 10770 -21007 10972 -20990
rect 10510 -21024 10526 -21007
rect 9938 -21040 10526 -21024
rect 10956 -21024 10972 -21007
rect 11528 -21007 11730 -20990
rect 11788 -20990 12748 -20952
rect 11788 -21007 11990 -20990
rect 11528 -21024 11544 -21007
rect 10956 -21040 11544 -21024
rect 11974 -21024 11990 -21007
rect 12546 -21007 12748 -20990
rect 12806 -20990 13766 -20952
rect 12806 -21007 13008 -20990
rect 12546 -21024 12562 -21007
rect 11974 -21040 12562 -21024
rect 12992 -21024 13008 -21007
rect 13564 -21007 13766 -20990
rect 13824 -20990 14784 -20952
rect 13824 -21007 14026 -20990
rect 13564 -21024 13580 -21007
rect 12992 -21040 13580 -21024
rect 14010 -21024 14026 -21007
rect 14582 -21007 14784 -20990
rect 14842 -20990 15802 -20952
rect 14842 -21007 15044 -20990
rect 14582 -21024 14598 -21007
rect 14010 -21040 14598 -21024
rect 15028 -21024 15044 -21007
rect 15600 -21007 15802 -20990
rect 15860 -20990 16820 -20952
rect 15860 -21007 16062 -20990
rect 15600 -21024 15616 -21007
rect 15028 -21040 15616 -21024
rect 16046 -21024 16062 -21007
rect 16618 -21007 16820 -20990
rect 16878 -20990 17838 -20952
rect 16878 -21007 17080 -20990
rect 16618 -21024 16634 -21007
rect 16046 -21040 16634 -21024
rect 17064 -21024 17080 -21007
rect 17636 -21007 17838 -20990
rect 17896 -20990 18856 -20952
rect 17896 -21007 18098 -20990
rect 17636 -21024 17652 -21007
rect 17064 -21040 17652 -21024
rect 18082 -21024 18098 -21007
rect 18654 -21007 18856 -20990
rect 18914 -20990 19874 -20952
rect 18914 -21007 19116 -20990
rect 18654 -21024 18670 -21007
rect 18082 -21040 18670 -21024
rect 19100 -21024 19116 -21007
rect 19672 -21007 19874 -20990
rect 19932 -20990 20892 -20952
rect 19932 -21007 20134 -20990
rect 19672 -21024 19688 -21007
rect 19100 -21040 19688 -21024
rect 20118 -21024 20134 -21007
rect 20690 -21007 20892 -20990
rect 20950 -20990 21910 -20952
rect 20950 -21007 21152 -20990
rect 20690 -21024 20706 -21007
rect 20118 -21040 20706 -21024
rect 21136 -21024 21152 -21007
rect 21708 -21007 21910 -20990
rect 21968 -20990 22928 -20952
rect 21968 -21007 22170 -20990
rect 21708 -21024 21724 -21007
rect 21136 -21040 21724 -21024
rect 22154 -21024 22170 -21007
rect 22726 -21007 22928 -20990
rect 22726 -21024 22742 -21007
rect 22154 -21040 22742 -21024
rect 2812 -21512 3400 -21496
rect 2812 -21529 2828 -21512
rect 2626 -21546 2828 -21529
rect 3384 -21529 3400 -21512
rect 3830 -21512 4418 -21496
rect 3830 -21529 3846 -21512
rect 3384 -21546 3586 -21529
rect 2626 -21584 3586 -21546
rect 3644 -21546 3846 -21529
rect 4402 -21529 4418 -21512
rect 4848 -21512 5436 -21496
rect 4848 -21529 4864 -21512
rect 4402 -21546 4604 -21529
rect 3644 -21584 4604 -21546
rect 4662 -21546 4864 -21529
rect 5420 -21529 5436 -21512
rect 5866 -21512 6454 -21496
rect 5866 -21529 5882 -21512
rect 5420 -21546 5622 -21529
rect 4662 -21584 5622 -21546
rect 5680 -21546 5882 -21529
rect 6438 -21529 6454 -21512
rect 6884 -21512 7472 -21496
rect 6884 -21529 6900 -21512
rect 6438 -21546 6640 -21529
rect 5680 -21584 6640 -21546
rect 6698 -21546 6900 -21529
rect 7456 -21529 7472 -21512
rect 7902 -21512 8490 -21496
rect 7902 -21529 7918 -21512
rect 7456 -21546 7658 -21529
rect 6698 -21584 7658 -21546
rect 7716 -21546 7918 -21529
rect 8474 -21529 8490 -21512
rect 8920 -21512 9508 -21496
rect 8920 -21529 8936 -21512
rect 8474 -21546 8676 -21529
rect 7716 -21584 8676 -21546
rect 8734 -21546 8936 -21529
rect 9492 -21529 9508 -21512
rect 9938 -21512 10526 -21496
rect 9938 -21529 9954 -21512
rect 9492 -21546 9694 -21529
rect 8734 -21584 9694 -21546
rect 9752 -21546 9954 -21529
rect 10510 -21529 10526 -21512
rect 10956 -21512 11544 -21496
rect 10956 -21529 10972 -21512
rect 10510 -21546 10712 -21529
rect 9752 -21584 10712 -21546
rect 10770 -21546 10972 -21529
rect 11528 -21529 11544 -21512
rect 11974 -21512 12562 -21496
rect 11974 -21529 11990 -21512
rect 11528 -21546 11730 -21529
rect 10770 -21584 11730 -21546
rect 11788 -21546 11990 -21529
rect 12546 -21529 12562 -21512
rect 12992 -21512 13580 -21496
rect 12992 -21529 13008 -21512
rect 12546 -21546 12748 -21529
rect 11788 -21584 12748 -21546
rect 12806 -21546 13008 -21529
rect 13564 -21529 13580 -21512
rect 14010 -21512 14598 -21496
rect 14010 -21529 14026 -21512
rect 13564 -21546 13766 -21529
rect 12806 -21584 13766 -21546
rect 13824 -21546 14026 -21529
rect 14582 -21529 14598 -21512
rect 15028 -21512 15616 -21496
rect 15028 -21529 15044 -21512
rect 14582 -21546 14784 -21529
rect 13824 -21584 14784 -21546
rect 14842 -21546 15044 -21529
rect 15600 -21529 15616 -21512
rect 16046 -21512 16634 -21496
rect 16046 -21529 16062 -21512
rect 15600 -21546 15802 -21529
rect 14842 -21584 15802 -21546
rect 15860 -21546 16062 -21529
rect 16618 -21529 16634 -21512
rect 17064 -21512 17652 -21496
rect 17064 -21529 17080 -21512
rect 16618 -21546 16820 -21529
rect 15860 -21584 16820 -21546
rect 16878 -21546 17080 -21529
rect 17636 -21529 17652 -21512
rect 18082 -21512 18670 -21496
rect 18082 -21529 18098 -21512
rect 17636 -21546 17838 -21529
rect 16878 -21584 17838 -21546
rect 17896 -21546 18098 -21529
rect 18654 -21529 18670 -21512
rect 19100 -21512 19688 -21496
rect 19100 -21529 19116 -21512
rect 18654 -21546 18856 -21529
rect 17896 -21584 18856 -21546
rect 18914 -21546 19116 -21529
rect 19672 -21529 19688 -21512
rect 20118 -21512 20706 -21496
rect 20118 -21529 20134 -21512
rect 19672 -21546 19874 -21529
rect 18914 -21584 19874 -21546
rect 19932 -21546 20134 -21529
rect 20690 -21529 20706 -21512
rect 21136 -21512 21724 -21496
rect 21136 -21529 21152 -21512
rect 20690 -21546 20892 -21529
rect 19932 -21584 20892 -21546
rect 20950 -21546 21152 -21529
rect 21708 -21529 21724 -21512
rect 22154 -21512 22742 -21496
rect 22154 -21529 22170 -21512
rect 21708 -21546 21910 -21529
rect 20950 -21584 21910 -21546
rect 21968 -21546 22170 -21529
rect 22726 -21529 22742 -21512
rect 22726 -21546 22928 -21529
rect 21968 -21584 22928 -21546
rect -9173 -21709 -8585 -21693
rect -9173 -21726 -9157 -21709
rect -9359 -21743 -9157 -21726
rect -8601 -21726 -8585 -21709
rect -8155 -21709 -7567 -21693
rect -8155 -21726 -8139 -21709
rect -8601 -21743 -8399 -21726
rect -9359 -21781 -8399 -21743
rect -8341 -21743 -8139 -21726
rect -7583 -21726 -7567 -21709
rect -7137 -21709 -6549 -21693
rect -7137 -21726 -7121 -21709
rect -7583 -21743 -7381 -21726
rect -8341 -21781 -7381 -21743
rect -7323 -21743 -7121 -21726
rect -6565 -21726 -6549 -21709
rect -6119 -21709 -5531 -21693
rect -6119 -21726 -6103 -21709
rect -6565 -21743 -6363 -21726
rect -7323 -21781 -6363 -21743
rect -6305 -21743 -6103 -21726
rect -5547 -21726 -5531 -21709
rect -5101 -21709 -4513 -21693
rect -5101 -21726 -5085 -21709
rect -5547 -21743 -5345 -21726
rect -6305 -21781 -5345 -21743
rect -5287 -21743 -5085 -21726
rect -4529 -21726 -4513 -21709
rect -4083 -21709 -3495 -21693
rect -4083 -21726 -4067 -21709
rect -4529 -21743 -4327 -21726
rect -5287 -21781 -4327 -21743
rect -4269 -21743 -4067 -21726
rect -3511 -21726 -3495 -21709
rect -2322 -21708 -2166 -21692
rect -2322 -21725 -2306 -21708
rect -3511 -21743 -3309 -21726
rect -4269 -21781 -3309 -21743
rect -2364 -21742 -2306 -21725
rect -2182 -21725 -2166 -21708
rect -2024 -21708 -1868 -21692
rect -2024 -21725 -2008 -21708
rect -2182 -21742 -2124 -21725
rect -2364 -21780 -2124 -21742
rect -2066 -21742 -2008 -21725
rect -1884 -21725 -1868 -21708
rect -1726 -21708 -1570 -21692
rect -1726 -21725 -1710 -21708
rect -1884 -21742 -1826 -21725
rect -2066 -21780 -1826 -21742
rect -1768 -21742 -1710 -21725
rect -1586 -21725 -1570 -21708
rect -1428 -21708 -1272 -21692
rect -1428 -21725 -1412 -21708
rect -1586 -21742 -1528 -21725
rect -1768 -21780 -1528 -21742
rect -1470 -21742 -1412 -21725
rect -1288 -21725 -1272 -21708
rect -1130 -21708 -974 -21692
rect -1130 -21725 -1114 -21708
rect -1288 -21742 -1230 -21725
rect -1470 -21780 -1230 -21742
rect -1172 -21742 -1114 -21725
rect -990 -21725 -974 -21708
rect -832 -21708 -676 -21692
rect -832 -21725 -816 -21708
rect -990 -21742 -932 -21725
rect -1172 -21780 -932 -21742
rect -874 -21742 -816 -21725
rect -692 -21725 -676 -21708
rect -534 -21708 -378 -21692
rect -534 -21725 -518 -21708
rect -692 -21742 -634 -21725
rect -874 -21780 -634 -21742
rect -576 -21742 -518 -21725
rect -394 -21725 -378 -21708
rect -236 -21708 -80 -21692
rect -236 -21725 -220 -21708
rect -394 -21742 -336 -21725
rect -576 -21780 -336 -21742
rect -278 -21742 -220 -21725
rect -96 -21725 -80 -21708
rect 62 -21708 218 -21692
rect 62 -21725 78 -21708
rect -96 -21742 -38 -21725
rect -278 -21780 -38 -21742
rect 20 -21742 78 -21725
rect 202 -21725 218 -21708
rect 360 -21708 516 -21692
rect 360 -21725 376 -21708
rect 202 -21742 260 -21725
rect 20 -21780 260 -21742
rect 318 -21742 376 -21725
rect 500 -21725 516 -21708
rect 658 -21708 814 -21692
rect 658 -21725 674 -21708
rect 500 -21742 558 -21725
rect 318 -21780 558 -21742
rect 616 -21742 674 -21725
rect 798 -21725 814 -21708
rect 798 -21742 856 -21725
rect 616 -21780 856 -21742
rect 2626 -22222 3586 -22184
rect 2626 -22239 2828 -22222
rect 2812 -22256 2828 -22239
rect 3384 -22239 3586 -22222
rect 3644 -22222 4604 -22184
rect 3644 -22239 3846 -22222
rect 3384 -22256 3400 -22239
rect 2812 -22272 3400 -22256
rect 3830 -22256 3846 -22239
rect 4402 -22239 4604 -22222
rect 4662 -22222 5622 -22184
rect 4662 -22239 4864 -22222
rect 4402 -22256 4418 -22239
rect 3830 -22272 4418 -22256
rect 4848 -22256 4864 -22239
rect 5420 -22239 5622 -22222
rect 5680 -22222 6640 -22184
rect 5680 -22239 5882 -22222
rect 5420 -22256 5436 -22239
rect 4848 -22272 5436 -22256
rect 5866 -22256 5882 -22239
rect 6438 -22239 6640 -22222
rect 6698 -22222 7658 -22184
rect 6698 -22239 6900 -22222
rect 6438 -22256 6454 -22239
rect 5866 -22272 6454 -22256
rect 6884 -22256 6900 -22239
rect 7456 -22239 7658 -22222
rect 7716 -22222 8676 -22184
rect 7716 -22239 7918 -22222
rect 7456 -22256 7472 -22239
rect 6884 -22272 7472 -22256
rect 7902 -22256 7918 -22239
rect 8474 -22239 8676 -22222
rect 8734 -22222 9694 -22184
rect 8734 -22239 8936 -22222
rect 8474 -22256 8490 -22239
rect 7902 -22272 8490 -22256
rect 8920 -22256 8936 -22239
rect 9492 -22239 9694 -22222
rect 9752 -22222 10712 -22184
rect 9752 -22239 9954 -22222
rect 9492 -22256 9508 -22239
rect 8920 -22272 9508 -22256
rect 9938 -22256 9954 -22239
rect 10510 -22239 10712 -22222
rect 10770 -22222 11730 -22184
rect 10770 -22239 10972 -22222
rect 10510 -22256 10526 -22239
rect 9938 -22272 10526 -22256
rect 10956 -22256 10972 -22239
rect 11528 -22239 11730 -22222
rect 11788 -22222 12748 -22184
rect 11788 -22239 11990 -22222
rect 11528 -22256 11544 -22239
rect 10956 -22272 11544 -22256
rect 11974 -22256 11990 -22239
rect 12546 -22239 12748 -22222
rect 12806 -22222 13766 -22184
rect 12806 -22239 13008 -22222
rect 12546 -22256 12562 -22239
rect 11974 -22272 12562 -22256
rect 12992 -22256 13008 -22239
rect 13564 -22239 13766 -22222
rect 13824 -22222 14784 -22184
rect 13824 -22239 14026 -22222
rect 13564 -22256 13580 -22239
rect 12992 -22272 13580 -22256
rect 14010 -22256 14026 -22239
rect 14582 -22239 14784 -22222
rect 14842 -22222 15802 -22184
rect 14842 -22239 15044 -22222
rect 14582 -22256 14598 -22239
rect 14010 -22272 14598 -22256
rect 15028 -22256 15044 -22239
rect 15600 -22239 15802 -22222
rect 15860 -22222 16820 -22184
rect 15860 -22239 16062 -22222
rect 15600 -22256 15616 -22239
rect 15028 -22272 15616 -22256
rect 16046 -22256 16062 -22239
rect 16618 -22239 16820 -22222
rect 16878 -22222 17838 -22184
rect 16878 -22239 17080 -22222
rect 16618 -22256 16634 -22239
rect 16046 -22272 16634 -22256
rect 17064 -22256 17080 -22239
rect 17636 -22239 17838 -22222
rect 17896 -22222 18856 -22184
rect 17896 -22239 18098 -22222
rect 17636 -22256 17652 -22239
rect 17064 -22272 17652 -22256
rect 18082 -22256 18098 -22239
rect 18654 -22239 18856 -22222
rect 18914 -22222 19874 -22184
rect 18914 -22239 19116 -22222
rect 18654 -22256 18670 -22239
rect 18082 -22272 18670 -22256
rect 19100 -22256 19116 -22239
rect 19672 -22239 19874 -22222
rect 19932 -22222 20892 -22184
rect 19932 -22239 20134 -22222
rect 19672 -22256 19688 -22239
rect 19100 -22272 19688 -22256
rect 20118 -22256 20134 -22239
rect 20690 -22239 20892 -22222
rect 20950 -22222 21910 -22184
rect 20950 -22239 21152 -22222
rect 20690 -22256 20706 -22239
rect 20118 -22272 20706 -22256
rect 21136 -22256 21152 -22239
rect 21708 -22239 21910 -22222
rect 21968 -22222 22928 -22184
rect 21968 -22239 22170 -22222
rect 21708 -22256 21724 -22239
rect 21136 -22272 21724 -22256
rect 22154 -22256 22170 -22239
rect 22726 -22239 22928 -22222
rect 22726 -22256 22742 -22239
rect 22154 -22272 22742 -22256
rect -9359 -22419 -8399 -22381
rect -9359 -22436 -9157 -22419
rect -9173 -22453 -9157 -22436
rect -8601 -22436 -8399 -22419
rect -8341 -22419 -7381 -22381
rect -8341 -22436 -8139 -22419
rect -8601 -22453 -8585 -22436
rect -9173 -22469 -8585 -22453
rect -8155 -22453 -8139 -22436
rect -7583 -22436 -7381 -22419
rect -7323 -22419 -6363 -22381
rect -7323 -22436 -7121 -22419
rect -7583 -22453 -7567 -22436
rect -8155 -22469 -7567 -22453
rect -7137 -22453 -7121 -22436
rect -6565 -22436 -6363 -22419
rect -6305 -22419 -5345 -22381
rect -6305 -22436 -6103 -22419
rect -6565 -22453 -6549 -22436
rect -7137 -22469 -6549 -22453
rect -6119 -22453 -6103 -22436
rect -5547 -22436 -5345 -22419
rect -5287 -22419 -4327 -22381
rect -5287 -22436 -5085 -22419
rect -5547 -22453 -5531 -22436
rect -6119 -22469 -5531 -22453
rect -5101 -22453 -5085 -22436
rect -4529 -22436 -4327 -22419
rect -4269 -22419 -3309 -22381
rect -4269 -22436 -4067 -22419
rect -4529 -22453 -4513 -22436
rect -5101 -22469 -4513 -22453
rect -4083 -22453 -4067 -22436
rect -3511 -22436 -3309 -22419
rect -2364 -22418 -2124 -22380
rect -2364 -22435 -2306 -22418
rect -3511 -22453 -3495 -22436
rect -4083 -22469 -3495 -22453
rect -2322 -22452 -2306 -22435
rect -2182 -22435 -2124 -22418
rect -2066 -22418 -1826 -22380
rect -2066 -22435 -2008 -22418
rect -2182 -22452 -2166 -22435
rect -2322 -22468 -2166 -22452
rect -2024 -22452 -2008 -22435
rect -1884 -22435 -1826 -22418
rect -1768 -22418 -1528 -22380
rect -1768 -22435 -1710 -22418
rect -1884 -22452 -1868 -22435
rect -2024 -22468 -1868 -22452
rect -1726 -22452 -1710 -22435
rect -1586 -22435 -1528 -22418
rect -1470 -22418 -1230 -22380
rect -1470 -22435 -1412 -22418
rect -1586 -22452 -1570 -22435
rect -1726 -22468 -1570 -22452
rect -1428 -22452 -1412 -22435
rect -1288 -22435 -1230 -22418
rect -1172 -22418 -932 -22380
rect -1172 -22435 -1114 -22418
rect -1288 -22452 -1272 -22435
rect -1428 -22468 -1272 -22452
rect -1130 -22452 -1114 -22435
rect -990 -22435 -932 -22418
rect -874 -22418 -634 -22380
rect -874 -22435 -816 -22418
rect -990 -22452 -974 -22435
rect -1130 -22468 -974 -22452
rect -832 -22452 -816 -22435
rect -692 -22435 -634 -22418
rect -576 -22418 -336 -22380
rect -576 -22435 -518 -22418
rect -692 -22452 -676 -22435
rect -832 -22468 -676 -22452
rect -534 -22452 -518 -22435
rect -394 -22435 -336 -22418
rect -278 -22418 -38 -22380
rect -278 -22435 -220 -22418
rect -394 -22452 -378 -22435
rect -534 -22468 -378 -22452
rect -236 -22452 -220 -22435
rect -96 -22435 -38 -22418
rect 20 -22418 260 -22380
rect 20 -22435 78 -22418
rect -96 -22452 -80 -22435
rect -236 -22468 -80 -22452
rect 62 -22452 78 -22435
rect 202 -22435 260 -22418
rect 318 -22418 558 -22380
rect 318 -22435 376 -22418
rect 202 -22452 218 -22435
rect 62 -22468 218 -22452
rect 360 -22452 376 -22435
rect 500 -22435 558 -22418
rect 616 -22418 856 -22380
rect 616 -22435 674 -22418
rect 500 -22452 516 -22435
rect 360 -22468 516 -22452
rect 658 -22452 674 -22435
rect 798 -22435 856 -22418
rect 798 -22452 814 -22435
rect 658 -22468 814 -22452
rect 2812 -22746 3400 -22730
rect 2812 -22763 2828 -22746
rect 2626 -22780 2828 -22763
rect 3384 -22763 3400 -22746
rect 3830 -22746 4418 -22730
rect 3830 -22763 3846 -22746
rect 3384 -22780 3586 -22763
rect -9174 -22822 -8586 -22806
rect -9174 -22839 -9158 -22822
rect -9360 -22856 -9158 -22839
rect -8602 -22839 -8586 -22822
rect -8156 -22822 -7568 -22806
rect -8156 -22839 -8140 -22822
rect -8602 -22856 -8400 -22839
rect -9360 -22894 -8400 -22856
rect -8342 -22856 -8140 -22839
rect -7584 -22839 -7568 -22822
rect -7138 -22822 -6550 -22806
rect -7138 -22839 -7122 -22822
rect -7584 -22856 -7382 -22839
rect -8342 -22894 -7382 -22856
rect -7324 -22856 -7122 -22839
rect -6566 -22839 -6550 -22822
rect -6120 -22822 -5532 -22806
rect -6120 -22839 -6104 -22822
rect -6566 -22856 -6364 -22839
rect -7324 -22894 -6364 -22856
rect -6306 -22856 -6104 -22839
rect -5548 -22839 -5532 -22822
rect -5102 -22822 -4514 -22806
rect -5102 -22839 -5086 -22822
rect -5548 -22856 -5346 -22839
rect -6306 -22894 -5346 -22856
rect -5288 -22856 -5086 -22839
rect -4530 -22839 -4514 -22822
rect -4084 -22822 -3496 -22806
rect -4084 -22839 -4068 -22822
rect -4530 -22856 -4328 -22839
rect -5288 -22894 -4328 -22856
rect -4270 -22856 -4068 -22839
rect -3512 -22839 -3496 -22822
rect -2322 -22820 -2166 -22804
rect -2322 -22837 -2306 -22820
rect -3512 -22856 -3310 -22839
rect -4270 -22894 -3310 -22856
rect -2364 -22854 -2306 -22837
rect -2182 -22837 -2166 -22820
rect -2024 -22820 -1868 -22804
rect -2024 -22837 -2008 -22820
rect -2182 -22854 -2124 -22837
rect -2364 -22892 -2124 -22854
rect -2066 -22854 -2008 -22837
rect -1884 -22837 -1868 -22820
rect -1726 -22820 -1570 -22804
rect -1726 -22837 -1710 -22820
rect -1884 -22854 -1826 -22837
rect -2066 -22892 -1826 -22854
rect -1768 -22854 -1710 -22837
rect -1586 -22837 -1570 -22820
rect -1428 -22820 -1272 -22804
rect -1428 -22837 -1412 -22820
rect -1586 -22854 -1528 -22837
rect -1768 -22892 -1528 -22854
rect -1470 -22854 -1412 -22837
rect -1288 -22837 -1272 -22820
rect -1130 -22820 -974 -22804
rect -1130 -22837 -1114 -22820
rect -1288 -22854 -1230 -22837
rect -1470 -22892 -1230 -22854
rect -1172 -22854 -1114 -22837
rect -990 -22837 -974 -22820
rect -832 -22820 -676 -22804
rect -832 -22837 -816 -22820
rect -990 -22854 -932 -22837
rect -1172 -22892 -932 -22854
rect -874 -22854 -816 -22837
rect -692 -22837 -676 -22820
rect -534 -22820 -378 -22804
rect -534 -22837 -518 -22820
rect -692 -22854 -634 -22837
rect -874 -22892 -634 -22854
rect -576 -22854 -518 -22837
rect -394 -22837 -378 -22820
rect -236 -22820 -80 -22804
rect -236 -22837 -220 -22820
rect -394 -22854 -336 -22837
rect -576 -22892 -336 -22854
rect -278 -22854 -220 -22837
rect -96 -22837 -80 -22820
rect 62 -22820 218 -22804
rect 62 -22837 78 -22820
rect -96 -22854 -38 -22837
rect -278 -22892 -38 -22854
rect 20 -22854 78 -22837
rect 202 -22837 218 -22820
rect 360 -22820 516 -22804
rect 360 -22837 376 -22820
rect 202 -22854 260 -22837
rect 20 -22892 260 -22854
rect 318 -22854 376 -22837
rect 500 -22837 516 -22820
rect 658 -22820 814 -22804
rect 2626 -22818 3586 -22780
rect 3644 -22780 3846 -22763
rect 4402 -22763 4418 -22746
rect 4848 -22746 5436 -22730
rect 4848 -22763 4864 -22746
rect 4402 -22780 4604 -22763
rect 3644 -22818 4604 -22780
rect 4662 -22780 4864 -22763
rect 5420 -22763 5436 -22746
rect 5866 -22746 6454 -22730
rect 5866 -22763 5882 -22746
rect 5420 -22780 5622 -22763
rect 4662 -22818 5622 -22780
rect 5680 -22780 5882 -22763
rect 6438 -22763 6454 -22746
rect 6884 -22746 7472 -22730
rect 6884 -22763 6900 -22746
rect 6438 -22780 6640 -22763
rect 5680 -22818 6640 -22780
rect 6698 -22780 6900 -22763
rect 7456 -22763 7472 -22746
rect 7902 -22746 8490 -22730
rect 7902 -22763 7918 -22746
rect 7456 -22780 7658 -22763
rect 6698 -22818 7658 -22780
rect 7716 -22780 7918 -22763
rect 8474 -22763 8490 -22746
rect 8920 -22746 9508 -22730
rect 8920 -22763 8936 -22746
rect 8474 -22780 8676 -22763
rect 7716 -22818 8676 -22780
rect 8734 -22780 8936 -22763
rect 9492 -22763 9508 -22746
rect 9938 -22746 10526 -22730
rect 9938 -22763 9954 -22746
rect 9492 -22780 9694 -22763
rect 8734 -22818 9694 -22780
rect 9752 -22780 9954 -22763
rect 10510 -22763 10526 -22746
rect 10956 -22746 11544 -22730
rect 10956 -22763 10972 -22746
rect 10510 -22780 10712 -22763
rect 9752 -22818 10712 -22780
rect 10770 -22780 10972 -22763
rect 11528 -22763 11544 -22746
rect 11974 -22746 12562 -22730
rect 11974 -22763 11990 -22746
rect 11528 -22780 11730 -22763
rect 10770 -22818 11730 -22780
rect 11788 -22780 11990 -22763
rect 12546 -22763 12562 -22746
rect 12992 -22746 13580 -22730
rect 12992 -22763 13008 -22746
rect 12546 -22780 12748 -22763
rect 11788 -22818 12748 -22780
rect 12806 -22780 13008 -22763
rect 13564 -22763 13580 -22746
rect 14010 -22746 14598 -22730
rect 14010 -22763 14026 -22746
rect 13564 -22780 13766 -22763
rect 12806 -22818 13766 -22780
rect 13824 -22780 14026 -22763
rect 14582 -22763 14598 -22746
rect 15028 -22746 15616 -22730
rect 15028 -22763 15044 -22746
rect 14582 -22780 14784 -22763
rect 13824 -22818 14784 -22780
rect 14842 -22780 15044 -22763
rect 15600 -22763 15616 -22746
rect 16046 -22746 16634 -22730
rect 16046 -22763 16062 -22746
rect 15600 -22780 15802 -22763
rect 14842 -22818 15802 -22780
rect 15860 -22780 16062 -22763
rect 16618 -22763 16634 -22746
rect 17064 -22746 17652 -22730
rect 17064 -22763 17080 -22746
rect 16618 -22780 16820 -22763
rect 15860 -22818 16820 -22780
rect 16878 -22780 17080 -22763
rect 17636 -22763 17652 -22746
rect 18082 -22746 18670 -22730
rect 18082 -22763 18098 -22746
rect 17636 -22780 17838 -22763
rect 16878 -22818 17838 -22780
rect 17896 -22780 18098 -22763
rect 18654 -22763 18670 -22746
rect 19100 -22746 19688 -22730
rect 19100 -22763 19116 -22746
rect 18654 -22780 18856 -22763
rect 17896 -22818 18856 -22780
rect 18914 -22780 19116 -22763
rect 19672 -22763 19688 -22746
rect 20118 -22746 20706 -22730
rect 20118 -22763 20134 -22746
rect 19672 -22780 19874 -22763
rect 18914 -22818 19874 -22780
rect 19932 -22780 20134 -22763
rect 20690 -22763 20706 -22746
rect 21136 -22746 21724 -22730
rect 21136 -22763 21152 -22746
rect 20690 -22780 20892 -22763
rect 19932 -22818 20892 -22780
rect 20950 -22780 21152 -22763
rect 21708 -22763 21724 -22746
rect 22154 -22746 22742 -22730
rect 22154 -22763 22170 -22746
rect 21708 -22780 21910 -22763
rect 20950 -22818 21910 -22780
rect 21968 -22780 22170 -22763
rect 22726 -22763 22742 -22746
rect 22726 -22780 22928 -22763
rect 21968 -22818 22928 -22780
rect 658 -22837 674 -22820
rect 500 -22854 558 -22837
rect 318 -22892 558 -22854
rect 616 -22854 674 -22837
rect 798 -22837 814 -22820
rect 798 -22854 856 -22837
rect 616 -22892 856 -22854
rect 2626 -23456 3586 -23418
rect 2626 -23473 2828 -23456
rect 2812 -23490 2828 -23473
rect 3384 -23473 3586 -23456
rect 3644 -23456 4604 -23418
rect 3644 -23473 3846 -23456
rect 3384 -23490 3400 -23473
rect -9360 -23532 -8400 -23494
rect -9360 -23549 -9158 -23532
rect -9174 -23566 -9158 -23549
rect -8602 -23549 -8400 -23532
rect -8342 -23532 -7382 -23494
rect -8342 -23549 -8140 -23532
rect -8602 -23566 -8586 -23549
rect -9174 -23582 -8586 -23566
rect -8156 -23566 -8140 -23549
rect -7584 -23549 -7382 -23532
rect -7324 -23532 -6364 -23494
rect -7324 -23549 -7122 -23532
rect -7584 -23566 -7568 -23549
rect -8156 -23582 -7568 -23566
rect -7138 -23566 -7122 -23549
rect -6566 -23549 -6364 -23532
rect -6306 -23532 -5346 -23494
rect -6306 -23549 -6104 -23532
rect -6566 -23566 -6550 -23549
rect -7138 -23582 -6550 -23566
rect -6120 -23566 -6104 -23549
rect -5548 -23549 -5346 -23532
rect -5288 -23532 -4328 -23494
rect -5288 -23549 -5086 -23532
rect -5548 -23566 -5532 -23549
rect -6120 -23582 -5532 -23566
rect -5102 -23566 -5086 -23549
rect -4530 -23549 -4328 -23532
rect -4270 -23532 -3310 -23494
rect -4270 -23549 -4068 -23532
rect -4530 -23566 -4514 -23549
rect -5102 -23582 -4514 -23566
rect -4084 -23566 -4068 -23549
rect -3512 -23549 -3310 -23532
rect -2364 -23530 -2124 -23492
rect -2364 -23547 -2306 -23530
rect -3512 -23566 -3496 -23549
rect -4084 -23582 -3496 -23566
rect -2322 -23564 -2306 -23547
rect -2182 -23547 -2124 -23530
rect -2066 -23530 -1826 -23492
rect -2066 -23547 -2008 -23530
rect -2182 -23564 -2166 -23547
rect -2322 -23580 -2166 -23564
rect -2024 -23564 -2008 -23547
rect -1884 -23547 -1826 -23530
rect -1768 -23530 -1528 -23492
rect -1768 -23547 -1710 -23530
rect -1884 -23564 -1868 -23547
rect -2024 -23580 -1868 -23564
rect -1726 -23564 -1710 -23547
rect -1586 -23547 -1528 -23530
rect -1470 -23530 -1230 -23492
rect -1470 -23547 -1412 -23530
rect -1586 -23564 -1570 -23547
rect -1726 -23580 -1570 -23564
rect -1428 -23564 -1412 -23547
rect -1288 -23547 -1230 -23530
rect -1172 -23530 -932 -23492
rect -1172 -23547 -1114 -23530
rect -1288 -23564 -1272 -23547
rect -1428 -23580 -1272 -23564
rect -1130 -23564 -1114 -23547
rect -990 -23547 -932 -23530
rect -874 -23530 -634 -23492
rect -874 -23547 -816 -23530
rect -990 -23564 -974 -23547
rect -1130 -23580 -974 -23564
rect -832 -23564 -816 -23547
rect -692 -23547 -634 -23530
rect -576 -23530 -336 -23492
rect -576 -23547 -518 -23530
rect -692 -23564 -676 -23547
rect -832 -23580 -676 -23564
rect -534 -23564 -518 -23547
rect -394 -23547 -336 -23530
rect -278 -23530 -38 -23492
rect -278 -23547 -220 -23530
rect -394 -23564 -378 -23547
rect -534 -23580 -378 -23564
rect -236 -23564 -220 -23547
rect -96 -23547 -38 -23530
rect 20 -23530 260 -23492
rect 20 -23547 78 -23530
rect -96 -23564 -80 -23547
rect -236 -23580 -80 -23564
rect 62 -23564 78 -23547
rect 202 -23547 260 -23530
rect 318 -23530 558 -23492
rect 318 -23547 376 -23530
rect 202 -23564 218 -23547
rect 62 -23580 218 -23564
rect 360 -23564 376 -23547
rect 500 -23547 558 -23530
rect 616 -23530 856 -23492
rect 2812 -23506 3400 -23490
rect 3830 -23490 3846 -23473
rect 4402 -23473 4604 -23456
rect 4662 -23456 5622 -23418
rect 4662 -23473 4864 -23456
rect 4402 -23490 4418 -23473
rect 3830 -23506 4418 -23490
rect 4848 -23490 4864 -23473
rect 5420 -23473 5622 -23456
rect 5680 -23456 6640 -23418
rect 5680 -23473 5882 -23456
rect 5420 -23490 5436 -23473
rect 4848 -23506 5436 -23490
rect 5866 -23490 5882 -23473
rect 6438 -23473 6640 -23456
rect 6698 -23456 7658 -23418
rect 6698 -23473 6900 -23456
rect 6438 -23490 6454 -23473
rect 5866 -23506 6454 -23490
rect 6884 -23490 6900 -23473
rect 7456 -23473 7658 -23456
rect 7716 -23456 8676 -23418
rect 7716 -23473 7918 -23456
rect 7456 -23490 7472 -23473
rect 6884 -23506 7472 -23490
rect 7902 -23490 7918 -23473
rect 8474 -23473 8676 -23456
rect 8734 -23456 9694 -23418
rect 8734 -23473 8936 -23456
rect 8474 -23490 8490 -23473
rect 7902 -23506 8490 -23490
rect 8920 -23490 8936 -23473
rect 9492 -23473 9694 -23456
rect 9752 -23456 10712 -23418
rect 9752 -23473 9954 -23456
rect 9492 -23490 9508 -23473
rect 8920 -23506 9508 -23490
rect 9938 -23490 9954 -23473
rect 10510 -23473 10712 -23456
rect 10770 -23456 11730 -23418
rect 10770 -23473 10972 -23456
rect 10510 -23490 10526 -23473
rect 9938 -23506 10526 -23490
rect 10956 -23490 10972 -23473
rect 11528 -23473 11730 -23456
rect 11788 -23456 12748 -23418
rect 11788 -23473 11990 -23456
rect 11528 -23490 11544 -23473
rect 10956 -23506 11544 -23490
rect 11974 -23490 11990 -23473
rect 12546 -23473 12748 -23456
rect 12806 -23456 13766 -23418
rect 12806 -23473 13008 -23456
rect 12546 -23490 12562 -23473
rect 11974 -23506 12562 -23490
rect 12992 -23490 13008 -23473
rect 13564 -23473 13766 -23456
rect 13824 -23456 14784 -23418
rect 13824 -23473 14026 -23456
rect 13564 -23490 13580 -23473
rect 12992 -23506 13580 -23490
rect 14010 -23490 14026 -23473
rect 14582 -23473 14784 -23456
rect 14842 -23456 15802 -23418
rect 14842 -23473 15044 -23456
rect 14582 -23490 14598 -23473
rect 14010 -23506 14598 -23490
rect 15028 -23490 15044 -23473
rect 15600 -23473 15802 -23456
rect 15860 -23456 16820 -23418
rect 15860 -23473 16062 -23456
rect 15600 -23490 15616 -23473
rect 15028 -23506 15616 -23490
rect 16046 -23490 16062 -23473
rect 16618 -23473 16820 -23456
rect 16878 -23456 17838 -23418
rect 16878 -23473 17080 -23456
rect 16618 -23490 16634 -23473
rect 16046 -23506 16634 -23490
rect 17064 -23490 17080 -23473
rect 17636 -23473 17838 -23456
rect 17896 -23456 18856 -23418
rect 17896 -23473 18098 -23456
rect 17636 -23490 17652 -23473
rect 17064 -23506 17652 -23490
rect 18082 -23490 18098 -23473
rect 18654 -23473 18856 -23456
rect 18914 -23456 19874 -23418
rect 18914 -23473 19116 -23456
rect 18654 -23490 18670 -23473
rect 18082 -23506 18670 -23490
rect 19100 -23490 19116 -23473
rect 19672 -23473 19874 -23456
rect 19932 -23456 20892 -23418
rect 19932 -23473 20134 -23456
rect 19672 -23490 19688 -23473
rect 19100 -23506 19688 -23490
rect 20118 -23490 20134 -23473
rect 20690 -23473 20892 -23456
rect 20950 -23456 21910 -23418
rect 20950 -23473 21152 -23456
rect 20690 -23490 20706 -23473
rect 20118 -23506 20706 -23490
rect 21136 -23490 21152 -23473
rect 21708 -23473 21910 -23456
rect 21968 -23456 22928 -23418
rect 21968 -23473 22170 -23456
rect 21708 -23490 21724 -23473
rect 21136 -23506 21724 -23490
rect 22154 -23490 22170 -23473
rect 22726 -23473 22928 -23456
rect 22726 -23490 22742 -23473
rect 22154 -23506 22742 -23490
rect 616 -23547 674 -23530
rect 500 -23564 516 -23547
rect 360 -23580 516 -23564
rect 658 -23564 674 -23547
rect 798 -23547 856 -23530
rect 798 -23564 814 -23547
rect 658 -23580 814 -23564
rect -9173 -23933 -8585 -23917
rect -9173 -23950 -9157 -23933
rect -9359 -23967 -9157 -23950
rect -8601 -23950 -8585 -23933
rect -8155 -23933 -7567 -23917
rect -8155 -23950 -8139 -23933
rect -8601 -23967 -8399 -23950
rect -9359 -24005 -8399 -23967
rect -8341 -23967 -8139 -23950
rect -7583 -23950 -7567 -23933
rect -7137 -23933 -6549 -23917
rect -7137 -23950 -7121 -23933
rect -7583 -23967 -7381 -23950
rect -8341 -24005 -7381 -23967
rect -7323 -23967 -7121 -23950
rect -6565 -23950 -6549 -23933
rect -6119 -23933 -5531 -23917
rect -6119 -23950 -6103 -23933
rect -6565 -23967 -6363 -23950
rect -7323 -24005 -6363 -23967
rect -6305 -23967 -6103 -23950
rect -5547 -23950 -5531 -23933
rect -5101 -23933 -4513 -23917
rect -5101 -23950 -5085 -23933
rect -5547 -23967 -5345 -23950
rect -6305 -24005 -5345 -23967
rect -5287 -23967 -5085 -23950
rect -4529 -23950 -4513 -23933
rect -4083 -23933 -3495 -23917
rect -4083 -23950 -4067 -23933
rect -4529 -23967 -4327 -23950
rect -5287 -24005 -4327 -23967
rect -4269 -23967 -4067 -23950
rect -3511 -23950 -3495 -23933
rect -2324 -23932 -2168 -23916
rect -2324 -23949 -2308 -23932
rect -3511 -23967 -3309 -23950
rect -4269 -24005 -3309 -23967
rect -2366 -23966 -2308 -23949
rect -2184 -23949 -2168 -23932
rect -2026 -23932 -1870 -23916
rect -2026 -23949 -2010 -23932
rect -2184 -23966 -2126 -23949
rect -2366 -24004 -2126 -23966
rect -2068 -23966 -2010 -23949
rect -1886 -23949 -1870 -23932
rect -1728 -23932 -1572 -23916
rect -1728 -23949 -1712 -23932
rect -1886 -23966 -1828 -23949
rect -2068 -24004 -1828 -23966
rect -1770 -23966 -1712 -23949
rect -1588 -23949 -1572 -23932
rect -1430 -23932 -1274 -23916
rect -1430 -23949 -1414 -23932
rect -1588 -23966 -1530 -23949
rect -1770 -24004 -1530 -23966
rect -1472 -23966 -1414 -23949
rect -1290 -23949 -1274 -23932
rect -1132 -23932 -976 -23916
rect -1132 -23949 -1116 -23932
rect -1290 -23966 -1232 -23949
rect -1472 -24004 -1232 -23966
rect -1174 -23966 -1116 -23949
rect -992 -23949 -976 -23932
rect -834 -23932 -678 -23916
rect -834 -23949 -818 -23932
rect -992 -23966 -934 -23949
rect -1174 -24004 -934 -23966
rect -876 -23966 -818 -23949
rect -694 -23949 -678 -23932
rect -536 -23932 -380 -23916
rect -536 -23949 -520 -23932
rect -694 -23966 -636 -23949
rect -876 -24004 -636 -23966
rect -578 -23966 -520 -23949
rect -396 -23949 -380 -23932
rect -238 -23932 -82 -23916
rect -238 -23949 -222 -23932
rect -396 -23966 -338 -23949
rect -578 -24004 -338 -23966
rect -280 -23966 -222 -23949
rect -98 -23949 -82 -23932
rect 60 -23932 216 -23916
rect 60 -23949 76 -23932
rect -98 -23966 -40 -23949
rect -280 -24004 -40 -23966
rect 18 -23966 76 -23949
rect 200 -23949 216 -23932
rect 358 -23932 514 -23916
rect 358 -23949 374 -23932
rect 200 -23966 258 -23949
rect 18 -24004 258 -23966
rect 316 -23966 374 -23949
rect 498 -23949 514 -23932
rect 656 -23932 812 -23916
rect 656 -23949 672 -23932
rect 498 -23966 556 -23949
rect 316 -24004 556 -23966
rect 614 -23966 672 -23949
rect 796 -23949 812 -23932
rect 796 -23966 854 -23949
rect 614 -24004 854 -23966
rect 2812 -23980 3400 -23964
rect 2812 -23997 2828 -23980
rect 2626 -24014 2828 -23997
rect 3384 -23997 3400 -23980
rect 3830 -23980 4418 -23964
rect 3830 -23997 3846 -23980
rect 3384 -24014 3586 -23997
rect 2626 -24052 3586 -24014
rect 3644 -24014 3846 -23997
rect 4402 -23997 4418 -23980
rect 4848 -23980 5436 -23964
rect 4848 -23997 4864 -23980
rect 4402 -24014 4604 -23997
rect 3644 -24052 4604 -24014
rect 4662 -24014 4864 -23997
rect 5420 -23997 5436 -23980
rect 5866 -23980 6454 -23964
rect 5866 -23997 5882 -23980
rect 5420 -24014 5622 -23997
rect 4662 -24052 5622 -24014
rect 5680 -24014 5882 -23997
rect 6438 -23997 6454 -23980
rect 6884 -23980 7472 -23964
rect 6884 -23997 6900 -23980
rect 6438 -24014 6640 -23997
rect 5680 -24052 6640 -24014
rect 6698 -24014 6900 -23997
rect 7456 -23997 7472 -23980
rect 7902 -23980 8490 -23964
rect 7902 -23997 7918 -23980
rect 7456 -24014 7658 -23997
rect 6698 -24052 7658 -24014
rect 7716 -24014 7918 -23997
rect 8474 -23997 8490 -23980
rect 8920 -23980 9508 -23964
rect 8920 -23997 8936 -23980
rect 8474 -24014 8676 -23997
rect 7716 -24052 8676 -24014
rect 8734 -24014 8936 -23997
rect 9492 -23997 9508 -23980
rect 9938 -23980 10526 -23964
rect 9938 -23997 9954 -23980
rect 9492 -24014 9694 -23997
rect 8734 -24052 9694 -24014
rect 9752 -24014 9954 -23997
rect 10510 -23997 10526 -23980
rect 10956 -23980 11544 -23964
rect 10956 -23997 10972 -23980
rect 10510 -24014 10712 -23997
rect 9752 -24052 10712 -24014
rect 10770 -24014 10972 -23997
rect 11528 -23997 11544 -23980
rect 11974 -23980 12562 -23964
rect 11974 -23997 11990 -23980
rect 11528 -24014 11730 -23997
rect 10770 -24052 11730 -24014
rect 11788 -24014 11990 -23997
rect 12546 -23997 12562 -23980
rect 12992 -23980 13580 -23964
rect 12992 -23997 13008 -23980
rect 12546 -24014 12748 -23997
rect 11788 -24052 12748 -24014
rect 12806 -24014 13008 -23997
rect 13564 -23997 13580 -23980
rect 14010 -23980 14598 -23964
rect 14010 -23997 14026 -23980
rect 13564 -24014 13766 -23997
rect 12806 -24052 13766 -24014
rect 13824 -24014 14026 -23997
rect 14582 -23997 14598 -23980
rect 15028 -23980 15616 -23964
rect 15028 -23997 15044 -23980
rect 14582 -24014 14784 -23997
rect 13824 -24052 14784 -24014
rect 14842 -24014 15044 -23997
rect 15600 -23997 15616 -23980
rect 16046 -23980 16634 -23964
rect 16046 -23997 16062 -23980
rect 15600 -24014 15802 -23997
rect 14842 -24052 15802 -24014
rect 15860 -24014 16062 -23997
rect 16618 -23997 16634 -23980
rect 17064 -23980 17652 -23964
rect 17064 -23997 17080 -23980
rect 16618 -24014 16820 -23997
rect 15860 -24052 16820 -24014
rect 16878 -24014 17080 -23997
rect 17636 -23997 17652 -23980
rect 18082 -23980 18670 -23964
rect 18082 -23997 18098 -23980
rect 17636 -24014 17838 -23997
rect 16878 -24052 17838 -24014
rect 17896 -24014 18098 -23997
rect 18654 -23997 18670 -23980
rect 19100 -23980 19688 -23964
rect 19100 -23997 19116 -23980
rect 18654 -24014 18856 -23997
rect 17896 -24052 18856 -24014
rect 18914 -24014 19116 -23997
rect 19672 -23997 19688 -23980
rect 20118 -23980 20706 -23964
rect 20118 -23997 20134 -23980
rect 19672 -24014 19874 -23997
rect 18914 -24052 19874 -24014
rect 19932 -24014 20134 -23997
rect 20690 -23997 20706 -23980
rect 21136 -23980 21724 -23964
rect 21136 -23997 21152 -23980
rect 20690 -24014 20892 -23997
rect 19932 -24052 20892 -24014
rect 20950 -24014 21152 -23997
rect 21708 -23997 21724 -23980
rect 22154 -23980 22742 -23964
rect 22154 -23997 22170 -23980
rect 21708 -24014 21910 -23997
rect 20950 -24052 21910 -24014
rect 21968 -24014 22170 -23997
rect 22726 -23997 22742 -23980
rect 22726 -24014 22928 -23997
rect 21968 -24052 22928 -24014
rect -9359 -24643 -8399 -24605
rect -9359 -24660 -9157 -24643
rect -9173 -24677 -9157 -24660
rect -8601 -24660 -8399 -24643
rect -8341 -24643 -7381 -24605
rect -8341 -24660 -8139 -24643
rect -8601 -24677 -8585 -24660
rect -9173 -24693 -8585 -24677
rect -8155 -24677 -8139 -24660
rect -7583 -24660 -7381 -24643
rect -7323 -24643 -6363 -24605
rect -7323 -24660 -7121 -24643
rect -7583 -24677 -7567 -24660
rect -8155 -24693 -7567 -24677
rect -7137 -24677 -7121 -24660
rect -6565 -24660 -6363 -24643
rect -6305 -24643 -5345 -24605
rect -6305 -24660 -6103 -24643
rect -6565 -24677 -6549 -24660
rect -7137 -24693 -6549 -24677
rect -6119 -24677 -6103 -24660
rect -5547 -24660 -5345 -24643
rect -5287 -24643 -4327 -24605
rect -5287 -24660 -5085 -24643
rect -5547 -24677 -5531 -24660
rect -6119 -24693 -5531 -24677
rect -5101 -24677 -5085 -24660
rect -4529 -24660 -4327 -24643
rect -4269 -24643 -3309 -24605
rect -4269 -24660 -4067 -24643
rect -4529 -24677 -4513 -24660
rect -5101 -24693 -4513 -24677
rect -4083 -24677 -4067 -24660
rect -3511 -24660 -3309 -24643
rect -2366 -24642 -2126 -24604
rect -2366 -24659 -2308 -24642
rect -3511 -24677 -3495 -24660
rect -4083 -24693 -3495 -24677
rect -2324 -24676 -2308 -24659
rect -2184 -24659 -2126 -24642
rect -2068 -24642 -1828 -24604
rect -2068 -24659 -2010 -24642
rect -2184 -24676 -2168 -24659
rect -2324 -24692 -2168 -24676
rect -2026 -24676 -2010 -24659
rect -1886 -24659 -1828 -24642
rect -1770 -24642 -1530 -24604
rect -1770 -24659 -1712 -24642
rect -1886 -24676 -1870 -24659
rect -2026 -24692 -1870 -24676
rect -1728 -24676 -1712 -24659
rect -1588 -24659 -1530 -24642
rect -1472 -24642 -1232 -24604
rect -1472 -24659 -1414 -24642
rect -1588 -24676 -1572 -24659
rect -1728 -24692 -1572 -24676
rect -1430 -24676 -1414 -24659
rect -1290 -24659 -1232 -24642
rect -1174 -24642 -934 -24604
rect -1174 -24659 -1116 -24642
rect -1290 -24676 -1274 -24659
rect -1430 -24692 -1274 -24676
rect -1132 -24676 -1116 -24659
rect -992 -24659 -934 -24642
rect -876 -24642 -636 -24604
rect -876 -24659 -818 -24642
rect -992 -24676 -976 -24659
rect -1132 -24692 -976 -24676
rect -834 -24676 -818 -24659
rect -694 -24659 -636 -24642
rect -578 -24642 -338 -24604
rect -578 -24659 -520 -24642
rect -694 -24676 -678 -24659
rect -834 -24692 -678 -24676
rect -536 -24676 -520 -24659
rect -396 -24659 -338 -24642
rect -280 -24642 -40 -24604
rect -280 -24659 -222 -24642
rect -396 -24676 -380 -24659
rect -536 -24692 -380 -24676
rect -238 -24676 -222 -24659
rect -98 -24659 -40 -24642
rect 18 -24642 258 -24604
rect 18 -24659 76 -24642
rect -98 -24676 -82 -24659
rect -238 -24692 -82 -24676
rect 60 -24676 76 -24659
rect 200 -24659 258 -24642
rect 316 -24642 556 -24604
rect 316 -24659 374 -24642
rect 200 -24676 216 -24659
rect 60 -24692 216 -24676
rect 358 -24676 374 -24659
rect 498 -24659 556 -24642
rect 614 -24642 854 -24604
rect 614 -24659 672 -24642
rect 498 -24676 514 -24659
rect 358 -24692 514 -24676
rect 656 -24676 672 -24659
rect 796 -24659 854 -24642
rect 796 -24676 812 -24659
rect 656 -24692 812 -24676
rect 2626 -24690 3586 -24652
rect 2626 -24707 2828 -24690
rect 2812 -24724 2828 -24707
rect 3384 -24707 3586 -24690
rect 3644 -24690 4604 -24652
rect 3644 -24707 3846 -24690
rect 3384 -24724 3400 -24707
rect 2812 -24740 3400 -24724
rect 3830 -24724 3846 -24707
rect 4402 -24707 4604 -24690
rect 4662 -24690 5622 -24652
rect 4662 -24707 4864 -24690
rect 4402 -24724 4418 -24707
rect 3830 -24740 4418 -24724
rect 4848 -24724 4864 -24707
rect 5420 -24707 5622 -24690
rect 5680 -24690 6640 -24652
rect 5680 -24707 5882 -24690
rect 5420 -24724 5436 -24707
rect 4848 -24740 5436 -24724
rect 5866 -24724 5882 -24707
rect 6438 -24707 6640 -24690
rect 6698 -24690 7658 -24652
rect 6698 -24707 6900 -24690
rect 6438 -24724 6454 -24707
rect 5866 -24740 6454 -24724
rect 6884 -24724 6900 -24707
rect 7456 -24707 7658 -24690
rect 7716 -24690 8676 -24652
rect 7716 -24707 7918 -24690
rect 7456 -24724 7472 -24707
rect 6884 -24740 7472 -24724
rect 7902 -24724 7918 -24707
rect 8474 -24707 8676 -24690
rect 8734 -24690 9694 -24652
rect 8734 -24707 8936 -24690
rect 8474 -24724 8490 -24707
rect 7902 -24740 8490 -24724
rect 8920 -24724 8936 -24707
rect 9492 -24707 9694 -24690
rect 9752 -24690 10712 -24652
rect 9752 -24707 9954 -24690
rect 9492 -24724 9508 -24707
rect 8920 -24740 9508 -24724
rect 9938 -24724 9954 -24707
rect 10510 -24707 10712 -24690
rect 10770 -24690 11730 -24652
rect 10770 -24707 10972 -24690
rect 10510 -24724 10526 -24707
rect 9938 -24740 10526 -24724
rect 10956 -24724 10972 -24707
rect 11528 -24707 11730 -24690
rect 11788 -24690 12748 -24652
rect 11788 -24707 11990 -24690
rect 11528 -24724 11544 -24707
rect 10956 -24740 11544 -24724
rect 11974 -24724 11990 -24707
rect 12546 -24707 12748 -24690
rect 12806 -24690 13766 -24652
rect 12806 -24707 13008 -24690
rect 12546 -24724 12562 -24707
rect 11974 -24740 12562 -24724
rect 12992 -24724 13008 -24707
rect 13564 -24707 13766 -24690
rect 13824 -24690 14784 -24652
rect 13824 -24707 14026 -24690
rect 13564 -24724 13580 -24707
rect 12992 -24740 13580 -24724
rect 14010 -24724 14026 -24707
rect 14582 -24707 14784 -24690
rect 14842 -24690 15802 -24652
rect 14842 -24707 15044 -24690
rect 14582 -24724 14598 -24707
rect 14010 -24740 14598 -24724
rect 15028 -24724 15044 -24707
rect 15600 -24707 15802 -24690
rect 15860 -24690 16820 -24652
rect 15860 -24707 16062 -24690
rect 15600 -24724 15616 -24707
rect 15028 -24740 15616 -24724
rect 16046 -24724 16062 -24707
rect 16618 -24707 16820 -24690
rect 16878 -24690 17838 -24652
rect 16878 -24707 17080 -24690
rect 16618 -24724 16634 -24707
rect 16046 -24740 16634 -24724
rect 17064 -24724 17080 -24707
rect 17636 -24707 17838 -24690
rect 17896 -24690 18856 -24652
rect 17896 -24707 18098 -24690
rect 17636 -24724 17652 -24707
rect 17064 -24740 17652 -24724
rect 18082 -24724 18098 -24707
rect 18654 -24707 18856 -24690
rect 18914 -24690 19874 -24652
rect 18914 -24707 19116 -24690
rect 18654 -24724 18670 -24707
rect 18082 -24740 18670 -24724
rect 19100 -24724 19116 -24707
rect 19672 -24707 19874 -24690
rect 19932 -24690 20892 -24652
rect 19932 -24707 20134 -24690
rect 19672 -24724 19688 -24707
rect 19100 -24740 19688 -24724
rect 20118 -24724 20134 -24707
rect 20690 -24707 20892 -24690
rect 20950 -24690 21910 -24652
rect 20950 -24707 21152 -24690
rect 20690 -24724 20706 -24707
rect 20118 -24740 20706 -24724
rect 21136 -24724 21152 -24707
rect 21708 -24707 21910 -24690
rect 21968 -24690 22928 -24652
rect 21968 -24707 22170 -24690
rect 21708 -24724 21724 -24707
rect 21136 -24740 21724 -24724
rect 22154 -24724 22170 -24707
rect 22726 -24707 22928 -24690
rect 22726 -24724 22742 -24707
rect 22154 -24740 22742 -24724
rect -9174 -25046 -8586 -25030
rect -9174 -25063 -9158 -25046
rect -9360 -25080 -9158 -25063
rect -8602 -25063 -8586 -25046
rect -8156 -25046 -7568 -25030
rect -8156 -25063 -8140 -25046
rect -8602 -25080 -8400 -25063
rect -9360 -25118 -8400 -25080
rect -8342 -25080 -8140 -25063
rect -7584 -25063 -7568 -25046
rect -7138 -25046 -6550 -25030
rect -7138 -25063 -7122 -25046
rect -7584 -25080 -7382 -25063
rect -8342 -25118 -7382 -25080
rect -7324 -25080 -7122 -25063
rect -6566 -25063 -6550 -25046
rect -6120 -25046 -5532 -25030
rect -6120 -25063 -6104 -25046
rect -6566 -25080 -6364 -25063
rect -7324 -25118 -6364 -25080
rect -6306 -25080 -6104 -25063
rect -5548 -25063 -5532 -25046
rect -5102 -25046 -4514 -25030
rect -5102 -25063 -5086 -25046
rect -5548 -25080 -5346 -25063
rect -6306 -25118 -5346 -25080
rect -5288 -25080 -5086 -25063
rect -4530 -25063 -4514 -25046
rect -4084 -25046 -3496 -25030
rect -4084 -25063 -4068 -25046
rect -4530 -25080 -4328 -25063
rect -5288 -25118 -4328 -25080
rect -4270 -25080 -4068 -25063
rect -3512 -25063 -3496 -25046
rect -2324 -25042 -2168 -25026
rect -2324 -25059 -2308 -25042
rect -3512 -25080 -3310 -25063
rect -4270 -25118 -3310 -25080
rect -2366 -25076 -2308 -25059
rect -2184 -25059 -2168 -25042
rect -2026 -25042 -1870 -25026
rect -2026 -25059 -2010 -25042
rect -2184 -25076 -2126 -25059
rect -2366 -25114 -2126 -25076
rect -2068 -25076 -2010 -25059
rect -1886 -25059 -1870 -25042
rect -1728 -25042 -1572 -25026
rect -1728 -25059 -1712 -25042
rect -1886 -25076 -1828 -25059
rect -2068 -25114 -1828 -25076
rect -1770 -25076 -1712 -25059
rect -1588 -25059 -1572 -25042
rect -1430 -25042 -1274 -25026
rect -1430 -25059 -1414 -25042
rect -1588 -25076 -1530 -25059
rect -1770 -25114 -1530 -25076
rect -1472 -25076 -1414 -25059
rect -1290 -25059 -1274 -25042
rect -1132 -25042 -976 -25026
rect -1132 -25059 -1116 -25042
rect -1290 -25076 -1232 -25059
rect -1472 -25114 -1232 -25076
rect -1174 -25076 -1116 -25059
rect -992 -25059 -976 -25042
rect -834 -25042 -678 -25026
rect -834 -25059 -818 -25042
rect -992 -25076 -934 -25059
rect -1174 -25114 -934 -25076
rect -876 -25076 -818 -25059
rect -694 -25059 -678 -25042
rect -536 -25042 -380 -25026
rect -536 -25059 -520 -25042
rect -694 -25076 -636 -25059
rect -876 -25114 -636 -25076
rect -578 -25076 -520 -25059
rect -396 -25059 -380 -25042
rect -238 -25042 -82 -25026
rect -238 -25059 -222 -25042
rect -396 -25076 -338 -25059
rect -578 -25114 -338 -25076
rect -280 -25076 -222 -25059
rect -98 -25059 -82 -25042
rect 60 -25042 216 -25026
rect 60 -25059 76 -25042
rect -98 -25076 -40 -25059
rect -280 -25114 -40 -25076
rect 18 -25076 76 -25059
rect 200 -25059 216 -25042
rect 358 -25042 514 -25026
rect 358 -25059 374 -25042
rect 200 -25076 258 -25059
rect 18 -25114 258 -25076
rect 316 -25076 374 -25059
rect 498 -25059 514 -25042
rect 656 -25042 812 -25026
rect 656 -25059 672 -25042
rect 498 -25076 556 -25059
rect 316 -25114 556 -25076
rect 614 -25076 672 -25059
rect 796 -25059 812 -25042
rect 796 -25076 854 -25059
rect 614 -25114 854 -25076
rect 2812 -25212 3400 -25196
rect 2812 -25229 2828 -25212
rect 2626 -25246 2828 -25229
rect 3384 -25229 3400 -25212
rect 3830 -25212 4418 -25196
rect 3830 -25229 3846 -25212
rect 3384 -25246 3586 -25229
rect 2626 -25284 3586 -25246
rect 3644 -25246 3846 -25229
rect 4402 -25229 4418 -25212
rect 4848 -25212 5436 -25196
rect 4848 -25229 4864 -25212
rect 4402 -25246 4604 -25229
rect 3644 -25284 4604 -25246
rect 4662 -25246 4864 -25229
rect 5420 -25229 5436 -25212
rect 5866 -25212 6454 -25196
rect 5866 -25229 5882 -25212
rect 5420 -25246 5622 -25229
rect 4662 -25284 5622 -25246
rect 5680 -25246 5882 -25229
rect 6438 -25229 6454 -25212
rect 6884 -25212 7472 -25196
rect 6884 -25229 6900 -25212
rect 6438 -25246 6640 -25229
rect 5680 -25284 6640 -25246
rect 6698 -25246 6900 -25229
rect 7456 -25229 7472 -25212
rect 7902 -25212 8490 -25196
rect 7902 -25229 7918 -25212
rect 7456 -25246 7658 -25229
rect 6698 -25284 7658 -25246
rect 7716 -25246 7918 -25229
rect 8474 -25229 8490 -25212
rect 8920 -25212 9508 -25196
rect 8920 -25229 8936 -25212
rect 8474 -25246 8676 -25229
rect 7716 -25284 8676 -25246
rect 8734 -25246 8936 -25229
rect 9492 -25229 9508 -25212
rect 9938 -25212 10526 -25196
rect 9938 -25229 9954 -25212
rect 9492 -25246 9694 -25229
rect 8734 -25284 9694 -25246
rect 9752 -25246 9954 -25229
rect 10510 -25229 10526 -25212
rect 10956 -25212 11544 -25196
rect 10956 -25229 10972 -25212
rect 10510 -25246 10712 -25229
rect 9752 -25284 10712 -25246
rect 10770 -25246 10972 -25229
rect 11528 -25229 11544 -25212
rect 11974 -25212 12562 -25196
rect 11974 -25229 11990 -25212
rect 11528 -25246 11730 -25229
rect 10770 -25284 11730 -25246
rect 11788 -25246 11990 -25229
rect 12546 -25229 12562 -25212
rect 12992 -25212 13580 -25196
rect 12992 -25229 13008 -25212
rect 12546 -25246 12748 -25229
rect 11788 -25284 12748 -25246
rect 12806 -25246 13008 -25229
rect 13564 -25229 13580 -25212
rect 14010 -25212 14598 -25196
rect 14010 -25229 14026 -25212
rect 13564 -25246 13766 -25229
rect 12806 -25284 13766 -25246
rect 13824 -25246 14026 -25229
rect 14582 -25229 14598 -25212
rect 15028 -25212 15616 -25196
rect 15028 -25229 15044 -25212
rect 14582 -25246 14784 -25229
rect 13824 -25284 14784 -25246
rect 14842 -25246 15044 -25229
rect 15600 -25229 15616 -25212
rect 16046 -25212 16634 -25196
rect 16046 -25229 16062 -25212
rect 15600 -25246 15802 -25229
rect 14842 -25284 15802 -25246
rect 15860 -25246 16062 -25229
rect 16618 -25229 16634 -25212
rect 17064 -25212 17652 -25196
rect 17064 -25229 17080 -25212
rect 16618 -25246 16820 -25229
rect 15860 -25284 16820 -25246
rect 16878 -25246 17080 -25229
rect 17636 -25229 17652 -25212
rect 18082 -25212 18670 -25196
rect 18082 -25229 18098 -25212
rect 17636 -25246 17838 -25229
rect 16878 -25284 17838 -25246
rect 17896 -25246 18098 -25229
rect 18654 -25229 18670 -25212
rect 19100 -25212 19688 -25196
rect 19100 -25229 19116 -25212
rect 18654 -25246 18856 -25229
rect 17896 -25284 18856 -25246
rect 18914 -25246 19116 -25229
rect 19672 -25229 19688 -25212
rect 20118 -25212 20706 -25196
rect 20118 -25229 20134 -25212
rect 19672 -25246 19874 -25229
rect 18914 -25284 19874 -25246
rect 19932 -25246 20134 -25229
rect 20690 -25229 20706 -25212
rect 21136 -25212 21724 -25196
rect 21136 -25229 21152 -25212
rect 20690 -25246 20892 -25229
rect 19932 -25284 20892 -25246
rect 20950 -25246 21152 -25229
rect 21708 -25229 21724 -25212
rect 22154 -25212 22742 -25196
rect 22154 -25229 22170 -25212
rect 21708 -25246 21910 -25229
rect 20950 -25284 21910 -25246
rect 21968 -25246 22170 -25229
rect 22726 -25229 22742 -25212
rect 22726 -25246 22928 -25229
rect 21968 -25284 22928 -25246
rect -9360 -25756 -8400 -25718
rect -9360 -25773 -9158 -25756
rect -9174 -25790 -9158 -25773
rect -8602 -25773 -8400 -25756
rect -8342 -25756 -7382 -25718
rect -8342 -25773 -8140 -25756
rect -8602 -25790 -8586 -25773
rect -9174 -25806 -8586 -25790
rect -8156 -25790 -8140 -25773
rect -7584 -25773 -7382 -25756
rect -7324 -25756 -6364 -25718
rect -7324 -25773 -7122 -25756
rect -7584 -25790 -7568 -25773
rect -8156 -25806 -7568 -25790
rect -7138 -25790 -7122 -25773
rect -6566 -25773 -6364 -25756
rect -6306 -25756 -5346 -25718
rect -6306 -25773 -6104 -25756
rect -6566 -25790 -6550 -25773
rect -7138 -25806 -6550 -25790
rect -6120 -25790 -6104 -25773
rect -5548 -25773 -5346 -25756
rect -5288 -25756 -4328 -25718
rect -5288 -25773 -5086 -25756
rect -5548 -25790 -5532 -25773
rect -6120 -25806 -5532 -25790
rect -5102 -25790 -5086 -25773
rect -4530 -25773 -4328 -25756
rect -4270 -25756 -3310 -25718
rect -4270 -25773 -4068 -25756
rect -4530 -25790 -4514 -25773
rect -5102 -25806 -4514 -25790
rect -4084 -25790 -4068 -25773
rect -3512 -25773 -3310 -25756
rect -2366 -25752 -2126 -25714
rect -2366 -25769 -2308 -25752
rect -3512 -25790 -3496 -25773
rect -4084 -25806 -3496 -25790
rect -2324 -25786 -2308 -25769
rect -2184 -25769 -2126 -25752
rect -2068 -25752 -1828 -25714
rect -2068 -25769 -2010 -25752
rect -2184 -25786 -2168 -25769
rect -2324 -25802 -2168 -25786
rect -2026 -25786 -2010 -25769
rect -1886 -25769 -1828 -25752
rect -1770 -25752 -1530 -25714
rect -1770 -25769 -1712 -25752
rect -1886 -25786 -1870 -25769
rect -2026 -25802 -1870 -25786
rect -1728 -25786 -1712 -25769
rect -1588 -25769 -1530 -25752
rect -1472 -25752 -1232 -25714
rect -1472 -25769 -1414 -25752
rect -1588 -25786 -1572 -25769
rect -1728 -25802 -1572 -25786
rect -1430 -25786 -1414 -25769
rect -1290 -25769 -1232 -25752
rect -1174 -25752 -934 -25714
rect -1174 -25769 -1116 -25752
rect -1290 -25786 -1274 -25769
rect -1430 -25802 -1274 -25786
rect -1132 -25786 -1116 -25769
rect -992 -25769 -934 -25752
rect -876 -25752 -636 -25714
rect -876 -25769 -818 -25752
rect -992 -25786 -976 -25769
rect -1132 -25802 -976 -25786
rect -834 -25786 -818 -25769
rect -694 -25769 -636 -25752
rect -578 -25752 -338 -25714
rect -578 -25769 -520 -25752
rect -694 -25786 -678 -25769
rect -834 -25802 -678 -25786
rect -536 -25786 -520 -25769
rect -396 -25769 -338 -25752
rect -280 -25752 -40 -25714
rect -280 -25769 -222 -25752
rect -396 -25786 -380 -25769
rect -536 -25802 -380 -25786
rect -238 -25786 -222 -25769
rect -98 -25769 -40 -25752
rect 18 -25752 258 -25714
rect 18 -25769 76 -25752
rect -98 -25786 -82 -25769
rect -238 -25802 -82 -25786
rect 60 -25786 76 -25769
rect 200 -25769 258 -25752
rect 316 -25752 556 -25714
rect 316 -25769 374 -25752
rect 200 -25786 216 -25769
rect 60 -25802 216 -25786
rect 358 -25786 374 -25769
rect 498 -25769 556 -25752
rect 614 -25752 854 -25714
rect 614 -25769 672 -25752
rect 498 -25786 514 -25769
rect 358 -25802 514 -25786
rect 656 -25786 672 -25769
rect 796 -25769 854 -25752
rect 796 -25786 812 -25769
rect 656 -25802 812 -25786
rect 2626 -25922 3586 -25884
rect 2626 -25939 2828 -25922
rect 2812 -25956 2828 -25939
rect 3384 -25939 3586 -25922
rect 3644 -25922 4604 -25884
rect 3644 -25939 3846 -25922
rect 3384 -25956 3400 -25939
rect 2812 -25972 3400 -25956
rect 3830 -25956 3846 -25939
rect 4402 -25939 4604 -25922
rect 4662 -25922 5622 -25884
rect 4662 -25939 4864 -25922
rect 4402 -25956 4418 -25939
rect 3830 -25972 4418 -25956
rect 4848 -25956 4864 -25939
rect 5420 -25939 5622 -25922
rect 5680 -25922 6640 -25884
rect 5680 -25939 5882 -25922
rect 5420 -25956 5436 -25939
rect 4848 -25972 5436 -25956
rect 5866 -25956 5882 -25939
rect 6438 -25939 6640 -25922
rect 6698 -25922 7658 -25884
rect 6698 -25939 6900 -25922
rect 6438 -25956 6454 -25939
rect 5866 -25972 6454 -25956
rect 6884 -25956 6900 -25939
rect 7456 -25939 7658 -25922
rect 7716 -25922 8676 -25884
rect 7716 -25939 7918 -25922
rect 7456 -25956 7472 -25939
rect 6884 -25972 7472 -25956
rect 7902 -25956 7918 -25939
rect 8474 -25939 8676 -25922
rect 8734 -25922 9694 -25884
rect 8734 -25939 8936 -25922
rect 8474 -25956 8490 -25939
rect 7902 -25972 8490 -25956
rect 8920 -25956 8936 -25939
rect 9492 -25939 9694 -25922
rect 9752 -25922 10712 -25884
rect 9752 -25939 9954 -25922
rect 9492 -25956 9508 -25939
rect 8920 -25972 9508 -25956
rect 9938 -25956 9954 -25939
rect 10510 -25939 10712 -25922
rect 10770 -25922 11730 -25884
rect 10770 -25939 10972 -25922
rect 10510 -25956 10526 -25939
rect 9938 -25972 10526 -25956
rect 10956 -25956 10972 -25939
rect 11528 -25939 11730 -25922
rect 11788 -25922 12748 -25884
rect 11788 -25939 11990 -25922
rect 11528 -25956 11544 -25939
rect 10956 -25972 11544 -25956
rect 11974 -25956 11990 -25939
rect 12546 -25939 12748 -25922
rect 12806 -25922 13766 -25884
rect 12806 -25939 13008 -25922
rect 12546 -25956 12562 -25939
rect 11974 -25972 12562 -25956
rect 12992 -25956 13008 -25939
rect 13564 -25939 13766 -25922
rect 13824 -25922 14784 -25884
rect 13824 -25939 14026 -25922
rect 13564 -25956 13580 -25939
rect 12992 -25972 13580 -25956
rect 14010 -25956 14026 -25939
rect 14582 -25939 14784 -25922
rect 14842 -25922 15802 -25884
rect 14842 -25939 15044 -25922
rect 14582 -25956 14598 -25939
rect 14010 -25972 14598 -25956
rect 15028 -25956 15044 -25939
rect 15600 -25939 15802 -25922
rect 15860 -25922 16820 -25884
rect 15860 -25939 16062 -25922
rect 15600 -25956 15616 -25939
rect 15028 -25972 15616 -25956
rect 16046 -25956 16062 -25939
rect 16618 -25939 16820 -25922
rect 16878 -25922 17838 -25884
rect 16878 -25939 17080 -25922
rect 16618 -25956 16634 -25939
rect 16046 -25972 16634 -25956
rect 17064 -25956 17080 -25939
rect 17636 -25939 17838 -25922
rect 17896 -25922 18856 -25884
rect 17896 -25939 18098 -25922
rect 17636 -25956 17652 -25939
rect 17064 -25972 17652 -25956
rect 18082 -25956 18098 -25939
rect 18654 -25939 18856 -25922
rect 18914 -25922 19874 -25884
rect 18914 -25939 19116 -25922
rect 18654 -25956 18670 -25939
rect 18082 -25972 18670 -25956
rect 19100 -25956 19116 -25939
rect 19672 -25939 19874 -25922
rect 19932 -25922 20892 -25884
rect 19932 -25939 20134 -25922
rect 19672 -25956 19688 -25939
rect 19100 -25972 19688 -25956
rect 20118 -25956 20134 -25939
rect 20690 -25939 20892 -25922
rect 20950 -25922 21910 -25884
rect 20950 -25939 21152 -25922
rect 20690 -25956 20706 -25939
rect 20118 -25972 20706 -25956
rect 21136 -25956 21152 -25939
rect 21708 -25939 21910 -25922
rect 21968 -25922 22928 -25884
rect 21968 -25939 22170 -25922
rect 21708 -25956 21724 -25939
rect 21136 -25972 21724 -25956
rect 22154 -25956 22170 -25939
rect 22726 -25939 22928 -25922
rect 22726 -25956 22742 -25939
rect 22154 -25972 22742 -25956
<< polycont >>
rect 3714 -4643 3790 -4609
rect 3932 -4643 4008 -4609
rect 4150 -4643 4226 -4609
rect 4368 -4643 4444 -4609
rect 4586 -4643 4662 -4609
rect 4804 -4643 4880 -4609
rect 5022 -4643 5098 -4609
rect 5240 -4643 5316 -4609
rect 5458 -4643 5534 -4609
rect 5676 -4643 5752 -4609
rect 3714 -5171 3790 -5137
rect 3932 -5171 4008 -5137
rect 4150 -5171 4226 -5137
rect 4368 -5171 4444 -5137
rect 4586 -5171 4662 -5137
rect 4804 -5171 4880 -5137
rect 5022 -5171 5098 -5137
rect 5240 -5171 5316 -5137
rect 5458 -5171 5534 -5137
rect 5676 -5171 5752 -5137
rect 3714 -5581 3790 -5547
rect 3932 -5581 4008 -5547
rect 4150 -5581 4226 -5547
rect 4368 -5581 4444 -5547
rect 4586 -5581 4662 -5547
rect 4804 -5581 4880 -5547
rect 5022 -5581 5098 -5547
rect 5240 -5581 5316 -5547
rect 5458 -5581 5534 -5547
rect 5676 -5581 5752 -5547
rect 3714 -6109 3790 -6075
rect 3932 -6109 4008 -6075
rect 4150 -6109 4226 -6075
rect 4368 -6109 4444 -6075
rect 4586 -6109 4662 -6075
rect 4804 -6109 4880 -6075
rect 5022 -6109 5098 -6075
rect 5240 -6109 5316 -6075
rect 5458 -6109 5534 -6075
rect 5676 -6109 5752 -6075
rect 3714 -6519 3790 -6485
rect 3932 -6519 4008 -6485
rect 4150 -6519 4226 -6485
rect 4368 -6519 4444 -6485
rect 4586 -6519 4662 -6485
rect 4804 -6519 4880 -6485
rect 5022 -6519 5098 -6485
rect 5240 -6519 5316 -6485
rect 5458 -6519 5534 -6485
rect 5676 -6519 5752 -6485
rect 3714 -7047 3790 -7013
rect 3932 -7047 4008 -7013
rect 4150 -7047 4226 -7013
rect 4368 -7047 4444 -7013
rect 4586 -7047 4662 -7013
rect 4804 -7047 4880 -7013
rect 5022 -7047 5098 -7013
rect 5240 -7047 5316 -7013
rect 5458 -7047 5534 -7013
rect 5676 -7047 5752 -7013
rect 3714 -7457 3790 -7423
rect 3932 -7457 4008 -7423
rect 4150 -7457 4226 -7423
rect 4368 -7457 4444 -7423
rect 4586 -7457 4662 -7423
rect 4804 -7457 4880 -7423
rect 5022 -7457 5098 -7423
rect 5240 -7457 5316 -7423
rect 5458 -7457 5534 -7423
rect 5676 -7457 5752 -7423
rect 3714 -7985 3790 -7951
rect 3932 -7985 4008 -7951
rect 4150 -7985 4226 -7951
rect 4368 -7985 4444 -7951
rect 4586 -7985 4662 -7951
rect 4804 -7985 4880 -7951
rect 5022 -7985 5098 -7951
rect 5240 -7985 5316 -7951
rect 5458 -7985 5534 -7951
rect 5676 -7985 5752 -7951
rect 2830 -11680 3386 -11646
rect 3848 -11680 4404 -11646
rect 4866 -11680 5422 -11646
rect 5884 -11680 6440 -11646
rect 6902 -11680 7458 -11646
rect 7920 -11680 8476 -11646
rect 8938 -11680 9494 -11646
rect 9956 -11680 10512 -11646
rect 10974 -11680 11530 -11646
rect 11992 -11680 12548 -11646
rect 13010 -11680 13566 -11646
rect 14028 -11680 14584 -11646
rect 15046 -11680 15602 -11646
rect 16064 -11680 16620 -11646
rect 17082 -11680 17638 -11646
rect 18100 -11680 18656 -11646
rect 19118 -11680 19674 -11646
rect 20136 -11680 20692 -11646
rect 21154 -11680 21710 -11646
rect 22172 -11680 22728 -11646
rect 2830 -12390 3386 -12356
rect 3848 -12390 4404 -12356
rect 4866 -12390 5422 -12356
rect 5884 -12390 6440 -12356
rect 6902 -12390 7458 -12356
rect 7920 -12390 8476 -12356
rect 8938 -12390 9494 -12356
rect 9956 -12390 10512 -12356
rect 10974 -12390 11530 -12356
rect 11992 -12390 12548 -12356
rect 13010 -12390 13566 -12356
rect 14028 -12390 14584 -12356
rect 15046 -12390 15602 -12356
rect 16064 -12390 16620 -12356
rect 17082 -12390 17638 -12356
rect 18100 -12390 18656 -12356
rect 19118 -12390 19674 -12356
rect 20136 -12390 20692 -12356
rect 21154 -12390 21710 -12356
rect 22172 -12390 22728 -12356
rect -8936 -12474 -8380 -12440
rect -7918 -12474 -7362 -12440
rect -6900 -12474 -6344 -12440
rect -5882 -12474 -5326 -12440
rect -4864 -12474 -4308 -12440
rect -3846 -12474 -3290 -12440
rect -2828 -12474 -2272 -12440
rect -1810 -12474 -1254 -12440
rect -792 -12474 -236 -12440
rect 2830 -12914 3386 -12880
rect 3848 -12914 4404 -12880
rect 4866 -12914 5422 -12880
rect 5884 -12914 6440 -12880
rect 6902 -12914 7458 -12880
rect 7920 -12914 8476 -12880
rect 8938 -12914 9494 -12880
rect 9956 -12914 10512 -12880
rect 10974 -12914 11530 -12880
rect 11992 -12914 12548 -12880
rect 13010 -12914 13566 -12880
rect 14028 -12914 14584 -12880
rect 15046 -12914 15602 -12880
rect 16064 -12914 16620 -12880
rect 17082 -12914 17638 -12880
rect 18100 -12914 18656 -12880
rect 19118 -12914 19674 -12880
rect 20136 -12914 20692 -12880
rect 21154 -12914 21710 -12880
rect 22172 -12914 22728 -12880
rect -8936 -13184 -8380 -13150
rect -7918 -13184 -7362 -13150
rect -6900 -13184 -6344 -13150
rect -5882 -13184 -5326 -13150
rect -4864 -13184 -4308 -13150
rect -3846 -13184 -3290 -13150
rect -2828 -13184 -2272 -13150
rect -1810 -13184 -1254 -13150
rect -792 -13184 -236 -13150
rect -8936 -13292 -8380 -13258
rect -7918 -13292 -7362 -13258
rect -6900 -13292 -6344 -13258
rect -5882 -13292 -5326 -13258
rect -4864 -13292 -4308 -13258
rect -3846 -13292 -3290 -13258
rect -2828 -13292 -2272 -13258
rect -1810 -13292 -1254 -13258
rect -792 -13292 -236 -13258
rect 2830 -13624 3386 -13590
rect 3848 -13624 4404 -13590
rect 4866 -13624 5422 -13590
rect 5884 -13624 6440 -13590
rect 6902 -13624 7458 -13590
rect 7920 -13624 8476 -13590
rect 8938 -13624 9494 -13590
rect 9956 -13624 10512 -13590
rect 10974 -13624 11530 -13590
rect 11992 -13624 12548 -13590
rect 13010 -13624 13566 -13590
rect 14028 -13624 14584 -13590
rect 15046 -13624 15602 -13590
rect 16064 -13624 16620 -13590
rect 17082 -13624 17638 -13590
rect 18100 -13624 18656 -13590
rect 19118 -13624 19674 -13590
rect 20136 -13624 20692 -13590
rect 21154 -13624 21710 -13590
rect 22172 -13624 22728 -13590
rect -8936 -14002 -8380 -13968
rect -7918 -14002 -7362 -13968
rect -6900 -14002 -6344 -13968
rect -5882 -14002 -5326 -13968
rect -4864 -14002 -4308 -13968
rect -3846 -14002 -3290 -13968
rect -2828 -14002 -2272 -13968
rect -1810 -14002 -1254 -13968
rect -792 -14002 -236 -13968
rect -8936 -14110 -8380 -14076
rect -7918 -14110 -7362 -14076
rect -6900 -14110 -6344 -14076
rect -5882 -14110 -5326 -14076
rect -4864 -14110 -4308 -14076
rect -3846 -14110 -3290 -14076
rect -2828 -14110 -2272 -14076
rect -1810 -14110 -1254 -14076
rect -792 -14110 -236 -14076
rect 2830 -14146 3386 -14112
rect 3848 -14146 4404 -14112
rect 4866 -14146 5422 -14112
rect 5884 -14146 6440 -14112
rect 6902 -14146 7458 -14112
rect 7920 -14146 8476 -14112
rect 8938 -14146 9494 -14112
rect 9956 -14146 10512 -14112
rect 10974 -14146 11530 -14112
rect 11992 -14146 12548 -14112
rect 13010 -14146 13566 -14112
rect 14028 -14146 14584 -14112
rect 15046 -14146 15602 -14112
rect 16064 -14146 16620 -14112
rect 17082 -14146 17638 -14112
rect 18100 -14146 18656 -14112
rect 19118 -14146 19674 -14112
rect 20136 -14146 20692 -14112
rect 21154 -14146 21710 -14112
rect 22172 -14146 22728 -14112
rect -8936 -14820 -8380 -14786
rect -7918 -14820 -7362 -14786
rect -6900 -14820 -6344 -14786
rect -5882 -14820 -5326 -14786
rect -4864 -14820 -4308 -14786
rect -3846 -14820 -3290 -14786
rect -2828 -14820 -2272 -14786
rect -1810 -14820 -1254 -14786
rect -792 -14820 -236 -14786
rect 2830 -14856 3386 -14822
rect 3848 -14856 4404 -14822
rect 4866 -14856 5422 -14822
rect 5884 -14856 6440 -14822
rect 6902 -14856 7458 -14822
rect 7920 -14856 8476 -14822
rect 8938 -14856 9494 -14822
rect 9956 -14856 10512 -14822
rect 10974 -14856 11530 -14822
rect 11992 -14856 12548 -14822
rect 13010 -14856 13566 -14822
rect 14028 -14856 14584 -14822
rect 15046 -14856 15602 -14822
rect 16064 -14856 16620 -14822
rect 17082 -14856 17638 -14822
rect 18100 -14856 18656 -14822
rect 19118 -14856 19674 -14822
rect 20136 -14856 20692 -14822
rect 21154 -14856 21710 -14822
rect 22172 -14856 22728 -14822
rect -8936 -14928 -8380 -14894
rect -7918 -14928 -7362 -14894
rect -6900 -14928 -6344 -14894
rect -5882 -14928 -5326 -14894
rect -4864 -14928 -4308 -14894
rect -3846 -14928 -3290 -14894
rect -2828 -14928 -2272 -14894
rect -1810 -14928 -1254 -14894
rect -792 -14928 -236 -14894
rect 2828 -15380 3384 -15346
rect 3846 -15380 4402 -15346
rect 4864 -15380 5420 -15346
rect 5882 -15380 6438 -15346
rect 6900 -15380 7456 -15346
rect 7918 -15380 8474 -15346
rect 8936 -15380 9492 -15346
rect 9954 -15380 10510 -15346
rect 10972 -15380 11528 -15346
rect 11990 -15380 12546 -15346
rect 13008 -15380 13564 -15346
rect 14026 -15380 14582 -15346
rect 15044 -15380 15600 -15346
rect 16062 -15380 16618 -15346
rect 17080 -15380 17636 -15346
rect 18098 -15380 18654 -15346
rect 19116 -15380 19672 -15346
rect 20134 -15380 20690 -15346
rect 21152 -15380 21708 -15346
rect 22170 -15380 22726 -15346
rect -8936 -15638 -8380 -15604
rect -7918 -15638 -7362 -15604
rect -6900 -15638 -6344 -15604
rect -5882 -15638 -5326 -15604
rect -4864 -15638 -4308 -15604
rect -3846 -15638 -3290 -15604
rect -2828 -15638 -2272 -15604
rect -1810 -15638 -1254 -15604
rect -792 -15638 -236 -15604
rect -8936 -15746 -8380 -15712
rect -7918 -15746 -7362 -15712
rect -6900 -15746 -6344 -15712
rect -5882 -15746 -5326 -15712
rect -4864 -15746 -4308 -15712
rect -3846 -15746 -3290 -15712
rect -2828 -15746 -2272 -15712
rect -1810 -15746 -1254 -15712
rect -792 -15746 -236 -15712
rect 2828 -16090 3384 -16056
rect 3846 -16090 4402 -16056
rect 4864 -16090 5420 -16056
rect 5882 -16090 6438 -16056
rect 6900 -16090 7456 -16056
rect 7918 -16090 8474 -16056
rect 8936 -16090 9492 -16056
rect 9954 -16090 10510 -16056
rect 10972 -16090 11528 -16056
rect 11990 -16090 12546 -16056
rect 13008 -16090 13564 -16056
rect 14026 -16090 14582 -16056
rect 15044 -16090 15600 -16056
rect 16062 -16090 16618 -16056
rect 17080 -16090 17636 -16056
rect 18098 -16090 18654 -16056
rect 19116 -16090 19672 -16056
rect 20134 -16090 20690 -16056
rect 21152 -16090 21708 -16056
rect 22170 -16090 22726 -16056
rect -8936 -16456 -8380 -16422
rect -7918 -16456 -7362 -16422
rect -6900 -16456 -6344 -16422
rect -5882 -16456 -5326 -16422
rect -4864 -16456 -4308 -16422
rect -3846 -16456 -3290 -16422
rect -2828 -16456 -2272 -16422
rect -1810 -16456 -1254 -16422
rect -792 -16456 -236 -16422
rect -8936 -16564 -8380 -16530
rect -7918 -16564 -7362 -16530
rect -6900 -16564 -6344 -16530
rect -5882 -16564 -5326 -16530
rect -4864 -16564 -4308 -16530
rect -3846 -16564 -3290 -16530
rect -2828 -16564 -2272 -16530
rect -1810 -16564 -1254 -16530
rect -792 -16564 -236 -16530
rect 2828 -16614 3384 -16580
rect 3846 -16614 4402 -16580
rect 4864 -16614 5420 -16580
rect 5882 -16614 6438 -16580
rect 6900 -16614 7456 -16580
rect 7918 -16614 8474 -16580
rect 8936 -16614 9492 -16580
rect 9954 -16614 10510 -16580
rect 10972 -16614 11528 -16580
rect 11990 -16614 12546 -16580
rect 13008 -16614 13564 -16580
rect 14026 -16614 14582 -16580
rect 15044 -16614 15600 -16580
rect 16062 -16614 16618 -16580
rect 17080 -16614 17636 -16580
rect 18098 -16614 18654 -16580
rect 19116 -16614 19672 -16580
rect 20134 -16614 20690 -16580
rect 21152 -16614 21708 -16580
rect 22170 -16614 22726 -16580
rect -8936 -17274 -8380 -17240
rect -7918 -17274 -7362 -17240
rect -6900 -17274 -6344 -17240
rect -5882 -17274 -5326 -17240
rect -4864 -17274 -4308 -17240
rect -3846 -17274 -3290 -17240
rect -2828 -17274 -2272 -17240
rect -1810 -17274 -1254 -17240
rect -792 -17274 -236 -17240
rect 2828 -17324 3384 -17290
rect -8936 -17382 -8380 -17348
rect -7918 -17382 -7362 -17348
rect -6900 -17382 -6344 -17348
rect -5882 -17382 -5326 -17348
rect -4864 -17382 -4308 -17348
rect -3846 -17382 -3290 -17348
rect -2828 -17382 -2272 -17348
rect -1810 -17382 -1254 -17348
rect 3846 -17324 4402 -17290
rect 4864 -17324 5420 -17290
rect 5882 -17324 6438 -17290
rect 6900 -17324 7456 -17290
rect 7918 -17324 8474 -17290
rect 8936 -17324 9492 -17290
rect 9954 -17324 10510 -17290
rect 10972 -17324 11528 -17290
rect 11990 -17324 12546 -17290
rect 13008 -17324 13564 -17290
rect 14026 -17324 14582 -17290
rect 15044 -17324 15600 -17290
rect 16062 -17324 16618 -17290
rect 17080 -17324 17636 -17290
rect 18098 -17324 18654 -17290
rect 19116 -17324 19672 -17290
rect 20134 -17324 20690 -17290
rect 21152 -17324 21708 -17290
rect 22170 -17324 22726 -17290
rect -792 -17382 -236 -17348
rect 2828 -17846 3384 -17812
rect 3846 -17846 4402 -17812
rect 4864 -17846 5420 -17812
rect 5882 -17846 6438 -17812
rect 6900 -17846 7456 -17812
rect 7918 -17846 8474 -17812
rect 8936 -17846 9492 -17812
rect 9954 -17846 10510 -17812
rect 10972 -17846 11528 -17812
rect 11990 -17846 12546 -17812
rect 13008 -17846 13564 -17812
rect 14026 -17846 14582 -17812
rect 15044 -17846 15600 -17812
rect 16062 -17846 16618 -17812
rect 17080 -17846 17636 -17812
rect 18098 -17846 18654 -17812
rect 19116 -17846 19672 -17812
rect 20134 -17846 20690 -17812
rect 21152 -17846 21708 -17812
rect 22170 -17846 22726 -17812
rect -8936 -18092 -8380 -18058
rect -7918 -18092 -7362 -18058
rect -6900 -18092 -6344 -18058
rect -5882 -18092 -5326 -18058
rect -4864 -18092 -4308 -18058
rect -3846 -18092 -3290 -18058
rect -2828 -18092 -2272 -18058
rect -1810 -18092 -1254 -18058
rect -792 -18092 -236 -18058
rect -8936 -18200 -8380 -18166
rect -7918 -18200 -7362 -18166
rect -6900 -18200 -6344 -18166
rect -5882 -18200 -5326 -18166
rect -4864 -18200 -4308 -18166
rect -3846 -18200 -3290 -18166
rect -2828 -18200 -2272 -18166
rect -1810 -18200 -1254 -18166
rect -792 -18200 -236 -18166
rect 2828 -18556 3384 -18522
rect 3846 -18556 4402 -18522
rect 4864 -18556 5420 -18522
rect 5882 -18556 6438 -18522
rect 6900 -18556 7456 -18522
rect 7918 -18556 8474 -18522
rect 8936 -18556 9492 -18522
rect 9954 -18556 10510 -18522
rect 10972 -18556 11528 -18522
rect 11990 -18556 12546 -18522
rect 13008 -18556 13564 -18522
rect 14026 -18556 14582 -18522
rect 15044 -18556 15600 -18522
rect 16062 -18556 16618 -18522
rect 17080 -18556 17636 -18522
rect 18098 -18556 18654 -18522
rect 19116 -18556 19672 -18522
rect 20134 -18556 20690 -18522
rect 21152 -18556 21708 -18522
rect 22170 -18556 22726 -18522
rect -8936 -18910 -8380 -18876
rect -7918 -18910 -7362 -18876
rect -6900 -18910 -6344 -18876
rect -5882 -18910 -5326 -18876
rect -4864 -18910 -4308 -18876
rect -3846 -18910 -3290 -18876
rect -2828 -18910 -2272 -18876
rect -1810 -18910 -1254 -18876
rect -792 -18910 -236 -18876
rect 2828 -19080 3384 -19046
rect 3846 -19080 4402 -19046
rect 4864 -19080 5420 -19046
rect 5882 -19080 6438 -19046
rect 6900 -19080 7456 -19046
rect 7918 -19080 8474 -19046
rect 8936 -19080 9492 -19046
rect 9954 -19080 10510 -19046
rect 10972 -19080 11528 -19046
rect 11990 -19080 12546 -19046
rect 13008 -19080 13564 -19046
rect 14026 -19080 14582 -19046
rect 15044 -19080 15600 -19046
rect 16062 -19080 16618 -19046
rect 17080 -19080 17636 -19046
rect 18098 -19080 18654 -19046
rect 19116 -19080 19672 -19046
rect 20134 -19080 20690 -19046
rect 21152 -19080 21708 -19046
rect 22170 -19080 22726 -19046
rect -2236 -19584 -2160 -19550
rect -2018 -19584 -1942 -19550
rect -1800 -19584 -1724 -19550
rect -1582 -19584 -1506 -19550
rect -1364 -19584 -1288 -19550
rect -1146 -19584 -1070 -19550
rect -928 -19584 -852 -19550
rect -710 -19584 -634 -19550
rect -492 -19584 -416 -19550
rect -274 -19584 -198 -19550
rect 2828 -19790 3384 -19756
rect 3846 -19790 4402 -19756
rect 4864 -19790 5420 -19756
rect 5882 -19790 6438 -19756
rect 6900 -19790 7456 -19756
rect 7918 -19790 8474 -19756
rect 8936 -19790 9492 -19756
rect 9954 -19790 10510 -19756
rect 10972 -19790 11528 -19756
rect 11990 -19790 12546 -19756
rect 13008 -19790 13564 -19756
rect 14026 -19790 14582 -19756
rect 15044 -19790 15600 -19756
rect 16062 -19790 16618 -19756
rect 17080 -19790 17636 -19756
rect 18098 -19790 18654 -19756
rect 19116 -19790 19672 -19756
rect 20134 -19790 20690 -19756
rect 21152 -19790 21708 -19756
rect 22170 -19790 22726 -19756
rect -2236 -19894 -2160 -19860
rect -2018 -19894 -1942 -19860
rect -1800 -19894 -1724 -19860
rect -1582 -19894 -1506 -19860
rect -1364 -19894 -1288 -19860
rect -1146 -19894 -1070 -19860
rect -928 -19894 -852 -19860
rect -710 -19894 -634 -19860
rect -492 -19894 -416 -19860
rect -274 -19894 -198 -19860
rect 2828 -20314 3384 -20280
rect 3846 -20314 4402 -20280
rect 4864 -20314 5420 -20280
rect 5882 -20314 6438 -20280
rect 6900 -20314 7456 -20280
rect 7918 -20314 8474 -20280
rect 8936 -20314 9492 -20280
rect 9954 -20314 10510 -20280
rect 10972 -20314 11528 -20280
rect 11990 -20314 12546 -20280
rect 13008 -20314 13564 -20280
rect 14026 -20314 14582 -20280
rect 15044 -20314 15600 -20280
rect 16062 -20314 16618 -20280
rect 17080 -20314 17636 -20280
rect 18098 -20314 18654 -20280
rect 19116 -20314 19672 -20280
rect 20134 -20314 20690 -20280
rect 21152 -20314 21708 -20280
rect 22170 -20314 22726 -20280
rect -2236 -20416 -2160 -20382
rect -2018 -20416 -1942 -20382
rect -1800 -20416 -1724 -20382
rect -1582 -20416 -1506 -20382
rect -1364 -20416 -1288 -20382
rect -1146 -20416 -1070 -20382
rect -928 -20416 -852 -20382
rect -710 -20416 -634 -20382
rect -492 -20416 -416 -20382
rect -274 -20416 -198 -20382
rect -2236 -20726 -2160 -20692
rect -2018 -20726 -1942 -20692
rect -1800 -20726 -1724 -20692
rect -1582 -20726 -1506 -20692
rect -1364 -20726 -1288 -20692
rect -1146 -20726 -1070 -20692
rect -928 -20726 -852 -20692
rect -710 -20726 -634 -20692
rect -492 -20726 -416 -20692
rect -274 -20726 -198 -20692
rect 2828 -21024 3384 -20990
rect 3846 -21024 4402 -20990
rect 4864 -21024 5420 -20990
rect 5882 -21024 6438 -20990
rect 6900 -21024 7456 -20990
rect 7918 -21024 8474 -20990
rect 8936 -21024 9492 -20990
rect 9954 -21024 10510 -20990
rect 10972 -21024 11528 -20990
rect 11990 -21024 12546 -20990
rect 13008 -21024 13564 -20990
rect 14026 -21024 14582 -20990
rect 15044 -21024 15600 -20990
rect 16062 -21024 16618 -20990
rect 17080 -21024 17636 -20990
rect 18098 -21024 18654 -20990
rect 19116 -21024 19672 -20990
rect 20134 -21024 20690 -20990
rect 21152 -21024 21708 -20990
rect 22170 -21024 22726 -20990
rect 2828 -21546 3384 -21512
rect 3846 -21546 4402 -21512
rect 4864 -21546 5420 -21512
rect 5882 -21546 6438 -21512
rect 6900 -21546 7456 -21512
rect 7918 -21546 8474 -21512
rect 8936 -21546 9492 -21512
rect 9954 -21546 10510 -21512
rect 10972 -21546 11528 -21512
rect 11990 -21546 12546 -21512
rect 13008 -21546 13564 -21512
rect 14026 -21546 14582 -21512
rect 15044 -21546 15600 -21512
rect 16062 -21546 16618 -21512
rect 17080 -21546 17636 -21512
rect 18098 -21546 18654 -21512
rect 19116 -21546 19672 -21512
rect 20134 -21546 20690 -21512
rect 21152 -21546 21708 -21512
rect 22170 -21546 22726 -21512
rect -9157 -21743 -8601 -21709
rect -8139 -21743 -7583 -21709
rect -7121 -21743 -6565 -21709
rect -6103 -21743 -5547 -21709
rect -5085 -21743 -4529 -21709
rect -4067 -21743 -3511 -21709
rect -2306 -21742 -2182 -21708
rect -2008 -21742 -1884 -21708
rect -1710 -21742 -1586 -21708
rect -1412 -21742 -1288 -21708
rect -1114 -21742 -990 -21708
rect -816 -21742 -692 -21708
rect -518 -21742 -394 -21708
rect -220 -21742 -96 -21708
rect 78 -21742 202 -21708
rect 376 -21742 500 -21708
rect 674 -21742 798 -21708
rect 2828 -22256 3384 -22222
rect 3846 -22256 4402 -22222
rect 4864 -22256 5420 -22222
rect 5882 -22256 6438 -22222
rect 6900 -22256 7456 -22222
rect 7918 -22256 8474 -22222
rect 8936 -22256 9492 -22222
rect 9954 -22256 10510 -22222
rect 10972 -22256 11528 -22222
rect 11990 -22256 12546 -22222
rect 13008 -22256 13564 -22222
rect 14026 -22256 14582 -22222
rect 15044 -22256 15600 -22222
rect 16062 -22256 16618 -22222
rect 17080 -22256 17636 -22222
rect 18098 -22256 18654 -22222
rect 19116 -22256 19672 -22222
rect 20134 -22256 20690 -22222
rect 21152 -22256 21708 -22222
rect 22170 -22256 22726 -22222
rect -9157 -22453 -8601 -22419
rect -8139 -22453 -7583 -22419
rect -7121 -22453 -6565 -22419
rect -6103 -22453 -5547 -22419
rect -5085 -22453 -4529 -22419
rect -4067 -22453 -3511 -22419
rect -2306 -22452 -2182 -22418
rect -2008 -22452 -1884 -22418
rect -1710 -22452 -1586 -22418
rect -1412 -22452 -1288 -22418
rect -1114 -22452 -990 -22418
rect -816 -22452 -692 -22418
rect -518 -22452 -394 -22418
rect -220 -22452 -96 -22418
rect 78 -22452 202 -22418
rect 376 -22452 500 -22418
rect 674 -22452 798 -22418
rect 2828 -22780 3384 -22746
rect -9158 -22856 -8602 -22822
rect -8140 -22856 -7584 -22822
rect -7122 -22856 -6566 -22822
rect -6104 -22856 -5548 -22822
rect -5086 -22856 -4530 -22822
rect -4068 -22856 -3512 -22822
rect -2306 -22854 -2182 -22820
rect -2008 -22854 -1884 -22820
rect -1710 -22854 -1586 -22820
rect -1412 -22854 -1288 -22820
rect -1114 -22854 -990 -22820
rect -816 -22854 -692 -22820
rect -518 -22854 -394 -22820
rect -220 -22854 -96 -22820
rect 78 -22854 202 -22820
rect 376 -22854 500 -22820
rect 3846 -22780 4402 -22746
rect 4864 -22780 5420 -22746
rect 5882 -22780 6438 -22746
rect 6900 -22780 7456 -22746
rect 7918 -22780 8474 -22746
rect 8936 -22780 9492 -22746
rect 9954 -22780 10510 -22746
rect 10972 -22780 11528 -22746
rect 11990 -22780 12546 -22746
rect 13008 -22780 13564 -22746
rect 14026 -22780 14582 -22746
rect 15044 -22780 15600 -22746
rect 16062 -22780 16618 -22746
rect 17080 -22780 17636 -22746
rect 18098 -22780 18654 -22746
rect 19116 -22780 19672 -22746
rect 20134 -22780 20690 -22746
rect 21152 -22780 21708 -22746
rect 22170 -22780 22726 -22746
rect 674 -22854 798 -22820
rect 2828 -23490 3384 -23456
rect -9158 -23566 -8602 -23532
rect -8140 -23566 -7584 -23532
rect -7122 -23566 -6566 -23532
rect -6104 -23566 -5548 -23532
rect -5086 -23566 -4530 -23532
rect -4068 -23566 -3512 -23532
rect -2306 -23564 -2182 -23530
rect -2008 -23564 -1884 -23530
rect -1710 -23564 -1586 -23530
rect -1412 -23564 -1288 -23530
rect -1114 -23564 -990 -23530
rect -816 -23564 -692 -23530
rect -518 -23564 -394 -23530
rect -220 -23564 -96 -23530
rect 78 -23564 202 -23530
rect 376 -23564 500 -23530
rect 3846 -23490 4402 -23456
rect 4864 -23490 5420 -23456
rect 5882 -23490 6438 -23456
rect 6900 -23490 7456 -23456
rect 7918 -23490 8474 -23456
rect 8936 -23490 9492 -23456
rect 9954 -23490 10510 -23456
rect 10972 -23490 11528 -23456
rect 11990 -23490 12546 -23456
rect 13008 -23490 13564 -23456
rect 14026 -23490 14582 -23456
rect 15044 -23490 15600 -23456
rect 16062 -23490 16618 -23456
rect 17080 -23490 17636 -23456
rect 18098 -23490 18654 -23456
rect 19116 -23490 19672 -23456
rect 20134 -23490 20690 -23456
rect 21152 -23490 21708 -23456
rect 22170 -23490 22726 -23456
rect 674 -23564 798 -23530
rect -9157 -23967 -8601 -23933
rect -8139 -23967 -7583 -23933
rect -7121 -23967 -6565 -23933
rect -6103 -23967 -5547 -23933
rect -5085 -23967 -4529 -23933
rect -4067 -23967 -3511 -23933
rect -2308 -23966 -2184 -23932
rect -2010 -23966 -1886 -23932
rect -1712 -23966 -1588 -23932
rect -1414 -23966 -1290 -23932
rect -1116 -23966 -992 -23932
rect -818 -23966 -694 -23932
rect -520 -23966 -396 -23932
rect -222 -23966 -98 -23932
rect 76 -23966 200 -23932
rect 374 -23966 498 -23932
rect 672 -23966 796 -23932
rect 2828 -24014 3384 -23980
rect 3846 -24014 4402 -23980
rect 4864 -24014 5420 -23980
rect 5882 -24014 6438 -23980
rect 6900 -24014 7456 -23980
rect 7918 -24014 8474 -23980
rect 8936 -24014 9492 -23980
rect 9954 -24014 10510 -23980
rect 10972 -24014 11528 -23980
rect 11990 -24014 12546 -23980
rect 13008 -24014 13564 -23980
rect 14026 -24014 14582 -23980
rect 15044 -24014 15600 -23980
rect 16062 -24014 16618 -23980
rect 17080 -24014 17636 -23980
rect 18098 -24014 18654 -23980
rect 19116 -24014 19672 -23980
rect 20134 -24014 20690 -23980
rect 21152 -24014 21708 -23980
rect 22170 -24014 22726 -23980
rect -9157 -24677 -8601 -24643
rect -8139 -24677 -7583 -24643
rect -7121 -24677 -6565 -24643
rect -6103 -24677 -5547 -24643
rect -5085 -24677 -4529 -24643
rect -4067 -24677 -3511 -24643
rect -2308 -24676 -2184 -24642
rect -2010 -24676 -1886 -24642
rect -1712 -24676 -1588 -24642
rect -1414 -24676 -1290 -24642
rect -1116 -24676 -992 -24642
rect -818 -24676 -694 -24642
rect -520 -24676 -396 -24642
rect -222 -24676 -98 -24642
rect 76 -24676 200 -24642
rect 374 -24676 498 -24642
rect 672 -24676 796 -24642
rect 2828 -24724 3384 -24690
rect 3846 -24724 4402 -24690
rect 4864 -24724 5420 -24690
rect 5882 -24724 6438 -24690
rect 6900 -24724 7456 -24690
rect 7918 -24724 8474 -24690
rect 8936 -24724 9492 -24690
rect 9954 -24724 10510 -24690
rect 10972 -24724 11528 -24690
rect 11990 -24724 12546 -24690
rect 13008 -24724 13564 -24690
rect 14026 -24724 14582 -24690
rect 15044 -24724 15600 -24690
rect 16062 -24724 16618 -24690
rect 17080 -24724 17636 -24690
rect 18098 -24724 18654 -24690
rect 19116 -24724 19672 -24690
rect 20134 -24724 20690 -24690
rect 21152 -24724 21708 -24690
rect 22170 -24724 22726 -24690
rect -9158 -25080 -8602 -25046
rect -8140 -25080 -7584 -25046
rect -7122 -25080 -6566 -25046
rect -6104 -25080 -5548 -25046
rect -5086 -25080 -4530 -25046
rect -4068 -25080 -3512 -25046
rect -2308 -25076 -2184 -25042
rect -2010 -25076 -1886 -25042
rect -1712 -25076 -1588 -25042
rect -1414 -25076 -1290 -25042
rect -1116 -25076 -992 -25042
rect -818 -25076 -694 -25042
rect -520 -25076 -396 -25042
rect -222 -25076 -98 -25042
rect 76 -25076 200 -25042
rect 374 -25076 498 -25042
rect 672 -25076 796 -25042
rect 2828 -25246 3384 -25212
rect 3846 -25246 4402 -25212
rect 4864 -25246 5420 -25212
rect 5882 -25246 6438 -25212
rect 6900 -25246 7456 -25212
rect 7918 -25246 8474 -25212
rect 8936 -25246 9492 -25212
rect 9954 -25246 10510 -25212
rect 10972 -25246 11528 -25212
rect 11990 -25246 12546 -25212
rect 13008 -25246 13564 -25212
rect 14026 -25246 14582 -25212
rect 15044 -25246 15600 -25212
rect 16062 -25246 16618 -25212
rect 17080 -25246 17636 -25212
rect 18098 -25246 18654 -25212
rect 19116 -25246 19672 -25212
rect 20134 -25246 20690 -25212
rect 21152 -25246 21708 -25212
rect 22170 -25246 22726 -25212
rect -9158 -25790 -8602 -25756
rect -8140 -25790 -7584 -25756
rect -7122 -25790 -6566 -25756
rect -6104 -25790 -5548 -25756
rect -5086 -25790 -4530 -25756
rect -4068 -25790 -3512 -25756
rect -2308 -25786 -2184 -25752
rect -2010 -25786 -1886 -25752
rect -1712 -25786 -1588 -25752
rect -1414 -25786 -1290 -25752
rect -1116 -25786 -992 -25752
rect -818 -25786 -694 -25752
rect -520 -25786 -396 -25752
rect -222 -25786 -98 -25752
rect 76 -25786 200 -25752
rect 374 -25786 498 -25752
rect 672 -25786 796 -25752
rect 2828 -25956 3384 -25922
rect 3846 -25956 4402 -25922
rect 4864 -25956 5420 -25922
rect 5882 -25956 6438 -25922
rect 6900 -25956 7456 -25922
rect 7918 -25956 8474 -25922
rect 8936 -25956 9492 -25922
rect 9954 -25956 10510 -25922
rect 10972 -25956 11528 -25922
rect 11990 -25956 12546 -25922
rect 13008 -25956 13564 -25922
rect 14026 -25956 14582 -25922
rect 15044 -25956 15600 -25922
rect 16062 -25956 16618 -25922
rect 17080 -25956 17636 -25922
rect 18098 -25956 18654 -25922
rect 19116 -25956 19672 -25922
rect 20134 -25956 20690 -25922
rect 21152 -25956 21708 -25922
rect 22170 -25956 22726 -25922
<< locali >>
rect 378 1560 478 1722
rect 24722 1560 24822 1722
rect 3698 -4643 3714 -4609
rect 3790 -4643 3806 -4609
rect 3916 -4643 3932 -4609
rect 4008 -4643 4024 -4609
rect 4134 -4643 4150 -4609
rect 4226 -4643 4242 -4609
rect 4352 -4643 4368 -4609
rect 4444 -4643 4460 -4609
rect 4570 -4643 4586 -4609
rect 4662 -4643 4678 -4609
rect 4788 -4643 4804 -4609
rect 4880 -4643 4896 -4609
rect 5006 -4643 5022 -4609
rect 5098 -4643 5114 -4609
rect 5224 -4643 5240 -4609
rect 5316 -4643 5332 -4609
rect 5442 -4643 5458 -4609
rect 5534 -4643 5550 -4609
rect 5660 -4643 5676 -4609
rect 5752 -4643 5768 -4609
rect 3626 -4702 3660 -4686
rect 3626 -5094 3660 -5078
rect 3844 -4702 3878 -4686
rect 3844 -5094 3878 -5078
rect 4062 -4702 4096 -4686
rect 4062 -5094 4096 -5078
rect 4280 -4702 4314 -4686
rect 4280 -5094 4314 -5078
rect 4498 -4702 4532 -4686
rect 4498 -5094 4532 -5078
rect 4716 -4702 4750 -4686
rect 4716 -5094 4750 -5078
rect 4934 -4702 4968 -4686
rect 4934 -5094 4968 -5078
rect 5152 -4702 5186 -4686
rect 5152 -5094 5186 -5078
rect 5370 -4702 5404 -4686
rect 5370 -5094 5404 -5078
rect 5588 -4702 5622 -4686
rect 5588 -5094 5622 -5078
rect 5806 -4702 5840 -4686
rect 5806 -5094 5840 -5078
rect 3944 -5137 4004 -5136
rect 3698 -5171 3714 -5137
rect 3790 -5171 3806 -5137
rect 3916 -5171 3932 -5137
rect 4008 -5171 4024 -5137
rect 4134 -5171 4150 -5137
rect 4226 -5171 4242 -5137
rect 4352 -5171 4368 -5137
rect 4444 -5171 4460 -5137
rect 4570 -5171 4586 -5137
rect 4662 -5171 4678 -5137
rect 4788 -5171 4804 -5137
rect 4880 -5171 4896 -5137
rect 5006 -5171 5022 -5137
rect 5098 -5171 5114 -5137
rect 5224 -5171 5240 -5137
rect 5316 -5171 5332 -5137
rect 5442 -5171 5458 -5137
rect 5534 -5171 5550 -5137
rect 5660 -5171 5676 -5137
rect 5752 -5171 5768 -5137
rect 3698 -5581 3714 -5547
rect 3790 -5581 3806 -5547
rect 3916 -5581 3932 -5547
rect 4008 -5581 4024 -5547
rect 4134 -5581 4150 -5547
rect 4226 -5581 4242 -5547
rect 4352 -5581 4368 -5547
rect 4444 -5581 4460 -5547
rect 4570 -5581 4586 -5547
rect 4662 -5581 4678 -5547
rect 4788 -5581 4804 -5547
rect 4880 -5581 4896 -5547
rect 5006 -5581 5022 -5547
rect 5098 -5581 5114 -5547
rect 5224 -5581 5240 -5547
rect 5316 -5581 5332 -5547
rect 5442 -5581 5458 -5547
rect 5534 -5581 5550 -5547
rect 5660 -5581 5676 -5547
rect 5752 -5581 5768 -5547
rect 3626 -5640 3660 -5624
rect 3626 -6032 3660 -6016
rect 3844 -5640 3878 -5624
rect 3844 -6032 3878 -6016
rect 4062 -5640 4096 -5624
rect 4062 -6032 4096 -6016
rect 4280 -5640 4314 -5624
rect 4280 -6032 4314 -6016
rect 4498 -5640 4532 -5624
rect 4498 -6032 4532 -6016
rect 4716 -5640 4750 -5624
rect 4716 -6032 4750 -6016
rect 4934 -5640 4968 -5624
rect 4934 -6032 4968 -6016
rect 5152 -5640 5186 -5624
rect 5152 -6032 5186 -6016
rect 5370 -5640 5404 -5624
rect 5370 -6032 5404 -6016
rect 5588 -5640 5622 -5624
rect 5588 -6032 5622 -6016
rect 5806 -5640 5840 -5624
rect 5806 -6032 5840 -6016
rect 4376 -6075 4436 -6074
rect 5248 -6075 5308 -6074
rect 3698 -6109 3714 -6075
rect 3790 -6109 3806 -6075
rect 3916 -6109 3932 -6075
rect 4008 -6109 4024 -6075
rect 4134 -6109 4150 -6075
rect 4226 -6109 4242 -6075
rect 4352 -6109 4368 -6075
rect 4444 -6109 4460 -6075
rect 4570 -6109 4586 -6075
rect 4662 -6109 4678 -6075
rect 4788 -6109 4804 -6075
rect 4880 -6109 4896 -6075
rect 5006 -6109 5022 -6075
rect 5098 -6109 5114 -6075
rect 5224 -6109 5240 -6075
rect 5316 -6109 5332 -6075
rect 5442 -6109 5458 -6075
rect 5534 -6109 5550 -6075
rect 5660 -6109 5676 -6075
rect 5752 -6109 5768 -6075
rect 3698 -6519 3714 -6485
rect 3790 -6519 3806 -6485
rect 3916 -6519 3932 -6485
rect 4008 -6519 4024 -6485
rect 4134 -6519 4150 -6485
rect 4226 -6519 4242 -6485
rect 4352 -6519 4368 -6485
rect 4444 -6519 4460 -6485
rect 4570 -6519 4586 -6485
rect 4662 -6519 4678 -6485
rect 4788 -6519 4804 -6485
rect 4880 -6519 4896 -6485
rect 5006 -6519 5022 -6485
rect 5098 -6519 5114 -6485
rect 5224 -6519 5240 -6485
rect 5316 -6519 5332 -6485
rect 5442 -6519 5458 -6485
rect 5534 -6519 5550 -6485
rect 5660 -6519 5676 -6485
rect 5752 -6519 5768 -6485
rect 3938 -6520 3998 -6519
rect 4376 -6520 4436 -6519
rect 3626 -6578 3660 -6562
rect 3626 -6970 3660 -6954
rect 3844 -6578 3878 -6562
rect 3844 -6970 3878 -6954
rect 4062 -6578 4096 -6562
rect 4062 -6970 4096 -6954
rect 4280 -6578 4314 -6562
rect 4280 -6970 4314 -6954
rect 4498 -6578 4532 -6562
rect 4498 -6970 4532 -6954
rect 4716 -6578 4750 -6562
rect 4716 -6970 4750 -6954
rect 4934 -6578 4968 -6562
rect 4934 -6970 4968 -6954
rect 5152 -6578 5186 -6562
rect 5152 -6970 5186 -6954
rect 5370 -6578 5404 -6562
rect 5370 -6970 5404 -6954
rect 5588 -6578 5622 -6562
rect 5588 -6970 5622 -6954
rect 5806 -6578 5840 -6562
rect 5806 -6970 5840 -6954
rect 3698 -7047 3714 -7013
rect 3790 -7047 3806 -7013
rect 3916 -7047 3932 -7013
rect 4008 -7047 4024 -7013
rect 4134 -7047 4150 -7013
rect 4226 -7047 4242 -7013
rect 4352 -7047 4368 -7013
rect 4444 -7047 4460 -7013
rect 4570 -7047 4586 -7013
rect 4662 -7047 4678 -7013
rect 4788 -7047 4804 -7013
rect 4880 -7047 4896 -7013
rect 5006 -7047 5022 -7013
rect 5098 -7047 5114 -7013
rect 5224 -7047 5240 -7013
rect 5316 -7047 5332 -7013
rect 5442 -7047 5458 -7013
rect 5534 -7047 5550 -7013
rect 5660 -7047 5676 -7013
rect 5752 -7047 5768 -7013
rect 3698 -7457 3714 -7423
rect 3790 -7457 3806 -7423
rect 3916 -7457 3932 -7423
rect 4008 -7457 4024 -7423
rect 4134 -7457 4150 -7423
rect 4226 -7457 4242 -7423
rect 4352 -7457 4368 -7423
rect 4444 -7457 4460 -7423
rect 4570 -7457 4586 -7423
rect 4662 -7457 4678 -7423
rect 4788 -7457 4804 -7423
rect 4880 -7457 4896 -7423
rect 5006 -7457 5022 -7423
rect 5098 -7457 5114 -7423
rect 5224 -7457 5240 -7423
rect 5316 -7457 5332 -7423
rect 5442 -7457 5458 -7423
rect 5534 -7457 5550 -7423
rect 5660 -7457 5676 -7423
rect 5752 -7457 5768 -7423
rect 4380 -7458 4440 -7457
rect 3626 -7516 3660 -7500
rect 3626 -7908 3660 -7892
rect 3844 -7516 3878 -7500
rect 3844 -7908 3878 -7892
rect 4062 -7516 4096 -7500
rect 4062 -7908 4096 -7892
rect 4280 -7516 4314 -7500
rect 4280 -7908 4314 -7892
rect 4498 -7516 4532 -7500
rect 4498 -7908 4532 -7892
rect 4716 -7516 4750 -7500
rect 4716 -7908 4750 -7892
rect 4934 -7516 4968 -7500
rect 4934 -7908 4968 -7892
rect 5152 -7516 5186 -7500
rect 5152 -7908 5186 -7892
rect 5370 -7516 5404 -7500
rect 5370 -7908 5404 -7892
rect 5588 -7516 5622 -7500
rect 5588 -7908 5622 -7892
rect 5806 -7516 5840 -7500
rect 5806 -7908 5840 -7892
rect 3698 -7985 3714 -7951
rect 3790 -7985 3806 -7951
rect 3916 -7985 3932 -7951
rect 4008 -7985 4024 -7951
rect 4134 -7985 4150 -7951
rect 4226 -7985 4242 -7951
rect 4352 -7985 4368 -7951
rect 4444 -7985 4460 -7951
rect 4570 -7985 4586 -7951
rect 4662 -7985 4678 -7951
rect 4788 -7985 4804 -7951
rect 4880 -7985 4896 -7951
rect 5006 -7985 5022 -7951
rect 5098 -7985 5114 -7951
rect 5224 -7985 5240 -7951
rect 5316 -7985 5332 -7951
rect 5442 -7985 5458 -7951
rect 5534 -7985 5550 -7951
rect 5660 -7985 5676 -7951
rect 5752 -7985 5768 -7951
rect 378 -8882 478 -8720
rect 24722 -8882 24822 -8720
rect -12322 -11340 -12222 -11178
rect 24822 -11340 24922 -11178
rect 2814 -11680 2830 -11646
rect 3386 -11680 3402 -11646
rect 2582 -11730 2616 -11714
rect 2582 -12322 2616 -12306
rect 3600 -12322 3634 -12306
rect 4618 -12322 4652 -12306
rect 5636 -12322 5670 -12306
rect 6654 -12322 6688 -12306
rect 7672 -12322 7706 -12306
rect 8690 -12322 8724 -12306
rect 9708 -12322 9742 -12306
rect 10726 -12322 10760 -12306
rect 11744 -12322 11778 -12306
rect 12762 -12322 12796 -12306
rect 13780 -12322 13814 -12306
rect 14798 -12322 14832 -12306
rect 15816 -12322 15850 -12306
rect 16834 -12322 16868 -12306
rect 17852 -12322 17886 -12306
rect 18870 -12322 18904 -12306
rect 19888 -12322 19922 -12306
rect 20906 -12322 20940 -12306
rect 21924 -12322 21958 -12306
rect 22942 -12322 22976 -12306
rect 4100 -12356 4160 -12354
rect 5114 -12356 5174 -12348
rect 6118 -12356 6178 -12342
rect 7144 -12356 7204 -12354
rect 8168 -12356 8228 -12348
rect 9188 -12356 9248 -12354
rect 11214 -12356 11274 -12348
rect 12238 -12356 12298 -12354
rect 13248 -12356 13308 -12354
rect 14268 -12356 14328 -12348
rect 15298 -12356 15358 -12354
rect 16302 -12356 16362 -12348
rect 17318 -12356 17378 -12348
rect 18348 -12356 18408 -12354
rect 19362 -12356 19422 -12354
rect 20378 -12356 20438 -12354
rect 21404 -12356 21464 -12354
rect 22426 -12356 22486 -12354
rect 2814 -12390 2830 -12356
rect 3386 -12390 3402 -12356
rect 3832 -12390 3848 -12356
rect 4404 -12390 4420 -12356
rect 4850 -12390 4866 -12356
rect 5422 -12390 5438 -12356
rect 5868 -12390 5884 -12356
rect 6440 -12390 6456 -12356
rect 6886 -12390 6902 -12356
rect 7458 -12390 7474 -12356
rect 7904 -12390 7920 -12356
rect 8476 -12390 8492 -12356
rect 8922 -12390 8938 -12356
rect 9494 -12390 9510 -12356
rect 9940 -12390 9956 -12356
rect 10512 -12390 10528 -12356
rect 10958 -12390 10974 -12356
rect 11530 -12390 11546 -12356
rect 11976 -12390 11992 -12356
rect 12548 -12390 12564 -12356
rect 12994 -12390 13010 -12356
rect 13566 -12390 13582 -12356
rect 14012 -12390 14028 -12356
rect 14584 -12390 14600 -12356
rect 15030 -12390 15046 -12356
rect 15602 -12390 15618 -12356
rect 16048 -12390 16064 -12356
rect 16620 -12390 16636 -12356
rect 17066 -12390 17082 -12356
rect 17638 -12390 17654 -12356
rect 18084 -12390 18100 -12356
rect 18656 -12390 18672 -12356
rect 19102 -12390 19118 -12356
rect 19674 -12390 19690 -12356
rect 20120 -12390 20136 -12356
rect 20692 -12390 20708 -12356
rect 21138 -12390 21154 -12356
rect 21710 -12390 21726 -12356
rect 22156 -12390 22172 -12356
rect 22728 -12390 22744 -12356
rect -8952 -12474 -8936 -12440
rect -8380 -12474 -8364 -12440
rect -7934 -12474 -7918 -12440
rect -7362 -12474 -7346 -12440
rect -6916 -12474 -6900 -12440
rect -6344 -12474 -6328 -12440
rect -5898 -12474 -5882 -12440
rect -5326 -12474 -5310 -12440
rect -4880 -12474 -4864 -12440
rect -4308 -12474 -4292 -12440
rect -3862 -12474 -3846 -12440
rect -3290 -12474 -3274 -12440
rect -2844 -12474 -2828 -12440
rect -2272 -12474 -2256 -12440
rect -1826 -12474 -1810 -12440
rect -1254 -12474 -1238 -12440
rect -808 -12474 -792 -12440
rect -236 -12474 -220 -12440
rect -9184 -12524 -9150 -12508
rect -9184 -13116 -9150 -13100
rect -8166 -12524 -8132 -12508
rect -8166 -13116 -8132 -13100
rect -7148 -12524 -7114 -12508
rect -7148 -13116 -7114 -13100
rect -6130 -12524 -6096 -12508
rect -6130 -13116 -6096 -13100
rect -5112 -12524 -5078 -12508
rect -5112 -13116 -5078 -13100
rect -4094 -12524 -4060 -12508
rect -4094 -13116 -4060 -13100
rect -3076 -12524 -3042 -12508
rect -3076 -13116 -3042 -13100
rect -2058 -12524 -2024 -12508
rect -2058 -13116 -2024 -13100
rect -1040 -12524 -1006 -12508
rect -1040 -13116 -1006 -13100
rect -22 -12524 12 -12508
rect 2814 -12914 2830 -12880
rect 3386 -12914 3402 -12880
rect 3832 -12914 3848 -12880
rect 4404 -12914 4420 -12880
rect 4850 -12914 4866 -12880
rect 5422 -12914 5438 -12880
rect 5868 -12914 5884 -12880
rect 6440 -12914 6456 -12880
rect 6886 -12914 6902 -12880
rect 7458 -12914 7474 -12880
rect 7904 -12914 7920 -12880
rect 8476 -12914 8492 -12880
rect 8922 -12914 8938 -12880
rect 9494 -12914 9510 -12880
rect 9940 -12914 9956 -12880
rect 10512 -12914 10528 -12880
rect 10958 -12914 10974 -12880
rect 11530 -12914 11546 -12880
rect 11976 -12914 11992 -12880
rect 12548 -12914 12564 -12880
rect 12994 -12914 13010 -12880
rect 13566 -12914 13582 -12880
rect 14012 -12914 14028 -12880
rect 14584 -12914 14600 -12880
rect 15030 -12914 15046 -12880
rect 15602 -12914 15618 -12880
rect 16048 -12914 16064 -12880
rect 16620 -12914 16636 -12880
rect 17066 -12914 17082 -12880
rect 17638 -12914 17654 -12880
rect 18084 -12914 18100 -12880
rect 18656 -12914 18672 -12880
rect 19102 -12914 19118 -12880
rect 19674 -12914 19690 -12880
rect 20120 -12914 20136 -12880
rect 20692 -12914 20708 -12880
rect 21138 -12914 21154 -12880
rect 21710 -12914 21726 -12880
rect 22156 -12914 22172 -12880
rect 22728 -12914 22744 -12880
rect 12238 -12920 12298 -12914
rect -22 -13116 12 -13100
rect 2582 -12964 2616 -12948
rect -8952 -13184 -8936 -13150
rect -8380 -13184 -8364 -13150
rect -7934 -13184 -7918 -13150
rect -7362 -13184 -7346 -13150
rect -6916 -13184 -6900 -13150
rect -6344 -13184 -6328 -13150
rect -5898 -13184 -5882 -13150
rect -5326 -13184 -5310 -13150
rect -4880 -13184 -4864 -13150
rect -4308 -13184 -4292 -13150
rect -3862 -13184 -3846 -13150
rect -3290 -13184 -3274 -13150
rect -2844 -13184 -2828 -13150
rect -2272 -13184 -2256 -13150
rect -1826 -13184 -1810 -13150
rect -1254 -13184 -1238 -13150
rect -808 -13184 -792 -13150
rect -236 -13184 -220 -13150
rect -8952 -13292 -8936 -13258
rect -8380 -13292 -8364 -13258
rect -7934 -13292 -7918 -13258
rect -7362 -13292 -7346 -13258
rect -6916 -13292 -6900 -13258
rect -6344 -13292 -6328 -13258
rect -5898 -13292 -5882 -13258
rect -5326 -13292 -5310 -13258
rect -4880 -13292 -4864 -13258
rect -4308 -13292 -4292 -13258
rect -3862 -13292 -3846 -13258
rect -3290 -13292 -3274 -13258
rect -2844 -13292 -2828 -13258
rect -2272 -13292 -2256 -13258
rect -1826 -13292 -1810 -13258
rect -1254 -13292 -1238 -13258
rect -808 -13292 -792 -13258
rect -236 -13292 -220 -13258
rect -3592 -13294 -3532 -13292
rect -9184 -13342 -9150 -13326
rect -9184 -13934 -9150 -13918
rect -8166 -13342 -8132 -13326
rect -8166 -13934 -8132 -13918
rect -7148 -13342 -7114 -13326
rect -7148 -13934 -7114 -13918
rect -6130 -13342 -6096 -13326
rect -6130 -13934 -6096 -13918
rect -5112 -13342 -5078 -13326
rect -5112 -13934 -5078 -13918
rect -4094 -13342 -4060 -13326
rect -4094 -13934 -4060 -13918
rect -3076 -13342 -3042 -13326
rect -3076 -13934 -3042 -13918
rect -2058 -13342 -2024 -13326
rect -2058 -13934 -2024 -13918
rect -1040 -13342 -1006 -13326
rect -1040 -13934 -1006 -13918
rect -22 -13342 12 -13326
rect 2582 -13556 2616 -13540
rect 3600 -12964 3634 -12948
rect 3600 -13556 3634 -13540
rect 4618 -12964 4652 -12948
rect 4618 -13556 4652 -13540
rect 5636 -12964 5670 -12948
rect 5636 -13556 5670 -13540
rect 6654 -12964 6688 -12948
rect 6654 -13556 6688 -13540
rect 7672 -12964 7706 -12948
rect 7672 -13556 7706 -13540
rect 8690 -12964 8724 -12948
rect 8690 -13556 8724 -13540
rect 9708 -12964 9742 -12948
rect 9708 -13556 9742 -13540
rect 10726 -12964 10760 -12948
rect 10726 -13556 10760 -13540
rect 11744 -12964 11778 -12948
rect 11744 -13556 11778 -13540
rect 12762 -12964 12796 -12948
rect 12762 -13556 12796 -13540
rect 13780 -12964 13814 -12948
rect 13780 -13556 13814 -13540
rect 14798 -12964 14832 -12948
rect 14798 -13556 14832 -13540
rect 15816 -12964 15850 -12948
rect 15816 -13556 15850 -13540
rect 16834 -12964 16868 -12948
rect 16834 -13556 16868 -13540
rect 17852 -12964 17886 -12948
rect 17852 -13556 17886 -13540
rect 18870 -12964 18904 -12948
rect 18870 -13556 18904 -13540
rect 19888 -12964 19922 -12948
rect 19888 -13556 19922 -13540
rect 20906 -12964 20940 -12948
rect 20906 -13556 20940 -13540
rect 21924 -12964 21958 -12948
rect 21924 -13556 21958 -13540
rect 22942 -12964 22976 -12948
rect 22942 -13556 22976 -13540
rect 8166 -13590 8226 -13584
rect 10202 -13590 10262 -13584
rect 11222 -13590 11282 -13584
rect 16294 -13590 16354 -13584
rect 2814 -13624 2830 -13590
rect 3386 -13624 3402 -13590
rect 3832 -13624 3848 -13590
rect 4404 -13624 4420 -13590
rect 4850 -13624 4866 -13590
rect 5422 -13624 5438 -13590
rect 5868 -13624 5884 -13590
rect 6440 -13624 6456 -13590
rect 6886 -13624 6902 -13590
rect 7458 -13624 7474 -13590
rect 7904 -13624 7920 -13590
rect 8476 -13624 8492 -13590
rect 8922 -13624 8938 -13590
rect 9494 -13624 9510 -13590
rect 9940 -13624 9956 -13590
rect 10512 -13624 10528 -13590
rect 10958 -13624 10974 -13590
rect 11530 -13624 11546 -13590
rect 11976 -13624 11992 -13590
rect 12548 -13624 12564 -13590
rect 12994 -13624 13010 -13590
rect 13566 -13624 13582 -13590
rect 14012 -13624 14028 -13590
rect 14584 -13624 14600 -13590
rect 15030 -13624 15046 -13590
rect 15602 -13624 15618 -13590
rect 16048 -13624 16064 -13590
rect 16620 -13624 16636 -13590
rect 17066 -13624 17082 -13590
rect 17638 -13624 17654 -13590
rect 18084 -13624 18100 -13590
rect 18656 -13624 18672 -13590
rect 19102 -13624 19118 -13590
rect 19674 -13624 19690 -13590
rect 20120 -13624 20136 -13590
rect 20692 -13624 20708 -13590
rect 21138 -13624 21154 -13590
rect 21710 -13624 21726 -13590
rect 22156 -13624 22172 -13590
rect 22728 -13624 22744 -13590
rect -22 -13934 12 -13918
rect -7660 -13968 -7600 -13966
rect -6646 -13968 -6586 -13966
rect -2572 -13968 -2512 -13966
rect -1556 -13968 -1496 -13966
rect -8952 -14002 -8936 -13968
rect -8380 -14002 -8364 -13968
rect -7934 -14002 -7918 -13968
rect -7362 -14002 -7346 -13968
rect -6916 -14002 -6900 -13968
rect -6344 -14002 -6328 -13968
rect -5898 -14002 -5882 -13968
rect -5326 -14002 -5310 -13968
rect -4880 -14002 -4864 -13968
rect -4308 -14002 -4292 -13968
rect -3862 -14002 -3846 -13968
rect -3290 -14002 -3274 -13968
rect -2844 -14002 -2828 -13968
rect -2272 -14002 -2256 -13968
rect -1826 -14002 -1810 -13968
rect -1254 -14002 -1238 -13968
rect -808 -14002 -792 -13968
rect -236 -14002 -220 -13968
rect -8952 -14110 -8936 -14076
rect -8380 -14110 -8364 -14076
rect -7934 -14110 -7918 -14076
rect -7362 -14110 -7346 -14076
rect -6916 -14110 -6900 -14076
rect -6344 -14110 -6328 -14076
rect -5898 -14110 -5882 -14076
rect -5326 -14110 -5310 -14076
rect -4880 -14110 -4864 -14076
rect -4308 -14110 -4292 -14076
rect -3862 -14110 -3846 -14076
rect -3290 -14110 -3274 -14076
rect -2844 -14110 -2828 -14076
rect -2272 -14110 -2256 -14076
rect -1826 -14110 -1810 -14076
rect -1254 -14110 -1238 -14076
rect -808 -14110 -792 -14076
rect -236 -14110 -220 -14076
rect -9184 -14160 -9150 -14144
rect -9184 -14752 -9150 -14736
rect -8166 -14160 -8132 -14144
rect -8166 -14752 -8132 -14736
rect -7148 -14160 -7114 -14144
rect -7148 -14752 -7114 -14736
rect -6130 -14160 -6096 -14144
rect -6130 -14752 -6096 -14736
rect -5112 -14160 -5078 -14144
rect -5112 -14752 -5078 -14736
rect -4094 -14160 -4060 -14144
rect -4094 -14752 -4060 -14736
rect -3076 -14160 -3042 -14144
rect -3076 -14752 -3042 -14736
rect -2058 -14160 -2024 -14144
rect -2058 -14752 -2024 -14736
rect -1040 -14160 -1006 -14144
rect -1040 -14752 -1006 -14736
rect -22 -14160 12 -14144
rect 2814 -14146 2830 -14112
rect 3386 -14146 3402 -14112
rect 3832 -14146 3848 -14112
rect 4404 -14146 4420 -14112
rect 4850 -14146 4866 -14112
rect 5422 -14146 5438 -14112
rect 5868 -14146 5884 -14112
rect 6440 -14146 6456 -14112
rect 6886 -14146 6902 -14112
rect 7458 -14146 7474 -14112
rect 7904 -14146 7920 -14112
rect 8476 -14146 8492 -14112
rect 8922 -14146 8938 -14112
rect 9494 -14146 9510 -14112
rect 9940 -14146 9956 -14112
rect 10512 -14146 10528 -14112
rect 10958 -14146 10974 -14112
rect 11530 -14146 11546 -14112
rect 11976 -14146 11992 -14112
rect 12548 -14146 12564 -14112
rect 12994 -14146 13010 -14112
rect 13566 -14146 13582 -14112
rect 14012 -14146 14028 -14112
rect 14584 -14146 14600 -14112
rect 15030 -14146 15046 -14112
rect 15602 -14146 15618 -14112
rect 16048 -14146 16064 -14112
rect 16620 -14146 16636 -14112
rect 17066 -14146 17082 -14112
rect 17638 -14146 17654 -14112
rect 18084 -14146 18100 -14112
rect 18656 -14146 18672 -14112
rect 19102 -14146 19118 -14112
rect 19674 -14146 19690 -14112
rect 20120 -14146 20136 -14112
rect 20692 -14146 20708 -14112
rect 21138 -14146 21154 -14112
rect 21710 -14146 21726 -14112
rect 22156 -14146 22172 -14112
rect 22728 -14146 22744 -14112
rect 4100 -14150 4160 -14146
rect 5116 -14150 5176 -14146
rect 9192 -14154 9252 -14146
rect 13258 -14150 13318 -14146
rect 15292 -14150 15352 -14146
rect 21404 -14150 21464 -14146
rect -22 -14752 12 -14736
rect 2582 -14196 2616 -14180
rect -7656 -14786 -7596 -14784
rect -6642 -14786 -6582 -14784
rect -2568 -14786 -2508 -14784
rect -1552 -14786 -1492 -14784
rect -8952 -14820 -8936 -14786
rect -8380 -14820 -8364 -14786
rect -7934 -14820 -7918 -14786
rect -7362 -14820 -7346 -14786
rect -6916 -14820 -6900 -14786
rect -6344 -14820 -6328 -14786
rect -5898 -14820 -5882 -14786
rect -5326 -14820 -5310 -14786
rect -4880 -14820 -4864 -14786
rect -4308 -14820 -4292 -14786
rect -3862 -14820 -3846 -14786
rect -3290 -14820 -3274 -14786
rect -2844 -14820 -2828 -14786
rect -2272 -14820 -2256 -14786
rect -1826 -14820 -1810 -14786
rect -1254 -14820 -1238 -14786
rect -808 -14820 -792 -14786
rect -236 -14820 -220 -14786
rect 2582 -14788 2616 -14772
rect 3600 -14196 3634 -14180
rect 3600 -14788 3634 -14772
rect 4618 -14196 4652 -14180
rect 4618 -14788 4652 -14772
rect 5636 -14196 5670 -14180
rect 5636 -14788 5670 -14772
rect 6654 -14196 6688 -14180
rect 6654 -14788 6688 -14772
rect 7672 -14196 7706 -14180
rect 7672 -14788 7706 -14772
rect 8690 -14196 8724 -14180
rect 8690 -14788 8724 -14772
rect 9708 -14196 9742 -14180
rect 9708 -14788 9742 -14772
rect 10726 -14196 10760 -14180
rect 10726 -14788 10760 -14772
rect 11744 -14196 11778 -14180
rect 11744 -14788 11778 -14772
rect 12762 -14196 12796 -14180
rect 12762 -14788 12796 -14772
rect 13780 -14196 13814 -14180
rect 13780 -14788 13814 -14772
rect 14798 -14196 14832 -14180
rect 14798 -14788 14832 -14772
rect 15816 -14196 15850 -14180
rect 15816 -14788 15850 -14772
rect 16834 -14196 16868 -14180
rect 16834 -14788 16868 -14772
rect 17852 -14196 17886 -14180
rect 17852 -14788 17886 -14772
rect 18870 -14196 18904 -14180
rect 18870 -14788 18904 -14772
rect 19888 -14196 19922 -14180
rect 19888 -14788 19922 -14772
rect 20906 -14196 20940 -14180
rect 20906 -14788 20940 -14772
rect 21924 -14196 21958 -14180
rect 21924 -14788 21958 -14772
rect 22942 -14196 22976 -14180
rect 22942 -14788 22976 -14772
rect 6126 -14822 6186 -14820
rect 2814 -14856 2830 -14822
rect 3386 -14856 3402 -14822
rect 3832 -14856 3848 -14822
rect 4404 -14856 4420 -14822
rect 4850 -14856 4866 -14822
rect 5422 -14856 5438 -14822
rect 5868 -14856 5884 -14822
rect 6440 -14856 6456 -14822
rect 6886 -14856 6902 -14822
rect 7458 -14856 7474 -14822
rect 7904 -14856 7920 -14822
rect 8476 -14856 8492 -14822
rect 8922 -14856 8938 -14822
rect 9494 -14856 9510 -14822
rect 9940 -14856 9956 -14822
rect 10512 -14856 10528 -14822
rect 10958 -14856 10974 -14822
rect 11530 -14856 11546 -14822
rect 11976 -14856 11992 -14822
rect 12548 -14856 12564 -14822
rect 12994 -14856 13010 -14822
rect 13566 -14856 13582 -14822
rect 14012 -14856 14028 -14822
rect 14584 -14856 14600 -14822
rect 15030 -14856 15046 -14822
rect 15602 -14856 15618 -14822
rect 16048 -14856 16064 -14822
rect 16620 -14856 16636 -14822
rect 17066 -14856 17082 -14822
rect 17638 -14856 17654 -14822
rect 18084 -14856 18100 -14822
rect 18656 -14856 18672 -14822
rect 19102 -14856 19118 -14822
rect 19674 -14856 19690 -14822
rect 20120 -14856 20136 -14822
rect 20692 -14856 20708 -14822
rect 21138 -14856 21154 -14822
rect 21710 -14856 21726 -14822
rect 22156 -14856 22172 -14822
rect 22728 -14856 22744 -14822
rect 8160 -14860 8220 -14856
rect 17318 -14870 17378 -14856
rect 18352 -14870 18412 -14856
rect -8952 -14928 -8936 -14894
rect -8380 -14928 -8364 -14894
rect -7934 -14928 -7918 -14894
rect -7362 -14928 -7346 -14894
rect -6916 -14928 -6900 -14894
rect -6344 -14928 -6328 -14894
rect -5898 -14928 -5882 -14894
rect -5326 -14928 -5310 -14894
rect -4880 -14928 -4864 -14894
rect -4308 -14928 -4292 -14894
rect -3862 -14928 -3846 -14894
rect -3290 -14928 -3274 -14894
rect -2844 -14928 -2828 -14894
rect -2272 -14928 -2256 -14894
rect -1826 -14928 -1810 -14894
rect -1254 -14928 -1238 -14894
rect -808 -14928 -792 -14894
rect -236 -14928 -220 -14894
rect -9184 -14978 -9150 -14962
rect -9184 -15570 -9150 -15554
rect -8166 -14978 -8132 -14962
rect -8166 -15570 -8132 -15554
rect -7148 -14978 -7114 -14962
rect -7148 -15570 -7114 -15554
rect -6130 -14978 -6096 -14962
rect -6130 -15570 -6096 -15554
rect -5112 -14978 -5078 -14962
rect -5112 -15570 -5078 -15554
rect -4094 -14978 -4060 -14962
rect -4094 -15570 -4060 -15554
rect -3076 -14978 -3042 -14962
rect -3076 -15570 -3042 -15554
rect -2058 -14978 -2024 -14962
rect -2058 -15570 -2024 -15554
rect -1040 -14978 -1006 -14962
rect -1040 -15570 -1006 -15554
rect -22 -14978 12 -14962
rect 2812 -15380 2828 -15346
rect 3384 -15380 3400 -15346
rect 3830 -15380 3846 -15346
rect 4402 -15380 4418 -15346
rect 4848 -15380 4864 -15346
rect 5420 -15380 5436 -15346
rect 5866 -15380 5882 -15346
rect 6438 -15380 6454 -15346
rect 6884 -15380 6900 -15346
rect 7456 -15380 7472 -15346
rect 7902 -15380 7918 -15346
rect 8474 -15380 8490 -15346
rect 8920 -15380 8936 -15346
rect 9492 -15380 9508 -15346
rect 9938 -15380 9954 -15346
rect 10510 -15380 10526 -15346
rect 10956 -15380 10972 -15346
rect 11528 -15380 11544 -15346
rect 11974 -15380 11990 -15346
rect 12546 -15380 12562 -15346
rect 12992 -15380 13008 -15346
rect 13564 -15380 13580 -15346
rect 14010 -15380 14026 -15346
rect 14582 -15380 14598 -15346
rect 15028 -15380 15044 -15346
rect 15600 -15380 15616 -15346
rect 16046 -15380 16062 -15346
rect 16618 -15380 16634 -15346
rect 17064 -15380 17080 -15346
rect 17636 -15380 17652 -15346
rect 18082 -15380 18098 -15346
rect 18654 -15380 18670 -15346
rect 19100 -15380 19116 -15346
rect 19672 -15380 19688 -15346
rect 20118 -15380 20134 -15346
rect 20690 -15380 20706 -15346
rect 21136 -15380 21152 -15346
rect 21708 -15380 21724 -15346
rect 22154 -15380 22170 -15346
rect 22726 -15380 22742 -15346
rect 5122 -15384 5182 -15380
rect -22 -15570 12 -15554
rect 2580 -15430 2614 -15414
rect -8952 -15638 -8936 -15604
rect -8380 -15638 -8364 -15604
rect -7934 -15638 -7918 -15604
rect -7362 -15638 -7346 -15604
rect -6916 -15638 -6900 -15604
rect -6344 -15638 -6328 -15604
rect -5898 -15638 -5882 -15604
rect -5326 -15638 -5310 -15604
rect -4880 -15638 -4864 -15604
rect -4308 -15638 -4292 -15604
rect -3862 -15638 -3846 -15604
rect -3290 -15638 -3274 -15604
rect -2844 -15638 -2828 -15604
rect -2272 -15638 -2256 -15604
rect -1826 -15638 -1810 -15604
rect -1254 -15638 -1238 -15604
rect -808 -15638 -792 -15604
rect -236 -15638 -220 -15604
rect -8952 -15746 -8936 -15712
rect -8380 -15746 -8364 -15712
rect -7934 -15746 -7918 -15712
rect -7362 -15746 -7346 -15712
rect -6916 -15746 -6900 -15712
rect -6344 -15746 -6328 -15712
rect -5898 -15746 -5882 -15712
rect -5326 -15746 -5310 -15712
rect -4880 -15746 -4864 -15712
rect -4308 -15746 -4292 -15712
rect -3862 -15746 -3846 -15712
rect -3290 -15746 -3274 -15712
rect -2844 -15746 -2828 -15712
rect -2272 -15746 -2256 -15712
rect -1826 -15746 -1810 -15712
rect -1254 -15746 -1238 -15712
rect -808 -15746 -792 -15712
rect -236 -15746 -220 -15712
rect -3596 -15748 -3536 -15746
rect -9184 -15796 -9150 -15780
rect -9184 -16388 -9150 -16372
rect -8166 -15796 -8132 -15780
rect -8166 -16388 -8132 -16372
rect -7148 -15796 -7114 -15780
rect -7148 -16388 -7114 -16372
rect -6130 -15796 -6096 -15780
rect -6130 -16388 -6096 -16372
rect -5112 -15796 -5078 -15780
rect -5112 -16388 -5078 -16372
rect -4094 -15796 -4060 -15780
rect -4094 -16388 -4060 -16372
rect -3076 -15796 -3042 -15780
rect -3076 -16388 -3042 -16372
rect -2058 -15796 -2024 -15780
rect -2058 -16388 -2024 -16372
rect -1040 -15796 -1006 -15780
rect -1040 -16388 -1006 -16372
rect -22 -15796 12 -15780
rect 2580 -16022 2614 -16006
rect 3598 -15430 3632 -15414
rect 3598 -16022 3632 -16006
rect 4616 -15430 4650 -15414
rect 4616 -16022 4650 -16006
rect 5634 -15430 5668 -15414
rect 5634 -16022 5668 -16006
rect 6652 -15430 6686 -15414
rect 6652 -16022 6686 -16006
rect 7670 -15430 7704 -15414
rect 7670 -16022 7704 -16006
rect 8688 -15430 8722 -15414
rect 8688 -16022 8722 -16006
rect 9706 -15430 9740 -15414
rect 9706 -16022 9740 -16006
rect 10724 -15430 10758 -15414
rect 10724 -16022 10758 -16006
rect 11742 -15430 11776 -15414
rect 11742 -16022 11776 -16006
rect 12760 -15430 12794 -15414
rect 12760 -16022 12794 -16006
rect 13778 -15430 13812 -15414
rect 13778 -16022 13812 -16006
rect 14796 -15430 14830 -15414
rect 14796 -16022 14830 -16006
rect 15814 -15430 15848 -15414
rect 15814 -16022 15848 -16006
rect 16832 -15430 16866 -15414
rect 16832 -16022 16866 -16006
rect 17850 -15430 17884 -15414
rect 17850 -16022 17884 -16006
rect 18868 -15430 18902 -15414
rect 18868 -16022 18902 -16006
rect 19886 -15430 19920 -15414
rect 19886 -16022 19920 -16006
rect 20904 -15430 20938 -15414
rect 20904 -16022 20938 -16006
rect 21922 -15430 21956 -15414
rect 21922 -16022 21956 -16006
rect 22940 -15430 22974 -15414
rect 22940 -16022 22974 -16006
rect 10190 -16056 10250 -16052
rect 11218 -16056 11278 -16054
rect 13262 -16056 13322 -16052
rect 2812 -16090 2828 -16056
rect 3384 -16090 3400 -16056
rect 3830 -16090 3846 -16056
rect 4402 -16090 4418 -16056
rect 4848 -16090 4864 -16056
rect 5420 -16090 5436 -16056
rect 5866 -16090 5882 -16056
rect 6438 -16090 6454 -16056
rect 6884 -16090 6900 -16056
rect 7456 -16090 7472 -16056
rect 7902 -16090 7918 -16056
rect 8474 -16090 8490 -16056
rect 8920 -16090 8936 -16056
rect 9492 -16090 9508 -16056
rect 9938 -16090 9954 -16056
rect 10510 -16090 10526 -16056
rect 10956 -16090 10972 -16056
rect 11528 -16090 11544 -16056
rect 11974 -16090 11990 -16056
rect 12546 -16090 12562 -16056
rect 12992 -16090 13008 -16056
rect 13564 -16090 13580 -16056
rect 14010 -16090 14026 -16056
rect 14582 -16090 14598 -16056
rect 15028 -16090 15044 -16056
rect 15600 -16090 15616 -16056
rect 16046 -16090 16062 -16056
rect 16618 -16090 16634 -16056
rect 17064 -16090 17080 -16056
rect 17636 -16090 17652 -16056
rect 18082 -16090 18098 -16056
rect 18654 -16090 18670 -16056
rect 19100 -16090 19116 -16056
rect 19672 -16090 19688 -16056
rect 20118 -16090 20134 -16056
rect 20690 -16090 20706 -16056
rect 21136 -16090 21152 -16056
rect 21708 -16090 21724 -16056
rect 22154 -16090 22170 -16056
rect 22726 -16090 22742 -16056
rect -22 -16388 12 -16372
rect -7670 -16422 -7610 -16420
rect -6656 -16422 -6596 -16420
rect -2582 -16422 -2522 -16420
rect -1566 -16422 -1506 -16420
rect -8952 -16456 -8936 -16422
rect -8380 -16456 -8364 -16422
rect -7934 -16456 -7918 -16422
rect -7362 -16456 -7346 -16422
rect -6916 -16456 -6900 -16422
rect -6344 -16456 -6328 -16422
rect -5898 -16456 -5882 -16422
rect -5326 -16456 -5310 -16422
rect -4880 -16456 -4864 -16422
rect -4308 -16456 -4292 -16422
rect -3862 -16456 -3846 -16422
rect -3290 -16456 -3274 -16422
rect -2844 -16456 -2828 -16422
rect -2272 -16456 -2256 -16422
rect -1826 -16456 -1810 -16422
rect -1254 -16456 -1238 -16422
rect -808 -16456 -792 -16422
rect -236 -16456 -220 -16422
rect -8952 -16564 -8936 -16530
rect -8380 -16564 -8364 -16530
rect -7934 -16564 -7918 -16530
rect -7362 -16564 -7346 -16530
rect -6916 -16564 -6900 -16530
rect -6344 -16564 -6328 -16530
rect -5898 -16564 -5882 -16530
rect -5326 -16564 -5310 -16530
rect -4880 -16564 -4864 -16530
rect -4308 -16564 -4292 -16530
rect -3862 -16564 -3846 -16530
rect -3290 -16564 -3274 -16530
rect -2844 -16564 -2828 -16530
rect -2272 -16564 -2256 -16530
rect -1826 -16564 -1810 -16530
rect -1254 -16564 -1238 -16530
rect -808 -16564 -792 -16530
rect -236 -16564 -220 -16530
rect -9184 -16614 -9150 -16598
rect -9184 -17206 -9150 -17190
rect -8166 -16614 -8132 -16598
rect -8166 -17206 -8132 -17190
rect -7148 -16614 -7114 -16598
rect -7148 -17206 -7114 -17190
rect -6130 -16614 -6096 -16598
rect -6130 -17206 -6096 -17190
rect -5112 -16614 -5078 -16598
rect -5112 -17206 -5078 -17190
rect -4094 -16614 -4060 -16598
rect -4094 -17206 -4060 -17190
rect -3076 -16614 -3042 -16598
rect -3076 -17206 -3042 -17190
rect -2058 -16614 -2024 -16598
rect -2058 -17206 -2024 -17190
rect -1040 -16614 -1006 -16598
rect -1040 -17206 -1006 -17190
rect -22 -16614 12 -16598
rect 2812 -16614 2828 -16580
rect 3384 -16614 3400 -16580
rect 3830 -16614 3846 -16580
rect 4402 -16614 4418 -16580
rect 4848 -16614 4864 -16580
rect 5420 -16614 5436 -16580
rect 5866 -16614 5882 -16580
rect 6438 -16614 6454 -16580
rect 6884 -16614 6900 -16580
rect 7456 -16614 7472 -16580
rect 7902 -16614 7918 -16580
rect 8474 -16614 8490 -16580
rect 8920 -16614 8936 -16580
rect 9492 -16614 9508 -16580
rect 9938 -16614 9954 -16580
rect 10510 -16614 10526 -16580
rect 10956 -16614 10972 -16580
rect 11528 -16614 11544 -16580
rect 11974 -16614 11990 -16580
rect 12546 -16614 12562 -16580
rect 12992 -16614 13008 -16580
rect 13564 -16614 13580 -16580
rect 14010 -16614 14026 -16580
rect 14582 -16614 14598 -16580
rect 15028 -16614 15044 -16580
rect 15600 -16614 15616 -16580
rect 16046 -16614 16062 -16580
rect 16618 -16614 16634 -16580
rect 17064 -16614 17080 -16580
rect 17636 -16614 17652 -16580
rect 18082 -16614 18098 -16580
rect 18654 -16614 18670 -16580
rect 19100 -16614 19116 -16580
rect 19672 -16614 19688 -16580
rect 20118 -16614 20134 -16580
rect 20690 -16614 20706 -16580
rect 21136 -16614 21152 -16580
rect 21708 -16614 21724 -16580
rect 22154 -16614 22170 -16580
rect 22726 -16614 22742 -16580
rect -22 -17206 12 -17190
rect 2580 -16664 2614 -16648
rect -7666 -17240 -7606 -17238
rect -6652 -17240 -6592 -17238
rect -2578 -17240 -2518 -17238
rect -1562 -17240 -1502 -17238
rect -8952 -17274 -8936 -17240
rect -8380 -17274 -8364 -17240
rect -7934 -17274 -7918 -17240
rect -7362 -17274 -7346 -17240
rect -6916 -17274 -6900 -17240
rect -6344 -17274 -6328 -17240
rect -5898 -17274 -5882 -17240
rect -5326 -17274 -5310 -17240
rect -4880 -17274 -4864 -17240
rect -4308 -17274 -4292 -17240
rect -3862 -17274 -3846 -17240
rect -3290 -17274 -3274 -17240
rect -2844 -17274 -2828 -17240
rect -2272 -17274 -2256 -17240
rect -1826 -17274 -1810 -17240
rect -1254 -17274 -1238 -17240
rect -808 -17274 -792 -17240
rect -236 -17274 -220 -17240
rect 2580 -17256 2614 -17240
rect 3598 -16664 3632 -16648
rect 3598 -17256 3632 -17240
rect 4616 -16664 4650 -16648
rect 4616 -17256 4650 -17240
rect 5634 -16664 5668 -16648
rect 5634 -17256 5668 -17240
rect 6652 -16664 6686 -16648
rect 6652 -17256 6686 -17240
rect 7670 -16664 7704 -16648
rect 7670 -17256 7704 -17240
rect 8688 -16664 8722 -16648
rect 8688 -17256 8722 -17240
rect 9706 -16664 9740 -16648
rect 9706 -17256 9740 -17240
rect 10724 -16664 10758 -16648
rect 10724 -17256 10758 -17240
rect 11742 -16664 11776 -16648
rect 11742 -17256 11776 -17240
rect 12760 -16664 12794 -16648
rect 12760 -17256 12794 -17240
rect 13778 -16664 13812 -16648
rect 13778 -17256 13812 -17240
rect 14796 -16664 14830 -16648
rect 14796 -17256 14830 -17240
rect 15814 -16664 15848 -16648
rect 15814 -17256 15848 -17240
rect 16832 -16664 16866 -16648
rect 16832 -17256 16866 -17240
rect 17850 -16664 17884 -16648
rect 17850 -17256 17884 -17240
rect 18868 -16664 18902 -16648
rect 18868 -17256 18902 -17240
rect 19886 -16664 19920 -16648
rect 19886 -17256 19920 -17240
rect 20904 -16664 20938 -16648
rect 20904 -17256 20938 -17240
rect 21922 -16664 21956 -16648
rect 21922 -17256 21956 -17240
rect 22940 -16664 22974 -16648
rect 22940 -17256 22974 -17240
rect 2812 -17324 2828 -17290
rect 3384 -17324 3400 -17290
rect 3830 -17324 3846 -17290
rect 4402 -17324 4418 -17290
rect 4848 -17324 4864 -17290
rect 5420 -17324 5436 -17290
rect 5866 -17324 5882 -17290
rect 6438 -17324 6454 -17290
rect 6884 -17324 6900 -17290
rect 7456 -17324 7472 -17290
rect 7902 -17324 7918 -17290
rect 8474 -17324 8490 -17290
rect 8920 -17324 8936 -17290
rect 9492 -17324 9508 -17290
rect 9938 -17324 9954 -17290
rect 10510 -17324 10526 -17290
rect 10956 -17324 10972 -17290
rect 11528 -17324 11544 -17290
rect 11974 -17324 11990 -17290
rect 12546 -17324 12562 -17290
rect 12992 -17324 13008 -17290
rect 13564 -17324 13580 -17290
rect 14010 -17324 14026 -17290
rect 14582 -17324 14598 -17290
rect 15028 -17324 15044 -17290
rect 15600 -17324 15616 -17290
rect 16046 -17324 16062 -17290
rect 16618 -17324 16634 -17290
rect 17064 -17324 17080 -17290
rect 17636 -17324 17652 -17290
rect 18082 -17324 18098 -17290
rect 18654 -17324 18670 -17290
rect 19100 -17324 19116 -17290
rect 19672 -17324 19688 -17290
rect 20118 -17324 20134 -17290
rect 20690 -17324 20706 -17290
rect 21136 -17324 21152 -17290
rect 21708 -17324 21724 -17290
rect 22154 -17324 22170 -17290
rect 22726 -17324 22742 -17290
rect -8952 -17382 -8936 -17348
rect -8380 -17382 -8364 -17348
rect -7934 -17382 -7918 -17348
rect -7362 -17382 -7346 -17348
rect -6916 -17382 -6900 -17348
rect -6344 -17382 -6328 -17348
rect -5898 -17382 -5882 -17348
rect -5326 -17382 -5310 -17348
rect -4880 -17382 -4864 -17348
rect -4308 -17382 -4292 -17348
rect -3862 -17382 -3846 -17348
rect -3290 -17382 -3274 -17348
rect -2844 -17382 -2828 -17348
rect -2272 -17382 -2256 -17348
rect -1826 -17382 -1810 -17348
rect -1254 -17382 -1238 -17348
rect -808 -17382 -792 -17348
rect -236 -17382 -220 -17348
rect -9184 -17432 -9150 -17416
rect -9184 -18024 -9150 -18008
rect -8166 -17432 -8132 -17416
rect -8166 -18024 -8132 -18008
rect -7148 -17432 -7114 -17416
rect -7148 -18024 -7114 -18008
rect -6130 -17432 -6096 -17416
rect -6130 -18024 -6096 -18008
rect -5112 -17432 -5078 -17416
rect -5112 -18024 -5078 -18008
rect -4094 -17432 -4060 -17416
rect -4094 -18024 -4060 -18008
rect -3076 -17432 -3042 -17416
rect -3076 -18024 -3042 -18008
rect -2058 -17432 -2024 -17416
rect -2058 -18024 -2024 -18008
rect -1040 -17432 -1006 -17416
rect -1040 -18024 -1006 -18008
rect -22 -17432 12 -17416
rect 2812 -17846 2828 -17812
rect 3384 -17846 3400 -17812
rect 3830 -17846 3846 -17812
rect 4402 -17846 4418 -17812
rect 4848 -17846 4864 -17812
rect 5420 -17846 5436 -17812
rect 5866 -17846 5882 -17812
rect 6438 -17846 6454 -17812
rect 6884 -17846 6900 -17812
rect 7456 -17846 7472 -17812
rect 7902 -17846 7918 -17812
rect 8474 -17846 8490 -17812
rect 8920 -17846 8936 -17812
rect 9492 -17846 9508 -17812
rect 9938 -17846 9954 -17812
rect 10510 -17846 10526 -17812
rect 10956 -17846 10972 -17812
rect 11528 -17846 11544 -17812
rect 11974 -17846 11990 -17812
rect 12546 -17846 12562 -17812
rect 12992 -17846 13008 -17812
rect 13564 -17846 13580 -17812
rect 14010 -17846 14026 -17812
rect 14582 -17846 14598 -17812
rect 15028 -17846 15044 -17812
rect 15600 -17846 15616 -17812
rect 16046 -17846 16062 -17812
rect 16618 -17846 16634 -17812
rect 17064 -17846 17080 -17812
rect 17636 -17846 17652 -17812
rect 18082 -17846 18098 -17812
rect 18654 -17846 18670 -17812
rect 19100 -17846 19116 -17812
rect 19672 -17846 19688 -17812
rect 20118 -17846 20134 -17812
rect 20690 -17846 20706 -17812
rect 21136 -17846 21152 -17812
rect 21708 -17846 21724 -17812
rect 22154 -17846 22170 -17812
rect 22726 -17846 22742 -17812
rect -22 -18024 12 -18008
rect 2580 -17896 2614 -17880
rect -8692 -18058 -8632 -18056
rect -7666 -18058 -7606 -18054
rect -6652 -18058 -6592 -18054
rect -5632 -18058 -5572 -18056
rect -4610 -18058 -4550 -18056
rect -2578 -18058 -2518 -18054
rect -1562 -18058 -1502 -18054
rect -542 -18058 -482 -18056
rect -8952 -18092 -8936 -18058
rect -8380 -18092 -8364 -18058
rect -7934 -18092 -7918 -18058
rect -7362 -18092 -7346 -18058
rect -6916 -18092 -6900 -18058
rect -6344 -18092 -6328 -18058
rect -5898 -18092 -5882 -18058
rect -5326 -18092 -5310 -18058
rect -4880 -18092 -4864 -18058
rect -4308 -18092 -4292 -18058
rect -3862 -18092 -3846 -18058
rect -3290 -18092 -3274 -18058
rect -2844 -18092 -2828 -18058
rect -2272 -18092 -2256 -18058
rect -1826 -18092 -1810 -18058
rect -1254 -18092 -1238 -18058
rect -808 -18092 -792 -18058
rect -236 -18092 -220 -18058
rect -8952 -18200 -8936 -18166
rect -8380 -18200 -8364 -18166
rect -7934 -18200 -7918 -18166
rect -7362 -18200 -7346 -18166
rect -6916 -18200 -6900 -18166
rect -6344 -18200 -6328 -18166
rect -5898 -18200 -5882 -18166
rect -5326 -18200 -5310 -18166
rect -4880 -18200 -4864 -18166
rect -4308 -18200 -4292 -18166
rect -3862 -18200 -3846 -18166
rect -3290 -18200 -3274 -18166
rect -2844 -18200 -2828 -18166
rect -2272 -18200 -2256 -18166
rect -1826 -18200 -1810 -18166
rect -1254 -18200 -1238 -18166
rect -808 -18200 -792 -18166
rect -236 -18200 -220 -18166
rect -9184 -18250 -9150 -18234
rect -9184 -18842 -9150 -18826
rect -8166 -18250 -8132 -18234
rect -8166 -18842 -8132 -18826
rect -7148 -18250 -7114 -18234
rect -7148 -18842 -7114 -18826
rect -6130 -18250 -6096 -18234
rect -6130 -18842 -6096 -18826
rect -5112 -18250 -5078 -18234
rect -5112 -18842 -5078 -18826
rect -4094 -18250 -4060 -18234
rect -4094 -18842 -4060 -18826
rect -3076 -18250 -3042 -18234
rect -3076 -18842 -3042 -18826
rect -2058 -18250 -2024 -18234
rect -2058 -18842 -2024 -18826
rect -1040 -18250 -1006 -18234
rect -1040 -18842 -1006 -18826
rect -22 -18250 12 -18234
rect 2580 -18488 2614 -18472
rect 3598 -17896 3632 -17880
rect 3598 -18488 3632 -18472
rect 4616 -17896 4650 -17880
rect 4616 -18488 4650 -18472
rect 5634 -17896 5668 -17880
rect 5634 -18488 5668 -18472
rect 6652 -17896 6686 -17880
rect 6652 -18488 6686 -18472
rect 7670 -17896 7704 -17880
rect 7670 -18488 7704 -18472
rect 8688 -17896 8722 -17880
rect 8688 -18488 8722 -18472
rect 9706 -17896 9740 -17880
rect 9706 -18488 9740 -18472
rect 10724 -17896 10758 -17880
rect 10724 -18488 10758 -18472
rect 11742 -17896 11776 -17880
rect 11742 -18488 11776 -18472
rect 12760 -17896 12794 -17880
rect 12760 -18488 12794 -18472
rect 13778 -17896 13812 -17880
rect 13778 -18488 13812 -18472
rect 14796 -17896 14830 -17880
rect 14796 -18488 14830 -18472
rect 15814 -17896 15848 -17880
rect 15814 -18488 15848 -18472
rect 16832 -17896 16866 -17880
rect 16832 -18488 16866 -18472
rect 17850 -17896 17884 -17880
rect 17850 -18488 17884 -18472
rect 18868 -17896 18902 -17880
rect 18868 -18488 18902 -18472
rect 19886 -17896 19920 -17880
rect 19886 -18488 19920 -18472
rect 20904 -17896 20938 -17880
rect 20904 -18488 20938 -18472
rect 21922 -17896 21956 -17880
rect 21922 -18488 21956 -18472
rect 22940 -17896 22974 -17880
rect 22940 -18488 22974 -18472
rect 11230 -18522 11290 -18520
rect 13274 -18522 13334 -18518
rect 21408 -18522 21468 -18520
rect 2812 -18556 2828 -18522
rect 3384 -18556 3400 -18522
rect 3830 -18556 3846 -18522
rect 4402 -18556 4418 -18522
rect 4848 -18556 4864 -18522
rect 5420 -18556 5436 -18522
rect 5866 -18556 5882 -18522
rect 6438 -18556 6454 -18522
rect 6884 -18556 6900 -18522
rect 7456 -18556 7472 -18522
rect 7902 -18556 7918 -18522
rect 8474 -18556 8490 -18522
rect 8920 -18556 8936 -18522
rect 9492 -18556 9508 -18522
rect 9938 -18556 9954 -18522
rect 10510 -18556 10526 -18522
rect 10956 -18556 10972 -18522
rect 11528 -18556 11544 -18522
rect 11974 -18556 11990 -18522
rect 12546 -18556 12562 -18522
rect 12992 -18556 13008 -18522
rect 13564 -18556 13580 -18522
rect 14010 -18556 14026 -18522
rect 14582 -18556 14598 -18522
rect 15028 -18556 15044 -18522
rect 15600 -18556 15616 -18522
rect 16046 -18556 16062 -18522
rect 16618 -18556 16634 -18522
rect 17064 -18556 17080 -18522
rect 17636 -18556 17652 -18522
rect 18082 -18556 18098 -18522
rect 18654 -18556 18670 -18522
rect 19100 -18556 19116 -18522
rect 19672 -18556 19688 -18522
rect 20118 -18556 20134 -18522
rect 20690 -18556 20706 -18522
rect 21136 -18556 21152 -18522
rect 21708 -18556 21724 -18522
rect 22154 -18556 22170 -18522
rect 22726 -18556 22742 -18522
rect -22 -18842 12 -18826
rect -8952 -18910 -8936 -18876
rect -8380 -18910 -8364 -18876
rect -7934 -18910 -7918 -18876
rect -7362 -18910 -7346 -18876
rect -6916 -18910 -6900 -18876
rect -6344 -18910 -6328 -18876
rect -5898 -18910 -5882 -18876
rect -5326 -18910 -5310 -18876
rect -4880 -18910 -4864 -18876
rect -4308 -18910 -4292 -18876
rect -3862 -18910 -3846 -18876
rect -3290 -18910 -3274 -18876
rect -2844 -18910 -2828 -18876
rect -2272 -18910 -2256 -18876
rect -1826 -18910 -1810 -18876
rect -1254 -18910 -1238 -18876
rect -808 -18910 -792 -18876
rect -236 -18910 -220 -18876
rect 2812 -19080 2828 -19046
rect 3384 -19080 3400 -19046
rect 3830 -19080 3846 -19046
rect 4402 -19080 4418 -19046
rect 4848 -19080 4864 -19046
rect 5420 -19080 5436 -19046
rect 5866 -19080 5882 -19046
rect 6438 -19080 6454 -19046
rect 6884 -19080 6900 -19046
rect 7456 -19080 7472 -19046
rect 7902 -19080 7918 -19046
rect 8474 -19080 8490 -19046
rect 8920 -19080 8936 -19046
rect 9492 -19080 9508 -19046
rect 9938 -19080 9954 -19046
rect 10510 -19080 10526 -19046
rect 10956 -19080 10972 -19046
rect 11528 -19080 11544 -19046
rect 11974 -19080 11990 -19046
rect 12546 -19080 12562 -19046
rect 12992 -19080 13008 -19046
rect 13564 -19080 13580 -19046
rect 14010 -19080 14026 -19046
rect 14582 -19080 14598 -19046
rect 15028 -19080 15044 -19046
rect 15600 -19080 15616 -19046
rect 16046 -19080 16062 -19046
rect 16618 -19080 16634 -19046
rect 17064 -19080 17080 -19046
rect 17636 -19080 17652 -19046
rect 18082 -19080 18098 -19046
rect 18654 -19080 18670 -19046
rect 19100 -19080 19116 -19046
rect 19672 -19080 19688 -19046
rect 20118 -19080 20134 -19046
rect 20690 -19080 20706 -19046
rect 21136 -19080 21152 -19046
rect 21708 -19080 21724 -19046
rect 22154 -19080 22170 -19046
rect 22726 -19080 22742 -19046
rect 2580 -19130 2614 -19114
rect -2252 -19584 -2236 -19550
rect -2160 -19584 -2144 -19550
rect -2034 -19584 -2018 -19550
rect -1942 -19584 -1926 -19550
rect -1816 -19584 -1800 -19550
rect -1724 -19584 -1708 -19550
rect -1598 -19584 -1582 -19550
rect -1506 -19584 -1490 -19550
rect -1380 -19584 -1364 -19550
rect -1288 -19584 -1272 -19550
rect -1162 -19584 -1146 -19550
rect -1070 -19584 -1054 -19550
rect -944 -19584 -928 -19550
rect -852 -19584 -836 -19550
rect -726 -19584 -710 -19550
rect -634 -19584 -618 -19550
rect -508 -19584 -492 -19550
rect -416 -19584 -400 -19550
rect -290 -19584 -274 -19550
rect -198 -19584 -182 -19550
rect -2324 -19634 -2290 -19618
rect -2324 -19826 -2290 -19810
rect -2106 -19634 -2072 -19618
rect -2106 -19826 -2072 -19810
rect -1888 -19634 -1854 -19618
rect -1888 -19826 -1854 -19810
rect -1670 -19634 -1636 -19618
rect -1670 -19826 -1636 -19810
rect -1452 -19634 -1418 -19618
rect -1452 -19826 -1418 -19810
rect -1234 -19634 -1200 -19618
rect -1234 -19826 -1200 -19810
rect -1016 -19634 -982 -19618
rect -1016 -19826 -982 -19810
rect -798 -19634 -764 -19618
rect -798 -19826 -764 -19810
rect -580 -19634 -546 -19618
rect -580 -19826 -546 -19810
rect -362 -19634 -328 -19618
rect -362 -19826 -328 -19810
rect -144 -19634 -110 -19618
rect 2580 -19722 2614 -19706
rect 3598 -19130 3632 -19114
rect 3598 -19722 3632 -19706
rect 4616 -19130 4650 -19114
rect 4616 -19722 4650 -19706
rect 5634 -19130 5668 -19114
rect 5634 -19722 5668 -19706
rect 6652 -19130 6686 -19114
rect 6652 -19722 6686 -19706
rect 7670 -19130 7704 -19114
rect 7670 -19722 7704 -19706
rect 8688 -19130 8722 -19114
rect 8688 -19722 8722 -19706
rect 9706 -19130 9740 -19114
rect 9706 -19722 9740 -19706
rect 10724 -19130 10758 -19114
rect 10724 -19722 10758 -19706
rect 11742 -19130 11776 -19114
rect 11742 -19722 11776 -19706
rect 12760 -19130 12794 -19114
rect 12760 -19722 12794 -19706
rect 13778 -19130 13812 -19114
rect 13778 -19722 13812 -19706
rect 14796 -19130 14830 -19114
rect 14796 -19722 14830 -19706
rect 15814 -19130 15848 -19114
rect 15814 -19722 15848 -19706
rect 16832 -19130 16866 -19114
rect 16832 -19722 16866 -19706
rect 17850 -19130 17884 -19114
rect 17850 -19722 17884 -19706
rect 18868 -19130 18902 -19114
rect 18868 -19722 18902 -19706
rect 19886 -19130 19920 -19114
rect 19886 -19722 19920 -19706
rect 20904 -19130 20938 -19114
rect 20904 -19722 20938 -19706
rect 21922 -19130 21956 -19114
rect 21922 -19722 21956 -19706
rect 22940 -19130 22974 -19114
rect 22940 -19722 22974 -19706
rect 5106 -19756 5166 -19752
rect 2812 -19790 2828 -19756
rect 3384 -19790 3400 -19756
rect 3830 -19790 3846 -19756
rect 4402 -19790 4418 -19756
rect 4848 -19790 4864 -19756
rect 5420 -19790 5436 -19756
rect 5866 -19790 5882 -19756
rect 6438 -19790 6454 -19756
rect 6884 -19790 6900 -19756
rect 7456 -19790 7472 -19756
rect 7902 -19790 7918 -19756
rect 8474 -19790 8490 -19756
rect 8920 -19790 8936 -19756
rect 9492 -19790 9508 -19756
rect 9938 -19790 9954 -19756
rect 10510 -19790 10526 -19756
rect 10956 -19790 10972 -19756
rect 11528 -19790 11544 -19756
rect 11974 -19790 11990 -19756
rect 12546 -19790 12562 -19756
rect 12992 -19790 13008 -19756
rect 13564 -19790 13580 -19756
rect 14010 -19790 14026 -19756
rect 14582 -19790 14598 -19756
rect 15028 -19790 15044 -19756
rect 15600 -19790 15616 -19756
rect 16046 -19790 16062 -19756
rect 16618 -19790 16634 -19756
rect 17064 -19790 17080 -19756
rect 17636 -19790 17652 -19756
rect 18082 -19790 18098 -19756
rect 18654 -19790 18670 -19756
rect 19100 -19790 19116 -19756
rect 19672 -19790 19688 -19756
rect 20118 -19790 20134 -19756
rect 20690 -19790 20706 -19756
rect 21136 -19790 21152 -19756
rect 21708 -19790 21724 -19756
rect 22154 -19790 22170 -19756
rect 22726 -19790 22742 -19756
rect -144 -19826 -110 -19810
rect -2252 -19894 -2236 -19860
rect -2160 -19894 -2144 -19860
rect -2034 -19894 -2018 -19860
rect -1942 -19894 -1926 -19860
rect -1816 -19894 -1800 -19860
rect -1724 -19894 -1708 -19860
rect -1598 -19894 -1582 -19860
rect -1506 -19894 -1490 -19860
rect -1380 -19894 -1364 -19860
rect -1288 -19894 -1272 -19860
rect -1162 -19894 -1146 -19860
rect -1070 -19894 -1054 -19860
rect -944 -19894 -928 -19860
rect -852 -19894 -836 -19860
rect -726 -19894 -710 -19860
rect -634 -19894 -618 -19860
rect -508 -19894 -492 -19860
rect -416 -19894 -400 -19860
rect -290 -19894 -274 -19860
rect -198 -19894 -182 -19860
rect 2812 -20314 2828 -20280
rect 3384 -20314 3400 -20280
rect 3830 -20314 3846 -20280
rect 4402 -20314 4418 -20280
rect 4848 -20314 4864 -20280
rect 5420 -20314 5436 -20280
rect 5866 -20314 5882 -20280
rect 6438 -20314 6454 -20280
rect 6884 -20314 6900 -20280
rect 7456 -20314 7472 -20280
rect 7902 -20314 7918 -20280
rect 8474 -20314 8490 -20280
rect 8920 -20314 8936 -20280
rect 9492 -20314 9508 -20280
rect 9938 -20314 9954 -20280
rect 10510 -20314 10526 -20280
rect 10956 -20314 10972 -20280
rect 11528 -20314 11544 -20280
rect 11974 -20314 11990 -20280
rect 12546 -20314 12562 -20280
rect 12992 -20314 13008 -20280
rect 13564 -20314 13580 -20280
rect 14010 -20314 14026 -20280
rect 14582 -20314 14598 -20280
rect 15028 -20314 15044 -20280
rect 15600 -20314 15616 -20280
rect 16046 -20314 16062 -20280
rect 16618 -20314 16634 -20280
rect 17064 -20314 17080 -20280
rect 17636 -20314 17652 -20280
rect 18082 -20314 18098 -20280
rect 18654 -20314 18670 -20280
rect 19100 -20314 19116 -20280
rect 19672 -20314 19688 -20280
rect 20118 -20314 20134 -20280
rect 20690 -20314 20706 -20280
rect 21136 -20314 21152 -20280
rect 21708 -20314 21724 -20280
rect 22154 -20314 22170 -20280
rect 22726 -20314 22742 -20280
rect 2580 -20364 2614 -20348
rect -2252 -20416 -2236 -20382
rect -2160 -20416 -2144 -20382
rect -2034 -20416 -2018 -20382
rect -1942 -20416 -1926 -20382
rect -1816 -20416 -1800 -20382
rect -1724 -20416 -1708 -20382
rect -1598 -20416 -1582 -20382
rect -1506 -20416 -1490 -20382
rect -1380 -20416 -1364 -20382
rect -1288 -20416 -1272 -20382
rect -1162 -20416 -1146 -20382
rect -1070 -20416 -1054 -20382
rect -944 -20416 -928 -20382
rect -852 -20416 -836 -20382
rect -726 -20416 -710 -20382
rect -634 -20416 -618 -20382
rect -508 -20416 -492 -20382
rect -416 -20416 -400 -20382
rect -290 -20416 -274 -20382
rect -198 -20416 -182 -20382
rect -2324 -20466 -2290 -20450
rect -2324 -20658 -2290 -20642
rect -2106 -20466 -2072 -20450
rect -2106 -20658 -2072 -20642
rect -1888 -20466 -1854 -20450
rect -1888 -20658 -1854 -20642
rect -1670 -20466 -1636 -20450
rect -1670 -20658 -1636 -20642
rect -1452 -20466 -1418 -20450
rect -1452 -20658 -1418 -20642
rect -1234 -20466 -1200 -20450
rect -1234 -20658 -1200 -20642
rect -1016 -20466 -982 -20450
rect -1016 -20658 -982 -20642
rect -798 -20466 -764 -20450
rect -798 -20658 -764 -20642
rect -580 -20466 -546 -20450
rect -580 -20658 -546 -20642
rect -362 -20466 -328 -20450
rect -362 -20658 -328 -20642
rect -144 -20466 -110 -20450
rect -144 -20658 -110 -20642
rect -2252 -20726 -2236 -20692
rect -2160 -20726 -2144 -20692
rect -2034 -20726 -2018 -20692
rect -1942 -20726 -1926 -20692
rect -1816 -20726 -1800 -20692
rect -1724 -20726 -1708 -20692
rect -1598 -20726 -1582 -20692
rect -1506 -20726 -1490 -20692
rect -1380 -20726 -1364 -20692
rect -1288 -20726 -1272 -20692
rect -1162 -20726 -1146 -20692
rect -1070 -20726 -1054 -20692
rect -944 -20726 -928 -20692
rect -852 -20726 -836 -20692
rect -726 -20726 -710 -20692
rect -634 -20726 -618 -20692
rect -508 -20726 -492 -20692
rect -416 -20726 -400 -20692
rect -290 -20726 -274 -20692
rect -198 -20726 -182 -20692
rect 2580 -20956 2614 -20940
rect 3598 -20364 3632 -20348
rect 3598 -20956 3632 -20940
rect 4616 -20364 4650 -20348
rect 4616 -20956 4650 -20940
rect 5634 -20364 5668 -20348
rect 5634 -20956 5668 -20940
rect 6652 -20364 6686 -20348
rect 6652 -20956 6686 -20940
rect 7670 -20364 7704 -20348
rect 7670 -20956 7704 -20940
rect 8688 -20364 8722 -20348
rect 8688 -20956 8722 -20940
rect 9706 -20364 9740 -20348
rect 9706 -20956 9740 -20940
rect 10724 -20364 10758 -20348
rect 10724 -20956 10758 -20940
rect 11742 -20364 11776 -20348
rect 11742 -20956 11776 -20940
rect 12760 -20364 12794 -20348
rect 12760 -20956 12794 -20940
rect 13778 -20364 13812 -20348
rect 13778 -20956 13812 -20940
rect 14796 -20364 14830 -20348
rect 14796 -20956 14830 -20940
rect 15814 -20364 15848 -20348
rect 15814 -20956 15848 -20940
rect 16832 -20364 16866 -20348
rect 16832 -20956 16866 -20940
rect 17850 -20364 17884 -20348
rect 17850 -20956 17884 -20940
rect 18868 -20364 18902 -20348
rect 18868 -20956 18902 -20940
rect 19886 -20364 19920 -20348
rect 19886 -20956 19920 -20940
rect 20904 -20364 20938 -20348
rect 20904 -20956 20938 -20940
rect 21922 -20364 21956 -20348
rect 21922 -20956 21956 -20940
rect 22940 -20364 22974 -20348
rect 22940 -20956 22974 -20940
rect 11230 -20990 11290 -20988
rect 13274 -20990 13334 -20986
rect 16312 -20990 16372 -20986
rect 2812 -21024 2828 -20990
rect 3384 -21024 3400 -20990
rect 3830 -21024 3846 -20990
rect 4402 -21024 4418 -20990
rect 4848 -21024 4864 -20990
rect 5420 -21024 5436 -20990
rect 5866 -21024 5882 -20990
rect 6438 -21024 6454 -20990
rect 6884 -21024 6900 -20990
rect 7456 -21024 7472 -20990
rect 7902 -21024 7918 -20990
rect 8474 -21024 8490 -20990
rect 8920 -21024 8936 -20990
rect 9492 -21024 9508 -20990
rect 9938 -21024 9954 -20990
rect 10510 -21024 10526 -20990
rect 10956 -21024 10972 -20990
rect 11528 -21024 11544 -20990
rect 11974 -21024 11990 -20990
rect 12546 -21024 12562 -20990
rect 12992 -21024 13008 -20990
rect 13564 -21024 13580 -20990
rect 14010 -21024 14026 -20990
rect 14582 -21024 14598 -20990
rect 15028 -21024 15044 -20990
rect 15600 -21024 15616 -20990
rect 16046 -21024 16062 -20990
rect 16618 -21024 16634 -20990
rect 17064 -21024 17080 -20990
rect 17636 -21024 17652 -20990
rect 18082 -21024 18098 -20990
rect 18654 -21024 18670 -20990
rect 19100 -21024 19116 -20990
rect 19672 -21024 19688 -20990
rect 20118 -21024 20134 -20990
rect 20690 -21024 20706 -20990
rect 21136 -21024 21152 -20990
rect 21708 -21024 21724 -20990
rect 22154 -21024 22170 -20990
rect 22726 -21024 22742 -20990
rect 2812 -21546 2828 -21512
rect 3384 -21546 3400 -21512
rect 3830 -21546 3846 -21512
rect 4402 -21546 4418 -21512
rect 4848 -21546 4864 -21512
rect 5420 -21546 5436 -21512
rect 5866 -21546 5882 -21512
rect 6438 -21546 6454 -21512
rect 6884 -21546 6900 -21512
rect 7456 -21546 7472 -21512
rect 7902 -21546 7918 -21512
rect 8474 -21546 8490 -21512
rect 8920 -21546 8936 -21512
rect 9492 -21546 9508 -21512
rect 9938 -21546 9954 -21512
rect 10510 -21546 10526 -21512
rect 10956 -21546 10972 -21512
rect 11528 -21546 11544 -21512
rect 11974 -21546 11990 -21512
rect 12546 -21546 12562 -21512
rect 12992 -21546 13008 -21512
rect 13564 -21546 13580 -21512
rect 14010 -21546 14026 -21512
rect 14582 -21546 14598 -21512
rect 15028 -21546 15044 -21512
rect 15600 -21546 15616 -21512
rect 16046 -21546 16062 -21512
rect 16618 -21546 16634 -21512
rect 17064 -21546 17080 -21512
rect 17636 -21546 17652 -21512
rect 18082 -21546 18098 -21512
rect 18654 -21546 18670 -21512
rect 19100 -21546 19116 -21512
rect 19672 -21546 19688 -21512
rect 20118 -21546 20134 -21512
rect 20690 -21546 20706 -21512
rect 21136 -21546 21152 -21512
rect 21708 -21546 21724 -21512
rect 22154 -21546 22170 -21512
rect 22726 -21546 22742 -21512
rect 6134 -21548 6194 -21546
rect 2580 -21596 2614 -21580
rect -9173 -21743 -9157 -21709
rect -8601 -21743 -8585 -21709
rect -8155 -21743 -8139 -21709
rect -7583 -21743 -7567 -21709
rect -7137 -21743 -7121 -21709
rect -6565 -21743 -6549 -21709
rect -6119 -21743 -6103 -21709
rect -5547 -21743 -5531 -21709
rect -5101 -21743 -5085 -21709
rect -4529 -21743 -4513 -21709
rect -4083 -21743 -4067 -21709
rect -3511 -21743 -3495 -21709
rect -2322 -21742 -2306 -21708
rect -2182 -21742 -2166 -21708
rect -2024 -21742 -2008 -21708
rect -1884 -21742 -1868 -21708
rect -1726 -21742 -1710 -21708
rect -1586 -21742 -1570 -21708
rect -1428 -21742 -1412 -21708
rect -1288 -21742 -1272 -21708
rect -1130 -21742 -1114 -21708
rect -990 -21742 -974 -21708
rect -832 -21742 -816 -21708
rect -692 -21742 -676 -21708
rect -534 -21742 -518 -21708
rect -394 -21742 -378 -21708
rect -236 -21742 -220 -21708
rect -96 -21742 -80 -21708
rect 62 -21742 78 -21708
rect 202 -21742 218 -21708
rect 360 -21742 376 -21708
rect 500 -21742 516 -21708
rect 658 -21742 674 -21708
rect 798 -21742 814 -21708
rect -9405 -21793 -9371 -21777
rect -9405 -22385 -9371 -22369
rect -8387 -21793 -8353 -21777
rect -8387 -22385 -8353 -22369
rect -7369 -21793 -7335 -21777
rect -7369 -22385 -7335 -22369
rect -6351 -21793 -6317 -21777
rect -6351 -22385 -6317 -22369
rect -5333 -21793 -5299 -21777
rect -5333 -22385 -5299 -22369
rect -4315 -21793 -4281 -21777
rect -4315 -22385 -4281 -22369
rect -3297 -21793 -3263 -21777
rect -3297 -22385 -3263 -22369
rect -2410 -21792 -2376 -21776
rect -2410 -22384 -2376 -22368
rect -2112 -21792 -2078 -21776
rect -2112 -22384 -2078 -22368
rect -1814 -21792 -1780 -21776
rect -1814 -22384 -1780 -22368
rect -1516 -21792 -1482 -21776
rect -1516 -22384 -1482 -22368
rect -1218 -21792 -1184 -21776
rect -1218 -22384 -1184 -22368
rect -920 -21792 -886 -21776
rect -920 -22384 -886 -22368
rect -622 -21792 -588 -21776
rect -622 -22384 -588 -22368
rect -324 -21792 -290 -21776
rect -324 -22384 -290 -22368
rect -26 -21792 8 -21776
rect -26 -22384 8 -22368
rect 272 -21792 306 -21776
rect 272 -22384 306 -22368
rect 570 -21792 604 -21776
rect 570 -22384 604 -22368
rect 868 -21792 902 -21776
rect 2580 -22188 2614 -22172
rect 3598 -21596 3632 -21580
rect 3598 -22188 3632 -22172
rect 4616 -21596 4650 -21580
rect 4616 -22188 4650 -22172
rect 5634 -21596 5668 -21580
rect 5634 -22188 5668 -22172
rect 6652 -21596 6686 -21580
rect 6652 -22188 6686 -22172
rect 7670 -21596 7704 -21580
rect 7670 -22188 7704 -22172
rect 8688 -21596 8722 -21580
rect 8688 -22188 8722 -22172
rect 9706 -21596 9740 -21580
rect 9706 -22188 9740 -22172
rect 10724 -21596 10758 -21580
rect 10724 -22188 10758 -22172
rect 11742 -21596 11776 -21580
rect 11742 -22188 11776 -22172
rect 12760 -21596 12794 -21580
rect 12760 -22188 12794 -22172
rect 13778 -21596 13812 -21580
rect 13778 -22188 13812 -22172
rect 14796 -21596 14830 -21580
rect 14796 -22188 14830 -22172
rect 15814 -21596 15848 -21580
rect 15814 -22188 15848 -22172
rect 16832 -21596 16866 -21580
rect 16832 -22188 16866 -22172
rect 17850 -21596 17884 -21580
rect 17850 -22188 17884 -22172
rect 18868 -21596 18902 -21580
rect 18868 -22188 18902 -22172
rect 19886 -21596 19920 -21580
rect 19886 -22188 19920 -22172
rect 20904 -21596 20938 -21580
rect 21922 -21596 21956 -21580
rect 22940 -21596 22974 -21580
rect 20904 -22188 20938 -22172
rect 22940 -22188 22974 -22172
rect 10206 -22222 10266 -22212
rect 2812 -22256 2828 -22222
rect 3384 -22256 3400 -22222
rect 3830 -22256 3846 -22222
rect 4402 -22256 4418 -22222
rect 4848 -22256 4864 -22222
rect 5420 -22256 5436 -22222
rect 5866 -22256 5882 -22222
rect 6438 -22256 6454 -22222
rect 6884 -22256 6900 -22222
rect 7456 -22256 7472 -22222
rect 7902 -22256 7918 -22222
rect 8474 -22256 8490 -22222
rect 8920 -22256 8936 -22222
rect 9492 -22256 9508 -22222
rect 9938 -22256 9954 -22222
rect 10510 -22256 10526 -22222
rect 10956 -22256 10972 -22222
rect 11528 -22256 11544 -22222
rect 11974 -22256 11990 -22222
rect 12546 -22256 12562 -22222
rect 12992 -22256 13008 -22222
rect 13564 -22256 13580 -22222
rect 14010 -22256 14026 -22222
rect 14582 -22256 14598 -22222
rect 15028 -22256 15044 -22222
rect 15600 -22256 15616 -22222
rect 16046 -22256 16062 -22222
rect 16618 -22256 16634 -22222
rect 17064 -22256 17080 -22222
rect 17636 -22256 17652 -22222
rect 18082 -22256 18098 -22222
rect 18654 -22256 18670 -22222
rect 19100 -22256 19116 -22222
rect 19672 -22256 19688 -22222
rect 20118 -22256 20134 -22222
rect 20690 -22256 20706 -22222
rect 21136 -22256 21152 -22222
rect 21708 -22256 21724 -22222
rect 22154 -22256 22170 -22222
rect 22726 -22256 22742 -22222
rect 868 -22384 902 -22368
rect -7892 -22419 -7832 -22418
rect -6882 -22419 -6822 -22418
rect -4834 -22419 -4774 -22418
rect -9173 -22453 -9157 -22419
rect -8601 -22453 -8585 -22419
rect -8155 -22453 -8139 -22419
rect -7583 -22453 -7567 -22419
rect -7137 -22453 -7121 -22419
rect -6565 -22453 -6549 -22419
rect -6119 -22453 -6103 -22419
rect -5547 -22453 -5531 -22419
rect -5101 -22453 -5085 -22419
rect -4529 -22453 -4513 -22419
rect -4083 -22453 -4067 -22419
rect -3511 -22453 -3495 -22419
rect -2322 -22452 -2306 -22418
rect -2182 -22452 -2166 -22418
rect -2024 -22452 -2008 -22418
rect -1884 -22452 -1868 -22418
rect -1726 -22452 -1710 -22418
rect -1586 -22452 -1570 -22418
rect -1428 -22452 -1412 -22418
rect -1288 -22452 -1272 -22418
rect -1130 -22452 -1114 -22418
rect -990 -22452 -974 -22418
rect -832 -22452 -816 -22418
rect -692 -22452 -676 -22418
rect -534 -22452 -518 -22418
rect -394 -22452 -378 -22418
rect -236 -22452 -220 -22418
rect -96 -22452 -80 -22418
rect 62 -22452 78 -22418
rect 202 -22452 218 -22418
rect 360 -22452 376 -22418
rect 500 -22452 516 -22418
rect 658 -22452 674 -22418
rect 798 -22452 814 -22418
rect -1974 -22472 -1914 -22452
rect 2812 -22780 2828 -22746
rect 3384 -22780 3400 -22746
rect 3830 -22780 3846 -22746
rect 4402 -22780 4418 -22746
rect 4848 -22780 4864 -22746
rect 5420 -22780 5436 -22746
rect 5866 -22780 5882 -22746
rect 6438 -22780 6454 -22746
rect 6884 -22780 6900 -22746
rect 7456 -22780 7472 -22746
rect 7902 -22780 7918 -22746
rect 8474 -22780 8490 -22746
rect 8920 -22780 8936 -22746
rect 9492 -22780 9508 -22746
rect 9938 -22780 9954 -22746
rect 10510 -22780 10526 -22746
rect 10956 -22780 10972 -22746
rect 11528 -22780 11544 -22746
rect 11974 -22780 11990 -22746
rect 12546 -22780 12562 -22746
rect 12992 -22780 13008 -22746
rect 13564 -22780 13580 -22746
rect 14010 -22780 14026 -22746
rect 14582 -22780 14598 -22746
rect 15028 -22780 15044 -22746
rect 15600 -22780 15616 -22746
rect 16046 -22780 16062 -22746
rect 16618 -22780 16634 -22746
rect 17064 -22780 17080 -22746
rect 17636 -22780 17652 -22746
rect 18082 -22780 18098 -22746
rect 18654 -22780 18670 -22746
rect 19100 -22780 19116 -22746
rect 19672 -22780 19688 -22746
rect 20118 -22780 20134 -22746
rect 20690 -22780 20706 -22746
rect 21136 -22780 21152 -22746
rect 21708 -22780 21724 -22746
rect 22154 -22780 22170 -22746
rect 22726 -22780 22742 -22746
rect 6120 -22782 6180 -22780
rect -9174 -22856 -9158 -22822
rect -8602 -22856 -8586 -22822
rect -8156 -22856 -8140 -22822
rect -7584 -22856 -7568 -22822
rect -7138 -22856 -7122 -22822
rect -6566 -22856 -6550 -22822
rect -6120 -22856 -6104 -22822
rect -5548 -22856 -5532 -22822
rect -5102 -22856 -5086 -22822
rect -4530 -22856 -4514 -22822
rect -4084 -22856 -4068 -22822
rect -3512 -22856 -3496 -22822
rect -2322 -22854 -2306 -22820
rect -2182 -22854 -2166 -22820
rect -2024 -22854 -2008 -22820
rect -1884 -22854 -1868 -22820
rect -1726 -22854 -1710 -22820
rect -1586 -22854 -1570 -22820
rect -1428 -22854 -1412 -22820
rect -1288 -22854 -1272 -22820
rect -1130 -22854 -1114 -22820
rect -990 -22854 -974 -22820
rect -832 -22854 -816 -22820
rect -692 -22854 -676 -22820
rect -534 -22854 -518 -22820
rect -394 -22854 -378 -22820
rect -236 -22854 -220 -22820
rect -96 -22854 -80 -22820
rect 62 -22854 78 -22820
rect 202 -22854 218 -22820
rect 360 -22854 376 -22820
rect 500 -22854 516 -22820
rect 658 -22854 674 -22820
rect 798 -22854 814 -22820
rect 2580 -22830 2614 -22814
rect -7892 -22858 -7832 -22856
rect -5856 -22858 -5796 -22856
rect -4834 -22858 -4774 -22856
rect -9406 -22906 -9372 -22890
rect -9406 -23498 -9372 -23482
rect -8388 -22906 -8354 -22890
rect -8388 -23498 -8354 -23482
rect -7370 -22906 -7336 -22890
rect -7370 -23498 -7336 -23482
rect -6352 -22906 -6318 -22890
rect -6352 -23498 -6318 -23482
rect -5334 -22906 -5300 -22890
rect -5334 -23498 -5300 -23482
rect -4316 -22906 -4282 -22890
rect -4316 -23498 -4282 -23482
rect -3298 -22906 -3264 -22890
rect -3298 -23498 -3264 -23482
rect -2410 -22904 -2376 -22888
rect -2410 -23496 -2376 -23480
rect -2112 -22904 -2078 -22888
rect -2112 -23496 -2078 -23480
rect -1814 -22904 -1780 -22888
rect -1814 -23496 -1780 -23480
rect -1516 -22904 -1482 -22888
rect -1516 -23496 -1482 -23480
rect -1218 -22904 -1184 -22888
rect -1218 -23496 -1184 -23480
rect -920 -22904 -886 -22888
rect -920 -23496 -886 -23480
rect -622 -22904 -588 -22888
rect -622 -23496 -588 -23480
rect -324 -22904 -290 -22888
rect -324 -23496 -290 -23480
rect -26 -22904 8 -22888
rect -26 -23496 8 -23480
rect 272 -22904 306 -22888
rect 272 -23496 306 -23480
rect 570 -22904 604 -22888
rect 570 -23496 604 -23480
rect 868 -22904 902 -22888
rect 2580 -23422 2614 -23406
rect 3598 -22830 3632 -22814
rect 3598 -23422 3632 -23406
rect 4616 -22830 4650 -22814
rect 4616 -23422 4650 -23406
rect 5634 -22830 5668 -22814
rect 5634 -23422 5668 -23406
rect 6652 -22830 6686 -22814
rect 6652 -23422 6686 -23406
rect 7670 -22830 7704 -22814
rect 7670 -23422 7704 -23406
rect 8688 -22830 8722 -22814
rect 8688 -23422 8722 -23406
rect 9706 -22830 9740 -22814
rect 9706 -23422 9740 -23406
rect 10724 -22830 10758 -22814
rect 10724 -23422 10758 -23406
rect 11742 -22830 11776 -22814
rect 11742 -23422 11776 -23406
rect 12760 -22830 12794 -22814
rect 12760 -23422 12794 -23406
rect 13778 -22830 13812 -22814
rect 13778 -23422 13812 -23406
rect 14796 -22830 14830 -22814
rect 14796 -23422 14830 -23406
rect 15814 -22830 15848 -22814
rect 15814 -23422 15848 -23406
rect 16832 -22830 16866 -22814
rect 16832 -23422 16866 -23406
rect 17850 -22830 17884 -22814
rect 17850 -23422 17884 -23406
rect 18868 -22830 18902 -22814
rect 18868 -23422 18902 -23406
rect 19886 -22830 19920 -22814
rect 19886 -23422 19920 -23406
rect 20904 -22830 20938 -22814
rect 20904 -23422 20938 -23406
rect 21922 -22830 21956 -22814
rect 21922 -23422 21956 -23406
rect 22940 -22830 22974 -22814
rect 22940 -23422 22974 -23406
rect 4088 -23456 4148 -23454
rect 10200 -23456 10260 -23454
rect 12234 -23456 12294 -23454
rect 16300 -23456 16360 -23450
rect 20376 -23456 20436 -23454
rect 21392 -23456 21452 -23454
rect 868 -23496 902 -23480
rect 2812 -23490 2828 -23456
rect 3384 -23490 3400 -23456
rect 3830 -23490 3846 -23456
rect 4402 -23490 4418 -23456
rect 4848 -23490 4864 -23456
rect 5420 -23490 5436 -23456
rect 5866 -23490 5882 -23456
rect 6438 -23490 6454 -23456
rect 6884 -23490 6900 -23456
rect 7456 -23490 7472 -23456
rect 7902 -23490 7918 -23456
rect 8474 -23490 8490 -23456
rect 8920 -23490 8936 -23456
rect 9492 -23490 9508 -23456
rect 9938 -23490 9954 -23456
rect 10510 -23490 10526 -23456
rect 10956 -23490 10972 -23456
rect 11528 -23490 11544 -23456
rect 11974 -23490 11990 -23456
rect 12546 -23490 12562 -23456
rect 12992 -23490 13008 -23456
rect 13564 -23490 13580 -23456
rect 14010 -23490 14026 -23456
rect 14582 -23490 14598 -23456
rect 15028 -23490 15044 -23456
rect 15600 -23490 15616 -23456
rect 16046 -23490 16062 -23456
rect 16618 -23490 16634 -23456
rect 17064 -23490 17080 -23456
rect 17636 -23490 17652 -23456
rect 18082 -23490 18098 -23456
rect 18654 -23490 18670 -23456
rect 19100 -23490 19116 -23456
rect 19672 -23490 19688 -23456
rect 20118 -23490 20134 -23456
rect 20690 -23490 20706 -23456
rect 21136 -23490 21152 -23456
rect 21708 -23490 21724 -23456
rect 22154 -23490 22170 -23456
rect 22726 -23490 22742 -23456
rect -7890 -23532 -7830 -23528
rect -6880 -23532 -6820 -23528
rect -4832 -23532 -4772 -23528
rect -9174 -23566 -9158 -23532
rect -8602 -23566 -8586 -23532
rect -8156 -23566 -8140 -23532
rect -7584 -23566 -7568 -23532
rect -7138 -23566 -7122 -23532
rect -6566 -23566 -6550 -23532
rect -6120 -23566 -6104 -23532
rect -5548 -23566 -5532 -23532
rect -5102 -23566 -5086 -23532
rect -4530 -23566 -4514 -23532
rect -4084 -23566 -4068 -23532
rect -3512 -23566 -3496 -23532
rect -2322 -23564 -2306 -23530
rect -2182 -23564 -2166 -23530
rect -2024 -23564 -2008 -23530
rect -1884 -23564 -1868 -23530
rect -1726 -23564 -1710 -23530
rect -1586 -23564 -1570 -23530
rect -1428 -23564 -1412 -23530
rect -1288 -23564 -1272 -23530
rect -1130 -23564 -1114 -23530
rect -990 -23564 -974 -23530
rect -832 -23564 -816 -23530
rect -692 -23564 -676 -23530
rect -534 -23564 -518 -23530
rect -394 -23564 -378 -23530
rect -236 -23564 -220 -23530
rect -96 -23564 -80 -23530
rect 62 -23564 78 -23530
rect 202 -23564 218 -23530
rect 360 -23564 376 -23530
rect 500 -23564 516 -23530
rect 658 -23564 674 -23530
rect 798 -23564 814 -23530
rect -9173 -23967 -9157 -23933
rect -8601 -23967 -8585 -23933
rect -8155 -23967 -8139 -23933
rect -7583 -23967 -7567 -23933
rect -7137 -23967 -7121 -23933
rect -6565 -23967 -6549 -23933
rect -6119 -23967 -6103 -23933
rect -5547 -23967 -5531 -23933
rect -5101 -23967 -5085 -23933
rect -4529 -23967 -4513 -23933
rect -4083 -23967 -4067 -23933
rect -3511 -23967 -3495 -23933
rect -2324 -23966 -2308 -23932
rect -2184 -23966 -2168 -23932
rect -2026 -23966 -2010 -23932
rect -1886 -23966 -1870 -23932
rect -1728 -23966 -1712 -23932
rect -1588 -23966 -1572 -23932
rect -1430 -23966 -1414 -23932
rect -1290 -23966 -1274 -23932
rect -1132 -23966 -1116 -23932
rect -992 -23966 -976 -23932
rect -834 -23966 -818 -23932
rect -694 -23966 -678 -23932
rect -536 -23966 -520 -23932
rect -396 -23966 -380 -23932
rect -238 -23966 -222 -23932
rect -98 -23966 -82 -23932
rect 60 -23966 76 -23932
rect 200 -23966 216 -23932
rect 358 -23966 374 -23932
rect 498 -23966 514 -23932
rect 656 -23966 672 -23932
rect 796 -23966 812 -23932
rect -7890 -23968 -7830 -23967
rect -5854 -23968 -5794 -23967
rect -4832 -23968 -4772 -23967
rect -9405 -24017 -9371 -24001
rect -9405 -24609 -9371 -24593
rect -8387 -24017 -8353 -24001
rect -8387 -24609 -8353 -24593
rect -7369 -24017 -7335 -24001
rect -7369 -24609 -7335 -24593
rect -6351 -24017 -6317 -24001
rect -6351 -24609 -6317 -24593
rect -5333 -24017 -5299 -24001
rect -5333 -24609 -5299 -24593
rect -4315 -24017 -4281 -24001
rect -4315 -24609 -4281 -24593
rect -3297 -24017 -3263 -24001
rect -3297 -24609 -3263 -24593
rect -2412 -24016 -2378 -24000
rect -2412 -24608 -2378 -24592
rect -2114 -24016 -2080 -24000
rect -2114 -24608 -2080 -24592
rect -1816 -24016 -1782 -24000
rect -1816 -24608 -1782 -24592
rect -1518 -24016 -1484 -24000
rect -1518 -24608 -1484 -24592
rect -1220 -24016 -1186 -24000
rect -1220 -24608 -1186 -24592
rect -922 -24016 -888 -24000
rect -922 -24608 -888 -24592
rect -624 -24016 -590 -24000
rect -624 -24608 -590 -24592
rect -326 -24016 -292 -24000
rect -326 -24608 -292 -24592
rect -28 -24016 6 -24000
rect -28 -24608 6 -24592
rect 270 -24016 304 -24000
rect 270 -24608 304 -24592
rect 568 -24016 602 -24000
rect 568 -24608 602 -24592
rect 866 -24016 900 -24000
rect 2812 -24014 2828 -23980
rect 3384 -24014 3400 -23980
rect 3830 -24014 3846 -23980
rect 4402 -24014 4418 -23980
rect 4848 -24014 4864 -23980
rect 5420 -24014 5436 -23980
rect 5866 -24014 5882 -23980
rect 6438 -24014 6454 -23980
rect 6884 -24014 6900 -23980
rect 7456 -24014 7472 -23980
rect 7902 -24014 7918 -23980
rect 8474 -24014 8490 -23980
rect 8920 -24014 8936 -23980
rect 9492 -24014 9508 -23980
rect 9938 -24014 9954 -23980
rect 10510 -24014 10526 -23980
rect 10956 -24014 10972 -23980
rect 11528 -24014 11544 -23980
rect 11974 -24014 11990 -23980
rect 12546 -24014 12562 -23980
rect 12992 -24014 13008 -23980
rect 13564 -24014 13580 -23980
rect 14010 -24014 14026 -23980
rect 14582 -24014 14598 -23980
rect 15028 -24014 15044 -23980
rect 15600 -24014 15616 -23980
rect 16046 -24014 16062 -23980
rect 16618 -24014 16634 -23980
rect 17064 -24014 17080 -23980
rect 17636 -24014 17652 -23980
rect 18082 -24014 18098 -23980
rect 18654 -24014 18670 -23980
rect 19100 -24014 19116 -23980
rect 19672 -24014 19688 -23980
rect 20118 -24014 20134 -23980
rect 20690 -24014 20706 -23980
rect 21136 -24014 21152 -23980
rect 21708 -24014 21724 -23980
rect 22154 -24014 22170 -23980
rect 22726 -24014 22742 -23980
rect 9198 -24020 9258 -24014
rect 14270 -24020 14330 -24014
rect 15290 -24020 15350 -24014
rect 17326 -24020 17386 -24014
rect 866 -24608 900 -24592
rect 2580 -24064 2614 -24048
rect -7888 -24643 -7828 -24638
rect -6878 -24643 -6818 -24638
rect -5852 -24643 -5792 -24642
rect -4830 -24643 -4770 -24638
rect -9173 -24677 -9157 -24643
rect -8601 -24677 -8585 -24643
rect -8155 -24677 -8139 -24643
rect -7583 -24677 -7567 -24643
rect -7137 -24677 -7121 -24643
rect -6565 -24677 -6549 -24643
rect -6119 -24677 -6103 -24643
rect -5547 -24677 -5531 -24643
rect -5101 -24677 -5085 -24643
rect -4529 -24677 -4513 -24643
rect -4083 -24677 -4067 -24643
rect -3511 -24677 -3495 -24643
rect -2324 -24676 -2308 -24642
rect -2184 -24676 -2168 -24642
rect -2026 -24676 -2010 -24642
rect -1886 -24676 -1870 -24642
rect -1728 -24676 -1712 -24642
rect -1588 -24676 -1572 -24642
rect -1430 -24676 -1414 -24642
rect -1290 -24676 -1274 -24642
rect -1132 -24676 -1116 -24642
rect -992 -24676 -976 -24642
rect -834 -24676 -818 -24642
rect -694 -24676 -678 -24642
rect -536 -24676 -520 -24642
rect -396 -24676 -380 -24642
rect -238 -24676 -222 -24642
rect -98 -24676 -82 -24642
rect 60 -24676 76 -24642
rect 200 -24676 216 -24642
rect 358 -24676 374 -24642
rect 498 -24676 514 -24642
rect 656 -24676 672 -24642
rect 796 -24676 812 -24642
rect 2580 -24656 2614 -24640
rect 3598 -24064 3632 -24048
rect 3598 -24656 3632 -24640
rect 4616 -24064 4650 -24048
rect 4616 -24656 4650 -24640
rect 5634 -24064 5668 -24048
rect 5634 -24656 5668 -24640
rect 6652 -24064 6686 -24048
rect 6652 -24656 6686 -24640
rect 7670 -24064 7704 -24048
rect 7670 -24656 7704 -24640
rect 8688 -24064 8722 -24048
rect 8688 -24656 8722 -24640
rect 9706 -24064 9740 -24048
rect 9706 -24656 9740 -24640
rect 10724 -24064 10758 -24048
rect 10724 -24656 10758 -24640
rect 11742 -24064 11776 -24048
rect 11742 -24656 11776 -24640
rect 12760 -24064 12794 -24048
rect 12760 -24656 12794 -24640
rect 13778 -24064 13812 -24048
rect 13778 -24656 13812 -24640
rect 14796 -24064 14830 -24048
rect 14796 -24656 14830 -24640
rect 15814 -24064 15848 -24048
rect 15814 -24656 15848 -24640
rect 16832 -24064 16866 -24048
rect 16832 -24656 16866 -24640
rect 17850 -24064 17884 -24048
rect 17850 -24656 17884 -24640
rect 18868 -24064 18902 -24048
rect 18868 -24656 18902 -24640
rect 19886 -24064 19920 -24048
rect 19886 -24656 19920 -24640
rect 20904 -24064 20938 -24048
rect 20904 -24656 20938 -24640
rect 21922 -24064 21956 -24048
rect 21922 -24656 21956 -24640
rect 22940 -24064 22974 -24048
rect 22940 -24656 22974 -24640
rect 13254 -24690 13314 -24684
rect 2812 -24724 2828 -24690
rect 3384 -24724 3400 -24690
rect 3830 -24724 3846 -24690
rect 4402 -24724 4418 -24690
rect 4848 -24724 4864 -24690
rect 5420 -24724 5436 -24690
rect 5866 -24724 5882 -24690
rect 6438 -24724 6454 -24690
rect 6884 -24724 6900 -24690
rect 7456 -24724 7472 -24690
rect 7902 -24724 7918 -24690
rect 8474 -24724 8490 -24690
rect 8920 -24724 8936 -24690
rect 9492 -24724 9508 -24690
rect 9938 -24724 9954 -24690
rect 10510 -24724 10526 -24690
rect 10956 -24724 10972 -24690
rect 11528 -24724 11544 -24690
rect 11974 -24724 11990 -24690
rect 12546 -24724 12562 -24690
rect 12992 -24724 13008 -24690
rect 13564 -24724 13580 -24690
rect 14010 -24724 14026 -24690
rect 14582 -24724 14598 -24690
rect 15028 -24724 15044 -24690
rect 15600 -24724 15616 -24690
rect 16046 -24724 16062 -24690
rect 16618 -24724 16634 -24690
rect 17064 -24724 17080 -24690
rect 17636 -24724 17652 -24690
rect 18082 -24724 18098 -24690
rect 18654 -24724 18670 -24690
rect 19100 -24724 19116 -24690
rect 19672 -24724 19688 -24690
rect 20118 -24724 20134 -24690
rect 20690 -24724 20706 -24690
rect 21136 -24724 21152 -24690
rect 21708 -24724 21724 -24690
rect 22154 -24724 22170 -24690
rect 22726 -24724 22742 -24690
rect -9174 -25080 -9158 -25046
rect -8602 -25080 -8586 -25046
rect -8156 -25080 -8140 -25046
rect -7584 -25080 -7568 -25046
rect -7138 -25080 -7122 -25046
rect -6566 -25080 -6550 -25046
rect -6120 -25080 -6104 -25046
rect -5548 -25080 -5532 -25046
rect -5102 -25080 -5086 -25046
rect -4530 -25080 -4514 -25046
rect -4084 -25080 -4068 -25046
rect -3512 -25080 -3496 -25046
rect -2324 -25076 -2308 -25042
rect -2184 -25076 -2168 -25042
rect -2026 -25076 -2010 -25042
rect -1886 -25076 -1870 -25042
rect -1728 -25076 -1712 -25042
rect -1588 -25076 -1572 -25042
rect -1430 -25076 -1414 -25042
rect -1290 -25076 -1274 -25042
rect -1132 -25076 -1116 -25042
rect -992 -25076 -976 -25042
rect -834 -25076 -818 -25042
rect -694 -25076 -678 -25042
rect -536 -25076 -520 -25042
rect -396 -25076 -380 -25042
rect -238 -25076 -222 -25042
rect -98 -25076 -82 -25042
rect 60 -25076 76 -25042
rect 200 -25076 216 -25042
rect 358 -25076 374 -25042
rect 498 -25076 514 -25042
rect 656 -25076 672 -25042
rect 796 -25076 812 -25042
rect -9406 -25130 -9372 -25114
rect -9406 -25722 -9372 -25706
rect -8388 -25130 -8354 -25114
rect -8388 -25722 -8354 -25706
rect -7370 -25130 -7336 -25114
rect -7370 -25722 -7336 -25706
rect -6352 -25130 -6318 -25114
rect -6352 -25722 -6318 -25706
rect -5334 -25130 -5300 -25114
rect -5334 -25722 -5300 -25706
rect -4316 -25130 -4282 -25114
rect -4316 -25722 -4282 -25706
rect -3298 -25130 -3264 -25114
rect -3298 -25722 -3264 -25706
rect -2412 -25126 -2378 -25110
rect -2412 -25718 -2378 -25702
rect -2114 -25126 -2080 -25110
rect -2114 -25718 -2080 -25702
rect -1816 -25126 -1782 -25110
rect -1816 -25718 -1782 -25702
rect -1518 -25126 -1484 -25110
rect -1518 -25718 -1484 -25702
rect -1220 -25126 -1186 -25110
rect -1220 -25718 -1186 -25702
rect -922 -25126 -888 -25110
rect -922 -25718 -888 -25702
rect -624 -25126 -590 -25110
rect -624 -25718 -590 -25702
rect -326 -25126 -292 -25110
rect -326 -25718 -292 -25702
rect -28 -25126 6 -25110
rect -28 -25718 6 -25702
rect 270 -25126 304 -25110
rect 270 -25718 304 -25702
rect 568 -25126 602 -25110
rect 568 -25718 602 -25702
rect 866 -25126 900 -25110
rect 2812 -25246 2828 -25212
rect 3384 -25246 3400 -25212
rect 3830 -25246 3846 -25212
rect 4402 -25246 4418 -25212
rect 4848 -25246 4864 -25212
rect 5420 -25246 5436 -25212
rect 5866 -25246 5882 -25212
rect 6438 -25246 6454 -25212
rect 6884 -25246 6900 -25212
rect 7456 -25246 7472 -25212
rect 7902 -25246 7918 -25212
rect 8474 -25246 8490 -25212
rect 8920 -25246 8936 -25212
rect 9492 -25246 9508 -25212
rect 9938 -25246 9954 -25212
rect 10510 -25246 10526 -25212
rect 10956 -25246 10972 -25212
rect 11528 -25246 11544 -25212
rect 11974 -25246 11990 -25212
rect 12546 -25246 12562 -25212
rect 12992 -25246 13008 -25212
rect 13564 -25246 13580 -25212
rect 14010 -25246 14026 -25212
rect 14582 -25246 14598 -25212
rect 15028 -25246 15044 -25212
rect 15600 -25246 15616 -25212
rect 16046 -25246 16062 -25212
rect 16618 -25246 16634 -25212
rect 17064 -25246 17080 -25212
rect 17636 -25246 17652 -25212
rect 18082 -25246 18098 -25212
rect 18654 -25246 18670 -25212
rect 19100 -25246 19116 -25212
rect 19672 -25246 19688 -25212
rect 20118 -25246 20134 -25212
rect 20690 -25246 20706 -25212
rect 21136 -25246 21152 -25212
rect 21708 -25246 21724 -25212
rect 22154 -25246 22170 -25212
rect 22726 -25246 22742 -25212
rect 3066 -25250 3126 -25246
rect 4088 -25250 4148 -25246
rect 5114 -25250 5174 -25246
rect 6130 -25250 6190 -25246
rect 7144 -25250 7204 -25246
rect 8174 -25256 8234 -25246
rect 9190 -25256 9250 -25246
rect 10194 -25250 10254 -25246
rect 11224 -25256 11284 -25246
rect 12244 -25250 12304 -25246
rect 13254 -25250 13314 -25246
rect 14278 -25256 14338 -25246
rect 16304 -25250 16364 -25246
rect 17324 -25256 17384 -25246
rect 18348 -25250 18408 -25246
rect 21392 -25250 21452 -25246
rect 22414 -25248 22474 -25246
rect 866 -25718 900 -25702
rect 2580 -25296 2614 -25280
rect -9174 -25790 -9158 -25756
rect -8602 -25790 -8586 -25756
rect -8156 -25790 -8140 -25756
rect -7584 -25790 -7568 -25756
rect -7138 -25790 -7122 -25756
rect -6566 -25790 -6550 -25756
rect -6120 -25790 -6104 -25756
rect -5548 -25790 -5532 -25756
rect -5102 -25790 -5086 -25756
rect -4530 -25790 -4514 -25756
rect -4084 -25790 -4068 -25756
rect -3512 -25790 -3496 -25756
rect -2324 -25786 -2308 -25752
rect -2184 -25786 -2168 -25752
rect -2026 -25786 -2010 -25752
rect -1886 -25786 -1870 -25752
rect -1728 -25786 -1712 -25752
rect -1588 -25786 -1572 -25752
rect -1430 -25786 -1414 -25752
rect -1290 -25786 -1274 -25752
rect -1132 -25786 -1116 -25752
rect -992 -25786 -976 -25752
rect -834 -25786 -818 -25752
rect -694 -25786 -678 -25752
rect -536 -25786 -520 -25752
rect -396 -25786 -380 -25752
rect -238 -25786 -222 -25752
rect -98 -25786 -82 -25752
rect 60 -25786 76 -25752
rect 200 -25786 216 -25752
rect 358 -25786 374 -25752
rect 498 -25786 514 -25752
rect 656 -25786 672 -25752
rect 796 -25786 812 -25752
rect 3598 -25296 3632 -25280
rect 3582 -25872 3598 -25832
rect 4616 -25296 4650 -25280
rect 3632 -25872 3642 -25832
rect 5634 -25296 5668 -25280
rect 6652 -25296 6686 -25280
rect 7670 -25296 7704 -25280
rect 7656 -25872 7670 -25828
rect 8688 -25296 8722 -25280
rect 7704 -25872 7716 -25828
rect 9706 -25296 9740 -25280
rect 10724 -25296 10758 -25280
rect 11742 -25296 11776 -25280
rect 12760 -25296 12794 -25280
rect 13778 -25296 13812 -25280
rect 13764 -25872 13778 -25826
rect 14796 -25296 14830 -25280
rect 13812 -25872 13824 -25826
rect 15814 -25296 15848 -25280
rect 16832 -25296 16866 -25280
rect 17850 -25296 17884 -25280
rect 17836 -25872 17850 -25836
rect 18868 -25296 18902 -25280
rect 17884 -25872 17896 -25836
rect 19886 -25296 19920 -25280
rect 20904 -25296 20938 -25280
rect 21922 -25296 21956 -25280
rect 21906 -25872 21922 -25834
rect 22940 -25296 22974 -25280
rect 21956 -25872 21966 -25834
rect 2580 -25888 2614 -25872
rect 4616 -25888 4650 -25872
rect 6652 -25888 6686 -25872
rect 8688 -25888 8722 -25872
rect 10724 -25888 10758 -25872
rect 12760 -25888 12794 -25872
rect 14796 -25888 14830 -25872
rect 16832 -25888 16866 -25872
rect 18868 -25888 18902 -25872
rect 20904 -25888 20938 -25872
rect 22940 -25888 22974 -25872
rect 9186 -25922 9246 -25920
rect 15298 -25922 15358 -25920
rect 20384 -25922 20444 -25920
rect 2812 -25956 2828 -25922
rect 3384 -25956 3400 -25922
rect 3830 -25956 3846 -25922
rect 4402 -25956 4418 -25922
rect 4848 -25956 4864 -25922
rect 5420 -25956 5436 -25922
rect 5866 -25956 5882 -25922
rect 6438 -25956 6454 -25922
rect 6884 -25956 6900 -25922
rect 7456 -25956 7472 -25922
rect 7902 -25956 7918 -25922
rect 8474 -25956 8490 -25922
rect 8920 -25956 8936 -25922
rect 9492 -25956 9508 -25922
rect 9938 -25956 9954 -25922
rect 10510 -25956 10526 -25922
rect 10956 -25956 10972 -25922
rect 11528 -25956 11544 -25922
rect 11974 -25956 11990 -25922
rect 12546 -25956 12562 -25922
rect 12992 -25956 13008 -25922
rect 13564 -25956 13580 -25922
rect 14010 -25956 14026 -25922
rect 14582 -25956 14598 -25922
rect 15028 -25956 15044 -25922
rect 15600 -25956 15616 -25922
rect 16046 -25956 16062 -25922
rect 16618 -25956 16634 -25922
rect 17064 -25956 17080 -25922
rect 17636 -25956 17652 -25922
rect 18082 -25956 18098 -25922
rect 18654 -25956 18670 -25922
rect 19100 -25956 19116 -25922
rect 19672 -25956 19688 -25922
rect 20118 -25956 20134 -25922
rect 20690 -25956 20706 -25922
rect 21136 -25956 21152 -25922
rect 21708 -25956 21724 -25922
rect 22154 -25956 22170 -25922
rect 22726 -25956 22742 -25922
rect -12322 -27222 -12222 -27060
rect 24822 -27222 24922 -27060
<< viali >>
rect 478 1622 540 1722
rect 540 1622 24660 1722
rect 24660 1622 24722 1722
rect 378 -8262 478 1102
rect 3720 -4643 3784 -4609
rect 3938 -4643 4002 -4609
rect 4156 -4643 4220 -4609
rect 4374 -4643 4438 -4609
rect 4592 -4643 4656 -4609
rect 4810 -4643 4874 -4609
rect 5028 -4643 5092 -4609
rect 5246 -4643 5310 -4609
rect 5464 -4643 5528 -4609
rect 5682 -4643 5746 -4609
rect 3626 -5078 3660 -4702
rect 3844 -5078 3878 -4702
rect 4062 -5078 4096 -4702
rect 4280 -5078 4314 -4702
rect 4498 -5078 4532 -4702
rect 4716 -5078 4750 -4702
rect 4934 -5078 4968 -4702
rect 5152 -5078 5186 -4702
rect 5370 -5078 5404 -4702
rect 5588 -5078 5622 -4702
rect 5806 -5078 5840 -4702
rect 3720 -5171 3784 -5137
rect 3938 -5171 4002 -5137
rect 4156 -5171 4220 -5137
rect 4374 -5171 4438 -5137
rect 4592 -5171 4656 -5137
rect 4810 -5171 4874 -5137
rect 5028 -5171 5092 -5137
rect 5246 -5171 5310 -5137
rect 5464 -5171 5528 -5137
rect 5682 -5171 5746 -5137
rect 3720 -5581 3784 -5547
rect 3938 -5581 4002 -5547
rect 4156 -5581 4220 -5547
rect 4374 -5581 4438 -5547
rect 4592 -5581 4656 -5547
rect 4810 -5581 4874 -5547
rect 5028 -5581 5092 -5547
rect 5246 -5581 5310 -5547
rect 5464 -5581 5528 -5547
rect 5682 -5581 5746 -5547
rect 3626 -6016 3660 -5640
rect 3844 -6016 3878 -5640
rect 4062 -6016 4096 -5640
rect 4280 -6016 4314 -5640
rect 4498 -6016 4532 -5640
rect 4716 -6016 4750 -5640
rect 4934 -6016 4968 -5640
rect 5152 -6016 5186 -5640
rect 5370 -6016 5404 -5640
rect 5588 -6016 5622 -5640
rect 5806 -6016 5840 -5640
rect 3720 -6109 3784 -6075
rect 3938 -6109 4002 -6075
rect 4156 -6109 4220 -6075
rect 4374 -6109 4438 -6075
rect 4592 -6109 4656 -6075
rect 4810 -6109 4874 -6075
rect 5028 -6109 5092 -6075
rect 5246 -6109 5310 -6075
rect 5464 -6109 5528 -6075
rect 5682 -6109 5746 -6075
rect 3720 -6519 3784 -6485
rect 3938 -6519 4002 -6485
rect 4156 -6519 4220 -6485
rect 4374 -6519 4438 -6485
rect 4592 -6519 4656 -6485
rect 4810 -6519 4874 -6485
rect 5028 -6519 5092 -6485
rect 5246 -6519 5310 -6485
rect 5464 -6519 5528 -6485
rect 5682 -6519 5746 -6485
rect 3626 -6954 3660 -6578
rect 3844 -6954 3878 -6578
rect 4062 -6954 4096 -6578
rect 4280 -6954 4314 -6578
rect 4498 -6954 4532 -6578
rect 4716 -6954 4750 -6578
rect 4934 -6954 4968 -6578
rect 5152 -6954 5186 -6578
rect 5370 -6954 5404 -6578
rect 5588 -6954 5622 -6578
rect 5806 -6954 5840 -6578
rect 3720 -7047 3784 -7013
rect 3938 -7047 4002 -7013
rect 4156 -7047 4220 -7013
rect 4374 -7047 4438 -7013
rect 4592 -7047 4656 -7013
rect 4810 -7047 4874 -7013
rect 5028 -7047 5092 -7013
rect 5246 -7047 5310 -7013
rect 5464 -7047 5528 -7013
rect 5682 -7047 5746 -7013
rect 3720 -7457 3784 -7423
rect 3938 -7457 4002 -7423
rect 4156 -7457 4220 -7423
rect 4374 -7457 4438 -7423
rect 4592 -7457 4656 -7423
rect 4810 -7457 4874 -7423
rect 5028 -7457 5092 -7423
rect 5246 -7457 5310 -7423
rect 5464 -7457 5528 -7423
rect 5682 -7457 5746 -7423
rect 3626 -7892 3660 -7516
rect 3844 -7892 3878 -7516
rect 4062 -7892 4096 -7516
rect 4280 -7892 4314 -7516
rect 4498 -7892 4532 -7516
rect 4716 -7892 4750 -7516
rect 4934 -7892 4968 -7516
rect 5152 -7892 5186 -7516
rect 5370 -7892 5404 -7516
rect 5588 -7892 5622 -7516
rect 5806 -7892 5840 -7516
rect 3720 -7985 3784 -7951
rect 3938 -7985 4002 -7951
rect 4156 -7985 4220 -7951
rect 4374 -7985 4438 -7951
rect 4592 -7985 4656 -7951
rect 4810 -7985 4874 -7951
rect 5028 -7985 5092 -7951
rect 5246 -7985 5310 -7951
rect 5464 -7985 5528 -7951
rect 5682 -7985 5746 -7951
rect 24722 -8262 24822 1102
rect 478 -8882 540 -8782
rect 540 -8882 24660 -8782
rect 24660 -8882 24722 -8782
rect -12222 -11278 -12160 -11178
rect -12160 -11278 24760 -11178
rect 24760 -11278 24822 -11178
rect 2876 -11680 3340 -11646
rect 3894 -11680 4358 -11646
rect 4912 -11680 5376 -11646
rect 5930 -11680 6394 -11646
rect 6948 -11680 7412 -11646
rect 7966 -11680 8430 -11646
rect 8984 -11680 9448 -11646
rect 10002 -11680 10466 -11646
rect 11020 -11680 11484 -11646
rect 12038 -11680 12502 -11646
rect 13056 -11680 13520 -11646
rect 14074 -11680 14538 -11646
rect 15092 -11680 15556 -11646
rect 16110 -11680 16574 -11646
rect 17128 -11680 17592 -11646
rect 18146 -11680 18610 -11646
rect 19164 -11680 19628 -11646
rect 20182 -11680 20646 -11646
rect 21200 -11680 21664 -11646
rect 22218 -11680 22682 -11646
rect -12322 -26330 -12222 -12070
rect 2582 -12306 2616 -11730
rect 3600 -12306 3634 -11730
rect 4618 -12306 4652 -11730
rect 5636 -12306 5670 -11730
rect 6654 -12306 6688 -11730
rect 7672 -12306 7706 -11730
rect 8690 -12306 8724 -11730
rect 9708 -12306 9742 -11730
rect 10726 -12306 10760 -11730
rect 11744 -12306 11778 -11730
rect 12762 -12306 12796 -11730
rect 13780 -12306 13814 -11730
rect 14798 -12306 14832 -11730
rect 15816 -12306 15850 -11730
rect 16834 -12306 16868 -11730
rect 17852 -12306 17886 -11730
rect 18870 -12306 18904 -11730
rect 19888 -12306 19922 -11730
rect 20906 -12306 20940 -11730
rect 21924 -12306 21958 -11730
rect 22942 -12306 22976 -11730
rect 2876 -12390 3340 -12356
rect 3894 -12390 4358 -12356
rect 4912 -12390 5376 -12356
rect 5930 -12390 6394 -12356
rect 6948 -12390 7412 -12356
rect 7966 -12390 8430 -12356
rect 8984 -12390 9448 -12356
rect 10002 -12390 10466 -12356
rect 11020 -12390 11484 -12356
rect 12038 -12390 12502 -12356
rect 13056 -12390 13520 -12356
rect 14074 -12390 14538 -12356
rect 15092 -12390 15556 -12356
rect 16110 -12390 16574 -12356
rect 17128 -12390 17592 -12356
rect 18146 -12390 18610 -12356
rect 19164 -12390 19628 -12356
rect 20182 -12390 20646 -12356
rect 21200 -12390 21664 -12356
rect 22218 -12390 22682 -12356
rect -8890 -12474 -8426 -12440
rect -7872 -12474 -7408 -12440
rect -6854 -12474 -6390 -12440
rect -5836 -12474 -5372 -12440
rect -4818 -12474 -4354 -12440
rect -3800 -12474 -3336 -12440
rect -2782 -12474 -2318 -12440
rect -1764 -12474 -1300 -12440
rect -746 -12474 -282 -12440
rect -9184 -13100 -9150 -12524
rect -8166 -13100 -8132 -12524
rect -7148 -13100 -7114 -12524
rect -6130 -13100 -6096 -12524
rect -5112 -13100 -5078 -12524
rect -4094 -13100 -4060 -12524
rect -3076 -13100 -3042 -12524
rect -2058 -13100 -2024 -12524
rect -1040 -13100 -1006 -12524
rect -22 -13100 12 -12524
rect 2876 -12914 3340 -12880
rect 3894 -12914 4358 -12880
rect 4912 -12914 5376 -12880
rect 5930 -12914 6394 -12880
rect 6948 -12914 7412 -12880
rect 7966 -12914 8430 -12880
rect 8984 -12914 9448 -12880
rect 10002 -12914 10466 -12880
rect 11020 -12914 11484 -12880
rect 12038 -12914 12502 -12880
rect 13056 -12914 13520 -12880
rect 14074 -12914 14538 -12880
rect 15092 -12914 15556 -12880
rect 16110 -12914 16574 -12880
rect 17128 -12914 17592 -12880
rect 18146 -12914 18610 -12880
rect 19164 -12914 19628 -12880
rect 20182 -12914 20646 -12880
rect 21200 -12914 21664 -12880
rect 22218 -12914 22682 -12880
rect -8890 -13184 -8426 -13150
rect -7872 -13184 -7408 -13150
rect -6854 -13184 -6390 -13150
rect -5836 -13184 -5372 -13150
rect -4818 -13184 -4354 -13150
rect -3800 -13184 -3336 -13150
rect -2782 -13184 -2318 -13150
rect -1764 -13184 -1300 -13150
rect -746 -13184 -282 -13150
rect -8890 -13292 -8426 -13258
rect -7872 -13292 -7408 -13258
rect -6854 -13292 -6390 -13258
rect -5836 -13292 -5372 -13258
rect -4818 -13292 -4354 -13258
rect -3800 -13292 -3336 -13258
rect -2782 -13292 -2318 -13258
rect -1764 -13292 -1300 -13258
rect -746 -13292 -282 -13258
rect -9184 -13918 -9150 -13342
rect -8166 -13918 -8132 -13342
rect -7148 -13918 -7114 -13342
rect -6130 -13918 -6096 -13342
rect -5112 -13918 -5078 -13342
rect -4094 -13918 -4060 -13342
rect -3076 -13918 -3042 -13342
rect -2058 -13918 -2024 -13342
rect -1040 -13918 -1006 -13342
rect -22 -13918 12 -13342
rect 2582 -13540 2616 -12964
rect 3600 -13540 3634 -12964
rect 4618 -13540 4652 -12964
rect 5636 -13540 5670 -12964
rect 6654 -13540 6688 -12964
rect 7672 -13540 7706 -12964
rect 8690 -13540 8724 -12964
rect 9708 -13540 9742 -12964
rect 10726 -13540 10760 -12964
rect 11744 -13540 11778 -12964
rect 12762 -13540 12796 -12964
rect 13780 -13540 13814 -12964
rect 14798 -13540 14832 -12964
rect 15816 -13540 15850 -12964
rect 16834 -13540 16868 -12964
rect 17852 -13540 17886 -12964
rect 18870 -13540 18904 -12964
rect 19888 -13540 19922 -12964
rect 20906 -13540 20940 -12964
rect 21924 -13540 21958 -12964
rect 22942 -13540 22976 -12964
rect 2876 -13624 3340 -13590
rect 3894 -13624 4358 -13590
rect 4912 -13624 5376 -13590
rect 5930 -13624 6394 -13590
rect 6948 -13624 7412 -13590
rect 7966 -13624 8430 -13590
rect 8984 -13624 9448 -13590
rect 10002 -13624 10466 -13590
rect 11020 -13624 11484 -13590
rect 12038 -13624 12502 -13590
rect 13056 -13624 13520 -13590
rect 14074 -13624 14538 -13590
rect 15092 -13624 15556 -13590
rect 16110 -13624 16574 -13590
rect 17128 -13624 17592 -13590
rect 18146 -13624 18610 -13590
rect 19164 -13624 19628 -13590
rect 20182 -13624 20646 -13590
rect 21200 -13624 21664 -13590
rect 22218 -13624 22682 -13590
rect -8890 -14002 -8426 -13968
rect -7872 -14002 -7408 -13968
rect -6854 -14002 -6390 -13968
rect -5836 -14002 -5372 -13968
rect -4818 -14002 -4354 -13968
rect -3800 -14002 -3336 -13968
rect -2782 -14002 -2318 -13968
rect -1764 -14002 -1300 -13968
rect -746 -14002 -282 -13968
rect -8890 -14110 -8426 -14076
rect -7872 -14110 -7408 -14076
rect -6854 -14110 -6390 -14076
rect -5836 -14110 -5372 -14076
rect -4818 -14110 -4354 -14076
rect -3800 -14110 -3336 -14076
rect -2782 -14110 -2318 -14076
rect -1764 -14110 -1300 -14076
rect -746 -14110 -282 -14076
rect -9184 -14736 -9150 -14160
rect -8166 -14736 -8132 -14160
rect -7148 -14736 -7114 -14160
rect -6130 -14736 -6096 -14160
rect -5112 -14736 -5078 -14160
rect -4094 -14736 -4060 -14160
rect -3076 -14736 -3042 -14160
rect -2058 -14736 -2024 -14160
rect -1040 -14736 -1006 -14160
rect 2876 -14146 3340 -14112
rect 3894 -14146 4358 -14112
rect 4912 -14146 5376 -14112
rect 5930 -14146 6394 -14112
rect 6948 -14146 7412 -14112
rect 7966 -14146 8430 -14112
rect 8984 -14146 9448 -14112
rect 10002 -14146 10466 -14112
rect 11020 -14146 11484 -14112
rect 12038 -14146 12502 -14112
rect 13056 -14146 13520 -14112
rect 14074 -14146 14538 -14112
rect 15092 -14146 15556 -14112
rect 16110 -14146 16574 -14112
rect 17128 -14146 17592 -14112
rect 18146 -14146 18610 -14112
rect 19164 -14146 19628 -14112
rect 20182 -14146 20646 -14112
rect 21200 -14146 21664 -14112
rect 22218 -14146 22682 -14112
rect -22 -14736 12 -14160
rect 2582 -14772 2616 -14196
rect -8890 -14820 -8426 -14786
rect -7872 -14820 -7408 -14786
rect -6854 -14820 -6390 -14786
rect -5836 -14820 -5372 -14786
rect -4818 -14820 -4354 -14786
rect -3800 -14820 -3336 -14786
rect -2782 -14820 -2318 -14786
rect -1764 -14820 -1300 -14786
rect -746 -14820 -282 -14786
rect 3600 -14772 3634 -14196
rect 4618 -14772 4652 -14196
rect 5636 -14772 5670 -14196
rect 6654 -14772 6688 -14196
rect 7672 -14772 7706 -14196
rect 8690 -14772 8724 -14196
rect 9708 -14772 9742 -14196
rect 10726 -14772 10760 -14196
rect 11744 -14772 11778 -14196
rect 12762 -14772 12796 -14196
rect 13780 -14772 13814 -14196
rect 14798 -14772 14832 -14196
rect 15816 -14772 15850 -14196
rect 16834 -14772 16868 -14196
rect 17852 -14772 17886 -14196
rect 18870 -14772 18904 -14196
rect 19888 -14772 19922 -14196
rect 20906 -14772 20940 -14196
rect 21924 -14772 21958 -14196
rect 22942 -14772 22976 -14196
rect 2876 -14856 3340 -14822
rect 3894 -14856 4358 -14822
rect 4912 -14856 5376 -14822
rect 5930 -14856 6394 -14822
rect 6948 -14856 7412 -14822
rect 7966 -14856 8430 -14822
rect 8984 -14856 9448 -14822
rect 10002 -14856 10466 -14822
rect 11020 -14856 11484 -14822
rect 12038 -14856 12502 -14822
rect 13056 -14856 13520 -14822
rect 14074 -14856 14538 -14822
rect 15092 -14856 15556 -14822
rect 16110 -14856 16574 -14822
rect 17128 -14854 17592 -14822
rect 17128 -14856 17318 -14854
rect 17378 -14856 17592 -14854
rect 18146 -14850 18610 -14822
rect 18146 -14856 18352 -14850
rect 18412 -14856 18610 -14850
rect 19164 -14856 19628 -14822
rect 20182 -14856 20646 -14822
rect 21200 -14856 21664 -14822
rect 22218 -14856 22682 -14822
rect -8890 -14928 -8426 -14894
rect -7872 -14928 -7408 -14894
rect -6854 -14928 -6390 -14894
rect -5836 -14928 -5372 -14894
rect -4818 -14928 -4354 -14894
rect -3800 -14928 -3336 -14894
rect -2782 -14928 -2318 -14894
rect -1764 -14928 -1300 -14894
rect -746 -14928 -282 -14894
rect -9184 -15554 -9150 -14978
rect -8166 -15554 -8132 -14978
rect -7148 -15554 -7114 -14978
rect -6130 -15554 -6096 -14978
rect -5112 -15554 -5078 -14978
rect -4094 -15554 -4060 -14978
rect -3076 -15554 -3042 -14978
rect -2058 -15554 -2024 -14978
rect -1040 -15554 -1006 -14978
rect -22 -15554 12 -14978
rect 2874 -15380 3338 -15346
rect 3892 -15380 4356 -15346
rect 4910 -15380 5374 -15346
rect 5928 -15380 6392 -15346
rect 6946 -15380 7410 -15346
rect 7964 -15380 8428 -15346
rect 8982 -15380 9446 -15346
rect 10000 -15380 10464 -15346
rect 11018 -15380 11482 -15346
rect 12036 -15380 12500 -15346
rect 13054 -15380 13518 -15346
rect 14072 -15380 14536 -15346
rect 15090 -15380 15554 -15346
rect 16108 -15380 16572 -15346
rect 17126 -15380 17590 -15346
rect 18144 -15380 18608 -15346
rect 19162 -15380 19626 -15346
rect 20180 -15380 20644 -15346
rect 21198 -15380 21662 -15346
rect 22216 -15380 22680 -15346
rect -8890 -15638 -8426 -15604
rect -7872 -15638 -7408 -15604
rect -6854 -15638 -6390 -15604
rect -5836 -15638 -5372 -15604
rect -4818 -15638 -4354 -15604
rect -3800 -15638 -3336 -15604
rect -2782 -15638 -2318 -15604
rect -1764 -15638 -1300 -15604
rect -746 -15638 -282 -15604
rect -8890 -15746 -8426 -15712
rect -7872 -15746 -7408 -15712
rect -6854 -15746 -6390 -15712
rect -5836 -15746 -5372 -15712
rect -4818 -15746 -4354 -15712
rect -3800 -15746 -3336 -15712
rect -2782 -15746 -2318 -15712
rect -1764 -15746 -1300 -15712
rect -746 -15746 -282 -15712
rect -9184 -16372 -9150 -15796
rect -8166 -16372 -8132 -15796
rect -7148 -16372 -7114 -15796
rect -6130 -16372 -6096 -15796
rect -5112 -16372 -5078 -15796
rect -4094 -16372 -4060 -15796
rect -3076 -16372 -3042 -15796
rect -2058 -16372 -2024 -15796
rect -1040 -16372 -1006 -15796
rect -22 -16372 12 -15796
rect 2580 -16006 2614 -15430
rect 3598 -16006 3632 -15430
rect 4616 -16006 4650 -15430
rect 5634 -16006 5668 -15430
rect 6652 -16006 6686 -15430
rect 7670 -16006 7704 -15430
rect 8688 -16006 8722 -15430
rect 9706 -16006 9740 -15430
rect 10724 -16006 10758 -15430
rect 11742 -16006 11776 -15430
rect 12760 -16006 12794 -15430
rect 13778 -16006 13812 -15430
rect 14796 -16006 14830 -15430
rect 15814 -16006 15848 -15430
rect 16832 -16006 16866 -15430
rect 17850 -16006 17884 -15430
rect 18868 -16006 18902 -15430
rect 19886 -16006 19920 -15430
rect 20904 -16006 20938 -15430
rect 21922 -16006 21956 -15430
rect 22940 -16006 22974 -15430
rect 2874 -16090 3338 -16056
rect 3892 -16090 4356 -16056
rect 4910 -16090 5374 -16056
rect 5928 -16090 6392 -16056
rect 6946 -16090 7410 -16056
rect 7964 -16090 8428 -16056
rect 8982 -16090 9446 -16056
rect 10000 -16090 10464 -16056
rect 11018 -16090 11482 -16056
rect 12036 -16090 12500 -16056
rect 13054 -16090 13518 -16056
rect 14072 -16090 14536 -16056
rect 15090 -16090 15554 -16056
rect 16108 -16090 16572 -16056
rect 17126 -16090 17590 -16056
rect 18144 -16090 18608 -16056
rect 19162 -16090 19626 -16056
rect 20180 -16090 20644 -16056
rect 21198 -16090 21662 -16056
rect 22216 -16090 22680 -16056
rect -8890 -16456 -8426 -16422
rect -7872 -16456 -7408 -16422
rect -6854 -16456 -6390 -16422
rect -5836 -16456 -5372 -16422
rect -4818 -16456 -4354 -16422
rect -3800 -16456 -3336 -16422
rect -2782 -16456 -2318 -16422
rect -1764 -16456 -1300 -16422
rect -746 -16456 -282 -16422
rect -8890 -16564 -8426 -16530
rect -7872 -16564 -7408 -16530
rect -6854 -16564 -6390 -16530
rect -5836 -16564 -5372 -16530
rect -4818 -16564 -4354 -16530
rect -3800 -16564 -3336 -16530
rect -2782 -16564 -2318 -16530
rect -1764 -16564 -1300 -16530
rect -746 -16564 -282 -16530
rect -9184 -17190 -9150 -16614
rect -8166 -17190 -8132 -16614
rect -7148 -17190 -7114 -16614
rect -6130 -17190 -6096 -16614
rect -5112 -17190 -5078 -16614
rect -4094 -17190 -4060 -16614
rect -3076 -17190 -3042 -16614
rect -2058 -17190 -2024 -16614
rect -1040 -17190 -1006 -16614
rect 2874 -16614 3338 -16580
rect 3892 -16614 4356 -16580
rect 4910 -16614 5374 -16580
rect 5928 -16614 6392 -16580
rect 6946 -16614 7410 -16580
rect 7964 -16614 8428 -16580
rect 8982 -16614 9446 -16580
rect 10000 -16614 10464 -16580
rect 11018 -16614 11482 -16580
rect 12036 -16614 12500 -16580
rect 13054 -16614 13518 -16580
rect 14072 -16614 14536 -16580
rect 15090 -16614 15554 -16580
rect 16108 -16614 16572 -16580
rect 17126 -16614 17590 -16580
rect 18144 -16614 18608 -16580
rect 19162 -16614 19626 -16580
rect 20180 -16614 20644 -16580
rect 21198 -16614 21662 -16580
rect 22216 -16614 22680 -16580
rect -22 -17190 12 -16614
rect 2580 -17240 2614 -16664
rect -8890 -17274 -8426 -17240
rect -7872 -17274 -7408 -17240
rect -6854 -17274 -6390 -17240
rect -5836 -17274 -5372 -17240
rect -4818 -17274 -4354 -17240
rect -3800 -17274 -3336 -17240
rect -2782 -17274 -2318 -17240
rect -1764 -17274 -1300 -17240
rect -746 -17274 -282 -17240
rect 3598 -17240 3632 -16664
rect 4616 -17240 4650 -16664
rect 5634 -17240 5668 -16664
rect 6652 -17240 6686 -16664
rect 7670 -17240 7704 -16664
rect 8688 -17240 8722 -16664
rect 9706 -17240 9740 -16664
rect 10724 -17240 10758 -16664
rect 11742 -17240 11776 -16664
rect 12760 -17240 12794 -16664
rect 13778 -17240 13812 -16664
rect 14796 -17240 14830 -16664
rect 15814 -17240 15848 -16664
rect 16832 -17240 16866 -16664
rect 17850 -17240 17884 -16664
rect 18868 -17240 18902 -16664
rect 19886 -17240 19920 -16664
rect 20904 -17240 20938 -16664
rect 21922 -17240 21956 -16664
rect 22940 -17240 22974 -16664
rect 2874 -17324 3338 -17290
rect 3892 -17324 4356 -17290
rect 4910 -17324 5374 -17290
rect 5928 -17324 6392 -17290
rect 6946 -17324 7410 -17290
rect 7964 -17324 8428 -17290
rect 8982 -17324 9446 -17290
rect 10000 -17324 10464 -17290
rect 11018 -17324 11482 -17290
rect 12036 -17324 12500 -17290
rect 13054 -17324 13518 -17290
rect 14072 -17324 14536 -17290
rect 15090 -17324 15554 -17290
rect 16108 -17324 16572 -17290
rect 17126 -17324 17590 -17290
rect 18144 -17324 18608 -17290
rect 19162 -17324 19626 -17290
rect 20180 -17324 20644 -17290
rect 21198 -17294 21662 -17290
rect 21198 -17324 21392 -17294
rect 21452 -17324 21662 -17294
rect 22216 -17324 22680 -17290
rect -8890 -17382 -8426 -17348
rect -7872 -17382 -7408 -17348
rect -6854 -17382 -6390 -17348
rect -5836 -17382 -5372 -17348
rect -4818 -17382 -4354 -17348
rect -3800 -17382 -3336 -17348
rect -2782 -17382 -2318 -17348
rect -1764 -17382 -1300 -17348
rect -746 -17382 -282 -17348
rect -9184 -18008 -9150 -17432
rect -8166 -18008 -8132 -17432
rect -7148 -18008 -7114 -17432
rect -6130 -18008 -6096 -17432
rect -5112 -18008 -5078 -17432
rect -4094 -18008 -4060 -17432
rect -3076 -18008 -3042 -17432
rect -2058 -18008 -2024 -17432
rect -1040 -18008 -1006 -17432
rect -22 -18008 12 -17432
rect 2874 -17846 3338 -17812
rect 3892 -17846 4356 -17812
rect 4910 -17846 5374 -17812
rect 5928 -17846 6392 -17812
rect 6946 -17846 7410 -17812
rect 7964 -17846 8428 -17812
rect 8982 -17846 9446 -17812
rect 10000 -17846 10464 -17812
rect 11018 -17846 11482 -17812
rect 12036 -17846 12500 -17812
rect 13054 -17846 13518 -17812
rect 14072 -17846 14536 -17812
rect 15090 -17846 15554 -17812
rect 16108 -17846 16572 -17812
rect 17126 -17846 17590 -17812
rect 18144 -17846 18608 -17812
rect 19162 -17846 19626 -17812
rect 20180 -17846 20644 -17812
rect 21198 -17846 21662 -17812
rect 22216 -17846 22680 -17812
rect -8890 -18092 -8426 -18058
rect -7872 -18092 -7408 -18058
rect -6854 -18092 -6390 -18058
rect -5836 -18092 -5372 -18058
rect -4818 -18092 -4354 -18058
rect -3800 -18092 -3336 -18058
rect -2782 -18092 -2318 -18058
rect -1764 -18092 -1300 -18058
rect -746 -18092 -282 -18058
rect -8890 -18200 -8426 -18166
rect -7872 -18200 -7408 -18166
rect -6854 -18200 -6390 -18166
rect -5836 -18200 -5372 -18166
rect -4818 -18200 -4354 -18166
rect -3800 -18200 -3336 -18166
rect -2782 -18200 -2318 -18166
rect -1764 -18200 -1300 -18166
rect -746 -18200 -282 -18166
rect -9184 -18826 -9150 -18250
rect -8166 -18826 -8132 -18250
rect -7148 -18826 -7114 -18250
rect -6130 -18826 -6096 -18250
rect -5112 -18826 -5078 -18250
rect -4094 -18826 -4060 -18250
rect -3076 -18826 -3042 -18250
rect -2058 -18826 -2024 -18250
rect -1040 -18826 -1006 -18250
rect -22 -18826 12 -18250
rect 2580 -18472 2614 -17896
rect 3598 -18472 3632 -17896
rect 4616 -18472 4650 -17896
rect 5634 -18472 5668 -17896
rect 6652 -18472 6686 -17896
rect 7670 -18472 7704 -17896
rect 8688 -18472 8722 -17896
rect 9706 -18472 9740 -17896
rect 10724 -18472 10758 -17896
rect 11742 -18472 11776 -17896
rect 12760 -18472 12794 -17896
rect 13778 -18472 13812 -17896
rect 14796 -18472 14830 -17896
rect 15814 -18472 15848 -17896
rect 16832 -18472 16866 -17896
rect 17850 -18472 17884 -17896
rect 18868 -18472 18902 -17896
rect 19886 -18472 19920 -17896
rect 20904 -18472 20938 -17896
rect 21922 -18472 21956 -17896
rect 22940 -18472 22974 -17896
rect 2874 -18556 3338 -18522
rect 3892 -18556 4356 -18522
rect 4910 -18556 5374 -18522
rect 5928 -18556 6392 -18522
rect 6946 -18556 7410 -18522
rect 7964 -18556 8428 -18522
rect 8982 -18556 9446 -18522
rect 10000 -18556 10464 -18522
rect 11018 -18556 11482 -18522
rect 12036 -18556 12500 -18522
rect 13054 -18556 13518 -18522
rect 14072 -18556 14536 -18522
rect 15090 -18556 15554 -18522
rect 16108 -18556 16572 -18522
rect 17126 -18556 17590 -18522
rect 18144 -18556 18608 -18522
rect 19162 -18556 19626 -18522
rect 20180 -18556 20644 -18522
rect 21198 -18556 21662 -18522
rect 22216 -18556 22680 -18522
rect -8890 -18910 -8426 -18876
rect -7872 -18910 -7408 -18876
rect -6854 -18910 -6390 -18876
rect -5836 -18910 -5372 -18876
rect -4818 -18910 -4354 -18876
rect -3800 -18910 -3336 -18876
rect -2782 -18910 -2318 -18876
rect -1764 -18910 -1300 -18876
rect -746 -18910 -282 -18876
rect 2874 -19080 3338 -19046
rect 3892 -19080 4356 -19046
rect 4910 -19080 5374 -19046
rect 5928 -19080 6392 -19046
rect 6946 -19080 7410 -19046
rect 7964 -19080 8428 -19046
rect 8982 -19080 9446 -19046
rect 10000 -19080 10464 -19046
rect 11018 -19080 11482 -19046
rect 12036 -19080 12500 -19046
rect 13054 -19080 13518 -19046
rect 14072 -19080 14536 -19046
rect 15090 -19080 15554 -19046
rect 16108 -19080 16572 -19046
rect 17126 -19080 17590 -19046
rect 18144 -19080 18608 -19046
rect 19162 -19080 19626 -19046
rect 20180 -19080 20644 -19046
rect 21198 -19080 21662 -19046
rect 22216 -19080 22680 -19046
rect -2230 -19584 -2166 -19550
rect -2012 -19584 -1948 -19550
rect -1794 -19584 -1730 -19550
rect -1576 -19584 -1512 -19550
rect -1358 -19584 -1294 -19550
rect -1140 -19584 -1076 -19550
rect -922 -19584 -858 -19550
rect -704 -19584 -640 -19550
rect -486 -19584 -422 -19550
rect -268 -19584 -204 -19550
rect -2324 -19810 -2290 -19634
rect -2106 -19810 -2072 -19634
rect -1888 -19810 -1854 -19634
rect -1670 -19810 -1636 -19634
rect -1452 -19810 -1418 -19634
rect -1234 -19810 -1200 -19634
rect -1016 -19810 -982 -19634
rect -798 -19810 -764 -19634
rect -580 -19810 -546 -19634
rect -362 -19810 -328 -19634
rect -144 -19810 -110 -19634
rect 2580 -19706 2614 -19130
rect 3598 -19706 3632 -19130
rect 4616 -19706 4650 -19130
rect 5634 -19706 5668 -19130
rect 6652 -19706 6686 -19130
rect 7670 -19706 7704 -19130
rect 8688 -19706 8722 -19130
rect 9706 -19706 9740 -19130
rect 10724 -19706 10758 -19130
rect 11742 -19706 11776 -19130
rect 12760 -19706 12794 -19130
rect 13778 -19706 13812 -19130
rect 14796 -19706 14830 -19130
rect 15814 -19706 15848 -19130
rect 16832 -19706 16866 -19130
rect 17850 -19706 17884 -19130
rect 18868 -19706 18902 -19130
rect 19886 -19706 19920 -19130
rect 20904 -19706 20938 -19130
rect 21922 -19706 21956 -19130
rect 22940 -19706 22974 -19130
rect 2874 -19790 3338 -19756
rect 3892 -19790 4356 -19756
rect 4910 -19790 5374 -19756
rect 5928 -19790 6392 -19756
rect 6946 -19790 7410 -19756
rect 7964 -19790 8428 -19756
rect 8982 -19790 9446 -19756
rect 10000 -19790 10464 -19756
rect 11018 -19790 11482 -19756
rect 12036 -19790 12500 -19756
rect 13054 -19790 13518 -19756
rect 14072 -19790 14536 -19756
rect 15090 -19790 15554 -19756
rect 16108 -19790 16572 -19756
rect 17126 -19790 17590 -19756
rect 18144 -19790 18608 -19756
rect 19162 -19790 19626 -19756
rect 20180 -19790 20644 -19756
rect 21198 -19790 21662 -19756
rect 22216 -19790 22680 -19756
rect -2230 -19894 -2166 -19860
rect -2012 -19894 -1948 -19860
rect -1794 -19894 -1730 -19860
rect -1576 -19894 -1512 -19860
rect -1358 -19894 -1294 -19860
rect -1140 -19894 -1076 -19860
rect -922 -19894 -858 -19860
rect -704 -19894 -640 -19860
rect -486 -19894 -422 -19860
rect -268 -19894 -204 -19860
rect 2874 -20314 3338 -20280
rect 3892 -20314 4356 -20280
rect 4910 -20314 5374 -20280
rect 5928 -20314 6392 -20280
rect 6946 -20314 7410 -20280
rect 7964 -20314 8428 -20280
rect 8982 -20314 9446 -20280
rect 10000 -20314 10464 -20280
rect 11018 -20314 11482 -20280
rect 12036 -20314 12500 -20280
rect 13054 -20314 13518 -20280
rect 14072 -20314 14536 -20280
rect 15090 -20314 15554 -20280
rect 16108 -20314 16572 -20280
rect 17126 -20314 17590 -20280
rect 18144 -20314 18608 -20280
rect 19162 -20314 19626 -20280
rect 20180 -20314 20644 -20280
rect 21198 -20314 21662 -20280
rect 22216 -20314 22680 -20280
rect -2230 -20416 -2166 -20382
rect -2012 -20416 -1948 -20382
rect -1794 -20416 -1730 -20382
rect -1576 -20416 -1512 -20382
rect -1358 -20416 -1294 -20382
rect -1140 -20416 -1076 -20382
rect -922 -20416 -858 -20382
rect -704 -20416 -640 -20382
rect -486 -20416 -422 -20382
rect -268 -20416 -204 -20382
rect -2324 -20642 -2290 -20466
rect -2106 -20642 -2072 -20466
rect -1888 -20642 -1854 -20466
rect -1670 -20642 -1636 -20466
rect -1452 -20642 -1418 -20466
rect -1234 -20642 -1200 -20466
rect -1016 -20642 -982 -20466
rect -798 -20642 -764 -20466
rect -580 -20642 -546 -20466
rect -362 -20642 -328 -20466
rect -144 -20642 -110 -20466
rect -2230 -20726 -2166 -20692
rect -2012 -20726 -1948 -20692
rect -1794 -20726 -1730 -20692
rect -1576 -20726 -1512 -20692
rect -1358 -20726 -1294 -20692
rect -1140 -20726 -1076 -20692
rect -922 -20726 -858 -20692
rect -704 -20726 -640 -20692
rect -486 -20726 -422 -20692
rect -268 -20726 -204 -20692
rect 2580 -20940 2614 -20364
rect 3598 -20940 3632 -20364
rect 4616 -20940 4650 -20364
rect 5634 -20940 5668 -20364
rect 6652 -20940 6686 -20364
rect 7670 -20940 7704 -20364
rect 8688 -20940 8722 -20364
rect 9706 -20940 9740 -20364
rect 10724 -20940 10758 -20364
rect 11742 -20940 11776 -20364
rect 12760 -20940 12794 -20364
rect 13778 -20940 13812 -20364
rect 14796 -20940 14830 -20364
rect 15814 -20940 15848 -20364
rect 16832 -20940 16866 -20364
rect 17850 -20940 17884 -20364
rect 18868 -20940 18902 -20364
rect 19886 -20940 19920 -20364
rect 20904 -20940 20938 -20364
rect 21922 -20940 21956 -20364
rect 22940 -20940 22974 -20364
rect 2874 -21024 3338 -20990
rect 3892 -21024 4356 -20990
rect 4910 -21024 5374 -20990
rect 5928 -21024 6392 -20990
rect 6946 -21024 7410 -20990
rect 7964 -21024 8428 -20990
rect 8982 -21024 9446 -20990
rect 10000 -21024 10464 -20990
rect 11018 -21024 11482 -20990
rect 12036 -21024 12500 -20990
rect 13054 -21024 13518 -20990
rect 14072 -21024 14536 -20990
rect 15090 -21024 15554 -20990
rect 16108 -21024 16572 -20990
rect 17126 -21024 17590 -20990
rect 18144 -21024 18608 -20990
rect 19162 -21024 19626 -20990
rect 20180 -21024 20644 -20990
rect 21198 -21024 21662 -20990
rect 22216 -21024 22680 -20990
rect 2874 -21546 3338 -21512
rect 3892 -21546 4356 -21512
rect 4910 -21546 5374 -21512
rect 5928 -21546 6392 -21512
rect 6946 -21546 7410 -21512
rect 7964 -21546 8428 -21512
rect 8982 -21546 9446 -21512
rect 10000 -21546 10464 -21512
rect 11018 -21546 11482 -21512
rect 12036 -21546 12500 -21512
rect 13054 -21546 13518 -21512
rect 14072 -21546 14536 -21512
rect 15090 -21546 15554 -21512
rect 16108 -21546 16572 -21512
rect 17126 -21546 17590 -21512
rect 18144 -21546 18608 -21512
rect 19162 -21546 19626 -21512
rect 20180 -21546 20644 -21512
rect 21198 -21546 21662 -21512
rect 22216 -21546 22680 -21512
rect -9111 -21743 -8647 -21709
rect -8093 -21743 -7629 -21709
rect -7075 -21743 -6611 -21709
rect -6057 -21743 -5593 -21709
rect -5039 -21743 -4575 -21709
rect -4021 -21743 -3557 -21709
rect -2296 -21742 -2192 -21708
rect -1998 -21742 -1894 -21708
rect -1700 -21742 -1596 -21708
rect -1402 -21742 -1298 -21708
rect -1104 -21742 -1000 -21708
rect -806 -21742 -702 -21708
rect -508 -21742 -404 -21708
rect -210 -21742 -106 -21708
rect 88 -21742 192 -21708
rect 386 -21742 490 -21708
rect 684 -21742 788 -21708
rect -9405 -22369 -9371 -21793
rect -8387 -22369 -8353 -21793
rect -7369 -22369 -7335 -21793
rect -6351 -22369 -6317 -21793
rect -5333 -22369 -5299 -21793
rect -4315 -22369 -4281 -21793
rect -3297 -22369 -3263 -21793
rect -2410 -22368 -2376 -21792
rect -2112 -22368 -2078 -21792
rect -1814 -22368 -1780 -21792
rect -1516 -22368 -1482 -21792
rect -1218 -22368 -1184 -21792
rect -920 -22368 -886 -21792
rect -622 -22368 -588 -21792
rect -324 -22368 -290 -21792
rect -26 -22368 8 -21792
rect 272 -22368 306 -21792
rect 570 -22368 604 -21792
rect 868 -22368 902 -21792
rect 2580 -22172 2614 -21596
rect 3598 -22172 3632 -21596
rect 4616 -22172 4650 -21596
rect 5634 -22172 5668 -21596
rect 6652 -22172 6686 -21596
rect 7670 -22172 7704 -21596
rect 8688 -22172 8722 -21596
rect 9706 -22172 9740 -21596
rect 10724 -22172 10758 -21596
rect 11742 -22172 11776 -21596
rect 12760 -22172 12794 -21596
rect 13778 -22172 13812 -21596
rect 14796 -22172 14830 -21596
rect 15814 -22172 15848 -21596
rect 16832 -22172 16866 -21596
rect 17850 -22172 17884 -21596
rect 18868 -22172 18902 -21596
rect 19886 -22172 19920 -21596
rect 20904 -22172 20938 -21596
rect 21922 -22172 21956 -21596
rect 22940 -22172 22974 -21596
rect 2874 -22256 3338 -22222
rect 3892 -22256 4356 -22222
rect 4910 -22256 5374 -22222
rect 5928 -22256 6392 -22222
rect 6946 -22256 7410 -22222
rect 7964 -22256 8428 -22222
rect 8982 -22256 9446 -22222
rect 10000 -22256 10464 -22222
rect 11018 -22256 11482 -22222
rect 12036 -22256 12500 -22222
rect 13054 -22256 13518 -22222
rect 14072 -22256 14536 -22222
rect 15090 -22256 15554 -22222
rect 16108 -22256 16572 -22222
rect 17126 -22256 17590 -22222
rect 18144 -22256 18608 -22222
rect 19162 -22256 19626 -22222
rect 20180 -22256 20644 -22222
rect 21198 -22228 21662 -22222
rect 21198 -22256 21408 -22228
rect 21468 -22256 21662 -22228
rect 22216 -22256 22680 -22222
rect -9111 -22453 -8647 -22419
rect -8093 -22453 -7629 -22419
rect -7075 -22453 -6611 -22419
rect -6057 -22453 -5593 -22419
rect -5039 -22453 -4575 -22419
rect -4021 -22453 -3557 -22419
rect -2296 -22452 -2192 -22418
rect -1998 -22452 -1894 -22418
rect -1700 -22452 -1596 -22418
rect -1402 -22452 -1298 -22418
rect -1104 -22452 -1000 -22418
rect -806 -22452 -702 -22418
rect -508 -22452 -404 -22418
rect -210 -22452 -106 -22418
rect 88 -22452 192 -22418
rect 386 -22452 490 -22418
rect 684 -22452 788 -22418
rect 2874 -22780 3338 -22746
rect 3892 -22780 4356 -22746
rect 4910 -22780 5374 -22746
rect 5928 -22780 6392 -22746
rect 6946 -22780 7410 -22746
rect 7964 -22780 8428 -22746
rect 8982 -22780 9446 -22746
rect 10000 -22780 10464 -22746
rect 11018 -22780 11482 -22746
rect 12036 -22780 12500 -22746
rect 13054 -22780 13518 -22746
rect 14072 -22780 14536 -22746
rect 15090 -22780 15554 -22746
rect 16108 -22780 16572 -22746
rect 17126 -22780 17590 -22746
rect 18144 -22780 18608 -22746
rect 19162 -22780 19626 -22746
rect 20180 -22780 20644 -22746
rect 21198 -22780 21662 -22746
rect 22216 -22780 22680 -22746
rect -9112 -22856 -8648 -22822
rect -8094 -22856 -7630 -22822
rect -7076 -22856 -6612 -22822
rect -6058 -22856 -5594 -22822
rect -5040 -22856 -4576 -22822
rect -4022 -22856 -3558 -22822
rect -2296 -22854 -2192 -22820
rect -1998 -22854 -1894 -22820
rect -1700 -22854 -1596 -22820
rect -1402 -22854 -1298 -22820
rect -1104 -22854 -1000 -22820
rect -806 -22854 -702 -22820
rect -508 -22854 -404 -22820
rect -210 -22854 -106 -22820
rect 88 -22854 192 -22820
rect 386 -22854 490 -22820
rect 684 -22854 788 -22820
rect -9406 -23482 -9372 -22906
rect -8388 -23482 -8354 -22906
rect -7370 -23482 -7336 -22906
rect -6352 -23482 -6318 -22906
rect -5334 -23482 -5300 -22906
rect -4316 -23482 -4282 -22906
rect -3298 -23482 -3264 -22906
rect -2410 -23480 -2376 -22904
rect -2112 -23480 -2078 -22904
rect -1814 -23480 -1780 -22904
rect -1516 -23480 -1482 -22904
rect -1218 -23480 -1184 -22904
rect -920 -23480 -886 -22904
rect -622 -23480 -588 -22904
rect -324 -23480 -290 -22904
rect -26 -23480 8 -22904
rect 272 -23480 306 -22904
rect 570 -23480 604 -22904
rect 868 -23480 902 -22904
rect 2580 -23406 2614 -22830
rect 3598 -23406 3632 -22830
rect 4616 -23406 4650 -22830
rect 5634 -23406 5668 -22830
rect 6652 -23406 6686 -22830
rect 7670 -23406 7704 -22830
rect 8688 -23406 8722 -22830
rect 9706 -23406 9740 -22830
rect 10724 -23406 10758 -22830
rect 11742 -23406 11776 -22830
rect 12760 -23406 12794 -22830
rect 13778 -23406 13812 -22830
rect 14796 -23406 14830 -22830
rect 15814 -23406 15848 -22830
rect 16832 -23406 16866 -22830
rect 17850 -23406 17884 -22830
rect 18868 -23406 18902 -22830
rect 19886 -23406 19920 -22830
rect 20904 -23406 20938 -22830
rect 21922 -23406 21956 -22830
rect 22940 -23406 22974 -22830
rect 2874 -23490 3338 -23456
rect 3892 -23490 4356 -23456
rect 4910 -23490 5374 -23456
rect 5928 -23490 6392 -23456
rect 6946 -23490 7410 -23456
rect 7964 -23490 8428 -23456
rect 8982 -23490 9446 -23456
rect 10000 -23490 10464 -23456
rect 11018 -23490 11482 -23456
rect 12036 -23490 12500 -23456
rect 13054 -23490 13518 -23456
rect 14072 -23490 14536 -23456
rect 15090 -23490 15554 -23456
rect 16108 -23490 16572 -23456
rect 17126 -23490 17590 -23456
rect 18144 -23490 18608 -23456
rect 19162 -23490 19626 -23456
rect 20180 -23490 20644 -23456
rect 21198 -23490 21662 -23456
rect 22216 -23490 22680 -23456
rect -9112 -23566 -8648 -23532
rect -8094 -23566 -7630 -23532
rect -7076 -23566 -6612 -23532
rect -6058 -23566 -5594 -23532
rect -5040 -23566 -4576 -23532
rect -4022 -23566 -3558 -23532
rect -2296 -23564 -2192 -23530
rect -1998 -23564 -1894 -23530
rect -1700 -23564 -1596 -23530
rect -1402 -23564 -1298 -23530
rect -1104 -23564 -1000 -23530
rect -806 -23564 -702 -23530
rect -508 -23564 -404 -23530
rect -210 -23564 -106 -23530
rect 88 -23564 192 -23530
rect 386 -23564 490 -23530
rect 684 -23564 788 -23530
rect -9111 -23967 -8647 -23933
rect -8093 -23967 -7629 -23933
rect -7075 -23967 -6611 -23933
rect -6057 -23967 -5593 -23933
rect -5039 -23967 -4575 -23933
rect -4021 -23967 -3557 -23933
rect -2298 -23966 -2194 -23932
rect -2000 -23966 -1896 -23932
rect -1702 -23966 -1598 -23932
rect -1404 -23966 -1300 -23932
rect -1106 -23966 -1002 -23932
rect -808 -23966 -704 -23932
rect -510 -23966 -406 -23932
rect -212 -23966 -108 -23932
rect 86 -23966 190 -23932
rect 384 -23966 488 -23932
rect 682 -23966 786 -23932
rect -9405 -24593 -9371 -24017
rect -8387 -24593 -8353 -24017
rect -7369 -24593 -7335 -24017
rect -6351 -24593 -6317 -24017
rect -5333 -24593 -5299 -24017
rect -4315 -24593 -4281 -24017
rect -3297 -24593 -3263 -24017
rect -2412 -24592 -2378 -24016
rect -2114 -24592 -2080 -24016
rect -1816 -24592 -1782 -24016
rect -1518 -24592 -1484 -24016
rect -1220 -24592 -1186 -24016
rect -922 -24592 -888 -24016
rect -624 -24592 -590 -24016
rect -326 -24592 -292 -24016
rect -28 -24592 6 -24016
rect 270 -24592 304 -24016
rect 568 -24592 602 -24016
rect 2874 -24014 3338 -23980
rect 3892 -24014 4356 -23980
rect 4910 -24014 5374 -23980
rect 5928 -24014 6392 -23980
rect 6946 -24014 7410 -23980
rect 7964 -24014 8428 -23980
rect 8982 -24014 9446 -23980
rect 10000 -24014 10464 -23980
rect 11018 -24014 11482 -23980
rect 12036 -24014 12500 -23980
rect 13054 -24014 13518 -23980
rect 14072 -24014 14536 -23980
rect 15090 -24014 15554 -23980
rect 16108 -24014 16572 -23980
rect 17126 -24014 17590 -23980
rect 18144 -24014 18608 -23980
rect 19162 -24014 19626 -23980
rect 20180 -24014 20644 -23980
rect 21198 -24014 21662 -23980
rect 22216 -24014 22680 -23980
rect 866 -24592 900 -24016
rect 2580 -24640 2614 -24064
rect -9111 -24677 -8647 -24643
rect -8093 -24677 -7629 -24643
rect -7075 -24677 -6611 -24643
rect -6057 -24677 -5593 -24643
rect -5039 -24677 -4575 -24643
rect -4021 -24677 -3557 -24643
rect -2298 -24676 -2194 -24642
rect -2000 -24676 -1896 -24642
rect -1702 -24676 -1598 -24642
rect -1404 -24676 -1300 -24642
rect -1106 -24676 -1002 -24642
rect -808 -24676 -704 -24642
rect -510 -24676 -406 -24642
rect -212 -24676 -108 -24642
rect 86 -24676 190 -24642
rect 384 -24676 488 -24642
rect 682 -24676 786 -24642
rect 3598 -24640 3632 -24064
rect 4616 -24640 4650 -24064
rect 5634 -24640 5668 -24064
rect 6652 -24640 6686 -24064
rect 7670 -24640 7704 -24064
rect 8688 -24640 8722 -24064
rect 9706 -24640 9740 -24064
rect 10724 -24640 10758 -24064
rect 11742 -24640 11776 -24064
rect 12760 -24640 12794 -24064
rect 13778 -24640 13812 -24064
rect 14796 -24640 14830 -24064
rect 15814 -24640 15848 -24064
rect 16832 -24640 16866 -24064
rect 17850 -24640 17884 -24064
rect 18868 -24640 18902 -24064
rect 19886 -24640 19920 -24064
rect 20904 -24640 20938 -24064
rect 21922 -24640 21956 -24064
rect 22940 -24640 22974 -24064
rect 2874 -24724 3338 -24690
rect 3892 -24724 4356 -24690
rect 4910 -24724 5374 -24690
rect 5928 -24724 6392 -24690
rect 6946 -24724 7410 -24690
rect 7964 -24724 8428 -24690
rect 8982 -24724 9446 -24690
rect 10000 -24724 10464 -24690
rect 11018 -24724 11482 -24690
rect 12036 -24724 12500 -24690
rect 13054 -24724 13518 -24690
rect 14072 -24724 14536 -24690
rect 15090 -24724 15554 -24690
rect 16108 -24724 16572 -24690
rect 17126 -24724 17590 -24690
rect 18144 -24724 18608 -24690
rect 19162 -24724 19626 -24690
rect 20180 -24724 20644 -24690
rect 21198 -24724 21662 -24690
rect 22216 -24724 22680 -24690
rect -9112 -25080 -8648 -25046
rect -8094 -25080 -7630 -25046
rect -7076 -25080 -6612 -25046
rect -6058 -25080 -5594 -25046
rect -5040 -25080 -4576 -25046
rect -4022 -25080 -3558 -25046
rect -2298 -25076 -2194 -25042
rect -2000 -25076 -1896 -25042
rect -1702 -25076 -1598 -25042
rect -1404 -25076 -1300 -25042
rect -1106 -25076 -1002 -25042
rect -808 -25076 -704 -25042
rect -510 -25076 -406 -25042
rect -212 -25076 -108 -25042
rect 86 -25076 190 -25042
rect 384 -25076 488 -25042
rect 682 -25076 786 -25042
rect -9406 -25706 -9372 -25130
rect -8388 -25706 -8354 -25130
rect -7370 -25706 -7336 -25130
rect -6352 -25706 -6318 -25130
rect -5334 -25706 -5300 -25130
rect -4316 -25706 -4282 -25130
rect -3298 -25706 -3264 -25130
rect -2412 -25702 -2378 -25126
rect -2114 -25702 -2080 -25126
rect -1816 -25702 -1782 -25126
rect -1518 -25702 -1484 -25126
rect -1220 -25702 -1186 -25126
rect -922 -25702 -888 -25126
rect -624 -25702 -590 -25126
rect -326 -25702 -292 -25126
rect -28 -25702 6 -25126
rect 270 -25702 304 -25126
rect 568 -25702 602 -25126
rect 866 -25702 900 -25126
rect 2874 -25246 3338 -25212
rect 3892 -25246 4356 -25212
rect 4910 -25246 5374 -25212
rect 5928 -25246 6392 -25212
rect 6946 -25246 7410 -25212
rect 7964 -25246 8428 -25212
rect 8982 -25246 9446 -25212
rect 10000 -25246 10464 -25212
rect 11018 -25246 11482 -25212
rect 12036 -25246 12500 -25212
rect 13054 -25246 13518 -25212
rect 14072 -25246 14536 -25212
rect 15090 -25246 15554 -25212
rect 16108 -25246 16572 -25212
rect 17126 -25246 17590 -25212
rect 18144 -25246 18608 -25212
rect 19162 -25246 19626 -25212
rect 20180 -25246 20644 -25212
rect 21198 -25246 21662 -25212
rect 22216 -25246 22680 -25212
rect -9112 -25790 -8648 -25756
rect -8094 -25790 -7630 -25756
rect -7076 -25790 -6612 -25756
rect -6058 -25790 -5594 -25756
rect -5040 -25790 -4576 -25756
rect -4022 -25790 -3558 -25756
rect -2298 -25786 -2194 -25752
rect -2000 -25786 -1896 -25752
rect -1702 -25786 -1598 -25752
rect -1404 -25786 -1300 -25752
rect -1106 -25786 -1002 -25752
rect -808 -25786 -704 -25752
rect -510 -25786 -406 -25752
rect -212 -25786 -108 -25752
rect 86 -25786 190 -25752
rect 384 -25786 488 -25752
rect 682 -25786 786 -25752
rect 2580 -25872 2614 -25296
rect 3598 -25872 3632 -25296
rect 4616 -25872 4650 -25296
rect 5634 -25872 5668 -25296
rect 6652 -25872 6686 -25296
rect 7670 -25872 7704 -25296
rect 8688 -25872 8722 -25296
rect 9706 -25872 9740 -25296
rect 10724 -25872 10758 -25296
rect 11742 -25872 11776 -25296
rect 12760 -25872 12794 -25296
rect 13778 -25872 13812 -25296
rect 14796 -25872 14830 -25296
rect 15814 -25872 15848 -25296
rect 16832 -25872 16866 -25296
rect 17850 -25872 17884 -25296
rect 18868 -25872 18902 -25296
rect 19886 -25872 19920 -25296
rect 20904 -25872 20938 -25296
rect 21922 -25872 21956 -25296
rect 22940 -25872 22974 -25296
rect 2874 -25956 3338 -25922
rect 3892 -25956 4356 -25922
rect 4910 -25956 5374 -25922
rect 5928 -25956 6392 -25922
rect 6946 -25956 7410 -25922
rect 7964 -25956 8428 -25922
rect 8982 -25956 9446 -25922
rect 10000 -25956 10464 -25922
rect 11018 -25956 11482 -25922
rect 12036 -25956 12500 -25922
rect 13054 -25956 13518 -25922
rect 14072 -25956 14536 -25922
rect 15090 -25956 15554 -25922
rect 16108 -25956 16572 -25922
rect 17126 -25956 17590 -25922
rect 18144 -25956 18608 -25922
rect 19162 -25956 19626 -25922
rect 20180 -25956 20644 -25922
rect 21198 -25956 21662 -25922
rect 22216 -25956 22680 -25922
rect 24822 -26330 24922 -12070
rect -12222 -27222 -12160 -27122
rect -12160 -27222 24760 -27122
rect 24760 -27222 24822 -27122
<< metal1 >>
rect 372 1722 24828 1728
rect 372 1622 478 1722
rect 24722 1622 24828 1722
rect 372 1616 24828 1622
rect 372 1102 484 1616
rect 1084 1316 1094 1616
rect 24106 1316 24116 1616
rect 372 -8262 378 1102
rect 478 -8262 484 1102
rect 3998 1234 20878 1266
rect 3998 1020 4061 1234
rect 20846 1020 20878 1234
rect 3998 1000 20878 1020
rect 24716 1102 24828 1616
rect 3998 998 8352 1000
rect 3614 -4562 4002 -4502
rect 3614 -4702 3674 -4562
rect 3716 -4603 3776 -4562
rect 3708 -4609 3796 -4603
rect 3708 -4643 3720 -4609
rect 3784 -4643 3796 -4609
rect 3708 -4649 3796 -4643
rect 3614 -4730 3626 -4702
rect 3620 -5078 3626 -4730
rect 3660 -4730 3674 -4702
rect 3832 -4702 3892 -4562
rect 3942 -4603 4002 -4562
rect 3926 -4609 4014 -4603
rect 3926 -4643 3938 -4609
rect 4002 -4643 4014 -4609
rect 3926 -4649 4014 -4643
rect 3660 -5078 3666 -4730
rect 3832 -4734 3844 -4702
rect 3838 -5048 3844 -4734
rect 3620 -5090 3666 -5078
rect 3832 -5078 3844 -5048
rect 3878 -4734 3892 -4702
rect 4048 -4702 4108 998
rect 4150 -4562 4156 -4502
rect 4216 -4562 4222 -4502
rect 4262 -4562 4268 -4502
rect 4328 -4562 4334 -4502
rect 4372 -4562 4378 -4502
rect 4438 -4562 4444 -4502
rect 4156 -4603 4216 -4562
rect 4144 -4609 4232 -4603
rect 4144 -4643 4156 -4609
rect 4220 -4643 4232 -4609
rect 4144 -4649 4232 -4643
rect 3878 -5048 3884 -4734
rect 3878 -5078 3892 -5048
rect 3708 -5137 3796 -5131
rect 3708 -5171 3720 -5137
rect 3784 -5171 3796 -5137
rect 3708 -5177 3796 -5171
rect 3832 -5214 3892 -5078
rect 4048 -5078 4062 -4702
rect 4096 -5078 4108 -4702
rect 4268 -4702 4328 -4562
rect 4378 -4603 4438 -4562
rect 4362 -4609 4376 -4603
rect 4378 -4609 4450 -4603
rect 4362 -4643 4374 -4609
rect 4438 -4643 4450 -4609
rect 4362 -4649 4450 -4643
rect 4268 -4728 4280 -4702
rect 3926 -5137 4014 -5131
rect 3926 -5171 3938 -5137
rect 4002 -5171 4014 -5137
rect 3926 -5177 4014 -5171
rect 3942 -5214 4002 -5177
rect 3486 -5274 3492 -5214
rect 3552 -5274 3558 -5214
rect 3826 -5274 3832 -5214
rect 3892 -5274 3898 -5214
rect 3936 -5274 3942 -5214
rect 4002 -5274 4008 -5214
rect 2104 -6220 2110 -6160
rect 2170 -6220 2176 -6160
rect 372 -8776 484 -8262
rect 2110 -8392 2170 -6220
rect 3492 -6998 3552 -5274
rect 4048 -5320 4108 -5078
rect 4274 -5078 4280 -4728
rect 4314 -4728 4328 -4702
rect 4484 -4702 4544 998
rect 4580 -4609 4668 -4603
rect 4580 -4643 4592 -4609
rect 4656 -4643 4668 -4609
rect 4580 -4649 4668 -4643
rect 4798 -4609 4886 -4603
rect 4798 -4643 4810 -4609
rect 4874 -4643 4886 -4609
rect 4798 -4649 4886 -4643
rect 4314 -5078 4320 -4728
rect 4274 -5090 4320 -5078
rect 4484 -5078 4498 -4702
rect 4532 -5078 4544 -4702
rect 4710 -4702 4756 -4690
rect 4710 -5046 4716 -4702
rect 4144 -5137 4232 -5131
rect 4144 -5171 4156 -5137
rect 4220 -5171 4232 -5137
rect 4144 -5177 4232 -5171
rect 4362 -5137 4450 -5131
rect 4362 -5171 4374 -5137
rect 4438 -5171 4450 -5137
rect 4362 -5177 4450 -5171
rect 4484 -5320 4544 -5078
rect 4704 -5078 4716 -5046
rect 4750 -5046 4756 -4702
rect 4922 -4702 4982 998
rect 5022 -4562 5028 -4502
rect 5088 -4562 5094 -4502
rect 5132 -4562 5138 -4502
rect 5198 -4562 5204 -4502
rect 5240 -4562 5246 -4502
rect 5306 -4562 5312 -4502
rect 5028 -4603 5088 -4562
rect 5016 -4609 5088 -4603
rect 5090 -4609 5104 -4603
rect 5016 -4643 5028 -4609
rect 5092 -4643 5104 -4609
rect 5016 -4649 5104 -4643
rect 4750 -5078 4764 -5046
rect 4580 -5137 4668 -5131
rect 4580 -5171 4592 -5137
rect 4656 -5171 4668 -5137
rect 4580 -5177 4668 -5171
rect 4592 -5214 4652 -5177
rect 4704 -5214 4764 -5078
rect 4922 -5078 4934 -4702
rect 4968 -5078 4982 -4702
rect 5138 -4702 5198 -4562
rect 5246 -4603 5306 -4562
rect 5234 -4609 5306 -4603
rect 5308 -4609 5322 -4603
rect 5234 -4643 5246 -4609
rect 5310 -4643 5322 -4609
rect 5234 -4649 5322 -4643
rect 5138 -4730 5152 -4702
rect 4798 -5137 4886 -5131
rect 4798 -5171 4810 -5137
rect 4874 -5171 4886 -5137
rect 4798 -5177 4886 -5171
rect 4812 -5214 4872 -5177
rect 4586 -5274 4592 -5214
rect 4652 -5274 4658 -5214
rect 4698 -5274 4704 -5214
rect 4764 -5274 4770 -5214
rect 4806 -5274 4812 -5214
rect 4872 -5274 4878 -5214
rect 4922 -5320 4982 -5078
rect 5146 -5078 5152 -4730
rect 5186 -4730 5198 -4702
rect 5356 -4702 5416 998
rect 7980 824 7986 884
rect 8046 824 8052 884
rect 6474 608 7552 668
rect 6474 388 6534 608
rect 6978 492 7038 608
rect 7492 402 7552 608
rect 7986 484 8046 824
rect 8512 638 8572 1000
rect 9062 824 9068 884
rect 9128 824 9134 884
rect 10020 824 10026 884
rect 10086 824 10092 884
rect 8506 578 8512 638
rect 8572 578 8578 638
rect 8512 404 8572 578
rect 9068 482 9128 824
rect 10026 478 10086 824
rect 10548 638 10608 1000
rect 11056 824 11062 884
rect 11122 824 11128 884
rect 12062 824 12068 884
rect 12128 824 12134 884
rect 10542 578 10548 638
rect 10608 578 10614 638
rect 10548 404 10608 578
rect 11062 478 11122 824
rect 11560 690 11566 750
rect 11626 690 11632 750
rect 11566 400 11626 690
rect 12068 488 12128 824
rect 12586 640 12646 1000
rect 13084 824 13090 884
rect 13150 824 13156 884
rect 14102 824 14108 884
rect 14168 824 14174 884
rect 12580 580 12586 640
rect 12646 580 12652 640
rect 12586 388 12646 580
rect 13090 488 13150 824
rect 14108 482 14168 824
rect 14618 640 14678 1000
rect 15126 824 15132 884
rect 15192 824 15198 884
rect 16138 824 16144 884
rect 16204 824 16210 884
rect 14610 580 14616 640
rect 14676 580 14682 640
rect 14618 388 14678 580
rect 15132 488 15192 824
rect 16144 488 16204 824
rect 16658 642 16718 1000
rect 17156 824 17162 884
rect 17222 824 17228 884
rect 18168 824 18174 884
rect 18234 824 18240 884
rect 16652 582 16658 642
rect 16718 582 16724 642
rect 16658 390 16718 582
rect 17162 488 17222 824
rect 17664 690 17670 750
rect 17730 690 17736 750
rect 17670 386 17730 690
rect 18174 482 18234 824
rect 18690 642 18750 1000
rect 19196 824 19202 884
rect 19262 824 19268 884
rect 20208 824 20214 884
rect 20274 824 20280 884
rect 18684 582 18690 642
rect 18750 582 18756 642
rect 18690 400 18750 582
rect 19202 488 19262 824
rect 20214 488 20274 824
rect 20726 642 20786 1000
rect 21226 824 21232 884
rect 21292 824 21298 884
rect 20720 582 20726 642
rect 20786 582 20792 642
rect 20726 396 20786 582
rect 21232 482 21292 824
rect 21746 590 22826 650
rect 21746 398 21806 590
rect 22248 488 22308 590
rect 22766 382 22826 590
rect 7494 -294 7554 -112
rect 6324 -354 6330 -294
rect 6390 -354 6396 -294
rect 7488 -354 7494 -294
rect 7554 -354 7560 -294
rect 6194 -558 6200 -498
rect 6260 -558 6266 -498
rect 6200 -3426 6260 -558
rect 6330 -2968 6390 -354
rect 7488 -558 7494 -498
rect 7554 -558 7560 -498
rect 7494 -746 7554 -558
rect 7998 -658 8058 -200
rect 8514 -748 8574 -108
rect 9020 -652 9080 -194
rect 9530 -398 9590 -120
rect 9524 -458 9530 -398
rect 9590 -458 9596 -398
rect 10050 -652 10110 -194
rect 10538 -738 10602 -90
rect 11050 -646 11110 -188
rect 11560 -458 11566 -398
rect 11626 -458 11632 -398
rect 11566 -746 11626 -458
rect 12068 -652 12128 -194
rect 12574 -742 12638 -94
rect 13092 -656 13152 -198
rect 13604 -294 13664 -108
rect 13598 -354 13604 -294
rect 13664 -354 13670 -294
rect 13594 -558 13600 -498
rect 13660 -558 13666 -498
rect 13600 -734 13660 -558
rect 14110 -650 14170 -192
rect 14616 -740 14680 -92
rect 15126 -658 15186 -195
rect 15638 -294 15698 -110
rect 15632 -354 15638 -294
rect 15698 -354 15704 -294
rect 15630 -558 15636 -498
rect 15696 -558 15702 -498
rect 15636 -740 15696 -558
rect 16138 -658 16198 -195
rect 16654 -756 16718 -108
rect 17144 -658 17204 -195
rect 17672 -300 17732 -116
rect 17672 -360 17874 -300
rect 17666 -458 17672 -398
rect 17732 -458 17738 -398
rect 17672 -732 17732 -458
rect 17814 -502 17874 -360
rect 17808 -562 17814 -502
rect 17874 -562 17880 -502
rect 18162 -658 18222 -195
rect 18690 -752 18750 -100
rect 19180 -658 19240 -195
rect 19706 -398 19766 -116
rect 19700 -458 19706 -398
rect 19766 -458 19772 -398
rect 19702 -562 19708 -502
rect 19768 -562 19774 -502
rect 19708 -736 19768 -562
rect 20180 -658 20240 -195
rect 20730 -744 20790 -110
rect 21210 -652 21270 -189
rect 21746 -294 21806 -108
rect 21740 -354 21746 -294
rect 21806 -354 21812 -294
rect 22878 -354 22884 -294
rect 22944 -354 22950 -294
rect 21750 -570 22820 -510
rect 21750 -736 21810 -570
rect 22256 -644 22316 -570
rect 22760 -742 22820 -570
rect 14618 -1238 14678 -1236
rect 6476 -1434 6536 -1248
rect 6988 -1434 7048 -1346
rect 7494 -1434 7554 -1254
rect 10546 -1258 10606 -1256
rect 6476 -1494 7554 -1434
rect 7488 -1642 7548 -1636
rect 6478 -1702 7548 -1642
rect 6478 -1876 6538 -1702
rect 6988 -1778 7048 -1702
rect 7488 -1876 7548 -1702
rect 7980 -1788 8040 -1330
rect 8510 -1432 8570 -1258
rect 8504 -1492 8510 -1432
rect 8570 -1492 8576 -1432
rect 8510 -1896 8570 -1492
rect 9026 -1788 9086 -1330
rect 9528 -1528 9588 -1264
rect 10546 -1432 10610 -1258
rect 10540 -1492 10546 -1432
rect 10606 -1492 10612 -1432
rect 9522 -1588 9528 -1528
rect 9588 -1588 9594 -1528
rect 10226 -1594 10232 -1530
rect 10296 -1594 10302 -1530
rect 10232 -1624 10296 -1594
rect 9530 -1688 10296 -1624
rect 9530 -1890 9594 -1688
rect 10546 -1892 10610 -1492
rect 11074 -1782 11134 -1324
rect 11564 -1530 11628 -1248
rect 12580 -1250 12640 -1248
rect 11398 -1594 11404 -1530
rect 11468 -1594 11628 -1530
rect 11560 -1698 11566 -1638
rect 11626 -1698 11632 -1638
rect 11566 -1880 11626 -1698
rect 12092 -1792 12152 -1334
rect 12580 -1432 12644 -1250
rect 12574 -1492 12580 -1432
rect 12640 -1492 12646 -1432
rect 12580 -1904 12644 -1492
rect 13092 -1788 13152 -1330
rect 14120 -1798 14180 -1340
rect 14618 -1434 14682 -1238
rect 16654 -1242 16714 -1240
rect 14612 -1494 14618 -1434
rect 14678 -1494 14684 -1434
rect 14618 -1884 14682 -1494
rect 15138 -1788 15198 -1325
rect 15638 -1532 15698 -1254
rect 15632 -1592 15638 -1532
rect 15698 -1592 15704 -1532
rect 16138 -1792 16198 -1329
rect 16654 -1434 16718 -1242
rect 16648 -1494 16654 -1434
rect 16714 -1494 16720 -1434
rect 16654 -1896 16718 -1494
rect 17144 -1792 17204 -1329
rect 17666 -1698 17672 -1638
rect 17732 -1698 17738 -1638
rect 17672 -1880 17732 -1698
rect 18186 -1792 18246 -1329
rect 18690 -1434 18750 -1248
rect 18684 -1494 18690 -1434
rect 18750 -1494 18756 -1434
rect 18690 -1898 18750 -1494
rect 19186 -1788 19246 -1325
rect 19708 -1638 19768 -1248
rect 20724 -1254 20784 -1252
rect 19702 -1698 19708 -1638
rect 19768 -1698 19774 -1638
rect 20212 -1792 20272 -1329
rect 20724 -1436 20788 -1254
rect 20718 -1496 20724 -1436
rect 20784 -1496 20790 -1436
rect 20724 -1890 20788 -1496
rect 21210 -1794 21270 -1331
rect 21746 -1532 21806 -1254
rect 21740 -1592 21746 -1532
rect 21806 -1592 21812 -1532
rect 21748 -1646 21808 -1644
rect 21748 -1706 22820 -1646
rect 21748 -1870 21808 -1706
rect 22252 -1782 22312 -1706
rect 22760 -1894 22820 -1706
rect 7488 -2818 7552 -2378
rect 8510 -2570 8570 -2384
rect 10546 -2396 10606 -2394
rect 8504 -2630 8510 -2570
rect 8570 -2630 8576 -2570
rect 9526 -2680 9590 -2396
rect 9520 -2744 9526 -2680
rect 9590 -2744 9596 -2680
rect 7482 -2882 7488 -2818
rect 7552 -2882 7558 -2818
rect 7312 -2968 7372 -2962
rect 6324 -3028 6330 -2968
rect 6390 -3028 6396 -2968
rect 6916 -3304 6976 -3298
rect 6200 -3486 6862 -3426
rect 5576 -4570 5856 -4510
rect 6042 -4562 6048 -4502
rect 6108 -4562 6114 -4502
rect 5452 -4609 5540 -4603
rect 5452 -4643 5464 -4609
rect 5528 -4643 5540 -4609
rect 5452 -4649 5540 -4643
rect 5186 -5078 5192 -4730
rect 5146 -5090 5192 -5078
rect 5356 -5078 5370 -4702
rect 5404 -5078 5416 -4702
rect 5576 -4702 5636 -4570
rect 5684 -4603 5744 -4570
rect 5670 -4609 5758 -4603
rect 5670 -4643 5682 -4609
rect 5746 -4643 5758 -4609
rect 5670 -4649 5758 -4643
rect 5576 -4726 5588 -4702
rect 5582 -5032 5588 -4726
rect 5016 -5137 5104 -5131
rect 5016 -5171 5028 -5137
rect 5092 -5171 5104 -5137
rect 5016 -5177 5104 -5171
rect 5234 -5137 5322 -5131
rect 5234 -5171 5246 -5137
rect 5310 -5171 5322 -5137
rect 5234 -5177 5322 -5171
rect 5356 -5320 5416 -5078
rect 5574 -5078 5588 -5032
rect 5622 -4726 5636 -4702
rect 5796 -4702 5856 -4570
rect 5622 -5032 5628 -4726
rect 5796 -4734 5806 -4702
rect 5622 -5078 5634 -5032
rect 5452 -5137 5540 -5131
rect 5452 -5171 5464 -5137
rect 5528 -5171 5540 -5137
rect 5452 -5177 5540 -5171
rect 5464 -5214 5524 -5177
rect 5574 -5214 5634 -5078
rect 5800 -5078 5806 -4734
rect 5840 -4734 5856 -4702
rect 5840 -5078 5846 -4734
rect 5800 -5090 5846 -5078
rect 5670 -5137 5758 -5131
rect 5670 -5171 5682 -5137
rect 5746 -5171 5758 -5137
rect 5670 -5177 5758 -5171
rect 5458 -5274 5464 -5214
rect 5524 -5274 5530 -5214
rect 5568 -5274 5574 -5214
rect 5634 -5274 5640 -5214
rect 4042 -5380 4048 -5320
rect 4108 -5380 4114 -5320
rect 4478 -5380 4484 -5320
rect 4544 -5380 4550 -5320
rect 4916 -5380 4922 -5320
rect 4982 -5380 4988 -5320
rect 5350 -5380 5356 -5320
rect 5416 -5380 5422 -5320
rect 3616 -5498 3892 -5438
rect 3616 -5640 3676 -5498
rect 3720 -5541 3780 -5498
rect 3708 -5547 3796 -5541
rect 3708 -5581 3720 -5547
rect 3784 -5581 3796 -5547
rect 3708 -5587 3796 -5581
rect 3616 -5674 3626 -5640
rect 3620 -6016 3626 -5674
rect 3660 -5674 3676 -5640
rect 3832 -5640 3892 -5498
rect 3926 -5547 4014 -5541
rect 3926 -5581 3938 -5547
rect 4002 -5581 4014 -5547
rect 3926 -5587 4014 -5581
rect 3832 -5670 3844 -5640
rect 3660 -6016 3666 -5674
rect 3838 -5982 3844 -5670
rect 3620 -6028 3666 -6016
rect 3832 -6016 3844 -5982
rect 3878 -5670 3892 -5640
rect 4048 -5640 4108 -5380
rect 4262 -5496 4268 -5436
rect 4328 -5496 4334 -5436
rect 4144 -5547 4232 -5541
rect 4144 -5581 4156 -5547
rect 4220 -5581 4232 -5547
rect 4144 -5587 4232 -5581
rect 4048 -5668 4062 -5640
rect 3878 -5982 3884 -5670
rect 4056 -5974 4062 -5668
rect 3878 -6016 3892 -5982
rect 3708 -6075 3796 -6069
rect 3708 -6109 3720 -6075
rect 3784 -6109 3796 -6075
rect 3708 -6115 3796 -6109
rect 3832 -6160 3892 -6016
rect 4048 -6016 4062 -5974
rect 4096 -5668 4108 -5640
rect 4268 -5640 4328 -5496
rect 4362 -5547 4450 -5541
rect 4362 -5581 4374 -5547
rect 4438 -5581 4450 -5547
rect 4362 -5587 4450 -5581
rect 4268 -5666 4280 -5640
rect 4096 -5974 4102 -5668
rect 4096 -6016 4108 -5974
rect 3926 -6075 4014 -6069
rect 3926 -6109 3938 -6075
rect 4002 -6109 4014 -6075
rect 3926 -6115 4014 -6109
rect 3826 -6220 3832 -6160
rect 3892 -6220 3898 -6160
rect 3942 -6358 4002 -6115
rect 4048 -6264 4108 -6016
rect 4274 -6016 4280 -5666
rect 4314 -5666 4328 -5640
rect 4484 -5640 4544 -5380
rect 4580 -5547 4668 -5541
rect 4580 -5581 4592 -5547
rect 4656 -5581 4668 -5547
rect 4580 -5587 4668 -5581
rect 4798 -5547 4886 -5541
rect 4798 -5581 4810 -5547
rect 4874 -5581 4886 -5547
rect 4798 -5587 4886 -5581
rect 4314 -6016 4320 -5666
rect 4484 -5670 4498 -5640
rect 4492 -5984 4498 -5670
rect 4274 -6028 4320 -6016
rect 4484 -6016 4498 -5984
rect 4532 -5670 4544 -5640
rect 4710 -5640 4756 -5628
rect 4532 -5984 4538 -5670
rect 4710 -5980 4716 -5640
rect 4532 -6016 4544 -5984
rect 4144 -6075 4232 -6069
rect 4144 -6109 4156 -6075
rect 4220 -6109 4232 -6075
rect 4144 -6115 4232 -6109
rect 4362 -6075 4450 -6069
rect 4362 -6109 4374 -6075
rect 4438 -6109 4450 -6075
rect 4362 -6115 4450 -6109
rect 4042 -6324 4048 -6264
rect 4108 -6324 4114 -6264
rect 3614 -6362 4002 -6358
rect 3614 -6418 3942 -6362
rect 3614 -6578 3674 -6418
rect 3720 -6479 3780 -6418
rect 3708 -6485 3796 -6479
rect 3708 -6519 3720 -6485
rect 3784 -6519 3796 -6485
rect 3708 -6525 3796 -6519
rect 3614 -6604 3626 -6578
rect 3620 -6954 3626 -6604
rect 3660 -6604 3674 -6578
rect 3834 -6578 3894 -6418
rect 3936 -6422 3942 -6418
rect 4002 -6422 4008 -6362
rect 3942 -6479 4002 -6422
rect 3926 -6485 4014 -6479
rect 3926 -6519 3938 -6485
rect 4002 -6519 4014 -6485
rect 3926 -6525 4014 -6519
rect 3660 -6954 3666 -6604
rect 3834 -6616 3844 -6578
rect 3838 -6928 3844 -6616
rect 3620 -6966 3666 -6954
rect 3832 -6954 3844 -6928
rect 3878 -6616 3894 -6578
rect 4048 -6578 4108 -6324
rect 4156 -6362 4216 -6115
rect 4260 -6220 4266 -6160
rect 4326 -6220 4332 -6160
rect 4150 -6422 4156 -6362
rect 4216 -6422 4222 -6362
rect 4156 -6479 4216 -6422
rect 4144 -6485 4232 -6479
rect 4144 -6519 4156 -6485
rect 4220 -6519 4232 -6485
rect 4144 -6525 4232 -6519
rect 4048 -6612 4062 -6578
rect 3878 -6928 3884 -6616
rect 3878 -6954 3892 -6928
rect 4056 -6930 4062 -6612
rect 3708 -7013 3796 -7007
rect 3708 -7047 3720 -7013
rect 3784 -7047 3796 -7013
rect 3708 -7053 3796 -7047
rect 3492 -7314 3552 -7058
rect 3832 -7098 3892 -6954
rect 4048 -6954 4062 -6930
rect 4096 -6612 4108 -6578
rect 4266 -6578 4326 -6220
rect 4376 -6362 4436 -6115
rect 4484 -6264 4544 -6016
rect 4702 -6016 4716 -5980
rect 4750 -5980 4756 -5640
rect 4922 -5640 4982 -5380
rect 5132 -5496 5138 -5436
rect 5198 -5496 5204 -5436
rect 5016 -5547 5104 -5541
rect 5016 -5581 5028 -5547
rect 5092 -5581 5104 -5547
rect 5016 -5587 5104 -5581
rect 4922 -5674 4934 -5640
rect 4750 -6016 4762 -5980
rect 4928 -5988 4934 -5674
rect 4580 -6075 4668 -6069
rect 4580 -6109 4592 -6075
rect 4656 -6109 4668 -6075
rect 4580 -6115 4668 -6109
rect 4478 -6324 4484 -6264
rect 4544 -6324 4550 -6264
rect 4370 -6422 4376 -6362
rect 4436 -6422 4442 -6362
rect 4376 -6479 4436 -6422
rect 4362 -6485 4450 -6479
rect 4362 -6519 4374 -6485
rect 4438 -6519 4450 -6485
rect 4362 -6525 4450 -6519
rect 4266 -6612 4280 -6578
rect 4096 -6930 4102 -6612
rect 4096 -6954 4108 -6930
rect 3926 -7013 4014 -7007
rect 3926 -7047 3938 -7013
rect 4002 -7047 4014 -7013
rect 3926 -7053 4014 -7047
rect 3826 -7158 3832 -7098
rect 3892 -7158 3898 -7098
rect 4048 -7196 4108 -6954
rect 4274 -6954 4280 -6612
rect 4314 -6612 4326 -6578
rect 4484 -6578 4544 -6324
rect 4594 -6362 4654 -6115
rect 4702 -6160 4762 -6016
rect 4922 -6016 4934 -5988
rect 4968 -5674 4982 -5640
rect 5138 -5640 5198 -5496
rect 5234 -5547 5322 -5541
rect 5234 -5581 5246 -5547
rect 5310 -5581 5322 -5547
rect 5234 -5587 5322 -5581
rect 5138 -5672 5152 -5640
rect 4968 -5988 4974 -5674
rect 4968 -6016 4982 -5988
rect 4798 -6075 4886 -6069
rect 4798 -6109 4810 -6075
rect 4874 -6109 4886 -6075
rect 4798 -6115 4886 -6109
rect 4696 -6220 4702 -6160
rect 4762 -6220 4768 -6160
rect 4810 -6362 4870 -6115
rect 4922 -6264 4982 -6016
rect 5146 -6016 5152 -5672
rect 5186 -5672 5198 -5640
rect 5356 -5640 5416 -5380
rect 5576 -5480 5856 -5420
rect 5452 -5547 5540 -5541
rect 5452 -5581 5464 -5547
rect 5528 -5581 5540 -5547
rect 5452 -5587 5540 -5581
rect 5356 -5662 5370 -5640
rect 5186 -6016 5192 -5672
rect 5364 -5986 5370 -5662
rect 5146 -6028 5192 -6016
rect 5356 -6016 5370 -5986
rect 5404 -5662 5416 -5640
rect 5576 -5640 5636 -5480
rect 5686 -5541 5746 -5480
rect 5670 -5547 5758 -5541
rect 5670 -5581 5682 -5547
rect 5746 -5581 5758 -5547
rect 5670 -5587 5758 -5581
rect 5404 -5986 5410 -5662
rect 5576 -5664 5588 -5640
rect 5582 -5980 5588 -5664
rect 5404 -6016 5416 -5986
rect 5016 -6075 5104 -6069
rect 5016 -6109 5028 -6075
rect 5092 -6109 5104 -6075
rect 5016 -6115 5104 -6109
rect 5234 -6075 5322 -6069
rect 5234 -6109 5246 -6075
rect 5310 -6109 5322 -6075
rect 5234 -6115 5322 -6109
rect 4916 -6324 4922 -6264
rect 4982 -6324 4988 -6264
rect 4588 -6422 4594 -6362
rect 4654 -6422 4660 -6362
rect 4698 -6422 4704 -6362
rect 4764 -6422 4770 -6362
rect 4804 -6422 4810 -6362
rect 4870 -6422 4876 -6362
rect 4594 -6479 4654 -6422
rect 4580 -6485 4668 -6479
rect 4580 -6519 4592 -6485
rect 4656 -6519 4668 -6485
rect 4580 -6525 4668 -6519
rect 4314 -6954 4320 -6612
rect 4484 -6614 4498 -6578
rect 4492 -6916 4498 -6614
rect 4274 -6966 4320 -6954
rect 4484 -6954 4498 -6916
rect 4532 -6614 4544 -6578
rect 4704 -6578 4764 -6422
rect 4810 -6479 4870 -6422
rect 4798 -6485 4886 -6479
rect 4798 -6519 4810 -6485
rect 4874 -6519 4886 -6485
rect 4798 -6525 4886 -6519
rect 4704 -6606 4716 -6578
rect 4532 -6916 4538 -6614
rect 4532 -6954 4544 -6916
rect 4710 -6924 4716 -6606
rect 4144 -7013 4232 -7007
rect 4144 -7047 4156 -7013
rect 4220 -7047 4232 -7013
rect 4144 -7053 4232 -7047
rect 4362 -7013 4450 -7007
rect 4362 -7047 4374 -7013
rect 4438 -7047 4450 -7013
rect 4362 -7053 4450 -7047
rect 4484 -7196 4544 -6954
rect 4702 -6954 4716 -6924
rect 4750 -6606 4764 -6578
rect 4922 -6578 4982 -6324
rect 5028 -6362 5088 -6115
rect 5132 -6220 5138 -6160
rect 5198 -6220 5204 -6160
rect 5022 -6422 5028 -6362
rect 5088 -6422 5094 -6362
rect 5028 -6479 5088 -6422
rect 5016 -6485 5104 -6479
rect 5016 -6519 5028 -6485
rect 5092 -6519 5104 -6485
rect 5016 -6525 5104 -6519
rect 4750 -6924 4756 -6606
rect 4922 -6618 4934 -6578
rect 4928 -6920 4934 -6618
rect 4750 -6954 4762 -6924
rect 4580 -7013 4668 -7007
rect 4580 -7047 4592 -7013
rect 4656 -7047 4668 -7013
rect 4580 -7053 4668 -7047
rect 4702 -7098 4762 -6954
rect 4922 -6954 4934 -6920
rect 4968 -6618 4982 -6578
rect 5138 -6578 5198 -6220
rect 5246 -6362 5306 -6115
rect 5356 -6264 5416 -6016
rect 5576 -6016 5588 -5980
rect 5622 -5664 5636 -5640
rect 5796 -5640 5856 -5480
rect 5926 -5496 5932 -5436
rect 5992 -5496 5998 -5436
rect 5622 -5980 5628 -5664
rect 5796 -5676 5806 -5640
rect 5622 -6016 5636 -5980
rect 5452 -6075 5540 -6069
rect 5452 -6109 5464 -6075
rect 5528 -6109 5540 -6075
rect 5452 -6115 5540 -6109
rect 5350 -6324 5356 -6264
rect 5416 -6324 5422 -6264
rect 5240 -6422 5246 -6362
rect 5306 -6422 5312 -6362
rect 5246 -6479 5306 -6422
rect 5234 -6485 5322 -6479
rect 5234 -6519 5246 -6485
rect 5310 -6519 5322 -6485
rect 5234 -6525 5322 -6519
rect 5138 -6604 5152 -6578
rect 4968 -6920 4974 -6618
rect 4968 -6954 4982 -6920
rect 4798 -7013 4886 -7007
rect 4798 -7047 4810 -7013
rect 4874 -7047 4886 -7013
rect 4798 -7053 4886 -7047
rect 4696 -7158 4702 -7098
rect 4762 -7158 4768 -7098
rect 4922 -7196 4982 -6954
rect 5146 -6954 5152 -6604
rect 5186 -6604 5198 -6578
rect 5356 -6578 5416 -6324
rect 5462 -6362 5522 -6115
rect 5576 -6160 5636 -6016
rect 5800 -6016 5806 -5676
rect 5840 -5676 5856 -5640
rect 5840 -6016 5846 -5676
rect 5800 -6028 5846 -6016
rect 5670 -6075 5758 -6069
rect 5670 -6109 5682 -6075
rect 5746 -6109 5758 -6075
rect 5670 -6115 5758 -6109
rect 5570 -6220 5576 -6160
rect 5636 -6220 5642 -6160
rect 5456 -6422 5462 -6362
rect 5522 -6422 5856 -6362
rect 5462 -6479 5522 -6422
rect 5452 -6485 5540 -6479
rect 5452 -6519 5464 -6485
rect 5528 -6519 5540 -6485
rect 5452 -6525 5540 -6519
rect 5186 -6954 5192 -6604
rect 5356 -6606 5370 -6578
rect 5364 -6920 5370 -6606
rect 5146 -6966 5192 -6954
rect 5356 -6954 5370 -6920
rect 5404 -6606 5416 -6578
rect 5574 -6578 5634 -6422
rect 5682 -6479 5742 -6422
rect 5670 -6485 5758 -6479
rect 5670 -6519 5682 -6485
rect 5746 -6519 5758 -6485
rect 5670 -6525 5758 -6519
rect 5574 -6596 5588 -6578
rect 5404 -6920 5410 -6606
rect 5582 -6920 5588 -6596
rect 5404 -6954 5416 -6920
rect 5016 -7013 5104 -7007
rect 5016 -7047 5028 -7013
rect 5092 -7047 5104 -7013
rect 5016 -7053 5104 -7047
rect 5234 -7013 5322 -7007
rect 5234 -7047 5246 -7013
rect 5310 -7047 5322 -7013
rect 5234 -7053 5322 -7047
rect 5356 -7196 5416 -6954
rect 5576 -6954 5588 -6920
rect 5622 -6596 5634 -6578
rect 5796 -6578 5856 -6422
rect 5622 -6920 5628 -6596
rect 5796 -6600 5806 -6578
rect 5622 -6954 5636 -6920
rect 5452 -7013 5540 -7007
rect 5452 -7047 5464 -7013
rect 5528 -7047 5540 -7013
rect 5452 -7053 5540 -7047
rect 5576 -7098 5636 -6954
rect 5800 -6954 5806 -6600
rect 5840 -6600 5856 -6578
rect 5840 -6954 5846 -6600
rect 5800 -6966 5846 -6954
rect 5670 -7013 5758 -7007
rect 5670 -7047 5682 -7013
rect 5746 -7047 5758 -7013
rect 5670 -7053 5758 -7047
rect 5932 -7098 5992 -5496
rect 5570 -7158 5576 -7098
rect 5636 -7158 5642 -7098
rect 5926 -7158 5932 -7098
rect 5992 -7158 5998 -7098
rect 4042 -7256 4048 -7196
rect 4108 -7256 4114 -7196
rect 4478 -7256 4484 -7196
rect 4544 -7256 4550 -7196
rect 4916 -7256 4922 -7196
rect 4982 -7256 4988 -7196
rect 5350 -7256 5356 -7196
rect 5416 -7256 5422 -7196
rect 3486 -7374 3492 -7314
rect 3552 -7374 3558 -7314
rect 3616 -7376 4002 -7316
rect 3616 -7516 3676 -7376
rect 3722 -7417 3782 -7376
rect 3708 -7423 3796 -7417
rect 3708 -7457 3720 -7423
rect 3784 -7457 3796 -7423
rect 3708 -7463 3796 -7457
rect 3616 -7546 3626 -7516
rect 3620 -7892 3626 -7546
rect 3660 -7546 3676 -7516
rect 3832 -7516 3892 -7376
rect 3942 -7417 4002 -7376
rect 3926 -7423 4014 -7417
rect 3926 -7457 3938 -7423
rect 4002 -7457 4014 -7423
rect 3926 -7463 4014 -7457
rect 3832 -7540 3844 -7516
rect 3660 -7892 3666 -7546
rect 3838 -7864 3844 -7540
rect 3620 -7904 3666 -7892
rect 3832 -7892 3844 -7864
rect 3878 -7540 3892 -7516
rect 4048 -7516 4108 -7256
rect 4152 -7374 4158 -7314
rect 4218 -7374 4224 -7314
rect 4260 -7374 4266 -7314
rect 4326 -7374 4332 -7314
rect 4368 -7374 4374 -7314
rect 4434 -7374 4440 -7314
rect 4158 -7417 4218 -7374
rect 4144 -7423 4232 -7417
rect 4144 -7457 4156 -7423
rect 4220 -7457 4232 -7423
rect 4144 -7463 4232 -7457
rect 3878 -7864 3884 -7540
rect 4048 -7544 4062 -7516
rect 3878 -7892 3892 -7864
rect 3708 -7951 3796 -7945
rect 3708 -7985 3720 -7951
rect 3784 -7985 3796 -7951
rect 3708 -7991 3796 -7985
rect 3832 -8034 3892 -7892
rect 4056 -7892 4062 -7544
rect 4096 -7544 4108 -7516
rect 4266 -7516 4326 -7374
rect 4374 -7417 4434 -7374
rect 4362 -7423 4450 -7417
rect 4362 -7457 4374 -7423
rect 4438 -7457 4450 -7423
rect 4362 -7463 4450 -7457
rect 4266 -7540 4280 -7516
rect 4096 -7892 4102 -7544
rect 4056 -7904 4102 -7892
rect 4274 -7892 4280 -7540
rect 4314 -7540 4326 -7516
rect 4484 -7516 4544 -7256
rect 4580 -7423 4668 -7417
rect 4580 -7457 4592 -7423
rect 4656 -7457 4668 -7423
rect 4580 -7463 4668 -7457
rect 4798 -7423 4886 -7417
rect 4798 -7457 4810 -7423
rect 4874 -7457 4886 -7423
rect 4798 -7463 4886 -7457
rect 4314 -7892 4320 -7540
rect 4484 -7546 4498 -7516
rect 4274 -7904 4320 -7892
rect 4492 -7892 4498 -7546
rect 4532 -7546 4544 -7516
rect 4710 -7516 4756 -7504
rect 4532 -7892 4538 -7546
rect 4710 -7862 4716 -7516
rect 4492 -7904 4538 -7892
rect 4702 -7892 4716 -7862
rect 4750 -7862 4756 -7516
rect 4922 -7516 4982 -7256
rect 5014 -7374 5020 -7314
rect 5080 -7374 5086 -7314
rect 5132 -7374 5138 -7314
rect 5198 -7374 5204 -7314
rect 5241 -7374 5247 -7316
rect 5305 -7374 5311 -7316
rect 5020 -7417 5080 -7374
rect 5016 -7423 5104 -7417
rect 5016 -7457 5028 -7423
rect 5092 -7457 5104 -7423
rect 5016 -7463 5104 -7457
rect 4922 -7550 4934 -7516
rect 4750 -7892 4762 -7862
rect 3926 -7951 4014 -7945
rect 3926 -7985 3938 -7951
rect 4002 -7985 4014 -7951
rect 3926 -7991 3940 -7985
rect 3942 -7991 4014 -7985
rect 4144 -7951 4232 -7945
rect 4144 -7985 4156 -7951
rect 4220 -7985 4232 -7951
rect 4144 -7991 4232 -7985
rect 4362 -7951 4450 -7945
rect 4362 -7985 4374 -7951
rect 4438 -7985 4450 -7951
rect 4362 -7991 4450 -7985
rect 4580 -7951 4668 -7945
rect 4580 -7991 4592 -7951
rect 4656 -7985 4668 -7951
rect 4596 -7991 4668 -7985
rect 3942 -8034 4002 -7991
rect 4596 -8034 4656 -7991
rect 4702 -8034 4762 -7892
rect 4928 -7892 4934 -7550
rect 4968 -7550 4982 -7516
rect 5138 -7516 5198 -7374
rect 5247 -7417 5305 -7374
rect 5234 -7423 5322 -7417
rect 5234 -7457 5246 -7423
rect 5310 -7457 5322 -7423
rect 5234 -7463 5322 -7457
rect 4968 -7892 4974 -7550
rect 5138 -7556 5152 -7516
rect 4928 -7904 4974 -7892
rect 5146 -7892 5152 -7556
rect 5186 -7556 5198 -7516
rect 5356 -7516 5416 -7256
rect 5576 -7366 5856 -7306
rect 5452 -7423 5540 -7417
rect 5452 -7457 5464 -7423
rect 5528 -7457 5540 -7423
rect 5452 -7463 5540 -7457
rect 5356 -7538 5370 -7516
rect 5186 -7892 5192 -7556
rect 5146 -7904 5192 -7892
rect 5364 -7892 5370 -7538
rect 5404 -7538 5416 -7516
rect 5576 -7516 5636 -7366
rect 5682 -7417 5742 -7366
rect 5670 -7423 5758 -7417
rect 5670 -7457 5682 -7423
rect 5746 -7457 5758 -7423
rect 5670 -7463 5758 -7457
rect 5404 -7892 5410 -7538
rect 5576 -7540 5588 -7516
rect 5582 -7858 5588 -7540
rect 5364 -7904 5410 -7892
rect 5576 -7892 5588 -7858
rect 5622 -7540 5636 -7516
rect 5796 -7516 5856 -7366
rect 5622 -7858 5628 -7540
rect 5796 -7544 5806 -7516
rect 5622 -7892 5636 -7858
rect 4798 -7951 4886 -7945
rect 4798 -7985 4810 -7951
rect 4798 -7991 4872 -7985
rect 4874 -7991 4886 -7951
rect 5016 -7951 5104 -7945
rect 5016 -7985 5028 -7951
rect 5092 -7985 5104 -7951
rect 5016 -7991 5104 -7985
rect 5234 -7951 5322 -7945
rect 5234 -7985 5246 -7951
rect 5310 -7985 5322 -7951
rect 5234 -7991 5322 -7985
rect 5452 -7951 5540 -7945
rect 5452 -7985 5464 -7951
rect 5528 -7985 5540 -7951
rect 5452 -7991 5540 -7985
rect 4812 -8034 4872 -7991
rect 5464 -8034 5524 -7991
rect 5576 -8034 5636 -7892
rect 5800 -7892 5806 -7544
rect 5840 -7544 5856 -7516
rect 5840 -7892 5846 -7544
rect 5800 -7904 5846 -7892
rect 5670 -7951 5758 -7945
rect 5670 -7985 5682 -7951
rect 5746 -7985 5758 -7951
rect 5670 -7991 5758 -7985
rect 6048 -8034 6108 -4562
rect 6802 -5608 6862 -3486
rect 6796 -5668 6802 -5608
rect 6862 -5668 6868 -5608
rect 6916 -5712 6976 -3364
rect 7312 -3404 7372 -3028
rect 9526 -3114 9590 -2744
rect 10032 -2752 10092 -2480
rect 10546 -2570 10610 -2396
rect 10540 -2630 10546 -2570
rect 10606 -2630 10612 -2570
rect 11074 -2752 11134 -2480
rect 10032 -2812 11134 -2752
rect 9520 -3178 9526 -3114
rect 9590 -3178 9596 -3114
rect 10032 -3216 10092 -2812
rect 9494 -3276 10092 -3216
rect 7306 -3464 7312 -3404
rect 7372 -3464 7378 -3404
rect 8472 -3464 8478 -3404
rect 8538 -3464 8544 -3404
rect 7038 -4510 7044 -4450
rect 7104 -4510 7110 -4450
rect 6910 -5772 6916 -5712
rect 6976 -5772 6982 -5712
rect 3826 -8094 3832 -8034
rect 3892 -8094 3898 -8034
rect 3936 -8094 3942 -8034
rect 4002 -8094 4008 -8034
rect 4590 -8094 4596 -8034
rect 4656 -8094 4662 -8034
rect 4696 -8094 4702 -8034
rect 4762 -8094 4768 -8034
rect 4806 -8094 4812 -8034
rect 4872 -8094 4878 -8034
rect 5458 -8094 5464 -8034
rect 5524 -8094 5530 -8034
rect 5570 -8094 5576 -8034
rect 5636 -8094 5642 -8034
rect 6042 -8094 6048 -8034
rect 6108 -8094 6114 -8034
rect 7044 -8122 7104 -4510
rect 7174 -4608 7180 -4548
rect 7240 -4608 7246 -4548
rect 7038 -8182 7044 -8122
rect 7104 -8182 7110 -8122
rect 7180 -8252 7240 -4608
rect 7312 -7072 7372 -3464
rect 8478 -3644 8538 -3464
rect 9494 -3664 9554 -3276
rect 11564 -3304 11624 -2372
rect 14618 -2376 14678 -2374
rect 12580 -2388 12640 -2386
rect 12580 -2566 12644 -2388
rect 12040 -2574 12100 -2568
rect 11558 -3364 11564 -3304
rect 11624 -3364 11630 -3304
rect 10508 -3464 10514 -3404
rect 10574 -3464 10580 -3404
rect 10514 -3642 10574 -3464
rect 12040 -3562 12100 -2634
rect 12548 -2570 12644 -2566
rect 12548 -2572 12580 -2570
rect 12640 -2630 12646 -2570
rect 13034 -2630 13040 -2570
rect 13100 -2630 13106 -2570
rect 7460 -4352 7520 -4158
rect 7974 -4352 8034 -4256
rect 8476 -4352 8536 -4170
rect 7460 -4412 8536 -4352
rect 8476 -4718 8482 -4658
rect 8542 -4718 8548 -4658
rect 8482 -4900 8542 -4718
rect 8966 -4816 9026 -4248
rect 9496 -4352 9556 -4170
rect 9490 -4412 9496 -4352
rect 9556 -4412 9562 -4352
rect 9496 -4548 9556 -4412
rect 9490 -4608 9496 -4548
rect 9556 -4608 9562 -4548
rect 10004 -4821 10064 -4247
rect 10510 -4606 10516 -4546
rect 10576 -4606 10582 -4546
rect 10516 -4658 10576 -4606
rect 10510 -4718 10516 -4658
rect 10576 -4718 10582 -4658
rect 10516 -4896 10576 -4718
rect 11010 -4821 11070 -4247
rect 11532 -4352 11592 -4166
rect 12042 -4348 12102 -4252
rect 12548 -4348 12608 -2632
rect 13040 -3558 13100 -2630
rect 13598 -2818 13662 -2388
rect 14618 -2562 14682 -2376
rect 16654 -2380 16714 -2378
rect 14084 -2568 14144 -2562
rect 13592 -2882 13598 -2818
rect 13662 -2882 13668 -2818
rect 13598 -3102 13662 -2882
rect 13598 -3172 13662 -3166
rect 14084 -3572 14144 -2628
rect 14586 -2568 14682 -2562
rect 14646 -2572 14682 -2568
rect 15100 -2568 15160 -2562
rect 14586 -2632 14618 -2628
rect 14678 -2632 14684 -2572
rect 13062 -4348 13122 -4256
rect 13568 -4348 13628 -4170
rect 14072 -4348 14132 -4254
rect 14586 -4348 14646 -2632
rect 15100 -3562 15160 -2628
rect 15634 -2818 15698 -2384
rect 16128 -2568 16188 -2562
rect 16654 -2568 16718 -2380
rect 18690 -2392 18750 -2390
rect 15628 -2882 15634 -2818
rect 15698 -2882 15704 -2818
rect 16128 -3562 16188 -2628
rect 16622 -2572 16718 -2568
rect 16622 -2574 16654 -2572
rect 16714 -2632 16720 -2572
rect 17150 -2578 17210 -2572
rect 15094 -4348 15154 -4256
rect 15602 -4348 15662 -4168
rect 16116 -4348 16176 -4256
rect 16622 -4348 16682 -2634
rect 17150 -3566 17210 -2638
rect 17638 -2574 17698 -2568
rect 17142 -4348 17202 -4255
rect 17638 -4348 17698 -2634
rect 18150 -2578 18210 -2572
rect 18690 -2574 18754 -2392
rect 18684 -2634 18690 -2574
rect 18750 -2634 18756 -2574
rect 18150 -3572 18210 -2638
rect 19706 -2680 19770 -2386
rect 20724 -2392 20784 -2390
rect 20724 -2574 20788 -2392
rect 20718 -2634 20724 -2574
rect 20784 -2634 20790 -2574
rect 19700 -2744 19706 -2680
rect 19770 -2744 19776 -2680
rect 21742 -2818 21806 -2390
rect 21736 -2882 21742 -2818
rect 21806 -2882 21812 -2818
rect 21714 -3098 21774 -3092
rect 21714 -3400 21774 -3158
rect 22884 -3104 22944 -354
rect 22884 -3170 22944 -3164
rect 18654 -3464 18660 -3404
rect 18720 -3464 18726 -3404
rect 20688 -3464 20694 -3404
rect 20754 -3464 20760 -3404
rect 21714 -3460 22790 -3400
rect 18660 -3646 18720 -3464
rect 20694 -3642 20754 -3464
rect 21714 -3654 21774 -3460
rect 22228 -3556 22288 -3460
rect 22730 -3642 22790 -3460
rect 23132 -3464 23138 -3404
rect 23198 -3464 23204 -3404
rect 18154 -4348 18214 -4258
rect 11526 -4412 11532 -4352
rect 11592 -4412 11598 -4352
rect 12042 -4408 18214 -4348
rect 12548 -4508 12608 -4408
rect 17638 -4508 17698 -4408
rect 12548 -4568 17698 -4508
rect 12548 -4918 12608 -4568
rect 13566 -4720 13572 -4660
rect 13632 -4720 13638 -4660
rect 14076 -4706 15134 -4646
rect 13572 -4902 13632 -4720
rect 14076 -4818 14136 -4706
rect 15076 -4744 15134 -4706
rect 15600 -4720 15606 -4660
rect 15666 -4720 15672 -4660
rect 15076 -4818 15136 -4744
rect 15606 -4904 15666 -4720
rect 17638 -4894 17698 -4568
rect 18656 -4720 18662 -4660
rect 18722 -4720 18728 -4660
rect 18662 -4902 18722 -4720
rect 19162 -4821 19222 -4247
rect 19676 -4352 19736 -4170
rect 19670 -4412 19676 -4352
rect 19736 -4412 19742 -4352
rect 20186 -4821 20246 -4247
rect 20690 -4720 20696 -4660
rect 20756 -4720 20762 -4660
rect 20696 -4898 20756 -4720
rect 21192 -4815 21252 -4241
rect 21712 -4352 21772 -4166
rect 21706 -4412 21712 -4352
rect 21772 -4412 21778 -4352
rect 22972 -4606 22978 -4546
rect 23038 -4606 23044 -4546
rect 21714 -4714 22790 -4654
rect 21714 -4908 21774 -4714
rect 22228 -4810 22288 -4714
rect 22730 -4896 22790 -4714
rect 7464 -5608 7524 -5414
rect 7978 -5608 8038 -5512
rect 8480 -5608 8540 -5426
rect 7464 -5668 8540 -5608
rect 7462 -5970 8538 -5910
rect 7462 -6164 7522 -5970
rect 7976 -6066 8036 -5970
rect 8478 -6152 8538 -5970
rect 8960 -6076 9020 -5502
rect 9498 -5712 9558 -5424
rect 9498 -5778 9558 -5772
rect 9492 -5976 9498 -5916
rect 9558 -5976 9564 -5916
rect 9498 -6154 9558 -5976
rect 9998 -6077 10058 -5502
rect 11004 -6077 11064 -5502
rect 11534 -5712 11594 -5420
rect 12054 -5604 12114 -5511
rect 12550 -5604 12610 -5420
rect 13066 -5604 13126 -5514
rect 12054 -5664 13126 -5604
rect 11528 -5772 11534 -5712
rect 11594 -5772 11600 -5712
rect 11526 -5874 11532 -5814
rect 11592 -5874 11598 -5814
rect 11532 -5916 11592 -5874
rect 11526 -5976 11532 -5916
rect 11592 -5976 11598 -5916
rect 11532 -6158 11592 -5976
rect 12550 -6168 12610 -5664
rect 13562 -5668 13568 -5608
rect 13628 -5668 13634 -5608
rect 13568 -6154 13628 -5668
rect 14070 -6082 14130 -5508
rect 14588 -5608 14648 -5426
rect 14582 -5668 14588 -5608
rect 14648 -5668 14654 -5608
rect 14582 -5974 14588 -5914
rect 14648 -5974 14654 -5914
rect 14588 -6152 14648 -5974
rect 15100 -6070 15160 -5496
rect 15606 -5914 15666 -5422
rect 15600 -5974 15606 -5914
rect 15666 -5974 15672 -5914
rect 16112 -6070 16172 -5496
rect 16624 -5608 16684 -5422
rect 17142 -5606 17202 -5513
rect 17638 -5606 17698 -5422
rect 18154 -5606 18214 -5516
rect 16618 -5668 16624 -5608
rect 16684 -5668 16690 -5608
rect 17142 -5666 18214 -5606
rect 16616 -5974 16622 -5914
rect 16682 -5974 16688 -5914
rect 16622 -6156 16682 -5974
rect 17638 -6160 17698 -5666
rect 18652 -5772 18658 -5712
rect 18718 -5772 18724 -5712
rect 18658 -6162 18718 -5772
rect 19156 -6077 19216 -5502
rect 19520 -5654 19526 -5594
rect 19586 -5654 19592 -5594
rect 19526 -5914 19586 -5654
rect 19674 -5704 19734 -5414
rect 19668 -5764 19674 -5704
rect 19734 -5764 19740 -5704
rect 19520 -5974 19526 -5914
rect 19586 -5974 19592 -5914
rect 19672 -5972 19678 -5912
rect 19738 -5972 19744 -5912
rect 19678 -6150 19738 -5972
rect 20180 -6077 20240 -5502
rect 20694 -5814 20754 -5422
rect 20688 -5874 20694 -5814
rect 20754 -5874 20760 -5814
rect 21186 -6071 21246 -5496
rect 21714 -5704 21774 -5410
rect 21708 -5764 21714 -5704
rect 21774 -5764 21780 -5704
rect 22840 -5764 22846 -5704
rect 22906 -5764 22912 -5704
rect 21706 -5972 21712 -5912
rect 21772 -5972 21778 -5912
rect 21712 -6154 21772 -5972
rect 8480 -6864 8540 -6678
rect 8474 -6924 8480 -6864
rect 8540 -6924 8546 -6864
rect 7306 -7132 7312 -7072
rect 7372 -7132 7378 -7072
rect 7462 -7230 8538 -7170
rect 7462 -7424 7522 -7230
rect 7976 -7326 8036 -7230
rect 8478 -7412 8538 -7230
rect 8972 -7326 9032 -6752
rect 9488 -7234 9494 -7174
rect 9554 -7234 9560 -7174
rect 9494 -7412 9554 -7234
rect 10010 -7326 10070 -6752
rect 10516 -6864 10576 -6682
rect 10510 -6924 10516 -6864
rect 10576 -6924 10582 -6864
rect 10516 -6972 10576 -6924
rect 10510 -7032 10516 -6972
rect 10576 -7032 10582 -6972
rect 11016 -7022 11076 -6752
rect 12052 -6856 12112 -6763
rect 12548 -6856 12608 -6672
rect 13064 -6856 13124 -6766
rect 12052 -6916 13124 -6856
rect 13570 -6862 13630 -6676
rect 11016 -7082 11792 -7022
rect 11016 -7326 11076 -7082
rect 11732 -7168 11792 -7082
rect 11522 -7234 11528 -7174
rect 11588 -7234 11594 -7174
rect 11726 -7228 11732 -7168
rect 11792 -7228 11798 -7168
rect 11528 -7416 11588 -7234
rect 12548 -7444 12608 -6916
rect 13564 -6922 13570 -6862
rect 13630 -6922 13636 -6862
rect 14080 -6994 14140 -6764
rect 15096 -6994 15156 -6756
rect 15606 -6862 15666 -6680
rect 15600 -6922 15606 -6862
rect 15666 -6922 15672 -6862
rect 16110 -6994 16170 -6760
rect 17140 -6858 17200 -6765
rect 17636 -6858 17696 -6674
rect 18152 -6858 18212 -6768
rect 17140 -6918 18212 -6858
rect 18660 -6860 18720 -6674
rect 14080 -7054 16894 -6994
rect 13566 -7168 13626 -7162
rect 14080 -7168 14140 -7054
rect 13626 -7228 14140 -7168
rect 13566 -7234 13626 -7228
rect 14580 -7232 14586 -7172
rect 14646 -7232 14652 -7172
rect 16614 -7232 16620 -7172
rect 16680 -7232 16686 -7172
rect 16834 -7176 16894 -7054
rect 14586 -7410 14646 -7232
rect 16620 -7414 16680 -7232
rect 16828 -7236 16834 -7176
rect 16894 -7236 16900 -7176
rect 17636 -7424 17696 -6918
rect 18654 -6920 18660 -6860
rect 18720 -6920 18726 -6860
rect 19168 -7170 19228 -6752
rect 19168 -7176 19230 -7170
rect 19168 -7236 19170 -7176
rect 19676 -7234 19682 -7174
rect 19742 -7234 19748 -7174
rect 19168 -7242 19230 -7236
rect 19168 -7326 19228 -7242
rect 19682 -7412 19742 -7234
rect 20192 -7326 20252 -6752
rect 20696 -6860 20756 -6678
rect 20690 -6920 20696 -6860
rect 20756 -6920 20762 -6860
rect 21198 -7320 21258 -6746
rect 21712 -6864 21772 -6670
rect 22226 -6864 22286 -6768
rect 22728 -6864 22788 -6682
rect 21712 -6924 22788 -6864
rect 22846 -6972 22906 -5764
rect 22978 -5912 23038 -4606
rect 22972 -5972 22978 -5912
rect 23038 -5972 23044 -5912
rect 22840 -7032 22846 -6972
rect 22906 -7032 22912 -6972
rect 21710 -7234 21716 -7174
rect 21776 -7234 21782 -7174
rect 21716 -7416 21776 -7234
rect 8476 -8122 8536 -7936
rect 8470 -8182 8476 -8122
rect 8536 -8182 8542 -8122
rect 8984 -8236 9044 -8024
rect 10008 -8236 10068 -8016
rect 10512 -8122 10572 -7940
rect 10506 -8182 10512 -8122
rect 10572 -8182 10578 -8122
rect 11014 -8236 11074 -8016
rect 7174 -8312 7180 -8252
rect 7240 -8312 7246 -8252
rect 8984 -8296 11074 -8236
rect 2104 -8452 2110 -8392
rect 2170 -8452 2176 -8392
rect 1954 -8498 2014 -8492
rect 7180 -8498 7240 -8312
rect 2014 -8558 7240 -8498
rect 1954 -8564 2014 -8558
rect 1184 -8616 1244 -8610
rect 8984 -8616 9044 -8296
rect 11014 -8546 11074 -8296
rect 11534 -8392 11594 -7926
rect 12052 -8116 12112 -8021
rect 12548 -8116 12608 -7930
rect 13064 -8116 13124 -8024
rect 13570 -8116 13630 -7918
rect 14080 -8116 14140 -8024
rect 14586 -8116 14646 -7938
rect 15096 -8116 15156 -8024
rect 15604 -8116 15664 -7924
rect 16106 -8116 16166 -8024
rect 16622 -8116 16682 -7934
rect 17140 -8116 17200 -8023
rect 17636 -8116 17696 -7932
rect 18152 -8116 18212 -8026
rect 12052 -8176 18212 -8116
rect 18664 -8122 18724 -7936
rect 18658 -8182 18664 -8122
rect 18724 -8182 18730 -8122
rect 19172 -8234 19232 -8008
rect 20192 -8234 20252 -8016
rect 20700 -8122 20760 -7940
rect 20694 -8182 20700 -8122
rect 20760 -8182 20766 -8122
rect 21194 -8234 21254 -8016
rect 21714 -8118 21774 -7924
rect 22228 -8118 22288 -8022
rect 22730 -8118 22790 -7936
rect 21714 -8178 22790 -8118
rect 19172 -8294 21254 -8234
rect 11528 -8452 11534 -8392
rect 11594 -8452 11600 -8392
rect 19172 -8546 19232 -8294
rect 23138 -8392 23198 -3464
rect 24716 -8262 24722 1102
rect 24822 -8262 24828 1102
rect 23132 -8452 23138 -8392
rect 23198 -8452 23204 -8392
rect 11014 -8606 19232 -8546
rect 1244 -8676 9044 -8616
rect 1184 -8682 1244 -8676
rect 24716 -8776 24828 -8262
rect 372 -8782 24828 -8776
rect 372 -8882 478 -8782
rect 24722 -8882 24828 -8782
rect 372 -8888 24828 -8882
rect -645 -11172 -523 -11167
rect -12328 -11176 24928 -11172
rect -12328 -11178 -5038 -11176
rect -4938 -11178 -2438 -11176
rect -2338 -11178 -634 -11176
rect -534 -11178 24928 -11176
rect -12328 -11278 -12222 -11178
rect 24822 -11278 24928 -11178
rect -12328 -11284 24928 -11278
rect -12328 -12070 -12216 -11284
rect 1948 -11408 1954 -11348
rect 2014 -11408 2020 -11348
rect 2104 -11408 2110 -11348
rect 2170 -11408 2176 -11348
rect 2336 -11356 2396 -11350
rect -12328 -26330 -12322 -12070
rect -12222 -26330 -12216 -12070
rect 1954 -12186 2014 -11408
rect -2072 -12246 2014 -12186
rect -2072 -12324 -2012 -12246
rect -9196 -12384 -2012 -12324
rect -9196 -12524 -9136 -12384
rect -8686 -12434 -8626 -12384
rect -8902 -12440 -8414 -12434
rect -8902 -12474 -8890 -12440
rect -8426 -12474 -8414 -12440
rect -8902 -12480 -8414 -12474
rect -9196 -12554 -9184 -12524
rect -9190 -13082 -9184 -12554
rect -9200 -13100 -9184 -13082
rect -9150 -12554 -9136 -12524
rect -8180 -12524 -8120 -12384
rect -7678 -12434 -7618 -12384
rect -6650 -12434 -6590 -12384
rect -7884 -12440 -7396 -12434
rect -7884 -12474 -7872 -12440
rect -7408 -12474 -7396 -12440
rect -7884 -12480 -7396 -12474
rect -6866 -12440 -6378 -12434
rect -6866 -12474 -6854 -12440
rect -6390 -12474 -6378 -12440
rect -6866 -12480 -6378 -12474
rect -8180 -12548 -8166 -12524
rect -9150 -13082 -9144 -12554
rect -8172 -13078 -8166 -12548
rect -9150 -13100 -9140 -13082
rect -9200 -13342 -9140 -13100
rect -8180 -13100 -8166 -13078
rect -8132 -12548 -8120 -12524
rect -7154 -12524 -7108 -12512
rect -8132 -13078 -8126 -12548
rect -7154 -13076 -7148 -12524
rect -8132 -13100 -8120 -13078
rect -8902 -13150 -8414 -13144
rect -8902 -13184 -8890 -13150
rect -8426 -13184 -8414 -13150
rect -8902 -13190 -8414 -13184
rect -8686 -13252 -8626 -13190
rect -8902 -13258 -8414 -13252
rect -8902 -13292 -8890 -13258
rect -8426 -13292 -8414 -13258
rect -8902 -13298 -8414 -13292
rect -9200 -13372 -9184 -13342
rect -9190 -13896 -9184 -13372
rect -9198 -13918 -9184 -13896
rect -9150 -13372 -9140 -13342
rect -8180 -13342 -8120 -13100
rect -7160 -13100 -7148 -13076
rect -7114 -13076 -7108 -12524
rect -6142 -12524 -6082 -12384
rect -5636 -12434 -5576 -12384
rect -4622 -12434 -4562 -12384
rect -5848 -12440 -5360 -12434
rect -5848 -12474 -5836 -12440
rect -5372 -12474 -5360 -12440
rect -5848 -12480 -5360 -12474
rect -4830 -12440 -4342 -12434
rect -4830 -12474 -4818 -12440
rect -4354 -12474 -4342 -12440
rect -4830 -12480 -4342 -12474
rect -6142 -12562 -6130 -12524
rect -7114 -13100 -7100 -13076
rect -6136 -13080 -6130 -12562
rect -7884 -13150 -7396 -13144
rect -7884 -13184 -7872 -13150
rect -7408 -13184 -7396 -13150
rect -7884 -13190 -7396 -13184
rect -7682 -13252 -7622 -13190
rect -7884 -13258 -7396 -13252
rect -7884 -13292 -7872 -13258
rect -7408 -13292 -7396 -13258
rect -7884 -13298 -7396 -13292
rect -8180 -13368 -8166 -13342
rect -9150 -13896 -9144 -13372
rect -8172 -13892 -8166 -13368
rect -9150 -13918 -9138 -13896
rect -9198 -14160 -9138 -13918
rect -8178 -13918 -8166 -13892
rect -8132 -13368 -8120 -13342
rect -7160 -13342 -7100 -13100
rect -6142 -13100 -6130 -13080
rect -6096 -12562 -6082 -12524
rect -5118 -12524 -5072 -12512
rect -4106 -12524 -4046 -12384
rect -3590 -12434 -3530 -12384
rect -2584 -12434 -2524 -12384
rect -3812 -12440 -3324 -12434
rect -3812 -12474 -3800 -12440
rect -3336 -12474 -3324 -12440
rect -3812 -12480 -3324 -12474
rect -2794 -12440 -2306 -12434
rect -2794 -12474 -2782 -12440
rect -2318 -12474 -2306 -12440
rect -2794 -12480 -2306 -12474
rect -6096 -13080 -6090 -12562
rect -5118 -13072 -5112 -12524
rect -6096 -13100 -6082 -13080
rect -6866 -13150 -6378 -13144
rect -6866 -13184 -6854 -13150
rect -6390 -13184 -6378 -13150
rect -6866 -13190 -6378 -13184
rect -6652 -13252 -6592 -13190
rect -6866 -13258 -6378 -13252
rect -6866 -13292 -6854 -13258
rect -6390 -13292 -6378 -13258
rect -6866 -13298 -6378 -13292
rect -7160 -13366 -7148 -13342
rect -8132 -13892 -8126 -13368
rect -7154 -13890 -7148 -13366
rect -8132 -13918 -8118 -13892
rect -8902 -13968 -8414 -13962
rect -8902 -14002 -8890 -13968
rect -8426 -14002 -8414 -13968
rect -8902 -14008 -8414 -14002
rect -8686 -14070 -8626 -14008
rect -8902 -14076 -8414 -14070
rect -8902 -14110 -8890 -14076
rect -8426 -14110 -8414 -14076
rect -8902 -14116 -8414 -14110
rect -9198 -14186 -9184 -14160
rect -9190 -14724 -9184 -14186
rect -9198 -14736 -9184 -14724
rect -9150 -14186 -9138 -14160
rect -8178 -14160 -8118 -13918
rect -7158 -13918 -7148 -13890
rect -7114 -13366 -7100 -13342
rect -6142 -13342 -6082 -13100
rect -5122 -13100 -5112 -13072
rect -5078 -13072 -5072 -12524
rect -4108 -12558 -4094 -12524
rect -4106 -12570 -4094 -12558
rect -5078 -13100 -5062 -13072
rect -4100 -13080 -4094 -12570
rect -5848 -13150 -5360 -13144
rect -5848 -13184 -5836 -13150
rect -5372 -13184 -5360 -13150
rect -5848 -13190 -5360 -13184
rect -5650 -13252 -5590 -13190
rect -5848 -13258 -5360 -13252
rect -5848 -13292 -5836 -13258
rect -5372 -13292 -5360 -13258
rect -5848 -13298 -5360 -13292
rect -7114 -13890 -7108 -13366
rect -6142 -13370 -6130 -13342
rect -7114 -13918 -7098 -13890
rect -6136 -13894 -6130 -13370
rect -7884 -13968 -7396 -13962
rect -7884 -14002 -7872 -13968
rect -7408 -14002 -7396 -13968
rect -7884 -14008 -7396 -14002
rect -7670 -14070 -7610 -14008
rect -7884 -14076 -7396 -14070
rect -7884 -14110 -7872 -14076
rect -7408 -14110 -7396 -14076
rect -7884 -14116 -7396 -14110
rect -8178 -14182 -8166 -14160
rect -9150 -14724 -9144 -14186
rect -8172 -14720 -8166 -14182
rect -9150 -14736 -9138 -14724
rect -9198 -14978 -9138 -14736
rect -8178 -14736 -8166 -14720
rect -8132 -14182 -8118 -14160
rect -7158 -14160 -7098 -13918
rect -6140 -13918 -6130 -13894
rect -6096 -13370 -6082 -13342
rect -5122 -13342 -5062 -13100
rect -4110 -13100 -4094 -13080
rect -4060 -12570 -4046 -12524
rect -3082 -12524 -3036 -12512
rect -4060 -13080 -4054 -12570
rect -3082 -13080 -3076 -12524
rect -4060 -13100 -4050 -13080
rect -4830 -13150 -4342 -13144
rect -4830 -13184 -4818 -13150
rect -4354 -13184 -4342 -13150
rect -4830 -13190 -4342 -13184
rect -4620 -13252 -4560 -13190
rect -4830 -13258 -4342 -13252
rect -4830 -13292 -4818 -13258
rect -4354 -13292 -4342 -13258
rect -4830 -13298 -4342 -13292
rect -5122 -13362 -5112 -13342
rect -6096 -13894 -6090 -13370
rect -5118 -13886 -5112 -13362
rect -6096 -13918 -6080 -13894
rect -6866 -13968 -6378 -13962
rect -6866 -14002 -6854 -13968
rect -6390 -14002 -6378 -13968
rect -6866 -14008 -6378 -14002
rect -6652 -14070 -6592 -14008
rect -6866 -14076 -6378 -14070
rect -6866 -14110 -6854 -14076
rect -6390 -14110 -6378 -14076
rect -6866 -14116 -6378 -14110
rect -7158 -14180 -7148 -14160
rect -8132 -14720 -8126 -14182
rect -7154 -14718 -7148 -14180
rect -8132 -14736 -8118 -14720
rect -8902 -14786 -8414 -14780
rect -8902 -14820 -8890 -14786
rect -8426 -14820 -8414 -14786
rect -8902 -14826 -8414 -14820
rect -8692 -14888 -8632 -14826
rect -8902 -14894 -8414 -14888
rect -8902 -14928 -8890 -14894
rect -8426 -14928 -8414 -14894
rect -8902 -14934 -8414 -14928
rect -9198 -15014 -9184 -14978
rect -9190 -15536 -9184 -15014
rect -9198 -15554 -9184 -15536
rect -9150 -15014 -9138 -14978
rect -8178 -14978 -8118 -14736
rect -7158 -14736 -7148 -14718
rect -7114 -14180 -7098 -14160
rect -6140 -14160 -6080 -13918
rect -5120 -13918 -5112 -13886
rect -5078 -13362 -5062 -13342
rect -4110 -13342 -4050 -13100
rect -3088 -13100 -3076 -13080
rect -3042 -13080 -3036 -12524
rect -2072 -12524 -2012 -12384
rect -1562 -12434 -1502 -12246
rect 1184 -12334 1244 -12328
rect -32 -12394 1184 -12334
rect -1776 -12440 -1288 -12434
rect -1776 -12474 -1764 -12440
rect -1300 -12474 -1288 -12440
rect -1776 -12480 -1288 -12474
rect -758 -12440 -270 -12434
rect -758 -12474 -746 -12440
rect -282 -12474 -270 -12440
rect -758 -12480 -270 -12474
rect -2072 -12560 -2058 -12524
rect -2064 -13080 -2058 -12560
rect -3042 -13100 -3028 -13080
rect -3812 -13150 -3324 -13144
rect -3812 -13184 -3800 -13150
rect -3336 -13184 -3324 -13150
rect -3812 -13190 -3324 -13184
rect -3604 -13252 -3544 -13190
rect -3812 -13258 -3324 -13252
rect -3812 -13292 -3800 -13258
rect -3336 -13292 -3324 -13258
rect -3812 -13298 -3324 -13292
rect -5078 -13886 -5072 -13362
rect -4110 -13370 -4094 -13342
rect -5078 -13918 -5060 -13886
rect -4100 -13894 -4094 -13370
rect -5848 -13968 -5360 -13962
rect -5848 -14002 -5836 -13968
rect -5372 -14002 -5360 -13968
rect -5848 -14008 -5360 -14002
rect -5650 -14070 -5590 -14008
rect -5848 -14076 -5360 -14070
rect -5848 -14110 -5836 -14076
rect -5372 -14110 -5360 -14076
rect -5848 -14116 -5360 -14110
rect -7114 -14718 -7108 -14180
rect -6140 -14184 -6130 -14160
rect -7114 -14736 -7098 -14718
rect -6136 -14722 -6130 -14184
rect -7884 -14786 -7396 -14780
rect -7884 -14820 -7872 -14786
rect -7408 -14820 -7396 -14786
rect -7884 -14826 -7396 -14820
rect -7670 -14888 -7610 -14826
rect -7884 -14894 -7396 -14888
rect -7884 -14928 -7872 -14894
rect -7408 -14928 -7396 -14894
rect -7884 -14934 -7396 -14928
rect -8178 -15010 -8166 -14978
rect -9150 -15536 -9144 -15014
rect -8172 -15532 -8166 -15010
rect -9150 -15554 -9138 -15536
rect -9198 -15796 -9138 -15554
rect -8178 -15554 -8166 -15532
rect -8132 -15010 -8118 -14978
rect -7158 -14978 -7098 -14736
rect -6140 -14736 -6130 -14722
rect -6096 -14184 -6080 -14160
rect -5120 -14160 -5060 -13918
rect -4108 -13918 -4094 -13894
rect -4060 -13370 -4050 -13342
rect -3088 -13342 -3028 -13100
rect -2068 -13100 -2058 -13080
rect -2024 -12560 -2012 -12524
rect -1046 -12524 -1000 -12512
rect -2024 -13080 -2018 -12560
rect -1046 -13076 -1040 -12524
rect -2024 -13100 -2008 -13080
rect -2794 -13150 -2306 -13144
rect -2794 -13184 -2782 -13150
rect -2318 -13184 -2306 -13150
rect -2794 -13190 -2306 -13184
rect -2582 -13252 -2522 -13190
rect -2794 -13258 -2306 -13252
rect -2794 -13292 -2782 -13258
rect -2318 -13292 -2306 -13258
rect -2794 -13298 -2306 -13292
rect -3088 -13370 -3076 -13342
rect -4060 -13894 -4054 -13370
rect -3082 -13894 -3076 -13370
rect -4060 -13918 -4048 -13894
rect -4830 -13968 -4342 -13962
rect -4830 -14002 -4818 -13968
rect -4354 -14002 -4342 -13968
rect -4830 -14008 -4342 -14002
rect -4620 -14070 -4560 -14008
rect -4830 -14076 -4342 -14070
rect -4830 -14110 -4818 -14076
rect -4354 -14110 -4342 -14076
rect -4830 -14116 -4342 -14110
rect -5120 -14176 -5112 -14160
rect -6096 -14722 -6090 -14184
rect -5118 -14714 -5112 -14176
rect -6096 -14736 -6080 -14722
rect -6866 -14786 -6378 -14780
rect -6866 -14820 -6854 -14786
rect -6390 -14820 -6378 -14786
rect -6866 -14826 -6378 -14820
rect -6658 -14888 -6598 -14826
rect -6866 -14894 -6378 -14888
rect -6866 -14928 -6854 -14894
rect -6390 -14928 -6378 -14894
rect -6866 -14934 -6378 -14928
rect -7158 -15008 -7148 -14978
rect -8132 -15532 -8126 -15010
rect -7154 -15530 -7148 -15008
rect -8132 -15554 -8118 -15532
rect -8902 -15604 -8414 -15598
rect -8902 -15638 -8890 -15604
rect -8426 -15638 -8414 -15604
rect -8902 -15644 -8414 -15638
rect -8694 -15706 -8634 -15644
rect -8902 -15712 -8414 -15706
rect -8902 -15746 -8890 -15712
rect -8426 -15746 -8414 -15712
rect -8902 -15752 -8414 -15746
rect -9198 -15826 -9184 -15796
rect -9190 -16356 -9184 -15826
rect -9198 -16372 -9184 -16356
rect -9150 -15826 -9138 -15796
rect -8178 -15796 -8118 -15554
rect -7158 -15554 -7148 -15530
rect -7114 -15008 -7098 -14978
rect -6140 -14978 -6080 -14736
rect -5120 -14736 -5112 -14714
rect -5078 -14176 -5060 -14160
rect -4108 -14160 -4048 -13918
rect -3086 -13918 -3076 -13894
rect -3042 -13370 -3028 -13342
rect -2068 -13342 -2008 -13100
rect -1052 -13100 -1040 -13076
rect -1006 -13076 -1000 -12524
rect -32 -12524 28 -12394
rect 1184 -12400 1244 -12394
rect 1844 -12508 1850 -12448
rect 1910 -12508 1916 -12448
rect -32 -12576 -22 -12524
rect -1006 -13100 -992 -13076
rect -28 -13080 -22 -12576
rect -1776 -13150 -1288 -13144
rect -1776 -13184 -1764 -13150
rect -1300 -13184 -1288 -13150
rect -1776 -13190 -1288 -13184
rect -1570 -13252 -1510 -13190
rect -1776 -13258 -1288 -13252
rect -1776 -13292 -1764 -13258
rect -1300 -13292 -1288 -13258
rect -1776 -13298 -1288 -13292
rect -2068 -13370 -2058 -13342
rect -3042 -13894 -3036 -13370
rect -2064 -13894 -2058 -13370
rect -3042 -13918 -3026 -13894
rect -3812 -13968 -3324 -13962
rect -3812 -14002 -3800 -13968
rect -3336 -14002 -3324 -13968
rect -3812 -14008 -3324 -14002
rect -3604 -14070 -3544 -14008
rect -3812 -14076 -3324 -14070
rect -3812 -14110 -3800 -14076
rect -3336 -14110 -3324 -14076
rect -3812 -14116 -3324 -14110
rect -5078 -14714 -5072 -14176
rect -4108 -14184 -4094 -14160
rect -5078 -14736 -5060 -14714
rect -4100 -14722 -4094 -14184
rect -5848 -14786 -5360 -14780
rect -5848 -14820 -5836 -14786
rect -5372 -14820 -5360 -14786
rect -5848 -14826 -5360 -14820
rect -5656 -14888 -5596 -14826
rect -5848 -14894 -5360 -14888
rect -5848 -14928 -5836 -14894
rect -5372 -14928 -5360 -14894
rect -5848 -14934 -5360 -14928
rect -7114 -15530 -7108 -15008
rect -6140 -15012 -6130 -14978
rect -7114 -15554 -7098 -15530
rect -6136 -15534 -6130 -15012
rect -7884 -15604 -7396 -15598
rect -7884 -15638 -7872 -15604
rect -7408 -15638 -7396 -15604
rect -7884 -15644 -7396 -15638
rect -7676 -15706 -7616 -15644
rect -7884 -15712 -7396 -15706
rect -7884 -15746 -7872 -15712
rect -7408 -15746 -7396 -15712
rect -7884 -15752 -7396 -15746
rect -8178 -15822 -8166 -15796
rect -9150 -16356 -9144 -15826
rect -8172 -16352 -8166 -15822
rect -9150 -16372 -9138 -16356
rect -9198 -16614 -9138 -16372
rect -8178 -16372 -8166 -16352
rect -8132 -15822 -8118 -15796
rect -7158 -15796 -7098 -15554
rect -6140 -15554 -6130 -15534
rect -6096 -15012 -6080 -14978
rect -5120 -14978 -5060 -14736
rect -4108 -14736 -4094 -14722
rect -4060 -14184 -4048 -14160
rect -3086 -14160 -3026 -13918
rect -2066 -13918 -2058 -13894
rect -2024 -13370 -2008 -13342
rect -1052 -13342 -992 -13100
rect -30 -13100 -22 -13080
rect 12 -12576 28 -12524
rect 12 -13080 18 -12576
rect 12 -13100 30 -13080
rect -758 -13150 -270 -13144
rect -758 -13184 -746 -13150
rect -282 -13184 -270 -13150
rect -758 -13190 -270 -13184
rect -550 -13252 -490 -13190
rect -758 -13258 -270 -13252
rect -758 -13292 -746 -13258
rect -282 -13292 -270 -13258
rect -758 -13298 -270 -13292
rect -1052 -13366 -1040 -13342
rect -2024 -13894 -2018 -13370
rect -1046 -13890 -1040 -13366
rect -2024 -13918 -2006 -13894
rect -2794 -13968 -2306 -13962
rect -2794 -14002 -2782 -13968
rect -2318 -14002 -2306 -13968
rect -2794 -14008 -2306 -14002
rect -2582 -14070 -2522 -14008
rect -2794 -14076 -2306 -14070
rect -2794 -14110 -2782 -14076
rect -2318 -14110 -2306 -14076
rect -2794 -14116 -2306 -14110
rect -3086 -14184 -3076 -14160
rect -4060 -14722 -4054 -14184
rect -3082 -14722 -3076 -14184
rect -4060 -14736 -4048 -14722
rect -4830 -14786 -4342 -14780
rect -4830 -14820 -4818 -14786
rect -4354 -14820 -4342 -14786
rect -4830 -14826 -4342 -14820
rect -4626 -14888 -4566 -14826
rect -4830 -14894 -4342 -14888
rect -4830 -14928 -4818 -14894
rect -4354 -14928 -4342 -14894
rect -4830 -14934 -4342 -14928
rect -5120 -15004 -5112 -14978
rect -6096 -15534 -6090 -15012
rect -5118 -15526 -5112 -15004
rect -6096 -15554 -6080 -15534
rect -6866 -15604 -6378 -15598
rect -6866 -15638 -6854 -15604
rect -6390 -15638 -6378 -15604
rect -6866 -15644 -6378 -15638
rect -6660 -15706 -6600 -15644
rect -6866 -15712 -6378 -15706
rect -6866 -15746 -6854 -15712
rect -6390 -15746 -6378 -15712
rect -6866 -15752 -6378 -15746
rect -7158 -15820 -7148 -15796
rect -8132 -16352 -8126 -15822
rect -7154 -16350 -7148 -15820
rect -8132 -16372 -8118 -16352
rect -8902 -16422 -8414 -16416
rect -8902 -16456 -8890 -16422
rect -8426 -16456 -8414 -16422
rect -8902 -16462 -8414 -16456
rect -8692 -16524 -8632 -16462
rect -8902 -16530 -8414 -16524
rect -8902 -16564 -8890 -16530
rect -8426 -16564 -8414 -16530
rect -8902 -16570 -8414 -16564
rect -9198 -16646 -9184 -16614
rect -9190 -17168 -9184 -16646
rect -9198 -17190 -9184 -17168
rect -9150 -16646 -9138 -16614
rect -8178 -16614 -8118 -16372
rect -7158 -16372 -7148 -16350
rect -7114 -15820 -7098 -15796
rect -6140 -15796 -6080 -15554
rect -5120 -15554 -5112 -15526
rect -5078 -15004 -5060 -14978
rect -4108 -14978 -4048 -14736
rect -3086 -14736 -3076 -14722
rect -3042 -14184 -3026 -14160
rect -2066 -14160 -2006 -13918
rect -1050 -13918 -1040 -13890
rect -1006 -13366 -992 -13342
rect -30 -13342 30 -13100
rect -1006 -13890 -1000 -13366
rect -30 -13370 -22 -13342
rect -1006 -13918 -990 -13890
rect -1776 -13968 -1288 -13962
rect -1776 -14002 -1764 -13968
rect -1300 -14002 -1288 -13968
rect -1776 -14008 -1288 -14002
rect -1570 -14070 -1510 -14008
rect -1776 -14076 -1288 -14070
rect -1776 -14110 -1764 -14076
rect -1300 -14110 -1288 -14076
rect -1776 -14116 -1288 -14110
rect -2066 -14184 -2058 -14160
rect -3042 -14722 -3036 -14184
rect -2064 -14722 -2058 -14184
rect -3042 -14736 -3026 -14722
rect -3812 -14786 -3324 -14780
rect -3812 -14820 -3800 -14786
rect -3336 -14820 -3324 -14786
rect -3812 -14826 -3324 -14820
rect -3610 -14888 -3550 -14826
rect -3812 -14894 -3324 -14888
rect -3812 -14928 -3800 -14894
rect -3336 -14928 -3324 -14894
rect -3812 -14934 -3324 -14928
rect -5078 -15526 -5072 -15004
rect -4108 -15012 -4094 -14978
rect -5078 -15554 -5060 -15526
rect -4100 -15534 -4094 -15012
rect -5848 -15604 -5360 -15598
rect -5848 -15638 -5836 -15604
rect -5372 -15638 -5360 -15604
rect -5848 -15644 -5360 -15638
rect -5658 -15706 -5598 -15644
rect -5848 -15712 -5360 -15706
rect -5848 -15746 -5836 -15712
rect -5372 -15746 -5360 -15712
rect -5848 -15752 -5360 -15746
rect -7114 -16350 -7108 -15820
rect -6140 -15824 -6130 -15796
rect -7114 -16372 -7098 -16350
rect -6136 -16354 -6130 -15824
rect -7884 -16422 -7396 -16416
rect -7884 -16456 -7872 -16422
rect -7408 -16456 -7396 -16422
rect -7884 -16462 -7396 -16456
rect -7678 -16524 -7618 -16462
rect -7884 -16530 -7396 -16524
rect -7884 -16564 -7872 -16530
rect -7408 -16564 -7396 -16530
rect -7884 -16570 -7396 -16564
rect -8178 -16642 -8166 -16614
rect -9150 -17168 -9144 -16646
rect -8172 -17164 -8166 -16642
rect -9150 -17190 -9138 -17168
rect -9198 -17432 -9138 -17190
rect -8178 -17190 -8166 -17164
rect -8132 -16642 -8118 -16614
rect -7158 -16614 -7098 -16372
rect -6140 -16372 -6130 -16354
rect -6096 -15824 -6080 -15796
rect -5120 -15796 -5060 -15554
rect -4108 -15554 -4094 -15534
rect -4060 -15012 -4048 -14978
rect -3086 -14978 -3026 -14736
rect -2066 -14736 -2058 -14722
rect -2024 -14184 -2006 -14160
rect -1050 -14160 -990 -13918
rect -28 -13918 -22 -13370
rect 12 -13370 30 -13342
rect 12 -13894 18 -13370
rect 12 -13918 32 -13894
rect -758 -13968 -270 -13962
rect -758 -14002 -746 -13968
rect -282 -14002 -270 -13968
rect -758 -14008 -270 -14002
rect -550 -14070 -490 -14008
rect -758 -14076 -270 -14070
rect -758 -14110 -746 -14076
rect -282 -14110 -270 -14076
rect -758 -14116 -270 -14110
rect -1050 -14180 -1040 -14160
rect -2024 -14722 -2018 -14184
rect -1046 -14718 -1040 -14180
rect -2024 -14736 -2006 -14722
rect -2794 -14786 -2306 -14780
rect -2794 -14820 -2782 -14786
rect -2318 -14820 -2306 -14786
rect -2794 -14826 -2306 -14820
rect -2588 -14888 -2528 -14826
rect -2794 -14894 -2306 -14888
rect -2794 -14928 -2782 -14894
rect -2318 -14928 -2306 -14894
rect -2794 -14934 -2306 -14928
rect -3086 -15012 -3076 -14978
rect -4060 -15534 -4054 -15012
rect -3082 -15534 -3076 -15012
rect -4060 -15554 -4048 -15534
rect -4830 -15604 -4342 -15598
rect -4830 -15638 -4818 -15604
rect -4354 -15638 -4342 -15604
rect -4830 -15644 -4342 -15638
rect -4628 -15706 -4568 -15644
rect -4830 -15712 -4342 -15706
rect -4830 -15746 -4818 -15712
rect -4354 -15746 -4342 -15712
rect -4830 -15752 -4342 -15746
rect -5120 -15816 -5112 -15796
rect -6096 -16354 -6090 -15824
rect -5118 -16346 -5112 -15816
rect -6096 -16372 -6080 -16354
rect -6866 -16422 -6378 -16416
rect -6866 -16456 -6854 -16422
rect -6390 -16456 -6378 -16422
rect -6866 -16462 -6378 -16456
rect -6658 -16524 -6598 -16462
rect -6866 -16530 -6378 -16524
rect -6866 -16564 -6854 -16530
rect -6390 -16564 -6378 -16530
rect -6866 -16570 -6378 -16564
rect -7158 -16640 -7148 -16614
rect -8132 -17164 -8126 -16642
rect -7154 -17162 -7148 -16640
rect -8132 -17190 -8118 -17164
rect -8902 -17240 -8414 -17234
rect -8902 -17274 -8890 -17240
rect -8426 -17274 -8414 -17240
rect -8902 -17280 -8414 -17274
rect -8690 -17342 -8630 -17280
rect -8902 -17348 -8414 -17342
rect -8902 -17382 -8890 -17348
rect -8426 -17382 -8414 -17348
rect -8902 -17388 -8414 -17382
rect -9198 -17458 -9184 -17432
rect -9190 -17986 -9184 -17458
rect -9198 -18008 -9184 -17986
rect -9150 -17458 -9138 -17432
rect -8178 -17432 -8118 -17190
rect -7158 -17190 -7148 -17162
rect -7114 -16640 -7098 -16614
rect -6140 -16614 -6080 -16372
rect -5120 -16372 -5112 -16346
rect -5078 -15816 -5060 -15796
rect -4108 -15796 -4048 -15554
rect -3086 -15554 -3076 -15534
rect -3042 -15012 -3026 -14978
rect -2066 -14978 -2006 -14736
rect -1050 -14736 -1040 -14718
rect -1006 -14180 -990 -14160
rect -28 -14160 32 -13918
rect -1006 -14718 -1000 -14180
rect -1006 -14736 -990 -14718
rect -1776 -14786 -1288 -14780
rect -1776 -14820 -1764 -14786
rect -1300 -14820 -1288 -14786
rect -1776 -14826 -1288 -14820
rect -1576 -14888 -1516 -14826
rect -1776 -14894 -1288 -14888
rect -1776 -14928 -1764 -14894
rect -1300 -14928 -1288 -14894
rect -1776 -14934 -1288 -14928
rect -2066 -15012 -2058 -14978
rect -3042 -15534 -3036 -15012
rect -2064 -15534 -2058 -15012
rect -3042 -15554 -3026 -15534
rect -3812 -15604 -3324 -15598
rect -3812 -15638 -3800 -15604
rect -3336 -15638 -3324 -15604
rect -3812 -15644 -3324 -15638
rect -3612 -15706 -3552 -15644
rect -3812 -15712 -3324 -15706
rect -3812 -15746 -3800 -15712
rect -3336 -15746 -3324 -15712
rect -3812 -15752 -3324 -15746
rect -5078 -16346 -5072 -15816
rect -4108 -15824 -4094 -15796
rect -5078 -16372 -5060 -16346
rect -4100 -16354 -4094 -15824
rect -5848 -16422 -5360 -16416
rect -5848 -16456 -5836 -16422
rect -5372 -16456 -5360 -16422
rect -5848 -16462 -5360 -16456
rect -5656 -16524 -5596 -16462
rect -5848 -16530 -5360 -16524
rect -5848 -16564 -5836 -16530
rect -5372 -16564 -5360 -16530
rect -5848 -16570 -5360 -16564
rect -7114 -17162 -7108 -16640
rect -6140 -16644 -6130 -16614
rect -7114 -17190 -7098 -17162
rect -6136 -17166 -6130 -16644
rect -7884 -17240 -7396 -17234
rect -7884 -17274 -7872 -17240
rect -7408 -17274 -7396 -17240
rect -7884 -17280 -7396 -17274
rect -7676 -17342 -7616 -17280
rect -7884 -17348 -7396 -17342
rect -7884 -17382 -7872 -17348
rect -7408 -17382 -7396 -17348
rect -7884 -17388 -7396 -17382
rect -8178 -17454 -8166 -17432
rect -9150 -17986 -9144 -17458
rect -8172 -17982 -8166 -17454
rect -9150 -18008 -9138 -17986
rect -9198 -18250 -9138 -18008
rect -8178 -18008 -8166 -17982
rect -8132 -17454 -8118 -17432
rect -7158 -17432 -7098 -17190
rect -6140 -17190 -6130 -17166
rect -6096 -16644 -6080 -16614
rect -5120 -16614 -5060 -16372
rect -4108 -16372 -4094 -16354
rect -4060 -15824 -4048 -15796
rect -3086 -15796 -3026 -15554
rect -2066 -15554 -2058 -15534
rect -2024 -15012 -2006 -14978
rect -1050 -14978 -990 -14736
rect -28 -14736 -22 -14160
rect 12 -14184 32 -14160
rect 12 -14722 18 -14184
rect 12 -14736 32 -14722
rect -758 -14786 -270 -14780
rect -758 -14820 -746 -14786
rect -282 -14820 -270 -14786
rect -758 -14826 -270 -14820
rect -556 -14888 -496 -14826
rect -758 -14894 -270 -14888
rect -758 -14928 -746 -14894
rect -282 -14928 -270 -14894
rect -758 -14934 -270 -14928
rect -1050 -15008 -1040 -14978
rect -2024 -15534 -2018 -15012
rect -1046 -15530 -1040 -15008
rect -2024 -15554 -2006 -15534
rect -2794 -15604 -2306 -15598
rect -2794 -15638 -2782 -15604
rect -2318 -15638 -2306 -15604
rect -2794 -15644 -2306 -15638
rect -2590 -15706 -2530 -15644
rect -2794 -15712 -2306 -15706
rect -2794 -15746 -2782 -15712
rect -2318 -15746 -2306 -15712
rect -2794 -15752 -2306 -15746
rect -3086 -15824 -3076 -15796
rect -4060 -16354 -4054 -15824
rect -3082 -16354 -3076 -15824
rect -4060 -16372 -4048 -16354
rect -4830 -16422 -4342 -16416
rect -4830 -16456 -4818 -16422
rect -4354 -16456 -4342 -16422
rect -4830 -16462 -4342 -16456
rect -4626 -16524 -4566 -16462
rect -4830 -16530 -4342 -16524
rect -4830 -16564 -4818 -16530
rect -4354 -16564 -4342 -16530
rect -4830 -16570 -4342 -16564
rect -5120 -16636 -5112 -16614
rect -6096 -17166 -6090 -16644
rect -5118 -17158 -5112 -16636
rect -6096 -17190 -6080 -17166
rect -6866 -17240 -6378 -17234
rect -6866 -17274 -6854 -17240
rect -6390 -17274 -6378 -17240
rect -6866 -17280 -6378 -17274
rect -6656 -17342 -6596 -17280
rect -6866 -17348 -6378 -17342
rect -6866 -17382 -6854 -17348
rect -6390 -17382 -6378 -17348
rect -6866 -17388 -6378 -17382
rect -7158 -17452 -7148 -17432
rect -8132 -17982 -8126 -17454
rect -7154 -17980 -7148 -17452
rect -8132 -18008 -8118 -17982
rect -8902 -18058 -8414 -18052
rect -8902 -18092 -8890 -18058
rect -8426 -18092 -8414 -18058
rect -8902 -18098 -8414 -18092
rect -8688 -18160 -8628 -18098
rect -8902 -18166 -8414 -18160
rect -8902 -18200 -8890 -18166
rect -8426 -18200 -8414 -18166
rect -8902 -18206 -8414 -18200
rect -9198 -18276 -9184 -18250
rect -9190 -18826 -9184 -18276
rect -9150 -18276 -9138 -18250
rect -8178 -18250 -8118 -18008
rect -7158 -18008 -7148 -17980
rect -7114 -17452 -7098 -17432
rect -6140 -17432 -6080 -17190
rect -5120 -17190 -5112 -17158
rect -5078 -16636 -5060 -16614
rect -4108 -16614 -4048 -16372
rect -3086 -16372 -3076 -16354
rect -3042 -15824 -3026 -15796
rect -2066 -15796 -2006 -15554
rect -1050 -15554 -1040 -15530
rect -1006 -15008 -990 -14978
rect -28 -14978 32 -14736
rect 1850 -14902 1910 -12508
rect 2110 -13782 2170 -11408
rect 2110 -13788 2172 -13782
rect 2110 -13848 2112 -13788
rect 2110 -13854 2172 -13848
rect 1970 -14060 1976 -14000
rect 2036 -14060 2042 -14000
rect 1844 -14962 1850 -14902
rect 1910 -14962 1916 -14902
rect -1006 -15530 -1000 -15008
rect -1006 -15554 -990 -15530
rect -1776 -15604 -1288 -15598
rect -1776 -15638 -1764 -15604
rect -1300 -15638 -1288 -15604
rect -1776 -15644 -1288 -15638
rect -1578 -15706 -1518 -15644
rect -1776 -15712 -1288 -15706
rect -1776 -15746 -1764 -15712
rect -1300 -15746 -1288 -15712
rect -1776 -15752 -1288 -15746
rect -2066 -15824 -2058 -15796
rect -3042 -16354 -3036 -15824
rect -2064 -16354 -2058 -15824
rect -3042 -16372 -3026 -16354
rect -3812 -16422 -3324 -16416
rect -3812 -16456 -3800 -16422
rect -3336 -16456 -3324 -16422
rect -3812 -16462 -3324 -16456
rect -3610 -16524 -3550 -16462
rect -3812 -16530 -3324 -16524
rect -3812 -16564 -3800 -16530
rect -3336 -16564 -3324 -16530
rect -3812 -16570 -3324 -16564
rect -5078 -17158 -5072 -16636
rect -4108 -16644 -4094 -16614
rect -5078 -17190 -5060 -17158
rect -4100 -17166 -4094 -16644
rect -5848 -17240 -5360 -17234
rect -5848 -17274 -5836 -17240
rect -5372 -17274 -5360 -17240
rect -5848 -17280 -5360 -17274
rect -5654 -17342 -5594 -17280
rect -5848 -17348 -5360 -17342
rect -5848 -17382 -5836 -17348
rect -5372 -17382 -5360 -17348
rect -5848 -17388 -5360 -17382
rect -7114 -17980 -7108 -17452
rect -6140 -17456 -6130 -17432
rect -7114 -18008 -7098 -17980
rect -6136 -17984 -6130 -17456
rect -7884 -18058 -7396 -18052
rect -7884 -18092 -7872 -18058
rect -7408 -18092 -7396 -18058
rect -7884 -18098 -7396 -18092
rect -7674 -18160 -7614 -18098
rect -7884 -18166 -7396 -18160
rect -7884 -18200 -7872 -18166
rect -7408 -18200 -7396 -18166
rect -7884 -18206 -7396 -18200
rect -8178 -18272 -8166 -18250
rect -9150 -18826 -9144 -18276
rect -9190 -18838 -9144 -18826
rect -8172 -18826 -8166 -18272
rect -8132 -18272 -8118 -18250
rect -7158 -18250 -7098 -18008
rect -6140 -18008 -6130 -17984
rect -6096 -17456 -6080 -17432
rect -5120 -17432 -5060 -17190
rect -4108 -17190 -4094 -17166
rect -4060 -16644 -4048 -16614
rect -3086 -16614 -3026 -16372
rect -2066 -16372 -2058 -16354
rect -2024 -15824 -2006 -15796
rect -1050 -15796 -990 -15554
rect -28 -15554 -22 -14978
rect 12 -15012 32 -14978
rect 12 -15534 18 -15012
rect 12 -15554 32 -15534
rect -758 -15604 -270 -15598
rect -758 -15638 -746 -15604
rect -282 -15638 -270 -15604
rect -758 -15644 -270 -15638
rect -558 -15706 -498 -15644
rect -758 -15712 -270 -15706
rect -758 -15746 -746 -15712
rect -282 -15746 -270 -15712
rect -758 -15752 -270 -15746
rect -1050 -15820 -1040 -15796
rect -2024 -16354 -2018 -15824
rect -1046 -16350 -1040 -15820
rect -2024 -16372 -2006 -16354
rect -2794 -16422 -2306 -16416
rect -2794 -16456 -2782 -16422
rect -2318 -16456 -2306 -16422
rect -2794 -16462 -2306 -16456
rect -2588 -16524 -2528 -16462
rect -2794 -16530 -2306 -16524
rect -2794 -16564 -2782 -16530
rect -2318 -16564 -2306 -16530
rect -2794 -16570 -2306 -16564
rect -3086 -16644 -3076 -16614
rect -4060 -17166 -4054 -16644
rect -3082 -17166 -3076 -16644
rect -4060 -17190 -4048 -17166
rect -4830 -17240 -4342 -17234
rect -4830 -17274 -4818 -17240
rect -4354 -17274 -4342 -17240
rect -4830 -17280 -4342 -17274
rect -4624 -17342 -4564 -17280
rect -4830 -17348 -4342 -17342
rect -4830 -17382 -4818 -17348
rect -4354 -17382 -4342 -17348
rect -4830 -17388 -4342 -17382
rect -5120 -17448 -5112 -17432
rect -6096 -17984 -6090 -17456
rect -5118 -17976 -5112 -17448
rect -6096 -18008 -6080 -17984
rect -6866 -18058 -6378 -18052
rect -6866 -18092 -6854 -18058
rect -6390 -18092 -6378 -18058
rect -6866 -18098 -6378 -18092
rect -6654 -18160 -6594 -18098
rect -6866 -18166 -6378 -18160
rect -6866 -18200 -6854 -18166
rect -6390 -18200 -6378 -18166
rect -6866 -18206 -6378 -18200
rect -7158 -18270 -7148 -18250
rect -8132 -18826 -8126 -18272
rect -7154 -18780 -7148 -18270
rect -8172 -18838 -8126 -18826
rect -7164 -18826 -7148 -18780
rect -7114 -18270 -7098 -18250
rect -6140 -18250 -6080 -18008
rect -5120 -18008 -5112 -17976
rect -5078 -17448 -5060 -17432
rect -4108 -17432 -4048 -17190
rect -3086 -17190 -3076 -17166
rect -3042 -16644 -3026 -16614
rect -2066 -16614 -2006 -16372
rect -1050 -16372 -1040 -16350
rect -1006 -15820 -990 -15796
rect -28 -15796 32 -15554
rect -1006 -16350 -1000 -15820
rect -1006 -16372 -990 -16350
rect -1776 -16422 -1288 -16416
rect -1776 -16456 -1764 -16422
rect -1300 -16456 -1288 -16422
rect -1776 -16462 -1288 -16456
rect -1576 -16524 -1516 -16462
rect -1776 -16530 -1288 -16524
rect -1776 -16564 -1764 -16530
rect -1300 -16564 -1288 -16530
rect -1776 -16570 -1288 -16564
rect -2066 -16644 -2058 -16614
rect -3042 -17166 -3036 -16644
rect -2064 -17166 -2058 -16644
rect -3042 -17190 -3026 -17166
rect -3812 -17240 -3324 -17234
rect -3812 -17274 -3800 -17240
rect -3336 -17274 -3324 -17240
rect -3812 -17280 -3324 -17274
rect -3608 -17342 -3548 -17280
rect -3812 -17348 -3324 -17342
rect -3812 -17382 -3800 -17348
rect -3336 -17382 -3324 -17348
rect -3812 -17388 -3324 -17382
rect -5078 -17976 -5072 -17448
rect -4108 -17456 -4094 -17432
rect -5078 -18008 -5060 -17976
rect -4100 -17984 -4094 -17456
rect -5848 -18058 -5360 -18052
rect -5848 -18092 -5836 -18058
rect -5372 -18092 -5360 -18058
rect -5848 -18098 -5360 -18092
rect -5652 -18160 -5592 -18098
rect -5848 -18166 -5360 -18160
rect -5848 -18200 -5836 -18166
rect -5372 -18200 -5360 -18166
rect -5848 -18206 -5360 -18200
rect -7114 -18780 -7108 -18270
rect -6140 -18274 -6130 -18250
rect -7114 -18826 -7104 -18780
rect -8902 -18876 -8414 -18870
rect -8902 -18910 -8890 -18876
rect -8426 -18910 -8414 -18876
rect -8902 -18916 -8414 -18910
rect -7884 -18876 -7396 -18870
rect -7884 -18910 -7872 -18876
rect -7408 -18910 -7396 -18876
rect -7884 -18916 -7672 -18910
rect -7612 -18916 -7396 -18910
rect -7164 -19000 -7104 -18826
rect -6136 -18826 -6130 -18274
rect -6096 -18274 -6080 -18250
rect -5120 -18250 -5060 -18008
rect -4108 -18008 -4094 -17984
rect -4060 -17456 -4048 -17432
rect -3086 -17432 -3026 -17190
rect -2066 -17190 -2058 -17166
rect -2024 -16644 -2006 -16614
rect -1050 -16614 -990 -16372
rect -28 -16372 -22 -15796
rect 12 -15824 32 -15796
rect 12 -16354 18 -15824
rect 12 -16372 32 -16354
rect -758 -16422 -270 -16416
rect -758 -16456 -746 -16422
rect -282 -16456 -270 -16422
rect -758 -16462 -270 -16456
rect -556 -16524 -496 -16462
rect -758 -16530 -270 -16524
rect -758 -16564 -746 -16530
rect -282 -16564 -270 -16530
rect -758 -16570 -270 -16564
rect -1050 -16640 -1040 -16614
rect -2024 -17166 -2018 -16644
rect -1046 -17162 -1040 -16640
rect -2024 -17190 -2006 -17166
rect -2794 -17240 -2306 -17234
rect -2794 -17274 -2782 -17240
rect -2318 -17274 -2306 -17240
rect -2794 -17280 -2306 -17274
rect -2586 -17342 -2526 -17280
rect -2794 -17348 -2306 -17342
rect -2794 -17382 -2782 -17348
rect -2318 -17382 -2306 -17348
rect -2794 -17388 -2306 -17382
rect -3086 -17456 -3076 -17432
rect -4060 -17984 -4054 -17456
rect -3082 -17984 -3076 -17456
rect -4060 -18008 -4048 -17984
rect -4830 -18058 -4342 -18052
rect -4830 -18092 -4818 -18058
rect -4354 -18092 -4342 -18058
rect -4830 -18098 -4342 -18092
rect -4622 -18160 -4562 -18098
rect -4830 -18166 -4342 -18160
rect -4830 -18200 -4818 -18166
rect -4354 -18200 -4342 -18166
rect -4830 -18206 -4342 -18200
rect -5120 -18266 -5112 -18250
rect -6096 -18826 -6090 -18274
rect -5118 -18778 -5112 -18266
rect -6136 -18838 -6090 -18826
rect -5126 -18826 -5112 -18778
rect -5078 -18266 -5060 -18250
rect -4108 -18250 -4048 -18008
rect -3086 -18008 -3076 -17984
rect -3042 -17456 -3026 -17432
rect -2066 -17432 -2006 -17190
rect -1050 -17190 -1040 -17162
rect -1006 -16640 -990 -16614
rect -28 -16614 32 -16372
rect -1006 -17162 -1000 -16640
rect -1006 -17190 -990 -17162
rect -1776 -17240 -1288 -17234
rect -1776 -17274 -1764 -17240
rect -1300 -17274 -1288 -17240
rect -1776 -17280 -1288 -17274
rect -1574 -17342 -1514 -17280
rect -1776 -17348 -1288 -17342
rect -1776 -17382 -1764 -17348
rect -1300 -17382 -1288 -17348
rect -1776 -17388 -1288 -17382
rect -2066 -17456 -2058 -17432
rect -3042 -17984 -3036 -17456
rect -2064 -17984 -2058 -17456
rect -3042 -18008 -3026 -17984
rect -3812 -18058 -3324 -18052
rect -3812 -18092 -3800 -18058
rect -3336 -18092 -3324 -18058
rect -3812 -18098 -3324 -18092
rect -3606 -18160 -3546 -18098
rect -3812 -18166 -3324 -18160
rect -3812 -18200 -3800 -18166
rect -3336 -18200 -3324 -18166
rect -3812 -18206 -3324 -18200
rect -5078 -18778 -5072 -18266
rect -4108 -18274 -4094 -18250
rect -5078 -18826 -5066 -18778
rect -6866 -18876 -6378 -18870
rect -6866 -18910 -6854 -18876
rect -6390 -18910 -6378 -18876
rect -6866 -18916 -6378 -18910
rect -5848 -18876 -5360 -18870
rect -5848 -18910 -5836 -18876
rect -5372 -18910 -5360 -18876
rect -5848 -18916 -5360 -18910
rect -5126 -19000 -5066 -18826
rect -4100 -18826 -4094 -18274
rect -4060 -18274 -4048 -18250
rect -3086 -18250 -3026 -18008
rect -2066 -18008 -2058 -17984
rect -2024 -17456 -2006 -17432
rect -1050 -17432 -990 -17190
rect -28 -17190 -22 -16614
rect 12 -16644 32 -16614
rect 12 -17166 18 -16644
rect 12 -17190 32 -17166
rect -758 -17240 -270 -17234
rect -758 -17274 -746 -17240
rect -282 -17274 -270 -17240
rect -758 -17280 -270 -17274
rect -554 -17342 -494 -17280
rect -758 -17348 -270 -17342
rect -758 -17382 -746 -17348
rect -282 -17382 -270 -17348
rect -758 -17388 -270 -17382
rect -1050 -17452 -1040 -17432
rect -2024 -17984 -2018 -17456
rect -1046 -17980 -1040 -17452
rect -2024 -18008 -2006 -17984
rect -2794 -18058 -2306 -18052
rect -2794 -18092 -2782 -18058
rect -2318 -18092 -2306 -18058
rect -2794 -18098 -2306 -18092
rect -2584 -18160 -2524 -18098
rect -2794 -18166 -2306 -18160
rect -2794 -18200 -2782 -18166
rect -2318 -18200 -2306 -18166
rect -2794 -18206 -2306 -18200
rect -3086 -18274 -3076 -18250
rect -4060 -18826 -4054 -18274
rect -3082 -18782 -3076 -18274
rect -4100 -18838 -4054 -18826
rect -3090 -18826 -3076 -18782
rect -3042 -18274 -3026 -18250
rect -2066 -18250 -2006 -18008
rect -1050 -18008 -1040 -17980
rect -1006 -17452 -990 -17432
rect -28 -17432 32 -17190
rect -1006 -17980 -1000 -17452
rect -1006 -18008 -990 -17980
rect -1776 -18058 -1288 -18052
rect -1776 -18092 -1764 -18058
rect -1300 -18092 -1288 -18058
rect -1776 -18098 -1288 -18092
rect -1572 -18160 -1512 -18098
rect -1776 -18166 -1288 -18160
rect -1776 -18200 -1764 -18166
rect -1300 -18200 -1288 -18166
rect -1776 -18206 -1288 -18200
rect -2066 -18274 -2058 -18250
rect -3042 -18782 -3036 -18274
rect -3042 -18826 -3030 -18782
rect -4830 -18876 -4342 -18870
rect -4830 -18910 -4818 -18876
rect -4354 -18910 -4342 -18876
rect -4830 -18916 -4342 -18910
rect -3812 -18876 -3324 -18870
rect -3812 -18910 -3800 -18876
rect -3336 -18910 -3324 -18876
rect -3812 -18916 -3324 -18910
rect -3090 -19000 -3030 -18826
rect -2064 -18826 -2058 -18274
rect -2024 -18274 -2006 -18250
rect -1050 -18250 -990 -18008
rect -28 -18008 -22 -17432
rect 12 -17456 32 -17432
rect 12 -17984 18 -17456
rect 12 -18008 32 -17984
rect -758 -18058 -270 -18052
rect -758 -18092 -746 -18058
rect -282 -18092 -270 -18058
rect -758 -18098 -270 -18092
rect -552 -18160 -492 -18098
rect -758 -18166 -270 -18160
rect -758 -18200 -746 -18166
rect -282 -18200 -270 -18166
rect -758 -18206 -270 -18200
rect -1050 -18270 -1040 -18250
rect -2024 -18826 -2018 -18274
rect -1046 -18784 -1040 -18270
rect -2064 -18838 -2018 -18826
rect -1054 -18826 -1040 -18784
rect -1006 -18270 -990 -18250
rect -28 -18250 32 -18008
rect -1006 -18784 -1000 -18270
rect -28 -18772 -22 -18250
rect -1006 -18826 -994 -18784
rect -2794 -18876 -2306 -18870
rect -2794 -18910 -2782 -18876
rect -2318 -18910 -2306 -18876
rect -2794 -18916 -2306 -18910
rect -1776 -18876 -1288 -18870
rect -1776 -18910 -1764 -18876
rect -1300 -18910 -1288 -18876
rect -1776 -18916 -1288 -18910
rect -1054 -19000 -994 -18826
rect -34 -18826 -22 -18772
rect 12 -18274 32 -18250
rect 12 -18772 18 -18274
rect 12 -18826 26 -18772
rect -758 -18876 -270 -18870
rect -758 -18910 -746 -18876
rect -282 -18910 -270 -18876
rect -758 -18916 -270 -18910
rect -540 -19000 -480 -18916
rect -34 -19000 26 -18826
rect 952 -18858 1012 -18852
rect -7164 -19060 26 -19000
rect 690 -18888 750 -18866
rect -2982 -20220 -2976 -20160
rect -2916 -20220 -2910 -20160
rect -9416 -21614 -8338 -21554
rect -9416 -21793 -9356 -21614
rect -8902 -21703 -8842 -21614
rect -9123 -21709 -8635 -21703
rect -9123 -21743 -9111 -21709
rect -8647 -21743 -8635 -21709
rect -9123 -21749 -8635 -21743
rect -9416 -21838 -9405 -21793
rect -9411 -22369 -9405 -21838
rect -9371 -21838 -9356 -21793
rect -8398 -21793 -8338 -21614
rect -7392 -21660 -7386 -21600
rect -7326 -21660 -7320 -21600
rect -6878 -21614 -5796 -21554
rect -2976 -21556 -2916 -20220
rect -8105 -21709 -7617 -21703
rect -8105 -21743 -8093 -21709
rect -7629 -21743 -7617 -21709
rect -8105 -21749 -7617 -21743
rect -9371 -22369 -9365 -21838
rect -8398 -21842 -8387 -21793
rect -8393 -22324 -8387 -21842
rect -9411 -22381 -9365 -22369
rect -8400 -22369 -8387 -22324
rect -8353 -21842 -8338 -21793
rect -7386 -21793 -7326 -21660
rect -6878 -21703 -6818 -21614
rect -7087 -21709 -6599 -21703
rect -7087 -21743 -7075 -21709
rect -6611 -21743 -6599 -21709
rect -7087 -21749 -6599 -21743
rect -8353 -22324 -8347 -21842
rect -8353 -22369 -8340 -22324
rect -9123 -22419 -8635 -22413
rect -9123 -22453 -9111 -22419
rect -8647 -22453 -8635 -22419
rect -9123 -22459 -8635 -22453
rect -8400 -22504 -8340 -22369
rect -7386 -22369 -7369 -21793
rect -7335 -22369 -7326 -21793
rect -6362 -21793 -6302 -21614
rect -5856 -21703 -5796 -21614
rect -5352 -21660 -5346 -21600
rect -5286 -21660 -5280 -21600
rect -4326 -21616 -2916 -21556
rect -6069 -21709 -5581 -21703
rect -6069 -21743 -6057 -21709
rect -5593 -21743 -5581 -21709
rect -6069 -21749 -5581 -21743
rect -6362 -21850 -6351 -21793
rect -6357 -22328 -6351 -21850
rect -8105 -22419 -7617 -22413
rect -8105 -22453 -8093 -22419
rect -7629 -22453 -7617 -22419
rect -8105 -22459 -7617 -22453
rect -9544 -22564 -9538 -22504
rect -9478 -22564 -9472 -22504
rect -8406 -22564 -8400 -22504
rect -8340 -22564 -8334 -22504
rect -9538 -24926 -9478 -22564
rect -9418 -22780 -8342 -22720
rect -9418 -22906 -9358 -22780
rect -8908 -22816 -8848 -22780
rect -9124 -22822 -8636 -22816
rect -9124 -22856 -9112 -22822
rect -8648 -22856 -8636 -22822
rect -9124 -22862 -8636 -22856
rect -9418 -22966 -9406 -22906
rect -9412 -23482 -9406 -22966
rect -9372 -22966 -9358 -22906
rect -8402 -22906 -8342 -22780
rect -7890 -22816 -7830 -22459
rect -7386 -22600 -7326 -22369
rect -6364 -22369 -6351 -22328
rect -6317 -21850 -6302 -21793
rect -5346 -21793 -5286 -21660
rect -5051 -21709 -4563 -21703
rect -5051 -21743 -5039 -21709
rect -4575 -21743 -4563 -21709
rect -5051 -21749 -4563 -21743
rect -5346 -21838 -5333 -21793
rect -6317 -22328 -6311 -21850
rect -6317 -22369 -6304 -22328
rect -5339 -22330 -5333 -21838
rect -7087 -22419 -6599 -22413
rect -7087 -22453 -7075 -22419
rect -6611 -22453 -6599 -22419
rect -7087 -22459 -6599 -22453
rect -7392 -22660 -7386 -22600
rect -7326 -22660 -7320 -22600
rect -8106 -22822 -7618 -22816
rect -8106 -22856 -8094 -22822
rect -7630 -22856 -7618 -22822
rect -8106 -22862 -7618 -22856
rect -8402 -22952 -8388 -22906
rect -9372 -23482 -9366 -22966
rect -8394 -23436 -8388 -22952
rect -9412 -23494 -9366 -23482
rect -8402 -23482 -8388 -23436
rect -8354 -22952 -8342 -22906
rect -7386 -22906 -7326 -22660
rect -6870 -22816 -6810 -22459
rect -6364 -22716 -6304 -22369
rect -5346 -22369 -5333 -22330
rect -5299 -21838 -5286 -21793
rect -4326 -21793 -4266 -21616
rect -3818 -21703 -3758 -21616
rect -4033 -21709 -3545 -21703
rect -4033 -21743 -4021 -21709
rect -3557 -21743 -3545 -21709
rect -4033 -21749 -3545 -21743
rect -5299 -22330 -5293 -21838
rect -4326 -21846 -4315 -21793
rect -4321 -22324 -4315 -21846
rect -5299 -22369 -5286 -22330
rect -6069 -22419 -5581 -22413
rect -6069 -22453 -6057 -22419
rect -5593 -22453 -5581 -22419
rect -6069 -22459 -5581 -22453
rect -6370 -22776 -6364 -22716
rect -6304 -22776 -6298 -22716
rect -5862 -22816 -5802 -22459
rect -5346 -22600 -5286 -22369
rect -4326 -22369 -4315 -22324
rect -4281 -21846 -4266 -21793
rect -3310 -21793 -3250 -21616
rect -3310 -21840 -3297 -21793
rect -4281 -22324 -4275 -21846
rect -4281 -22369 -4266 -22324
rect -5051 -22419 -4563 -22413
rect -5051 -22453 -5039 -22419
rect -4575 -22453 -4563 -22419
rect -5051 -22459 -4563 -22453
rect -5352 -22660 -5346 -22600
rect -5286 -22660 -5280 -22600
rect -7088 -22822 -6600 -22816
rect -7088 -22856 -7076 -22822
rect -6612 -22856 -6600 -22822
rect -7088 -22862 -6600 -22856
rect -6070 -22822 -5582 -22816
rect -6070 -22856 -6058 -22822
rect -5594 -22856 -5582 -22822
rect -6070 -22862 -5582 -22856
rect -7386 -22952 -7370 -22906
rect -8354 -23436 -8348 -22952
rect -8354 -23482 -8342 -23436
rect -7376 -23440 -7370 -22952
rect -9124 -23532 -8636 -23526
rect -9124 -23566 -9112 -23532
rect -8648 -23566 -8636 -23532
rect -9124 -23572 -8636 -23566
rect -8402 -23724 -8342 -23482
rect -7384 -23482 -7370 -23440
rect -7336 -22952 -7326 -22906
rect -6358 -22906 -6312 -22894
rect -7336 -23440 -7330 -22952
rect -6358 -23430 -6352 -22906
rect -7336 -23482 -7324 -23440
rect -8106 -23532 -7618 -23526
rect -8106 -23566 -8094 -23532
rect -7630 -23566 -7618 -23532
rect -8106 -23572 -7618 -23566
rect -8260 -23676 -8254 -23616
rect -8194 -23676 -8188 -23616
rect -8408 -23784 -8402 -23724
rect -8342 -23784 -8336 -23724
rect -8254 -23826 -8194 -23676
rect -9418 -23886 -8194 -23826
rect -9418 -24017 -9358 -23886
rect -8902 -23927 -8842 -23886
rect -9123 -23933 -8635 -23927
rect -9123 -23967 -9111 -23933
rect -8647 -23967 -8635 -23933
rect -9123 -23973 -8635 -23967
rect -9418 -24058 -9405 -24017
rect -9411 -24593 -9405 -24058
rect -9371 -24058 -9358 -24017
rect -8400 -24017 -8340 -23886
rect -7884 -23927 -7824 -23572
rect -7384 -23836 -7324 -23482
rect -6368 -23482 -6352 -23430
rect -6318 -23430 -6312 -22906
rect -5346 -22906 -5286 -22660
rect -4840 -22816 -4780 -22459
rect -4326 -22504 -4266 -22369
rect -3303 -22369 -3297 -21840
rect -3263 -21840 -3250 -21793
rect -3263 -22369 -3257 -21840
rect -3303 -22381 -3257 -22369
rect -4033 -22419 -3545 -22413
rect -4033 -22453 -4021 -22419
rect -3557 -22453 -3545 -22419
rect -4033 -22459 -3545 -22453
rect -4332 -22564 -4326 -22504
rect -4266 -22564 -4260 -22504
rect -2846 -22610 -2786 -19060
rect -820 -19184 -814 -19124
rect -754 -19184 -748 -19124
rect 92 -19184 98 -19124
rect 158 -19184 164 -19124
rect -1690 -19294 -1684 -19234
rect -1624 -19294 -1618 -19234
rect -2604 -19402 -2598 -19342
rect -2538 -19402 -2532 -19342
rect -2598 -20896 -2538 -19402
rect -2474 -19510 -2468 -19450
rect -2408 -19510 -2402 -19450
rect -2468 -20774 -2408 -19510
rect -2242 -19550 -2154 -19544
rect -2242 -19584 -2230 -19550
rect -2166 -19584 -2154 -19550
rect -2242 -19590 -2154 -19584
rect -2024 -19550 -1936 -19544
rect -2024 -19584 -2012 -19550
rect -1948 -19584 -1936 -19550
rect -2024 -19590 -1936 -19584
rect -1806 -19550 -1718 -19544
rect -1806 -19584 -1794 -19550
rect -1730 -19584 -1718 -19550
rect -1806 -19590 -1718 -19584
rect -2330 -19634 -2284 -19622
rect -2330 -19780 -2324 -19634
rect -2338 -19810 -2324 -19780
rect -2290 -19780 -2284 -19634
rect -2112 -19634 -2066 -19622
rect -2290 -19810 -2278 -19780
rect -2112 -19788 -2106 -19634
rect -2338 -19960 -2278 -19810
rect -2118 -19810 -2106 -19788
rect -2072 -19788 -2066 -19634
rect -1894 -19634 -1848 -19622
rect -2072 -19810 -2058 -19788
rect -1894 -19798 -1888 -19634
rect -2242 -19860 -2154 -19854
rect -2242 -19894 -2230 -19860
rect -2166 -19894 -2154 -19860
rect -2242 -19900 -2154 -19894
rect -2230 -19960 -2170 -19900
rect -2118 -19960 -2058 -19810
rect -1902 -19810 -1888 -19798
rect -1854 -19798 -1848 -19634
rect -1684 -19634 -1624 -19294
rect -926 -19402 -920 -19342
rect -860 -19402 -854 -19342
rect -1144 -19510 -1138 -19450
rect -1078 -19510 -1072 -19450
rect -1138 -19544 -1078 -19510
rect -920 -19544 -860 -19402
rect -1588 -19550 -1500 -19544
rect -1588 -19584 -1576 -19550
rect -1512 -19584 -1500 -19550
rect -1588 -19590 -1500 -19584
rect -1370 -19550 -1282 -19544
rect -1370 -19584 -1358 -19550
rect -1294 -19584 -1282 -19550
rect -1370 -19590 -1282 -19584
rect -1152 -19550 -1064 -19544
rect -1152 -19584 -1140 -19550
rect -1076 -19584 -1064 -19550
rect -1152 -19590 -1064 -19584
rect -934 -19550 -846 -19544
rect -934 -19584 -922 -19550
rect -858 -19584 -846 -19550
rect -934 -19590 -846 -19584
rect -1684 -19650 -1670 -19634
rect -1854 -19810 -1842 -19798
rect -2024 -19860 -1936 -19854
rect -2024 -19894 -2012 -19860
rect -1948 -19894 -1936 -19860
rect -2024 -19900 -1936 -19894
rect -2010 -19950 -1950 -19900
rect -2338 -20020 -2058 -19960
rect -2016 -20010 -2010 -19950
rect -1950 -20010 -1944 -19950
rect -2118 -20278 -2058 -20020
rect -1902 -20050 -1842 -19810
rect -1676 -19810 -1670 -19650
rect -1636 -19650 -1624 -19634
rect -1458 -19634 -1412 -19622
rect -1636 -19810 -1630 -19650
rect -1458 -19784 -1452 -19634
rect -1676 -19822 -1630 -19810
rect -1464 -19810 -1452 -19784
rect -1418 -19784 -1412 -19634
rect -1240 -19634 -1194 -19622
rect -1240 -19774 -1234 -19634
rect -1418 -19810 -1404 -19784
rect -1806 -19860 -1718 -19854
rect -1806 -19894 -1794 -19860
rect -1730 -19894 -1718 -19860
rect -1806 -19900 -1718 -19894
rect -1588 -19860 -1500 -19854
rect -1588 -19894 -1576 -19860
rect -1512 -19894 -1500 -19860
rect -1588 -19900 -1500 -19894
rect -1908 -20110 -1902 -20050
rect -1842 -20110 -1836 -20050
rect -1906 -20220 -1900 -20160
rect -1840 -20220 -1834 -20160
rect -2336 -20338 -2058 -20278
rect -2336 -20466 -2276 -20338
rect -2226 -20376 -2166 -20338
rect -2242 -20382 -2154 -20376
rect -2242 -20416 -2230 -20382
rect -2166 -20416 -2154 -20382
rect -2242 -20422 -2154 -20416
rect -2336 -20492 -2324 -20466
rect -2330 -20642 -2324 -20492
rect -2290 -20492 -2276 -20466
rect -2118 -20466 -2058 -20338
rect -2024 -20382 -1936 -20376
rect -2024 -20416 -2012 -20382
rect -1948 -20416 -1936 -20382
rect -2024 -20422 -1936 -20416
rect -2290 -20642 -2284 -20492
rect -2330 -20654 -2284 -20642
rect -2118 -20642 -2106 -20466
rect -2072 -20642 -2058 -20466
rect -1900 -20466 -1840 -20220
rect -1792 -20270 -1732 -19900
rect -1572 -20270 -1512 -19900
rect -1464 -20050 -1404 -19810
rect -1248 -19810 -1234 -19774
rect -1200 -19774 -1194 -19634
rect -1022 -19634 -976 -19622
rect -1200 -19810 -1188 -19774
rect -1022 -19776 -1016 -19634
rect -1370 -19860 -1282 -19854
rect -1370 -19894 -1358 -19860
rect -1294 -19894 -1282 -19860
rect -1370 -19900 -1282 -19894
rect -1354 -19950 -1294 -19900
rect -1360 -20010 -1354 -19950
rect -1294 -20010 -1288 -19950
rect -1470 -20110 -1464 -20050
rect -1404 -20110 -1398 -20050
rect -1472 -20220 -1466 -20160
rect -1406 -20220 -1400 -20160
rect -1798 -20330 -1792 -20270
rect -1732 -20330 -1726 -20270
rect -1578 -20330 -1572 -20270
rect -1512 -20330 -1506 -20270
rect -1792 -20376 -1732 -20330
rect -1572 -20376 -1512 -20330
rect -1806 -20382 -1718 -20376
rect -1806 -20416 -1794 -20382
rect -1730 -20416 -1718 -20382
rect -1806 -20422 -1718 -20416
rect -1588 -20382 -1500 -20376
rect -1588 -20416 -1576 -20382
rect -1512 -20416 -1500 -20382
rect -1588 -20422 -1500 -20416
rect -1900 -20502 -1888 -20466
rect -2242 -20692 -2154 -20686
rect -2242 -20726 -2230 -20692
rect -2166 -20726 -2154 -20692
rect -2242 -20732 -2154 -20726
rect -2474 -20834 -2468 -20774
rect -2408 -20834 -2402 -20774
rect -2604 -20956 -2598 -20896
rect -2538 -20956 -2532 -20896
rect -2118 -21020 -2058 -20642
rect -1894 -20642 -1888 -20502
rect -1854 -20502 -1840 -20466
rect -1676 -20466 -1630 -20454
rect -1854 -20642 -1848 -20502
rect -1676 -20602 -1670 -20466
rect -1894 -20654 -1848 -20642
rect -1680 -20642 -1670 -20602
rect -1636 -20602 -1630 -20466
rect -1466 -20466 -1406 -20220
rect -1370 -20382 -1282 -20376
rect -1370 -20416 -1358 -20382
rect -1294 -20416 -1282 -20382
rect -1370 -20422 -1282 -20416
rect -1466 -20496 -1452 -20466
rect -1636 -20642 -1620 -20602
rect -2024 -20692 -1936 -20686
rect -2024 -20726 -2012 -20692
rect -1948 -20726 -1936 -20692
rect -2024 -20732 -1936 -20726
rect -1806 -20692 -1718 -20686
rect -1806 -20726 -1794 -20692
rect -1730 -20726 -1718 -20692
rect -1806 -20732 -1718 -20726
rect -2010 -20774 -1950 -20732
rect -2016 -20834 -2010 -20774
rect -1950 -20834 -1944 -20774
rect -1792 -20896 -1732 -20732
rect -1798 -20956 -1792 -20896
rect -1732 -20956 -1726 -20896
rect -2124 -21080 -2118 -21020
rect -2058 -21080 -2052 -21020
rect -1680 -21146 -1620 -20642
rect -1458 -20642 -1452 -20496
rect -1418 -20496 -1406 -20466
rect -1248 -20466 -1188 -19810
rect -1028 -19810 -1016 -19776
rect -982 -19776 -976 -19634
rect -814 -19634 -754 -19184
rect -28 -19294 -22 -19234
rect 38 -19294 44 -19234
rect -708 -19402 -702 -19342
rect -642 -19402 -636 -19342
rect -702 -19544 -642 -19402
rect -490 -19510 -484 -19450
rect -424 -19510 -418 -19450
rect -484 -19544 -424 -19510
rect -716 -19550 -628 -19544
rect -716 -19584 -704 -19550
rect -640 -19584 -628 -19550
rect -716 -19590 -628 -19584
rect -498 -19550 -410 -19544
rect -498 -19584 -486 -19550
rect -422 -19584 -410 -19550
rect -498 -19590 -410 -19584
rect -280 -19550 -192 -19544
rect -280 -19584 -268 -19550
rect -204 -19584 -192 -19550
rect -280 -19590 -192 -19584
rect -814 -19680 -798 -19634
rect -982 -19810 -968 -19776
rect -1152 -19860 -1064 -19854
rect -1152 -19894 -1140 -19860
rect -1076 -19894 -1064 -19860
rect -1152 -19900 -1064 -19894
rect -1028 -20050 -968 -19810
rect -804 -19810 -798 -19680
rect -764 -19680 -754 -19634
rect -586 -19634 -540 -19622
rect -764 -19810 -758 -19680
rect -586 -19784 -580 -19634
rect -804 -19822 -758 -19810
rect -592 -19810 -580 -19784
rect -546 -19784 -540 -19634
rect -368 -19634 -322 -19622
rect -546 -19810 -532 -19784
rect -368 -19792 -362 -19634
rect -934 -19860 -846 -19854
rect -934 -19894 -922 -19860
rect -858 -19894 -846 -19860
rect -934 -19900 -846 -19894
rect -716 -19860 -628 -19854
rect -716 -19894 -704 -19860
rect -640 -19894 -628 -19860
rect -716 -19900 -628 -19894
rect -592 -20050 -532 -19810
rect -374 -19810 -362 -19792
rect -328 -19792 -322 -19634
rect -150 -19634 -104 -19622
rect -150 -19774 -144 -19634
rect -328 -19810 -314 -19792
rect -498 -19860 -410 -19854
rect -498 -19894 -486 -19860
rect -422 -19894 -410 -19860
rect -498 -19900 -410 -19894
rect -490 -20010 -484 -19950
rect -424 -20010 -418 -19950
rect -374 -19952 -314 -19810
rect -156 -19810 -144 -19774
rect -110 -19774 -104 -19634
rect -22 -19724 38 -19294
rect -110 -19810 -96 -19774
rect -280 -19860 -192 -19854
rect -280 -19894 -268 -19860
rect -204 -19894 -192 -19860
rect -280 -19900 -192 -19894
rect -266 -19952 -206 -19900
rect -156 -19952 -96 -19810
rect -1138 -20110 -532 -20050
rect -1138 -20160 -1078 -20110
rect -1144 -20220 -1138 -20160
rect -1078 -20220 -1072 -20160
rect -1034 -20220 -1028 -20160
rect -968 -20220 -962 -20160
rect -598 -20220 -592 -20160
rect -532 -20220 -526 -20160
rect -1152 -20382 -1064 -20376
rect -1152 -20416 -1140 -20382
rect -1076 -20416 -1064 -20382
rect -1152 -20422 -1064 -20416
rect -1418 -20642 -1412 -20496
rect -1458 -20654 -1412 -20642
rect -1248 -20642 -1234 -20466
rect -1200 -20642 -1188 -20466
rect -1028 -20466 -968 -20220
rect -924 -20330 -918 -20270
rect -858 -20330 -852 -20270
rect -708 -20330 -702 -20270
rect -642 -20330 -636 -20270
rect -918 -20376 -858 -20330
rect -702 -20376 -642 -20330
rect -934 -20382 -846 -20376
rect -934 -20416 -922 -20382
rect -858 -20416 -846 -20382
rect -934 -20422 -846 -20416
rect -716 -20382 -628 -20376
rect -716 -20416 -704 -20382
rect -640 -20416 -628 -20382
rect -716 -20422 -628 -20416
rect -1028 -20484 -1016 -20466
rect -1588 -20692 -1500 -20686
rect -1588 -20726 -1576 -20692
rect -1512 -20726 -1500 -20692
rect -1588 -20732 -1500 -20726
rect -1370 -20692 -1282 -20686
rect -1370 -20726 -1358 -20692
rect -1294 -20726 -1282 -20692
rect -1370 -20732 -1282 -20726
rect -1574 -20896 -1514 -20732
rect -1354 -20774 -1294 -20732
rect -1360 -20834 -1354 -20774
rect -1294 -20834 -1288 -20774
rect -1580 -20956 -1574 -20896
rect -1514 -20956 -1508 -20896
rect -1686 -21206 -1680 -21146
rect -1620 -21206 -1614 -21146
rect -1344 -21260 -1296 -20834
rect -1248 -21020 -1188 -20642
rect -1022 -20642 -1016 -20484
rect -982 -20484 -968 -20466
rect -804 -20466 -758 -20454
rect -982 -20642 -976 -20484
rect -804 -20620 -798 -20466
rect -1022 -20654 -976 -20642
rect -810 -20642 -798 -20620
rect -764 -20620 -758 -20466
rect -592 -20466 -532 -20220
rect -484 -20376 -424 -20010
rect -374 -20012 -96 -19952
rect -374 -20070 -314 -20012
rect -380 -20130 -374 -20070
rect -314 -20130 -308 -20070
rect -374 -20268 -314 -20130
rect -374 -20328 -96 -20268
rect -498 -20382 -410 -20376
rect -498 -20416 -486 -20382
rect -422 -20416 -410 -20382
rect -498 -20422 -410 -20416
rect -592 -20498 -580 -20466
rect -764 -20642 -750 -20620
rect -1152 -20692 -1064 -20686
rect -1152 -20726 -1140 -20692
rect -1076 -20726 -1064 -20692
rect -1152 -20732 -1064 -20726
rect -934 -20692 -846 -20686
rect -934 -20726 -922 -20692
rect -858 -20726 -846 -20692
rect -934 -20732 -846 -20726
rect -1138 -20894 -1078 -20732
rect -810 -20774 -750 -20642
rect -586 -20642 -580 -20498
rect -546 -20498 -532 -20466
rect -374 -20466 -314 -20328
rect -266 -20376 -206 -20328
rect -280 -20382 -192 -20376
rect -280 -20416 -268 -20382
rect -204 -20416 -192 -20382
rect -280 -20422 -192 -20416
rect -374 -20484 -362 -20466
rect -546 -20642 -540 -20498
rect -368 -20612 -362 -20484
rect -586 -20654 -540 -20642
rect -376 -20642 -362 -20612
rect -328 -20484 -314 -20466
rect -156 -20466 -96 -20328
rect -328 -20612 -322 -20484
rect -156 -20486 -144 -20466
rect -328 -20642 -316 -20612
rect -716 -20692 -628 -20686
rect -716 -20726 -704 -20692
rect -640 -20726 -628 -20692
rect -716 -20732 -628 -20726
rect -498 -20692 -410 -20686
rect -498 -20726 -486 -20692
rect -422 -20726 -410 -20692
rect -498 -20732 -410 -20726
rect -816 -20834 -810 -20774
rect -750 -20834 -744 -20774
rect -482 -20894 -422 -20732
rect -1144 -20954 -1138 -20894
rect -1078 -20954 -1072 -20894
rect -488 -20954 -482 -20894
rect -422 -20954 -416 -20894
rect -376 -21020 -316 -20642
rect -150 -20642 -144 -20486
rect -110 -20486 -96 -20466
rect -110 -20642 -104 -20486
rect -150 -20654 -104 -20642
rect -280 -20692 -192 -20686
rect -280 -20726 -268 -20692
rect -204 -20726 -192 -20692
rect -280 -20732 -192 -20726
rect -22 -20774 38 -19784
rect -28 -20834 -22 -20774
rect 38 -20834 44 -20774
rect -1254 -21080 -1248 -21020
rect -1188 -21080 -1182 -21020
rect -382 -21080 -376 -21020
rect -316 -21080 -310 -21020
rect 98 -21146 158 -19184
rect 214 -20010 220 -19950
rect 280 -20010 286 -19950
rect 220 -20196 280 -20010
rect 220 -20264 280 -20256
rect 92 -21206 98 -21146
rect 158 -21206 164 -21146
rect -1352 -21312 -1346 -21260
rect -1294 -21312 -1288 -21260
rect 690 -21340 750 -18948
rect -2538 -21400 750 -21340
rect -2676 -21640 -2670 -21580
rect -2610 -21640 -2604 -21580
rect -4328 -22670 -2786 -22610
rect -5052 -22822 -4564 -22816
rect -5052 -22856 -5040 -22822
rect -4576 -22856 -4564 -22822
rect -5052 -22862 -4564 -22856
rect -5346 -22940 -5334 -22906
rect -6318 -23482 -6308 -23430
rect -5340 -23448 -5334 -22940
rect -7088 -23532 -6600 -23526
rect -7088 -23566 -7076 -23532
rect -6612 -23566 -6600 -23532
rect -7088 -23572 -6600 -23566
rect -7390 -23896 -7384 -23836
rect -7324 -23896 -7318 -23836
rect -8105 -23933 -7617 -23927
rect -8105 -23967 -8093 -23933
rect -7629 -23967 -7617 -23933
rect -8105 -23973 -7617 -23967
rect -8400 -24058 -8387 -24017
rect -9371 -24593 -9365 -24058
rect -9411 -24605 -9365 -24593
rect -8393 -24593 -8387 -24058
rect -8353 -24058 -8340 -24017
rect -7384 -24017 -7324 -23896
rect -6870 -23927 -6810 -23572
rect -6368 -23616 -6308 -23482
rect -5344 -23482 -5334 -23448
rect -5300 -22940 -5286 -22906
rect -4328 -22906 -4268 -22670
rect -3818 -22816 -3758 -22670
rect -4034 -22822 -3546 -22816
rect -4034 -22856 -4022 -22822
rect -3558 -22856 -3546 -22822
rect -4034 -22862 -3546 -22856
rect -3312 -22906 -3252 -22670
rect -3208 -22776 -3202 -22716
rect -3142 -22776 -3136 -22716
rect -5300 -23448 -5294 -22940
rect -4328 -22952 -4316 -22906
rect -4326 -22954 -4316 -22952
rect -4322 -23444 -4316 -22954
rect -5300 -23482 -5284 -23448
rect -6070 -23532 -5582 -23526
rect -6070 -23566 -6058 -23532
rect -5594 -23566 -5582 -23532
rect -6070 -23572 -5582 -23566
rect -6374 -23676 -6368 -23616
rect -6308 -23676 -6302 -23616
rect -6372 -23784 -6366 -23724
rect -6306 -23784 -6300 -23724
rect -7087 -23933 -6599 -23927
rect -7087 -23967 -7075 -23933
rect -6611 -23967 -6599 -23933
rect -7087 -23973 -6599 -23967
rect -7384 -24046 -7369 -24017
rect -8353 -24593 -8347 -24058
rect -7375 -24556 -7369 -24046
rect -8393 -24605 -8347 -24593
rect -7382 -24593 -7369 -24556
rect -7335 -24046 -7324 -24017
rect -6366 -24017 -6306 -23784
rect -5842 -23927 -5782 -23572
rect -5344 -23830 -5284 -23482
rect -4330 -23482 -4316 -23444
rect -4282 -22954 -4266 -22906
rect -3312 -22936 -3298 -22906
rect -3310 -22938 -3298 -22936
rect -4282 -23444 -4276 -22954
rect -4282 -23482 -4270 -23444
rect -5052 -23532 -4564 -23526
rect -5052 -23566 -5040 -23532
rect -4576 -23566 -4564 -23532
rect -5052 -23572 -4564 -23566
rect -5346 -23836 -5284 -23830
rect -5286 -23896 -5284 -23836
rect -5346 -23902 -5284 -23896
rect -6069 -23933 -5581 -23927
rect -6069 -23967 -6057 -23933
rect -5593 -23967 -5581 -23933
rect -6069 -23973 -5581 -23967
rect -7335 -24556 -7329 -24046
rect -6366 -24060 -6351 -24017
rect -7335 -24593 -7322 -24556
rect -9123 -24643 -8635 -24637
rect -9123 -24677 -9111 -24643
rect -8647 -24677 -8635 -24643
rect -9123 -24683 -8635 -24677
rect -8105 -24643 -7617 -24637
rect -8105 -24677 -8093 -24643
rect -7629 -24677 -7617 -24643
rect -8105 -24683 -7617 -24677
rect -8406 -24880 -8400 -24820
rect -8340 -24880 -8334 -24820
rect -9544 -24986 -9538 -24926
rect -9478 -24986 -9472 -24926
rect -9124 -25046 -8636 -25040
rect -9124 -25080 -9112 -25046
rect -8648 -25080 -8636 -25046
rect -9124 -25086 -8636 -25080
rect -9412 -25130 -9366 -25118
rect -9412 -25666 -9406 -25130
rect -9418 -25706 -9406 -25666
rect -9372 -25666 -9366 -25130
rect -8400 -25130 -8340 -24880
rect -7876 -25040 -7816 -24683
rect -7382 -24718 -7322 -24593
rect -6357 -24593 -6351 -24060
rect -6317 -24060 -6306 -24017
rect -5344 -24017 -5284 -23902
rect -4832 -23927 -4772 -23572
rect -4504 -23676 -4498 -23616
rect -4438 -23676 -4432 -23616
rect -4498 -23826 -4438 -23676
rect -4330 -23724 -4270 -23482
rect -3304 -23482 -3298 -22938
rect -3264 -22938 -3250 -22906
rect -3264 -23482 -3258 -22938
rect -3304 -23494 -3258 -23482
rect -4034 -23532 -3546 -23526
rect -4034 -23566 -4022 -23532
rect -3558 -23566 -3546 -23532
rect -4034 -23572 -3546 -23566
rect -4336 -23784 -4330 -23724
rect -4270 -23784 -4264 -23724
rect -4498 -23886 -3254 -23826
rect -5051 -23933 -4563 -23927
rect -5051 -23967 -5039 -23933
rect -4575 -23967 -4563 -23933
rect -5051 -23973 -4563 -23967
rect -5344 -24054 -5333 -24017
rect -6317 -24593 -6311 -24060
rect -5339 -24560 -5333 -24054
rect -6357 -24605 -6311 -24593
rect -5348 -24593 -5333 -24560
rect -5299 -24054 -5284 -24017
rect -4328 -24017 -4268 -23886
rect -3810 -23927 -3750 -23886
rect -4033 -23933 -3545 -23927
rect -4033 -23967 -4021 -23933
rect -3557 -23967 -3545 -23933
rect -4033 -23973 -3545 -23967
rect -5299 -24560 -5293 -24054
rect -4328 -24058 -4315 -24017
rect -5299 -24593 -5288 -24560
rect -7087 -24643 -6599 -24637
rect -7087 -24677 -7075 -24643
rect -6611 -24677 -6599 -24643
rect -7087 -24683 -6599 -24677
rect -6069 -24643 -5581 -24637
rect -6069 -24677 -6057 -24643
rect -5593 -24677 -5581 -24643
rect -6069 -24683 -5581 -24677
rect -7388 -24778 -7382 -24718
rect -7322 -24778 -7316 -24718
rect -8106 -25046 -7618 -25040
rect -8106 -25080 -8094 -25046
rect -7630 -25080 -7618 -25046
rect -8106 -25086 -7618 -25080
rect -8400 -25174 -8388 -25130
rect -9372 -25706 -9358 -25666
rect -8394 -25672 -8388 -25174
rect -9418 -25870 -9358 -25706
rect -8402 -25706 -8388 -25672
rect -8354 -25174 -8340 -25130
rect -7382 -25130 -7322 -24778
rect -6876 -25040 -6816 -24683
rect -6372 -24986 -6366 -24926
rect -6306 -24986 -6300 -24926
rect -7088 -25046 -6600 -25040
rect -7088 -25080 -7076 -25046
rect -6612 -25080 -6600 -25046
rect -7088 -25086 -6600 -25080
rect -8354 -25672 -8348 -25174
rect -8354 -25706 -8342 -25672
rect -9124 -25756 -8636 -25750
rect -9124 -25790 -9112 -25756
rect -8648 -25790 -8636 -25756
rect -9124 -25796 -8636 -25790
rect -8910 -25870 -8850 -25796
rect -8402 -25870 -8342 -25706
rect -7382 -25706 -7370 -25130
rect -7336 -25706 -7322 -25130
rect -6366 -25130 -6306 -24986
rect -5852 -25040 -5792 -24683
rect -5348 -24712 -5288 -24593
rect -4321 -24593 -4315 -24058
rect -4281 -24058 -4268 -24017
rect -3314 -24017 -3254 -23886
rect -3314 -24052 -3297 -24017
rect -4281 -24593 -4275 -24058
rect -4321 -24605 -4275 -24593
rect -3303 -24593 -3297 -24052
rect -3263 -24052 -3254 -24017
rect -3263 -24593 -3257 -24052
rect -3303 -24605 -3257 -24593
rect -5051 -24643 -4563 -24637
rect -5051 -24677 -5039 -24643
rect -4575 -24677 -4563 -24643
rect -5051 -24683 -4563 -24677
rect -4033 -24643 -3545 -24637
rect -4033 -24677 -4021 -24643
rect -3557 -24677 -3545 -24643
rect -4033 -24683 -3545 -24677
rect -5352 -24718 -5288 -24712
rect -5292 -24778 -5288 -24718
rect -5352 -24784 -5288 -24778
rect -6070 -25046 -5582 -25040
rect -6070 -25080 -6058 -25046
rect -5594 -25080 -5582 -25046
rect -6070 -25086 -5582 -25080
rect -6366 -25182 -6352 -25130
rect -8106 -25756 -7618 -25750
rect -8106 -25790 -8094 -25756
rect -7630 -25790 -7618 -25756
rect -8106 -25796 -7618 -25790
rect -7896 -25870 -7836 -25796
rect -9418 -25930 -7896 -25870
rect -7836 -25930 -7830 -25870
rect -12328 -27116 -12216 -26330
rect -7382 -26430 -7322 -25706
rect -6358 -25706 -6352 -25182
rect -6318 -25182 -6306 -25130
rect -5348 -25130 -5288 -24784
rect -4836 -25040 -4776 -24683
rect -3202 -24820 -3142 -22776
rect -2670 -23620 -2610 -21640
rect -2538 -22614 -2478 -21400
rect -2122 -21480 -2062 -21474
rect 952 -21480 1012 -18918
rect -2124 -21540 -2122 -21534
rect -938 -21540 -932 -21480
rect -872 -21540 -866 -21480
rect 256 -21540 262 -21480
rect 322 -21540 328 -21480
rect 946 -21540 952 -21480
rect 1012 -21540 1018 -21480
rect -2124 -21575 -2062 -21540
rect -2427 -21637 -2062 -21575
rect -2427 -21792 -2365 -21637
rect -2275 -21702 -2213 -21637
rect -2308 -21708 -2180 -21702
rect -2308 -21742 -2296 -21708
rect -2192 -21742 -2180 -21708
rect -2308 -21748 -2180 -21742
rect -2124 -21792 -2062 -21637
rect -1684 -21640 -1678 -21580
rect -1618 -21640 -1612 -21580
rect -1386 -21640 -1380 -21580
rect -1320 -21640 -1314 -21580
rect -1678 -21702 -1618 -21640
rect -1380 -21702 -1320 -21640
rect -2010 -21708 -1882 -21702
rect -2010 -21742 -1998 -21708
rect -1894 -21742 -1882 -21708
rect -2010 -21748 -1882 -21742
rect -1712 -21708 -1584 -21702
rect -1712 -21742 -1700 -21708
rect -1596 -21742 -1584 -21708
rect -1712 -21748 -1584 -21742
rect -1414 -21708 -1286 -21702
rect -1414 -21742 -1402 -21708
rect -1298 -21742 -1286 -21708
rect -1414 -21748 -1286 -21742
rect -1116 -21708 -988 -21702
rect -1116 -21742 -1104 -21708
rect -1000 -21742 -988 -21708
rect -1116 -21748 -988 -21742
rect -1522 -21792 -1476 -21780
rect -2427 -21825 -2410 -21792
rect -2416 -22368 -2410 -21825
rect -2376 -21824 -2362 -21792
rect -2376 -21825 -2365 -21824
rect -2376 -22368 -2370 -21825
rect -2124 -21832 -2112 -21792
rect -2122 -21844 -2112 -21832
rect -2416 -22380 -2370 -22368
rect -2118 -22368 -2112 -21844
rect -2078 -21844 -2062 -21792
rect -2078 -22368 -2072 -21844
rect -1820 -22319 -1814 -21832
rect -2118 -22380 -2072 -22368
rect -1829 -22368 -1814 -22319
rect -1780 -22319 -1774 -21832
rect -1522 -22312 -1516 -21792
rect -1780 -22368 -1771 -22319
rect -1530 -22332 -1516 -22312
rect -2308 -22418 -2180 -22412
rect -2308 -22452 -2296 -22418
rect -2192 -22452 -2180 -22418
rect -2308 -22458 -2180 -22452
rect -2126 -22614 -2066 -22608
rect -2548 -22674 -2542 -22614
rect -2482 -22674 -2476 -22614
rect -2066 -22674 -2064 -22664
rect -2126 -22704 -2064 -22674
rect -2422 -22764 -2064 -22704
rect -1974 -22722 -1914 -22452
rect -1829 -22483 -1771 -22368
rect -1532 -22368 -1516 -22332
rect -1482 -22312 -1476 -21792
rect -1224 -21792 -1178 -21786
rect -1482 -22368 -1470 -22312
rect -1224 -22354 -1218 -21792
rect -1230 -22368 -1218 -22354
rect -1184 -22354 -1178 -21792
rect -932 -21792 -872 -21540
rect -490 -21640 -484 -21580
rect -424 -21640 -418 -21580
rect -194 -21640 -188 -21580
rect -128 -21640 -122 -21580
rect -484 -21702 -424 -21640
rect -188 -21702 -128 -21640
rect -818 -21708 -690 -21702
rect -818 -21742 -806 -21708
rect -702 -21742 -690 -21708
rect -818 -21748 -690 -21742
rect -520 -21708 -392 -21702
rect -520 -21742 -508 -21708
rect -404 -21742 -392 -21708
rect -520 -21748 -392 -21742
rect -222 -21708 -94 -21702
rect -222 -21742 -210 -21708
rect -106 -21742 -94 -21708
rect -222 -21748 -94 -21742
rect 76 -21708 204 -21702
rect 76 -21742 88 -21708
rect 192 -21742 204 -21708
rect 76 -21748 204 -21742
rect -330 -21792 -284 -21780
rect 262 -21792 322 -21540
rect 374 -21708 502 -21702
rect 374 -21742 386 -21708
rect 490 -21742 502 -21708
rect 374 -21748 502 -21742
rect 672 -21708 800 -21702
rect 672 -21742 684 -21708
rect 788 -21742 800 -21708
rect 672 -21748 800 -21742
rect -932 -21852 -920 -21792
rect -1184 -22361 -1170 -22354
rect -1184 -22368 -1167 -22361
rect -1712 -22418 -1584 -22412
rect -1712 -22452 -1700 -22418
rect -1596 -22452 -1584 -22418
rect -1712 -22458 -1584 -22452
rect -1835 -22541 -1829 -22483
rect -1771 -22541 -1765 -22483
rect -2422 -22904 -2362 -22764
rect -2274 -22814 -2214 -22764
rect -2308 -22820 -2180 -22814
rect -2308 -22854 -2296 -22820
rect -2192 -22854 -2180 -22820
rect -2308 -22860 -2180 -22854
rect -2422 -22952 -2410 -22904
rect -2416 -23480 -2410 -22952
rect -2376 -22952 -2362 -22904
rect -2126 -22904 -2064 -22764
rect -1980 -22782 -1974 -22722
rect -1914 -22782 -1908 -22722
rect -2010 -22820 -1882 -22814
rect -2010 -22854 -1998 -22820
rect -1894 -22854 -1882 -22820
rect -2010 -22860 -1882 -22854
rect -2126 -22942 -2112 -22904
rect -2376 -23480 -2370 -22952
rect -2124 -22954 -2112 -22942
rect -2118 -23440 -2112 -22954
rect -2416 -23492 -2370 -23480
rect -2126 -23480 -2112 -23440
rect -2078 -22954 -2064 -22904
rect -1829 -22904 -1771 -22541
rect -1532 -22614 -1472 -22368
rect -1414 -22418 -1286 -22412
rect -1414 -22452 -1402 -22418
rect -1298 -22452 -1286 -22418
rect -1414 -22458 -1286 -22452
rect -1230 -22483 -1167 -22368
rect -926 -22368 -920 -21852
rect -886 -21852 -872 -21792
rect -886 -22368 -880 -21852
rect -628 -22345 -622 -21878
rect -926 -22380 -880 -22368
rect -634 -22368 -622 -22345
rect -588 -22345 -582 -21878
rect -330 -22310 -324 -21792
rect -338 -22326 -324 -22310
rect -588 -22368 -576 -22345
rect -1116 -22418 -988 -22412
rect -1116 -22452 -1104 -22418
rect -1000 -22452 -988 -22418
rect -1116 -22458 -988 -22452
rect -818 -22418 -690 -22412
rect -818 -22452 -806 -22418
rect -702 -22452 -690 -22418
rect -818 -22458 -690 -22452
rect -1231 -22541 -1225 -22483
rect -1167 -22541 -1161 -22483
rect -1538 -22674 -1532 -22614
rect -1472 -22674 -1466 -22614
rect -1682 -22782 -1676 -22722
rect -1616 -22782 -1610 -22722
rect -1382 -22782 -1376 -22722
rect -1316 -22782 -1310 -22722
rect -1676 -22814 -1616 -22782
rect -1376 -22814 -1316 -22782
rect -1704 -22820 -1584 -22814
rect -1704 -22854 -1700 -22820
rect -1596 -22854 -1584 -22820
rect -1704 -22860 -1584 -22854
rect -1414 -22820 -1286 -22814
rect -1414 -22854 -1402 -22820
rect -1298 -22854 -1286 -22820
rect -1414 -22860 -1286 -22854
rect -1829 -22935 -1814 -22904
rect -2078 -23440 -2072 -22954
rect -1820 -23440 -1814 -23002
rect -2078 -23480 -2066 -23440
rect -2308 -23530 -2180 -23524
rect -2308 -23564 -2296 -23530
rect -2192 -23564 -2180 -23530
rect -2308 -23570 -2180 -23564
rect -2676 -23680 -2670 -23620
rect -2610 -23680 -2604 -23620
rect -4338 -24880 -4332 -24820
rect -4272 -24880 -4266 -24820
rect -3208 -24880 -3202 -24820
rect -3142 -24880 -3136 -24820
rect -5052 -25046 -4564 -25040
rect -5052 -25080 -5040 -25046
rect -4576 -25080 -4564 -25046
rect -5052 -25086 -4564 -25080
rect -6318 -25706 -6312 -25182
rect -6358 -25718 -6312 -25706
rect -5348 -25706 -5334 -25130
rect -5300 -25706 -5288 -25130
rect -4332 -25130 -4272 -24880
rect -4034 -25046 -3546 -25040
rect -4034 -25080 -4022 -25046
rect -3558 -25080 -3546 -25046
rect -4034 -25086 -3546 -25080
rect -4332 -25170 -4316 -25130
rect -4322 -25650 -4316 -25170
rect -7088 -25756 -6600 -25750
rect -7088 -25790 -7076 -25756
rect -6612 -25790 -6600 -25756
rect -7088 -25796 -6600 -25790
rect -6070 -25756 -5582 -25750
rect -6070 -25790 -6058 -25756
rect -5594 -25790 -5582 -25756
rect -6070 -25796 -5582 -25790
rect -6870 -25870 -6810 -25796
rect -5846 -25870 -5786 -25796
rect -6876 -25930 -6870 -25870
rect -6810 -25930 -6804 -25870
rect -5852 -25930 -5846 -25870
rect -5786 -25930 -5780 -25870
rect -5348 -26430 -5288 -25706
rect -4328 -25706 -4316 -25650
rect -4282 -25170 -4272 -25130
rect -3304 -25130 -3258 -25118
rect -4282 -25650 -4276 -25170
rect -4282 -25706 -4268 -25650
rect -3304 -25666 -3298 -25130
rect -5052 -25756 -4564 -25750
rect -5052 -25790 -5040 -25756
rect -4576 -25790 -4564 -25756
rect -5052 -25796 -4564 -25790
rect -4946 -25870 -4886 -25864
rect -4844 -25870 -4784 -25796
rect -4328 -25870 -4268 -25706
rect -3312 -25706 -3298 -25666
rect -3264 -25666 -3258 -25130
rect -3264 -25706 -3252 -25666
rect -4034 -25756 -3546 -25750
rect -4034 -25790 -4022 -25756
rect -3558 -25790 -3546 -25756
rect -4034 -25796 -3546 -25790
rect -3820 -25870 -3760 -25796
rect -3312 -25870 -3252 -25706
rect -2670 -25840 -2610 -23680
rect -2310 -23932 -2182 -23926
rect -2310 -23966 -2298 -23932
rect -2194 -23966 -2182 -23932
rect -2310 -23972 -2182 -23966
rect -2418 -24016 -2372 -24004
rect -2418 -24544 -2412 -24016
rect -2424 -24592 -2412 -24544
rect -2378 -24544 -2372 -24016
rect -2126 -24016 -2066 -23480
rect -1828 -23480 -1814 -23440
rect -1780 -22935 -1771 -22904
rect -1522 -22904 -1476 -22892
rect -1780 -23440 -1774 -23002
rect -1522 -23440 -1516 -22904
rect -1780 -23480 -1768 -23440
rect -1972 -23524 -1924 -23522
rect -2010 -23530 -1882 -23524
rect -2010 -23564 -1998 -23530
rect -1894 -23564 -1882 -23530
rect -2010 -23570 -1882 -23564
rect -1976 -23620 -1916 -23570
rect -1982 -23680 -1976 -23620
rect -1916 -23680 -1910 -23620
rect -1976 -23926 -1916 -23680
rect -2012 -23932 -1884 -23926
rect -2012 -23966 -2000 -23932
rect -1896 -23966 -1884 -23932
rect -2012 -23972 -1884 -23966
rect -2126 -24054 -2114 -24016
rect -2378 -24592 -2364 -24544
rect -2120 -24546 -2114 -24054
rect -2424 -24740 -2364 -24592
rect -2128 -24592 -2114 -24546
rect -2080 -24054 -2066 -24016
rect -1828 -24016 -1768 -23480
rect -1530 -23480 -1516 -23440
rect -1482 -23440 -1476 -22904
rect -1230 -22904 -1167 -22541
rect -1082 -22722 -1022 -22458
rect -940 -22674 -934 -22614
rect -874 -22674 -868 -22614
rect -1088 -22782 -1082 -22722
rect -1022 -22782 -1016 -22722
rect -1116 -22820 -988 -22814
rect -1116 -22854 -1104 -22820
rect -1000 -22854 -988 -22820
rect -1116 -22860 -988 -22854
rect -1230 -22917 -1218 -22904
rect -1482 -23480 -1470 -23440
rect -1224 -23480 -1218 -22962
rect -1184 -22917 -1167 -22904
rect -934 -22904 -874 -22674
rect -786 -22722 -726 -22458
rect -634 -22483 -576 -22368
rect -340 -22368 -324 -22326
rect -290 -22310 -284 -21792
rect -290 -22368 -278 -22310
rect -32 -22317 -26 -21878
rect -37 -22338 -26 -22317
rect -38 -22368 -26 -22338
rect 262 -21848 272 -21792
rect 8 -22317 14 -21878
rect 8 -22338 21 -22317
rect 8 -22368 22 -22338
rect -520 -22418 -392 -22412
rect -520 -22452 -508 -22418
rect -404 -22452 -392 -22418
rect -520 -22458 -392 -22452
rect -640 -22541 -634 -22483
rect -576 -22541 -570 -22483
rect -792 -22782 -786 -22722
rect -726 -22782 -720 -22722
rect -818 -22820 -690 -22814
rect -818 -22854 -806 -22820
rect -702 -22854 -690 -22820
rect -818 -22860 -690 -22854
rect -934 -22954 -920 -22904
rect -1184 -23480 -1178 -22962
rect -926 -23480 -920 -22954
rect -886 -22954 -874 -22904
rect -634 -22904 -576 -22541
rect -340 -22614 -280 -22368
rect -222 -22418 -94 -22412
rect -222 -22452 -210 -22418
rect -106 -22452 -94 -22418
rect -222 -22458 -94 -22452
rect -38 -22483 22 -22368
rect 266 -22368 272 -21848
rect 306 -21848 322 -21792
rect 564 -21792 610 -21780
rect 306 -22368 312 -21848
rect 564 -22323 570 -21792
rect 559 -22330 570 -22323
rect 266 -22380 312 -22368
rect 556 -22368 570 -22330
rect 604 -22323 610 -21792
rect 862 -21792 908 -21780
rect 604 -22368 617 -22323
rect 862 -22328 868 -21792
rect 76 -22418 204 -22412
rect 76 -22452 88 -22418
rect 192 -22452 204 -22418
rect 76 -22458 204 -22452
rect 374 -22418 502 -22412
rect 374 -22452 386 -22418
rect 490 -22452 502 -22418
rect 374 -22458 502 -22452
rect -38 -22541 -37 -22483
rect 21 -22541 22 -22483
rect -346 -22674 -340 -22614
rect -280 -22674 -274 -22614
rect -492 -22782 -486 -22722
rect -426 -22782 -420 -22722
rect -190 -22782 -184 -22722
rect -124 -22782 -118 -22722
rect -486 -22814 -426 -22782
rect -184 -22814 -124 -22782
rect -520 -22820 -392 -22814
rect -520 -22854 -508 -22820
rect -404 -22854 -392 -22820
rect -520 -22860 -392 -22854
rect -222 -22820 -94 -22814
rect -222 -22854 -210 -22820
rect -106 -22854 -94 -22820
rect -222 -22860 -94 -22854
rect -330 -22904 -284 -22892
rect -634 -22933 -622 -22904
rect -886 -23480 -880 -22954
rect -628 -23396 -622 -22933
rect -1712 -23530 -1584 -23524
rect -1712 -23564 -1700 -23530
rect -1596 -23564 -1584 -23530
rect -1712 -23570 -1584 -23564
rect -1530 -23728 -1470 -23480
rect -1414 -23530 -1286 -23524
rect -1414 -23564 -1402 -23530
rect -1298 -23564 -1286 -23530
rect -1414 -23570 -1286 -23564
rect -1536 -23788 -1530 -23728
rect -1470 -23788 -1464 -23728
rect -1714 -23932 -1586 -23926
rect -1714 -23966 -1702 -23932
rect -1598 -23966 -1586 -23932
rect -1714 -23972 -1586 -23966
rect -1828 -24054 -1816 -24016
rect -2080 -24542 -2074 -24054
rect -1822 -24534 -1816 -24054
rect -2080 -24592 -2060 -24542
rect -1828 -24592 -1816 -24538
rect -1782 -24054 -1768 -24016
rect -1530 -24016 -1470 -23788
rect -1416 -23932 -1288 -23926
rect -1416 -23966 -1404 -23932
rect -1300 -23966 -1288 -23932
rect -1416 -23972 -1288 -23966
rect -1230 -24016 -1170 -23480
rect -926 -23492 -880 -23480
rect -636 -23480 -622 -23474
rect -588 -22932 -572 -22904
rect -588 -22933 -576 -22932
rect -588 -23396 -582 -22933
rect -330 -23424 -324 -22904
rect -336 -23438 -324 -23424
rect -588 -23480 -576 -23474
rect -338 -23480 -324 -23438
rect -290 -23424 -284 -22904
rect -38 -22904 22 -22541
rect 106 -22722 166 -22458
rect 252 -22674 258 -22614
rect 318 -22674 324 -22614
rect 100 -22782 106 -22722
rect 166 -22782 172 -22722
rect 76 -22820 204 -22814
rect 76 -22854 88 -22820
rect 192 -22854 204 -22820
rect 76 -22860 204 -22854
rect -38 -22924 -26 -22904
rect -32 -23416 -26 -22974
rect -290 -23480 -276 -23424
rect 8 -22924 22 -22904
rect 258 -22904 318 -22674
rect 410 -22722 470 -22458
rect 556 -22483 617 -22368
rect 854 -22368 868 -22328
rect 902 -22328 908 -21792
rect 902 -22368 914 -22328
rect 672 -22418 800 -22412
rect 672 -22452 684 -22418
rect 788 -22452 800 -22418
rect 672 -22458 800 -22452
rect 556 -22492 559 -22483
rect 558 -22541 559 -22492
rect 710 -22486 770 -22458
rect 854 -22486 914 -22368
rect 617 -22541 914 -22486
rect 558 -22546 914 -22541
rect 558 -22698 618 -22546
rect 404 -22782 410 -22722
rect 470 -22782 476 -22722
rect 558 -22758 916 -22698
rect 374 -22820 502 -22814
rect 374 -22854 386 -22820
rect 490 -22854 502 -22820
rect 374 -22860 502 -22854
rect 258 -22954 272 -22904
rect 8 -23416 14 -22974
rect 266 -23480 272 -22954
rect 306 -22954 318 -22904
rect 558 -22904 618 -22758
rect 706 -22814 766 -22758
rect 672 -22820 800 -22814
rect 672 -22854 684 -22820
rect 788 -22854 800 -22820
rect 672 -22860 800 -22854
rect 558 -22936 570 -22904
rect 306 -23480 312 -22954
rect 564 -23402 570 -22936
rect -1116 -23530 -988 -23524
rect -1116 -23564 -1104 -23530
rect -1000 -23564 -988 -23530
rect -1116 -23570 -988 -23564
rect -818 -23530 -690 -23524
rect -818 -23564 -806 -23530
rect -702 -23564 -690 -23530
rect -818 -23570 -690 -23564
rect -1080 -23620 -1020 -23570
rect -786 -23620 -726 -23570
rect -1086 -23680 -1080 -23620
rect -1020 -23680 -1014 -23620
rect -792 -23680 -786 -23620
rect -726 -23680 -720 -23620
rect -1076 -23926 -1020 -23680
rect -786 -23926 -730 -23680
rect -1118 -23932 -990 -23926
rect -1118 -23966 -1106 -23932
rect -1002 -23966 -990 -23932
rect -1118 -23972 -990 -23966
rect -820 -23932 -692 -23926
rect -820 -23966 -808 -23932
rect -704 -23966 -692 -23932
rect -820 -23972 -692 -23966
rect -928 -24016 -882 -24004
rect -636 -24010 -576 -23480
rect -512 -23530 -392 -23524
rect -512 -23564 -508 -23530
rect -404 -23564 -392 -23530
rect -512 -23570 -392 -23564
rect -336 -23728 -276 -23480
rect -222 -23530 -96 -23524
rect -222 -23564 -210 -23530
rect -106 -23564 -96 -23530
rect -222 -23570 -96 -23564
rect -342 -23788 -336 -23728
rect -276 -23788 -270 -23728
rect -522 -23932 -394 -23926
rect -522 -23966 -510 -23932
rect -406 -23966 -394 -23932
rect -522 -23972 -394 -23966
rect -336 -24016 -276 -23788
rect -224 -23932 -96 -23926
rect -224 -23966 -212 -23932
rect -108 -23966 -96 -23932
rect -224 -23972 -96 -23966
rect -1530 -24054 -1518 -24016
rect -1782 -24534 -1776 -24054
rect -1524 -24534 -1518 -24054
rect -1782 -24592 -1768 -24538
rect -1484 -24054 -1470 -24016
rect -1484 -24534 -1478 -24054
rect -1226 -24532 -1220 -24056
rect -1234 -24592 -1220 -24532
rect -1186 -24532 -1180 -24056
rect -1186 -24592 -1174 -24532
rect -928 -24544 -922 -24016
rect -2310 -24642 -2182 -24636
rect -2310 -24676 -2298 -24642
rect -2194 -24676 -2182 -24642
rect -2310 -24682 -2182 -24676
rect -2278 -24740 -2218 -24682
rect -2128 -24740 -2068 -24592
rect -2012 -24642 -1884 -24636
rect -2012 -24676 -2000 -24642
rect -1896 -24676 -1884 -24642
rect -2012 -24682 -1884 -24676
rect -1828 -24712 -1768 -24592
rect -1714 -24642 -1586 -24636
rect -1714 -24676 -1702 -24642
rect -1598 -24676 -1586 -24642
rect -1714 -24682 -1586 -24676
rect -1416 -24642 -1288 -24636
rect -1416 -24676 -1404 -24642
rect -1300 -24676 -1288 -24642
rect -1416 -24682 -1288 -24676
rect -2424 -24800 -2068 -24740
rect -1834 -24772 -1828 -24712
rect -1768 -24772 -1762 -24712
rect -2426 -24806 -2364 -24800
rect -2366 -24860 -2364 -24806
rect -2426 -24872 -2366 -24866
rect -1984 -24974 -1978 -24914
rect -1918 -24974 -1912 -24914
rect -1978 -25036 -1918 -24974
rect -2310 -25042 -2182 -25036
rect -2310 -25076 -2298 -25042
rect -2194 -25076 -2182 -25042
rect -2310 -25082 -2182 -25076
rect -2012 -25042 -1884 -25036
rect -2012 -25076 -2000 -25042
rect -1896 -25076 -1884 -25042
rect -2012 -25082 -1884 -25076
rect -2418 -25126 -2372 -25114
rect -2418 -25650 -2412 -25126
rect -2426 -25702 -2412 -25650
rect -2378 -25650 -2372 -25126
rect -2120 -25126 -2074 -25114
rect -2378 -25702 -2366 -25650
rect -2120 -25654 -2114 -25126
rect -2426 -25840 -2366 -25702
rect -2126 -25702 -2114 -25654
rect -2080 -25654 -2074 -25126
rect -1828 -25126 -1768 -24772
rect -1680 -24914 -1620 -24682
rect -1540 -24866 -1534 -24806
rect -1474 -24866 -1468 -24806
rect -1686 -24974 -1680 -24914
rect -1620 -24974 -1614 -24914
rect -1714 -25042 -1586 -25036
rect -1714 -25076 -1702 -25042
rect -1598 -25076 -1586 -25042
rect -1714 -25082 -1586 -25076
rect -1828 -25170 -1816 -25126
rect -1822 -25654 -1816 -25170
rect -2080 -25702 -2066 -25654
rect -1782 -25170 -1768 -25126
rect -1534 -25126 -1474 -24866
rect -1384 -24914 -1324 -24682
rect -1234 -24712 -1174 -24592
rect -936 -24592 -922 -24544
rect -888 -24544 -882 -24016
rect -888 -24550 -876 -24544
rect -888 -24592 -870 -24550
rect -630 -24562 -624 -24044
rect -634 -24592 -624 -24562
rect -590 -24562 -584 -24044
rect -338 -24054 -326 -24016
rect -590 -24592 -574 -24562
rect -1118 -24642 -990 -24636
rect -1118 -24676 -1106 -24642
rect -1002 -24676 -990 -24642
rect -1118 -24682 -990 -24676
rect -1240 -24772 -1234 -24712
rect -1174 -24772 -1168 -24712
rect -1390 -24974 -1384 -24914
rect -1324 -24974 -1318 -24914
rect -1416 -25042 -1288 -25036
rect -1416 -25076 -1404 -25042
rect -1300 -25076 -1288 -25042
rect -1416 -25082 -1288 -25076
rect -1234 -25126 -1174 -24772
rect -936 -24806 -876 -24592
rect -820 -24642 -692 -24636
rect -820 -24676 -808 -24642
rect -704 -24676 -692 -24642
rect -820 -24682 -692 -24676
rect -634 -24712 -574 -24592
rect -332 -24592 -326 -24054
rect -292 -24054 -276 -24016
rect -42 -24016 18 -23480
rect 266 -23492 312 -23480
rect 554 -23480 570 -23436
rect 604 -22936 618 -22904
rect 856 -22904 916 -22758
rect 604 -23402 610 -22936
rect 856 -22940 868 -22904
rect 604 -23480 614 -23436
rect 862 -23440 868 -22940
rect 856 -23480 868 -23440
rect 902 -22940 916 -22904
rect 902 -23440 908 -22940
rect 902 -23480 916 -23440
rect 76 -23530 204 -23524
rect 76 -23564 88 -23530
rect 192 -23564 204 -23530
rect 76 -23570 204 -23564
rect 374 -23530 502 -23524
rect 374 -23564 386 -23530
rect 490 -23564 502 -23530
rect 374 -23570 502 -23564
rect 108 -23620 168 -23570
rect 410 -23620 470 -23570
rect 102 -23680 108 -23620
rect 168 -23680 174 -23620
rect 404 -23680 410 -23620
rect 470 -23680 476 -23620
rect 112 -23926 168 -23680
rect 414 -23926 470 -23680
rect 74 -23932 202 -23926
rect 74 -23966 86 -23932
rect 190 -23966 202 -23932
rect 74 -23972 202 -23966
rect 372 -23932 500 -23926
rect 372 -23966 384 -23932
rect 488 -23966 500 -23932
rect 372 -23972 500 -23966
rect -42 -24044 -28 -24016
rect -292 -24592 -286 -24054
rect -34 -24502 -28 -24044
rect -332 -24604 -286 -24592
rect -40 -24592 -28 -24538
rect 6 -24044 18 -24016
rect 264 -24016 310 -24004
rect 6 -24502 12 -24044
rect 6 -24592 20 -24538
rect 264 -24542 270 -24016
rect -522 -24642 -394 -24636
rect -522 -24676 -510 -24642
rect -406 -24676 -394 -24642
rect -522 -24682 -394 -24676
rect -224 -24642 -96 -24636
rect -224 -24676 -212 -24642
rect -108 -24676 -96 -24642
rect -224 -24682 -96 -24676
rect -640 -24772 -634 -24712
rect -574 -24772 -568 -24712
rect -942 -24866 -936 -24806
rect -876 -24866 -870 -24806
rect -1086 -24974 -1080 -24914
rect -1020 -24974 -1014 -24914
rect -790 -24974 -784 -24914
rect -724 -24974 -718 -24914
rect -1080 -25042 -1020 -24974
rect -784 -25042 -724 -24974
rect -634 -25126 -574 -24772
rect -486 -24914 -426 -24682
rect -344 -24866 -338 -24806
rect -278 -24866 -272 -24806
rect -492 -24974 -486 -24914
rect -426 -24974 -420 -24914
rect -522 -25042 -394 -25036
rect -522 -25076 -510 -25042
rect -406 -25076 -394 -25042
rect -522 -25082 -394 -25076
rect -1534 -25160 -1518 -25126
rect -1782 -25654 -1776 -25170
rect -1526 -25184 -1518 -25160
rect -1524 -25654 -1518 -25184
rect -1484 -25184 -1466 -25126
rect -1234 -25160 -1220 -25126
rect -1484 -25654 -1478 -25184
rect -1226 -25654 -1220 -25170
rect -1186 -25160 -1174 -25126
rect -1186 -25654 -1180 -25170
rect -928 -25662 -922 -25170
rect -936 -25664 -922 -25662
rect -938 -25702 -922 -25664
rect -634 -25158 -624 -25126
rect -888 -25662 -882 -25170
rect -630 -25638 -624 -25170
rect -888 -25702 -876 -25662
rect -590 -25158 -574 -25126
rect -338 -25126 -278 -24866
rect -190 -24914 -130 -24682
rect -40 -24712 20 -24592
rect 262 -24592 270 -24542
rect 304 -24542 310 -24016
rect 554 -24016 614 -23480
rect 672 -23530 800 -23524
rect 672 -23564 684 -23530
rect 788 -23564 800 -23530
rect 672 -23570 708 -23564
rect 768 -23570 800 -23564
rect 952 -23728 1012 -21540
rect 670 -23932 798 -23926
rect 670 -23966 682 -23932
rect 786 -23966 798 -23932
rect 670 -23972 798 -23966
rect 304 -24592 322 -24542
rect 74 -24642 202 -24636
rect 74 -24676 86 -24642
rect 190 -24676 202 -24642
rect 74 -24682 202 -24676
rect -46 -24772 -40 -24712
rect 20 -24772 26 -24712
rect -196 -24974 -190 -24914
rect -130 -24974 -124 -24914
rect -224 -25042 -96 -25036
rect -224 -25076 -212 -25042
rect -108 -25076 -96 -25042
rect -224 -25082 -96 -25076
rect -40 -25126 20 -24772
rect 262 -24806 322 -24592
rect 554 -24592 568 -24016
rect 602 -24052 618 -24016
rect 852 -24048 866 -24016
rect 602 -24592 614 -24052
rect 860 -24540 866 -24048
rect 852 -24562 866 -24540
rect 850 -24592 866 -24562
rect 900 -24048 912 -24016
rect 900 -24540 906 -24048
rect 900 -24592 912 -24540
rect 372 -24642 500 -24636
rect 372 -24676 384 -24642
rect 488 -24676 500 -24642
rect 372 -24682 500 -24676
rect 554 -24712 614 -24592
rect 670 -24642 798 -24636
rect 670 -24676 682 -24642
rect 786 -24676 798 -24642
rect 670 -24682 762 -24676
rect 764 -24682 798 -24676
rect 548 -24772 554 -24712
rect 614 -24716 620 -24712
rect 702 -24716 762 -24682
rect 852 -24716 912 -24592
rect 614 -24772 912 -24716
rect 554 -24776 912 -24772
rect 256 -24866 262 -24806
rect 322 -24866 328 -24806
rect 100 -24974 106 -24914
rect 166 -24974 172 -24914
rect 404 -24974 410 -24914
rect 470 -24974 476 -24914
rect 554 -24938 614 -24776
rect 106 -25036 166 -24974
rect 410 -25036 470 -24974
rect 554 -24998 914 -24938
rect 74 -25042 202 -25036
rect 74 -25076 86 -25042
rect 190 -25076 202 -25042
rect 74 -25082 202 -25076
rect 372 -25042 500 -25036
rect 372 -25076 384 -25042
rect 488 -25076 500 -25042
rect 372 -25082 500 -25076
rect -338 -25164 -326 -25126
rect -590 -25638 -584 -25170
rect -334 -25186 -326 -25164
rect -332 -25638 -326 -25186
rect -292 -25186 -274 -25126
rect -40 -25152 -28 -25126
rect -292 -25638 -286 -25186
rect -34 -25638 -28 -25152
rect 6 -25152 20 -25126
rect 264 -25126 310 -25114
rect 6 -25638 12 -25152
rect 264 -25654 270 -25126
rect 256 -25702 270 -25654
rect 304 -25654 310 -25126
rect 554 -25126 614 -24998
rect 704 -25036 764 -24998
rect 670 -25042 798 -25036
rect 670 -25076 682 -25042
rect 786 -25076 798 -25042
rect 670 -25082 798 -25076
rect 554 -25182 568 -25126
rect 304 -25666 316 -25654
rect 304 -25702 318 -25666
rect -2310 -25752 -2182 -25746
rect -2310 -25786 -2298 -25752
rect -2194 -25786 -2182 -25752
rect -2310 -25792 -2218 -25786
rect -2216 -25792 -2182 -25786
rect -2278 -25840 -2218 -25792
rect -2126 -25840 -2066 -25702
rect -2012 -25752 -1884 -25746
rect -1118 -25752 -990 -25746
rect -2012 -25786 -2000 -25752
rect -1896 -25786 -1884 -25752
rect -2012 -25792 -1884 -25786
rect -1714 -25786 -1702 -25758
rect -1598 -25786 -1586 -25758
rect -1714 -25792 -1586 -25786
rect -1416 -25786 -1404 -25758
rect -1300 -25786 -1288 -25758
rect -1416 -25792 -1288 -25786
rect -1118 -25786 -1106 -25752
rect -1002 -25786 -990 -25752
rect -1118 -25792 -990 -25786
rect -1680 -25840 -1620 -25792
rect -1382 -25840 -1322 -25792
rect -4886 -25930 -3252 -25870
rect -2676 -25900 -2670 -25840
rect -2610 -25900 -2604 -25840
rect -2426 -25900 -2066 -25840
rect -1686 -25900 -1680 -25840
rect -1620 -25900 -1614 -25840
rect -1388 -25900 -1382 -25840
rect -1322 -25900 -1316 -25840
rect -4946 -25936 -4886 -25930
rect -2126 -25940 -2066 -25900
rect -938 -25940 -878 -25702
rect -820 -25752 -692 -25746
rect -486 -25752 -426 -25750
rect 74 -25752 202 -25746
rect -820 -25786 -808 -25752
rect -704 -25786 -692 -25752
rect -820 -25792 -692 -25786
rect -522 -25786 -510 -25780
rect -406 -25786 -394 -25780
rect -522 -25792 -394 -25786
rect -224 -25786 -212 -25780
rect -108 -25786 -96 -25780
rect -224 -25792 -96 -25786
rect 74 -25786 86 -25752
rect 190 -25786 202 -25752
rect 74 -25792 202 -25786
rect -486 -25840 -426 -25792
rect -184 -25840 -124 -25792
rect -492 -25900 -486 -25840
rect -426 -25900 -420 -25840
rect -190 -25900 -184 -25840
rect -124 -25900 -118 -25840
rect 258 -25940 318 -25702
rect 562 -25702 568 -25182
rect 602 -25182 614 -25126
rect 854 -25126 914 -24998
rect 854 -25152 866 -25126
rect 602 -25702 608 -25182
rect 562 -25714 608 -25702
rect 860 -25702 866 -25152
rect 900 -25152 914 -25126
rect 900 -25702 906 -25152
rect 860 -25714 906 -25702
rect 372 -25752 500 -25746
rect 372 -25786 384 -25752
rect 488 -25786 500 -25752
rect 372 -25792 500 -25786
rect 670 -25752 798 -25746
rect 670 -25786 682 -25752
rect 786 -25786 798 -25752
rect 670 -25792 798 -25786
rect 952 -25940 1012 -23788
rect 1076 -22722 1136 -22716
rect 1076 -24914 1136 -22782
rect 1976 -23544 2036 -14060
rect 1970 -23604 1976 -23544
rect 2036 -23604 2042 -23544
rect 2110 -23762 2170 -13854
rect 2336 -15116 2396 -11416
rect 3070 -11594 22482 -11534
rect 3070 -11640 3130 -11594
rect 2864 -11646 3352 -11640
rect 2864 -11680 2876 -11646
rect 3340 -11680 3352 -11646
rect 2864 -11686 3352 -11680
rect 2576 -11730 2622 -11718
rect 2576 -12272 2582 -11730
rect 2568 -12306 2582 -12272
rect 2616 -12272 2622 -11730
rect 3586 -11730 3646 -11594
rect 4098 -11640 4158 -11594
rect 5106 -11640 5166 -11594
rect 3882 -11646 4370 -11640
rect 3882 -11680 3894 -11646
rect 4358 -11680 4370 -11646
rect 3882 -11686 4370 -11680
rect 4900 -11646 5388 -11640
rect 4900 -11680 4912 -11646
rect 5376 -11680 5388 -11646
rect 4900 -11686 5388 -11680
rect 2616 -12306 2628 -12272
rect 2568 -12448 2628 -12306
rect 3586 -12306 3600 -11730
rect 3634 -12306 3646 -11730
rect 4612 -11730 4658 -11718
rect 4612 -12268 4618 -11730
rect 2864 -12356 3352 -12350
rect 2864 -12390 2876 -12356
rect 3340 -12390 3352 -12356
rect 2864 -12396 3352 -12390
rect 2562 -12508 2568 -12448
rect 2628 -12508 2634 -12448
rect 2568 -12964 2628 -12508
rect 3076 -12874 3136 -12396
rect 3586 -12546 3646 -12306
rect 4604 -12306 4618 -12268
rect 4652 -12268 4658 -11730
rect 5624 -11730 5684 -11594
rect 6116 -11640 6176 -11594
rect 7128 -11640 7188 -11594
rect 5918 -11646 6406 -11640
rect 5918 -11680 5930 -11646
rect 6394 -11680 6406 -11646
rect 5918 -11686 6406 -11680
rect 6936 -11646 7424 -11640
rect 6936 -11680 6948 -11646
rect 7412 -11680 7424 -11646
rect 6936 -11686 7424 -11680
rect 4652 -12306 4664 -12268
rect 3882 -12356 4370 -12350
rect 3882 -12390 3894 -12356
rect 4358 -12390 4370 -12356
rect 3882 -12396 4370 -12390
rect 3580 -12606 3586 -12546
rect 3646 -12606 3652 -12546
rect 2864 -12880 3352 -12874
rect 2864 -12914 2876 -12880
rect 3340 -12914 3352 -12880
rect 2864 -12920 3352 -12914
rect 2568 -12998 2582 -12964
rect 2576 -13540 2582 -12998
rect 2616 -12998 2628 -12964
rect 3586 -12964 3646 -12606
rect 4078 -12874 4138 -12396
rect 4604 -12448 4664 -12306
rect 5624 -12306 5636 -11730
rect 5670 -12306 5684 -11730
rect 6648 -11730 6694 -11718
rect 6648 -12276 6654 -11730
rect 5100 -12350 5160 -12348
rect 4900 -12356 5388 -12350
rect 4900 -12390 4912 -12356
rect 5376 -12390 5388 -12356
rect 4900 -12396 5388 -12390
rect 4598 -12508 4604 -12448
rect 4664 -12508 4670 -12448
rect 3882 -12880 4370 -12874
rect 3882 -12914 3894 -12880
rect 4358 -12914 4370 -12880
rect 3882 -12920 4370 -12914
rect 2616 -13540 2622 -12998
rect 3586 -13012 3600 -12964
rect 2576 -13552 2622 -13540
rect 3594 -13540 3600 -13012
rect 3634 -13012 3646 -12964
rect 4604 -12964 4664 -12508
rect 5100 -12874 5160 -12396
rect 5624 -12546 5684 -12306
rect 6638 -12306 6654 -12276
rect 6688 -12276 6694 -11730
rect 7658 -11730 7718 -11594
rect 8176 -11640 8236 -11594
rect 9164 -11640 9224 -11594
rect 7954 -11646 8442 -11640
rect 7954 -11680 7966 -11646
rect 8430 -11680 8442 -11646
rect 7954 -11686 8442 -11680
rect 8972 -11646 9460 -11640
rect 8972 -11680 8984 -11646
rect 9448 -11680 9460 -11646
rect 8972 -11686 9460 -11680
rect 6688 -12306 6698 -12276
rect 5918 -12356 6406 -12350
rect 5918 -12390 5930 -12356
rect 6394 -12390 6406 -12356
rect 5918 -12396 6406 -12390
rect 6638 -12448 6698 -12306
rect 7658 -12306 7672 -11730
rect 7706 -12306 7718 -11730
rect 8684 -11730 8730 -11718
rect 8684 -12262 8690 -11730
rect 6936 -12356 7424 -12350
rect 6936 -12390 6948 -12356
rect 7412 -12390 7424 -12356
rect 6936 -12396 7424 -12390
rect 6632 -12508 6638 -12448
rect 6698 -12508 6704 -12448
rect 7658 -12546 7718 -12306
rect 8678 -12306 8690 -12262
rect 8724 -12262 8730 -11730
rect 9692 -11730 9752 -11594
rect 10208 -11640 10268 -11594
rect 11210 -11640 11270 -11594
rect 9990 -11646 10478 -11640
rect 9990 -11680 10002 -11646
rect 10466 -11680 10478 -11646
rect 9990 -11686 10478 -11680
rect 11008 -11646 11496 -11640
rect 11008 -11680 11020 -11646
rect 11484 -11680 11496 -11646
rect 11008 -11686 11496 -11680
rect 8724 -12306 8738 -12262
rect 7954 -12356 8442 -12350
rect 7954 -12390 7966 -12356
rect 8430 -12390 8442 -12356
rect 7954 -12396 8442 -12390
rect 8678 -12448 8738 -12306
rect 9692 -12306 9708 -11730
rect 9742 -12306 9752 -11730
rect 10720 -11730 10766 -11718
rect 10720 -12266 10726 -11730
rect 8972 -12356 9460 -12350
rect 8972 -12390 8984 -12356
rect 9448 -12390 9460 -12356
rect 8972 -12396 9460 -12390
rect 8672 -12508 8678 -12448
rect 8738 -12508 8744 -12448
rect 9692 -12546 9752 -12306
rect 10714 -12306 10726 -12266
rect 10760 -12266 10766 -11730
rect 11732 -11730 11792 -11594
rect 12238 -11640 12298 -11594
rect 13256 -11640 13316 -11594
rect 12026 -11646 12514 -11640
rect 12026 -11680 12038 -11646
rect 12502 -11680 12514 -11646
rect 12026 -11686 12514 -11680
rect 13044 -11646 13532 -11640
rect 13044 -11680 13056 -11646
rect 13520 -11680 13532 -11646
rect 13044 -11686 13532 -11680
rect 12238 -11688 12298 -11686
rect 10760 -12306 10774 -12266
rect 9990 -12356 10478 -12350
rect 9990 -12390 10002 -12356
rect 10466 -12390 10478 -12356
rect 9990 -12396 10478 -12390
rect 10714 -12448 10774 -12306
rect 11732 -12306 11744 -11730
rect 11778 -12306 11792 -11730
rect 12756 -11730 12802 -11718
rect 12756 -12266 12762 -11730
rect 11008 -12356 11496 -12350
rect 11008 -12390 11020 -12356
rect 11484 -12390 11496 -12356
rect 11008 -12396 11496 -12390
rect 10708 -12508 10714 -12448
rect 10774 -12508 10780 -12448
rect 11732 -12546 11792 -12306
rect 12748 -12306 12762 -12266
rect 12796 -12266 12802 -11730
rect 13766 -11730 13826 -11594
rect 14274 -11640 14334 -11594
rect 15294 -11640 15354 -11594
rect 14062 -11646 14550 -11640
rect 14062 -11680 14074 -11646
rect 14538 -11680 14550 -11646
rect 14062 -11686 14550 -11680
rect 15080 -11646 15568 -11640
rect 15080 -11680 15092 -11646
rect 15556 -11680 15568 -11646
rect 15080 -11686 15568 -11680
rect 12796 -12306 12808 -12266
rect 12026 -12356 12514 -12350
rect 12026 -12390 12038 -12356
rect 12502 -12390 12514 -12356
rect 12026 -12396 12514 -12390
rect 12748 -12448 12808 -12306
rect 13766 -12306 13780 -11730
rect 13814 -12306 13826 -11730
rect 14792 -11730 14838 -11718
rect 14792 -12260 14798 -11730
rect 13044 -12356 13532 -12350
rect 13044 -12390 13056 -12356
rect 13520 -12390 13532 -12356
rect 13044 -12396 13532 -12390
rect 12742 -12508 12748 -12448
rect 12808 -12508 12814 -12448
rect 13766 -12546 13826 -12306
rect 14784 -12306 14798 -12260
rect 14832 -12260 14838 -11730
rect 15804 -11730 15864 -11594
rect 16302 -11640 16362 -11594
rect 17330 -11640 17390 -11594
rect 16098 -11646 16586 -11640
rect 16098 -11680 16110 -11646
rect 16574 -11680 16586 -11646
rect 16098 -11686 16586 -11680
rect 17116 -11646 17604 -11640
rect 17116 -11680 17128 -11646
rect 17592 -11680 17604 -11646
rect 17116 -11686 17604 -11680
rect 14832 -12306 14844 -12260
rect 14062 -12356 14550 -12350
rect 14062 -12390 14074 -12356
rect 14538 -12390 14550 -12356
rect 14062 -12396 14550 -12390
rect 14784 -12448 14844 -12306
rect 15804 -12306 15816 -11730
rect 15850 -12306 15864 -11730
rect 16828 -11730 16874 -11718
rect 16828 -12258 16834 -11730
rect 15080 -12356 15568 -12350
rect 15080 -12390 15092 -12356
rect 15556 -12390 15568 -12356
rect 15080 -12396 15568 -12390
rect 14778 -12508 14784 -12448
rect 14844 -12508 14850 -12448
rect 15804 -12546 15864 -12306
rect 16820 -12306 16834 -12258
rect 16868 -12258 16874 -11730
rect 17836 -11730 17896 -11594
rect 18332 -11640 18392 -11594
rect 19362 -11640 19422 -11594
rect 18134 -11646 18622 -11640
rect 18134 -11680 18146 -11646
rect 18610 -11680 18622 -11646
rect 18134 -11686 18622 -11680
rect 19152 -11646 19640 -11640
rect 19152 -11680 19164 -11646
rect 19628 -11680 19640 -11646
rect 19152 -11686 19640 -11680
rect 16868 -12306 16880 -12258
rect 16098 -12356 16586 -12350
rect 16098 -12390 16110 -12356
rect 16574 -12390 16586 -12356
rect 16098 -12396 16586 -12390
rect 16820 -12448 16880 -12306
rect 17836 -12306 17852 -11730
rect 17886 -12306 17896 -11730
rect 18864 -11730 18910 -11718
rect 18864 -12252 18870 -11730
rect 17116 -12356 17604 -12350
rect 17116 -12390 17128 -12356
rect 17592 -12390 17604 -12356
rect 17116 -12396 17604 -12390
rect 16814 -12508 16820 -12448
rect 16880 -12508 16886 -12448
rect 17836 -12546 17896 -12306
rect 18856 -12306 18870 -12252
rect 18904 -12252 18910 -11730
rect 19874 -11730 19934 -11594
rect 20410 -11640 20470 -11594
rect 21384 -11640 21444 -11594
rect 20170 -11646 20658 -11640
rect 20170 -11680 20182 -11646
rect 20646 -11680 20658 -11646
rect 20170 -11686 20658 -11680
rect 21188 -11646 21676 -11640
rect 21188 -11680 21200 -11646
rect 21664 -11680 21676 -11646
rect 21188 -11686 21676 -11680
rect 18904 -12306 18916 -12252
rect 18134 -12356 18622 -12350
rect 18134 -12390 18146 -12356
rect 18610 -12390 18622 -12356
rect 18134 -12396 18622 -12390
rect 18856 -12448 18916 -12306
rect 19874 -12306 19888 -11730
rect 19922 -12306 19934 -11730
rect 20900 -11730 20946 -11718
rect 20900 -12260 20906 -11730
rect 19152 -12356 19640 -12350
rect 19152 -12390 19164 -12356
rect 19628 -12390 19640 -12356
rect 19152 -12396 19640 -12390
rect 18850 -12508 18856 -12448
rect 18916 -12508 18922 -12448
rect 19874 -12546 19934 -12306
rect 20894 -12306 20906 -12260
rect 20940 -12260 20946 -11730
rect 21912 -11730 21972 -11594
rect 22422 -11640 22482 -11594
rect 22206 -11646 22694 -11640
rect 22206 -11680 22218 -11646
rect 22682 -11680 22694 -11646
rect 22206 -11686 22694 -11680
rect 20940 -12306 20954 -12260
rect 20170 -12356 20658 -12350
rect 20170 -12390 20182 -12356
rect 20646 -12390 20658 -12356
rect 20170 -12396 20658 -12390
rect 5618 -12606 5624 -12546
rect 5684 -12606 5690 -12546
rect 7652 -12606 7658 -12546
rect 7718 -12606 7724 -12546
rect 9686 -12606 9692 -12546
rect 9752 -12606 9758 -12546
rect 11726 -12606 11732 -12546
rect 11792 -12606 11798 -12546
rect 13760 -12606 13766 -12546
rect 13826 -12606 13832 -12546
rect 15798 -12606 15804 -12546
rect 15864 -12606 15870 -12546
rect 17830 -12606 17836 -12546
rect 17896 -12606 17902 -12546
rect 19868 -12606 19874 -12546
rect 19934 -12606 19940 -12546
rect 12218 -12660 12278 -12652
rect 12218 -12720 14326 -12660
rect 9190 -12838 10260 -12778
rect 11726 -12818 11732 -12758
rect 11792 -12818 11798 -12758
rect 9190 -12874 9250 -12838
rect 4900 -12880 5388 -12874
rect 4900 -12914 4912 -12880
rect 5376 -12914 5388 -12880
rect 4900 -12920 5388 -12914
rect 5918 -12880 6406 -12874
rect 5918 -12914 5930 -12880
rect 6394 -12914 6406 -12880
rect 5918 -12920 6406 -12914
rect 6936 -12880 7424 -12874
rect 6936 -12914 6948 -12880
rect 7412 -12914 7424 -12880
rect 6936 -12920 7424 -12914
rect 7954 -12880 8162 -12874
rect 8222 -12880 8442 -12874
rect 7954 -12914 7966 -12880
rect 8430 -12914 8442 -12880
rect 7954 -12920 8442 -12914
rect 8972 -12880 9460 -12874
rect 8972 -12914 8984 -12880
rect 9448 -12914 9460 -12880
rect 8972 -12920 9460 -12914
rect 4604 -12996 4618 -12964
rect 3634 -13540 3640 -13012
rect 3594 -13552 3640 -13540
rect 4612 -13540 4618 -12996
rect 4652 -12996 4664 -12964
rect 5630 -12964 5676 -12952
rect 4652 -13540 4658 -12996
rect 5630 -13512 5636 -12964
rect 4612 -13552 4658 -13540
rect 5624 -13540 5636 -13512
rect 5670 -13512 5676 -12964
rect 6648 -12964 6694 -12952
rect 8684 -12964 8730 -12952
rect 6648 -13492 6654 -12964
rect 5670 -13540 5684 -13512
rect 2864 -13590 3352 -13584
rect 2864 -13624 2876 -13590
rect 3340 -13624 3352 -13590
rect 2864 -13630 3352 -13624
rect 3882 -13590 4370 -13584
rect 3882 -13624 3894 -13590
rect 4358 -13624 4370 -13590
rect 3882 -13630 4370 -13624
rect 4900 -13590 5388 -13584
rect 4900 -13624 4912 -13590
rect 5376 -13624 5388 -13590
rect 4900 -13630 5388 -13624
rect 5624 -13682 5684 -13540
rect 6642 -13540 6654 -13492
rect 6688 -13492 6694 -12964
rect 7656 -12998 7672 -12964
rect 7666 -13464 7672 -12998
rect 6688 -13540 6702 -13492
rect 5918 -13590 6406 -13584
rect 5918 -13624 5930 -13590
rect 6394 -13624 6406 -13590
rect 5918 -13630 6406 -13624
rect 6272 -13678 6332 -13630
rect 6642 -13678 6702 -13540
rect 7656 -13540 7672 -13464
rect 7706 -12998 7716 -12964
rect 7706 -13464 7712 -12998
rect 7706 -13480 7716 -13464
rect 7706 -13540 7720 -13480
rect 8684 -13484 8690 -12964
rect 8676 -13540 8690 -13484
rect 8724 -13484 8730 -12964
rect 9696 -12964 9756 -12838
rect 10200 -12874 10260 -12838
rect 9990 -12880 10478 -12874
rect 9990 -12914 10002 -12880
rect 10466 -12914 10478 -12880
rect 9990 -12920 10478 -12914
rect 11008 -12880 11496 -12874
rect 11008 -12914 11020 -12880
rect 11484 -12914 11496 -12880
rect 11008 -12920 11496 -12914
rect 9696 -13014 9708 -12964
rect 8724 -13540 8736 -13484
rect 9702 -13490 9708 -13014
rect 9696 -13504 9708 -13490
rect 6936 -13590 7424 -13584
rect 6936 -13624 6948 -13590
rect 7412 -13624 7424 -13590
rect 6936 -13630 7424 -13624
rect 7144 -13678 7204 -13630
rect 7656 -13678 7716 -13540
rect 7954 -13590 8442 -13584
rect 7954 -13624 7966 -13590
rect 8430 -13624 8442 -13590
rect 7954 -13630 8442 -13624
rect 8184 -13678 8244 -13630
rect 8676 -13678 8736 -13540
rect 9694 -13540 9708 -13504
rect 9742 -13014 9756 -12964
rect 10720 -12964 10766 -12952
rect 9742 -13490 9748 -13014
rect 10720 -13464 10726 -12964
rect 9742 -13540 9756 -13490
rect 10708 -13540 10726 -13464
rect 10760 -13464 10766 -12964
rect 11732 -12964 11792 -12818
rect 12218 -12874 12278 -12720
rect 13252 -12874 13312 -12720
rect 13758 -12818 13764 -12758
rect 13824 -12818 13830 -12758
rect 12026 -12880 12514 -12874
rect 12026 -12914 12038 -12880
rect 12502 -12914 12514 -12880
rect 12026 -12920 12514 -12914
rect 13044 -12880 13532 -12874
rect 13044 -12914 13056 -12880
rect 13520 -12914 13532 -12880
rect 13044 -12920 13532 -12914
rect 11732 -12998 11744 -12964
rect 10760 -13540 10768 -13464
rect 11738 -13478 11744 -12998
rect 11732 -13482 11744 -13478
rect 8972 -13590 9460 -13584
rect 8972 -13624 8984 -13590
rect 9448 -13624 9460 -13590
rect 8972 -13630 9460 -13624
rect 5624 -13742 6196 -13682
rect 6266 -13738 6272 -13678
rect 6332 -13738 6338 -13678
rect 6636 -13738 6642 -13678
rect 6702 -13738 6708 -13678
rect 7138 -13738 7144 -13678
rect 7204 -13738 7210 -13678
rect 7650 -13738 7656 -13678
rect 7716 -13738 7722 -13678
rect 8178 -13738 8184 -13678
rect 8244 -13738 8250 -13678
rect 8670 -13738 8676 -13678
rect 8736 -13738 8742 -13678
rect 4090 -13848 4096 -13788
rect 4156 -13848 4162 -13788
rect 5112 -13848 5118 -13788
rect 5178 -13848 5184 -13788
rect 2566 -14060 2572 -14000
rect 2632 -14060 2638 -14000
rect 3064 -14060 3070 -14000
rect 3130 -14060 3136 -14000
rect 3576 -14060 3582 -14000
rect 3642 -14060 3648 -14000
rect 2572 -14196 2632 -14060
rect 3070 -14106 3130 -14060
rect 2864 -14112 3352 -14106
rect 2864 -14146 2876 -14112
rect 3340 -14146 3352 -14112
rect 2864 -14152 3352 -14146
rect 2572 -14236 2582 -14196
rect 2576 -14772 2582 -14236
rect 2616 -14236 2632 -14196
rect 3582 -14196 3642 -14060
rect 4096 -14106 4156 -13848
rect 5118 -14106 5178 -13848
rect 6136 -13886 6196 -13742
rect 6136 -13892 6198 -13886
rect 6136 -13952 6138 -13892
rect 6136 -13958 6198 -13952
rect 5618 -14060 5624 -14000
rect 5684 -14060 5690 -14000
rect 3882 -14112 4370 -14106
rect 3882 -14146 3894 -14112
rect 4358 -14146 4370 -14112
rect 3882 -14152 4370 -14146
rect 4900 -14112 5388 -14106
rect 4900 -14146 4912 -14112
rect 5376 -14146 5388 -14112
rect 4900 -14152 5388 -14146
rect 2616 -14772 2622 -14236
rect 3582 -14242 3600 -14196
rect 2576 -14784 2622 -14772
rect 3594 -14772 3600 -14242
rect 3634 -14242 3642 -14196
rect 4612 -14196 4658 -14184
rect 3634 -14772 3640 -14242
rect 4612 -14714 4618 -14196
rect 3594 -14784 3640 -14772
rect 4598 -14772 4618 -14714
rect 4652 -14772 4658 -14196
rect 5624 -14196 5684 -14060
rect 6136 -14106 6196 -13958
rect 5918 -14112 6406 -14106
rect 5918 -14146 5930 -14112
rect 6394 -14146 6406 -14112
rect 5918 -14152 6406 -14146
rect 5624 -14248 5636 -14196
rect 2864 -14822 3352 -14816
rect 2864 -14856 2876 -14822
rect 3340 -14856 3352 -14822
rect 2864 -14862 3352 -14856
rect 3882 -14822 4370 -14816
rect 3882 -14856 3894 -14822
rect 4358 -14856 4370 -14822
rect 3882 -14862 4370 -14856
rect 4080 -14962 4086 -14902
rect 4146 -14962 4152 -14902
rect 2330 -15176 2336 -15116
rect 2396 -15176 2402 -15116
rect 2336 -16358 2396 -15176
rect 2568 -15272 3646 -15212
rect 2568 -15430 2628 -15272
rect 3076 -15340 3136 -15272
rect 2862 -15346 3350 -15340
rect 2862 -15380 2874 -15346
rect 3338 -15380 3350 -15346
rect 2862 -15386 3350 -15380
rect 2568 -15456 2580 -15430
rect 2574 -16006 2580 -15456
rect 2614 -15456 2628 -15430
rect 3586 -15430 3646 -15272
rect 4086 -15340 4146 -14962
rect 4598 -14994 4658 -14772
rect 5630 -14772 5636 -14248
rect 5670 -14248 5684 -14196
rect 6642 -14196 6702 -13738
rect 7132 -13952 7138 -13892
rect 7198 -13952 7204 -13892
rect 8152 -13952 8158 -13892
rect 8218 -13952 8224 -13892
rect 7138 -14106 7198 -13952
rect 7652 -14060 7658 -14000
rect 7718 -14060 7724 -14000
rect 6936 -14112 7424 -14106
rect 6936 -14146 6948 -14112
rect 7412 -14146 7424 -14112
rect 6936 -14152 7424 -14146
rect 5670 -14772 5676 -14248
rect 6642 -14260 6654 -14196
rect 6648 -14708 6654 -14260
rect 5630 -14784 5676 -14772
rect 6634 -14772 6654 -14708
rect 6688 -14260 6702 -14196
rect 7658 -14196 7718 -14060
rect 8158 -14106 8218 -13952
rect 7954 -14112 8442 -14106
rect 7954 -14146 7966 -14112
rect 8430 -14146 8442 -14112
rect 7954 -14152 8442 -14146
rect 7658 -14230 7672 -14196
rect 6688 -14772 6694 -14260
rect 4900 -14822 5388 -14816
rect 4900 -14856 4912 -14822
rect 5376 -14856 5388 -14822
rect 4900 -14862 5388 -14856
rect 5918 -14822 6120 -14816
rect 6122 -14822 6406 -14816
rect 5918 -14856 5930 -14822
rect 6394 -14856 6406 -14822
rect 5918 -14862 6120 -14856
rect 6122 -14862 6406 -14856
rect 6122 -14890 6182 -14862
rect 5096 -14950 5102 -14890
rect 5162 -14950 5168 -14890
rect 6116 -14950 6122 -14890
rect 6182 -14950 6188 -14890
rect 4592 -15054 4598 -14994
rect 4658 -15054 4664 -14994
rect 4598 -15288 4604 -15228
rect 4664 -15288 4670 -15228
rect 3880 -15346 4368 -15340
rect 3880 -15380 3892 -15346
rect 4356 -15380 4368 -15346
rect 3880 -15386 4368 -15380
rect 2614 -16006 2620 -15456
rect 3586 -15462 3598 -15430
rect 3592 -15962 3598 -15462
rect 2574 -16018 2620 -16006
rect 3586 -16006 3598 -15962
rect 3632 -15462 3646 -15430
rect 4604 -15430 4664 -15288
rect 5102 -15340 5162 -14950
rect 5616 -15054 5622 -14994
rect 5682 -15054 5688 -14994
rect 4898 -15346 5386 -15340
rect 4898 -15380 4910 -15346
rect 5374 -15380 5386 -15346
rect 4898 -15386 5386 -15380
rect 4604 -15456 4616 -15430
rect 3632 -15962 3638 -15462
rect 3632 -16006 3646 -15962
rect 2862 -16056 3350 -16050
rect 2862 -16090 2874 -16056
rect 3338 -16090 3350 -16056
rect 2862 -16096 3350 -16090
rect 3586 -16158 3646 -16006
rect 4610 -16006 4616 -15456
rect 4650 -15456 4664 -15430
rect 5622 -15430 5682 -15054
rect 6122 -15340 6182 -14950
rect 6634 -14994 6694 -14772
rect 7666 -14772 7672 -14230
rect 7706 -14230 7718 -14196
rect 8676 -14196 8736 -13738
rect 9190 -13788 9250 -13630
rect 9694 -13788 9754 -13540
rect 9990 -13590 10478 -13584
rect 9990 -13624 10002 -13590
rect 10466 -13624 10478 -13590
rect 9990 -13630 10478 -13624
rect 10210 -13788 10270 -13630
rect 10708 -13678 10768 -13540
rect 11730 -13540 11744 -13482
rect 11778 -12998 11792 -12964
rect 12756 -12964 12802 -12952
rect 11778 -13478 11784 -12998
rect 12756 -13474 12762 -12964
rect 11778 -13540 11792 -13478
rect 12744 -13540 12762 -13474
rect 12796 -13474 12802 -12964
rect 13764 -12964 13824 -12818
rect 14266 -12874 14326 -12720
rect 15290 -12808 16372 -12748
rect 15290 -12874 15350 -12808
rect 14062 -12880 14550 -12874
rect 14062 -12914 14074 -12880
rect 14538 -12914 14550 -12880
rect 14062 -12920 14550 -12914
rect 15080 -12880 15568 -12874
rect 15080 -12914 15092 -12880
rect 15556 -12914 15568 -12880
rect 15080 -12920 15568 -12914
rect 13764 -12998 13780 -12964
rect 12796 -13540 12804 -13474
rect 13774 -13514 13780 -12998
rect 11008 -13590 11496 -13584
rect 11008 -13624 11020 -13590
rect 11484 -13624 11496 -13590
rect 11008 -13630 11496 -13624
rect 10702 -13738 10708 -13678
rect 10768 -13738 10774 -13678
rect 9184 -13848 9190 -13788
rect 9250 -13848 9256 -13788
rect 9688 -13848 9694 -13788
rect 9754 -13848 9760 -13788
rect 10204 -13848 10210 -13788
rect 10270 -13848 10276 -13788
rect 9190 -14106 9250 -13848
rect 9686 -14060 9692 -14000
rect 9752 -14060 9758 -14000
rect 8972 -14112 9460 -14106
rect 8972 -14146 8984 -14112
rect 9448 -14146 9460 -14112
rect 8972 -14152 9460 -14146
rect 7706 -14772 7712 -14230
rect 8676 -14238 8690 -14196
rect 8684 -14730 8690 -14238
rect 7666 -14784 7712 -14772
rect 8676 -14772 8690 -14730
rect 8724 -14238 8736 -14196
rect 9692 -14196 9752 -14060
rect 10210 -14106 10270 -13848
rect 9990 -14112 10478 -14106
rect 9990 -14146 10002 -14112
rect 10466 -14146 10478 -14112
rect 9990 -14152 10478 -14146
rect 8724 -14730 8730 -14238
rect 9692 -14258 9708 -14196
rect 8724 -14772 8736 -14730
rect 6936 -14822 7424 -14816
rect 6936 -14856 6948 -14822
rect 7412 -14856 7424 -14822
rect 6936 -14862 7132 -14856
rect 7134 -14862 7424 -14856
rect 7954 -14822 8442 -14816
rect 7954 -14856 7966 -14822
rect 8430 -14856 8442 -14822
rect 7954 -14862 8442 -14856
rect 7134 -14890 7194 -14862
rect 8160 -14890 8220 -14862
rect 7128 -14950 7134 -14890
rect 7194 -14950 7200 -14890
rect 8154 -14950 8160 -14890
rect 8220 -14950 8226 -14890
rect 6628 -15054 6634 -14994
rect 6694 -15054 6700 -14994
rect 6634 -15288 6640 -15228
rect 6700 -15288 6706 -15228
rect 5916 -15346 6120 -15340
rect 6122 -15346 6404 -15340
rect 5916 -15380 5928 -15346
rect 6392 -15380 6404 -15346
rect 5916 -15386 6404 -15380
rect 4650 -16006 4656 -15456
rect 5622 -15462 5634 -15430
rect 5628 -15966 5634 -15462
rect 4610 -16018 4656 -16006
rect 5620 -16006 5634 -15966
rect 5668 -15462 5682 -15430
rect 6640 -15430 6700 -15288
rect 7134 -15340 7194 -14950
rect 7648 -15054 7654 -14994
rect 7714 -15054 7720 -14994
rect 6934 -15346 7132 -15340
rect 7134 -15346 7422 -15340
rect 6934 -15380 6946 -15346
rect 7410 -15380 7422 -15346
rect 6934 -15386 7422 -15380
rect 6640 -15460 6652 -15430
rect 5668 -15966 5674 -15462
rect 5668 -16006 5680 -15966
rect 3880 -16056 4368 -16050
rect 3880 -16090 3892 -16056
rect 4356 -16090 4368 -16056
rect 3880 -16096 4368 -16090
rect 4898 -16056 5386 -16050
rect 4898 -16090 4910 -16056
rect 5374 -16090 5386 -16056
rect 4898 -16096 5386 -16090
rect 2442 -16218 2448 -16158
rect 2508 -16218 2514 -16158
rect 3580 -16218 3586 -16158
rect 3646 -16218 3652 -16158
rect 2330 -16418 2336 -16358
rect 2396 -16418 2402 -16358
rect 2224 -16520 2230 -16460
rect 2290 -16520 2296 -16460
rect 2230 -19950 2290 -16520
rect 2336 -17594 2396 -16418
rect 2330 -17654 2336 -17594
rect 2396 -17654 2402 -17594
rect 2224 -20010 2230 -19950
rect 2290 -20010 2296 -19950
rect 2230 -21254 2290 -20010
rect 2336 -20196 2396 -17654
rect 2448 -18932 2508 -16218
rect 3578 -16418 3584 -16358
rect 3644 -16418 3650 -16358
rect 3584 -16462 3644 -16418
rect 2568 -16522 3644 -16462
rect 2568 -16524 3132 -16522
rect 2568 -16664 2628 -16524
rect 3072 -16574 3132 -16524
rect 2862 -16580 3350 -16574
rect 2862 -16614 2874 -16580
rect 3338 -16614 3350 -16580
rect 2862 -16620 3350 -16614
rect 2568 -16696 2580 -16664
rect 2574 -17240 2580 -16696
rect 2614 -16696 2628 -16664
rect 3584 -16664 3644 -16522
rect 4088 -16574 4148 -16096
rect 4596 -16298 4602 -16238
rect 4662 -16298 4668 -16238
rect 3880 -16580 4368 -16574
rect 3880 -16614 3892 -16580
rect 4356 -16614 4368 -16580
rect 3880 -16620 4368 -16614
rect 2614 -17240 2620 -16696
rect 3584 -16700 3598 -16664
rect 2574 -17252 2620 -17240
rect 3592 -17240 3598 -16700
rect 3632 -16700 3644 -16664
rect 4602 -16664 4662 -16298
rect 5116 -16352 5176 -16096
rect 5620 -16134 5680 -16006
rect 6646 -16006 6652 -15460
rect 6686 -15460 6700 -15430
rect 7654 -15430 7714 -15054
rect 8160 -15340 8220 -14950
rect 8676 -14994 8736 -14772
rect 9702 -14772 9708 -14258
rect 9742 -14258 9752 -14196
rect 10708 -14196 10768 -13738
rect 11230 -13788 11290 -13630
rect 11730 -13676 11790 -13540
rect 12026 -13590 12514 -13584
rect 12026 -13624 12038 -13590
rect 12502 -13624 12514 -13590
rect 12026 -13630 12514 -13624
rect 11730 -13736 11908 -13676
rect 11224 -13848 11230 -13788
rect 11290 -13848 11296 -13788
rect 11726 -13848 11732 -13788
rect 11792 -13848 11798 -13788
rect 11230 -14106 11290 -13848
rect 11008 -14112 11496 -14106
rect 11008 -14146 11020 -14112
rect 11484 -14146 11496 -14112
rect 11008 -14152 11496 -14146
rect 11732 -14196 11792 -13848
rect 11848 -14000 11908 -13736
rect 12226 -13848 12232 -13788
rect 12292 -13848 12298 -13788
rect 11848 -14066 11908 -14060
rect 12232 -14106 12292 -13848
rect 12372 -13892 12432 -13630
rect 12744 -13678 12804 -13540
rect 13766 -13540 13780 -13514
rect 13814 -12998 13824 -12964
rect 14792 -12964 14838 -12952
rect 13814 -13514 13820 -12998
rect 14792 -13480 14798 -12964
rect 13814 -13540 13826 -13514
rect 13044 -13590 13532 -13584
rect 13044 -13624 13056 -13590
rect 13520 -13624 13532 -13590
rect 13044 -13630 13532 -13624
rect 12738 -13738 12744 -13678
rect 12804 -13738 12810 -13678
rect 12366 -13952 12372 -13892
rect 12432 -13952 12438 -13892
rect 12026 -14112 12514 -14106
rect 12026 -14146 12038 -14112
rect 12502 -14146 12514 -14112
rect 12026 -14152 12514 -14146
rect 10708 -14252 10726 -14196
rect 9742 -14772 9748 -14258
rect 10720 -14730 10726 -14252
rect 9702 -14784 9748 -14772
rect 10712 -14772 10726 -14730
rect 10760 -14252 10768 -14196
rect 11728 -14248 11744 -14196
rect 10760 -14730 10766 -14252
rect 11738 -14648 11744 -14248
rect 10760 -14772 10772 -14730
rect 8972 -14822 9460 -14816
rect 8972 -14856 8984 -14822
rect 9448 -14856 9460 -14822
rect 8972 -14862 9460 -14856
rect 9990 -14822 10478 -14816
rect 9990 -14856 10002 -14822
rect 10466 -14856 10478 -14822
rect 9990 -14862 10478 -14856
rect 10712 -14994 10772 -14772
rect 11730 -14772 11744 -14724
rect 11778 -14240 11792 -14196
rect 12744 -14196 12804 -13738
rect 13252 -13848 13258 -13788
rect 13318 -13848 13324 -13788
rect 13258 -14106 13318 -13848
rect 13380 -13892 13440 -13630
rect 13766 -13676 13826 -13540
rect 14780 -13540 14798 -13480
rect 14832 -13480 14838 -12964
rect 15802 -12964 15862 -12808
rect 16312 -12874 16372 -12808
rect 17328 -12808 17900 -12748
rect 17328 -12874 17388 -12808
rect 16098 -12880 16586 -12874
rect 16098 -12914 16110 -12880
rect 16574 -12914 16586 -12880
rect 16098 -12920 16586 -12914
rect 17116 -12880 17604 -12874
rect 17116 -12914 17128 -12880
rect 17592 -12914 17604 -12880
rect 17116 -12920 17604 -12914
rect 15802 -13004 15816 -12964
rect 15810 -13474 15816 -13004
rect 14832 -13540 14840 -13480
rect 14062 -13590 14550 -13584
rect 14062 -13624 14074 -13590
rect 14538 -13624 14550 -13590
rect 14062 -13630 14550 -13624
rect 13572 -13736 13826 -13676
rect 13374 -13952 13380 -13892
rect 13440 -13952 13446 -13892
rect 13572 -14002 13632 -13736
rect 13762 -13848 13768 -13788
rect 13828 -13848 13834 -13788
rect 14270 -13848 14276 -13788
rect 14336 -13848 14342 -13788
rect 13572 -14068 13632 -14062
rect 13044 -14112 13532 -14106
rect 13044 -14146 13056 -14112
rect 13520 -14146 13532 -14112
rect 13044 -14152 13532 -14146
rect 13768 -14196 13828 -13848
rect 14276 -14106 14336 -13848
rect 14422 -13892 14482 -13630
rect 14780 -13678 14840 -13540
rect 15806 -13540 15816 -13474
rect 15850 -13004 15862 -12964
rect 16828 -12964 16874 -12952
rect 15850 -13474 15856 -13004
rect 15850 -13540 15866 -13474
rect 16828 -13490 16834 -12964
rect 15080 -13590 15568 -13584
rect 15080 -13624 15092 -13590
rect 15556 -13624 15568 -13590
rect 15080 -13630 15568 -13624
rect 14774 -13738 14780 -13678
rect 14840 -13738 14846 -13678
rect 14416 -13952 14422 -13892
rect 14482 -13952 14488 -13892
rect 14062 -14112 14550 -14106
rect 14062 -14146 14074 -14112
rect 14538 -14146 14550 -14112
rect 14062 -14152 14550 -14146
rect 14780 -14196 14840 -13738
rect 15284 -13788 15344 -13630
rect 15806 -13788 15866 -13540
rect 16818 -13540 16834 -13490
rect 16868 -13490 16874 -12964
rect 17840 -12964 17900 -12808
rect 18134 -12880 18622 -12874
rect 18134 -12914 18146 -12880
rect 18610 -12914 18622 -12880
rect 18134 -12920 18622 -12914
rect 19152 -12880 19640 -12874
rect 19152 -12914 19164 -12880
rect 19628 -12914 19640 -12880
rect 19152 -12920 19640 -12914
rect 17840 -12990 17852 -12964
rect 17846 -13484 17852 -12990
rect 16868 -13540 16878 -13490
rect 17838 -13540 17852 -13484
rect 17886 -12990 17900 -12964
rect 18864 -12964 18910 -12952
rect 17886 -13484 17892 -12990
rect 17886 -13486 17898 -13484
rect 17886 -13540 17900 -13486
rect 18864 -13504 18870 -12964
rect 16296 -13584 16356 -13582
rect 16098 -13590 16586 -13584
rect 16098 -13624 16110 -13590
rect 16574 -13624 16586 -13590
rect 16098 -13630 16586 -13624
rect 16296 -13788 16356 -13630
rect 16818 -13678 16878 -13540
rect 17328 -13584 17388 -13582
rect 17116 -13590 17604 -13584
rect 17116 -13624 17128 -13590
rect 17592 -13624 17604 -13590
rect 17116 -13630 17604 -13624
rect 16812 -13738 16818 -13678
rect 16878 -13738 16884 -13678
rect 15278 -13848 15284 -13788
rect 15344 -13848 15350 -13788
rect 15800 -13848 15806 -13788
rect 15866 -13848 15872 -13788
rect 16290 -13848 16296 -13788
rect 16356 -13848 16362 -13788
rect 15284 -14106 15344 -13848
rect 15800 -14060 15806 -14000
rect 15866 -14060 15872 -14000
rect 15080 -14112 15568 -14106
rect 15080 -14146 15092 -14112
rect 15556 -14146 15568 -14112
rect 15080 -14152 15568 -14146
rect 11778 -14248 11788 -14240
rect 12744 -14244 12762 -14196
rect 11778 -14648 11784 -14248
rect 12756 -14724 12762 -14244
rect 11778 -14772 11790 -14724
rect 11008 -14822 11176 -14816
rect 11008 -14856 11020 -14822
rect 11008 -14862 11176 -14856
rect 11212 -14922 11272 -14856
rect 11730 -14922 11790 -14772
rect 12750 -14772 12762 -14724
rect 12796 -14244 12804 -14196
rect 13764 -14236 13780 -14196
rect 12796 -14724 12802 -14244
rect 13774 -14658 13780 -14236
rect 12796 -14772 12810 -14724
rect 12424 -14822 12514 -14816
rect 12502 -14856 12514 -14822
rect 12232 -14922 12292 -14856
rect 12424 -14862 12514 -14856
rect 11212 -14982 12292 -14922
rect 12750 -14994 12810 -14772
rect 13768 -14772 13780 -14754
rect 13814 -14234 13830 -14196
rect 13814 -14236 13828 -14234
rect 13814 -14658 13820 -14236
rect 14780 -14242 14798 -14196
rect 14792 -14718 14798 -14242
rect 13814 -14772 13828 -14754
rect 13044 -14822 13236 -14816
rect 13044 -14856 13056 -14822
rect 13044 -14862 13236 -14856
rect 13256 -14918 13316 -14856
rect 13768 -14918 13828 -14772
rect 14780 -14772 14798 -14718
rect 14832 -14242 14840 -14196
rect 15806 -14196 15866 -14060
rect 16296 -14106 16356 -13848
rect 16098 -14112 16586 -14106
rect 16098 -14146 16110 -14112
rect 16574 -14146 16586 -14112
rect 16098 -14152 16586 -14146
rect 15806 -14238 15816 -14196
rect 14832 -14718 14838 -14242
rect 14832 -14772 14840 -14718
rect 14062 -14822 14550 -14816
rect 14538 -14856 14550 -14822
rect 14062 -14862 14550 -14856
rect 14258 -14918 14318 -14862
rect 13256 -14978 14318 -14918
rect 14780 -14994 14840 -14772
rect 15810 -14772 15816 -14238
rect 15850 -14238 15866 -14196
rect 16818 -14196 16878 -13738
rect 17328 -13788 17388 -13630
rect 17840 -13788 17900 -13540
rect 18856 -13540 18870 -13504
rect 18904 -13504 18910 -12964
rect 19874 -12964 19934 -12606
rect 20378 -12874 20438 -12396
rect 20894 -12448 20954 -12306
rect 21912 -12306 21924 -11730
rect 21958 -12306 21972 -11730
rect 22936 -11730 22982 -11718
rect 22936 -12252 22942 -11730
rect 21188 -12356 21676 -12350
rect 21188 -12390 21200 -12356
rect 21664 -12390 21676 -12356
rect 21188 -12396 21676 -12390
rect 20888 -12508 20894 -12448
rect 20954 -12508 20960 -12448
rect 20170 -12880 20658 -12874
rect 20170 -12914 20182 -12880
rect 20646 -12914 20658 -12880
rect 20170 -12920 20658 -12914
rect 19874 -13004 19888 -12964
rect 18904 -13540 18916 -13504
rect 18134 -13590 18622 -13584
rect 18134 -13624 18146 -13590
rect 18610 -13624 18622 -13590
rect 18134 -13630 18622 -13624
rect 18342 -13678 18402 -13630
rect 18856 -13678 18916 -13540
rect 19882 -13540 19888 -13004
rect 19922 -13004 19934 -12964
rect 20894 -12964 20954 -12508
rect 21404 -12874 21464 -12396
rect 21912 -12546 21972 -12306
rect 22924 -12306 22942 -12252
rect 22976 -12252 22982 -11730
rect 24816 -12070 24928 -11284
rect 22976 -12306 22984 -12252
rect 22206 -12356 22694 -12350
rect 22206 -12390 22218 -12356
rect 22682 -12390 22694 -12356
rect 22206 -12396 22694 -12390
rect 21906 -12606 21912 -12546
rect 21972 -12606 21978 -12546
rect 21188 -12880 21676 -12874
rect 21188 -12914 21200 -12880
rect 21664 -12914 21676 -12880
rect 21188 -12920 21676 -12914
rect 20894 -12996 20906 -12964
rect 19922 -13540 19928 -13004
rect 19882 -13552 19928 -13540
rect 20900 -13540 20906 -12996
rect 20940 -12996 20954 -12964
rect 21912 -12964 21972 -12606
rect 22426 -12874 22486 -12396
rect 22924 -12448 22984 -12306
rect 22918 -12508 22924 -12448
rect 22984 -12508 22990 -12448
rect 22206 -12880 22694 -12874
rect 22206 -12914 22218 -12880
rect 22682 -12914 22694 -12880
rect 22206 -12920 22694 -12914
rect 21912 -12992 21924 -12964
rect 20940 -13540 20946 -12996
rect 20900 -13552 20946 -13540
rect 21918 -13540 21924 -12992
rect 21958 -12992 21972 -12964
rect 22924 -12964 22984 -12508
rect 23642 -12606 23648 -12546
rect 23708 -12606 23714 -12546
rect 22924 -12990 22942 -12964
rect 21958 -13540 21964 -12992
rect 21918 -13552 21964 -13540
rect 22936 -13540 22942 -12990
rect 22976 -12990 22984 -12964
rect 22976 -13540 22982 -12990
rect 22936 -13552 22982 -13540
rect 19152 -13590 19640 -13584
rect 19152 -13624 19164 -13590
rect 19628 -13624 19640 -13590
rect 19152 -13630 19640 -13624
rect 20170 -13590 20658 -13584
rect 20170 -13624 20182 -13590
rect 20646 -13624 20658 -13590
rect 20170 -13630 20658 -13624
rect 21188 -13590 21676 -13584
rect 21188 -13624 21200 -13590
rect 21664 -13624 21676 -13590
rect 21188 -13630 21676 -13624
rect 22206 -13590 22694 -13584
rect 22206 -13624 22218 -13590
rect 22682 -13624 22694 -13590
rect 22206 -13630 22694 -13624
rect 19364 -13678 19424 -13630
rect 18850 -13738 18856 -13678
rect 18916 -13738 18922 -13678
rect 19358 -13738 19364 -13678
rect 19424 -13738 19430 -13678
rect 18342 -13744 18402 -13738
rect 17322 -13848 17328 -13788
rect 17388 -13848 17394 -13788
rect 17834 -13848 17840 -13788
rect 17900 -13848 17906 -13788
rect 17308 -13952 17314 -13892
rect 17374 -13952 17380 -13892
rect 18346 -13952 18352 -13892
rect 18412 -13952 18418 -13892
rect 17314 -14106 17374 -13952
rect 17832 -14060 17838 -14000
rect 17898 -14060 17904 -14000
rect 17116 -14112 17604 -14106
rect 17116 -14146 17128 -14112
rect 17592 -14146 17604 -14112
rect 17116 -14152 17604 -14146
rect 15850 -14772 15856 -14238
rect 15810 -14784 15856 -14772
rect 16818 -14772 16834 -14196
rect 16868 -14772 16878 -14196
rect 17838 -14196 17898 -14060
rect 18352 -14106 18412 -13952
rect 18134 -14112 18622 -14106
rect 18134 -14146 18146 -14112
rect 18610 -14146 18622 -14112
rect 18134 -14152 18622 -14146
rect 17838 -14238 17852 -14196
rect 15080 -14822 15568 -14816
rect 15080 -14856 15092 -14822
rect 15556 -14856 15568 -14822
rect 15080 -14862 15568 -14856
rect 16098 -14822 16586 -14816
rect 16098 -14856 16110 -14822
rect 16574 -14856 16586 -14822
rect 16098 -14862 16586 -14856
rect 15304 -14964 16366 -14904
rect 8670 -15054 8676 -14994
rect 8736 -15054 8742 -14994
rect 10706 -15054 10712 -14994
rect 10772 -15054 10778 -14994
rect 12744 -15054 12750 -14994
rect 12810 -15054 12816 -14994
rect 14774 -15054 14780 -14994
rect 14840 -15054 14846 -14994
rect 9690 -15176 9696 -15116
rect 9756 -15176 9762 -15116
rect 11724 -15176 11730 -15116
rect 11790 -15176 11796 -15116
rect 13754 -15176 13760 -15116
rect 13820 -15176 13826 -15116
rect 7952 -15346 8440 -15340
rect 7952 -15380 7964 -15346
rect 8428 -15380 8440 -15346
rect 7952 -15386 8440 -15380
rect 8970 -15346 9458 -15340
rect 8970 -15380 8982 -15346
rect 9446 -15380 9458 -15346
rect 8970 -15386 9458 -15380
rect 6686 -16006 6692 -15460
rect 7654 -15474 7670 -15430
rect 7664 -15956 7670 -15474
rect 6646 -16018 6692 -16006
rect 7656 -16006 7670 -15956
rect 7704 -15474 7714 -15430
rect 8682 -15430 8728 -15418
rect 7704 -15956 7710 -15474
rect 7704 -16006 7716 -15956
rect 8682 -15970 8688 -15430
rect 5916 -16056 6404 -16050
rect 5916 -16090 5928 -16056
rect 6392 -16090 6404 -16056
rect 5916 -16096 6404 -16090
rect 6934 -16056 7422 -16050
rect 6934 -16090 6946 -16056
rect 7410 -16090 7422 -16056
rect 6934 -16096 7422 -16090
rect 5614 -16194 5620 -16134
rect 5680 -16194 5686 -16134
rect 5110 -16412 5116 -16352
rect 5176 -16412 5182 -16352
rect 5116 -16574 5176 -16412
rect 4898 -16580 5386 -16574
rect 4898 -16614 4910 -16580
rect 5374 -16614 5386 -16580
rect 4898 -16620 5386 -16614
rect 3632 -17240 3638 -16700
rect 4602 -16706 4616 -16664
rect 4610 -17182 4616 -16706
rect 3592 -17252 3638 -17240
rect 4604 -17240 4616 -17182
rect 4650 -16706 4662 -16664
rect 5620 -16664 5680 -16194
rect 6118 -16346 6178 -16096
rect 6636 -16298 6642 -16238
rect 6702 -16298 6708 -16238
rect 6118 -16352 6180 -16346
rect 6118 -16412 6120 -16352
rect 6118 -16418 6180 -16412
rect 6118 -16574 6178 -16418
rect 5916 -16580 6404 -16574
rect 5916 -16614 5928 -16580
rect 6392 -16614 6404 -16580
rect 5916 -16620 6404 -16614
rect 4650 -17182 4656 -16706
rect 5620 -16708 5634 -16664
rect 4650 -17240 4664 -17182
rect 5628 -17192 5634 -16708
rect 2862 -17290 3350 -17284
rect 2862 -17324 2874 -17290
rect 3338 -17324 3350 -17290
rect 2862 -17330 3350 -17324
rect 3880 -17290 4368 -17284
rect 3880 -17324 3892 -17290
rect 4356 -17324 4368 -17290
rect 3880 -17330 4368 -17324
rect 3578 -17450 3584 -17390
rect 3644 -17450 3650 -17390
rect 2862 -17812 3350 -17806
rect 2862 -17846 2874 -17812
rect 3338 -17846 3350 -17812
rect 2862 -17852 3350 -17846
rect 2574 -17896 2620 -17884
rect 2574 -18426 2580 -17896
rect 2564 -18472 2580 -18426
rect 2614 -18426 2620 -17896
rect 3584 -17896 3644 -17450
rect 4090 -17492 4150 -17330
rect 4084 -17552 4090 -17492
rect 4150 -17552 4156 -17492
rect 4604 -17694 4664 -17240
rect 5622 -17240 5634 -17192
rect 5668 -16708 5680 -16664
rect 6642 -16664 6702 -16298
rect 7134 -16346 7194 -16096
rect 7656 -16134 7716 -16006
rect 8674 -16006 8688 -15970
rect 8722 -15970 8728 -15430
rect 9696 -15430 9756 -15176
rect 9988 -15346 10476 -15340
rect 9988 -15380 10000 -15346
rect 10464 -15380 10476 -15346
rect 9988 -15386 10476 -15380
rect 11006 -15346 11494 -15340
rect 11006 -15380 11018 -15346
rect 11482 -15380 11494 -15346
rect 11006 -15386 11494 -15380
rect 9696 -15486 9706 -15430
rect 8722 -16006 8734 -15970
rect 7952 -16056 8440 -16050
rect 7952 -16090 7964 -16056
rect 8428 -16090 8440 -16056
rect 7952 -16096 8440 -16090
rect 7650 -16194 7656 -16134
rect 7716 -16194 7722 -16134
rect 7132 -16352 7194 -16346
rect 7192 -16412 7194 -16352
rect 7132 -16418 7194 -16412
rect 7134 -16574 7194 -16418
rect 6934 -16580 7422 -16574
rect 6934 -16614 6946 -16580
rect 7410 -16614 7422 -16580
rect 6934 -16620 7422 -16614
rect 6642 -16706 6652 -16664
rect 5668 -17192 5674 -16708
rect 5668 -17240 5682 -17192
rect 4898 -17290 5386 -17284
rect 4898 -17324 4910 -17290
rect 5374 -17324 5386 -17290
rect 4898 -17330 5386 -17324
rect 5622 -17390 5682 -17240
rect 6646 -17240 6652 -16706
rect 6686 -16706 6702 -16664
rect 7656 -16664 7716 -16194
rect 8152 -16352 8212 -16096
rect 8674 -16238 8734 -16006
rect 9700 -16006 9706 -15486
rect 9740 -15486 9756 -15430
rect 10718 -15430 10764 -15418
rect 9740 -16006 9746 -15486
rect 10718 -15976 10724 -15430
rect 9700 -16018 9746 -16006
rect 10708 -16006 10724 -15976
rect 10758 -15976 10764 -15430
rect 11730 -15430 11790 -15176
rect 12024 -15346 12512 -15340
rect 12024 -15380 12036 -15346
rect 12500 -15380 12512 -15346
rect 12024 -15386 12512 -15380
rect 13042 -15346 13530 -15340
rect 13042 -15380 13054 -15346
rect 13518 -15380 13530 -15346
rect 13042 -15386 13530 -15380
rect 11730 -15480 11742 -15430
rect 10758 -16006 10768 -15976
rect 8970 -16056 9458 -16050
rect 8970 -16090 8982 -16056
rect 9446 -16090 9458 -16056
rect 8970 -16096 9458 -16090
rect 9988 -16056 10476 -16050
rect 9988 -16090 10000 -16056
rect 10464 -16090 10476 -16056
rect 9988 -16096 10476 -16090
rect 8668 -16298 8674 -16238
rect 8734 -16298 8740 -16238
rect 9164 -16294 9224 -16096
rect 10206 -16294 10266 -16096
rect 10708 -16238 10768 -16006
rect 11736 -16006 11742 -15480
rect 11776 -15480 11790 -15430
rect 12754 -15430 12800 -15418
rect 11776 -16006 11782 -15480
rect 12754 -15964 12760 -15430
rect 11736 -16018 11782 -16006
rect 12748 -16006 12760 -15964
rect 12794 -15964 12800 -15430
rect 13760 -15430 13820 -15176
rect 15304 -15340 15364 -14964
rect 15794 -15054 15800 -14994
rect 15860 -15054 15866 -14994
rect 14060 -15346 14548 -15340
rect 14060 -15380 14072 -15346
rect 14536 -15380 14548 -15346
rect 14060 -15386 14548 -15380
rect 15078 -15346 15566 -15340
rect 15078 -15380 15090 -15346
rect 15554 -15380 15566 -15346
rect 15078 -15386 15566 -15380
rect 13760 -15474 13778 -15430
rect 12794 -16006 12808 -15964
rect 11006 -16056 11494 -16050
rect 11006 -16090 11018 -16056
rect 11482 -16090 11494 -16056
rect 11006 -16096 11494 -16090
rect 12024 -16056 12512 -16050
rect 12024 -16090 12036 -16056
rect 12500 -16090 12512 -16056
rect 12024 -16096 12512 -16090
rect 8668 -16410 8674 -16350
rect 8734 -16410 8740 -16350
rect 9164 -16354 10266 -16294
rect 10702 -16298 10708 -16238
rect 10768 -16298 10774 -16238
rect 8152 -16574 8212 -16412
rect 7952 -16580 8440 -16574
rect 7952 -16614 7964 -16580
rect 8428 -16614 8440 -16580
rect 7952 -16620 8440 -16614
rect 6686 -17240 6692 -16706
rect 7656 -16712 7670 -16664
rect 7664 -17190 7670 -16712
rect 6646 -17252 6692 -17240
rect 7658 -17240 7670 -17190
rect 7704 -16712 7716 -16664
rect 8674 -16664 8734 -16410
rect 9164 -16574 9224 -16354
rect 9686 -16520 9692 -16460
rect 9752 -16520 9758 -16460
rect 8970 -16580 9458 -16574
rect 8970 -16614 8982 -16580
rect 9446 -16614 9458 -16580
rect 8970 -16620 9458 -16614
rect 7704 -17190 7710 -16712
rect 8674 -16722 8688 -16664
rect 7704 -17240 7718 -17190
rect 5916 -17290 6404 -17284
rect 5916 -17324 5928 -17290
rect 6392 -17324 6404 -17290
rect 5916 -17330 6404 -17324
rect 6934 -17290 7422 -17284
rect 6934 -17324 6946 -17290
rect 7410 -17324 7422 -17290
rect 6934 -17330 7422 -17324
rect 5616 -17450 5622 -17390
rect 5682 -17450 5688 -17390
rect 5614 -17654 5620 -17594
rect 5680 -17654 5686 -17594
rect 6128 -17600 6188 -17330
rect 7150 -17600 7210 -17330
rect 7658 -17390 7718 -17240
rect 8682 -17240 8688 -16722
rect 8722 -16722 8734 -16664
rect 9692 -16664 9752 -16520
rect 10206 -16574 10266 -16354
rect 10704 -16410 10710 -16350
rect 10770 -16410 10776 -16350
rect 9988 -16580 10476 -16574
rect 9988 -16614 10000 -16580
rect 10464 -16614 10476 -16580
rect 9988 -16620 10476 -16614
rect 9692 -16710 9706 -16664
rect 8722 -17240 8728 -16722
rect 8682 -17252 8728 -17240
rect 9700 -17240 9706 -16710
rect 9740 -16710 9752 -16664
rect 10710 -16664 10770 -16410
rect 11206 -16574 11266 -16096
rect 11720 -16520 11726 -16460
rect 11786 -16520 11792 -16460
rect 11006 -16580 11494 -16574
rect 11006 -16614 11018 -16580
rect 11482 -16614 11494 -16580
rect 11006 -16620 11494 -16614
rect 9740 -17240 9746 -16710
rect 10710 -16732 10724 -16664
rect 9700 -17252 9746 -17240
rect 10718 -17240 10724 -16732
rect 10758 -16732 10770 -16664
rect 11726 -16664 11786 -16520
rect 12240 -16574 12300 -16096
rect 12748 -16238 12808 -16006
rect 13772 -16006 13778 -15474
rect 13812 -15474 13820 -15430
rect 14790 -15430 14836 -15418
rect 13812 -16006 13818 -15474
rect 14790 -15954 14796 -15430
rect 13772 -16018 13818 -16006
rect 14782 -16006 14796 -15954
rect 14830 -15954 14836 -15430
rect 15800 -15430 15860 -15054
rect 16306 -15170 16366 -14964
rect 16818 -14994 16878 -14772
rect 17846 -14772 17852 -14238
rect 17886 -14238 17898 -14196
rect 18856 -14196 18916 -13738
rect 20378 -13848 20384 -13788
rect 20444 -13848 20450 -13788
rect 21398 -13848 21404 -13788
rect 21464 -13848 21470 -13788
rect 19346 -13952 19352 -13892
rect 19412 -13952 19418 -13892
rect 19352 -14106 19412 -13952
rect 19864 -14060 19870 -14000
rect 19930 -14060 19936 -14000
rect 19152 -14112 19640 -14106
rect 19152 -14146 19164 -14112
rect 19628 -14146 19640 -14112
rect 19152 -14152 19640 -14146
rect 19352 -14164 19412 -14152
rect 17886 -14772 17892 -14238
rect 18856 -14254 18870 -14196
rect 18864 -14724 18870 -14254
rect 17846 -14784 17892 -14772
rect 18854 -14772 18870 -14724
rect 18904 -14254 18916 -14196
rect 19870 -14196 19930 -14060
rect 20384 -14106 20444 -13848
rect 21404 -14106 21464 -13848
rect 21906 -14060 21912 -14000
rect 21972 -14060 21978 -14000
rect 22410 -14060 22416 -14000
rect 22476 -14060 22482 -14000
rect 22920 -14060 22926 -14000
rect 22986 -14060 22992 -14000
rect 20170 -14112 20658 -14106
rect 20170 -14146 20182 -14112
rect 20646 -14146 20658 -14112
rect 20170 -14152 20658 -14146
rect 21188 -14112 21676 -14106
rect 21188 -14146 21200 -14112
rect 21664 -14146 21676 -14112
rect 21188 -14152 21676 -14146
rect 19870 -14242 19888 -14196
rect 18904 -14724 18910 -14254
rect 18904 -14772 18914 -14724
rect 17116 -14822 17604 -14816
rect 17116 -14856 17128 -14822
rect 17318 -14856 17378 -14854
rect 17592 -14856 17604 -14822
rect 17116 -14862 17604 -14856
rect 18134 -14822 18622 -14816
rect 18134 -14856 18146 -14822
rect 18352 -14856 18412 -14850
rect 18610 -14856 18622 -14822
rect 18134 -14862 18622 -14856
rect 17318 -14890 17378 -14862
rect 18352 -14890 18412 -14862
rect 17310 -14950 17316 -14890
rect 17376 -14950 17382 -14890
rect 18346 -14950 18352 -14890
rect 18412 -14950 18418 -14890
rect 16812 -15054 16818 -14994
rect 16878 -15054 16884 -14994
rect 17318 -15170 17378 -14950
rect 17832 -15054 17838 -14994
rect 17898 -15054 17904 -14994
rect 16306 -15230 17378 -15170
rect 16306 -15340 16366 -15230
rect 17318 -15340 17378 -15230
rect 16096 -15346 16584 -15340
rect 16096 -15380 16108 -15346
rect 16572 -15380 16584 -15346
rect 16096 -15386 16584 -15380
rect 17114 -15346 17602 -15340
rect 17114 -15380 17126 -15346
rect 17590 -15380 17602 -15346
rect 17114 -15386 17602 -15380
rect 15800 -15478 15814 -15430
rect 14830 -16006 14842 -15954
rect 15808 -15974 15814 -15478
rect 13042 -16056 13530 -16050
rect 13042 -16090 13054 -16056
rect 13518 -16090 13530 -16056
rect 13042 -16096 13530 -16090
rect 14060 -16056 14548 -16050
rect 14060 -16090 14072 -16056
rect 14536 -16090 14548 -16056
rect 14060 -16096 14548 -16090
rect 12742 -16298 12748 -16238
rect 12808 -16298 12814 -16238
rect 13262 -16294 13322 -16096
rect 14270 -16294 14330 -16096
rect 14782 -16238 14842 -16006
rect 15800 -16006 15814 -15974
rect 15848 -15478 15860 -15430
rect 16826 -15430 16872 -15418
rect 15848 -15974 15854 -15478
rect 16826 -15970 16832 -15430
rect 15848 -16006 15860 -15974
rect 15078 -16056 15566 -16050
rect 15078 -16090 15090 -16056
rect 15554 -16090 15566 -16056
rect 15078 -16096 15566 -16090
rect 12740 -16410 12746 -16350
rect 12806 -16410 12812 -16350
rect 13262 -16354 14330 -16294
rect 14776 -16298 14782 -16238
rect 14842 -16298 14848 -16238
rect 14972 -16302 14978 -16242
rect 15038 -16302 15044 -16242
rect 12024 -16580 12512 -16574
rect 12024 -16614 12036 -16580
rect 12500 -16614 12512 -16580
rect 12024 -16620 12512 -16614
rect 11726 -16712 11742 -16664
rect 10758 -17240 10764 -16732
rect 10718 -17252 10764 -17240
rect 11736 -17240 11742 -16712
rect 11776 -16712 11786 -16664
rect 12746 -16664 12806 -16410
rect 13262 -16574 13322 -16354
rect 13760 -16520 13766 -16460
rect 13826 -16520 13832 -16460
rect 13042 -16580 13530 -16574
rect 13042 -16614 13054 -16580
rect 13518 -16614 13530 -16580
rect 13042 -16620 13530 -16614
rect 11776 -17240 11782 -16712
rect 12746 -16714 12760 -16664
rect 11736 -17252 11782 -17240
rect 12754 -17240 12760 -16714
rect 12794 -16714 12806 -16664
rect 13766 -16664 13826 -16520
rect 14270 -16574 14330 -16354
rect 14776 -16410 14782 -16350
rect 14842 -16410 14848 -16350
rect 14060 -16580 14548 -16574
rect 14060 -16614 14072 -16580
rect 14536 -16614 14548 -16580
rect 14060 -16620 14548 -16614
rect 13766 -16702 13778 -16664
rect 12794 -17240 12800 -16714
rect 13772 -17194 13778 -16702
rect 12754 -17252 12800 -17240
rect 13766 -17240 13778 -17194
rect 13812 -16702 13826 -16664
rect 14782 -16664 14842 -16410
rect 14978 -16460 15038 -16302
rect 15272 -16458 15332 -16096
rect 15800 -16134 15860 -16006
rect 16816 -16006 16832 -15970
rect 16866 -15970 16872 -15430
rect 17838 -15430 17898 -15054
rect 18352 -15178 18412 -14950
rect 18854 -14994 18914 -14772
rect 19882 -14772 19888 -14242
rect 19922 -14242 19930 -14196
rect 20900 -14196 20946 -14184
rect 19922 -14772 19928 -14242
rect 20900 -14714 20906 -14196
rect 19882 -14784 19928 -14772
rect 20890 -14772 20906 -14714
rect 20940 -14714 20946 -14196
rect 21912 -14196 21972 -14060
rect 22416 -14106 22476 -14060
rect 22206 -14112 22694 -14106
rect 22206 -14146 22218 -14112
rect 22682 -14146 22694 -14112
rect 22206 -14152 22694 -14146
rect 21912 -14252 21924 -14196
rect 20940 -14772 20950 -14714
rect 19152 -14822 19640 -14816
rect 19152 -14856 19164 -14822
rect 19628 -14856 19640 -14822
rect 19152 -14862 19640 -14856
rect 20170 -14822 20658 -14816
rect 20170 -14856 20182 -14822
rect 20646 -14856 20658 -14822
rect 20170 -14862 20658 -14856
rect 19368 -14890 19428 -14862
rect 19362 -14950 19368 -14890
rect 19428 -14950 19434 -14890
rect 20890 -14994 20950 -14772
rect 21918 -14772 21924 -14252
rect 21958 -14252 21972 -14196
rect 22926 -14196 22986 -14060
rect 22926 -14232 22942 -14196
rect 21958 -14772 21964 -14252
rect 21918 -14784 21964 -14772
rect 22936 -14772 22942 -14232
rect 22976 -14232 22986 -14196
rect 22976 -14772 22982 -14232
rect 22936 -14784 22982 -14772
rect 21188 -14822 21676 -14816
rect 21188 -14856 21200 -14822
rect 21664 -14856 21676 -14822
rect 21188 -14862 21676 -14856
rect 22206 -14822 22694 -14816
rect 22206 -14856 22218 -14822
rect 22682 -14856 22694 -14822
rect 22206 -14862 22694 -14856
rect 18848 -15054 18854 -14994
rect 18914 -15054 18920 -14994
rect 20884 -15054 20890 -14994
rect 20950 -15054 20956 -14994
rect 18352 -15238 21440 -15178
rect 18352 -15340 18412 -15238
rect 21380 -15340 21440 -15238
rect 22418 -15264 22986 -15204
rect 22418 -15340 22478 -15264
rect 18132 -15346 18620 -15340
rect 18132 -15380 18144 -15346
rect 18608 -15380 18620 -15346
rect 18132 -15386 18620 -15380
rect 19150 -15346 19638 -15340
rect 19150 -15380 19162 -15346
rect 19626 -15380 19638 -15346
rect 19150 -15386 19638 -15380
rect 20168 -15346 20656 -15340
rect 20168 -15380 20180 -15346
rect 20644 -15380 20656 -15346
rect 20168 -15386 20656 -15380
rect 21186 -15346 21674 -15340
rect 21186 -15380 21198 -15346
rect 21662 -15380 21674 -15346
rect 21186 -15386 21674 -15380
rect 22204 -15346 22692 -15340
rect 22204 -15380 22216 -15346
rect 22680 -15380 22692 -15346
rect 22204 -15386 22692 -15380
rect 17838 -15488 17850 -15430
rect 17844 -15960 17850 -15488
rect 16866 -16006 16876 -15970
rect 16096 -16056 16584 -16050
rect 16096 -16090 16108 -16056
rect 16572 -16090 16584 -16056
rect 16096 -16096 16584 -16090
rect 15794 -16194 15800 -16134
rect 15860 -16194 15866 -16134
rect 14972 -16520 14978 -16460
rect 15038 -16520 15044 -16460
rect 15266 -16518 15272 -16458
rect 15332 -16518 15338 -16458
rect 15272 -16574 15332 -16518
rect 15078 -16580 15566 -16574
rect 15078 -16614 15090 -16580
rect 15554 -16614 15566 -16580
rect 15078 -16620 15566 -16614
rect 13812 -17194 13818 -16702
rect 14782 -16708 14796 -16664
rect 13812 -17240 13826 -17194
rect 7952 -17290 8440 -17284
rect 7952 -17324 7964 -17290
rect 8428 -17324 8440 -17290
rect 7952 -17330 8440 -17324
rect 8970 -17290 9458 -17284
rect 8970 -17324 8982 -17290
rect 9446 -17324 9458 -17290
rect 8970 -17330 9458 -17324
rect 9988 -17290 10476 -17284
rect 9988 -17324 10000 -17290
rect 10464 -17324 10476 -17290
rect 9988 -17330 10476 -17324
rect 11006 -17290 11494 -17284
rect 11006 -17324 11018 -17290
rect 11482 -17324 11494 -17290
rect 11006 -17330 11494 -17324
rect 12024 -17290 12512 -17284
rect 12024 -17324 12036 -17290
rect 12500 -17324 12512 -17290
rect 12024 -17330 12238 -17324
rect 12240 -17330 12512 -17324
rect 13042 -17290 13530 -17284
rect 13042 -17324 13054 -17290
rect 13518 -17324 13530 -17290
rect 13042 -17330 13264 -17324
rect 13268 -17330 13530 -17324
rect 7652 -17450 7658 -17390
rect 7718 -17450 7724 -17390
rect 4598 -17754 4604 -17694
rect 4664 -17754 4670 -17694
rect 3880 -17812 4368 -17806
rect 3880 -17846 3892 -17812
rect 4356 -17846 4368 -17812
rect 3880 -17852 4368 -17846
rect 3584 -17934 3598 -17896
rect 2614 -18472 2624 -18426
rect 3592 -18430 3598 -17934
rect 2564 -18634 2624 -18472
rect 3582 -18472 3598 -18430
rect 3632 -17934 3644 -17896
rect 4604 -17896 4664 -17754
rect 4898 -17812 5386 -17806
rect 4898 -17846 4910 -17812
rect 5374 -17846 5386 -17812
rect 4898 -17852 5386 -17846
rect 3632 -18430 3638 -17934
rect 4604 -17936 4616 -17896
rect 3632 -18472 3642 -18430
rect 2862 -18522 3350 -18516
rect 2862 -18556 2874 -18522
rect 3338 -18556 3350 -18522
rect 2862 -18562 3350 -18556
rect 3076 -18634 3136 -18562
rect 3582 -18634 3642 -18472
rect 4610 -18472 4616 -17936
rect 4650 -17936 4664 -17896
rect 5620 -17896 5680 -17654
rect 6122 -17660 6128 -17600
rect 6188 -17660 6194 -17600
rect 7144 -17660 7150 -17600
rect 7210 -17660 7216 -17600
rect 6632 -17754 6638 -17694
rect 6698 -17754 6704 -17694
rect 5916 -17812 6404 -17806
rect 5916 -17846 5928 -17812
rect 6392 -17846 6404 -17812
rect 5916 -17852 6404 -17846
rect 4650 -18472 4656 -17936
rect 5620 -17948 5634 -17896
rect 4610 -18484 4656 -18472
rect 5628 -18472 5634 -17948
rect 5668 -17948 5680 -17896
rect 6638 -17896 6698 -17754
rect 7150 -17806 7210 -17660
rect 6934 -17812 7422 -17806
rect 6934 -17846 6946 -17812
rect 7410 -17846 7422 -17812
rect 6934 -17852 7422 -17846
rect 6638 -17940 6652 -17896
rect 5668 -18472 5674 -17948
rect 6646 -18436 6652 -17940
rect 5628 -18484 5674 -18472
rect 6638 -18472 6652 -18436
rect 6686 -17940 6698 -17896
rect 7658 -17896 7718 -17450
rect 8164 -17600 8224 -17330
rect 9182 -17492 9242 -17330
rect 10202 -17380 10262 -17330
rect 11202 -17380 11262 -17330
rect 12240 -17380 12300 -17330
rect 13268 -17380 13328 -17330
rect 9684 -17450 9690 -17390
rect 9750 -17450 9756 -17390
rect 10202 -17440 13328 -17380
rect 9176 -17552 9182 -17492
rect 9242 -17552 9248 -17492
rect 8158 -17660 8164 -17600
rect 8224 -17660 8230 -17600
rect 9176 -17660 9182 -17600
rect 9242 -17660 9248 -17600
rect 8164 -17806 8224 -17660
rect 8668 -17754 8674 -17694
rect 8734 -17754 8740 -17694
rect 7952 -17812 8440 -17806
rect 7952 -17846 7964 -17812
rect 8428 -17846 8440 -17812
rect 7952 -17852 8440 -17846
rect 6686 -18436 6692 -17940
rect 6686 -18472 6698 -18436
rect 3880 -18522 4368 -18516
rect 3880 -18556 3892 -18522
rect 4356 -18556 4368 -18522
rect 3880 -18562 4368 -18556
rect 4898 -18522 5386 -18516
rect 4898 -18556 4910 -18522
rect 5374 -18556 5386 -18522
rect 4898 -18562 5386 -18556
rect 5916 -18522 6404 -18516
rect 5916 -18556 5928 -18522
rect 6392 -18556 6404 -18522
rect 5916 -18562 6404 -18556
rect 4086 -18618 4146 -18562
rect 2564 -18694 3642 -18634
rect 4080 -18678 4086 -18618
rect 4146 -18678 4152 -18618
rect 4990 -18678 4996 -18618
rect 5056 -18678 5062 -18618
rect 4080 -18894 4086 -18834
rect 4146 -18894 4152 -18834
rect 4086 -18900 4148 -18894
rect 2448 -18938 2510 -18932
rect 2448 -18998 2450 -18938
rect 2448 -19004 2510 -18998
rect 2330 -20256 2336 -20196
rect 2396 -20256 2402 -20196
rect 2230 -21260 2294 -21254
rect 2230 -21312 2242 -21260
rect 2230 -21318 2294 -21312
rect 2230 -22440 2290 -21318
rect 2336 -22314 2396 -20256
rect 2448 -21182 2508 -19004
rect 4088 -19040 4148 -18900
rect 4996 -19040 5056 -18678
rect 5124 -18834 5184 -18562
rect 5992 -18678 5998 -18618
rect 6058 -18678 6064 -18618
rect 5124 -18900 5184 -18894
rect 5998 -19040 6058 -18678
rect 6138 -18834 6198 -18562
rect 6638 -18720 6698 -18472
rect 7658 -18472 7670 -17896
rect 7704 -18472 7718 -17896
rect 8674 -17896 8734 -17754
rect 9182 -17806 9242 -17660
rect 8970 -17812 9458 -17806
rect 8970 -17846 8982 -17812
rect 9446 -17846 9458 -17812
rect 8970 -17852 9458 -17846
rect 8674 -17932 8688 -17896
rect 6934 -18522 7422 -18516
rect 6934 -18556 6946 -18522
rect 7410 -18556 7422 -18522
rect 6934 -18562 7126 -18556
rect 7150 -18562 7422 -18556
rect 7150 -18618 7210 -18562
rect 7144 -18678 7150 -18618
rect 7210 -18678 7216 -18618
rect 6632 -18780 6638 -18720
rect 6698 -18780 6704 -18720
rect 6132 -18894 6138 -18834
rect 6198 -18894 6204 -18834
rect 7150 -19040 7210 -18678
rect 2862 -19046 3350 -19040
rect 2862 -19080 2874 -19046
rect 3338 -19080 3350 -19046
rect 2862 -19086 3350 -19080
rect 3880 -19046 4368 -19040
rect 3880 -19080 3892 -19046
rect 4356 -19080 4368 -19046
rect 3880 -19086 4368 -19080
rect 4898 -19046 5386 -19040
rect 4898 -19080 4910 -19046
rect 5374 -19080 5386 -19046
rect 4898 -19086 5386 -19080
rect 5916 -19046 6404 -19040
rect 5916 -19080 5928 -19046
rect 6392 -19080 6404 -19046
rect 5916 -19086 6404 -19080
rect 6934 -19046 7422 -19040
rect 6934 -19080 6946 -19046
rect 7410 -19080 7422 -19046
rect 6934 -19086 7422 -19080
rect 2574 -19130 2620 -19118
rect 2574 -19668 2580 -19130
rect 2568 -19706 2580 -19668
rect 2614 -19668 2620 -19130
rect 3592 -19130 3638 -19118
rect 3592 -19668 3598 -19130
rect 2614 -19706 2628 -19668
rect 2568 -19836 2628 -19706
rect 3586 -19706 3598 -19668
rect 3632 -19668 3638 -19130
rect 4610 -19130 4656 -19118
rect 4610 -19656 4616 -19130
rect 3632 -19706 3646 -19668
rect 2862 -19756 3350 -19750
rect 2862 -19790 2874 -19756
rect 3338 -19790 3350 -19756
rect 2862 -19796 3350 -19790
rect 3066 -19836 3126 -19796
rect 3586 -19836 3646 -19706
rect 4602 -19706 4616 -19656
rect 4650 -19656 4656 -19130
rect 5628 -19130 5674 -19118
rect 5628 -19648 5634 -19130
rect 4650 -19706 4662 -19656
rect 3880 -19756 4368 -19750
rect 3880 -19790 3892 -19756
rect 4356 -19790 4368 -19756
rect 3880 -19796 4368 -19790
rect 2568 -19896 3646 -19836
rect 3586 -19950 3646 -19896
rect 4078 -19906 4084 -19846
rect 4144 -19906 4150 -19846
rect 3580 -20010 3586 -19950
rect 3646 -20010 3652 -19950
rect 3576 -20220 3582 -20160
rect 3642 -20220 3648 -20160
rect 2862 -20280 3350 -20274
rect 2862 -20314 2874 -20280
rect 3338 -20314 3350 -20280
rect 2862 -20320 3350 -20314
rect 2574 -20364 2620 -20352
rect 2574 -20906 2580 -20364
rect 2564 -20940 2580 -20906
rect 2614 -20906 2620 -20364
rect 3582 -20364 3642 -20220
rect 4084 -20274 4144 -19906
rect 4602 -20062 4662 -19706
rect 5620 -19706 5634 -19648
rect 5668 -19648 5674 -19130
rect 6646 -19130 6692 -19118
rect 5668 -19706 5680 -19648
rect 6646 -19660 6652 -19130
rect 4898 -19756 5386 -19750
rect 4898 -19790 4910 -19756
rect 5374 -19790 5386 -19756
rect 4898 -19796 5386 -19790
rect 5092 -19846 5152 -19796
rect 5086 -19906 5092 -19846
rect 5152 -19906 5158 -19846
rect 4596 -20122 4602 -20062
rect 4662 -20122 4668 -20062
rect 5620 -20160 5680 -19706
rect 6640 -19706 6652 -19660
rect 6686 -19660 6692 -19130
rect 7658 -19130 7718 -18472
rect 8682 -18472 8688 -17932
rect 8722 -17932 8734 -17896
rect 9690 -17896 9750 -17450
rect 10196 -17660 10202 -17600
rect 10262 -17660 10268 -17600
rect 13268 -17616 13328 -17440
rect 13766 -17506 13826 -17240
rect 14790 -17240 14796 -16708
rect 14830 -16708 14842 -16664
rect 15800 -16664 15860 -16194
rect 16302 -16452 16362 -16096
rect 16816 -16350 16876 -16006
rect 17836 -16006 17850 -15960
rect 17884 -15488 17898 -15430
rect 18862 -15430 18908 -15418
rect 17884 -15960 17890 -15488
rect 18862 -15950 18868 -15430
rect 17884 -16006 17896 -15960
rect 17114 -16056 17602 -16050
rect 17114 -16090 17126 -16056
rect 17590 -16090 17602 -16056
rect 17114 -16096 17602 -16090
rect 16810 -16410 16816 -16350
rect 16876 -16410 16882 -16350
rect 16300 -16458 16362 -16452
rect 16360 -16518 16362 -16458
rect 16300 -16524 16362 -16518
rect 16812 -16524 16818 -16464
rect 16878 -16524 16884 -16464
rect 16302 -16574 16362 -16524
rect 16096 -16580 16584 -16574
rect 16096 -16614 16108 -16580
rect 16572 -16614 16584 -16580
rect 16096 -16620 16584 -16614
rect 15800 -16708 15814 -16664
rect 14830 -17240 14836 -16708
rect 14790 -17252 14836 -17240
rect 15808 -17240 15814 -16708
rect 15848 -16708 15860 -16664
rect 16818 -16664 16878 -16524
rect 17326 -16574 17386 -16096
rect 17836 -16134 17896 -16006
rect 18854 -16006 18868 -15950
rect 18902 -15950 18908 -15430
rect 19880 -15430 19926 -15418
rect 18902 -16006 18914 -15950
rect 19880 -15962 19886 -15430
rect 18132 -16056 18620 -16050
rect 18132 -16090 18144 -16056
rect 18608 -16090 18620 -16056
rect 18132 -16096 18620 -16090
rect 17830 -16194 17836 -16134
rect 17896 -16194 17902 -16134
rect 17114 -16580 17602 -16574
rect 17114 -16614 17126 -16580
rect 17590 -16614 17602 -16580
rect 17114 -16620 17602 -16614
rect 16818 -16694 16832 -16664
rect 15848 -17240 15854 -16708
rect 16826 -17200 16832 -16694
rect 15808 -17252 15854 -17240
rect 16818 -17240 16832 -17200
rect 16866 -16694 16878 -16664
rect 17836 -16664 17896 -16194
rect 18352 -16574 18412 -16096
rect 18854 -16350 18914 -16006
rect 19870 -16006 19886 -15962
rect 19920 -15962 19926 -15430
rect 20898 -15430 20944 -15418
rect 20898 -15962 20904 -15430
rect 19920 -16006 19930 -15962
rect 19150 -16056 19638 -16050
rect 19150 -16090 19162 -16056
rect 19626 -16090 19638 -16056
rect 19150 -16096 19638 -16090
rect 18848 -16410 18854 -16350
rect 18914 -16410 18920 -16350
rect 19360 -16400 19420 -16096
rect 19870 -16242 19930 -16006
rect 20894 -16006 20904 -15962
rect 20938 -15962 20944 -15430
rect 21916 -15430 21962 -15418
rect 21916 -15956 21922 -15430
rect 20938 -16006 20954 -15962
rect 20168 -16056 20656 -16050
rect 20168 -16090 20180 -16056
rect 20644 -16090 20656 -16056
rect 20168 -16096 20656 -16090
rect 20376 -16240 20436 -16096
rect 19864 -16302 19870 -16242
rect 19930 -16302 19936 -16242
rect 20374 -16246 20436 -16240
rect 20434 -16306 20436 -16246
rect 20374 -16312 20436 -16306
rect 20376 -16400 20436 -16312
rect 20894 -16350 20954 -16006
rect 21910 -16006 21922 -15956
rect 21956 -15956 21962 -15430
rect 22926 -15430 22986 -15264
rect 23028 -15288 23034 -15228
rect 23094 -15288 23100 -15228
rect 22926 -15458 22940 -15430
rect 22934 -15948 22940 -15458
rect 21956 -16006 21970 -15956
rect 21186 -16056 21674 -16050
rect 21186 -16090 21198 -16056
rect 21662 -16090 21674 -16056
rect 21186 -16096 21674 -16090
rect 19360 -16460 20436 -16400
rect 20888 -16410 20894 -16350
rect 20954 -16410 20960 -16350
rect 18848 -16524 18854 -16464
rect 18914 -16524 18920 -16464
rect 18132 -16580 18620 -16574
rect 18132 -16614 18144 -16580
rect 18608 -16614 18620 -16580
rect 18132 -16620 18620 -16614
rect 16866 -17200 16872 -16694
rect 17836 -16704 17850 -16664
rect 16866 -17240 16878 -17200
rect 17844 -17206 17850 -16704
rect 14060 -17290 14548 -17284
rect 14060 -17324 14072 -17290
rect 14536 -17324 14548 -17290
rect 14060 -17330 14548 -17324
rect 15078 -17290 15566 -17284
rect 15078 -17324 15090 -17290
rect 15554 -17324 15566 -17290
rect 15078 -17330 15566 -17324
rect 16096 -17290 16584 -17284
rect 16096 -17324 16108 -17290
rect 16572 -17324 16584 -17290
rect 16096 -17330 16584 -17324
rect 14272 -17378 14332 -17330
rect 13760 -17566 13766 -17506
rect 13826 -17566 13832 -17506
rect 14272 -17616 14332 -17438
rect 10202 -17806 10262 -17660
rect 13268 -17676 14332 -17616
rect 15796 -17764 15802 -17704
rect 15862 -17764 15868 -17704
rect 9988 -17812 10476 -17806
rect 9988 -17846 10000 -17812
rect 10464 -17846 10476 -17812
rect 9988 -17852 10476 -17846
rect 11006 -17812 11494 -17806
rect 11006 -17846 11018 -17812
rect 11482 -17846 11494 -17812
rect 11006 -17852 11494 -17846
rect 12024 -17812 12512 -17806
rect 12024 -17846 12036 -17812
rect 12500 -17846 12512 -17812
rect 12024 -17852 12512 -17846
rect 13042 -17812 13530 -17806
rect 13042 -17846 13054 -17812
rect 13518 -17846 13530 -17812
rect 13042 -17852 13530 -17846
rect 14060 -17812 14548 -17806
rect 14060 -17846 14072 -17812
rect 14536 -17846 14548 -17812
rect 14060 -17852 14548 -17846
rect 15078 -17812 15566 -17806
rect 15078 -17846 15090 -17812
rect 15554 -17846 15566 -17812
rect 15078 -17852 15566 -17846
rect 8722 -18472 8728 -17932
rect 9690 -17934 9706 -17896
rect 8682 -18484 8728 -18472
rect 9700 -18472 9706 -17934
rect 9740 -17934 9750 -17896
rect 10718 -17896 10764 -17884
rect 9740 -18472 9746 -17934
rect 10718 -18430 10724 -17896
rect 9700 -18484 9746 -18472
rect 10710 -18472 10724 -18430
rect 10758 -18430 10764 -17896
rect 11736 -17896 11782 -17884
rect 10758 -18472 10770 -18430
rect 11736 -18434 11742 -17896
rect 7952 -18522 8440 -18516
rect 7952 -18556 7964 -18522
rect 8428 -18556 8440 -18522
rect 7952 -18562 8220 -18556
rect 8224 -18562 8440 -18556
rect 8970 -18522 9458 -18516
rect 8970 -18556 8982 -18522
rect 9446 -18556 9458 -18522
rect 8970 -18562 9458 -18556
rect 9988 -18522 10476 -18516
rect 9988 -18556 10000 -18522
rect 10464 -18556 10476 -18522
rect 9988 -18562 10476 -18556
rect 8160 -18618 8220 -18562
rect 9166 -18618 9226 -18562
rect 10210 -18618 10270 -18562
rect 10710 -18612 10770 -18472
rect 11730 -18472 11742 -18434
rect 11776 -18434 11782 -17896
rect 12754 -17896 12800 -17884
rect 11776 -18472 11790 -18434
rect 12754 -18440 12760 -17896
rect 11006 -18522 11494 -18516
rect 11006 -18556 11018 -18522
rect 11482 -18556 11494 -18522
rect 11006 -18562 11494 -18556
rect 8154 -18678 8160 -18618
rect 8220 -18678 8226 -18618
rect 9160 -18678 9166 -18618
rect 9226 -18678 9232 -18618
rect 10204 -18678 10210 -18618
rect 10270 -18678 10276 -18618
rect 10704 -18672 10710 -18612
rect 10770 -18672 10776 -18612
rect 8160 -19040 8220 -18678
rect 9158 -18894 9164 -18834
rect 9224 -18894 9230 -18834
rect 10198 -18894 10204 -18834
rect 10264 -18894 10270 -18834
rect 9164 -19040 9224 -18894
rect 9682 -18998 9688 -18938
rect 9748 -18998 9754 -18938
rect 7952 -19046 8440 -19040
rect 7952 -19080 7964 -19046
rect 8428 -19080 8440 -19046
rect 7952 -19086 8440 -19080
rect 8970 -19046 9458 -19040
rect 8970 -19080 8982 -19046
rect 9446 -19080 9458 -19046
rect 8970 -19086 9458 -19080
rect 7658 -19212 7670 -19130
rect 7664 -19660 7670 -19212
rect 6686 -19706 6700 -19660
rect 5916 -19756 6404 -19750
rect 5916 -19790 5928 -19756
rect 6392 -19790 6404 -19756
rect 5916 -19796 6404 -19790
rect 6106 -19846 6166 -19796
rect 6100 -19906 6106 -19846
rect 6166 -19906 6172 -19846
rect 6640 -20062 6700 -19706
rect 7660 -19706 7670 -19660
rect 7704 -19212 7718 -19130
rect 8682 -19130 8728 -19118
rect 7704 -19660 7710 -19212
rect 7704 -19706 7720 -19660
rect 8682 -19662 8688 -19130
rect 6934 -19756 7422 -19750
rect 6934 -19790 6946 -19756
rect 7410 -19790 7422 -19756
rect 6934 -19796 7422 -19790
rect 7144 -19846 7204 -19796
rect 7138 -19906 7144 -19846
rect 7204 -19906 7210 -19846
rect 6634 -20122 6640 -20062
rect 6700 -20122 6706 -20062
rect 5614 -20220 5620 -20160
rect 5680 -20220 5686 -20160
rect 7144 -20274 7204 -19906
rect 7660 -20160 7720 -19706
rect 8678 -19706 8688 -19662
rect 8722 -19662 8728 -19130
rect 9688 -19130 9748 -18998
rect 10204 -19040 10264 -18894
rect 9988 -19046 10476 -19040
rect 9988 -19080 10000 -19046
rect 10464 -19080 10476 -19046
rect 9988 -19086 10476 -19080
rect 9688 -19194 9706 -19130
rect 8722 -19706 8738 -19662
rect 7952 -19756 8440 -19750
rect 7952 -19790 7964 -19756
rect 8428 -19790 8440 -19756
rect 7952 -19796 8222 -19790
rect 8230 -19796 8440 -19790
rect 8162 -19846 8222 -19796
rect 8678 -19840 8738 -19706
rect 9700 -19706 9706 -19194
rect 9740 -19194 9748 -19130
rect 10710 -19130 10770 -18672
rect 11218 -18834 11278 -18562
rect 11212 -18894 11218 -18834
rect 11278 -18894 11284 -18834
rect 11218 -19040 11278 -18894
rect 11730 -18938 11790 -18472
rect 12746 -18472 12760 -18440
rect 12794 -18440 12800 -17896
rect 13772 -17896 13818 -17884
rect 13772 -18438 13778 -17896
rect 12794 -18472 12806 -18440
rect 12024 -18522 12512 -18516
rect 12024 -18556 12036 -18522
rect 12500 -18556 12512 -18522
rect 12024 -18562 12512 -18556
rect 12226 -18834 12286 -18562
rect 12746 -18612 12806 -18472
rect 13768 -18472 13778 -18438
rect 13812 -18438 13818 -17896
rect 14790 -17896 14836 -17884
rect 13812 -18472 13828 -18438
rect 14790 -18440 14796 -17896
rect 13042 -18522 13530 -18516
rect 13042 -18556 13054 -18522
rect 13518 -18556 13530 -18522
rect 13042 -18562 13530 -18556
rect 12740 -18672 12746 -18612
rect 12806 -18672 12812 -18612
rect 13270 -18834 13330 -18562
rect 12220 -18894 12226 -18834
rect 12286 -18894 12292 -18834
rect 13264 -18894 13270 -18834
rect 13330 -18894 13336 -18834
rect 11724 -18998 11730 -18938
rect 11790 -18998 11796 -18938
rect 11006 -19046 11494 -19040
rect 11006 -19080 11018 -19046
rect 11482 -19080 11494 -19046
rect 11006 -19086 11494 -19080
rect 10710 -19166 10724 -19130
rect 9740 -19706 9746 -19194
rect 10718 -19648 10724 -19166
rect 9700 -19718 9746 -19706
rect 10714 -19706 10724 -19648
rect 10758 -19166 10770 -19130
rect 11730 -19130 11790 -18998
rect 12226 -19040 12286 -18894
rect 13270 -19040 13330 -18894
rect 13768 -18938 13828 -18472
rect 14782 -18472 14796 -18440
rect 14830 -18440 14836 -17896
rect 15802 -17896 15862 -17764
rect 16096 -17812 16584 -17806
rect 16096 -17846 16108 -17812
rect 16572 -17846 16584 -17812
rect 16096 -17852 16584 -17846
rect 14830 -18472 14842 -18440
rect 14060 -18522 14548 -18516
rect 14060 -18556 14072 -18522
rect 14536 -18556 14548 -18522
rect 14060 -18562 14548 -18556
rect 14260 -18834 14320 -18562
rect 14782 -18612 14842 -18472
rect 15802 -18472 15814 -17896
rect 15848 -18472 15862 -17896
rect 16818 -17896 16878 -17240
rect 17838 -17240 17850 -17206
rect 17884 -16704 17896 -16664
rect 18854 -16664 18914 -16524
rect 19360 -16574 19420 -16460
rect 20376 -16574 20436 -16460
rect 20886 -16524 20892 -16464
rect 20952 -16524 20958 -16464
rect 19150 -16580 19638 -16574
rect 19150 -16614 19162 -16580
rect 19626 -16614 19638 -16580
rect 19150 -16620 19638 -16614
rect 20168 -16580 20656 -16574
rect 20168 -16614 20180 -16580
rect 20644 -16614 20656 -16580
rect 20168 -16620 20656 -16614
rect 17884 -17206 17890 -16704
rect 18854 -16706 18868 -16664
rect 17884 -17240 17898 -17206
rect 17114 -17290 17602 -17284
rect 17114 -17324 17126 -17290
rect 17590 -17324 17602 -17290
rect 17114 -17330 17602 -17324
rect 17314 -17600 17374 -17330
rect 17308 -17660 17314 -17600
rect 17374 -17660 17380 -17600
rect 17314 -17806 17374 -17660
rect 17114 -17812 17602 -17806
rect 17114 -17846 17126 -17812
rect 17590 -17846 17602 -17812
rect 17114 -17852 17602 -17846
rect 16818 -17936 16832 -17896
rect 16826 -18440 16832 -17936
rect 15078 -18522 15566 -18516
rect 15078 -18556 15090 -18522
rect 15554 -18556 15566 -18522
rect 15078 -18562 15566 -18556
rect 14776 -18672 14782 -18612
rect 14842 -18672 14848 -18612
rect 15278 -18834 15338 -18562
rect 14254 -18894 14260 -18834
rect 14320 -18894 14326 -18834
rect 15272 -18894 15278 -18834
rect 15338 -18894 15344 -18834
rect 13762 -18998 13768 -18938
rect 13828 -18998 13834 -18938
rect 12024 -19046 12512 -19040
rect 12024 -19080 12036 -19046
rect 12500 -19080 12512 -19046
rect 12024 -19086 12512 -19080
rect 13042 -19046 13530 -19040
rect 13042 -19080 13054 -19046
rect 13518 -19080 13530 -19046
rect 13042 -19086 13530 -19080
rect 10758 -19648 10764 -19166
rect 11730 -19168 11742 -19130
rect 10758 -19706 10774 -19648
rect 8970 -19756 9458 -19750
rect 8970 -19790 8982 -19756
rect 9446 -19790 9458 -19756
rect 8970 -19796 9458 -19790
rect 9988 -19756 10476 -19750
rect 9988 -19790 10000 -19756
rect 10464 -19790 10476 -19756
rect 9988 -19796 10476 -19790
rect 10714 -19840 10774 -19706
rect 11736 -19706 11742 -19168
rect 11776 -19168 11790 -19130
rect 12754 -19130 12800 -19118
rect 11776 -19706 11782 -19168
rect 12754 -19656 12760 -19130
rect 11736 -19718 11782 -19706
rect 12746 -19706 12760 -19656
rect 12794 -19656 12800 -19130
rect 13768 -19130 13828 -18998
rect 14260 -19040 14320 -18894
rect 15802 -18938 15862 -18472
rect 16820 -18472 16832 -18440
rect 16866 -17936 16878 -17896
rect 17838 -17896 17898 -17240
rect 18862 -17240 18868 -16706
rect 18902 -16706 18914 -16664
rect 19880 -16664 19926 -16652
rect 18902 -17240 18908 -16706
rect 19880 -17182 19886 -16664
rect 18862 -17252 18908 -17240
rect 19872 -17240 19886 -17182
rect 19920 -17182 19926 -16664
rect 20892 -16664 20952 -16524
rect 21394 -16574 21454 -16096
rect 21910 -16134 21970 -16006
rect 22928 -16006 22940 -15948
rect 22974 -15458 22986 -15430
rect 22974 -15948 22980 -15458
rect 22974 -16006 22988 -15948
rect 22204 -16056 22692 -16050
rect 22204 -16090 22216 -16056
rect 22680 -16090 22692 -16056
rect 22204 -16096 22692 -16090
rect 22928 -16116 22988 -16006
rect 21904 -16194 21910 -16134
rect 21970 -16194 21976 -16134
rect 22922 -16176 22928 -16116
rect 22988 -16176 22994 -16116
rect 21910 -16412 21970 -16194
rect 21910 -16472 22984 -16412
rect 23034 -16464 23094 -15288
rect 23522 -16306 23528 -16246
rect 23588 -16306 23594 -16246
rect 23272 -16410 23278 -16350
rect 23338 -16410 23344 -16350
rect 21186 -16580 21674 -16574
rect 21186 -16614 21198 -16580
rect 21662 -16614 21674 -16580
rect 21186 -16620 21674 -16614
rect 20892 -16706 20904 -16664
rect 19920 -17240 19932 -17182
rect 18344 -17284 18404 -17282
rect 18132 -17290 18620 -17284
rect 18132 -17324 18144 -17290
rect 18608 -17324 18620 -17290
rect 18132 -17330 18620 -17324
rect 19150 -17290 19638 -17284
rect 19150 -17324 19162 -17290
rect 19626 -17324 19638 -17290
rect 19150 -17330 19638 -17324
rect 18344 -17600 18404 -17330
rect 19366 -17378 19426 -17330
rect 19360 -17438 19366 -17378
rect 19426 -17438 19432 -17378
rect 19498 -17434 19504 -17374
rect 19564 -17434 19570 -17374
rect 19504 -17600 19564 -17434
rect 19872 -17600 19932 -17240
rect 20898 -17240 20904 -16706
rect 20938 -16706 20952 -16664
rect 21910 -16664 21970 -16472
rect 22414 -16574 22474 -16472
rect 22204 -16580 22692 -16574
rect 22204 -16614 22216 -16580
rect 22680 -16614 22692 -16580
rect 22204 -16620 22692 -16614
rect 21910 -16698 21922 -16664
rect 20938 -17240 20944 -16706
rect 21916 -17200 21922 -16698
rect 20898 -17252 20944 -17240
rect 21910 -17240 21922 -17200
rect 21956 -16698 21970 -16664
rect 22924 -16664 22984 -16472
rect 23028 -16524 23034 -16464
rect 23094 -16524 23100 -16464
rect 22924 -16688 22940 -16664
rect 21956 -17200 21962 -16698
rect 21956 -17240 21970 -17200
rect 20168 -17290 20656 -17284
rect 20168 -17324 20180 -17290
rect 20644 -17324 20656 -17290
rect 20168 -17330 20656 -17324
rect 21186 -17290 21674 -17284
rect 21186 -17324 21198 -17290
rect 21392 -17324 21452 -17294
rect 21662 -17324 21674 -17290
rect 21186 -17330 21674 -17324
rect 21392 -17374 21452 -17330
rect 20380 -17434 20386 -17374
rect 20446 -17434 20452 -17374
rect 21386 -17434 21392 -17374
rect 21452 -17434 21458 -17374
rect 21910 -17378 21970 -17240
rect 22934 -17240 22940 -16688
rect 22974 -16688 22984 -16664
rect 22974 -17240 22980 -16688
rect 22934 -17252 22980 -17240
rect 22204 -17290 22692 -17284
rect 22204 -17324 22216 -17290
rect 22680 -17324 22692 -17290
rect 22204 -17330 22692 -17324
rect 18338 -17660 18344 -17600
rect 18404 -17660 18410 -17600
rect 19498 -17660 19504 -17600
rect 19564 -17660 19570 -17600
rect 19866 -17660 19872 -17600
rect 19932 -17660 19938 -17600
rect 18344 -17806 18404 -17660
rect 19504 -17806 19564 -17660
rect 19872 -17704 19932 -17660
rect 19866 -17764 19872 -17704
rect 19932 -17764 19938 -17704
rect 20386 -17806 20446 -17434
rect 21904 -17438 21910 -17378
rect 21970 -17438 21976 -17378
rect 21904 -17566 21910 -17506
rect 21970 -17566 21976 -17506
rect 20882 -17762 20888 -17702
rect 20948 -17762 20954 -17702
rect 18132 -17812 18620 -17806
rect 18132 -17846 18144 -17812
rect 18608 -17846 18620 -17812
rect 18132 -17852 18620 -17846
rect 19150 -17812 19638 -17806
rect 19150 -17846 19162 -17812
rect 19626 -17846 19638 -17812
rect 19150 -17852 19638 -17846
rect 20168 -17812 20656 -17806
rect 20168 -17846 20180 -17812
rect 20644 -17846 20656 -17812
rect 20168 -17852 20656 -17846
rect 20386 -17854 20446 -17852
rect 16866 -18440 16872 -17936
rect 17838 -17942 17850 -17896
rect 17844 -18428 17850 -17942
rect 16866 -18472 16880 -18440
rect 16096 -18522 16584 -18516
rect 16096 -18556 16108 -18522
rect 16572 -18556 16584 -18522
rect 16096 -18562 16584 -18556
rect 16312 -18834 16372 -18562
rect 16820 -18612 16880 -18472
rect 17836 -18472 17850 -18428
rect 17884 -17942 17898 -17896
rect 18862 -17896 18908 -17884
rect 17884 -18428 17890 -17942
rect 17884 -18472 17896 -18428
rect 18862 -18432 18868 -17896
rect 17114 -18522 17602 -18516
rect 17114 -18556 17126 -18522
rect 17590 -18556 17602 -18522
rect 17114 -18562 17602 -18556
rect 16814 -18672 16820 -18612
rect 16880 -18672 16886 -18612
rect 16806 -18780 16812 -18720
rect 16872 -18780 16878 -18720
rect 16306 -18894 16312 -18834
rect 16372 -18894 16378 -18834
rect 15796 -18998 15802 -18938
rect 15862 -18998 15868 -18938
rect 16308 -19002 16314 -18942
rect 16374 -19002 16380 -18942
rect 16314 -19040 16374 -19002
rect 14060 -19046 14548 -19040
rect 14060 -19080 14072 -19046
rect 14536 -19080 14548 -19046
rect 14060 -19086 14548 -19080
rect 15078 -19046 15566 -19040
rect 15078 -19080 15090 -19046
rect 15554 -19080 15566 -19046
rect 15078 -19086 15566 -19080
rect 16096 -19046 16584 -19040
rect 16096 -19080 16108 -19046
rect 16572 -19080 16584 -19046
rect 16096 -19086 16584 -19080
rect 13768 -19166 13778 -19130
rect 12794 -19706 12806 -19656
rect 11006 -19756 11494 -19750
rect 11006 -19790 11018 -19756
rect 11482 -19790 11494 -19756
rect 11006 -19796 11494 -19790
rect 12024 -19756 12512 -19750
rect 12024 -19790 12036 -19756
rect 12500 -19790 12512 -19756
rect 12024 -19796 12512 -19790
rect 12746 -19840 12806 -19706
rect 13772 -19706 13778 -19166
rect 13812 -19166 13828 -19130
rect 14790 -19130 14836 -19118
rect 13812 -19706 13818 -19166
rect 14790 -19644 14796 -19130
rect 13772 -19718 13818 -19706
rect 14780 -19706 14796 -19644
rect 14830 -19644 14836 -19130
rect 15808 -19130 15854 -19118
rect 14830 -19706 14840 -19644
rect 15808 -19664 15814 -19130
rect 13042 -19756 13530 -19750
rect 13042 -19790 13054 -19756
rect 13518 -19790 13530 -19756
rect 13042 -19796 13530 -19790
rect 14060 -19756 14548 -19750
rect 14060 -19790 14072 -19756
rect 14536 -19790 14548 -19756
rect 14060 -19796 14548 -19790
rect 14780 -19840 14840 -19706
rect 15802 -19706 15814 -19664
rect 15848 -19664 15854 -19130
rect 16812 -19130 16872 -18780
rect 17336 -18942 17396 -18562
rect 17836 -18936 17896 -18472
rect 18856 -18472 18868 -18432
rect 18902 -18432 18908 -17896
rect 19880 -17896 19926 -17884
rect 19880 -18428 19886 -17896
rect 18902 -18472 18916 -18432
rect 18132 -18522 18620 -18516
rect 18132 -18556 18144 -18522
rect 18608 -18556 18620 -18522
rect 18132 -18562 18620 -18556
rect 17330 -19002 17336 -18942
rect 17396 -19002 17402 -18942
rect 17830 -18996 17836 -18936
rect 17896 -18996 17902 -18936
rect 17336 -19040 17396 -19002
rect 17114 -19046 17602 -19040
rect 17114 -19080 17126 -19046
rect 17590 -19080 17602 -19046
rect 17114 -19086 17602 -19080
rect 16812 -19166 16832 -19130
rect 15848 -19706 15862 -19664
rect 15078 -19756 15566 -19750
rect 15078 -19790 15090 -19756
rect 15554 -19790 15566 -19756
rect 15078 -19796 15566 -19790
rect 8156 -19906 8162 -19846
rect 8222 -19906 8228 -19846
rect 8672 -19900 8678 -19840
rect 8738 -19900 8744 -19840
rect 12740 -19900 12746 -19840
rect 12806 -19900 12812 -19840
rect 14774 -19900 14780 -19840
rect 14840 -19900 14846 -19840
rect 7654 -20220 7660 -20160
rect 7720 -20220 7726 -20160
rect 3880 -20280 4368 -20274
rect 3880 -20314 3892 -20280
rect 4356 -20314 4368 -20280
rect 3880 -20320 4368 -20314
rect 4898 -20280 5386 -20274
rect 4898 -20314 4910 -20280
rect 5374 -20314 5386 -20280
rect 4898 -20320 5386 -20314
rect 5916 -20280 6404 -20274
rect 5916 -20314 5928 -20280
rect 6392 -20314 6404 -20280
rect 5916 -20320 6404 -20314
rect 6934 -20280 7422 -20274
rect 6934 -20314 6946 -20280
rect 7410 -20314 7422 -20280
rect 6934 -20320 7422 -20314
rect 3582 -20418 3598 -20364
rect 2614 -20940 2624 -20906
rect 3592 -20910 3598 -20418
rect 2564 -21072 2624 -20940
rect 3588 -20940 3598 -20910
rect 3632 -20418 3642 -20364
rect 4610 -20364 4656 -20352
rect 3632 -20910 3638 -20418
rect 4610 -20894 4616 -20364
rect 3632 -20940 3648 -20910
rect 2862 -20990 3350 -20984
rect 2862 -21024 2874 -20990
rect 3338 -21024 3350 -20990
rect 2862 -21030 3350 -21024
rect 3084 -21072 3144 -21030
rect 3588 -21072 3648 -20940
rect 4602 -20940 4616 -20894
rect 4650 -20894 4656 -20364
rect 5628 -20364 5674 -20352
rect 4650 -20940 4662 -20894
rect 5628 -20910 5634 -20364
rect 3880 -20990 4368 -20984
rect 3880 -21024 3892 -20990
rect 4356 -21024 4368 -20990
rect 3880 -21030 4368 -21024
rect 2564 -21132 3648 -21072
rect 2442 -21242 2448 -21182
rect 2508 -21242 2514 -21182
rect 3588 -21278 3648 -21132
rect 2564 -21338 3648 -21278
rect 2564 -21596 2624 -21338
rect 3076 -21506 3136 -21338
rect 3588 -21398 3648 -21338
rect 3582 -21458 3588 -21398
rect 3648 -21458 3654 -21398
rect 2862 -21512 3350 -21506
rect 2862 -21546 2874 -21512
rect 3338 -21546 3350 -21512
rect 2862 -21552 3350 -21546
rect 2564 -21632 2580 -21596
rect 2574 -22172 2580 -21632
rect 2614 -21632 2624 -21596
rect 3588 -21596 3648 -21458
rect 4080 -21506 4140 -21030
rect 4602 -21084 4662 -20940
rect 5620 -20940 5634 -20910
rect 5668 -20910 5674 -20364
rect 6646 -20364 6692 -20352
rect 6646 -20898 6652 -20364
rect 5668 -20940 5680 -20910
rect 4898 -20990 5386 -20984
rect 4898 -21024 4910 -20990
rect 5374 -21024 5386 -20990
rect 4898 -21030 5386 -21024
rect 4596 -21144 4602 -21084
rect 4662 -21144 4668 -21084
rect 4600 -21338 4606 -21278
rect 4666 -21338 4672 -21278
rect 3880 -21512 4368 -21506
rect 3880 -21546 3892 -21512
rect 4356 -21546 4368 -21512
rect 3880 -21552 4368 -21546
rect 2614 -22172 2620 -21632
rect 3588 -21636 3598 -21596
rect 2574 -22184 2620 -22172
rect 3592 -22172 3598 -21636
rect 3632 -21636 3648 -21596
rect 4606 -21596 4666 -21338
rect 5100 -21342 5160 -21030
rect 5620 -21182 5680 -20940
rect 6638 -20940 6652 -20898
rect 6686 -20898 6692 -20364
rect 7660 -20364 7720 -20220
rect 8162 -20274 8222 -19906
rect 7952 -20280 8440 -20274
rect 7952 -20314 7964 -20280
rect 8428 -20314 8440 -20280
rect 7952 -20320 8440 -20314
rect 7660 -20394 7670 -20364
rect 7664 -20876 7670 -20394
rect 6686 -20940 6698 -20898
rect 5916 -20990 6404 -20984
rect 5916 -21024 5928 -20990
rect 6392 -21024 6404 -20990
rect 5916 -21030 6404 -21024
rect 5614 -21242 5620 -21182
rect 5680 -21242 5686 -21182
rect 6134 -21342 6194 -21030
rect 6638 -21084 6698 -20940
rect 7656 -20940 7670 -20876
rect 7704 -20394 7720 -20364
rect 8678 -20364 8738 -19900
rect 10714 -19906 10774 -19900
rect 11724 -20010 11730 -19950
rect 11790 -20010 11796 -19950
rect 13760 -20010 13766 -19950
rect 13826 -20010 13832 -19950
rect 10706 -20122 10712 -20062
rect 10772 -20122 10778 -20062
rect 9690 -20220 9696 -20160
rect 9756 -20220 9762 -20160
rect 8970 -20280 9458 -20274
rect 8970 -20314 8982 -20280
rect 9446 -20314 9458 -20280
rect 8970 -20320 9458 -20314
rect 7704 -20876 7710 -20394
rect 8678 -20406 8688 -20364
rect 7704 -20940 7716 -20876
rect 8682 -20900 8688 -20406
rect 6934 -20990 7422 -20984
rect 6934 -21024 6946 -20990
rect 7410 -21024 7422 -20990
rect 6934 -21030 7422 -21024
rect 6632 -21144 6638 -21084
rect 6698 -21144 6704 -21084
rect 7144 -21182 7204 -21030
rect 7138 -21242 7144 -21182
rect 7204 -21242 7210 -21182
rect 6636 -21338 6642 -21278
rect 6702 -21338 6708 -21278
rect 5100 -21402 6194 -21342
rect 5100 -21506 5160 -21402
rect 6134 -21506 6194 -21402
rect 4898 -21512 5386 -21506
rect 4898 -21546 4910 -21512
rect 5374 -21546 5386 -21512
rect 4898 -21552 5386 -21546
rect 5916 -21512 6404 -21506
rect 5916 -21546 5928 -21512
rect 6392 -21546 6404 -21512
rect 5916 -21552 6404 -21546
rect 3632 -22172 3638 -21636
rect 4606 -21640 4616 -21596
rect 3592 -22184 3638 -22172
rect 4610 -22172 4616 -21640
rect 4650 -21640 4666 -21596
rect 5628 -21596 5674 -21584
rect 4650 -22172 4656 -21640
rect 5628 -22130 5634 -21596
rect 4610 -22184 4656 -22172
rect 5620 -22172 5634 -22130
rect 5668 -22130 5674 -21596
rect 6642 -21596 6702 -21338
rect 7144 -21506 7204 -21242
rect 7656 -21398 7716 -20940
rect 8676 -20940 8688 -20900
rect 8722 -20406 8738 -20364
rect 9696 -20364 9756 -20220
rect 9988 -20280 10476 -20274
rect 9988 -20314 10000 -20280
rect 10464 -20314 10476 -20280
rect 9988 -20320 10476 -20314
rect 9696 -20400 9706 -20364
rect 8722 -20900 8728 -20406
rect 8722 -20940 8736 -20900
rect 9700 -20906 9706 -20400
rect 7952 -20990 8440 -20984
rect 7952 -21024 7964 -20990
rect 8428 -21024 8440 -20990
rect 7952 -21030 8440 -21024
rect 8166 -21182 8226 -21030
rect 8676 -21084 8736 -20940
rect 9690 -20940 9706 -20906
rect 9740 -20400 9756 -20364
rect 10712 -20364 10772 -20122
rect 11006 -20280 11494 -20274
rect 11006 -20314 11018 -20280
rect 11482 -20314 11494 -20280
rect 11006 -20320 11494 -20314
rect 10712 -20390 10724 -20364
rect 9740 -20906 9746 -20400
rect 10718 -20884 10724 -20390
rect 9740 -20940 9750 -20906
rect 8970 -20990 9458 -20984
rect 8970 -21024 8982 -20990
rect 9446 -21024 9458 -20990
rect 8970 -21030 9458 -21024
rect 8670 -21144 8676 -21084
rect 8736 -21144 8742 -21084
rect 9190 -21176 9250 -21030
rect 7650 -21458 7656 -21398
rect 7716 -21458 7722 -21398
rect 6934 -21512 7422 -21506
rect 6934 -21546 6946 -21512
rect 7410 -21546 7422 -21512
rect 6934 -21552 7422 -21546
rect 6642 -21648 6652 -21596
rect 5668 -22172 5680 -22130
rect 2862 -22222 3350 -22216
rect 2862 -22256 2874 -22222
rect 3338 -22256 3350 -22222
rect 2862 -22262 3350 -22256
rect 3880 -22222 4368 -22216
rect 3880 -22256 3892 -22222
rect 4356 -22256 4368 -22222
rect 3880 -22262 4368 -22256
rect 4898 -22222 5386 -22216
rect 4898 -22256 4910 -22222
rect 5374 -22256 5386 -22222
rect 4898 -22262 5386 -22256
rect 2330 -22374 2336 -22314
rect 2396 -22374 2402 -22314
rect 5620 -22440 5680 -22172
rect 6646 -22172 6652 -21648
rect 6686 -21648 6702 -21596
rect 7656 -21596 7716 -21458
rect 8166 -21506 8226 -21242
rect 9188 -21182 9250 -21176
rect 9248 -21242 9250 -21182
rect 9188 -21248 9250 -21242
rect 8664 -21338 8670 -21278
rect 8730 -21338 8736 -21278
rect 7952 -21512 8440 -21506
rect 7952 -21546 7964 -21512
rect 8428 -21546 8440 -21512
rect 7952 -21552 8440 -21546
rect 7656 -21636 7670 -21596
rect 6686 -22172 6692 -21648
rect 7664 -22118 7670 -21636
rect 6646 -22184 6692 -22172
rect 7658 -22172 7670 -22118
rect 7704 -21636 7716 -21596
rect 8670 -21596 8730 -21338
rect 9190 -21506 9250 -21248
rect 9690 -21398 9750 -20940
rect 10708 -20940 10724 -20884
rect 10758 -20390 10772 -20364
rect 11730 -20364 11790 -20010
rect 12024 -20280 12512 -20274
rect 12024 -20314 12036 -20280
rect 12500 -20314 12512 -20280
rect 12024 -20320 12512 -20314
rect 13042 -20280 13530 -20274
rect 13042 -20314 13054 -20280
rect 13518 -20314 13530 -20280
rect 13042 -20320 13530 -20314
rect 10758 -20884 10764 -20390
rect 11730 -20396 11742 -20364
rect 10758 -20940 10768 -20884
rect 9988 -20990 10476 -20984
rect 9988 -21024 10000 -20990
rect 10464 -21024 10476 -20990
rect 9988 -21030 10252 -21024
rect 10264 -21030 10476 -21024
rect 10192 -21182 10252 -21030
rect 10538 -21064 10598 -21058
rect 10708 -21064 10768 -20940
rect 11736 -20940 11742 -20396
rect 11776 -20396 11790 -20364
rect 12754 -20364 12800 -20352
rect 11776 -20940 11782 -20396
rect 12754 -20870 12760 -20364
rect 11736 -20952 11782 -20940
rect 12750 -20940 12760 -20870
rect 12794 -20870 12800 -20364
rect 13766 -20364 13826 -20010
rect 15308 -20048 15368 -19796
rect 15802 -19838 15862 -19706
rect 16826 -19706 16832 -19166
rect 16866 -19706 16872 -19130
rect 17836 -19130 17896 -18996
rect 18314 -19040 18374 -18562
rect 18856 -18612 18916 -18472
rect 19870 -18472 19886 -18428
rect 19920 -18428 19926 -17896
rect 20888 -17896 20948 -17762
rect 21186 -17812 21674 -17806
rect 21186 -17846 21198 -17812
rect 21662 -17846 21674 -17812
rect 21186 -17852 21674 -17846
rect 20888 -17946 20904 -17896
rect 19920 -18472 19930 -18428
rect 20898 -18444 20904 -17946
rect 19150 -18522 19638 -18516
rect 19150 -18556 19162 -18522
rect 19626 -18556 19638 -18522
rect 19150 -18562 19638 -18556
rect 18850 -18672 18856 -18612
rect 18916 -18672 18922 -18612
rect 18846 -18780 18852 -18720
rect 18912 -18780 18918 -18720
rect 18132 -19046 18620 -19040
rect 18132 -19080 18144 -19046
rect 18608 -19080 18620 -19046
rect 18132 -19086 18620 -19080
rect 17836 -19224 17850 -19130
rect 17844 -19664 17850 -19224
rect 16826 -19718 16872 -19706
rect 17836 -19706 17850 -19664
rect 17884 -19224 17896 -19130
rect 18852 -19130 18912 -18780
rect 19338 -18894 19344 -18834
rect 19404 -18894 19410 -18834
rect 19344 -19040 19404 -18894
rect 19870 -18936 19930 -18472
rect 20894 -18472 20904 -18444
rect 20938 -17946 20948 -17896
rect 21910 -17896 21970 -17566
rect 22204 -17812 22692 -17806
rect 22204 -17846 22216 -17812
rect 22680 -17846 22692 -17812
rect 22204 -17852 22692 -17846
rect 20938 -18444 20944 -17946
rect 21910 -17948 21922 -17896
rect 21916 -18444 21922 -17948
rect 20938 -18472 20954 -18444
rect 20168 -18522 20656 -18516
rect 20168 -18556 20180 -18522
rect 20644 -18556 20656 -18522
rect 20168 -18562 20656 -18556
rect 20894 -18612 20954 -18472
rect 21910 -18472 21922 -18444
rect 21956 -17948 21970 -17896
rect 22934 -17896 22980 -17884
rect 21956 -18444 21962 -17948
rect 22934 -18438 22940 -17896
rect 21956 -18472 21970 -18444
rect 21186 -18522 21674 -18516
rect 21186 -18556 21198 -18522
rect 21662 -18556 21674 -18522
rect 21186 -18562 21674 -18556
rect 20888 -18672 20894 -18612
rect 20954 -18672 20960 -18612
rect 20884 -18780 20890 -18720
rect 20950 -18780 20956 -18720
rect 20376 -18894 20382 -18834
rect 20442 -18894 20448 -18834
rect 19864 -18996 19870 -18936
rect 19930 -18996 19936 -18936
rect 20382 -19040 20442 -18894
rect 19150 -19046 19638 -19040
rect 19150 -19080 19162 -19046
rect 19626 -19080 19638 -19046
rect 19150 -19086 19638 -19080
rect 20168 -19046 20656 -19040
rect 20168 -19080 20180 -19046
rect 20644 -19080 20656 -19046
rect 20168 -19086 20656 -19080
rect 18852 -19196 18868 -19130
rect 17884 -19664 17890 -19224
rect 17884 -19706 17896 -19664
rect 16096 -19756 16584 -19750
rect 16096 -19790 16108 -19756
rect 16572 -19790 16584 -19756
rect 16096 -19796 16584 -19790
rect 17114 -19756 17602 -19750
rect 17114 -19790 17126 -19756
rect 17590 -19790 17602 -19756
rect 17114 -19796 17602 -19790
rect 15796 -19898 15802 -19838
rect 15862 -19898 15868 -19838
rect 16150 -19898 16156 -19838
rect 16216 -19898 16222 -19838
rect 15792 -20010 15798 -19950
rect 15858 -20010 15864 -19950
rect 15302 -20108 15308 -20048
rect 15368 -20108 15374 -20048
rect 14060 -20280 14548 -20274
rect 14060 -20314 14072 -20280
rect 14536 -20314 14548 -20280
rect 14060 -20320 14548 -20314
rect 15078 -20280 15566 -20274
rect 15078 -20314 15090 -20280
rect 15554 -20314 15566 -20280
rect 15078 -20320 15566 -20314
rect 13766 -20402 13778 -20364
rect 12794 -20940 12810 -20870
rect 11006 -20990 11494 -20984
rect 11006 -21024 11018 -20990
rect 11482 -21024 11494 -20990
rect 11006 -21030 11494 -21024
rect 12024 -20990 12512 -20984
rect 12024 -21024 12036 -20990
rect 12500 -21024 12512 -20990
rect 12024 -21030 12512 -21024
rect 10702 -21124 10708 -21064
rect 10768 -21124 10774 -21064
rect 10186 -21242 10192 -21182
rect 10252 -21242 10258 -21182
rect 9684 -21458 9690 -21398
rect 9750 -21458 9756 -21398
rect 8970 -21512 9458 -21506
rect 8970 -21546 8982 -21512
rect 9446 -21546 9458 -21512
rect 8970 -21552 9458 -21546
rect 7704 -22118 7710 -21636
rect 8670 -21656 8688 -21596
rect 7704 -22172 7718 -22118
rect 5916 -22222 6404 -22216
rect 5916 -22256 5928 -22222
rect 6392 -22256 6404 -22222
rect 5916 -22262 6256 -22256
rect 6316 -22262 6404 -22256
rect 6934 -22222 7422 -22216
rect 6934 -22256 6946 -22222
rect 7410 -22256 7422 -22222
rect 6934 -22262 7422 -22256
rect 6140 -22428 6200 -22262
rect 2224 -22500 2230 -22440
rect 2290 -22500 2296 -22440
rect 5614 -22500 5620 -22440
rect 5680 -22500 5686 -22440
rect 6134 -22488 6140 -22428
rect 6200 -22488 6206 -22428
rect 4596 -22610 4602 -22550
rect 4662 -22610 4668 -22550
rect 6632 -22610 6638 -22550
rect 6698 -22610 6704 -22550
rect 2862 -22746 3350 -22740
rect 2862 -22780 2874 -22746
rect 3338 -22780 3350 -22746
rect 2862 -22786 3350 -22780
rect 3880 -22746 4368 -22740
rect 3880 -22780 3892 -22746
rect 4356 -22780 4368 -22746
rect 3880 -22786 4368 -22780
rect 2574 -22830 2620 -22818
rect 2574 -23380 2580 -22830
rect 2568 -23406 2580 -23380
rect 2614 -23380 2620 -22830
rect 3592 -22830 3638 -22818
rect 3592 -23352 3598 -22830
rect 2614 -23406 2628 -23380
rect 2568 -23544 2628 -23406
rect 3580 -23406 3598 -23352
rect 3632 -23352 3638 -22830
rect 4602 -22830 4662 -22610
rect 6250 -22704 6256 -22644
rect 6316 -22704 6322 -22644
rect 6256 -22740 6316 -22704
rect 4898 -22746 5386 -22740
rect 4898 -22780 4910 -22746
rect 5374 -22780 5386 -22746
rect 4898 -22786 5386 -22780
rect 5916 -22746 6404 -22740
rect 5916 -22780 5928 -22746
rect 6392 -22780 6404 -22746
rect 5916 -22786 6404 -22780
rect 4602 -22890 4616 -22830
rect 3632 -23406 3640 -23352
rect 2862 -23456 3350 -23450
rect 2862 -23490 2874 -23456
rect 3338 -23490 3350 -23456
rect 2862 -23496 3350 -23490
rect 3082 -23544 3142 -23496
rect 3580 -23544 3640 -23406
rect 4610 -23406 4616 -22890
rect 4650 -22890 4662 -22830
rect 5628 -22830 5674 -22818
rect 4650 -23406 4656 -22890
rect 5628 -23362 5634 -22830
rect 4610 -23418 4656 -23406
rect 5622 -23406 5634 -23362
rect 5668 -23362 5674 -22830
rect 6638 -22830 6698 -22610
rect 7140 -22644 7200 -22262
rect 7658 -22550 7718 -22172
rect 8682 -22172 8688 -21656
rect 8722 -21656 8730 -21596
rect 9690 -21596 9750 -21458
rect 10192 -21506 10252 -21242
rect 10538 -21278 10598 -21124
rect 10532 -21338 10538 -21278
rect 10598 -21338 10604 -21278
rect 10708 -21332 10714 -21272
rect 10774 -21332 10780 -21272
rect 9988 -21512 10252 -21506
rect 10264 -21512 10476 -21506
rect 9988 -21546 10000 -21512
rect 10464 -21546 10476 -21512
rect 9988 -21552 10476 -21546
rect 9690 -21636 9706 -21596
rect 8722 -22172 8728 -21656
rect 9700 -22106 9706 -21636
rect 8682 -22184 8728 -22172
rect 9694 -22172 9706 -22106
rect 9740 -21636 9750 -21596
rect 10714 -21596 10774 -21332
rect 11230 -21334 11290 -21030
rect 12244 -21170 12304 -21030
rect 12750 -21064 12810 -20940
rect 13772 -20940 13778 -20402
rect 13812 -20402 13826 -20364
rect 14790 -20364 14836 -20352
rect 13812 -20940 13818 -20402
rect 14790 -20870 14796 -20364
rect 13772 -20952 13818 -20940
rect 14782 -20940 14796 -20870
rect 14830 -20870 14836 -20364
rect 15798 -20364 15858 -20010
rect 16156 -20156 16216 -19898
rect 16346 -20048 16406 -19796
rect 17322 -20048 17382 -19796
rect 16340 -20108 16346 -20048
rect 16406 -20108 16412 -20048
rect 17316 -20108 17322 -20048
rect 17382 -20108 17388 -20048
rect 17836 -20160 17896 -19706
rect 18862 -19706 18868 -19196
rect 18902 -19196 18912 -19130
rect 19880 -19130 19926 -19118
rect 18902 -19706 18908 -19196
rect 19880 -19662 19886 -19130
rect 18862 -19718 18908 -19706
rect 19874 -19706 19886 -19662
rect 19920 -19662 19926 -19130
rect 20890 -19130 20950 -18780
rect 21408 -18834 21468 -18562
rect 21910 -18654 21970 -18472
rect 22924 -18472 22940 -18438
rect 22974 -18438 22980 -17896
rect 22974 -18472 22984 -18438
rect 22204 -18522 22692 -18516
rect 22204 -18556 22216 -18522
rect 22680 -18556 22692 -18522
rect 22204 -18562 22692 -18556
rect 22418 -18654 22478 -18562
rect 22924 -18654 22984 -18472
rect 21910 -18714 22984 -18654
rect 21402 -18894 21408 -18834
rect 21468 -18894 21474 -18834
rect 21906 -18996 21912 -18936
rect 21972 -18996 21978 -18936
rect 21186 -19046 21674 -19040
rect 21186 -19080 21198 -19046
rect 21662 -19080 21674 -19046
rect 21186 -19086 21674 -19080
rect 20890 -19182 20904 -19130
rect 20898 -19656 20904 -19182
rect 19920 -19706 19934 -19662
rect 18132 -19756 18620 -19750
rect 18132 -19790 18144 -19756
rect 18608 -19790 18620 -19756
rect 18132 -19796 18620 -19790
rect 19150 -19756 19638 -19750
rect 19150 -19790 19162 -19756
rect 19626 -19790 19638 -19756
rect 19150 -19796 19638 -19790
rect 18338 -20048 18398 -19796
rect 19874 -19838 19934 -19706
rect 20892 -19706 20904 -19656
rect 20938 -19182 20950 -19130
rect 21912 -19130 21972 -18996
rect 22204 -19046 22692 -19040
rect 22204 -19080 22216 -19046
rect 22680 -19080 22692 -19046
rect 22204 -19086 22692 -19080
rect 21912 -19164 21922 -19130
rect 20938 -19656 20944 -19182
rect 20938 -19706 20952 -19656
rect 21916 -19662 21922 -19164
rect 20168 -19756 20656 -19750
rect 20168 -19790 20180 -19756
rect 20644 -19790 20656 -19756
rect 20168 -19796 20656 -19790
rect 19868 -19898 19874 -19838
rect 19934 -19898 19940 -19838
rect 18332 -20108 18338 -20048
rect 18398 -20108 18404 -20048
rect 20358 -20108 20364 -20048
rect 20424 -20108 20430 -20048
rect 16156 -20222 16216 -20216
rect 17830 -20220 17836 -20160
rect 17896 -20220 17902 -20160
rect 19866 -20220 19872 -20160
rect 19932 -20220 19938 -20160
rect 16096 -20280 16584 -20274
rect 16096 -20314 16108 -20280
rect 16572 -20314 16584 -20280
rect 16096 -20320 16584 -20314
rect 17114 -20280 17602 -20274
rect 17114 -20314 17126 -20280
rect 17590 -20314 17602 -20280
rect 17114 -20320 17602 -20314
rect 15798 -20406 15814 -20364
rect 14830 -20940 14842 -20870
rect 13042 -20990 13530 -20984
rect 13042 -21024 13054 -20990
rect 13518 -21024 13530 -20990
rect 13042 -21030 13530 -21024
rect 14060 -20990 14548 -20984
rect 14060 -21024 14072 -20990
rect 14536 -21024 14548 -20990
rect 14060 -21030 14548 -21024
rect 12744 -21124 12750 -21064
rect 12810 -21124 12816 -21064
rect 13266 -21170 13326 -21030
rect 14280 -21170 14340 -21030
rect 14782 -21064 14842 -20940
rect 15808 -20940 15814 -20406
rect 15848 -20406 15858 -20364
rect 16826 -20364 16872 -20352
rect 15848 -20940 15854 -20406
rect 16826 -20904 16832 -20364
rect 15808 -20952 15854 -20940
rect 16822 -20940 16832 -20904
rect 16866 -20904 16872 -20364
rect 17836 -20364 17896 -20220
rect 18132 -20280 18620 -20274
rect 18132 -20314 18144 -20280
rect 18608 -20314 18620 -20280
rect 18132 -20320 18620 -20314
rect 19150 -20280 19638 -20274
rect 19150 -20314 19162 -20280
rect 19626 -20314 19638 -20280
rect 19150 -20320 19638 -20314
rect 17836 -20402 17850 -20364
rect 17844 -20888 17850 -20402
rect 16866 -20940 16882 -20904
rect 15078 -20990 15566 -20984
rect 15078 -21024 15090 -20990
rect 15554 -21024 15566 -20990
rect 15078 -21030 15566 -21024
rect 16096 -20990 16584 -20984
rect 16096 -21024 16108 -20990
rect 16572 -21024 16584 -20990
rect 16096 -21030 16584 -21024
rect 14776 -21124 14782 -21064
rect 14842 -21124 14848 -21064
rect 15282 -21070 15342 -21030
rect 16308 -21070 16368 -21030
rect 16822 -21064 16882 -20940
rect 17840 -20940 17850 -20888
rect 17884 -20402 17896 -20364
rect 18862 -20364 18908 -20352
rect 17884 -20888 17890 -20402
rect 17884 -20940 17900 -20888
rect 18862 -20896 18868 -20364
rect 17114 -20990 17602 -20984
rect 17114 -21024 17126 -20990
rect 17590 -21024 17602 -20990
rect 17114 -21030 17602 -21024
rect 15282 -21130 16368 -21070
rect 16816 -21124 16822 -21064
rect 16882 -21124 16888 -21064
rect 15282 -21170 15342 -21130
rect 12244 -21230 15342 -21170
rect 15794 -21222 15800 -21162
rect 15860 -21222 15866 -21162
rect 12244 -21334 12304 -21230
rect 12736 -21332 12742 -21272
rect 12802 -21332 12808 -21272
rect 11230 -21394 12304 -21334
rect 11230 -21506 11290 -21394
rect 12244 -21506 12304 -21394
rect 11006 -21512 11494 -21506
rect 11006 -21546 11018 -21512
rect 11482 -21546 11494 -21512
rect 11006 -21552 11494 -21546
rect 12024 -21512 12512 -21506
rect 12024 -21546 12036 -21512
rect 12500 -21546 12512 -21512
rect 12024 -21552 12512 -21546
rect 9740 -22106 9746 -21636
rect 10714 -21640 10724 -21596
rect 9740 -22172 9754 -22106
rect 7952 -22222 8440 -22216
rect 7952 -22256 7964 -22222
rect 8428 -22256 8440 -22222
rect 7952 -22262 8440 -22256
rect 8970 -22222 9458 -22216
rect 8970 -22256 8982 -22222
rect 9446 -22256 9458 -22222
rect 8970 -22262 9458 -22256
rect 7652 -22610 7658 -22550
rect 7718 -22610 7724 -22550
rect 8162 -22644 8222 -22262
rect 9694 -22550 9754 -22172
rect 10718 -22172 10724 -21640
rect 10758 -21640 10774 -21596
rect 11736 -21596 11782 -21584
rect 10758 -22172 10764 -21640
rect 11736 -22120 11742 -21596
rect 10718 -22184 10764 -22172
rect 11724 -22172 11742 -22120
rect 11776 -22120 11782 -21596
rect 12742 -21596 12802 -21332
rect 13266 -21506 13326 -21230
rect 14280 -21506 14340 -21230
rect 14780 -21332 14786 -21272
rect 14846 -21332 14852 -21272
rect 13042 -21512 13530 -21506
rect 13042 -21546 13054 -21512
rect 13518 -21546 13530 -21512
rect 13042 -21552 13530 -21546
rect 14060 -21512 14548 -21506
rect 14060 -21546 14072 -21512
rect 14536 -21546 14548 -21512
rect 14060 -21552 14548 -21546
rect 12742 -21640 12760 -21596
rect 11776 -22172 11784 -22120
rect 9988 -22222 10476 -22216
rect 9988 -22256 10000 -22222
rect 10464 -22256 10476 -22222
rect 9988 -22262 10476 -22256
rect 11006 -22222 11494 -22216
rect 11006 -22256 11018 -22222
rect 11482 -22256 11494 -22222
rect 11006 -22262 11494 -22256
rect 8668 -22610 8674 -22550
rect 8734 -22610 8740 -22550
rect 9688 -22610 9694 -22550
rect 9754 -22610 9760 -22550
rect 7134 -22704 7140 -22644
rect 7200 -22704 7206 -22644
rect 8156 -22704 8162 -22644
rect 8222 -22704 8228 -22644
rect 7140 -22740 7200 -22704
rect 8162 -22740 8222 -22704
rect 6934 -22746 7422 -22740
rect 6934 -22780 6946 -22746
rect 7410 -22780 7422 -22746
rect 6934 -22786 7422 -22780
rect 7952 -22746 8440 -22740
rect 7952 -22780 7964 -22746
rect 8428 -22780 8440 -22746
rect 7952 -22786 8440 -22780
rect 6638 -22880 6652 -22830
rect 6646 -23344 6652 -22880
rect 5668 -23406 5682 -23362
rect 3880 -23456 4368 -23450
rect 3880 -23490 3892 -23456
rect 4356 -23490 4368 -23456
rect 3880 -23496 4368 -23490
rect 4898 -23456 5386 -23450
rect 4898 -23490 4910 -23456
rect 5374 -23490 5386 -23456
rect 4898 -23496 5386 -23490
rect 2562 -23604 2568 -23544
rect 2628 -23604 2634 -23544
rect 3076 -23604 3082 -23544
rect 3142 -23604 3148 -23544
rect 3574 -23604 3580 -23544
rect 3640 -23604 3646 -23544
rect 4096 -23762 4156 -23496
rect 5118 -23762 5178 -23496
rect 5622 -23544 5682 -23406
rect 6636 -23406 6652 -23344
rect 6686 -22880 6698 -22830
rect 7664 -22830 7710 -22818
rect 6686 -23344 6692 -22880
rect 6686 -23406 6696 -23344
rect 7664 -23366 7670 -22830
rect 5916 -23456 6404 -23450
rect 5916 -23490 5928 -23456
rect 6392 -23490 6404 -23456
rect 5916 -23496 6404 -23490
rect 5616 -23604 5622 -23544
rect 5682 -23604 5688 -23544
rect 6130 -23656 6190 -23496
rect 6124 -23716 6130 -23656
rect 6190 -23716 6196 -23656
rect 2104 -23822 2110 -23762
rect 2170 -23822 2176 -23762
rect 4090 -23822 4096 -23762
rect 4156 -23822 4162 -23762
rect 5112 -23822 5118 -23762
rect 5178 -23822 5184 -23762
rect 6636 -23866 6696 -23406
rect 7654 -23406 7670 -23366
rect 7704 -23366 7710 -22830
rect 8674 -22830 8734 -22610
rect 10204 -22644 10264 -22262
rect 11220 -22428 11280 -22262
rect 11724 -22314 11784 -22172
rect 12754 -22172 12760 -21640
rect 12794 -21640 12802 -21596
rect 13772 -21596 13818 -21584
rect 12794 -22172 12800 -21640
rect 13772 -22120 13778 -21596
rect 12754 -22184 12800 -22172
rect 13766 -22172 13778 -22120
rect 13812 -22120 13818 -21596
rect 14786 -21596 14846 -21332
rect 15282 -21506 15342 -21230
rect 15078 -21512 15566 -21506
rect 15078 -21546 15090 -21512
rect 15554 -21546 15566 -21512
rect 15078 -21552 15566 -21546
rect 14786 -21644 14796 -21596
rect 13812 -22172 13826 -22120
rect 12024 -22222 12512 -22216
rect 12024 -22256 12036 -22222
rect 12500 -22256 12512 -22222
rect 12024 -22262 12512 -22256
rect 13042 -22222 13530 -22216
rect 13042 -22256 13054 -22222
rect 13518 -22256 13530 -22222
rect 13042 -22262 13530 -22256
rect 13766 -22314 13826 -22172
rect 14790 -22172 14796 -21644
rect 14830 -21644 14846 -21596
rect 15800 -21596 15860 -21222
rect 16308 -21506 16368 -21130
rect 16808 -21332 16814 -21272
rect 16874 -21332 16880 -21272
rect 16096 -21512 16584 -21506
rect 16096 -21546 16108 -21512
rect 16572 -21546 16584 -21512
rect 16096 -21552 16584 -21546
rect 15800 -21632 15814 -21596
rect 14830 -22172 14836 -21644
rect 15808 -22128 15814 -21632
rect 14790 -22184 14836 -22172
rect 15802 -22172 15814 -22128
rect 15848 -21632 15860 -21596
rect 16814 -21596 16874 -21332
rect 17328 -21506 17388 -21030
rect 17840 -21398 17900 -20940
rect 18852 -20940 18868 -20896
rect 18902 -20896 18908 -20364
rect 19872 -20364 19932 -20220
rect 20364 -20274 20424 -20108
rect 20168 -20280 20656 -20274
rect 20168 -20314 20180 -20280
rect 20644 -20314 20656 -20280
rect 20168 -20320 20656 -20314
rect 19872 -20422 19886 -20364
rect 18902 -20940 18912 -20896
rect 19880 -20900 19886 -20422
rect 18132 -20990 18620 -20984
rect 18132 -21024 18144 -20990
rect 18608 -21024 18620 -20990
rect 18132 -21030 18620 -21024
rect 17834 -21458 17840 -21398
rect 17900 -21458 17906 -21398
rect 17114 -21512 17602 -21506
rect 17114 -21546 17126 -21512
rect 17590 -21546 17602 -21512
rect 17114 -21552 17602 -21546
rect 15848 -22128 15854 -21632
rect 16814 -21644 16832 -21596
rect 15848 -22172 15862 -22128
rect 14060 -22222 14548 -22216
rect 14060 -22256 14072 -22222
rect 14536 -22256 14548 -22222
rect 14060 -22262 14548 -22256
rect 15078 -22222 15566 -22216
rect 15078 -22256 15090 -22222
rect 15554 -22256 15566 -22222
rect 15078 -22262 15566 -22256
rect 15802 -22314 15862 -22172
rect 16826 -22172 16832 -21644
rect 16866 -21644 16874 -21596
rect 17840 -21596 17900 -21458
rect 18344 -21506 18404 -21030
rect 18852 -21272 18912 -20940
rect 19870 -20940 19886 -20900
rect 19920 -20422 19932 -20364
rect 20892 -20364 20952 -19706
rect 21908 -19706 21922 -19662
rect 21956 -19164 21972 -19130
rect 22934 -19130 22980 -19118
rect 21956 -19662 21962 -19164
rect 21956 -19706 21968 -19662
rect 22934 -19676 22940 -19130
rect 21186 -19756 21674 -19750
rect 21186 -19790 21198 -19756
rect 21662 -19790 21674 -19756
rect 21186 -19796 21674 -19790
rect 21394 -20048 21454 -19796
rect 21908 -19888 21968 -19706
rect 22924 -19706 22940 -19676
rect 22974 -19676 22980 -19130
rect 22974 -19706 22984 -19676
rect 22204 -19756 22692 -19750
rect 22204 -19790 22216 -19756
rect 22680 -19790 22692 -19756
rect 22204 -19796 22692 -19790
rect 22414 -19888 22474 -19796
rect 22924 -19888 22984 -19706
rect 21908 -19948 22984 -19888
rect 21388 -20108 21394 -20048
rect 21454 -20108 21460 -20048
rect 21908 -20160 21968 -19948
rect 21902 -20220 21908 -20160
rect 21968 -20220 21974 -20160
rect 21186 -20280 21674 -20274
rect 21186 -20314 21198 -20280
rect 21662 -20314 21674 -20280
rect 21186 -20320 21674 -20314
rect 22204 -20280 22692 -20274
rect 22204 -20314 22216 -20280
rect 22680 -20314 22692 -20280
rect 22204 -20320 22692 -20314
rect 20892 -20406 20904 -20364
rect 19920 -20900 19926 -20422
rect 20898 -20886 20904 -20406
rect 19920 -20940 19930 -20900
rect 19150 -20990 19638 -20984
rect 19150 -21024 19162 -20990
rect 19626 -21024 19638 -20990
rect 19150 -21030 19638 -21024
rect 18846 -21332 18852 -21272
rect 18912 -21332 18918 -21272
rect 19378 -21506 19438 -21030
rect 19870 -21398 19930 -20940
rect 20892 -20940 20904 -20886
rect 20938 -20406 20952 -20364
rect 21916 -20364 21962 -20352
rect 20938 -20886 20944 -20406
rect 20938 -20940 20952 -20886
rect 21916 -20894 21922 -20364
rect 20168 -20990 20656 -20984
rect 20168 -21024 20180 -20990
rect 20644 -21024 20656 -20990
rect 20168 -21030 20656 -21024
rect 20396 -21396 20456 -21030
rect 20892 -21272 20952 -20940
rect 21906 -20940 21922 -20894
rect 21956 -20894 21962 -20364
rect 22934 -20364 22980 -20352
rect 21956 -20940 21966 -20894
rect 22934 -20912 22940 -20364
rect 21186 -20990 21674 -20984
rect 21186 -21024 21198 -20990
rect 21662 -21024 21674 -20990
rect 21186 -21030 21674 -21024
rect 21410 -21268 21470 -21030
rect 21906 -21066 21966 -20940
rect 22926 -20940 22940 -20912
rect 22974 -20912 22980 -20364
rect 22974 -20940 22986 -20912
rect 22204 -20990 22692 -20984
rect 22204 -21024 22216 -20990
rect 22680 -21024 22692 -20990
rect 22204 -21030 22692 -21024
rect 22412 -21064 22472 -21030
rect 22926 -21064 22986 -20940
rect 22412 -21066 22986 -21064
rect 21906 -21126 22986 -21066
rect 21906 -21162 21966 -21126
rect 21900 -21222 21906 -21162
rect 21966 -21222 21972 -21162
rect 20886 -21332 20892 -21272
rect 20952 -21332 20958 -21272
rect 21404 -21328 21410 -21268
rect 21470 -21328 21476 -21268
rect 19864 -21458 19870 -21398
rect 19930 -21458 19936 -21398
rect 18132 -21512 18620 -21506
rect 18132 -21546 18144 -21512
rect 18608 -21546 18620 -21512
rect 18132 -21552 18620 -21546
rect 19150 -21512 19638 -21506
rect 19150 -21546 19162 -21512
rect 19626 -21546 19638 -21512
rect 19150 -21552 19638 -21546
rect 17840 -21642 17850 -21596
rect 16866 -22172 16872 -21644
rect 17844 -22112 17850 -21642
rect 16826 -22184 16872 -22172
rect 17838 -22172 17850 -22112
rect 17884 -21642 17900 -21596
rect 18862 -21596 18908 -21584
rect 17884 -22112 17890 -21642
rect 17884 -22172 17898 -22112
rect 18862 -22128 18868 -21596
rect 16096 -22222 16584 -22216
rect 16096 -22256 16108 -22222
rect 16572 -22256 16584 -22222
rect 16096 -22262 16584 -22256
rect 17114 -22222 17602 -22216
rect 17114 -22256 17126 -22222
rect 17590 -22256 17602 -22222
rect 17114 -22262 17602 -22256
rect 11718 -22374 11724 -22314
rect 11784 -22374 11790 -22314
rect 13760 -22374 13766 -22314
rect 13826 -22374 13832 -22314
rect 15796 -22374 15802 -22314
rect 15862 -22374 15868 -22314
rect 16308 -22424 16368 -22262
rect 11214 -22488 11220 -22428
rect 11280 -22488 11286 -22428
rect 16302 -22484 16308 -22424
rect 16368 -22484 16374 -22424
rect 10706 -22610 10712 -22550
rect 10772 -22610 10778 -22550
rect 12736 -22610 12742 -22550
rect 12802 -22610 12808 -22550
rect 14774 -22610 14780 -22550
rect 14840 -22610 14846 -22550
rect 16810 -22610 16816 -22550
rect 16876 -22610 16882 -22550
rect 10198 -22704 10204 -22644
rect 10264 -22704 10270 -22644
rect 8970 -22746 9458 -22740
rect 8970 -22780 8982 -22746
rect 9446 -22780 9458 -22746
rect 8970 -22786 9458 -22780
rect 9988 -22746 10476 -22740
rect 9988 -22780 10000 -22746
rect 10464 -22780 10476 -22746
rect 9988 -22786 10476 -22780
rect 7704 -23406 7714 -23366
rect 6934 -23456 7422 -23450
rect 6934 -23490 6946 -23456
rect 7410 -23490 7422 -23456
rect 6934 -23496 7422 -23490
rect 7142 -23656 7202 -23496
rect 7654 -23544 7714 -23406
rect 8674 -23406 8688 -22830
rect 8722 -23406 8734 -22830
rect 9700 -22830 9746 -22818
rect 9700 -23366 9706 -22830
rect 7952 -23456 8440 -23450
rect 7952 -23490 7964 -23456
rect 8428 -23490 8440 -23456
rect 7952 -23496 8440 -23490
rect 7648 -23604 7654 -23544
rect 7714 -23604 7720 -23544
rect 8156 -23656 8216 -23496
rect 7136 -23716 7142 -23656
rect 7202 -23716 7208 -23656
rect 8150 -23716 8156 -23656
rect 8216 -23716 8222 -23656
rect 7650 -23822 7656 -23762
rect 7716 -23822 7722 -23762
rect 8162 -23822 8168 -23762
rect 8228 -23822 8234 -23762
rect 1698 -23926 1704 -23866
rect 1764 -23926 1770 -23866
rect 6126 -23926 6132 -23866
rect 6192 -23926 6198 -23866
rect 6630 -23926 6636 -23866
rect 6696 -23926 6702 -23866
rect 7146 -23926 7152 -23866
rect 7212 -23926 7218 -23866
rect 1070 -24974 1076 -24914
rect 1136 -24974 1142 -24914
rect -2132 -26000 -2126 -25940
rect -2066 -26000 -2060 -25940
rect -944 -26000 -938 -25940
rect -878 -26000 -872 -25940
rect 252 -26000 258 -25940
rect 318 -26000 324 -25940
rect 946 -26000 952 -25940
rect 1012 -26000 1018 -25940
rect 1704 -26430 1764 -23926
rect 6132 -23974 6192 -23926
rect 2862 -23980 3350 -23974
rect 2862 -24014 2874 -23980
rect 3338 -24014 3350 -23980
rect 2862 -24020 3350 -24014
rect 3880 -23980 4368 -23974
rect 3880 -24014 3892 -23980
rect 4356 -24014 4368 -23980
rect 3880 -24020 4368 -24014
rect 4898 -23980 5386 -23974
rect 4898 -24014 4910 -23980
rect 5374 -24014 5386 -23980
rect 4898 -24020 5386 -24014
rect 5916 -23980 6404 -23974
rect 5916 -24014 5928 -23980
rect 6392 -24014 6404 -23980
rect 5916 -24020 6404 -24014
rect 2574 -24064 2620 -24052
rect 2574 -24614 2580 -24064
rect 2568 -24640 2580 -24614
rect 2614 -24614 2620 -24064
rect 3592 -24064 3638 -24052
rect 3592 -24612 3598 -24064
rect 2614 -24640 2628 -24614
rect 2568 -25096 2628 -24640
rect 3580 -24640 3598 -24612
rect 3632 -24612 3638 -24064
rect 4610 -24064 4656 -24052
rect 4610 -24608 4616 -24064
rect 3632 -24640 3640 -24612
rect 2862 -24690 3350 -24684
rect 2862 -24724 2874 -24690
rect 3338 -24724 3350 -24690
rect 2862 -24730 3350 -24724
rect 2562 -25156 2568 -25096
rect 2628 -25156 2634 -25096
rect 2568 -25296 2628 -25156
rect 3066 -25206 3126 -24730
rect 3580 -24998 3640 -24640
rect 4598 -24640 4616 -24608
rect 4650 -24608 4656 -24064
rect 5628 -24064 5674 -24052
rect 5628 -24600 5634 -24064
rect 4650 -24640 4658 -24608
rect 3880 -24690 4368 -24684
rect 3880 -24724 3892 -24690
rect 4356 -24724 4368 -24690
rect 3880 -24730 4368 -24724
rect 3574 -25058 3580 -24998
rect 3640 -25058 3646 -24998
rect 2862 -25212 3350 -25206
rect 2862 -25246 2874 -25212
rect 3338 -25246 3350 -25212
rect 2862 -25252 3350 -25246
rect 2568 -25352 2580 -25296
rect 2574 -25872 2580 -25352
rect 2614 -25352 2628 -25296
rect 3580 -25296 3640 -25058
rect 4088 -25206 4148 -24730
rect 4598 -25096 4658 -24640
rect 5618 -24640 5634 -24600
rect 5668 -24600 5674 -24064
rect 6636 -24064 6696 -23926
rect 7152 -23974 7212 -23926
rect 6934 -23980 7422 -23974
rect 6934 -24014 6946 -23980
rect 7410 -24014 7422 -23980
rect 6934 -24020 7422 -24014
rect 7656 -24064 7716 -23822
rect 8168 -23974 8228 -23822
rect 8674 -23866 8734 -23406
rect 9686 -23406 9706 -23366
rect 9740 -23406 9746 -22830
rect 10712 -22830 10772 -22610
rect 11218 -22686 12288 -22626
rect 11218 -22740 11278 -22686
rect 11006 -22746 11494 -22740
rect 11006 -22780 11018 -22746
rect 11482 -22780 11494 -22746
rect 11006 -22786 11494 -22780
rect 10712 -22886 10724 -22830
rect 10718 -23354 10724 -22886
rect 8970 -23456 9458 -23450
rect 8970 -23490 8982 -23456
rect 9446 -23490 9458 -23456
rect 8970 -23496 9458 -23490
rect 9186 -23762 9246 -23496
rect 9686 -23544 9746 -23406
rect 10712 -23406 10724 -23354
rect 10758 -22886 10772 -22830
rect 11730 -22830 11790 -22686
rect 12228 -22740 12288 -22686
rect 12024 -22746 12512 -22740
rect 12024 -22780 12036 -22746
rect 12500 -22780 12512 -22746
rect 12024 -22786 12512 -22780
rect 11730 -22866 11742 -22830
rect 10758 -23354 10764 -22886
rect 10758 -23406 10772 -23354
rect 11736 -23362 11742 -22866
rect 11728 -23370 11742 -23362
rect 11722 -23406 11742 -23370
rect 11776 -22866 11790 -22830
rect 12742 -22830 12802 -22610
rect 13242 -22682 14330 -22622
rect 13242 -22740 13302 -22682
rect 13042 -22746 13530 -22740
rect 13042 -22780 13054 -22746
rect 13518 -22780 13530 -22746
rect 13042 -22786 13530 -22780
rect 11776 -23362 11782 -22866
rect 12742 -22880 12760 -22830
rect 12754 -23356 12760 -22880
rect 11776 -23406 11788 -23362
rect 9988 -23456 10476 -23450
rect 9988 -23490 10000 -23456
rect 10464 -23490 10476 -23456
rect 9988 -23496 10476 -23490
rect 9680 -23604 9686 -23544
rect 9746 -23604 9752 -23544
rect 10198 -23762 10258 -23496
rect 9180 -23822 9186 -23762
rect 9246 -23822 9252 -23762
rect 9686 -23822 9692 -23762
rect 9752 -23822 9758 -23762
rect 10192 -23822 10198 -23762
rect 10258 -23822 10264 -23762
rect 8668 -23926 8674 -23866
rect 8734 -23926 8740 -23866
rect 7952 -23980 8440 -23974
rect 7952 -24014 7964 -23980
rect 8428 -24014 8440 -23980
rect 7952 -24020 8440 -24014
rect 6636 -24116 6652 -24064
rect 5668 -24640 5678 -24600
rect 4898 -24690 5386 -24684
rect 4898 -24724 4910 -24690
rect 5374 -24724 5386 -24690
rect 4898 -24730 5386 -24724
rect 4592 -25156 4598 -25096
rect 4658 -25156 4664 -25096
rect 3880 -25212 4368 -25206
rect 3880 -25246 3892 -25212
rect 4356 -25246 4368 -25212
rect 3880 -25252 4368 -25246
rect 3580 -25334 3598 -25296
rect 2614 -25872 2620 -25352
rect 3592 -25822 3598 -25334
rect 2574 -25884 2620 -25872
rect 3582 -25872 3598 -25822
rect 3632 -25334 3640 -25296
rect 4598 -25296 4658 -25156
rect 5114 -25206 5174 -24730
rect 5618 -24998 5678 -24640
rect 6646 -24640 6652 -24116
rect 6686 -24116 6696 -24064
rect 6686 -24640 6692 -24116
rect 7654 -24120 7670 -24064
rect 7664 -24598 7670 -24120
rect 6646 -24652 6692 -24640
rect 7654 -24640 7670 -24598
rect 7704 -24116 7716 -24064
rect 8674 -24064 8734 -23926
rect 9186 -23974 9246 -23822
rect 8970 -23980 9458 -23974
rect 8970 -24014 8982 -23980
rect 9446 -24014 9458 -23980
rect 8970 -24020 9458 -24014
rect 9692 -24064 9752 -23822
rect 10198 -23974 10258 -23822
rect 10712 -23866 10772 -23406
rect 11006 -23456 11494 -23450
rect 11006 -23490 11018 -23456
rect 11482 -23490 11494 -23456
rect 11006 -23496 11494 -23490
rect 11062 -23716 11068 -23656
rect 11128 -23716 11134 -23656
rect 10706 -23926 10712 -23866
rect 10772 -23926 10778 -23866
rect 9988 -23980 10476 -23974
rect 9988 -24014 10000 -23980
rect 10464 -24014 10476 -23980
rect 9988 -24020 10476 -24014
rect 8674 -24114 8688 -24064
rect 7704 -24120 7714 -24116
rect 7704 -24598 7710 -24120
rect 7704 -24640 7714 -24598
rect 5916 -24690 6404 -24684
rect 5916 -24724 5928 -24690
rect 6392 -24724 6404 -24690
rect 5916 -24730 6404 -24724
rect 6934 -24690 7422 -24684
rect 6934 -24724 6946 -24690
rect 7410 -24724 7422 -24690
rect 6934 -24730 7422 -24724
rect 7654 -24784 7714 -24640
rect 8682 -24640 8688 -24114
rect 8722 -24114 8734 -24064
rect 8722 -24640 8728 -24114
rect 9686 -24130 9706 -24064
rect 9700 -24606 9706 -24130
rect 8682 -24652 8728 -24640
rect 9692 -24640 9706 -24606
rect 9740 -24104 9752 -24064
rect 10712 -24064 10772 -23926
rect 11068 -23974 11128 -23716
rect 11210 -23762 11270 -23496
rect 11590 -23544 11650 -23538
rect 11204 -23822 11210 -23762
rect 11270 -23822 11276 -23762
rect 11590 -23774 11650 -23604
rect 11728 -23654 11788 -23406
rect 12748 -23406 12760 -23356
rect 12794 -22880 12802 -22830
rect 13766 -22830 13826 -22682
rect 14270 -22740 14330 -22682
rect 14060 -22746 14548 -22740
rect 14060 -22780 14072 -22746
rect 14536 -22780 14548 -22746
rect 14060 -22786 14548 -22780
rect 13766 -22862 13778 -22830
rect 12794 -23356 12800 -22880
rect 13772 -23352 13778 -22862
rect 12794 -23406 12808 -23356
rect 12024 -23456 12512 -23450
rect 12024 -23490 12036 -23456
rect 12500 -23490 12512 -23456
rect 12024 -23496 12512 -23490
rect 11722 -23714 11728 -23654
rect 11788 -23714 11794 -23654
rect 12230 -23762 12290 -23496
rect 12350 -23718 12356 -23658
rect 12416 -23718 12422 -23658
rect 11590 -23834 11790 -23774
rect 12224 -23822 12230 -23762
rect 12290 -23822 12296 -23762
rect 11006 -23980 11494 -23974
rect 11006 -24014 11018 -23980
rect 11482 -24014 11494 -23980
rect 11006 -24020 11494 -24014
rect 9740 -24606 9746 -24104
rect 10712 -24124 10724 -24064
rect 9740 -24640 9752 -24606
rect 7952 -24690 8440 -24684
rect 7952 -24724 7964 -24690
rect 8428 -24724 8440 -24690
rect 7952 -24730 8440 -24724
rect 8970 -24690 9458 -24684
rect 8970 -24724 8982 -24690
rect 9446 -24724 9458 -24690
rect 8970 -24730 9458 -24724
rect 8158 -24784 8218 -24730
rect 7654 -24844 8218 -24784
rect 9174 -24792 9234 -24730
rect 9692 -24792 9752 -24640
rect 10718 -24640 10724 -24124
rect 10758 -24124 10772 -24064
rect 11730 -24064 11790 -23834
rect 12356 -23974 12416 -23718
rect 12748 -23866 12808 -23406
rect 13764 -23406 13778 -23352
rect 13812 -22862 13826 -22830
rect 14780 -22830 14840 -22610
rect 15078 -22746 15566 -22740
rect 15078 -22780 15090 -22746
rect 15554 -22780 15566 -22746
rect 15078 -22786 15566 -22780
rect 16096 -22746 16584 -22740
rect 16096 -22780 16108 -22746
rect 16572 -22780 16584 -22746
rect 16096 -22786 16584 -22780
rect 13812 -23352 13818 -22862
rect 14780 -22874 14796 -22830
rect 13812 -23406 13824 -23352
rect 14790 -23368 14796 -22874
rect 13042 -23456 13530 -23450
rect 13042 -23490 13054 -23456
rect 13518 -23490 13530 -23456
rect 13042 -23496 13530 -23490
rect 13252 -23762 13312 -23496
rect 13396 -23718 13402 -23658
rect 13462 -23718 13468 -23658
rect 13246 -23822 13252 -23762
rect 13312 -23822 13318 -23762
rect 12742 -23926 12748 -23866
rect 12808 -23926 12814 -23866
rect 12024 -23980 12512 -23974
rect 12024 -24014 12036 -23980
rect 12500 -24014 12512 -23980
rect 12024 -24020 12512 -24014
rect 11730 -24092 11742 -24064
rect 10758 -24640 10764 -24124
rect 11736 -24616 11742 -24092
rect 10718 -24652 10764 -24640
rect 11730 -24640 11742 -24616
rect 11776 -24092 11790 -24064
rect 12748 -24064 12808 -23926
rect 13402 -23974 13462 -23718
rect 13764 -23762 13824 -23406
rect 14784 -23406 14796 -23368
rect 14830 -22874 14840 -22830
rect 15808 -22830 15854 -22818
rect 14830 -23368 14836 -22874
rect 15808 -23346 15814 -22830
rect 14830 -23406 14844 -23368
rect 14060 -23456 14548 -23450
rect 14060 -23490 14072 -23456
rect 14536 -23490 14548 -23456
rect 14060 -23496 14548 -23490
rect 13950 -23542 14010 -23536
rect 13758 -23822 13764 -23762
rect 13824 -23822 13830 -23762
rect 13950 -23870 14010 -23602
rect 14270 -23762 14330 -23496
rect 14264 -23822 14270 -23762
rect 14330 -23822 14336 -23762
rect 13766 -23930 14010 -23870
rect 13042 -23980 13530 -23974
rect 13042 -24014 13054 -23980
rect 13518 -24014 13530 -23980
rect 13042 -24020 13530 -24014
rect 11776 -24616 11782 -24092
rect 12748 -24130 12760 -24064
rect 11776 -24640 11790 -24616
rect 9988 -24690 10476 -24684
rect 9988 -24724 10000 -24690
rect 10464 -24724 10476 -24690
rect 9988 -24730 10476 -24724
rect 11006 -24690 11494 -24684
rect 11006 -24724 11018 -24690
rect 11482 -24724 11494 -24690
rect 11006 -24730 11494 -24724
rect 10200 -24792 10260 -24730
rect 9174 -24852 10260 -24792
rect 11220 -24902 11280 -24730
rect 11730 -24798 11790 -24640
rect 12754 -24640 12760 -24130
rect 12794 -24130 12808 -24064
rect 13766 -24064 13826 -23930
rect 14270 -23974 14330 -23822
rect 14784 -23866 14844 -23406
rect 15800 -23406 15814 -23346
rect 15848 -23346 15854 -22830
rect 16816 -22830 16876 -22610
rect 17326 -22644 17386 -22262
rect 17838 -22550 17898 -22172
rect 18856 -22172 18868 -22128
rect 18902 -22128 18908 -21596
rect 19870 -21596 19930 -21458
rect 20396 -21506 20456 -21456
rect 21410 -21506 21470 -21328
rect 21908 -21396 22986 -21338
rect 21902 -21456 21908 -21396
rect 21968 -21398 22986 -21396
rect 21968 -21456 21974 -21398
rect 20168 -21512 20656 -21506
rect 20168 -21546 20180 -21512
rect 20644 -21546 20656 -21512
rect 20168 -21552 20656 -21546
rect 21186 -21512 21674 -21506
rect 21186 -21546 21198 -21512
rect 21662 -21546 21674 -21512
rect 21186 -21552 21674 -21546
rect 19870 -21642 19886 -21596
rect 19880 -22124 19886 -21642
rect 18902 -22172 18916 -22128
rect 18132 -22222 18620 -22216
rect 18132 -22256 18144 -22222
rect 18608 -22256 18620 -22222
rect 18132 -22262 18620 -22256
rect 17832 -22610 17838 -22550
rect 17898 -22610 17904 -22550
rect 18346 -22644 18406 -22262
rect 18856 -22314 18916 -22172
rect 19872 -22172 19886 -22124
rect 19920 -21642 19930 -21596
rect 20898 -21596 20944 -21584
rect 19920 -22124 19926 -21642
rect 19920 -22172 19932 -22124
rect 20898 -22128 20904 -21596
rect 19150 -22222 19638 -22216
rect 19150 -22256 19162 -22222
rect 19626 -22256 19638 -22222
rect 19150 -22262 19638 -22256
rect 18850 -22374 18856 -22314
rect 18916 -22374 18922 -22314
rect 18852 -22610 18858 -22550
rect 18918 -22610 18924 -22550
rect 17320 -22704 17326 -22644
rect 17386 -22704 17392 -22644
rect 18340 -22704 18346 -22644
rect 18406 -22704 18412 -22644
rect 17326 -22740 17386 -22704
rect 18346 -22740 18406 -22704
rect 17114 -22746 17602 -22740
rect 17114 -22780 17126 -22746
rect 17590 -22780 17602 -22746
rect 17114 -22786 17602 -22780
rect 18132 -22746 18620 -22740
rect 18132 -22780 18144 -22746
rect 18608 -22780 18620 -22746
rect 18132 -22786 18620 -22780
rect 16816 -22874 16832 -22830
rect 15848 -23406 15860 -23346
rect 16826 -23352 16832 -22874
rect 15078 -23456 15566 -23450
rect 15078 -23490 15090 -23456
rect 15554 -23490 15566 -23456
rect 15078 -23496 15566 -23490
rect 15288 -23762 15348 -23496
rect 15800 -23544 15860 -23406
rect 16816 -23406 16832 -23352
rect 16866 -22874 16876 -22830
rect 17844 -22830 17890 -22818
rect 16866 -23352 16872 -22874
rect 16866 -23406 16876 -23352
rect 17844 -23374 17850 -22830
rect 16096 -23456 16584 -23450
rect 16096 -23490 16108 -23456
rect 16572 -23490 16584 -23456
rect 16096 -23496 16584 -23490
rect 15794 -23604 15800 -23544
rect 15860 -23604 15866 -23544
rect 16308 -23762 16368 -23496
rect 15282 -23822 15288 -23762
rect 15348 -23822 15354 -23762
rect 15794 -23822 15800 -23762
rect 15860 -23822 15866 -23762
rect 16302 -23822 16308 -23762
rect 16368 -23822 16374 -23762
rect 14778 -23926 14784 -23866
rect 14844 -23926 14850 -23866
rect 14060 -23980 14548 -23974
rect 14060 -24014 14072 -23980
rect 14536 -24014 14548 -23980
rect 14060 -24020 14548 -24014
rect 13766 -24098 13778 -24064
rect 12794 -24640 12800 -24130
rect 13772 -24574 13778 -24098
rect 12754 -24652 12800 -24640
rect 13766 -24640 13778 -24574
rect 13812 -24098 13826 -24064
rect 14784 -24064 14844 -23926
rect 15288 -23974 15348 -23822
rect 15078 -23980 15566 -23974
rect 15078 -24014 15090 -23980
rect 15554 -24014 15566 -23980
rect 15078 -24020 15566 -24014
rect 15800 -24064 15860 -23822
rect 16308 -23974 16368 -23822
rect 16816 -23866 16876 -23406
rect 17834 -23406 17850 -23374
rect 17884 -23374 17890 -22830
rect 18858 -22830 18918 -22610
rect 19360 -22644 19420 -22262
rect 19872 -22550 19932 -22172
rect 20888 -22172 20904 -22128
rect 20938 -22128 20944 -21596
rect 21908 -21596 21968 -21456
rect 22410 -21506 22470 -21398
rect 22204 -21512 22692 -21506
rect 22204 -21546 22216 -21512
rect 22680 -21546 22692 -21512
rect 22204 -21552 22692 -21546
rect 21908 -21630 21922 -21596
rect 20938 -22172 20948 -22128
rect 20168 -22222 20656 -22216
rect 20168 -22256 20180 -22222
rect 20644 -22256 20656 -22222
rect 20168 -22262 20656 -22256
rect 19866 -22610 19872 -22550
rect 19932 -22610 19938 -22550
rect 20396 -22644 20456 -22262
rect 20888 -22314 20948 -22172
rect 21916 -22172 21922 -21630
rect 21956 -21630 21968 -21596
rect 22926 -21596 22986 -21398
rect 21956 -22172 21962 -21630
rect 22926 -21634 22940 -21596
rect 21916 -22184 21962 -22172
rect 22934 -22172 22940 -21634
rect 22974 -21634 22986 -21596
rect 22974 -22172 22980 -21634
rect 22934 -22184 22980 -22172
rect 21186 -22222 21674 -22216
rect 21186 -22256 21198 -22222
rect 21408 -22256 21468 -22228
rect 21662 -22256 21674 -22222
rect 21186 -22262 21674 -22256
rect 22204 -22222 22692 -22216
rect 22204 -22256 22216 -22222
rect 22680 -22256 22692 -22222
rect 22204 -22262 22692 -22256
rect 20882 -22374 20888 -22314
rect 20948 -22374 20954 -22314
rect 21408 -22424 21468 -22262
rect 23034 -22314 23094 -16524
rect 23156 -17438 23162 -17378
rect 23222 -17438 23228 -17378
rect 23162 -18936 23222 -17438
rect 23278 -17702 23338 -16410
rect 23394 -17660 23400 -17600
rect 23460 -17660 23466 -17600
rect 23272 -17762 23278 -17702
rect 23338 -17762 23344 -17702
rect 23156 -18996 23162 -18936
rect 23222 -18996 23228 -18936
rect 23152 -19898 23158 -19838
rect 23218 -19898 23224 -19838
rect 23158 -21162 23218 -19898
rect 23278 -21064 23338 -17762
rect 23272 -21124 23278 -21064
rect 23338 -21124 23344 -21064
rect 23152 -21222 23158 -21162
rect 23218 -21222 23224 -21162
rect 23400 -21396 23460 -17660
rect 23528 -18828 23588 -16306
rect 23526 -18834 23588 -18828
rect 23586 -18894 23588 -18834
rect 23526 -18900 23588 -18894
rect 23528 -21268 23588 -18900
rect 23522 -21328 23528 -21268
rect 23588 -21328 23594 -21268
rect 23394 -21456 23400 -21396
rect 23460 -21456 23466 -21396
rect 23028 -22374 23034 -22314
rect 23094 -22374 23100 -22314
rect 21402 -22484 21408 -22424
rect 21468 -22484 21474 -22424
rect 21408 -22548 21468 -22484
rect 20888 -22610 20894 -22550
rect 20954 -22610 20960 -22550
rect 21408 -22608 23154 -22548
rect 19354 -22704 19360 -22644
rect 19420 -22704 19426 -22644
rect 20390 -22704 20396 -22644
rect 20456 -22704 20462 -22644
rect 19360 -22740 19420 -22704
rect 19150 -22746 19420 -22740
rect 19428 -22746 19638 -22740
rect 19150 -22780 19162 -22746
rect 19626 -22780 19638 -22746
rect 19150 -22786 19638 -22780
rect 20168 -22746 20656 -22740
rect 20168 -22780 20180 -22746
rect 20644 -22780 20656 -22746
rect 20168 -22786 20656 -22780
rect 19368 -22790 19428 -22786
rect 18858 -22896 18868 -22830
rect 18862 -23358 18868 -22896
rect 17884 -23406 17894 -23374
rect 17114 -23456 17602 -23450
rect 17114 -23490 17126 -23456
rect 17590 -23490 17602 -23456
rect 17114 -23496 17602 -23490
rect 17330 -23658 17390 -23496
rect 17834 -23544 17894 -23406
rect 18854 -23406 18868 -23358
rect 18902 -22896 18918 -22830
rect 19880 -22830 19926 -22818
rect 18902 -23358 18908 -22896
rect 19880 -23356 19886 -22830
rect 18902 -23406 18914 -23358
rect 18132 -23456 18620 -23450
rect 18132 -23490 18144 -23456
rect 18608 -23490 18620 -23456
rect 18132 -23496 18620 -23490
rect 17828 -23604 17834 -23544
rect 17894 -23604 17900 -23544
rect 18348 -23658 18408 -23496
rect 17324 -23718 17330 -23658
rect 17390 -23718 17396 -23658
rect 18342 -23718 18348 -23658
rect 18408 -23718 18414 -23658
rect 18854 -23866 18914 -23406
rect 19868 -23406 19886 -23356
rect 19920 -23356 19926 -22830
rect 20894 -22830 20954 -22610
rect 21186 -22746 21674 -22740
rect 21186 -22780 21198 -22746
rect 21662 -22780 21674 -22746
rect 21186 -22786 21674 -22780
rect 22204 -22746 22692 -22740
rect 22204 -22780 22216 -22746
rect 22680 -22780 22692 -22746
rect 22204 -22786 22692 -22780
rect 20894 -22890 20904 -22830
rect 19920 -23406 19928 -23356
rect 19150 -23456 19638 -23450
rect 19150 -23490 19162 -23456
rect 19626 -23490 19638 -23456
rect 19150 -23496 19638 -23490
rect 19356 -23652 19416 -23496
rect 19868 -23544 19928 -23406
rect 20898 -23406 20904 -22890
rect 20938 -22890 20954 -22830
rect 21916 -22830 21962 -22818
rect 20938 -23406 20944 -22890
rect 21916 -23362 21922 -22830
rect 20898 -23418 20944 -23406
rect 21910 -23406 21922 -23362
rect 21956 -23362 21962 -22830
rect 22934 -22830 22980 -22818
rect 21956 -23406 21970 -23362
rect 22934 -23364 22940 -22830
rect 20168 -23456 20656 -23450
rect 20168 -23490 20180 -23456
rect 20644 -23490 20656 -23456
rect 20168 -23496 20656 -23490
rect 21186 -23456 21674 -23450
rect 21186 -23490 21198 -23456
rect 21662 -23490 21674 -23456
rect 21186 -23496 21674 -23490
rect 19862 -23604 19868 -23544
rect 19928 -23604 19934 -23544
rect 19356 -23658 19418 -23652
rect 19356 -23718 19358 -23658
rect 19356 -23724 19418 -23718
rect 16810 -23926 16816 -23866
rect 16876 -23926 16882 -23866
rect 17332 -23926 17338 -23866
rect 17398 -23926 17404 -23866
rect 17832 -23926 17838 -23866
rect 17898 -23926 17904 -23866
rect 18340 -23926 18346 -23866
rect 18406 -23926 18412 -23866
rect 18848 -23926 18854 -23866
rect 18914 -23926 18920 -23866
rect 19198 -23926 19204 -23866
rect 19264 -23926 19270 -23866
rect 19356 -23868 19416 -23724
rect 20380 -23762 20440 -23496
rect 21382 -23762 21442 -23496
rect 21910 -23544 21970 -23406
rect 22928 -23406 22940 -23364
rect 22974 -23364 22980 -22830
rect 22974 -23406 22988 -23364
rect 22204 -23456 22692 -23450
rect 22204 -23490 22216 -23456
rect 22680 -23490 22692 -23456
rect 22204 -23496 22692 -23490
rect 22422 -23544 22482 -23496
rect 22928 -23544 22988 -23406
rect 21904 -23604 21910 -23544
rect 21970 -23604 21976 -23544
rect 22416 -23604 22422 -23544
rect 22482 -23604 22488 -23544
rect 22922 -23604 22928 -23544
rect 22988 -23604 22994 -23544
rect 20374 -23822 20380 -23762
rect 20440 -23822 20446 -23762
rect 21376 -23822 21382 -23762
rect 21442 -23822 21448 -23762
rect 16096 -23980 16584 -23974
rect 16096 -24014 16108 -23980
rect 16572 -24014 16584 -23980
rect 16096 -24020 16584 -24014
rect 13812 -24574 13818 -24098
rect 14784 -24140 14796 -24064
rect 13812 -24640 13826 -24574
rect 12024 -24690 12512 -24684
rect 12024 -24724 12036 -24690
rect 12500 -24724 12512 -24690
rect 12024 -24730 12512 -24724
rect 13042 -24690 13530 -24684
rect 13042 -24724 13054 -24690
rect 13518 -24724 13530 -24690
rect 13042 -24730 13530 -24724
rect 11724 -24858 11730 -24798
rect 11790 -24858 11796 -24798
rect 12232 -24902 12292 -24730
rect 13258 -24902 13318 -24730
rect 13766 -24798 13826 -24640
rect 14790 -24640 14796 -24140
rect 14830 -24140 14844 -24064
rect 15796 -24114 15814 -24064
rect 14830 -24640 14836 -24140
rect 15808 -24608 15814 -24114
rect 14790 -24652 14836 -24640
rect 15798 -24640 15814 -24608
rect 15848 -24112 15860 -24064
rect 16816 -24064 16876 -23926
rect 17338 -23974 17398 -23926
rect 17114 -23980 17602 -23974
rect 17114 -24014 17126 -23980
rect 17590 -24014 17602 -23980
rect 17114 -24020 17602 -24014
rect 17338 -24026 17398 -24020
rect 17838 -24064 17898 -23926
rect 18346 -23974 18406 -23926
rect 18132 -23980 18620 -23974
rect 18132 -24014 18144 -23980
rect 18608 -24014 18620 -23980
rect 18132 -24020 18620 -24014
rect 15848 -24114 15856 -24112
rect 15848 -24608 15854 -24114
rect 16816 -24120 16832 -24064
rect 15848 -24640 15858 -24608
rect 14060 -24690 14548 -24684
rect 14060 -24724 14072 -24690
rect 14536 -24724 14548 -24690
rect 14060 -24730 14548 -24724
rect 15078 -24690 15566 -24684
rect 15078 -24724 15090 -24690
rect 15554 -24724 15566 -24690
rect 15078 -24730 15566 -24724
rect 15286 -24790 15346 -24730
rect 15798 -24790 15858 -24640
rect 16826 -24640 16832 -24120
rect 16866 -24120 16876 -24064
rect 16866 -24640 16872 -24120
rect 17832 -24124 17850 -24064
rect 17844 -24602 17850 -24124
rect 17834 -24640 17850 -24602
rect 17884 -24124 17898 -24064
rect 18854 -24064 18914 -23926
rect 19204 -23974 19264 -23926
rect 19356 -23928 19934 -23868
rect 19150 -23980 19638 -23974
rect 19150 -24014 19162 -23980
rect 19626 -24014 19638 -23980
rect 19150 -24020 19638 -24014
rect 18854 -24098 18868 -24064
rect 17884 -24602 17890 -24124
rect 17884 -24640 17894 -24602
rect 18862 -24640 18868 -24098
rect 18902 -24098 18914 -24064
rect 19874 -24064 19934 -23928
rect 23094 -23930 23154 -22608
rect 20168 -23980 20656 -23974
rect 20168 -24014 20180 -23980
rect 20644 -24014 20656 -23980
rect 20168 -24020 20656 -24014
rect 21186 -23980 21674 -23974
rect 21186 -24014 21198 -23980
rect 21662 -24014 21674 -23980
rect 21186 -24020 21674 -24014
rect 22204 -23980 22692 -23974
rect 22204 -24014 22216 -23980
rect 22680 -24014 22692 -23980
rect 22204 -24020 22692 -24014
rect 22934 -23990 23154 -23930
rect 18902 -24640 18908 -24098
rect 19874 -24102 19886 -24064
rect 16826 -24652 16872 -24640
rect 18862 -24652 18908 -24640
rect 19880 -24640 19886 -24102
rect 19920 -24102 19934 -24064
rect 20898 -24064 20944 -24052
rect 19920 -24640 19926 -24102
rect 20898 -24608 20904 -24064
rect 19880 -24652 19926 -24640
rect 20888 -24640 20904 -24608
rect 20938 -24608 20944 -24064
rect 21916 -24064 21962 -24052
rect 21916 -24592 21922 -24064
rect 20938 -24640 20948 -24608
rect 16096 -24690 16584 -24684
rect 16096 -24724 16108 -24690
rect 16572 -24724 16584 -24690
rect 16096 -24730 16584 -24724
rect 17114 -24690 17602 -24684
rect 17114 -24724 17126 -24690
rect 17590 -24724 17602 -24690
rect 17114 -24730 17330 -24724
rect 17390 -24730 17602 -24724
rect 18132 -24690 18620 -24684
rect 18132 -24724 18144 -24690
rect 18608 -24724 18620 -24690
rect 18132 -24730 18620 -24724
rect 19150 -24690 19638 -24684
rect 19150 -24724 19162 -24690
rect 19626 -24724 19638 -24690
rect 19150 -24730 19638 -24724
rect 20168 -24690 20656 -24684
rect 20168 -24724 20180 -24690
rect 20644 -24724 20656 -24690
rect 20168 -24730 20656 -24724
rect 16304 -24790 16364 -24730
rect 13760 -24858 13766 -24798
rect 13826 -24858 13832 -24798
rect 15286 -24850 16364 -24790
rect 11220 -24962 13318 -24902
rect 5612 -25058 5618 -24998
rect 5678 -25058 5684 -24998
rect 7650 -25058 7656 -24998
rect 7716 -25058 7722 -24998
rect 9682 -25058 9688 -24998
rect 9748 -25058 9754 -24998
rect 11720 -25058 11726 -24998
rect 11786 -25058 11792 -24998
rect 13754 -25058 13760 -24998
rect 13820 -25058 13826 -24998
rect 15794 -25058 15800 -24998
rect 15860 -25058 15866 -24998
rect 17828 -25058 17834 -24998
rect 17894 -25058 17900 -24998
rect 19862 -25058 19868 -24998
rect 19928 -25058 19934 -24998
rect 4898 -25212 5386 -25206
rect 4898 -25246 4910 -25212
rect 5374 -25246 5386 -25212
rect 4898 -25252 5386 -25246
rect 3632 -25822 3638 -25334
rect 4598 -25344 4616 -25296
rect 3632 -25872 3642 -25822
rect 2862 -25922 3350 -25916
rect 2862 -25956 2874 -25922
rect 3338 -25956 3350 -25922
rect 2862 -25962 3350 -25956
rect 3066 -26028 3126 -25962
rect 3582 -26028 3642 -25872
rect 4610 -25872 4616 -25344
rect 4650 -25344 4658 -25296
rect 5618 -25296 5678 -25058
rect 6630 -25156 6636 -25096
rect 6696 -25156 6702 -25096
rect 5916 -25212 6404 -25206
rect 5916 -25246 5928 -25212
rect 6392 -25246 6404 -25212
rect 5916 -25252 6404 -25246
rect 5618 -25328 5634 -25296
rect 4650 -25872 4656 -25344
rect 5628 -25782 5634 -25328
rect 4610 -25884 4656 -25872
rect 5620 -25872 5634 -25844
rect 5668 -25328 5678 -25296
rect 6636 -25296 6696 -25156
rect 6934 -25212 7422 -25206
rect 6934 -25246 6946 -25212
rect 7410 -25246 7422 -25212
rect 6934 -25252 7422 -25246
rect 5668 -25782 5674 -25328
rect 6636 -25352 6652 -25296
rect 5668 -25872 5680 -25844
rect 3880 -25922 4368 -25916
rect 3880 -25956 3892 -25922
rect 4356 -25956 4368 -25922
rect 3880 -25962 4368 -25956
rect 4898 -25922 5386 -25916
rect 4898 -25956 4910 -25922
rect 5374 -25956 5386 -25922
rect 4898 -25962 5386 -25956
rect 4114 -26028 4174 -25962
rect 5104 -26028 5164 -25962
rect 5620 -26028 5680 -25872
rect 6646 -25872 6652 -25352
rect 6686 -25352 6696 -25296
rect 7656 -25296 7716 -25058
rect 8666 -25156 8672 -25096
rect 8732 -25156 8738 -25096
rect 7952 -25212 8440 -25206
rect 7952 -25246 7964 -25212
rect 8428 -25246 8440 -25212
rect 7952 -25252 8440 -25246
rect 7656 -25342 7670 -25296
rect 6686 -25872 6692 -25352
rect 7664 -25844 7670 -25342
rect 6646 -25884 6692 -25872
rect 7656 -25872 7670 -25844
rect 7704 -25342 7716 -25296
rect 8672 -25296 8732 -25156
rect 8970 -25212 9458 -25206
rect 8970 -25246 8982 -25212
rect 9446 -25246 9458 -25212
rect 8970 -25252 9458 -25246
rect 7704 -25844 7710 -25342
rect 8672 -25346 8688 -25296
rect 7704 -25872 7716 -25844
rect 5916 -25922 6404 -25916
rect 5916 -25956 5928 -25922
rect 6392 -25956 6404 -25922
rect 5916 -25962 6404 -25956
rect 6934 -25922 7422 -25916
rect 6934 -25956 6946 -25922
rect 7410 -25956 7422 -25922
rect 6934 -25962 7422 -25956
rect 6126 -26028 6186 -25962
rect 7148 -26028 7208 -25962
rect 7656 -26028 7716 -25872
rect 8682 -25872 8688 -25346
rect 8722 -25346 8732 -25296
rect 9688 -25296 9748 -25058
rect 10702 -25156 10708 -25096
rect 10768 -25156 10774 -25096
rect 9988 -25212 10476 -25206
rect 9988 -25246 10000 -25212
rect 10464 -25246 10476 -25212
rect 9988 -25252 10476 -25246
rect 8722 -25872 8728 -25346
rect 9688 -25352 9706 -25296
rect 9700 -25838 9706 -25352
rect 8682 -25884 8728 -25872
rect 9690 -25872 9706 -25838
rect 9740 -25352 9748 -25296
rect 10708 -25296 10768 -25156
rect 11006 -25212 11494 -25206
rect 11006 -25246 11018 -25212
rect 11482 -25246 11494 -25212
rect 11006 -25252 11494 -25246
rect 10708 -25344 10724 -25296
rect 9740 -25838 9746 -25352
rect 9740 -25872 9750 -25838
rect 7952 -25922 8440 -25916
rect 7952 -25956 7964 -25922
rect 8428 -25956 8440 -25922
rect 7952 -25962 8440 -25956
rect 8970 -25922 9458 -25916
rect 8970 -25956 8982 -25922
rect 9446 -25956 9458 -25922
rect 8970 -25962 9458 -25956
rect 8170 -26028 8230 -25962
rect 9180 -26028 9240 -25962
rect 9690 -26028 9750 -25872
rect 10718 -25872 10724 -25344
rect 10758 -25344 10768 -25296
rect 11726 -25296 11786 -25058
rect 12738 -25156 12744 -25096
rect 12804 -25156 12810 -25096
rect 12024 -25212 12512 -25206
rect 12024 -25246 12036 -25212
rect 12500 -25246 12512 -25212
rect 12024 -25252 12512 -25246
rect 11726 -25340 11742 -25296
rect 10758 -25872 10764 -25344
rect 11736 -25814 11742 -25340
rect 10718 -25884 10764 -25872
rect 11730 -25872 11742 -25814
rect 11776 -25340 11786 -25296
rect 12744 -25296 12804 -25156
rect 13042 -25212 13530 -25206
rect 13042 -25246 13054 -25212
rect 13518 -25246 13530 -25212
rect 13042 -25252 13530 -25246
rect 12744 -25338 12760 -25296
rect 11776 -25814 11782 -25340
rect 11776 -25872 11790 -25814
rect 9988 -25922 10476 -25916
rect 9988 -25956 10000 -25922
rect 10464 -25956 10476 -25922
rect 9988 -25962 10476 -25956
rect 11006 -25922 11494 -25916
rect 11006 -25956 11018 -25922
rect 11482 -25956 11494 -25922
rect 11006 -25962 11494 -25956
rect 10208 -26028 10268 -25962
rect 11226 -26028 11286 -25962
rect 11730 -26028 11790 -25872
rect 12754 -25872 12760 -25338
rect 12794 -25338 12804 -25296
rect 13760 -25296 13820 -25058
rect 14772 -25156 14778 -25096
rect 14838 -25156 14844 -25096
rect 14060 -25212 14548 -25206
rect 14060 -25246 14072 -25212
rect 14536 -25246 14548 -25212
rect 14060 -25252 14548 -25246
rect 12794 -25872 12800 -25338
rect 13760 -25352 13778 -25296
rect 13772 -25842 13778 -25352
rect 12754 -25884 12800 -25872
rect 13768 -25872 13778 -25842
rect 13812 -25352 13820 -25296
rect 14778 -25296 14838 -25156
rect 15078 -25212 15566 -25206
rect 15078 -25246 15090 -25212
rect 15554 -25246 15566 -25212
rect 15078 -25252 15566 -25246
rect 14778 -25338 14796 -25296
rect 13812 -25842 13818 -25352
rect 13812 -25872 13828 -25842
rect 12024 -25922 12512 -25916
rect 12024 -25956 12036 -25922
rect 12500 -25956 12512 -25922
rect 12024 -25962 12512 -25956
rect 13042 -25922 13530 -25916
rect 13042 -25956 13054 -25922
rect 13518 -25956 13530 -25922
rect 13042 -25962 13530 -25956
rect 12242 -26028 12302 -25962
rect 13264 -26028 13324 -25962
rect 13768 -26028 13828 -25872
rect 14790 -25872 14796 -25338
rect 14830 -25338 14838 -25296
rect 15800 -25296 15860 -25058
rect 16808 -25156 16814 -25096
rect 16874 -25156 16880 -25096
rect 16096 -25212 16584 -25206
rect 16096 -25246 16108 -25212
rect 16572 -25246 16584 -25212
rect 16096 -25252 16584 -25246
rect 14830 -25872 14836 -25338
rect 15800 -25342 15814 -25296
rect 15808 -25828 15814 -25342
rect 14790 -25884 14836 -25872
rect 15802 -25872 15814 -25828
rect 15848 -25342 15860 -25296
rect 16814 -25296 16874 -25156
rect 17114 -25212 17602 -25206
rect 17114 -25246 17126 -25212
rect 17590 -25246 17602 -25212
rect 17114 -25252 17602 -25246
rect 16814 -25342 16832 -25296
rect 15848 -25828 15854 -25342
rect 15848 -25872 15862 -25828
rect 14060 -25922 14548 -25916
rect 14060 -25956 14072 -25922
rect 14536 -25956 14548 -25922
rect 14060 -25962 14548 -25956
rect 15078 -25922 15566 -25916
rect 15078 -25956 15090 -25922
rect 15554 -25956 15566 -25922
rect 15078 -25962 15566 -25956
rect 14286 -26028 14346 -25962
rect 15294 -26028 15354 -25962
rect 15802 -26028 15862 -25872
rect 16826 -25872 16832 -25342
rect 16866 -25342 16874 -25296
rect 17834 -25296 17894 -25058
rect 18848 -25156 18854 -25096
rect 18914 -25156 18920 -25096
rect 18132 -25212 18620 -25206
rect 18132 -25246 18144 -25212
rect 18608 -25246 18620 -25212
rect 18132 -25252 18620 -25246
rect 16866 -25872 16872 -25342
rect 17834 -25354 17850 -25296
rect 17844 -25832 17850 -25354
rect 16826 -25884 16872 -25872
rect 17838 -25872 17850 -25832
rect 17884 -25354 17894 -25296
rect 18854 -25296 18914 -25156
rect 19150 -25212 19638 -25206
rect 19150 -25246 19162 -25212
rect 19626 -25246 19638 -25212
rect 19150 -25252 19638 -25246
rect 18854 -25328 18868 -25296
rect 17884 -25832 17890 -25354
rect 17884 -25872 17898 -25832
rect 16298 -25916 16358 -25914
rect 16096 -25922 16584 -25916
rect 16096 -25956 16108 -25922
rect 16572 -25956 16584 -25922
rect 16096 -25962 16584 -25956
rect 17114 -25922 17602 -25916
rect 17114 -25956 17126 -25922
rect 17590 -25956 17602 -25922
rect 17114 -25962 17602 -25956
rect 16298 -26028 16358 -25962
rect 17344 -26028 17404 -25962
rect 17838 -26028 17898 -25872
rect 18862 -25872 18868 -25328
rect 18902 -25328 18914 -25296
rect 19868 -25296 19928 -25058
rect 20366 -25206 20426 -24730
rect 20888 -25096 20948 -24640
rect 21906 -24640 21922 -24592
rect 21956 -24592 21962 -24064
rect 22934 -24064 22994 -23990
rect 21956 -24640 21966 -24592
rect 22934 -24606 22940 -24064
rect 21186 -24690 21674 -24684
rect 21186 -24724 21198 -24690
rect 21662 -24724 21674 -24690
rect 21186 -24730 21674 -24724
rect 20882 -25156 20888 -25096
rect 20948 -25156 20954 -25096
rect 20168 -25212 20656 -25206
rect 20168 -25246 20180 -25212
rect 20644 -25246 20656 -25212
rect 20168 -25252 20656 -25246
rect 18902 -25872 18908 -25328
rect 19868 -25338 19886 -25296
rect 19880 -25838 19886 -25338
rect 18862 -25884 18908 -25872
rect 19876 -25872 19886 -25838
rect 19920 -25338 19928 -25296
rect 20888 -25296 20948 -25156
rect 21394 -25206 21454 -24730
rect 21906 -24998 21966 -24640
rect 22924 -24640 22940 -24606
rect 22974 -24140 22994 -24064
rect 22974 -24606 22980 -24140
rect 22974 -24640 22984 -24606
rect 22204 -24690 22692 -24684
rect 22204 -24724 22216 -24690
rect 22680 -24724 22692 -24690
rect 22204 -24730 22692 -24724
rect 21900 -25058 21906 -24998
rect 21966 -25058 21972 -24998
rect 21186 -25212 21674 -25206
rect 21186 -25246 21198 -25212
rect 21662 -25246 21674 -25212
rect 21186 -25252 21674 -25246
rect 20888 -25336 20904 -25296
rect 19920 -25838 19926 -25338
rect 19920 -25872 19936 -25838
rect 18132 -25922 18620 -25916
rect 18132 -25956 18144 -25922
rect 18608 -25956 18620 -25922
rect 18132 -25962 18620 -25956
rect 19150 -25922 19638 -25916
rect 19150 -25956 19162 -25922
rect 19626 -25956 19638 -25922
rect 19150 -25962 19638 -25956
rect 18342 -26028 18402 -25962
rect 19354 -26028 19414 -25962
rect 19876 -26028 19936 -25872
rect 20898 -25872 20904 -25336
rect 20938 -25336 20948 -25296
rect 21906 -25296 21966 -25058
rect 22386 -25206 22446 -24730
rect 22924 -25096 22984 -24640
rect 23648 -24998 23708 -12606
rect 23800 -23926 23806 -23866
rect 23866 -23926 23872 -23866
rect 23642 -25058 23648 -24998
rect 23708 -25058 23714 -24998
rect 22918 -25156 22924 -25096
rect 22984 -25156 22990 -25096
rect 22204 -25212 22692 -25206
rect 22204 -25246 22216 -25212
rect 22680 -25246 22692 -25212
rect 22204 -25252 22692 -25246
rect 22386 -25254 22446 -25252
rect 21906 -25326 21922 -25296
rect 20938 -25872 20944 -25336
rect 21916 -25844 21922 -25326
rect 20898 -25884 20944 -25872
rect 21904 -25872 21922 -25844
rect 21956 -25326 21966 -25296
rect 22924 -25296 22984 -25156
rect 21956 -25844 21962 -25326
rect 22924 -25332 22940 -25296
rect 21956 -25872 21964 -25844
rect 20168 -25922 20656 -25916
rect 20168 -25956 20180 -25922
rect 20644 -25956 20656 -25922
rect 20168 -25962 20656 -25956
rect 21186 -25922 21674 -25916
rect 21186 -25956 21198 -25922
rect 21662 -25956 21674 -25922
rect 21186 -25962 21674 -25956
rect 20376 -26028 20436 -25962
rect 21442 -26028 21502 -25962
rect 21904 -26028 21964 -25872
rect 22934 -25872 22940 -25332
rect 22974 -25332 22984 -25296
rect 22974 -25872 22980 -25332
rect 22934 -25884 22980 -25872
rect 22204 -25922 22692 -25916
rect 22204 -25956 22216 -25922
rect 22680 -25956 22692 -25922
rect 22204 -25962 22692 -25956
rect 22404 -26028 22464 -25962
rect 3066 -26088 22464 -26028
rect 23806 -26430 23866 -23926
rect 24816 -26330 24822 -12070
rect 24922 -26330 24928 -12070
rect -7518 -26476 23968 -26430
rect -7518 -26630 -7472 -26476
rect 23928 -26630 23968 -26476
rect -7518 -26676 23968 -26630
rect -11616 -27116 -11606 -26816
rect 24206 -27116 24216 -26816
rect 24816 -27116 24928 -26330
rect -12328 -27122 24928 -27116
rect -12328 -27222 -12222 -27122
rect 24822 -27222 24928 -27122
rect -12328 -27228 24928 -27222
<< via1 >>
rect 484 1316 1084 1616
rect 24116 1316 24716 1616
rect 4061 1020 20846 1234
rect 4156 -4562 4216 -4502
rect 4268 -4562 4328 -4502
rect 4378 -4562 4438 -4502
rect 3492 -5274 3552 -5214
rect 3832 -5274 3892 -5214
rect 3942 -5274 4002 -5214
rect 2110 -6220 2170 -6160
rect 5028 -4562 5088 -4502
rect 5138 -4562 5198 -4502
rect 5246 -4562 5306 -4502
rect 4592 -5274 4652 -5214
rect 4704 -5274 4764 -5214
rect 4812 -5274 4872 -5214
rect 7986 824 8046 884
rect 9068 824 9128 884
rect 10026 824 10086 884
rect 8512 578 8572 638
rect 11062 824 11122 884
rect 12068 824 12128 884
rect 10548 578 10608 638
rect 11566 690 11626 750
rect 13090 824 13150 884
rect 14108 824 14168 884
rect 12586 580 12646 640
rect 15132 824 15192 884
rect 16144 824 16204 884
rect 14616 580 14676 640
rect 17162 824 17222 884
rect 18174 824 18234 884
rect 16658 582 16718 642
rect 17670 690 17730 750
rect 19202 824 19262 884
rect 20214 824 20274 884
rect 18690 582 18750 642
rect 21232 824 21292 884
rect 20726 582 20786 642
rect 6330 -354 6390 -294
rect 7494 -354 7554 -294
rect 6200 -558 6260 -498
rect 7494 -558 7554 -498
rect 9530 -458 9590 -398
rect 11566 -458 11626 -398
rect 13604 -354 13664 -294
rect 13600 -558 13660 -498
rect 15638 -354 15698 -294
rect 15636 -558 15696 -498
rect 17672 -458 17732 -398
rect 17814 -562 17874 -502
rect 19706 -458 19766 -398
rect 19708 -562 19768 -502
rect 21746 -354 21806 -294
rect 22884 -354 22944 -294
rect 8510 -1492 8570 -1432
rect 10546 -1492 10606 -1432
rect 9528 -1588 9588 -1528
rect 10232 -1594 10296 -1530
rect 11404 -1594 11468 -1530
rect 11566 -1698 11626 -1638
rect 12580 -1492 12640 -1432
rect 14618 -1494 14678 -1434
rect 15638 -1592 15698 -1532
rect 16654 -1494 16714 -1434
rect 17672 -1698 17732 -1638
rect 18690 -1494 18750 -1434
rect 19708 -1698 19768 -1638
rect 20724 -1496 20784 -1436
rect 21746 -1592 21806 -1532
rect 8510 -2630 8570 -2570
rect 9526 -2744 9590 -2680
rect 7488 -2882 7552 -2818
rect 6330 -3028 6390 -2968
rect 7312 -3028 7372 -2968
rect 6916 -3364 6976 -3304
rect 6048 -4562 6108 -4502
rect 5464 -5274 5524 -5214
rect 5574 -5274 5634 -5214
rect 4048 -5380 4108 -5320
rect 4484 -5380 4544 -5320
rect 4922 -5380 4982 -5320
rect 5356 -5380 5416 -5320
rect 4268 -5496 4328 -5436
rect 3832 -6220 3892 -6160
rect 4048 -6324 4108 -6264
rect 3942 -6422 4002 -6362
rect 4266 -6220 4326 -6160
rect 4156 -6422 4216 -6362
rect 3492 -7058 3552 -6998
rect 5138 -5496 5198 -5436
rect 4484 -6324 4544 -6264
rect 4376 -6422 4436 -6362
rect 3832 -7158 3892 -7098
rect 4702 -6220 4762 -6160
rect 4922 -6324 4982 -6264
rect 4594 -6422 4654 -6362
rect 4704 -6422 4764 -6362
rect 4810 -6422 4870 -6362
rect 5138 -6220 5198 -6160
rect 5028 -6422 5088 -6362
rect 5932 -5496 5992 -5436
rect 5356 -6324 5416 -6264
rect 5246 -6422 5306 -6362
rect 4702 -7158 4762 -7098
rect 5576 -6220 5636 -6160
rect 5462 -6422 5522 -6362
rect 5576 -7158 5636 -7098
rect 5932 -7158 5992 -7098
rect 4048 -7256 4108 -7196
rect 4484 -7256 4544 -7196
rect 4922 -7256 4982 -7196
rect 5356 -7256 5416 -7196
rect 3492 -7374 3552 -7314
rect 4158 -7374 4218 -7314
rect 4266 -7374 4326 -7314
rect 4374 -7374 4434 -7314
rect 5020 -7374 5080 -7314
rect 5138 -7374 5198 -7314
rect 5247 -7374 5305 -7316
rect 6802 -5668 6862 -5608
rect 10546 -2630 10606 -2570
rect 9526 -3178 9590 -3114
rect 7312 -3464 7372 -3404
rect 8478 -3464 8538 -3404
rect 7044 -4510 7104 -4450
rect 6916 -5772 6976 -5712
rect 3832 -8094 3892 -8034
rect 3942 -8094 4002 -8034
rect 4596 -8094 4656 -8034
rect 4702 -8094 4762 -8034
rect 4812 -8094 4872 -8034
rect 5464 -8094 5524 -8034
rect 5576 -8094 5636 -8034
rect 6048 -8094 6108 -8034
rect 7180 -4608 7240 -4548
rect 7044 -8182 7104 -8122
rect 12040 -2634 12100 -2574
rect 11564 -3364 11624 -3304
rect 10514 -3464 10574 -3404
rect 12580 -2572 12640 -2570
rect 12548 -2630 12640 -2572
rect 13040 -2630 13100 -2570
rect 12548 -2632 12608 -2630
rect 8482 -4718 8542 -4658
rect 9496 -4412 9556 -4352
rect 9496 -4608 9556 -4548
rect 10516 -4606 10576 -4546
rect 10516 -4718 10576 -4658
rect 14084 -2628 14144 -2568
rect 13598 -2882 13662 -2818
rect 13598 -3166 13662 -3102
rect 14586 -2572 14646 -2568
rect 14586 -2628 14678 -2572
rect 14618 -2632 14678 -2628
rect 15100 -2628 15160 -2568
rect 16128 -2628 16188 -2568
rect 15634 -2882 15698 -2818
rect 16654 -2574 16714 -2572
rect 16622 -2632 16714 -2574
rect 16622 -2634 16682 -2632
rect 17150 -2638 17210 -2578
rect 17638 -2634 17698 -2574
rect 18150 -2638 18210 -2578
rect 18690 -2634 18750 -2574
rect 20724 -2634 20784 -2574
rect 19706 -2744 19770 -2680
rect 21742 -2882 21806 -2818
rect 21714 -3158 21774 -3098
rect 22884 -3164 22944 -3104
rect 18660 -3464 18720 -3404
rect 20694 -3464 20754 -3404
rect 23138 -3464 23198 -3404
rect 11532 -4412 11592 -4352
rect 13572 -4720 13632 -4660
rect 15606 -4720 15666 -4660
rect 18662 -4720 18722 -4660
rect 19676 -4412 19736 -4352
rect 20696 -4720 20756 -4660
rect 21712 -4412 21772 -4352
rect 22978 -4606 23038 -4546
rect 9498 -5772 9558 -5712
rect 9498 -5976 9558 -5916
rect 11534 -5772 11594 -5712
rect 11532 -5874 11592 -5814
rect 11532 -5976 11592 -5916
rect 13568 -5668 13628 -5608
rect 14588 -5668 14648 -5608
rect 14588 -5974 14648 -5914
rect 15606 -5974 15666 -5914
rect 16624 -5668 16684 -5608
rect 16622 -5974 16682 -5914
rect 18658 -5772 18718 -5712
rect 19526 -5654 19586 -5594
rect 19674 -5764 19734 -5704
rect 19526 -5974 19586 -5914
rect 19678 -5972 19738 -5912
rect 20694 -5874 20754 -5814
rect 21714 -5764 21774 -5704
rect 22846 -5764 22906 -5704
rect 21712 -5972 21772 -5912
rect 8480 -6924 8540 -6864
rect 7312 -7132 7372 -7072
rect 9494 -7234 9554 -7174
rect 10516 -6924 10576 -6864
rect 10516 -7032 10576 -6972
rect 11528 -7234 11588 -7174
rect 11732 -7228 11792 -7168
rect 13570 -6922 13630 -6862
rect 15606 -6922 15666 -6862
rect 13566 -7228 13626 -7168
rect 14586 -7232 14646 -7172
rect 16620 -7232 16680 -7172
rect 16834 -7236 16894 -7176
rect 18660 -6920 18720 -6860
rect 19170 -7236 19230 -7176
rect 19682 -7234 19742 -7174
rect 20696 -6920 20756 -6860
rect 22978 -5972 23038 -5912
rect 22846 -7032 22906 -6972
rect 21716 -7234 21776 -7174
rect 8476 -8182 8536 -8122
rect 10512 -8182 10572 -8122
rect 7180 -8312 7240 -8252
rect 2110 -8452 2170 -8392
rect 1954 -8558 2014 -8498
rect 18664 -8182 18724 -8122
rect 20700 -8182 20760 -8122
rect 11534 -8452 11594 -8392
rect 23138 -8452 23198 -8392
rect 1184 -8676 1244 -8616
rect -5038 -11178 -4938 -11176
rect -2438 -11178 -2338 -11176
rect -634 -11178 -534 -11176
rect -12032 -11278 -11932 -11178
rect -10238 -11278 -10138 -11178
rect -7638 -11278 -7538 -11178
rect -5038 -11276 -4938 -11178
rect -2438 -11276 -2338 -11178
rect -634 -11276 -534 -11178
rect 1954 -11408 2014 -11348
rect 2110 -11408 2170 -11348
rect 1184 -12394 1244 -12334
rect 1850 -12508 1910 -12448
rect 2336 -11416 2396 -11356
rect 2112 -13848 2172 -13788
rect 1976 -14060 2036 -14000
rect 1850 -14962 1910 -14902
rect 690 -18948 750 -18888
rect -2976 -20220 -2916 -20160
rect -7386 -21660 -7326 -21600
rect -5346 -21660 -5286 -21600
rect -9538 -22564 -9478 -22504
rect -8400 -22564 -8340 -22504
rect -7386 -22660 -7326 -22600
rect -6364 -22776 -6304 -22716
rect -5346 -22660 -5286 -22600
rect -8254 -23676 -8194 -23616
rect -8402 -23784 -8342 -23724
rect -4326 -22564 -4266 -22504
rect -814 -19184 -754 -19124
rect 98 -19184 158 -19124
rect -1684 -19294 -1624 -19234
rect -2598 -19402 -2538 -19342
rect -2468 -19510 -2408 -19450
rect -920 -19402 -860 -19342
rect -1138 -19510 -1078 -19450
rect -2010 -20010 -1950 -19950
rect -1902 -20110 -1842 -20050
rect -1900 -20220 -1840 -20160
rect -1354 -20010 -1294 -19950
rect -1464 -20110 -1404 -20050
rect -1466 -20220 -1406 -20160
rect -1792 -20330 -1732 -20270
rect -1572 -20330 -1512 -20270
rect -2468 -20834 -2408 -20774
rect -2598 -20956 -2538 -20896
rect -2010 -20834 -1950 -20774
rect -1792 -20956 -1732 -20896
rect -2118 -21080 -2058 -21020
rect -22 -19294 38 -19234
rect -702 -19402 -642 -19342
rect -484 -19510 -424 -19450
rect -484 -20010 -424 -19950
rect -1138 -20220 -1078 -20160
rect -1028 -20220 -968 -20160
rect -592 -20220 -532 -20160
rect -918 -20330 -858 -20270
rect -702 -20330 -642 -20270
rect -1354 -20834 -1294 -20774
rect -1574 -20956 -1514 -20896
rect -1680 -21206 -1620 -21146
rect -22 -19784 38 -19724
rect -374 -20130 -314 -20070
rect -810 -20834 -750 -20774
rect -1138 -20954 -1078 -20894
rect -482 -20954 -422 -20894
rect -22 -20834 38 -20774
rect -1248 -21080 -1188 -21020
rect -376 -21080 -316 -21020
rect 220 -20010 280 -19950
rect 220 -20256 280 -20196
rect 98 -21206 158 -21146
rect -1346 -21312 -1294 -21260
rect 952 -18918 1012 -18858
rect -2670 -21640 -2610 -21580
rect -7384 -23896 -7324 -23836
rect -3202 -22776 -3142 -22716
rect -6368 -23676 -6308 -23616
rect -6366 -23784 -6306 -23724
rect -5346 -23896 -5286 -23836
rect -8400 -24880 -8340 -24820
rect -9538 -24986 -9478 -24926
rect -4498 -23676 -4438 -23616
rect -4330 -23784 -4270 -23724
rect -7382 -24778 -7322 -24718
rect -6366 -24986 -6306 -24926
rect -5352 -24778 -5292 -24718
rect -7896 -25930 -7836 -25870
rect -2122 -21540 -2062 -21480
rect -932 -21540 -872 -21480
rect 262 -21540 322 -21480
rect 952 -21540 1012 -21480
rect -1678 -21640 -1618 -21580
rect -1380 -21640 -1320 -21580
rect -2542 -22674 -2482 -22614
rect -2126 -22674 -2066 -22614
rect -484 -21640 -424 -21580
rect -188 -21640 -128 -21580
rect -1829 -22541 -1771 -22483
rect -1974 -22782 -1914 -22722
rect -1225 -22541 -1167 -22483
rect -1532 -22674 -1472 -22614
rect -1676 -22782 -1616 -22722
rect -1376 -22782 -1316 -22722
rect -2670 -23680 -2610 -23620
rect -4332 -24880 -4272 -24820
rect -3202 -24880 -3142 -24820
rect -6870 -25930 -6810 -25870
rect -5846 -25930 -5786 -25870
rect -1976 -23680 -1916 -23620
rect -934 -22674 -874 -22614
rect -1082 -22782 -1022 -22722
rect -634 -22541 -576 -22483
rect -786 -22782 -726 -22722
rect -37 -22541 21 -22483
rect -340 -22674 -280 -22614
rect -486 -22782 -426 -22722
rect -184 -22782 -124 -22722
rect -1530 -23788 -1470 -23728
rect 258 -22674 318 -22614
rect 106 -22782 166 -22722
rect 559 -22541 617 -22483
rect 410 -22782 470 -22722
rect -1080 -23680 -1020 -23620
rect -786 -23680 -726 -23620
rect -336 -23788 -276 -23728
rect -1828 -24772 -1768 -24712
rect -2426 -24866 -2366 -24806
rect -1978 -24974 -1918 -24914
rect -1534 -24866 -1474 -24806
rect -1680 -24974 -1620 -24914
rect -1234 -24772 -1174 -24712
rect -1384 -24974 -1324 -24914
rect 108 -23680 168 -23620
rect 410 -23680 470 -23620
rect -634 -24772 -574 -24712
rect -936 -24866 -876 -24806
rect -1080 -24974 -1020 -24914
rect -784 -24974 -724 -24914
rect -338 -24866 -278 -24806
rect -486 -24974 -426 -24914
rect 952 -23788 1012 -23728
rect -40 -24772 20 -24712
rect -190 -24974 -130 -24914
rect 554 -24772 614 -24712
rect 262 -24866 322 -24806
rect 106 -24974 166 -24914
rect 410 -24974 470 -24914
rect -4946 -25930 -4886 -25870
rect -2670 -25900 -2610 -25840
rect -1680 -25900 -1620 -25840
rect -1382 -25900 -1322 -25840
rect -486 -25900 -426 -25840
rect -184 -25900 -124 -25840
rect 1076 -22782 1136 -22722
rect 1976 -23604 2036 -23544
rect 2568 -12508 2628 -12448
rect 3586 -12606 3646 -12546
rect 4604 -12508 4664 -12448
rect 6638 -12508 6698 -12448
rect 8678 -12508 8738 -12448
rect 10714 -12508 10774 -12448
rect 12748 -12508 12808 -12448
rect 14784 -12508 14844 -12448
rect 16820 -12508 16880 -12448
rect 18856 -12508 18916 -12448
rect 5624 -12606 5684 -12546
rect 7658 -12606 7718 -12546
rect 9692 -12606 9752 -12546
rect 11732 -12606 11792 -12546
rect 13766 -12606 13826 -12546
rect 15804 -12606 15864 -12546
rect 17836 -12606 17896 -12546
rect 19874 -12606 19934 -12546
rect 11732 -12818 11792 -12758
rect 13764 -12818 13824 -12758
rect 6272 -13738 6332 -13678
rect 6642 -13738 6702 -13678
rect 7144 -13738 7204 -13678
rect 7656 -13738 7716 -13678
rect 8184 -13738 8244 -13678
rect 8676 -13738 8736 -13678
rect 4096 -13848 4156 -13788
rect 5118 -13848 5178 -13788
rect 2572 -14060 2632 -14000
rect 3070 -14060 3130 -14000
rect 3582 -14060 3642 -14000
rect 6138 -13952 6198 -13892
rect 5624 -14060 5684 -14000
rect 4086 -14962 4146 -14902
rect 2336 -15176 2396 -15116
rect 7138 -13952 7198 -13892
rect 8158 -13952 8218 -13892
rect 7658 -14060 7718 -14000
rect 5102 -14950 5162 -14890
rect 6122 -14950 6182 -14890
rect 4598 -15054 4658 -14994
rect 4604 -15288 4664 -15228
rect 5622 -15054 5682 -14994
rect 10708 -13738 10768 -13678
rect 9190 -13848 9250 -13788
rect 9694 -13848 9754 -13788
rect 10210 -13848 10270 -13788
rect 9692 -14060 9752 -14000
rect 7134 -14950 7194 -14890
rect 8160 -14950 8220 -14890
rect 6634 -15054 6694 -14994
rect 6640 -15288 6700 -15228
rect 7654 -15054 7714 -14994
rect 2448 -16218 2508 -16158
rect 3586 -16218 3646 -16158
rect 2336 -16418 2396 -16358
rect 2230 -16520 2290 -16460
rect 2336 -17654 2396 -17594
rect 2230 -20010 2290 -19950
rect 3584 -16418 3644 -16358
rect 4602 -16298 4662 -16238
rect 11230 -13848 11290 -13788
rect 11732 -13848 11792 -13788
rect 12232 -13848 12292 -13788
rect 11848 -14060 11908 -14000
rect 12744 -13738 12804 -13678
rect 12372 -13952 12432 -13892
rect 13258 -13848 13318 -13788
rect 13380 -13952 13440 -13892
rect 13768 -13848 13828 -13788
rect 14276 -13848 14336 -13788
rect 13572 -14062 13632 -14002
rect 14780 -13738 14840 -13678
rect 14422 -13952 14482 -13892
rect 16818 -13738 16878 -13678
rect 15284 -13848 15344 -13788
rect 15806 -13848 15866 -13788
rect 16296 -13848 16356 -13788
rect 15806 -14060 15866 -14000
rect 20894 -12508 20954 -12448
rect 21912 -12606 21972 -12546
rect 22924 -12508 22984 -12448
rect 23648 -12606 23708 -12546
rect 18342 -13738 18402 -13678
rect 18856 -13738 18916 -13678
rect 19364 -13738 19424 -13678
rect 17328 -13848 17388 -13788
rect 17840 -13848 17900 -13788
rect 17314 -13952 17374 -13892
rect 18352 -13952 18412 -13892
rect 17838 -14060 17898 -14000
rect 8676 -15054 8736 -14994
rect 10712 -15054 10772 -14994
rect 12750 -15054 12810 -14994
rect 14780 -15054 14840 -14994
rect 9696 -15176 9756 -15116
rect 11730 -15176 11790 -15116
rect 13760 -15176 13820 -15116
rect 5620 -16194 5680 -16134
rect 5116 -16412 5176 -16352
rect 6642 -16298 6702 -16238
rect 6120 -16412 6180 -16352
rect 3584 -17450 3644 -17390
rect 4090 -17552 4150 -17492
rect 7656 -16194 7716 -16134
rect 7132 -16412 7192 -16352
rect 8674 -16298 8734 -16238
rect 15800 -15054 15860 -14994
rect 8152 -16412 8212 -16352
rect 8674 -16410 8734 -16350
rect 10708 -16298 10768 -16238
rect 9692 -16520 9752 -16460
rect 5622 -17450 5682 -17390
rect 5620 -17654 5680 -17594
rect 10710 -16410 10770 -16350
rect 11726 -16520 11786 -16460
rect 20384 -13848 20444 -13788
rect 21404 -13848 21464 -13788
rect 19352 -13952 19412 -13892
rect 19870 -14060 19930 -14000
rect 21912 -14060 21972 -14000
rect 22416 -14060 22476 -14000
rect 22926 -14060 22986 -14000
rect 17316 -14950 17376 -14890
rect 18352 -14950 18412 -14890
rect 16818 -15054 16878 -14994
rect 17838 -15054 17898 -14994
rect 12748 -16298 12808 -16238
rect 12746 -16410 12806 -16350
rect 14782 -16298 14842 -16238
rect 14978 -16302 15038 -16242
rect 13766 -16520 13826 -16460
rect 14782 -16410 14842 -16350
rect 19368 -14950 19428 -14890
rect 18854 -15054 18914 -14994
rect 20890 -15054 20950 -14994
rect 15800 -16194 15860 -16134
rect 14978 -16520 15038 -16460
rect 15272 -16518 15332 -16458
rect 7658 -17450 7718 -17390
rect 4604 -17754 4664 -17694
rect 6128 -17660 6188 -17600
rect 7150 -17660 7210 -17600
rect 6638 -17754 6698 -17694
rect 9690 -17450 9750 -17390
rect 9182 -17552 9242 -17492
rect 8164 -17660 8224 -17600
rect 9182 -17660 9242 -17600
rect 8674 -17754 8734 -17694
rect 4086 -18678 4146 -18618
rect 4996 -18678 5056 -18618
rect 4086 -18894 4146 -18834
rect 2450 -18998 2510 -18938
rect 2336 -20256 2396 -20196
rect 2242 -21312 2294 -21260
rect 5998 -18678 6058 -18618
rect 5124 -18894 5184 -18834
rect 7150 -18678 7210 -18618
rect 6638 -18780 6698 -18720
rect 6138 -18894 6198 -18834
rect 4084 -19906 4144 -19846
rect 3586 -20010 3646 -19950
rect 3582 -20220 3642 -20160
rect 5092 -19906 5152 -19846
rect 4602 -20122 4662 -20062
rect 10202 -17660 10262 -17600
rect 16816 -16410 16876 -16350
rect 16300 -16518 16360 -16458
rect 16818 -16524 16878 -16464
rect 17836 -16194 17896 -16134
rect 18854 -16410 18914 -16350
rect 19870 -16302 19930 -16242
rect 20374 -16306 20434 -16246
rect 23034 -15288 23094 -15228
rect 20894 -16410 20954 -16350
rect 18854 -16524 18914 -16464
rect 14272 -17438 14332 -17378
rect 13766 -17566 13826 -17506
rect 15802 -17764 15862 -17704
rect 8160 -18678 8220 -18618
rect 9166 -18678 9226 -18618
rect 10210 -18678 10270 -18618
rect 10710 -18672 10770 -18612
rect 9164 -18894 9224 -18834
rect 10204 -18894 10264 -18834
rect 9688 -18998 9748 -18938
rect 6106 -19906 6166 -19846
rect 7144 -19906 7204 -19846
rect 6640 -20122 6700 -20062
rect 5620 -20220 5680 -20160
rect 11218 -18894 11278 -18834
rect 12746 -18672 12806 -18612
rect 12226 -18894 12286 -18834
rect 13270 -18894 13330 -18834
rect 11730 -18998 11790 -18938
rect 20892 -16524 20952 -16464
rect 17314 -17660 17374 -17600
rect 14782 -18672 14842 -18612
rect 14260 -18894 14320 -18834
rect 15278 -18894 15338 -18834
rect 13768 -18998 13828 -18938
rect 21910 -16194 21970 -16134
rect 22928 -16176 22988 -16116
rect 23528 -16306 23588 -16246
rect 23278 -16410 23338 -16350
rect 19366 -17438 19426 -17378
rect 19504 -17434 19564 -17374
rect 23034 -16524 23094 -16464
rect 20386 -17434 20446 -17374
rect 21392 -17434 21452 -17374
rect 18344 -17660 18404 -17600
rect 19504 -17660 19564 -17600
rect 19872 -17660 19932 -17600
rect 19872 -17764 19932 -17704
rect 21910 -17438 21970 -17378
rect 21910 -17566 21970 -17506
rect 20888 -17762 20948 -17702
rect 16820 -18672 16880 -18612
rect 16812 -18780 16872 -18720
rect 16312 -18894 16372 -18834
rect 15802 -18998 15862 -18938
rect 16314 -19002 16374 -18942
rect 17336 -19002 17396 -18942
rect 17836 -18996 17896 -18936
rect 8162 -19906 8222 -19846
rect 8678 -19900 8738 -19840
rect 10714 -19900 10774 -19840
rect 12746 -19900 12806 -19840
rect 14780 -19900 14840 -19840
rect 7660 -20220 7720 -20160
rect 2448 -21242 2508 -21182
rect 3588 -21458 3648 -21398
rect 4602 -21144 4662 -21084
rect 4606 -21338 4666 -21278
rect 5620 -21242 5680 -21182
rect 11730 -20010 11790 -19950
rect 13766 -20010 13826 -19950
rect 10712 -20122 10772 -20062
rect 9696 -20220 9756 -20160
rect 6638 -21144 6698 -21084
rect 7144 -21242 7204 -21182
rect 6642 -21338 6702 -21278
rect 8676 -21144 8736 -21084
rect 8166 -21242 8226 -21182
rect 7656 -21458 7716 -21398
rect 2336 -22374 2396 -22314
rect 9188 -21242 9248 -21182
rect 8670 -21338 8730 -21278
rect 18856 -18672 18916 -18612
rect 18852 -18780 18912 -18720
rect 19344 -18894 19404 -18834
rect 20894 -18672 20954 -18612
rect 20890 -18780 20950 -18720
rect 20382 -18894 20442 -18834
rect 19870 -18996 19930 -18936
rect 15802 -19898 15862 -19838
rect 16156 -19898 16216 -19838
rect 15798 -20010 15858 -19950
rect 15308 -20108 15368 -20048
rect 10538 -21124 10598 -21064
rect 10708 -21124 10768 -21064
rect 10192 -21242 10252 -21182
rect 9690 -21458 9750 -21398
rect 2230 -22500 2290 -22440
rect 5620 -22500 5680 -22440
rect 6140 -22488 6200 -22428
rect 4602 -22610 4662 -22550
rect 6638 -22610 6698 -22550
rect 6256 -22704 6316 -22644
rect 10538 -21338 10598 -21278
rect 10714 -21332 10774 -21272
rect 16346 -20108 16406 -20048
rect 17322 -20108 17382 -20048
rect 16156 -20216 16216 -20156
rect 21408 -18894 21468 -18834
rect 21912 -18996 21972 -18936
rect 19874 -19898 19934 -19838
rect 18338 -20108 18398 -20048
rect 20364 -20108 20424 -20048
rect 17836 -20220 17896 -20160
rect 19872 -20220 19932 -20160
rect 12750 -21124 12810 -21064
rect 14782 -21124 14842 -21064
rect 16822 -21124 16882 -21064
rect 15800 -21222 15860 -21162
rect 12742 -21332 12802 -21272
rect 7658 -22610 7718 -22550
rect 14786 -21332 14846 -21272
rect 8674 -22610 8734 -22550
rect 9694 -22610 9754 -22550
rect 7140 -22704 7200 -22644
rect 8162 -22704 8222 -22644
rect 2568 -23604 2628 -23544
rect 3082 -23604 3142 -23544
rect 3580 -23604 3640 -23544
rect 5622 -23604 5682 -23544
rect 6130 -23716 6190 -23656
rect 2110 -23822 2170 -23762
rect 4096 -23822 4156 -23762
rect 5118 -23822 5178 -23762
rect 16814 -21332 16874 -21272
rect 17840 -21458 17900 -21398
rect 21394 -20108 21454 -20048
rect 21908 -20220 21968 -20160
rect 18852 -21332 18912 -21272
rect 21906 -21222 21966 -21162
rect 20892 -21332 20952 -21272
rect 21410 -21328 21470 -21268
rect 19870 -21458 19930 -21398
rect 20396 -21456 20456 -21396
rect 11724 -22374 11784 -22314
rect 13766 -22374 13826 -22314
rect 15802 -22374 15862 -22314
rect 11220 -22488 11280 -22428
rect 16308 -22484 16368 -22424
rect 10712 -22610 10772 -22550
rect 12742 -22610 12802 -22550
rect 14780 -22610 14840 -22550
rect 16816 -22610 16876 -22550
rect 10204 -22704 10264 -22644
rect 7654 -23604 7714 -23544
rect 7142 -23716 7202 -23656
rect 8156 -23716 8216 -23656
rect 7656 -23822 7716 -23762
rect 8168 -23822 8228 -23762
rect 1704 -23926 1764 -23866
rect 6132 -23926 6192 -23866
rect 6636 -23926 6696 -23866
rect 7152 -23926 7212 -23866
rect 1076 -24974 1136 -24914
rect -2126 -26000 -2066 -25940
rect -938 -26000 -878 -25940
rect 258 -26000 318 -25940
rect 952 -26000 1012 -25940
rect 2568 -25156 2628 -25096
rect 3580 -25058 3640 -24998
rect 9686 -23604 9746 -23544
rect 9186 -23822 9246 -23762
rect 9692 -23822 9752 -23762
rect 10198 -23822 10258 -23762
rect 8674 -23926 8734 -23866
rect 4598 -25156 4658 -25096
rect 11068 -23716 11128 -23656
rect 10712 -23926 10772 -23866
rect 11590 -23604 11650 -23544
rect 11210 -23822 11270 -23762
rect 11728 -23714 11788 -23654
rect 12356 -23718 12416 -23658
rect 12230 -23822 12290 -23762
rect 13402 -23718 13462 -23658
rect 13252 -23822 13312 -23762
rect 12748 -23926 12808 -23866
rect 13950 -23602 14010 -23542
rect 13764 -23822 13824 -23762
rect 14270 -23822 14330 -23762
rect 21908 -21456 21968 -21396
rect 17838 -22610 17898 -22550
rect 18856 -22374 18916 -22314
rect 18858 -22610 18918 -22550
rect 17326 -22704 17386 -22644
rect 18346 -22704 18406 -22644
rect 15800 -23604 15860 -23544
rect 15288 -23822 15348 -23762
rect 15800 -23822 15860 -23762
rect 16308 -23822 16368 -23762
rect 14784 -23926 14844 -23866
rect 19872 -22610 19932 -22550
rect 20888 -22374 20948 -22314
rect 23162 -17438 23222 -17378
rect 23400 -17660 23460 -17600
rect 23278 -17762 23338 -17702
rect 23162 -18996 23222 -18936
rect 23158 -19898 23218 -19838
rect 23278 -21124 23338 -21064
rect 23158 -21222 23218 -21162
rect 23526 -18894 23586 -18834
rect 23528 -21328 23588 -21268
rect 23400 -21456 23460 -21396
rect 23034 -22374 23094 -22314
rect 21408 -22484 21468 -22424
rect 20894 -22610 20954 -22550
rect 19360 -22704 19420 -22644
rect 20396 -22704 20456 -22644
rect 17834 -23604 17894 -23544
rect 17330 -23718 17390 -23658
rect 18348 -23718 18408 -23658
rect 19868 -23604 19928 -23544
rect 19358 -23718 19418 -23658
rect 16816 -23926 16876 -23866
rect 17338 -23926 17398 -23866
rect 17838 -23926 17898 -23866
rect 18346 -23926 18406 -23866
rect 18854 -23926 18914 -23866
rect 19204 -23926 19264 -23866
rect 21910 -23604 21970 -23544
rect 22422 -23604 22482 -23544
rect 22928 -23604 22988 -23544
rect 20380 -23822 20440 -23762
rect 21382 -23822 21442 -23762
rect 11730 -24858 11790 -24798
rect 13766 -24858 13826 -24798
rect 5618 -25058 5678 -24998
rect 7656 -25058 7716 -24998
rect 9688 -25058 9748 -24998
rect 11726 -25058 11786 -24998
rect 13760 -25058 13820 -24998
rect 15800 -25058 15860 -24998
rect 17834 -25058 17894 -24998
rect 19868 -25058 19928 -24998
rect 6636 -25156 6696 -25096
rect 8672 -25156 8732 -25096
rect 10708 -25156 10768 -25096
rect 12744 -25156 12804 -25096
rect 14778 -25156 14838 -25096
rect 16814 -25156 16874 -25096
rect 18854 -25156 18914 -25096
rect 20888 -25156 20948 -25096
rect 21906 -25058 21966 -24998
rect 23806 -23926 23866 -23866
rect 23648 -25058 23708 -24998
rect 22924 -25156 22984 -25096
rect -7472 -26630 23928 -26476
rect -12216 -27116 -11616 -26816
rect 24216 -27116 24816 -26816
<< metal2 >>
rect 484 1616 1084 1626
rect 484 1306 1084 1316
rect 24116 1616 24716 1626
rect 24116 1306 24716 1316
rect 3998 1234 20878 1266
rect 3998 1020 4061 1234
rect 20846 1020 20878 1234
rect 3998 1000 20878 1020
rect 3998 998 8352 1000
rect 7986 884 8046 890
rect 9068 884 9128 890
rect 10026 884 10086 890
rect 11062 884 11122 890
rect 12068 884 12128 890
rect 13090 884 13150 890
rect 14108 884 14168 890
rect 15132 884 15192 890
rect 16144 884 16204 890
rect 17162 884 17222 890
rect 18174 884 18234 890
rect 19202 884 19262 890
rect 20214 884 20274 890
rect 21232 884 21292 890
rect 8046 824 9068 884
rect 9128 824 10026 884
rect 10086 824 11062 884
rect 11122 824 12068 884
rect 12128 824 13090 884
rect 13150 824 14108 884
rect 14168 824 15132 884
rect 15192 824 16144 884
rect 16204 824 17162 884
rect 17222 824 18174 884
rect 18234 824 19202 884
rect 19262 824 20214 884
rect 20274 824 21232 884
rect 7986 818 8046 824
rect 9068 818 9128 824
rect 10026 818 10086 824
rect 11062 818 11122 824
rect 12068 818 12128 824
rect 13090 818 13150 824
rect 14108 818 14168 824
rect 15132 818 15192 824
rect 16144 818 16204 824
rect 17162 818 17222 824
rect 18174 818 18234 824
rect 19202 818 19262 824
rect 20214 818 20274 824
rect 21232 818 21292 824
rect 11566 750 11626 756
rect 17670 750 17730 756
rect 11626 690 17670 750
rect 11566 684 11626 690
rect 17670 684 17730 690
rect 8512 638 8572 644
rect 10548 638 10608 644
rect 12586 640 12646 646
rect 14616 640 14676 646
rect 16658 642 16718 648
rect 18690 642 18750 648
rect 20726 642 20786 648
rect 8572 578 10548 638
rect 10608 580 12586 638
rect 12646 580 14616 640
rect 14676 582 16658 640
rect 16718 582 18690 642
rect 18750 582 20726 642
rect 14676 580 16856 582
rect 10608 578 12768 580
rect 8512 572 8572 578
rect 10548 572 10608 578
rect 12586 574 12646 578
rect 14616 574 14676 580
rect 16658 576 16718 580
rect 18690 576 18750 582
rect 20726 576 20786 582
rect 6330 -294 6390 -288
rect 7494 -294 7554 -288
rect 13604 -294 13664 -288
rect 6390 -354 7494 -294
rect 7554 -354 13604 -294
rect 6330 -360 6390 -354
rect 7494 -360 7554 -354
rect 13604 -360 13664 -354
rect 15638 -294 15698 -288
rect 21746 -294 21806 -288
rect 22884 -294 22944 -288
rect 15698 -354 21746 -294
rect 21806 -354 22884 -294
rect 15638 -360 15698 -354
rect 21746 -360 21806 -354
rect 22884 -360 22944 -354
rect 9530 -398 9590 -392
rect 11566 -398 11626 -392
rect 17672 -398 17732 -392
rect 19706 -398 19766 -392
rect 9590 -458 11566 -398
rect 11626 -406 12044 -398
rect 12260 -406 17672 -398
rect 11626 -452 17672 -406
rect 11626 -456 14060 -452
rect 11626 -458 13034 -456
rect 13272 -458 14060 -456
rect 14276 -458 17672 -452
rect 17732 -458 19706 -398
rect 9530 -464 9590 -458
rect 11566 -464 11626 -458
rect 17672 -464 17732 -458
rect 19706 -464 19766 -458
rect 6200 -498 6260 -492
rect 7494 -498 7554 -492
rect 13600 -498 13660 -492
rect 15636 -498 15696 -492
rect 6260 -558 7494 -498
rect 7554 -558 13600 -498
rect 13660 -558 15636 -498
rect 6200 -564 6260 -558
rect 7494 -564 7554 -558
rect 13600 -564 13660 -558
rect 15636 -564 15696 -558
rect 17814 -502 17874 -496
rect 19708 -502 19768 -496
rect 17874 -562 19708 -502
rect 17814 -568 17874 -562
rect 19708 -568 19768 -562
rect 8510 -1432 8570 -1426
rect 10546 -1432 10606 -1426
rect 12580 -1432 12640 -1426
rect 14618 -1432 14678 -1428
rect 8570 -1492 10546 -1432
rect 10606 -1492 12580 -1432
rect 12640 -1434 14822 -1432
rect 16654 -1434 16714 -1428
rect 18690 -1434 18750 -1428
rect 12640 -1492 14618 -1434
rect 8510 -1498 8570 -1492
rect 10546 -1498 10606 -1492
rect 12580 -1498 12640 -1492
rect 14678 -1494 16654 -1434
rect 16714 -1494 18690 -1434
rect 18750 -1436 19560 -1434
rect 20724 -1436 20784 -1430
rect 18750 -1494 20724 -1436
rect 14618 -1500 14678 -1494
rect 16654 -1500 16714 -1494
rect 18589 -1496 19104 -1494
rect 19354 -1496 20724 -1494
rect 18690 -1500 18750 -1496
rect 20724 -1502 20784 -1496
rect 9528 -1528 9588 -1522
rect 9588 -1588 10100 -1528
rect 9528 -1594 9588 -1588
rect 10040 -1638 10100 -1588
rect 10232 -1530 10296 -1524
rect 11404 -1530 11468 -1524
rect 10296 -1594 11404 -1530
rect 10232 -1600 10296 -1594
rect 11404 -1600 11468 -1594
rect 15638 -1532 15698 -1526
rect 21746 -1532 21806 -1526
rect 15698 -1592 21746 -1532
rect 15638 -1598 15698 -1592
rect 21746 -1598 21806 -1592
rect 11566 -1638 11626 -1632
rect 17672 -1638 17732 -1632
rect 19708 -1638 19768 -1632
rect 10040 -1698 11566 -1638
rect 11626 -1698 17672 -1638
rect 17732 -1698 19708 -1638
rect 11566 -1704 11626 -1698
rect 17672 -1704 17732 -1698
rect 19708 -1704 19768 -1698
rect 8510 -2570 8570 -2564
rect 10546 -2570 10606 -2564
rect 12580 -2570 12640 -2564
rect 13040 -2570 13100 -2564
rect 14618 -2568 14678 -2566
rect 14078 -2570 14084 -2568
rect 8570 -2630 10546 -2570
rect 10606 -2572 12580 -2570
rect 10606 -2574 12548 -2572
rect 10606 -2630 12040 -2574
rect 8510 -2636 8570 -2630
rect 10546 -2636 10606 -2630
rect 12034 -2634 12040 -2630
rect 12100 -2630 12548 -2574
rect 12640 -2630 13040 -2570
rect 13100 -2628 14084 -2570
rect 14144 -2570 14150 -2568
rect 14580 -2570 14586 -2568
rect 14144 -2628 14586 -2570
rect 14646 -2570 14678 -2568
rect 15094 -2570 15100 -2568
rect 14646 -2572 15100 -2570
rect 14678 -2628 15100 -2572
rect 15160 -2570 15166 -2568
rect 16122 -2570 16128 -2568
rect 15160 -2628 16128 -2570
rect 16188 -2570 16194 -2568
rect 16188 -2572 16500 -2570
rect 16654 -2572 16714 -2566
rect 18690 -2572 18750 -2568
rect 16188 -2574 16654 -2572
rect 16714 -2574 18878 -2572
rect 20724 -2574 20784 -2568
rect 16188 -2628 16622 -2574
rect 13100 -2630 14618 -2628
rect 12100 -2634 12106 -2630
rect 12542 -2632 12548 -2630
rect 12608 -2632 12640 -2630
rect 12580 -2636 12640 -2632
rect 13040 -2636 13100 -2630
rect 14678 -2630 16622 -2628
rect 14678 -2632 15066 -2630
rect 15272 -2632 16086 -2630
rect 16292 -2632 16622 -2630
rect 16714 -2578 17638 -2574
rect 16714 -2632 17150 -2578
rect 14618 -2638 14678 -2632
rect 16616 -2634 16622 -2632
rect 16682 -2634 16714 -2632
rect 16654 -2638 16714 -2634
rect 17144 -2638 17150 -2632
rect 17210 -2632 17638 -2578
rect 17210 -2638 17216 -2632
rect 17632 -2634 17638 -2632
rect 17698 -2578 18690 -2574
rect 17698 -2632 18150 -2578
rect 17698 -2634 17704 -2632
rect 18144 -2638 18150 -2632
rect 18210 -2632 18690 -2578
rect 18210 -2638 18216 -2632
rect 18750 -2634 20724 -2574
rect 18690 -2640 18750 -2634
rect 20724 -2640 20784 -2634
rect 9526 -2680 9590 -2674
rect 19706 -2680 19770 -2674
rect 9590 -2744 19706 -2680
rect 19770 -2744 23354 -2680
rect 9526 -2750 9590 -2744
rect 19706 -2750 19770 -2744
rect 7488 -2818 7552 -2812
rect 13598 -2818 13662 -2812
rect 7552 -2882 13598 -2818
rect 7488 -2888 7552 -2882
rect 13598 -2888 13662 -2882
rect 15634 -2818 15698 -2812
rect 21742 -2818 21806 -2812
rect 15698 -2826 18074 -2818
rect 18456 -2826 21742 -2818
rect 15698 -2882 21742 -2826
rect 15634 -2888 15698 -2882
rect 6330 -2968 6390 -2962
rect 15838 -2968 15898 -2882
rect 21742 -2888 21806 -2882
rect 6390 -3028 7312 -2968
rect 7372 -3028 15898 -2968
rect 6330 -3034 6390 -3028
rect 21708 -3100 21714 -3098
rect 13598 -3102 21714 -3100
rect 9526 -3114 9590 -3108
rect 690 -3178 9526 -3114
rect 13592 -3166 13598 -3102
rect 13662 -3158 21714 -3102
rect 21774 -3100 21780 -3098
rect 21774 -3104 22944 -3100
rect 21774 -3158 22884 -3104
rect 13662 -3164 22884 -3158
rect 22944 -3164 22950 -3104
rect 13662 -3166 13668 -3164
rect -12032 -11178 -11932 -11172
rect -10238 -11178 -10138 -11172
rect -7638 -11178 -7538 -11172
rect -5038 -11176 -4938 -11170
rect -2438 -11176 -2338 -11170
rect -634 -11176 -534 -11170
rect -12036 -11273 -12032 -11183
rect -11932 -11273 -11928 -11183
rect -10242 -11273 -10238 -11183
rect -10138 -11273 -10134 -11183
rect -7642 -11273 -7638 -11183
rect -7538 -11273 -7534 -11183
rect -5042 -11271 -5038 -11181
rect -4938 -11271 -4934 -11181
rect -2442 -11271 -2438 -11181
rect -2338 -11271 -2334 -11181
rect -638 -11271 -634 -11181
rect -534 -11271 -530 -11181
rect -12032 -11284 -11932 -11278
rect -10238 -11284 -10138 -11278
rect -7638 -11284 -7538 -11278
rect -5038 -11282 -4938 -11276
rect -2438 -11282 -2338 -11276
rect -634 -11282 -534 -11276
rect 690 -18888 750 -3178
rect 9526 -3184 9590 -3178
rect 11564 -3304 11624 -3298
rect 952 -3364 6916 -3304
rect 6976 -3364 11564 -3304
rect 952 -18858 1012 -3364
rect 11564 -3370 11624 -3364
rect 7312 -3404 7372 -3398
rect 8478 -3404 8538 -3398
rect 10514 -3404 10574 -3398
rect 7372 -3464 8478 -3404
rect 8538 -3464 10514 -3404
rect 7312 -3470 7372 -3464
rect 8478 -3470 8538 -3464
rect 10514 -3470 10574 -3464
rect 18660 -3404 18720 -3398
rect 20694 -3404 20754 -3398
rect 23138 -3404 23198 -3398
rect 18720 -3464 20694 -3404
rect 20754 -3464 23138 -3404
rect 18660 -3470 18720 -3464
rect 20694 -3470 20754 -3464
rect 23138 -3470 23198 -3464
rect 9496 -4352 9556 -4346
rect 11532 -4352 11592 -4346
rect 9556 -4412 11532 -4352
rect 9496 -4418 9556 -4412
rect 11532 -4418 11592 -4412
rect 19676 -4352 19736 -4346
rect 21712 -4352 21772 -4346
rect 19736 -4412 21712 -4352
rect 19676 -4418 19736 -4412
rect 7044 -4450 7104 -4444
rect 19784 -4450 19844 -4412
rect 21712 -4418 21772 -4412
rect 4156 -4502 4216 -4496
rect 4268 -4502 4328 -4496
rect 4378 -4502 4438 -4496
rect 5028 -4502 5088 -4496
rect 5138 -4502 5198 -4496
rect 5246 -4502 5306 -4496
rect 6048 -4502 6108 -4496
rect 1330 -4562 4156 -4502
rect 4216 -4562 4268 -4502
rect 4328 -4562 4378 -4502
rect 4438 -4562 5028 -4502
rect 5088 -4562 5138 -4502
rect 5198 -4562 5246 -4502
rect 5306 -4562 6048 -4502
rect 7104 -4510 19844 -4450
rect 7044 -4516 7104 -4510
rect 1178 -8676 1184 -8616
rect 1244 -8676 1250 -8616
rect 1184 -12334 1244 -8676
rect 1178 -12394 1184 -12334
rect 1244 -12394 1250 -12334
rect 684 -18948 690 -18888
rect 750 -18948 756 -18888
rect 946 -18918 952 -18858
rect 1012 -18918 1018 -18858
rect -814 -19124 -754 -19118
rect 98 -19124 158 -19118
rect 1330 -19124 1390 -4562
rect 4156 -4568 4216 -4562
rect 4268 -4568 4328 -4562
rect 4378 -4568 4438 -4562
rect 5028 -4568 5088 -4562
rect 5138 -4568 5198 -4562
rect 5246 -4568 5306 -4562
rect 6048 -4568 6108 -4562
rect 7180 -4548 7240 -4542
rect 9496 -4548 9556 -4542
rect 7240 -4608 9496 -4548
rect 7180 -4614 7240 -4608
rect 9496 -4614 9556 -4608
rect 10516 -4546 10576 -4540
rect 22978 -4546 23038 -4540
rect 10576 -4606 22978 -4546
rect 10516 -4612 10576 -4606
rect 22978 -4612 23038 -4606
rect 8482 -4658 8542 -4652
rect 10516 -4658 10576 -4652
rect 8542 -4718 10516 -4658
rect 8482 -4724 8542 -4718
rect 10516 -4724 10576 -4718
rect 13572 -4660 13632 -4654
rect 15606 -4660 15666 -4654
rect 13632 -4720 15606 -4660
rect 13572 -4726 13632 -4720
rect 15606 -4726 15666 -4720
rect 18662 -4660 18722 -4654
rect 20696 -4658 20756 -4654
rect 23290 -4658 23354 -2744
rect 20628 -4660 23354 -4658
rect 18722 -4720 20696 -4660
rect 20756 -4720 23354 -4660
rect 18662 -4726 18722 -4720
rect 20628 -4722 23354 -4720
rect 20696 -4726 20756 -4722
rect 3492 -5214 3552 -5208
rect 3832 -5214 3892 -5208
rect 3942 -5214 4002 -5208
rect 4592 -5214 4652 -5208
rect 4704 -5214 4764 -5208
rect 4812 -5214 4872 -5208
rect 5464 -5214 5524 -5208
rect 5574 -5214 5634 -5208
rect 3552 -5274 3832 -5214
rect 3892 -5274 3942 -5214
rect 4002 -5274 4592 -5214
rect 4652 -5274 4704 -5214
rect 4764 -5274 4812 -5214
rect 4872 -5274 5464 -5214
rect 5524 -5274 5574 -5214
rect 3492 -5280 3552 -5274
rect 3832 -5280 3892 -5274
rect 3942 -5280 4002 -5274
rect 4592 -5280 4652 -5274
rect 4704 -5280 4764 -5274
rect 4812 -5280 4872 -5274
rect 5464 -5280 5524 -5274
rect 5574 -5280 5634 -5274
rect 4048 -5320 4108 -5314
rect 4484 -5320 4544 -5314
rect 4922 -5320 4982 -5314
rect 5356 -5320 5416 -5314
rect 4108 -5380 4484 -5320
rect 4544 -5380 4922 -5320
rect 4982 -5380 5356 -5320
rect 4048 -5386 4108 -5380
rect 4484 -5386 4544 -5380
rect 4922 -5386 4982 -5380
rect 5356 -5386 5416 -5380
rect 4268 -5436 4328 -5430
rect 5138 -5436 5198 -5430
rect 5932 -5436 5992 -5430
rect 4328 -5496 5138 -5436
rect 5198 -5496 5932 -5436
rect 4268 -5502 4328 -5496
rect 5138 -5502 5198 -5496
rect 5932 -5502 5992 -5496
rect 19526 -5594 19586 -5588
rect 6802 -5608 6862 -5602
rect 13568 -5608 13628 -5602
rect 14588 -5608 14648 -5602
rect 16624 -5608 16684 -5602
rect 6862 -5668 13568 -5608
rect 13628 -5668 14588 -5608
rect 14648 -5668 16624 -5608
rect 19586 -5654 23948 -5594
rect 19526 -5660 19586 -5654
rect 6802 -5674 6862 -5668
rect 13568 -5674 13628 -5668
rect 14588 -5674 14648 -5668
rect 16624 -5674 16684 -5668
rect 19674 -5704 19734 -5698
rect 21714 -5704 21774 -5698
rect 22846 -5704 22906 -5698
rect 6916 -5712 6976 -5706
rect 11534 -5712 11594 -5706
rect 18658 -5712 18718 -5706
rect 6976 -5772 9498 -5712
rect 9558 -5772 11534 -5712
rect 11594 -5772 18658 -5712
rect 19734 -5764 21714 -5704
rect 21774 -5764 22846 -5704
rect 19674 -5770 19734 -5764
rect 21714 -5770 21774 -5764
rect 22846 -5770 22906 -5764
rect 6916 -5778 6976 -5772
rect 11534 -5778 11594 -5772
rect 18658 -5778 18718 -5772
rect 11532 -5814 11592 -5808
rect 20694 -5814 20754 -5808
rect 11592 -5874 20694 -5814
rect 11532 -5880 11592 -5874
rect 20694 -5880 20754 -5874
rect 9498 -5916 9558 -5910
rect 11532 -5916 11592 -5910
rect 9558 -5976 11532 -5916
rect 9498 -5982 9558 -5976
rect 11532 -5982 11592 -5976
rect 14588 -5914 14648 -5908
rect 15606 -5914 15666 -5908
rect 16622 -5914 16682 -5908
rect 19526 -5914 19586 -5908
rect 14648 -5974 15606 -5914
rect 15666 -5974 16622 -5914
rect 16682 -5974 19526 -5914
rect 14588 -5980 14648 -5974
rect 15606 -5980 15666 -5974
rect 16622 -5980 16682 -5974
rect 19526 -5980 19586 -5974
rect 19678 -5912 19738 -5906
rect 21712 -5912 21772 -5906
rect 22978 -5912 23038 -5906
rect 19738 -5972 21712 -5912
rect 21772 -5972 22978 -5912
rect 23038 -5972 23820 -5912
rect 19678 -5978 19738 -5972
rect 21712 -5978 21772 -5972
rect 22978 -5978 23038 -5972
rect 2110 -6160 2170 -6154
rect 3832 -6160 3892 -6154
rect 4266 -6160 4326 -6154
rect 4702 -6160 4762 -6154
rect 5138 -6160 5198 -6154
rect 5576 -6160 5636 -6154
rect 2170 -6220 3832 -6160
rect 3892 -6220 4266 -6160
rect 4326 -6220 4702 -6160
rect 4762 -6220 5138 -6160
rect 5198 -6220 5576 -6160
rect 2110 -6226 2170 -6220
rect 3832 -6226 3892 -6220
rect 4266 -6226 4326 -6220
rect 4702 -6226 4762 -6220
rect 5138 -6226 5198 -6220
rect 5576 -6226 5636 -6220
rect 4048 -6264 4108 -6258
rect 4484 -6264 4544 -6258
rect 4922 -6264 4982 -6258
rect 5356 -6264 5416 -6258
rect 4108 -6324 4484 -6264
rect 4544 -6324 4922 -6264
rect 4982 -6324 5356 -6264
rect 4048 -6330 4108 -6324
rect 4484 -6330 4544 -6324
rect 4922 -6330 4982 -6324
rect 5356 -6330 5416 -6324
rect 3942 -6362 4002 -6356
rect 4156 -6362 4216 -6356
rect 4376 -6362 4436 -6356
rect 4594 -6362 4654 -6356
rect 4704 -6362 4764 -6356
rect 4810 -6362 4870 -6356
rect 5028 -6362 5088 -6356
rect 5246 -6362 5306 -6356
rect 5462 -6362 5522 -6356
rect 4002 -6422 4156 -6362
rect 4216 -6422 4376 -6362
rect 4436 -6422 4594 -6362
rect 4654 -6422 4704 -6362
rect 4764 -6422 4810 -6362
rect 4870 -6422 5028 -6362
rect 5088 -6422 5246 -6362
rect 5306 -6422 5462 -6362
rect 3942 -6428 4002 -6422
rect 4156 -6428 4216 -6422
rect 4376 -6428 4436 -6422
rect 4594 -6428 4654 -6422
rect 4704 -6428 4764 -6422
rect 4810 -6428 4870 -6422
rect 5028 -6428 5088 -6422
rect 5246 -6428 5306 -6422
rect 5462 -6428 5522 -6422
rect 8480 -6864 8540 -6858
rect 10516 -6864 10576 -6858
rect 6914 -6924 8480 -6864
rect 8540 -6924 10516 -6864
rect -754 -19184 98 -19124
rect 158 -19184 1390 -19124
rect 1468 -7058 3492 -6998
rect 3552 -7058 3558 -6998
rect -814 -19190 -754 -19184
rect 98 -19190 158 -19184
rect -1684 -19234 -1624 -19228
rect -22 -19234 38 -19228
rect -1624 -19294 -22 -19234
rect -1684 -19300 -1624 -19294
rect -22 -19300 38 -19294
rect -2598 -19342 -2538 -19336
rect -920 -19342 -860 -19336
rect -702 -19342 -642 -19336
rect -2538 -19402 -920 -19342
rect -860 -19402 -702 -19342
rect -2598 -19408 -2538 -19402
rect -920 -19408 -860 -19402
rect -702 -19408 -642 -19402
rect -2468 -19450 -2408 -19444
rect -1138 -19450 -1078 -19444
rect -484 -19450 -424 -19444
rect -2408 -19510 -1138 -19450
rect -1078 -19510 -484 -19450
rect -2468 -19516 -2408 -19510
rect -1138 -19516 -1078 -19510
rect -484 -19516 -424 -19510
rect 1468 -19724 1528 -7058
rect 3832 -7098 3892 -7092
rect 4702 -7098 4762 -7092
rect 5576 -7098 5636 -7092
rect 5932 -7098 5992 -7092
rect -28 -19784 -22 -19724
rect 38 -19784 1528 -19724
rect 1586 -7158 3832 -7098
rect 3892 -7158 4702 -7098
rect 4762 -7158 5576 -7098
rect 5636 -7158 5932 -7098
rect -2010 -19950 -1950 -19944
rect -1354 -19950 -1294 -19944
rect -484 -19950 -424 -19944
rect 220 -19950 280 -19944
rect -1950 -20010 -1354 -19950
rect -1294 -20010 -484 -19950
rect -424 -20010 220 -19950
rect -2010 -20016 -1950 -20010
rect -1354 -20016 -1294 -20010
rect -484 -20016 -424 -20010
rect 220 -20016 280 -20010
rect -1902 -20050 -1842 -20044
rect -1464 -20050 -1404 -20044
rect -3096 -20110 -1902 -20050
rect -1842 -20110 -1464 -20050
rect -1404 -20110 -968 -20050
rect -7386 -21600 -7326 -21594
rect -5346 -21600 -5286 -21594
rect -7326 -21660 -5346 -21600
rect -7386 -21666 -7326 -21660
rect -5346 -21666 -5286 -21660
rect -9538 -22504 -9478 -22498
rect -8400 -22504 -8340 -22498
rect -4326 -22504 -4266 -22498
rect -9478 -22564 -8400 -22504
rect -8340 -22564 -4326 -22504
rect -9538 -22570 -9478 -22564
rect -8400 -22570 -8340 -22564
rect -4326 -22570 -4266 -22564
rect -7386 -22600 -7326 -22594
rect -5346 -22600 -5286 -22594
rect -7326 -22660 -5346 -22600
rect -7386 -22666 -7326 -22660
rect -5346 -22666 -5286 -22660
rect -6364 -22716 -6304 -22710
rect -3202 -22716 -3142 -22710
rect -6304 -22776 -3202 -22716
rect -6364 -22782 -6304 -22776
rect -3202 -22782 -3142 -22776
rect -8254 -23616 -8194 -23610
rect -6368 -23616 -6308 -23610
rect -4498 -23616 -4438 -23610
rect -3096 -23616 -3036 -20110
rect -1902 -20116 -1842 -20110
rect -1464 -20116 -1404 -20110
rect -2976 -20160 -2916 -20154
rect -1900 -20160 -1840 -20154
rect -1466 -20160 -1406 -20154
rect -1138 -20160 -1078 -20154
rect -2916 -20220 -1900 -20160
rect -1840 -20220 -1466 -20160
rect -1406 -20220 -1138 -20160
rect -2976 -20226 -2916 -20220
rect -1900 -20226 -1840 -20220
rect -1466 -20226 -1406 -20220
rect -1138 -20226 -1078 -20220
rect -1028 -20160 -968 -20110
rect -374 -20070 -314 -20064
rect 1586 -20070 1646 -7158
rect 3832 -7164 3892 -7158
rect 4702 -7164 4762 -7158
rect 5576 -7164 5636 -7158
rect 5932 -7164 5992 -7158
rect 4048 -7196 4108 -7190
rect 4484 -7196 4544 -7190
rect 4922 -7196 4982 -7190
rect 5356 -7196 5416 -7190
rect 4108 -7256 4484 -7196
rect 4544 -7256 4922 -7196
rect 4982 -7256 5356 -7196
rect 4048 -7262 4108 -7256
rect 4484 -7262 4544 -7256
rect 4922 -7262 4982 -7256
rect 5356 -7262 5416 -7256
rect 3492 -7314 3552 -7308
rect 4158 -7314 4218 -7308
rect 4266 -7314 4326 -7308
rect 4374 -7314 4434 -7308
rect 5020 -7314 5080 -7308
rect 5138 -7314 5198 -7308
rect 3552 -7374 4158 -7314
rect 4218 -7374 4266 -7314
rect 4326 -7374 4374 -7314
rect 4434 -7374 5020 -7314
rect 5080 -7374 5138 -7314
rect 5247 -7316 5305 -7310
rect 5198 -7374 5247 -7316
rect 3492 -7380 3552 -7374
rect 4158 -7380 4218 -7374
rect 4266 -7380 4326 -7374
rect 4374 -7380 4434 -7374
rect 5020 -7380 5080 -7374
rect 5138 -7380 5198 -7374
rect 5247 -7380 5305 -7374
rect 2318 -7717 2327 -7627
rect 2417 -7717 2426 -7627
rect 2110 -8392 2170 -8386
rect 1948 -8558 1954 -8498
rect 2014 -8558 2020 -8498
rect 1696 -10213 1705 -10123
rect 1795 -10213 1804 -10123
rect 1720 -11476 1780 -10213
rect 1954 -11348 2014 -8558
rect 1954 -11414 2014 -11408
rect 2110 -11348 2170 -8452
rect 2336 -11356 2396 -7717
rect 3832 -8034 3892 -8028
rect 3942 -8034 4002 -8028
rect 4596 -8034 4656 -8028
rect 4702 -8034 4762 -8028
rect 4812 -8034 4872 -8028
rect 5464 -8034 5524 -8028
rect 5576 -8034 5636 -8028
rect 6048 -8034 6108 -8028
rect 3892 -8094 3942 -8034
rect 4002 -8094 4596 -8034
rect 4656 -8094 4702 -8034
rect 4762 -8094 4812 -8034
rect 4872 -8094 5464 -8034
rect 5524 -8094 5576 -8034
rect 5636 -8094 6048 -8034
rect 3832 -8100 3892 -8094
rect 3942 -8100 4002 -8094
rect 4596 -8100 4656 -8094
rect 4702 -8100 4762 -8094
rect 4812 -8100 4872 -8094
rect 5464 -8100 5524 -8094
rect 5576 -8100 5636 -8094
rect 6048 -8100 6108 -8094
rect 2110 -11414 2170 -11408
rect 2330 -11416 2336 -11356
rect 2396 -11416 2402 -11356
rect 6914 -11476 6974 -6924
rect 8480 -6930 8540 -6924
rect 10516 -6930 10576 -6924
rect 13570 -6862 13630 -6856
rect 15606 -6862 15666 -6856
rect 13630 -6922 15606 -6862
rect 13570 -6928 13630 -6922
rect 15606 -6928 15666 -6922
rect 18660 -6860 18720 -6854
rect 20696 -6860 20756 -6854
rect 18720 -6920 20696 -6860
rect 18660 -6926 18720 -6920
rect 20696 -6926 20756 -6920
rect 10516 -6972 10576 -6966
rect 22846 -6972 22906 -6966
rect 10576 -7032 22846 -6972
rect 10516 -7038 10576 -7032
rect 22846 -7038 22906 -7032
rect 7312 -7072 7372 -7066
rect 7372 -7132 19896 -7072
rect 7312 -7138 7372 -7132
rect 11732 -7168 11792 -7162
rect 9494 -7174 9554 -7168
rect 11528 -7174 11588 -7168
rect 9554 -7234 11528 -7174
rect 11792 -7228 13566 -7168
rect 13626 -7228 13632 -7168
rect 14586 -7172 14646 -7166
rect 16620 -7172 16680 -7166
rect 11732 -7234 11792 -7228
rect 14646 -7232 16620 -7172
rect 9494 -7240 9554 -7234
rect 11528 -7240 11588 -7234
rect 14586 -7238 14646 -7232
rect 16620 -7238 16680 -7232
rect 16834 -7176 16894 -7170
rect 19682 -7174 19742 -7168
rect 19836 -7174 19896 -7132
rect 21716 -7174 21776 -7168
rect 16894 -7236 19170 -7176
rect 19230 -7236 19236 -7176
rect 19742 -7234 21716 -7174
rect 16834 -7242 16894 -7236
rect 19682 -7240 19742 -7234
rect 21716 -7240 21776 -7234
rect 7044 -8122 7104 -8116
rect 8476 -8122 8536 -8116
rect 10512 -8122 10572 -8116
rect 7104 -8182 8476 -8122
rect 8536 -8182 10512 -8122
rect 7044 -8188 7104 -8182
rect 8476 -8188 8536 -8182
rect 10512 -8188 10572 -8182
rect 18664 -8122 18724 -8116
rect 20700 -8122 20760 -8116
rect 18724 -8182 20700 -8122
rect 18664 -8188 18724 -8182
rect 7180 -8252 7240 -8246
rect 18794 -8252 18854 -8182
rect 20700 -8188 20760 -8182
rect 7240 -8312 18854 -8252
rect 7180 -8318 7240 -8312
rect 11534 -8392 11594 -8386
rect 23138 -8392 23198 -8386
rect 11594 -8452 23138 -8392
rect 11534 -8458 11594 -8452
rect 1720 -11536 6974 -11476
rect 1720 -16460 1780 -11536
rect 1850 -12448 1910 -12442
rect 2568 -12448 2628 -12442
rect 4604 -12448 4664 -12442
rect 6638 -12448 6698 -12442
rect 8678 -12448 8738 -12442
rect 10714 -12448 10774 -12442
rect 12748 -12448 12808 -12442
rect 14784 -12448 14844 -12442
rect 16820 -12448 16880 -12442
rect 18856 -12448 18916 -12442
rect 20894 -12448 20954 -12442
rect 22924 -12448 22984 -12442
rect 1910 -12508 2568 -12448
rect 2628 -12508 4604 -12448
rect 4664 -12508 6638 -12448
rect 6698 -12508 8678 -12448
rect 8738 -12508 10714 -12448
rect 10774 -12508 12748 -12448
rect 12808 -12508 14784 -12448
rect 14844 -12508 16820 -12448
rect 16880 -12508 18856 -12448
rect 18916 -12508 20894 -12448
rect 20954 -12508 22924 -12448
rect 1850 -12514 1910 -12508
rect 2568 -12514 2628 -12508
rect 4604 -12514 4664 -12508
rect 6638 -12514 6698 -12508
rect 8678 -12514 8738 -12508
rect 10714 -12514 10774 -12508
rect 12748 -12514 12808 -12508
rect 14784 -12514 14844 -12508
rect 16820 -12514 16880 -12508
rect 18856 -12514 18916 -12508
rect 20894 -12514 20954 -12508
rect 22924 -12514 22984 -12508
rect 3586 -12546 3646 -12540
rect 5624 -12546 5684 -12540
rect 7658 -12546 7718 -12540
rect 9692 -12546 9752 -12540
rect 11732 -12546 11792 -12540
rect 13766 -12546 13826 -12540
rect 15804 -12546 15864 -12540
rect 17836 -12546 17896 -12540
rect 19874 -12546 19934 -12540
rect 21912 -12546 21972 -12540
rect 23046 -12546 23106 -8452
rect 23138 -8458 23198 -8452
rect 23648 -12546 23708 -12540
rect 3646 -12606 5624 -12546
rect 5684 -12606 7658 -12546
rect 7718 -12606 9692 -12546
rect 9752 -12606 11732 -12546
rect 11792 -12606 13766 -12546
rect 13826 -12606 15804 -12546
rect 15864 -12606 17836 -12546
rect 17896 -12606 19874 -12546
rect 19934 -12606 21912 -12546
rect 21972 -12606 23648 -12546
rect 3586 -12612 3646 -12606
rect 5624 -12612 5684 -12606
rect 7658 -12612 7718 -12606
rect 9692 -12612 9752 -12606
rect 11732 -12612 11792 -12606
rect 13766 -12612 13826 -12606
rect 15804 -12612 15864 -12606
rect 17836 -12612 17896 -12606
rect 19874 -12612 19934 -12606
rect 21912 -12612 21972 -12606
rect 23648 -12612 23708 -12606
rect 11732 -12758 11792 -12752
rect 13764 -12758 13824 -12752
rect 11792 -12818 13764 -12758
rect 11732 -12824 11792 -12818
rect 13764 -12824 13824 -12818
rect 6272 -13678 6332 -13672
rect 6642 -13678 6702 -13672
rect 7144 -13678 7204 -13672
rect 7656 -13678 7716 -13672
rect 8184 -13678 8244 -13672
rect 8676 -13678 8736 -13672
rect 10708 -13678 10768 -13672
rect 12744 -13678 12804 -13672
rect 14780 -13678 14840 -13672
rect 16818 -13678 16878 -13672
rect 18856 -13678 18916 -13672
rect 19364 -13678 19424 -13672
rect 6332 -13738 6642 -13678
rect 6702 -13738 7144 -13678
rect 7204 -13738 7656 -13678
rect 7716 -13738 8184 -13678
rect 8244 -13738 8676 -13678
rect 8736 -13738 10708 -13678
rect 10768 -13738 12744 -13678
rect 12804 -13738 14780 -13678
rect 14840 -13738 16818 -13678
rect 16878 -13738 18342 -13678
rect 18402 -13738 18856 -13678
rect 18916 -13738 19364 -13678
rect 6272 -13744 6332 -13738
rect 6642 -13744 6702 -13738
rect 7144 -13744 7204 -13738
rect 7656 -13744 7716 -13738
rect 8184 -13744 8244 -13738
rect 8676 -13744 8736 -13738
rect 10708 -13744 10768 -13738
rect 12744 -13744 12804 -13738
rect 14780 -13744 14840 -13738
rect 16818 -13744 16878 -13738
rect 18856 -13744 18916 -13738
rect 19364 -13744 19424 -13738
rect 4096 -13788 4156 -13782
rect 5118 -13788 5178 -13782
rect 9190 -13788 9250 -13782
rect 9694 -13788 9754 -13782
rect 10210 -13788 10270 -13782
rect 11230 -13788 11290 -13782
rect 11732 -13788 11792 -13782
rect 12232 -13788 12292 -13782
rect 13258 -13788 13318 -13782
rect 13768 -13788 13828 -13782
rect 14276 -13788 14336 -13782
rect 15284 -13788 15344 -13782
rect 15806 -13788 15866 -13782
rect 16296 -13788 16356 -13782
rect 17328 -13788 17388 -13782
rect 17840 -13788 17900 -13782
rect 20384 -13788 20444 -13782
rect 21404 -13788 21464 -13782
rect 2106 -13848 2112 -13788
rect 2172 -13848 4096 -13788
rect 4156 -13848 5118 -13788
rect 5178 -13848 9190 -13788
rect 9250 -13848 9694 -13788
rect 9754 -13848 10210 -13788
rect 10270 -13848 11230 -13788
rect 11290 -13848 11732 -13788
rect 11792 -13848 12232 -13788
rect 12292 -13848 13258 -13788
rect 13318 -13848 13768 -13788
rect 13828 -13848 14276 -13788
rect 14336 -13848 15284 -13788
rect 15344 -13848 15806 -13788
rect 15866 -13848 16296 -13788
rect 16356 -13848 17328 -13788
rect 17388 -13848 17840 -13788
rect 17900 -13848 20384 -13788
rect 20444 -13848 21404 -13788
rect 4096 -13854 4156 -13848
rect 5118 -13854 5178 -13848
rect 9190 -13854 9250 -13848
rect 9694 -13854 9754 -13848
rect 10210 -13854 10270 -13848
rect 11230 -13854 11290 -13848
rect 11732 -13854 11792 -13848
rect 12232 -13854 12292 -13848
rect 13258 -13854 13318 -13848
rect 13768 -13854 13828 -13848
rect 14276 -13854 14336 -13848
rect 15284 -13854 15344 -13848
rect 15806 -13854 15866 -13848
rect 16296 -13854 16356 -13848
rect 17328 -13854 17388 -13848
rect 17840 -13854 17900 -13848
rect 20384 -13854 20444 -13848
rect 21404 -13854 21464 -13848
rect 7138 -13892 7198 -13886
rect 8158 -13892 8218 -13886
rect 12372 -13892 12432 -13886
rect 13380 -13892 13440 -13886
rect 14422 -13892 14482 -13886
rect 17314 -13892 17374 -13886
rect 18352 -13892 18412 -13886
rect 19352 -13892 19412 -13886
rect 6132 -13952 6138 -13892
rect 6198 -13952 7138 -13892
rect 7198 -13952 8158 -13892
rect 8218 -13952 12372 -13892
rect 12432 -13952 13380 -13892
rect 13440 -13952 14422 -13892
rect 14482 -13952 17314 -13892
rect 17374 -13952 18352 -13892
rect 18412 -13952 19352 -13892
rect 7138 -13958 7198 -13952
rect 8158 -13958 8218 -13952
rect 12372 -13958 12432 -13952
rect 13380 -13958 13440 -13952
rect 14422 -13958 14482 -13952
rect 17314 -13958 17374 -13952
rect 18352 -13958 18412 -13952
rect 19352 -13958 19412 -13952
rect 1976 -14000 2036 -13994
rect 2572 -14000 2632 -13994
rect 3070 -14000 3130 -13994
rect 3582 -14000 3642 -13994
rect 5624 -14000 5684 -13994
rect 7658 -14000 7718 -13994
rect 9692 -14000 9752 -13994
rect 15806 -14000 15866 -13994
rect 17838 -14000 17898 -13994
rect 19870 -14000 19930 -13994
rect 21912 -14000 21972 -13994
rect 22416 -14000 22476 -13994
rect 22926 -14000 22986 -13994
rect 2036 -14060 2572 -14000
rect 2632 -14060 3070 -14000
rect 3130 -14060 3582 -14000
rect 3642 -14060 5624 -14000
rect 5684 -14060 7658 -14000
rect 7718 -14060 9692 -14000
rect 9752 -14060 11848 -14000
rect 11908 -14002 15806 -14000
rect 11908 -14060 13572 -14002
rect 1976 -14066 2036 -14060
rect 2572 -14066 2632 -14060
rect 3070 -14066 3130 -14060
rect 3582 -14066 3642 -14060
rect 5624 -14066 5684 -14060
rect 7658 -14066 7718 -14060
rect 9692 -14066 9752 -14060
rect 13566 -14062 13572 -14060
rect 13632 -14060 15806 -14002
rect 15866 -14060 17838 -14000
rect 17898 -14060 19870 -14000
rect 19930 -14060 21912 -14000
rect 21972 -14060 22416 -14000
rect 22476 -14060 22926 -14000
rect 13632 -14062 13638 -14060
rect 15806 -14066 15866 -14060
rect 17838 -14066 17898 -14060
rect 19870 -14066 19930 -14060
rect 21912 -14066 21972 -14060
rect 22416 -14066 22476 -14060
rect 22926 -14066 22986 -14060
rect 5102 -14890 5162 -14884
rect 6122 -14890 6182 -14884
rect 7134 -14890 7194 -14884
rect 8160 -14890 8220 -14884
rect 17316 -14890 17376 -14884
rect 18352 -14890 18412 -14884
rect 19368 -14890 19428 -14884
rect 1850 -14902 1910 -14896
rect 4086 -14902 4146 -14896
rect 1910 -14962 4086 -14902
rect 5162 -14950 6122 -14890
rect 6182 -14950 7134 -14890
rect 7194 -14950 8160 -14890
rect 8220 -14950 17316 -14890
rect 17376 -14950 18352 -14890
rect 18412 -14950 19368 -14890
rect 5102 -14956 5162 -14950
rect 6122 -14956 6182 -14950
rect 7134 -14956 7194 -14950
rect 8160 -14956 8220 -14950
rect 17316 -14956 17376 -14950
rect 18352 -14956 18412 -14950
rect 19368 -14956 19428 -14950
rect 1850 -14968 1910 -14962
rect 4086 -14968 4146 -14962
rect 4598 -14994 4658 -14988
rect 5622 -14994 5682 -14988
rect 6634 -14994 6694 -14988
rect 7654 -14994 7714 -14988
rect 8676 -14994 8736 -14988
rect 10712 -14994 10772 -14988
rect 12750 -14994 12810 -14988
rect 14780 -14994 14840 -14988
rect 15800 -14994 15860 -14988
rect 16818 -14994 16878 -14988
rect 17838 -14994 17898 -14988
rect 18854 -14994 18914 -14988
rect 20890 -14994 20950 -14988
rect 4658 -15054 5622 -14994
rect 5682 -15054 6634 -14994
rect 6694 -15054 7654 -14994
rect 7714 -15054 8676 -14994
rect 8736 -15054 10712 -14994
rect 10772 -15054 12750 -14994
rect 12810 -15054 14780 -14994
rect 14840 -15054 15800 -14994
rect 15860 -15054 16818 -14994
rect 16878 -15054 17838 -14994
rect 17898 -15054 18854 -14994
rect 18914 -15054 20890 -14994
rect 4598 -15060 4658 -15054
rect 5622 -15060 5682 -15054
rect 6634 -15060 6694 -15054
rect 7654 -15060 7714 -15054
rect 8676 -15060 8736 -15054
rect 10712 -15060 10772 -15054
rect 12750 -15060 12810 -15054
rect 14780 -15060 14840 -15054
rect 15800 -15060 15860 -15054
rect 16818 -15060 16878 -15054
rect 17838 -15060 17898 -15054
rect 18854 -15060 18914 -15054
rect 20890 -15060 20950 -15054
rect 2336 -15116 2396 -15110
rect 9696 -15116 9756 -15110
rect 11730 -15116 11790 -15110
rect 13760 -15116 13820 -15110
rect 23760 -15116 23820 -5972
rect 2396 -15176 9696 -15116
rect 9756 -15176 11730 -15116
rect 11790 -15176 13760 -15116
rect 13820 -15176 23820 -15116
rect 2336 -15182 2396 -15176
rect 9696 -15182 9756 -15176
rect 11730 -15182 11790 -15176
rect 13760 -15182 13820 -15176
rect 4604 -15228 4664 -15222
rect 6640 -15228 6700 -15222
rect 23034 -15228 23094 -15222
rect 4664 -15288 6640 -15228
rect 6700 -15288 23034 -15228
rect 4604 -15294 4664 -15288
rect 6640 -15294 6700 -15288
rect 23034 -15294 23094 -15288
rect 22928 -16116 22988 -16110
rect 23888 -16116 23948 -5654
rect 5620 -16134 5680 -16128
rect 7656 -16134 7716 -16128
rect 15800 -16134 15860 -16128
rect 17836 -16134 17896 -16128
rect 21910 -16134 21970 -16128
rect 2448 -16158 2508 -16152
rect 3586 -16158 3646 -16152
rect 2508 -16218 3586 -16158
rect 3646 -16218 4468 -16158
rect 5680 -16194 7656 -16134
rect 7716 -16194 15800 -16134
rect 15860 -16194 17836 -16134
rect 17896 -16194 21910 -16134
rect 22988 -16176 23948 -16116
rect 22928 -16182 22988 -16176
rect 5620 -16200 5680 -16194
rect 7656 -16200 7716 -16194
rect 15800 -16200 15860 -16194
rect 17836 -16200 17896 -16194
rect 21910 -16200 21970 -16194
rect 2448 -16224 2508 -16218
rect 3586 -16224 3646 -16218
rect 2336 -16358 2396 -16352
rect 3584 -16358 3644 -16352
rect 2396 -16418 3584 -16358
rect 4408 -16354 4468 -16218
rect 4602 -16238 4662 -16232
rect 6642 -16238 6702 -16232
rect 8674 -16238 8734 -16232
rect 10708 -16238 10768 -16232
rect 12748 -16238 12808 -16232
rect 14782 -16238 14842 -16232
rect 4662 -16298 6642 -16238
rect 6702 -16298 8674 -16238
rect 8734 -16298 10708 -16238
rect 10768 -16298 12748 -16238
rect 12808 -16298 14782 -16238
rect 4602 -16304 4662 -16298
rect 6642 -16304 6702 -16298
rect 8674 -16304 8734 -16298
rect 10708 -16304 10768 -16298
rect 12748 -16304 12808 -16298
rect 14782 -16304 14842 -16298
rect 14978 -16242 15038 -16236
rect 19870 -16242 19930 -16236
rect 15038 -16302 19870 -16242
rect 23528 -16246 23588 -16240
rect 14978 -16308 15038 -16302
rect 19870 -16308 19930 -16302
rect 20368 -16306 20374 -16246
rect 20434 -16306 23528 -16246
rect 23528 -16312 23588 -16306
rect 5116 -16352 5176 -16346
rect 8674 -16350 8734 -16344
rect 10710 -16350 10770 -16344
rect 12746 -16350 12806 -16344
rect 14782 -16350 14842 -16344
rect 16816 -16350 16876 -16344
rect 18854 -16350 18914 -16344
rect 20894 -16350 20954 -16344
rect 23278 -16350 23338 -16344
rect 4408 -16412 5116 -16354
rect 5176 -16412 6120 -16352
rect 6180 -16412 7132 -16352
rect 7192 -16412 8152 -16352
rect 8212 -16412 8218 -16352
rect 8734 -16410 10710 -16350
rect 10770 -16410 12746 -16350
rect 12806 -16410 14782 -16350
rect 14842 -16410 16816 -16350
rect 16876 -16410 18854 -16350
rect 18914 -16410 20894 -16350
rect 20954 -16410 23278 -16350
rect 4408 -16414 5458 -16412
rect 5116 -16418 5176 -16414
rect 8674 -16416 8734 -16410
rect 10710 -16416 10770 -16410
rect 12746 -16416 12806 -16410
rect 14782 -16416 14842 -16410
rect 16816 -16416 16876 -16410
rect 18854 -16416 18914 -16410
rect 20894 -16416 20954 -16410
rect 23278 -16416 23338 -16410
rect 2336 -16424 2396 -16418
rect 3584 -16424 3644 -16418
rect 2230 -16460 2290 -16454
rect 9692 -16460 9752 -16454
rect 11726 -16460 11786 -16454
rect 13766 -16460 13826 -16454
rect 14978 -16460 15038 -16454
rect 1720 -16520 2230 -16460
rect 2290 -16520 9692 -16460
rect 9752 -16520 11726 -16460
rect 11786 -16520 13766 -16460
rect 13826 -16520 14978 -16460
rect 2230 -16526 2290 -16520
rect 9692 -16526 9752 -16520
rect 11726 -16526 11786 -16520
rect 13766 -16526 13826 -16520
rect 14978 -16526 15038 -16520
rect 15272 -16458 15332 -16452
rect 15332 -16518 16300 -16458
rect 16360 -16518 16366 -16458
rect 16818 -16464 16878 -16458
rect 18854 -16464 18914 -16458
rect 20892 -16464 20952 -16458
rect 23034 -16464 23094 -16458
rect 15272 -16524 15332 -16518
rect 16878 -16524 18854 -16464
rect 18914 -16524 20892 -16464
rect 20952 -16524 23034 -16464
rect 16818 -16530 16878 -16524
rect 18854 -16530 18914 -16524
rect 20892 -16530 20952 -16524
rect 23034 -16530 23094 -16524
rect 19366 -17378 19426 -17372
rect 3584 -17390 3644 -17384
rect 5622 -17390 5682 -17384
rect 7658 -17390 7718 -17384
rect 9690 -17390 9750 -17384
rect 3644 -17450 5622 -17390
rect 5682 -17450 7658 -17390
rect 7718 -17450 9690 -17390
rect 14266 -17438 14272 -17378
rect 14332 -17438 19366 -17378
rect 19366 -17444 19426 -17438
rect 19504 -17374 19564 -17368
rect 20386 -17374 20446 -17368
rect 21392 -17374 21452 -17368
rect 19564 -17434 20386 -17374
rect 20446 -17434 21392 -17374
rect 19504 -17440 19564 -17434
rect 20386 -17440 20446 -17434
rect 21392 -17440 21452 -17434
rect 21910 -17378 21970 -17372
rect 23162 -17378 23222 -17372
rect 21970 -17438 23162 -17378
rect 21910 -17444 21970 -17438
rect 23162 -17444 23222 -17438
rect 3584 -17456 3644 -17450
rect 5622 -17456 5682 -17450
rect 7658 -17456 7718 -17450
rect 9690 -17456 9750 -17450
rect 4090 -17492 4150 -17486
rect 9182 -17492 9242 -17486
rect 4150 -17552 9182 -17492
rect 4090 -17558 4150 -17552
rect 9182 -17558 9242 -17552
rect 13766 -17506 13826 -17500
rect 21910 -17506 21970 -17500
rect 13826 -17566 21910 -17506
rect 13766 -17572 13826 -17566
rect 21910 -17572 21970 -17566
rect 2336 -17594 2396 -17588
rect 5620 -17594 5680 -17588
rect 2396 -17654 5620 -17594
rect 2336 -17660 2396 -17654
rect 5620 -17660 5680 -17654
rect 6128 -17600 6188 -17594
rect 7150 -17600 7210 -17594
rect 8164 -17600 8224 -17594
rect 9182 -17600 9242 -17594
rect 10202 -17600 10262 -17594
rect 17314 -17600 17374 -17594
rect 18344 -17600 18404 -17594
rect 19504 -17600 19564 -17594
rect 6188 -17660 7150 -17600
rect 7210 -17660 8164 -17600
rect 8224 -17660 9182 -17600
rect 9242 -17660 10202 -17600
rect 10262 -17660 17314 -17600
rect 17374 -17660 18344 -17600
rect 18404 -17660 19504 -17600
rect 6128 -17666 6188 -17660
rect 7150 -17666 7210 -17660
rect 8164 -17666 8224 -17660
rect 9182 -17666 9242 -17660
rect 10202 -17666 10262 -17660
rect 17314 -17666 17374 -17660
rect 18344 -17666 18404 -17660
rect 19504 -17666 19564 -17660
rect 19872 -17600 19932 -17594
rect 23400 -17600 23460 -17594
rect 19932 -17660 23400 -17600
rect 19872 -17666 19932 -17660
rect 23400 -17666 23460 -17660
rect 4604 -17694 4664 -17688
rect 6638 -17694 6698 -17688
rect 8674 -17694 8734 -17688
rect 4664 -17754 6638 -17694
rect 6698 -17754 8674 -17694
rect 4604 -17760 4664 -17754
rect 6638 -17760 6698 -17754
rect 8674 -17760 8734 -17754
rect 15802 -17704 15862 -17698
rect 19872 -17704 19932 -17698
rect 15862 -17764 19872 -17704
rect 15802 -17770 15862 -17764
rect 19872 -17770 19932 -17764
rect 20888 -17702 20948 -17696
rect 23278 -17702 23338 -17696
rect 20948 -17762 23278 -17702
rect 20888 -17768 20948 -17762
rect 23278 -17768 23338 -17762
rect 10710 -18612 10770 -18606
rect 12746 -18612 12806 -18606
rect 14782 -18612 14842 -18606
rect 16820 -18612 16880 -18606
rect 4086 -18618 4146 -18612
rect 4996 -18618 5056 -18612
rect 5998 -18618 6058 -18612
rect 7150 -18618 7210 -18612
rect 8160 -18618 8220 -18612
rect 9166 -18618 9226 -18612
rect 10210 -18618 10270 -18612
rect 4146 -18678 4996 -18618
rect 5056 -18678 5998 -18618
rect 6058 -18678 7150 -18618
rect 7210 -18678 8160 -18618
rect 8220 -18678 9166 -18618
rect 9226 -18678 10210 -18618
rect 10770 -18672 12746 -18612
rect 12806 -18672 14782 -18612
rect 14842 -18672 16820 -18612
rect 10710 -18678 10770 -18672
rect 12746 -18678 12806 -18672
rect 14782 -18678 14842 -18672
rect 16820 -18678 16880 -18672
rect 18856 -18612 18916 -18606
rect 20894 -18612 20954 -18606
rect 18916 -18672 20894 -18612
rect 18856 -18678 18916 -18672
rect 20894 -18678 20954 -18672
rect 4086 -18684 4146 -18678
rect 4996 -18684 5056 -18678
rect 5998 -18684 6058 -18678
rect 7150 -18684 7210 -18678
rect 8160 -18684 8220 -18678
rect 9166 -18684 9226 -18678
rect 10210 -18684 10270 -18678
rect 6638 -18720 6698 -18714
rect 16812 -18720 16872 -18714
rect 18852 -18720 18912 -18714
rect 20890 -18720 20950 -18714
rect 6698 -18780 16812 -18720
rect 16872 -18780 18852 -18720
rect 18912 -18780 20890 -18720
rect 6638 -18786 6698 -18780
rect 16812 -18786 16872 -18780
rect 18852 -18786 18912 -18780
rect 20890 -18786 20950 -18780
rect 4086 -18834 4146 -18828
rect 6138 -18834 6198 -18828
rect 9164 -18834 9224 -18828
rect 10204 -18834 10264 -18828
rect 11218 -18834 11278 -18828
rect 12226 -18834 12286 -18828
rect 13270 -18834 13330 -18828
rect 14260 -18834 14320 -18828
rect 15278 -18834 15338 -18828
rect 16312 -18834 16372 -18828
rect 19344 -18834 19404 -18828
rect 20382 -18834 20442 -18828
rect 21408 -18834 21468 -18828
rect 4146 -18894 5124 -18834
rect 5184 -18894 6138 -18834
rect 6198 -18894 9164 -18834
rect 9224 -18894 10204 -18834
rect 10264 -18894 11218 -18834
rect 11278 -18894 12226 -18834
rect 12286 -18894 13270 -18834
rect 13330 -18894 14260 -18834
rect 14320 -18894 15278 -18834
rect 15338 -18894 16312 -18834
rect 16372 -18894 19344 -18834
rect 19404 -18894 20382 -18834
rect 20442 -18894 21408 -18834
rect 21468 -18894 23526 -18834
rect 23586 -18894 23592 -18834
rect 4086 -18900 4146 -18894
rect 6138 -18900 6198 -18894
rect 9164 -18900 9224 -18894
rect 10204 -18900 10264 -18894
rect 11218 -18900 11278 -18894
rect 12226 -18900 12286 -18894
rect 13270 -18900 13330 -18894
rect 14260 -18900 14320 -18894
rect 15278 -18900 15338 -18894
rect 16312 -18900 16372 -18894
rect 19344 -18900 19404 -18894
rect 20382 -18900 20442 -18894
rect 21408 -18900 21468 -18894
rect 9688 -18938 9748 -18932
rect 11730 -18938 11790 -18932
rect 13768 -18938 13828 -18932
rect 15802 -18938 15862 -18932
rect 17836 -18936 17896 -18930
rect 19870 -18936 19930 -18930
rect 21912 -18936 21972 -18930
rect 23162 -18936 23222 -18930
rect 2444 -18998 2450 -18938
rect 2510 -18998 9688 -18938
rect 9748 -18998 11730 -18938
rect 11790 -18998 13768 -18938
rect 13828 -18998 15802 -18938
rect 9688 -19004 9748 -18998
rect 11730 -19004 11790 -18998
rect 13768 -19004 13828 -18998
rect 15802 -19004 15862 -18998
rect 16314 -18942 16374 -18936
rect 17336 -18942 17396 -18936
rect 16374 -19002 17336 -18942
rect 17896 -18996 19870 -18936
rect 19930 -18996 21912 -18936
rect 21972 -18996 23162 -18936
rect 17836 -19002 17896 -18996
rect 19870 -19002 19930 -18996
rect 21912 -19002 21972 -18996
rect 23162 -19002 23222 -18996
rect 16314 -19008 16374 -19002
rect 17336 -19008 17396 -19002
rect 8678 -19840 8738 -19834
rect 12746 -19840 12806 -19834
rect 14780 -19840 14840 -19834
rect 4084 -19846 4144 -19840
rect 5092 -19846 5152 -19840
rect 6106 -19846 6166 -19840
rect 7144 -19846 7204 -19840
rect 8162 -19846 8222 -19840
rect 4144 -19906 5092 -19846
rect 5152 -19906 6106 -19846
rect 6166 -19906 7144 -19846
rect 7204 -19906 8162 -19846
rect 8738 -19900 10714 -19840
rect 10774 -19900 12746 -19840
rect 12806 -19900 14780 -19840
rect 8678 -19906 8738 -19900
rect 12746 -19906 12806 -19900
rect 14780 -19906 14840 -19900
rect 15802 -19838 15862 -19832
rect 16156 -19838 16216 -19832
rect 15862 -19898 16156 -19838
rect 15802 -19904 15862 -19898
rect 16156 -19904 16216 -19898
rect 19874 -19838 19934 -19832
rect 23158 -19838 23218 -19832
rect 19934 -19898 23158 -19838
rect 19874 -19904 19934 -19898
rect 23158 -19904 23218 -19898
rect 4084 -19912 4144 -19906
rect 5092 -19912 5152 -19906
rect 6106 -19912 6166 -19906
rect 7144 -19912 7204 -19906
rect 8162 -19912 8222 -19906
rect 2230 -19950 2290 -19944
rect 3586 -19950 3646 -19944
rect 11730 -19950 11790 -19944
rect 13766 -19950 13826 -19944
rect 15798 -19950 15858 -19944
rect 2290 -20010 3586 -19950
rect 3646 -20010 11730 -19950
rect 11790 -20010 13766 -19950
rect 13826 -20010 15798 -19950
rect 2230 -20016 2290 -20010
rect 3586 -20016 3646 -20010
rect 11730 -20016 11790 -20010
rect 13766 -20016 13826 -20010
rect 15798 -20016 15858 -20010
rect 15308 -20048 15368 -20042
rect 16346 -20048 16406 -20042
rect 17322 -20048 17382 -20042
rect 18338 -20048 18398 -20042
rect 20364 -20048 20424 -20042
rect 21394 -20048 21454 -20042
rect -314 -20130 1646 -20070
rect 4602 -20062 4662 -20056
rect 6640 -20062 6700 -20056
rect 10712 -20062 10772 -20056
rect 4662 -20122 6640 -20062
rect 6700 -20122 10712 -20062
rect 15368 -20108 16346 -20048
rect 16406 -20108 17322 -20048
rect 17382 -20108 18338 -20048
rect 18398 -20108 20364 -20048
rect 20424 -20108 21394 -20048
rect 15308 -20114 15368 -20108
rect 16346 -20114 16406 -20108
rect 17322 -20114 17382 -20108
rect 18338 -20114 18398 -20108
rect 20364 -20114 20424 -20108
rect 21394 -20114 21454 -20108
rect 4602 -20128 4662 -20122
rect 6640 -20128 6700 -20122
rect 10712 -20128 10772 -20122
rect -374 -20136 -314 -20130
rect -592 -20160 -532 -20154
rect -968 -20220 -592 -20160
rect 3582 -20160 3642 -20154
rect 5620 -20160 5680 -20154
rect 7660 -20160 7720 -20154
rect 9696 -20160 9756 -20154
rect 15800 -20160 15860 -20154
rect 16150 -20160 16156 -20156
rect 2336 -20196 2396 -20190
rect -1028 -20226 -968 -20220
rect -592 -20226 -532 -20220
rect 214 -20256 220 -20196
rect 280 -20256 2336 -20196
rect 3642 -20220 5620 -20160
rect 5680 -20220 7660 -20160
rect 7720 -20220 9696 -20160
rect 9756 -20216 16156 -20160
rect 16216 -20160 16222 -20156
rect 17836 -20160 17896 -20154
rect 19872 -20160 19932 -20154
rect 21908 -20160 21968 -20154
rect 16216 -20216 17836 -20160
rect 9756 -20220 17836 -20216
rect 17896 -20220 19872 -20160
rect 19932 -20220 21908 -20160
rect 3582 -20226 3642 -20220
rect 5620 -20226 5680 -20220
rect 7660 -20226 7720 -20220
rect 9696 -20226 9756 -20220
rect 15800 -20226 15860 -20220
rect 17836 -20226 17896 -20220
rect 19872 -20226 19932 -20220
rect 21908 -20226 21968 -20220
rect 2336 -20262 2396 -20256
rect -1792 -20270 -1732 -20264
rect -1572 -20270 -1512 -20264
rect -918 -20270 -858 -20264
rect -702 -20270 -642 -20264
rect -1732 -20330 -1572 -20270
rect -1512 -20330 -918 -20270
rect -858 -20330 -702 -20270
rect -1792 -20336 -1732 -20330
rect -1572 -20336 -1512 -20330
rect -918 -20336 -858 -20330
rect -702 -20336 -642 -20330
rect -2468 -20774 -2408 -20768
rect -2010 -20774 -1950 -20768
rect -1354 -20774 -1294 -20768
rect -2408 -20834 -2010 -20774
rect -1950 -20834 -1354 -20774
rect -2468 -20840 -2408 -20834
rect -2010 -20840 -1950 -20834
rect -1354 -20840 -1294 -20834
rect -810 -20774 -750 -20768
rect -22 -20774 38 -20768
rect -750 -20834 -22 -20774
rect -810 -20840 -750 -20834
rect -22 -20840 38 -20834
rect -2598 -20896 -2538 -20890
rect -1792 -20896 -1732 -20890
rect -1574 -20896 -1514 -20890
rect -2538 -20956 -1792 -20896
rect -1732 -20956 -1574 -20896
rect -2598 -20962 -2538 -20956
rect -1792 -20962 -1732 -20956
rect -1574 -20962 -1514 -20956
rect -1138 -20894 -1078 -20888
rect -482 -20894 -422 -20888
rect -1078 -20954 -482 -20894
rect -1138 -20960 -1078 -20954
rect -482 -20960 -422 -20954
rect -2118 -21020 -2058 -21014
rect -1248 -21020 -1188 -21014
rect -376 -21020 -316 -21014
rect -2058 -21080 -1248 -21020
rect -1188 -21080 -376 -21020
rect 10708 -21064 10768 -21058
rect 12750 -21064 12810 -21058
rect 14782 -21064 14842 -21058
rect 16822 -21064 16882 -21058
rect 23278 -21064 23338 -21058
rect -2118 -21086 -2058 -21080
rect -1248 -21086 -1188 -21080
rect -376 -21086 -316 -21080
rect 4602 -21084 4662 -21078
rect 6638 -21084 6698 -21078
rect 8676 -21084 8736 -21078
rect -1680 -21146 -1620 -21140
rect 98 -21146 158 -21140
rect -1620 -21206 98 -21146
rect 4662 -21144 6638 -21084
rect 6698 -21144 8676 -21084
rect 10532 -21124 10538 -21064
rect 10598 -21124 10708 -21064
rect 10768 -21124 12750 -21064
rect 12810 -21124 14782 -21064
rect 14842 -21124 16822 -21064
rect 16882 -21124 23278 -21064
rect 10708 -21130 10768 -21124
rect 12750 -21130 12810 -21124
rect 14782 -21130 14842 -21124
rect 16822 -21130 16882 -21124
rect 23278 -21130 23338 -21124
rect 4602 -21150 4662 -21144
rect 6638 -21150 6698 -21144
rect 8676 -21150 8736 -21144
rect 15800 -21162 15860 -21156
rect 21906 -21162 21966 -21156
rect 23158 -21162 23218 -21156
rect -1680 -21212 -1620 -21206
rect 98 -21212 158 -21206
rect 2448 -21182 2508 -21176
rect 5620 -21182 5680 -21176
rect 2508 -21242 5620 -21182
rect 2448 -21248 2508 -21242
rect 5620 -21248 5680 -21242
rect 7144 -21182 7204 -21176
rect 10192 -21182 10252 -21176
rect 7204 -21242 8166 -21182
rect 8226 -21242 9188 -21182
rect 9248 -21242 10192 -21182
rect 15860 -21222 21906 -21162
rect 21966 -21222 23158 -21162
rect 15800 -21228 15860 -21222
rect 21906 -21228 21966 -21222
rect 23158 -21228 23218 -21222
rect 7144 -21248 7204 -21242
rect 10192 -21248 10252 -21242
rect -1346 -21260 -1294 -21254
rect 2236 -21262 2242 -21260
rect -1294 -21310 2242 -21262
rect 2236 -21312 2242 -21310
rect 2294 -21312 2300 -21260
rect 10714 -21272 10774 -21266
rect 12742 -21272 12802 -21266
rect 14786 -21272 14846 -21266
rect 16814 -21272 16874 -21266
rect 18852 -21272 18912 -21266
rect 20892 -21272 20952 -21266
rect 4606 -21278 4666 -21272
rect 6642 -21278 6702 -21272
rect 8670 -21278 8730 -21272
rect 10538 -21278 10598 -21272
rect -1346 -21318 -1294 -21312
rect 4666 -21338 6642 -21278
rect 6702 -21338 8670 -21278
rect 8730 -21338 10538 -21278
rect 10774 -21332 12742 -21272
rect 12802 -21332 14786 -21272
rect 14846 -21332 16814 -21272
rect 16874 -21332 18852 -21272
rect 18912 -21332 20892 -21272
rect 10714 -21338 10774 -21332
rect 12742 -21338 12802 -21332
rect 14786 -21338 14846 -21332
rect 16814 -21338 16874 -21332
rect 18852 -21338 18912 -21332
rect 20892 -21338 20952 -21332
rect 21410 -21268 21470 -21262
rect 23528 -21268 23588 -21262
rect 21470 -21328 23528 -21268
rect 21410 -21334 21470 -21328
rect 23528 -21334 23588 -21328
rect 4606 -21344 4666 -21338
rect 6642 -21344 6702 -21338
rect 8670 -21344 8730 -21338
rect 10538 -21344 10598 -21338
rect 3588 -21398 3648 -21392
rect 7656 -21398 7716 -21392
rect 9690 -21398 9750 -21392
rect 17840 -21398 17900 -21392
rect 19870 -21398 19930 -21392
rect 21908 -21396 21968 -21390
rect 23400 -21396 23460 -21390
rect 3648 -21458 7656 -21398
rect 7716 -21458 9690 -21398
rect 9750 -21458 17840 -21398
rect 17900 -21458 19870 -21398
rect 20390 -21456 20396 -21396
rect 20456 -21456 21908 -21396
rect 21968 -21456 23400 -21396
rect 3588 -21464 3648 -21458
rect 7656 -21464 7716 -21458
rect 9690 -21464 9750 -21458
rect 17840 -21464 17900 -21458
rect 19870 -21464 19930 -21458
rect 21908 -21462 21968 -21456
rect 23400 -21462 23460 -21456
rect -932 -21480 -872 -21474
rect 262 -21480 322 -21474
rect 952 -21480 1012 -21474
rect -2128 -21540 -2122 -21480
rect -2062 -21540 -932 -21480
rect -872 -21540 262 -21480
rect 322 -21540 952 -21480
rect -932 -21546 -872 -21540
rect 262 -21546 322 -21540
rect 952 -21546 1012 -21540
rect -2670 -21580 -2610 -21574
rect -1678 -21580 -1618 -21574
rect -1380 -21580 -1320 -21574
rect -484 -21580 -424 -21574
rect -188 -21580 -128 -21574
rect -2610 -21640 -1678 -21580
rect -1618 -21640 -1380 -21580
rect -1320 -21640 -484 -21580
rect -424 -21640 -188 -21580
rect -2670 -21646 -2610 -21640
rect -1678 -21646 -1618 -21640
rect -1380 -21646 -1320 -21640
rect -484 -21646 -424 -21640
rect -188 -21646 -128 -21640
rect 2336 -22314 2396 -22308
rect 11724 -22314 11784 -22308
rect 13766 -22314 13826 -22308
rect 15802 -22314 15862 -22308
rect 2396 -22374 11724 -22314
rect 11784 -22374 13766 -22314
rect 13826 -22374 15802 -22314
rect 2336 -22380 2396 -22374
rect 11724 -22380 11784 -22374
rect 13766 -22380 13826 -22374
rect 15802 -22380 15862 -22374
rect 18856 -22314 18916 -22308
rect 20888 -22314 20948 -22308
rect 23034 -22314 23094 -22308
rect 18916 -22374 20888 -22314
rect 20948 -22374 23034 -22314
rect 18856 -22380 18916 -22374
rect 20888 -22380 20948 -22374
rect 23034 -22380 23094 -22374
rect 6140 -22428 6200 -22422
rect 11220 -22428 11280 -22422
rect 2230 -22440 2290 -22434
rect 5620 -22440 5680 -22434
rect -1829 -22483 -1771 -22477
rect -1225 -22483 -1167 -22477
rect -634 -22483 -576 -22477
rect -1771 -22541 -1225 -22483
rect -1167 -22541 -634 -22483
rect -576 -22541 -37 -22483
rect 21 -22541 559 -22483
rect 617 -22541 623 -22483
rect 2290 -22500 5620 -22440
rect 6200 -22488 11220 -22428
rect 6140 -22494 6200 -22488
rect 11220 -22494 11280 -22488
rect 16308 -22424 16368 -22418
rect 21408 -22424 21468 -22418
rect 16368 -22484 21408 -22424
rect 16308 -22490 16368 -22484
rect 21408 -22490 21468 -22484
rect 2230 -22506 2290 -22500
rect 5620 -22506 5680 -22500
rect -1829 -22547 -1771 -22541
rect -1225 -22547 -1167 -22541
rect -634 -22547 -576 -22541
rect 4602 -22550 4662 -22544
rect 6638 -22550 6698 -22544
rect 7658 -22550 7718 -22544
rect 8674 -22550 8734 -22544
rect 9694 -22550 9754 -22544
rect 10712 -22550 10772 -22544
rect 12742 -22550 12802 -22544
rect 14780 -22550 14840 -22544
rect 16816 -22550 16876 -22544
rect 17838 -22550 17898 -22544
rect 18858 -22550 18918 -22544
rect 19872 -22550 19932 -22544
rect 20894 -22550 20954 -22544
rect -2542 -22614 -2482 -22608
rect -1532 -22614 -1472 -22608
rect -934 -22614 -874 -22608
rect -340 -22614 -280 -22608
rect 258 -22614 318 -22608
rect -2482 -22674 -2126 -22614
rect -2066 -22674 -1532 -22614
rect -1472 -22674 -934 -22614
rect -874 -22674 -340 -22614
rect -280 -22674 258 -22614
rect 4662 -22610 6638 -22550
rect 6698 -22610 7658 -22550
rect 7718 -22610 8674 -22550
rect 8734 -22610 9694 -22550
rect 9754 -22610 10712 -22550
rect 10772 -22610 12742 -22550
rect 12802 -22610 14780 -22550
rect 14840 -22610 16816 -22550
rect 16876 -22610 17838 -22550
rect 17898 -22610 18858 -22550
rect 18918 -22610 19872 -22550
rect 19932 -22610 20894 -22550
rect 4602 -22616 4662 -22610
rect 6638 -22616 6698 -22610
rect 7658 -22616 7718 -22610
rect 8674 -22616 8734 -22610
rect 9694 -22616 9754 -22610
rect 10712 -22616 10772 -22610
rect 12742 -22616 12802 -22610
rect 14780 -22616 14840 -22610
rect 16816 -22616 16876 -22610
rect 17838 -22616 17898 -22610
rect 18858 -22616 18918 -22610
rect 19872 -22616 19932 -22610
rect 20894 -22616 20954 -22610
rect -2542 -22680 -2482 -22674
rect -1532 -22680 -1472 -22674
rect -934 -22680 -874 -22674
rect -340 -22680 -280 -22674
rect 258 -22680 318 -22674
rect 6256 -22644 6316 -22638
rect 7140 -22644 7200 -22638
rect 8162 -22644 8222 -22638
rect 10204 -22644 10264 -22638
rect 6316 -22704 7140 -22644
rect 7200 -22704 8162 -22644
rect 8222 -22704 10204 -22644
rect 6256 -22710 6316 -22704
rect 7140 -22710 7200 -22704
rect 8162 -22710 8222 -22704
rect 10204 -22710 10264 -22704
rect 17326 -22644 17386 -22638
rect 18346 -22644 18406 -22638
rect 19360 -22644 19420 -22638
rect 20396 -22644 20456 -22638
rect 17386 -22704 18346 -22644
rect 18406 -22704 19360 -22644
rect 19420 -22704 20396 -22644
rect 17326 -22710 17386 -22704
rect 18346 -22710 18406 -22704
rect 19360 -22710 19420 -22704
rect 20396 -22710 20456 -22704
rect -1974 -22722 -1914 -22716
rect -1676 -22722 -1616 -22716
rect -1376 -22722 -1316 -22716
rect -1082 -22722 -1022 -22716
rect -786 -22722 -726 -22716
rect -486 -22722 -426 -22716
rect -184 -22722 -124 -22716
rect 106 -22722 166 -22716
rect 410 -22722 470 -22716
rect -1914 -22782 -1676 -22722
rect -1616 -22782 -1376 -22722
rect -1316 -22782 -1082 -22722
rect -1022 -22782 -786 -22722
rect -726 -22782 -486 -22722
rect -426 -22782 -184 -22722
rect -124 -22782 106 -22722
rect 166 -22782 410 -22722
rect 470 -22782 1076 -22722
rect 1136 -22782 1142 -22722
rect -1974 -22788 -1914 -22782
rect -1676 -22788 -1616 -22782
rect -1376 -22788 -1316 -22782
rect -1082 -22788 -1022 -22782
rect -786 -22788 -726 -22782
rect -486 -22788 -426 -22782
rect -184 -22788 -124 -22782
rect 106 -22788 166 -22782
rect 410 -22788 470 -22782
rect 1976 -23544 2036 -23538
rect 2568 -23544 2628 -23538
rect 3082 -23544 3142 -23538
rect 3580 -23544 3640 -23538
rect 5622 -23544 5682 -23538
rect 7654 -23544 7714 -23538
rect 9686 -23544 9746 -23538
rect 13944 -23544 13950 -23542
rect 1544 -23546 1976 -23544
rect 1400 -23604 1976 -23546
rect 2036 -23604 2568 -23544
rect 2628 -23604 3082 -23544
rect 3142 -23604 3580 -23544
rect 3640 -23604 5622 -23544
rect 5682 -23604 7654 -23544
rect 7714 -23604 9686 -23544
rect 9746 -23604 11590 -23544
rect 11650 -23602 13950 -23544
rect 14010 -23544 14016 -23542
rect 15800 -23544 15860 -23538
rect 17834 -23544 17894 -23538
rect 19868 -23544 19928 -23538
rect 21910 -23544 21970 -23538
rect 22422 -23544 22482 -23538
rect 22928 -23544 22988 -23538
rect 14010 -23602 15800 -23544
rect 11650 -23604 15800 -23602
rect 15860 -23604 17834 -23544
rect 17894 -23604 19868 -23544
rect 19928 -23604 21910 -23544
rect 21970 -23604 22422 -23544
rect 22482 -23604 22928 -23544
rect 1400 -23606 1636 -23604
rect -8194 -23676 -6368 -23616
rect -6308 -23676 -4498 -23616
rect -4438 -23676 -3036 -23616
rect -2670 -23620 -2610 -23614
rect -1976 -23620 -1916 -23614
rect -1080 -23620 -1020 -23614
rect -786 -23620 -726 -23614
rect 108 -23620 168 -23614
rect 410 -23620 470 -23614
rect -8254 -23682 -8194 -23676
rect -6368 -23682 -6308 -23676
rect -4498 -23682 -4438 -23676
rect -2610 -23680 -1976 -23620
rect -1916 -23680 -1080 -23620
rect -1020 -23680 -786 -23620
rect -726 -23680 108 -23620
rect 168 -23680 410 -23620
rect -2670 -23686 -2610 -23680
rect -1976 -23686 -1916 -23680
rect -1080 -23686 -1020 -23680
rect -786 -23686 -726 -23680
rect 108 -23686 168 -23680
rect 410 -23686 470 -23680
rect -8402 -23724 -8342 -23718
rect -6366 -23724 -6306 -23718
rect -4330 -23724 -4270 -23718
rect -8342 -23784 -6366 -23724
rect -6306 -23784 -4330 -23724
rect -8402 -23790 -8342 -23784
rect -6366 -23790 -6306 -23784
rect -4330 -23790 -4270 -23784
rect -1530 -23728 -1470 -23722
rect -336 -23728 -276 -23722
rect -1470 -23788 -336 -23728
rect -276 -23788 952 -23728
rect 1012 -23788 1018 -23728
rect -1530 -23794 -1470 -23788
rect -336 -23794 -276 -23788
rect -7384 -23836 -7324 -23830
rect -7324 -23896 -5346 -23836
rect -5286 -23896 -5280 -23836
rect -7384 -23902 -7324 -23896
rect -1828 -24712 -1768 -24706
rect -1234 -24712 -1174 -24706
rect -634 -24712 -574 -24706
rect -40 -24712 20 -24706
rect 554 -24712 614 -24706
rect 1400 -24712 1460 -23606
rect 1976 -23610 2036 -23604
rect 2568 -23610 2628 -23604
rect 3082 -23610 3142 -23604
rect 3580 -23610 3640 -23604
rect 5622 -23610 5682 -23604
rect 7654 -23610 7714 -23604
rect 9686 -23610 9746 -23604
rect 15800 -23610 15860 -23604
rect 17834 -23610 17894 -23604
rect 19868 -23610 19928 -23604
rect 21910 -23610 21970 -23604
rect 22422 -23610 22482 -23604
rect 22928 -23610 22988 -23604
rect 6130 -23656 6190 -23650
rect 7142 -23656 7202 -23650
rect 8156 -23656 8216 -23650
rect 11068 -23656 11128 -23650
rect 6190 -23716 7142 -23656
rect 7202 -23716 8156 -23656
rect 8216 -23716 11068 -23656
rect 6130 -23722 6190 -23716
rect 7142 -23722 7202 -23716
rect 8156 -23722 8216 -23716
rect 11068 -23722 11128 -23716
rect 11728 -23654 11788 -23648
rect 2110 -23762 2170 -23756
rect 4096 -23762 4156 -23756
rect 5118 -23762 5178 -23756
rect 7656 -23762 7716 -23756
rect 8168 -23762 8228 -23756
rect 9186 -23762 9246 -23756
rect 9692 -23762 9752 -23756
rect 10198 -23762 10258 -23756
rect 11210 -23762 11270 -23756
rect 11728 -23762 11788 -23714
rect 12356 -23658 12416 -23652
rect 13402 -23658 13462 -23652
rect 17330 -23658 17390 -23652
rect 18348 -23658 18408 -23652
rect 12416 -23718 13402 -23658
rect 13462 -23718 17330 -23658
rect 17390 -23718 18348 -23658
rect 18408 -23718 19358 -23658
rect 19418 -23718 19424 -23658
rect 12356 -23724 12416 -23718
rect 13402 -23724 13462 -23718
rect 17330 -23724 17390 -23718
rect 18348 -23724 18408 -23718
rect 12230 -23762 12290 -23756
rect 13252 -23762 13312 -23756
rect 13764 -23762 13824 -23756
rect 14270 -23762 14330 -23756
rect 15288 -23762 15348 -23756
rect 15800 -23762 15860 -23756
rect 16308 -23762 16368 -23756
rect 20380 -23762 20440 -23756
rect 21382 -23762 21442 -23756
rect 2170 -23822 4096 -23762
rect 4156 -23822 5118 -23762
rect 5178 -23822 7656 -23762
rect 7716 -23822 8168 -23762
rect 8228 -23822 9186 -23762
rect 9246 -23822 9692 -23762
rect 9752 -23822 10198 -23762
rect 10258 -23822 11210 -23762
rect 11270 -23822 12230 -23762
rect 12290 -23822 13252 -23762
rect 13312 -23822 13764 -23762
rect 13824 -23822 14270 -23762
rect 14330 -23822 15288 -23762
rect 15348 -23822 15800 -23762
rect 15860 -23822 16308 -23762
rect 16368 -23822 20380 -23762
rect 20440 -23822 21382 -23762
rect 2110 -23828 2170 -23822
rect 4096 -23828 4156 -23822
rect 5118 -23828 5178 -23822
rect 7656 -23828 7716 -23822
rect 8168 -23828 8228 -23822
rect 9186 -23828 9246 -23822
rect 9692 -23828 9752 -23822
rect 10198 -23828 10258 -23822
rect 11210 -23828 11270 -23822
rect 12230 -23828 12290 -23822
rect 13252 -23828 13312 -23822
rect 13764 -23828 13824 -23822
rect 14270 -23828 14330 -23822
rect 15288 -23828 15348 -23822
rect 15800 -23828 15860 -23822
rect 16308 -23828 16368 -23822
rect 20380 -23828 20440 -23822
rect 21382 -23828 21442 -23822
rect 1704 -23866 1764 -23860
rect 6132 -23866 6192 -23860
rect 6636 -23866 6696 -23860
rect 7152 -23866 7212 -23860
rect 8674 -23866 8734 -23860
rect 10712 -23866 10772 -23860
rect 12748 -23866 12808 -23860
rect 14784 -23866 14844 -23860
rect 16816 -23866 16876 -23860
rect 17338 -23866 17398 -23860
rect 17838 -23866 17898 -23860
rect 18346 -23866 18406 -23860
rect 18854 -23866 18914 -23860
rect 19204 -23866 19264 -23860
rect 23806 -23866 23866 -23860
rect 1764 -23926 6132 -23866
rect 6192 -23926 6636 -23866
rect 6696 -23926 7152 -23866
rect 7212 -23926 8674 -23866
rect 8734 -23926 10712 -23866
rect 10772 -23926 12748 -23866
rect 12808 -23926 14784 -23866
rect 14844 -23926 16816 -23866
rect 16876 -23926 17338 -23866
rect 17398 -23926 17838 -23866
rect 17898 -23926 18346 -23866
rect 18406 -23926 18854 -23866
rect 18914 -23926 19204 -23866
rect 19264 -23926 23806 -23866
rect 1704 -23932 1764 -23926
rect 6132 -23932 6192 -23926
rect 6636 -23932 6696 -23926
rect 7152 -23932 7212 -23926
rect 8674 -23932 8734 -23926
rect 10712 -23932 10772 -23926
rect 12748 -23932 12808 -23926
rect 14784 -23932 14844 -23926
rect 16816 -23932 16876 -23926
rect 17338 -23932 17398 -23926
rect 17838 -23932 17898 -23926
rect 18346 -23932 18406 -23926
rect 18854 -23932 18914 -23926
rect 19204 -23932 19264 -23926
rect 23806 -23932 23866 -23926
rect -7382 -24718 -7322 -24712
rect -7322 -24778 -5352 -24718
rect -5292 -24778 -5286 -24718
rect -1768 -24772 -1234 -24712
rect -1174 -24772 -634 -24712
rect -574 -24772 -40 -24712
rect 20 -24772 554 -24712
rect 614 -24772 1460 -24712
rect -1828 -24778 -1768 -24772
rect -1234 -24778 -1174 -24772
rect -634 -24778 -574 -24772
rect -40 -24778 20 -24772
rect 554 -24778 614 -24772
rect -7382 -24784 -7322 -24778
rect 11730 -24798 11790 -24792
rect 13766 -24798 13826 -24792
rect -1534 -24806 -1474 -24800
rect -936 -24806 -876 -24800
rect -338 -24806 -278 -24800
rect 262 -24806 322 -24800
rect -8400 -24820 -8340 -24814
rect -4332 -24820 -4272 -24814
rect -3202 -24820 -3142 -24814
rect -8340 -24880 -4332 -24820
rect -4272 -24880 -3202 -24820
rect -2432 -24866 -2426 -24806
rect -2366 -24866 -1534 -24806
rect -1474 -24866 -936 -24806
rect -876 -24866 -338 -24806
rect -278 -24866 262 -24806
rect 11790 -24858 13766 -24798
rect 11730 -24864 11790 -24858
rect 13766 -24864 13826 -24858
rect -1534 -24872 -1474 -24866
rect -936 -24872 -876 -24866
rect -338 -24872 -278 -24866
rect 262 -24872 322 -24866
rect -8400 -24886 -8340 -24880
rect -4332 -24886 -4272 -24880
rect -3202 -24886 -3142 -24880
rect -1978 -24914 -1918 -24908
rect -1680 -24914 -1620 -24908
rect -1384 -24914 -1324 -24908
rect -1080 -24914 -1020 -24908
rect -784 -24914 -724 -24908
rect -486 -24914 -426 -24908
rect -190 -24914 -130 -24908
rect 106 -24914 166 -24908
rect 410 -24914 470 -24908
rect 1076 -24914 1136 -24908
rect -9538 -24926 -9478 -24920
rect -6366 -24926 -6306 -24920
rect -9478 -24986 -6366 -24926
rect -1918 -24974 -1680 -24914
rect -1620 -24974 -1384 -24914
rect -1324 -24974 -1080 -24914
rect -1020 -24974 -784 -24914
rect -724 -24974 -486 -24914
rect -426 -24974 -190 -24914
rect -130 -24974 106 -24914
rect 166 -24974 410 -24914
rect 470 -24974 1076 -24914
rect -1978 -24980 -1918 -24974
rect -1680 -24980 -1620 -24974
rect -1384 -24980 -1324 -24974
rect -1080 -24980 -1020 -24974
rect -784 -24980 -724 -24974
rect -486 -24980 -426 -24974
rect -190 -24980 -130 -24974
rect 106 -24980 166 -24974
rect 410 -24980 470 -24974
rect 1076 -24980 1136 -24974
rect -9538 -24992 -9478 -24986
rect -6366 -24992 -6306 -24986
rect 3580 -24998 3640 -24992
rect 5618 -24998 5678 -24992
rect 7656 -24998 7716 -24992
rect 9688 -24998 9748 -24992
rect 11726 -24998 11786 -24992
rect 13760 -24998 13820 -24992
rect 15800 -24998 15860 -24992
rect 17834 -24998 17894 -24992
rect 19868 -24998 19928 -24992
rect 21906 -24998 21966 -24992
rect 23648 -24998 23708 -24992
rect 3640 -25058 5618 -24998
rect 5678 -25058 7656 -24998
rect 7716 -25058 9688 -24998
rect 9748 -25058 11726 -24998
rect 11786 -25058 13760 -24998
rect 13820 -25058 15800 -24998
rect 15860 -25058 17834 -24998
rect 17894 -25058 19868 -24998
rect 19928 -25058 21906 -24998
rect 21966 -25058 23648 -24998
rect 3580 -25064 3640 -25058
rect 5618 -25064 5678 -25058
rect 7656 -25064 7716 -25058
rect 9688 -25064 9748 -25058
rect 11726 -25064 11786 -25058
rect 13760 -25064 13820 -25058
rect 15800 -25064 15860 -25058
rect 17834 -25064 17894 -25058
rect 19868 -25064 19928 -25058
rect 21906 -25064 21966 -25058
rect 23648 -25064 23708 -25058
rect 2568 -25096 2628 -25090
rect 4598 -25096 4658 -25090
rect 6636 -25096 6696 -25090
rect 8672 -25096 8732 -25090
rect 10708 -25096 10768 -25090
rect 12744 -25096 12804 -25090
rect 14778 -25096 14838 -25090
rect 16814 -25096 16874 -25090
rect 18854 -25096 18914 -25090
rect 20888 -25096 20948 -25090
rect 22924 -25096 22984 -25090
rect 2628 -25156 4598 -25096
rect 4658 -25156 6636 -25096
rect 6696 -25156 8672 -25096
rect 8732 -25156 10708 -25096
rect 10768 -25156 12744 -25096
rect 12804 -25156 14778 -25096
rect 14838 -25156 16814 -25096
rect 16874 -25156 18854 -25096
rect 18914 -25156 20888 -25096
rect 20948 -25156 22924 -25096
rect 2568 -25162 2628 -25156
rect 4598 -25162 4658 -25156
rect 6636 -25162 6696 -25156
rect 8672 -25162 8732 -25156
rect 10708 -25162 10768 -25156
rect 12744 -25162 12804 -25156
rect 14778 -25162 14838 -25156
rect 16814 -25162 16874 -25156
rect 18854 -25162 18914 -25156
rect 20888 -25162 20948 -25156
rect 22924 -25162 22984 -25156
rect -2670 -25840 -2610 -25834
rect -1680 -25840 -1620 -25834
rect -1382 -25840 -1322 -25834
rect -486 -25840 -426 -25834
rect -184 -25840 -124 -25834
rect -7896 -25870 -7836 -25864
rect -6870 -25870 -6810 -25864
rect -5846 -25870 -5786 -25864
rect -7836 -25930 -6870 -25870
rect -6810 -25930 -5846 -25870
rect -5786 -25930 -4946 -25870
rect -4886 -25930 -4880 -25870
rect -2610 -25900 -1680 -25840
rect -1620 -25900 -1382 -25840
rect -1322 -25900 -486 -25840
rect -426 -25900 -184 -25840
rect -2670 -25906 -2610 -25900
rect -1680 -25906 -1620 -25900
rect -1382 -25906 -1322 -25900
rect -486 -25906 -426 -25900
rect -184 -25906 -124 -25900
rect -7896 -25936 -7836 -25930
rect -6870 -25936 -6810 -25930
rect -5846 -25936 -5786 -25930
rect -2126 -25940 -2066 -25934
rect -938 -25940 -878 -25934
rect 258 -25940 318 -25934
rect 952 -25940 1012 -25934
rect -2066 -26000 -938 -25940
rect -878 -26000 258 -25940
rect 318 -26000 952 -25940
rect -2126 -26006 -2066 -26000
rect -938 -26006 -878 -26000
rect 258 -26006 318 -26000
rect 952 -26006 1012 -26000
rect -7518 -26476 23968 -26430
rect -7518 -26630 -7472 -26476
rect 23928 -26630 23968 -26476
rect -7518 -26676 23968 -26630
rect -12216 -26816 -11616 -26806
rect -12216 -27126 -11616 -27116
rect 24216 -26816 24816 -26806
rect 24216 -27126 24816 -27116
<< via2 >>
rect 484 1316 1084 1616
rect 24116 1316 24716 1616
rect 4061 1020 20846 1234
rect -12027 -11273 -11937 -11183
rect -10233 -11273 -10143 -11183
rect -7633 -11273 -7543 -11183
rect -5033 -11271 -4943 -11181
rect -2433 -11271 -2343 -11181
rect -629 -11271 -539 -11181
rect 2327 -7717 2417 -7627
rect 1705 -10213 1795 -10123
rect -7472 -26630 23928 -26476
rect -12216 -27116 -11616 -26816
rect 24216 -27116 24816 -26816
<< metal3 >>
rect 474 1616 1094 1621
rect 474 1316 484 1616
rect 1084 1316 1094 1616
rect 474 1311 1094 1316
rect 24106 1616 24726 1621
rect 24106 1316 24116 1616
rect 24716 1316 24726 1616
rect 24106 1311 24726 1316
rect 3998 1234 20878 1266
rect 3998 1020 4061 1234
rect 20846 1020 20878 1234
rect 3998 1000 20878 1020
rect 3998 998 8352 1000
rect -10238 -1378 -10138 32
rect -11658 -1478 -8642 -1378
rect -10238 -2894 -10138 -1478
rect -7638 -2894 -7538 48
rect -6524 -1478 -6042 -1378
rect -5038 -2894 -4938 26
rect -2438 -1378 -2338 22
rect -3924 -1478 -818 -1378
rect -2438 -2894 -2338 -1478
rect -11678 -3978 -8642 -3878
rect -6524 -3978 -6042 -3878
rect -3924 -3978 -812 -3878
rect -10238 -5394 -10138 -4982
rect -7638 -5394 -7538 -4982
rect -5038 -5394 -4938 -4982
rect -2438 -5394 -2338 -4982
rect -11678 -6478 -8642 -6378
rect -6524 -6478 -6042 -6378
rect -3924 -6478 -850 -6378
rect -10238 -8878 -10138 -7482
rect -11674 -8978 -8642 -8878
rect -12032 -11183 -11932 -10854
rect -12032 -11273 -12027 -11183
rect -11937 -11273 -11932 -11183
rect -12032 -11278 -11932 -11273
rect -10238 -11183 -10138 -8978
rect -10238 -11273 -10233 -11183
rect -10143 -11273 -10138 -11183
rect -10238 -11278 -10138 -11273
rect -7638 -11183 -7538 -7482
rect -6524 -8978 -6042 -8878
rect -7638 -11273 -7633 -11183
rect -7543 -11273 -7538 -11183
rect -7638 -11278 -7538 -11273
rect -5038 -11181 -4938 -7482
rect -2438 -8878 -2338 -7482
rect -1749 -7622 -1651 -7617
rect -1750 -7623 2422 -7622
rect -1750 -7721 -1749 -7623
rect -1651 -7627 2422 -7623
rect -1651 -7717 2327 -7627
rect 2417 -7717 2422 -7627
rect -1651 -7721 2422 -7717
rect -1750 -7722 2422 -7721
rect -1749 -7727 -1651 -7722
rect -3924 -8978 -844 -8878
rect -5038 -11271 -5033 -11181
rect -4943 -11271 -4938 -11181
rect -5038 -11276 -4938 -11271
rect -2438 -11181 -2338 -8978
rect -1089 -10118 -991 -10113
rect -1090 -10119 1800 -10118
rect -1090 -10217 -1089 -10119
rect -991 -10123 1800 -10119
rect -991 -10213 1705 -10123
rect 1795 -10213 1800 -10123
rect -991 -10217 1800 -10213
rect -1090 -10218 1800 -10217
rect -1089 -10223 -991 -10218
rect -2438 -11271 -2433 -11181
rect -2343 -11271 -2338 -11181
rect -2438 -11276 -2338 -11271
rect -634 -11181 -534 -10856
rect -634 -11271 -629 -11181
rect -539 -11271 -534 -11181
rect -634 -11276 -534 -11271
rect -7518 -26476 23968 -26430
rect -7518 -26630 -7472 -26476
rect 23928 -26630 23968 -26476
rect -7518 -26676 23968 -26630
rect -12226 -26816 -11606 -26811
rect -12226 -27116 -12216 -26816
rect -11616 -27116 -11606 -26816
rect -12226 -27121 -11606 -27116
rect 24206 -26816 24826 -26811
rect 24206 -27116 24216 -26816
rect 24816 -27116 24826 -26816
rect 24206 -27121 24826 -27116
<< via3 >>
rect 484 1316 1084 1616
rect 24116 1316 24716 1616
rect 4061 1020 20846 1234
rect -1749 -7721 -1651 -7623
rect -1089 -10217 -991 -10119
rect -7472 -26630 23928 -26476
rect -12216 -27116 -11616 -26816
rect 24216 -27116 24816 -26816
<< metal4 >>
rect -12400 1616 25000 1800
rect -12400 1316 484 1616
rect 1084 1316 24116 1616
rect 24716 1316 25000 1616
rect -12400 1234 25000 1316
rect -12400 1020 4061 1234
rect 20846 1020 25000 1234
rect -12400 1000 25000 1020
rect -12032 226 -186 326
rect -12032 -10566 -11932 226
rect -11680 -10566 -11580 226
rect -10230 -220 -992 -120
rect -10230 -542 -10130 -220
rect -5000 -566 -4900 -220
rect -7608 -2622 -7508 -2200
rect -2424 -2622 -2324 -2240
rect -11478 -2722 -2324 -2622
rect -11478 -7622 -11378 -2722
rect -10238 -3078 -10138 -2722
rect -5000 -3078 -4900 -2722
rect -7622 -5122 -7522 -4754
rect -2432 -5122 -2332 -4746
rect -1092 -5122 -992 -220
rect -10246 -5222 -992 -5122
rect -10246 -5600 -10146 -5222
rect -5008 -5592 -4908 -5222
rect -7630 -7622 -7530 -7266
rect -2440 -7622 -2340 -7242
rect -11478 -7623 -1650 -7622
rect -11478 -7721 -1749 -7623
rect -1651 -7721 -1650 -7623
rect -11478 -7722 -1650 -7721
rect -10254 -8080 -10154 -7722
rect -5008 -8096 -4908 -7722
rect -7646 -10118 -7546 -9780
rect -2440 -10118 -2340 -9786
rect -1092 -10118 -992 -5222
rect -7646 -10119 -990 -10118
rect -7646 -10217 -1089 -10119
rect -991 -10217 -990 -10119
rect -7646 -10218 -990 -10217
rect -636 -10566 -536 226
rect -286 -10566 -186 226
rect -12032 -10666 -186 -10566
rect -12032 -10668 -11932 -10666
rect -11680 -10668 -11580 -10666
rect -636 -10668 -536 -10666
rect -286 -10668 -186 -10666
rect -12400 -26476 25000 -26400
rect -12400 -26630 -7472 -26476
rect 23928 -26630 25000 -26476
rect -12400 -26816 25000 -26630
rect -12400 -27116 -12216 -26816
rect -11616 -27116 24216 -26816
rect 24816 -27116 25000 -26816
rect -12400 -27200 25000 -27116
use sky130_fd_pr__nfet_01v8_Y4K3TH  sky130_fd_pr__nfet_01v8_Y4K3TH_3
timestamp 1624477805
transform 1 0 -6335 0 1 -25418
box -3083 -388 3083 388
use ptap  ptap_272 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/ptap
timestamp 1624477805
transform 1 0 -7994 0 1 -26218
box 70 126 186 240
use ptap  ptap_273
timestamp 1624477805
transform 1 0 -9012 0 1 -26218
box 70 126 186 240
use ptap  ptap_271
timestamp 1624477805
transform 1 0 -6976 0 1 -26218
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_lvt_DHUKXE  sky130_fd_pr__nfet_01v8_lvt_DHUKXE_3
timestamp 1624477805
transform 1 0 -756 0 1 -25414
box -1668 -388 1668 388
use ptap  ptap_270
timestamp 1624477805
transform 1 0 -5958 0 1 -26218
box 70 126 186 240
use ptap  ptap_268
timestamp 1624477805
transform 1 0 -3922 0 1 -26218
box 70 126 186 240
use ptap  ptap_269
timestamp 1624477805
transform 1 0 -4940 0 1 -26218
box 70 126 186 240
use ptap  ptap_234
timestamp 1624477805
transform 1 0 -1402 0 1 -26272
box 70 126 186 240
use ptap  ptap_235
timestamp 1624477805
transform 1 0 -2420 0 1 -26272
box 70 126 186 240
use ptap  ptap_233
timestamp 1624477805
transform 1 0 -384 0 1 -26272
box 70 126 186 240
use ptap  ptap_232
timestamp 1624477805
transform 1 0 634 0 1 -26272
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_11 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/se_fold_casc_wide_swing_ota
timestamp 1624477805
transform 1 0 12777 0 1 -25584
box -10209 -388 10209 388
use sky130_fd_pr__nfet_01v8_Y4K3TH  sky130_fd_pr__nfet_01v8_Y4K3TH_2
timestamp 1624477805
transform 1 0 -6334 0 1 -24305
box -3083 -388 3083 388
use ptap  ptap_265
timestamp 1624477805
transform 1 0 -6950 0 1 -25024
box 70 126 186 240
use ptap  ptap_266
timestamp 1624477805
transform 1 0 -7968 0 1 -25024
box 70 126 186 240
use ptap  ptap_267
timestamp 1624477805
transform 1 0 -8986 0 1 -25024
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_lvt_DHUKXE  sky130_fd_pr__nfet_01v8_lvt_DHUKXE_2
timestamp 1624477805
transform 1 0 -756 0 1 -24304
box -1668 -388 1668 388
use ptap  ptap_263
timestamp 1624477805
transform 1 0 -4914 0 1 -25024
box 70 126 186 240
use ptap  ptap_264
timestamp 1624477805
transform 1 0 -5932 0 1 -25024
box 70 126 186 240
use ptap  ptap_229
timestamp 1624477805
transform 1 0 -358 0 1 -25038
box 70 126 186 240
use ptap  ptap_230
timestamp 1624477805
transform 1 0 -1376 0 1 -25038
box 70 126 186 240
use ptap  ptap_231
timestamp 1624477805
transform 1 0 -2394 0 1 -25038
box 70 126 186 240
use ptap  ptap_262
timestamp 1624477805
transform 1 0 -3896 0 1 -25024
box 70 126 186 240
use ptap  ptap_228
timestamp 1624477805
transform 1 0 660 0 1 -25038
box 70 126 186 240
use ptap  ptap_214
timestamp 1624477805
transform 1 0 2978 0 1 -25132
box 70 126 186 240
use ptap  ptap_215
timestamp 1624477805
transform 1 0 3996 0 1 -25132
box 70 126 186 240
use ptap  ptap_216
timestamp 1624477805
transform 1 0 5014 0 1 -25132
box 70 126 186 240
use ptap  ptap_217
timestamp 1624477805
transform 1 0 6032 0 1 -25132
box 70 126 186 240
use ptap  ptap_218
timestamp 1624477805
transform 1 0 7050 0 1 -25132
box 70 126 186 240
use ptap  ptap_219
timestamp 1624477805
transform 1 0 8068 0 1 -25132
box 70 126 186 240
use ptap  ptap_200
timestamp 1624477805
transform 1 0 9086 0 1 -25132
box 70 126 186 240
use ptap  ptap_201
timestamp 1624477805
transform 1 0 10104 0 1 -25132
box 70 126 186 240
use ptap  ptap_202
timestamp 1624477805
transform 1 0 11122 0 1 -25132
box 70 126 186 240
use ptap  ptap_203
timestamp 1624477805
transform 1 0 12140 0 1 -25132
box 70 126 186 240
use ptap  ptap_204
timestamp 1624477805
transform 1 0 13158 0 1 -25132
box 70 126 186 240
use ptap  ptap_205
timestamp 1624477805
transform 1 0 14176 0 1 -25132
box 70 126 186 240
use ptap  ptap_206
timestamp 1624477805
transform 1 0 15194 0 1 -25132
box 70 126 186 240
use ptap  ptap_207
timestamp 1624477805
transform 1 0 16212 0 1 -25132
box 70 126 186 240
use ptap  ptap_208
timestamp 1624477805
transform 1 0 17230 0 1 -25132
box 70 126 186 240
use ptap  ptap_209
timestamp 1624477805
transform 1 0 18248 0 1 -25132
box 70 126 186 240
use ptap  ptap_210
timestamp 1624477805
transform 1 0 19266 0 1 -25132
box 70 126 186 240
use ptap  ptap_211
timestamp 1624477805
transform 1 0 20284 0 1 -25132
box 70 126 186 240
use ptap  ptap_212
timestamp 1624477805
transform 1 0 21302 0 1 -25132
box 70 126 186 240
use ptap  ptap_213
timestamp 1624477805
transform 1 0 22320 0 1 -25132
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_10
timestamp 1624477805
transform 1 0 12777 0 1 -24352
box -10209 -388 10209 388
use sky130_fd_pr__nfet_01v8_Y4K3TH  sky130_fd_pr__nfet_01v8_Y4K3TH_1
timestamp 1624477805
transform 1 0 -6335 0 1 -23194
box -3083 -388 3083 388
use ptap  ptap_259
timestamp 1624477805
transform 1 0 -6976 0 1 -23926
box 70 126 186 240
use ptap  ptap_260
timestamp 1624477805
transform 1 0 -7994 0 1 -23926
box 70 126 186 240
use ptap  ptap_261
timestamp 1624477805
transform 1 0 -9012 0 1 -23926
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_lvt_DHUKXE  sky130_fd_pr__nfet_01v8_lvt_DHUKXE_1
timestamp 1624477805
transform 1 0 -754 0 1 -23192
box -1668 -388 1668 388
use ptap  ptap_257
timestamp 1624477805
transform 1 0 -4940 0 1 -23926
box 70 126 186 240
use ptap  ptap_258
timestamp 1624477805
transform 1 0 -5958 0 1 -23926
box 70 126 186 240
use ptap  ptap_225
timestamp 1624477805
transform 1 0 -412 0 1 -23926
box 70 126 186 240
use ptap  ptap_226
timestamp 1624477805
transform 1 0 -1430 0 1 -23926
box 70 126 186 240
use ptap  ptap_227
timestamp 1624477805
transform 1 0 -2448 0 1 -23926
box 70 126 186 240
use ptap  ptap_256
timestamp 1624477805
transform 1 0 -3922 0 1 -23926
box 70 126 186 240
use ptap  ptap_224
timestamp 1624477805
transform 1 0 606 0 1 -23926
box 70 126 186 240
use ptap  ptap_194
timestamp 1624477805
transform 1 0 2978 0 1 -23912
box 70 126 186 240
use ptap  ptap_196
timestamp 1624477805
transform 1 0 5014 0 1 -23912
box 70 126 186 240
use ptap  ptap_195
timestamp 1624477805
transform 1 0 3996 0 1 -23912
box 70 126 186 240
use ptap  ptap_197
timestamp 1624477805
transform 1 0 6032 0 1 -23912
box 70 126 186 240
use ptap  ptap_198
timestamp 1624477805
transform 1 0 7050 0 1 -23912
box 70 126 186 240
use ptap  ptap_199
timestamp 1624477805
transform 1 0 8068 0 1 -23912
box 70 126 186 240
use ptap  ptap_180
timestamp 1624477805
transform 1 0 9086 0 1 -23912
box 70 126 186 240
use ptap  ptap_181
timestamp 1624477805
transform 1 0 10104 0 1 -23912
box 70 126 186 240
use ptap  ptap_182
timestamp 1624477805
transform 1 0 11122 0 1 -23912
box 70 126 186 240
use ptap  ptap_183
timestamp 1624477805
transform 1 0 12140 0 1 -23912
box 70 126 186 240
use ptap  ptap_184
timestamp 1624477805
transform 1 0 13158 0 1 -23912
box 70 126 186 240
use ptap  ptap_185
timestamp 1624477805
transform 1 0 14176 0 1 -23912
box 70 126 186 240
use ptap  ptap_186
timestamp 1624477805
transform 1 0 15194 0 1 -23912
box 70 126 186 240
use ptap  ptap_187
timestamp 1624477805
transform 1 0 16212 0 1 -23912
box 70 126 186 240
use ptap  ptap_188
timestamp 1624477805
transform 1 0 17230 0 1 -23912
box 70 126 186 240
use ptap  ptap_189
timestamp 1624477805
transform 1 0 18248 0 1 -23912
box 70 126 186 240
use ptap  ptap_190
timestamp 1624477805
transform 1 0 19266 0 1 -23912
box 70 126 186 240
use ptap  ptap_191
timestamp 1624477805
transform 1 0 20284 0 1 -23912
box 70 126 186 240
use ptap  ptap_192
timestamp 1624477805
transform 1 0 21302 0 1 -23912
box 70 126 186 240
use ptap  ptap_193
timestamp 1624477805
transform 1 0 22320 0 1 -23912
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_9
timestamp 1624477805
transform 1 0 12777 0 1 -23118
box -10209 -388 10209 388
use sky130_fd_pr__nfet_01v8_Y4K3TH  sky130_fd_pr__nfet_01v8_Y4K3TH_0
timestamp 1624477805
transform 1 0 -6334 0 1 -22081
box -3083 -388 3083 388
use ptap  ptap_255
timestamp 1624477805
transform 1 0 -8986 0 1 -22800
box 70 126 186 240
use ptap  ptap_254
timestamp 1624477805
transform 1 0 -7968 0 1 -22800
box 70 126 186 240
use ptap  ptap_253
timestamp 1624477805
transform 1 0 -6950 0 1 -22800
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_lvt_DHUKXE  sky130_fd_pr__nfet_01v8_lvt_DHUKXE_0
timestamp 1624477805
transform 1 0 -754 0 1 -22080
box -1668 -388 1668 388
use ptap  ptap_252
timestamp 1624477805
transform 1 0 -5932 0 1 -22800
box 70 126 186 240
use ptap  ptap_251
timestamp 1624477805
transform 1 0 -4914 0 1 -22800
box 70 126 186 240
use ptap  ptap_250
timestamp 1624477805
transform 1 0 -3896 0 1 -22800
box 70 126 186 240
use ptap  ptap_223
timestamp 1624477805
transform 1 0 -2448 0 1 -22812
box 70 126 186 240
use ptap  ptap_222
timestamp 1624477805
transform 1 0 -1430 0 1 -22812
box 70 126 186 240
use ptap  ptap_221
timestamp 1624477805
transform 1 0 -412 0 1 -22812
box 70 126 186 240
use ptap  ptap_220
timestamp 1624477805
transform 1 0 606 0 1 -22812
box 70 126 186 240
use ptap  ptap_174
timestamp 1624477805
transform 1 0 2992 0 1 -22690
box 70 126 186 240
use ptap  ptap_175
timestamp 1624477805
transform 1 0 4010 0 1 -22690
box 70 126 186 240
use ptap  ptap_176
timestamp 1624477805
transform 1 0 5028 0 1 -22690
box 70 126 186 240
use ptap  ptap_177
timestamp 1624477805
transform 1 0 6046 0 1 -22690
box 70 126 186 240
use ptap  ptap_178
timestamp 1624477805
transform 1 0 7064 0 1 -22690
box 70 126 186 240
use ptap  ptap_179
timestamp 1624477805
transform 1 0 8082 0 1 -22690
box 70 126 186 240
use ptap  ptap_160
timestamp 1624477805
transform 1 0 9100 0 1 -22690
box 70 126 186 240
use ptap  ptap_161
timestamp 1624477805
transform 1 0 10118 0 1 -22690
box 70 126 186 240
use ptap  ptap_162
timestamp 1624477805
transform 1 0 11136 0 1 -22690
box 70 126 186 240
use ptap  ptap_163
timestamp 1624477805
transform 1 0 12154 0 1 -22690
box 70 126 186 240
use ptap  ptap_164
timestamp 1624477805
transform 1 0 13172 0 1 -22690
box 70 126 186 240
use ptap  ptap_165
timestamp 1624477805
transform 1 0 14190 0 1 -22690
box 70 126 186 240
use ptap  ptap_166
timestamp 1624477805
transform 1 0 15208 0 1 -22690
box 70 126 186 240
use ptap  ptap_167
timestamp 1624477805
transform 1 0 16226 0 1 -22690
box 70 126 186 240
use ptap  ptap_168
timestamp 1624477805
transform 1 0 17244 0 1 -22690
box 70 126 186 240
use ptap  ptap_169
timestamp 1624477805
transform 1 0 18262 0 1 -22690
box 70 126 186 240
use ptap  ptap_170
timestamp 1624477805
transform 1 0 19280 0 1 -22690
box 70 126 186 240
use ptap  ptap_171
timestamp 1624477805
transform 1 0 20298 0 1 -22690
box 70 126 186 240
use ptap  ptap_172
timestamp 1624477805
transform 1 0 21316 0 1 -22690
box 70 126 186 240
use ptap  ptap_173
timestamp 1624477805
transform 1 0 22334 0 1 -22690
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_5
timestamp 1624477805
transform 1 0 12777 0 1 -21884
box -10209 -388 10209 388
use ptap  ptap_249
timestamp 1624477805
transform 1 0 -9000 0 1 -21674
box 70 126 186 240
use ptap  ptap_247
timestamp 1624477805
transform 1 0 -6964 0 1 -21674
box 70 126 186 240
use ptap  ptap_246
timestamp 1624477805
transform 1 0 -5946 0 1 -21674
box 70 126 186 240
use ptap  ptap_248
timestamp 1624477805
transform 1 0 -7982 0 1 -21674
box 70 126 186 240
use ptap  ptap_239
timestamp 1624477805
transform 1 0 -2408 0 1 -21618
box 70 126 186 240
use ptap  ptap_245
timestamp 1624477805
transform 1 0 -4928 0 1 -21674
box 70 126 186 240
use ptap  ptap_244
timestamp 1624477805
transform 1 0 -3910 0 1 -21674
box 70 126 186 240
use ptap  ptap_236
timestamp 1624477805
transform 1 0 646 0 1 -21618
box 70 126 186 240
use ptap  ptap_238
timestamp 1624477805
transform 1 0 -1390 0 1 -21618
box 70 126 186 240
use ptap  ptap_237
timestamp 1624477805
transform 1 0 -372 0 1 -21618
box 70 126 186 240
use ptap  ptap_154
timestamp 1624477805
transform 1 0 2992 0 1 -21442
box 70 126 186 240
use ptap  ptap_155
timestamp 1624477805
transform 1 0 4010 0 1 -21442
box 70 126 186 240
use ptap  ptap_156
timestamp 1624477805
transform 1 0 5028 0 1 -21442
box 70 126 186 240
use ptap  ptap_157
timestamp 1624477805
transform 1 0 6046 0 1 -21442
box 70 126 186 240
use ptap  ptap_158
timestamp 1624477805
transform 1 0 7064 0 1 -21442
box 70 126 186 240
use ptap  ptap_159
timestamp 1624477805
transform 1 0 8082 0 1 -21442
box 70 126 186 240
use ptap  ptap_140
timestamp 1624477805
transform 1 0 9100 0 1 -21442
box 70 126 186 240
use ptap  ptap_141
timestamp 1624477805
transform 1 0 10118 0 1 -21442
box 70 126 186 240
use ptap  ptap_142
timestamp 1624477805
transform 1 0 11136 0 1 -21442
box 70 126 186 240
use ptap  ptap_143
timestamp 1624477805
transform 1 0 12154 0 1 -21442
box 70 126 186 240
use ptap  ptap_144
timestamp 1624477805
transform 1 0 13172 0 1 -21442
box 70 126 186 240
use ptap  ptap_145
timestamp 1624477805
transform 1 0 14190 0 1 -21442
box 70 126 186 240
use ptap  ptap_146
timestamp 1624477805
transform 1 0 15208 0 1 -21442
box 70 126 186 240
use ptap  ptap_147
timestamp 1624477805
transform 1 0 16226 0 1 -21442
box 70 126 186 240
use ptap  ptap_148
timestamp 1624477805
transform 1 0 17244 0 1 -21442
box 70 126 186 240
use ptap  ptap_149
timestamp 1624477805
transform 1 0 18262 0 1 -21442
box 70 126 186 240
use ptap  ptap_150
timestamp 1624477805
transform 1 0 19280 0 1 -21442
box 70 126 186 240
use ptap  ptap_151
timestamp 1624477805
transform 1 0 20298 0 1 -21442
box 70 126 186 240
use ptap  ptap_152
timestamp 1624477805
transform 1 0 21316 0 1 -21442
box 70 126 186 240
use ptap  ptap_153
timestamp 1624477805
transform 1 0 22334 0 1 -21442
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_lvt_LYGCX9  sky130_fd_pr__nfet_01v8_lvt_LYGCX9_1
timestamp 1624477805
transform 1 0 -1217 0 1 -20554
box -1119 -188 1119 188
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_4
timestamp 1624477805
transform 1 0 12777 0 1 -20652
box -10209 -388 10209 388
use ptap  ptap_242
timestamp 1624477805
transform 1 0 -1688 0 1 -20330
box 70 126 186 240
use ptap  ptap_243
timestamp 1624477805
transform 1 0 -2706 0 1 -20330
box 70 126 186 240
use ptap  ptap_240
timestamp 1624477805
transform 1 0 348 0 1 -20330
box 70 126 186 240
use ptap  ptap_241
timestamp 1624477805
transform 1 0 -670 0 1 -20330
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_lvt_LYGCX9  sky130_fd_pr__nfet_01v8_lvt_LYGCX9_0
timestamp 1624477805
transform 1 0 -1217 0 1 -19722
box -1119 -188 1119 188
use ptap  ptap_134
timestamp 1624477805
transform 1 0 2978 0 1 -20222
box 70 126 186 240
use ptap  ptap_136
timestamp 1624477805
transform 1 0 5014 0 1 -20222
box 70 126 186 240
use ptap  ptap_135
timestamp 1624477805
transform 1 0 3996 0 1 -20222
box 70 126 186 240
use ptap  ptap_138
timestamp 1624477805
transform 1 0 7050 0 1 -20222
box 70 126 186 240
use ptap  ptap_137
timestamp 1624477805
transform 1 0 6032 0 1 -20222
box 70 126 186 240
use ptap  ptap_120
timestamp 1624477805
transform 1 0 9086 0 1 -20222
box 70 126 186 240
use ptap  ptap_139
timestamp 1624477805
transform 1 0 8068 0 1 -20222
box 70 126 186 240
use ptap  ptap_123
timestamp 1624477805
transform 1 0 12140 0 1 -20222
box 70 126 186 240
use ptap  ptap_122
timestamp 1624477805
transform 1 0 11122 0 1 -20222
box 70 126 186 240
use ptap  ptap_121
timestamp 1624477805
transform 1 0 10104 0 1 -20222
box 70 126 186 240
use ptap  ptap_125
timestamp 1624477805
transform 1 0 14176 0 1 -20222
box 70 126 186 240
use ptap  ptap_124
timestamp 1624477805
transform 1 0 13158 0 1 -20222
box 70 126 186 240
use ptap  ptap_127
timestamp 1624477805
transform 1 0 16212 0 1 -20222
box 70 126 186 240
use ptap  ptap_126
timestamp 1624477805
transform 1 0 15194 0 1 -20222
box 70 126 186 240
use ptap  ptap_129
timestamp 1624477805
transform 1 0 18248 0 1 -20222
box 70 126 186 240
use ptap  ptap_128
timestamp 1624477805
transform 1 0 17230 0 1 -20222
box 70 126 186 240
use ptap  ptap_131
timestamp 1624477805
transform 1 0 20284 0 1 -20222
box 70 126 186 240
use ptap  ptap_130
timestamp 1624477805
transform 1 0 19266 0 1 -20222
box 70 126 186 240
use ptap  ptap_133
timestamp 1624477805
transform 1 0 22320 0 1 -20222
box 70 126 186 240
use ptap  ptap_132
timestamp 1624477805
transform 1 0 21302 0 1 -20222
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_3
timestamp 1624477805
transform 1 0 12777 0 1 -19418
box -10209 -388 10209 388
use ptap  ptap_282
timestamp 1624477805
transform 1 0 -8784 0 1 -19354
box 70 126 186 240
use ptap  ptap_281
timestamp 1624477805
transform 1 0 -7766 0 1 -19354
box 70 126 186 240
use ptap  ptap_280
timestamp 1624477805
transform 1 0 -6748 0 1 -19354
box 70 126 186 240
use ptap  ptap_279
timestamp 1624477805
transform 1 0 -5730 0 1 -19354
box 70 126 186 240
use ptap  ptap_278
timestamp 1624477805
transform 1 0 -4712 0 1 -19354
box 70 126 186 240
use ptap  ptap_277
timestamp 1624477805
transform 1 0 -3694 0 1 -19354
box 70 126 186 240
use ptap  ptap_276
timestamp 1624477805
transform 1 0 -2676 0 1 -19354
box 70 126 186 240
use ptap  ptap_275
timestamp 1624477805
transform 1 0 -1658 0 1 -19354
box 70 126 186 240
use ptap  ptap_274
timestamp 1624477805
transform 1 0 -640 0 1 -19354
box 70 126 186 240
use ptap  ptap_114
timestamp 1624477805
transform 1 0 2978 0 1 -18974
box 70 126 186 240
use ptap  ptap_115
timestamp 1624477805
transform 1 0 3996 0 1 -18974
box 70 126 186 240
use ptap  ptap_116
timestamp 1624477805
transform 1 0 5014 0 1 -18974
box 70 126 186 240
use ptap  ptap_117
timestamp 1624477805
transform 1 0 6032 0 1 -18974
box 70 126 186 240
use ptap  ptap_118
timestamp 1624477805
transform 1 0 7050 0 1 -18974
box 70 126 186 240
use ptap  ptap_119
timestamp 1624477805
transform 1 0 8068 0 1 -18974
box 70 126 186 240
use ptap  ptap_100
timestamp 1624477805
transform 1 0 9086 0 1 -18974
box 70 126 186 240
use ptap  ptap_101
timestamp 1624477805
transform 1 0 10104 0 1 -18974
box 70 126 186 240
use ptap  ptap_102
timestamp 1624477805
transform 1 0 11122 0 1 -18974
box 70 126 186 240
use ptap  ptap_103
timestamp 1624477805
transform 1 0 12140 0 1 -18974
box 70 126 186 240
use ptap  ptap_104
timestamp 1624477805
transform 1 0 13158 0 1 -18974
box 70 126 186 240
use ptap  ptap_106
timestamp 1624477805
transform 1 0 15194 0 1 -18974
box 70 126 186 240
use ptap  ptap_105
timestamp 1624477805
transform 1 0 14176 0 1 -18974
box 70 126 186 240
use ptap  ptap_108
timestamp 1624477805
transform 1 0 17230 0 1 -18974
box 70 126 186 240
use ptap  ptap_107
timestamp 1624477805
transform 1 0 16212 0 1 -18974
box 70 126 186 240
use ptap  ptap_110
timestamp 1624477805
transform 1 0 19266 0 1 -18974
box 70 126 186 240
use ptap  ptap_109
timestamp 1624477805
transform 1 0 18248 0 1 -18974
box 70 126 186 240
use ptap  ptap_111
timestamp 1624477805
transform 1 0 20284 0 1 -18974
box 70 126 186 240
use ptap  ptap_113
timestamp 1624477805
transform 1 0 22320 0 1 -18974
box 70 126 186 240
use ptap  ptap_112
timestamp 1624477805
transform 1 0 21302 0 1 -18974
box 70 126 186 240
use ptap  ptap_352
timestamp 1624477805
transform 1 0 -9294 0 1 -18312
box 70 126 186 240
use ptap  ptap_355
timestamp 1624477805
transform 1 0 -6240 0 1 -18312
box 70 126 186 240
use ptap  ptap_354
timestamp 1624477805
transform 1 0 -7258 0 1 -18312
box 70 126 186 240
use ptap  ptap_353
timestamp 1624477805
transform 1 0 -8276 0 1 -18312
box 70 126 186 240
use ptap  ptap_359
timestamp 1624477805
transform 1 0 -2168 0 1 -18312
box 70 126 186 240
use ptap  ptap_358
timestamp 1624477805
transform 1 0 -3186 0 1 -18312
box 70 126 186 240
use ptap  ptap_357
timestamp 1624477805
transform 1 0 -4204 0 1 -18312
box 70 126 186 240
use ptap  ptap_356
timestamp 1624477805
transform 1 0 -5222 0 1 -18312
box 70 126 186 240
use ptap  ptap_361
timestamp 1624477805
transform 1 0 -132 0 1 -18312
box 70 126 186 240
use ptap  ptap_360
timestamp 1624477805
transform 1 0 -1150 0 1 -18312
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_2
timestamp 1624477805
transform 1 0 12777 0 1 -18184
box -10209 -388 10209 388
use ptap  ptap_342
timestamp 1624477805
transform 1 0 -9294 0 1 -17494
box 70 126 186 240
use ptap  ptap_343
timestamp 1624477805
transform 1 0 -8276 0 1 -17494
box 70 126 186 240
use ptap  ptap_344
timestamp 1624477805
transform 1 0 -7258 0 1 -17494
box 70 126 186 240
use ptap  ptap_345
timestamp 1624477805
transform 1 0 -6240 0 1 -17494
box 70 126 186 240
use ptap  ptap_347
timestamp 1624477805
transform 1 0 -4204 0 1 -17494
box 70 126 186 240
use ptap  ptap_346
timestamp 1624477805
transform 1 0 -5222 0 1 -17494
box 70 126 186 240
use ptap  ptap_348
timestamp 1624477805
transform 1 0 -3186 0 1 -17494
box 70 126 186 240
use ptap  ptap_349
timestamp 1624477805
transform 1 0 -2168 0 1 -17494
box 70 126 186 240
use ptap  ptap_350
timestamp 1624477805
transform 1 0 -1150 0 1 -17494
box 70 126 186 240
use ptap  ptap_351
timestamp 1624477805
transform 1 0 -132 0 1 -17494
box 70 126 186 240
use ptap  ptap_95
timestamp 1624477805
transform 1 0 4010 0 1 -17752
box 70 126 186 240
use ptap  ptap_94
timestamp 1624477805
transform 1 0 2992 0 1 -17752
box 70 126 186 240
use ptap  ptap_96
timestamp 1624477805
transform 1 0 5028 0 1 -17752
box 70 126 186 240
use ptap  ptap_97
timestamp 1624477805
transform 1 0 6046 0 1 -17752
box 70 126 186 240
use ptap  ptap_98
timestamp 1624477805
transform 1 0 7064 0 1 -17752
box 70 126 186 240
use ptap  ptap_99
timestamp 1624477805
transform 1 0 8082 0 1 -17752
box 70 126 186 240
use ptap  ptap_80
timestamp 1624477805
transform 1 0 9100 0 1 -17752
box 70 126 186 240
use ptap  ptap_82
timestamp 1624477805
transform 1 0 11136 0 1 -17752
box 70 126 186 240
use ptap  ptap_81
timestamp 1624477805
transform 1 0 10118 0 1 -17752
box 70 126 186 240
use ptap  ptap_83
timestamp 1624477805
transform 1 0 12154 0 1 -17752
box 70 126 186 240
use ptap  ptap_84
timestamp 1624477805
transform 1 0 13172 0 1 -17752
box 70 126 186 240
use ptap  ptap_85
timestamp 1624477805
transform 1 0 14190 0 1 -17752
box 70 126 186 240
use ptap  ptap_86
timestamp 1624477805
transform 1 0 15208 0 1 -17752
box 70 126 186 240
use ptap  ptap_87
timestamp 1624477805
transform 1 0 16226 0 1 -17752
box 70 126 186 240
use ptap  ptap_88
timestamp 1624477805
transform 1 0 17244 0 1 -17752
box 70 126 186 240
use ptap  ptap_90
timestamp 1624477805
transform 1 0 19280 0 1 -17752
box 70 126 186 240
use ptap  ptap_89
timestamp 1624477805
transform 1 0 18262 0 1 -17752
box 70 126 186 240
use ptap  ptap_91
timestamp 1624477805
transform 1 0 20298 0 1 -17752
box 70 126 186 240
use ptap  ptap_92
timestamp 1624477805
transform 1 0 21316 0 1 -17752
box 70 126 186 240
use ptap  ptap_93
timestamp 1624477805
transform 1 0 22334 0 1 -17752
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_1
timestamp 1624477805
transform 1 0 12777 0 1 -16952
box -10209 -388 10209 388
use ptap  ptap_332
timestamp 1624477805
transform 1 0 -9294 0 1 -16676
box 70 126 186 240
use ptap  ptap_333
timestamp 1624477805
transform 1 0 -8276 0 1 -16676
box 70 126 186 240
use ptap  ptap_334
timestamp 1624477805
transform 1 0 -7258 0 1 -16676
box 70 126 186 240
use ptap  ptap_335
timestamp 1624477805
transform 1 0 -6240 0 1 -16676
box 70 126 186 240
use ptap  ptap_336
timestamp 1624477805
transform 1 0 -5222 0 1 -16676
box 70 126 186 240
use ptap  ptap_337
timestamp 1624477805
transform 1 0 -4204 0 1 -16676
box 70 126 186 240
use ptap  ptap_338
timestamp 1624477805
transform 1 0 -3186 0 1 -16676
box 70 126 186 240
use ptap  ptap_339
timestamp 1624477805
transform 1 0 -2168 0 1 -16676
box 70 126 186 240
use ptap  ptap_340
timestamp 1624477805
transform 1 0 -1150 0 1 -16676
box 70 126 186 240
use ptap  ptap_341
timestamp 1624477805
transform 1 0 -132 0 1 -16676
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_lvt_XH9Q8F  sky130_fd_pr__nfet_01v8_lvt_XH9Q8F_1 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/se_fold_casc_wide_swing_ota
timestamp 1624477805
transform 1 0 -4586 0 1 -17311
box -4610 -1615 4610 1615
use ptap  ptap_74
timestamp 1624477805
transform 1 0 2978 0 1 -16504
box 70 126 186 240
use ptap  ptap_76
timestamp 1624477805
transform 1 0 5014 0 1 -16504
box 70 126 186 240
use ptap  ptap_75
timestamp 1624477805
transform 1 0 3996 0 1 -16504
box 70 126 186 240
use ptap  ptap_77
timestamp 1624477805
transform 1 0 6032 0 1 -16504
box 70 126 186 240
use ptap  ptap_79
timestamp 1624477805
transform 1 0 8068 0 1 -16504
box 70 126 186 240
use ptap  ptap_78
timestamp 1624477805
transform 1 0 7050 0 1 -16504
box 70 126 186 240
use ptap  ptap_61
timestamp 1624477805
transform 1 0 10104 0 1 -16504
box 70 126 186 240
use ptap  ptap_60
timestamp 1624477805
transform 1 0 9086 0 1 -16504
box 70 126 186 240
use ptap  ptap_63
timestamp 1624477805
transform 1 0 12140 0 1 -16504
box 70 126 186 240
use ptap  ptap_62
timestamp 1624477805
transform 1 0 11122 0 1 -16504
box 70 126 186 240
use ptap  ptap_64
timestamp 1624477805
transform 1 0 13158 0 1 -16504
box 70 126 186 240
use ptap  ptap_66
timestamp 1624477805
transform 1 0 15194 0 1 -16504
box 70 126 186 240
use ptap  ptap_65
timestamp 1624477805
transform 1 0 14176 0 1 -16504
box 70 126 186 240
use ptap  ptap_68
timestamp 1624477805
transform 1 0 17230 0 1 -16504
box 70 126 186 240
use ptap  ptap_67
timestamp 1624477805
transform 1 0 16212 0 1 -16504
box 70 126 186 240
use ptap  ptap_70
timestamp 1624477805
transform 1 0 19266 0 1 -16504
box 70 126 186 240
use ptap  ptap_69
timestamp 1624477805
transform 1 0 18248 0 1 -16504
box 70 126 186 240
use ptap  ptap_71
timestamp 1624477805
transform 1 0 20284 0 1 -16504
box 70 126 186 240
use ptap  ptap_73
timestamp 1624477805
transform 1 0 22320 0 1 -16504
box 70 126 186 240
use ptap  ptap_72
timestamp 1624477805
transform 1 0 21302 0 1 -16504
box 70 126 186 240
use ptap  ptap_322
timestamp 1624477805
transform 1 0 -9294 0 1 -15858
box 70 126 186 240
use ptap  ptap_325
timestamp 1624477805
transform 1 0 -6240 0 1 -15858
box 70 126 186 240
use ptap  ptap_324
timestamp 1624477805
transform 1 0 -7258 0 1 -15858
box 70 126 186 240
use ptap  ptap_323
timestamp 1624477805
transform 1 0 -8276 0 1 -15858
box 70 126 186 240
use ptap  ptap_329
timestamp 1624477805
transform 1 0 -2168 0 1 -15858
box 70 126 186 240
use ptap  ptap_328
timestamp 1624477805
transform 1 0 -3186 0 1 -15858
box 70 126 186 240
use ptap  ptap_327
timestamp 1624477805
transform 1 0 -4204 0 1 -15858
box 70 126 186 240
use ptap  ptap_326
timestamp 1624477805
transform 1 0 -5222 0 1 -15858
box 70 126 186 240
use ptap  ptap_331
timestamp 1624477805
transform 1 0 -132 0 1 -15858
box 70 126 186 240
use ptap  ptap_330
timestamp 1624477805
transform 1 0 -1150 0 1 -15858
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_0
timestamp 1624477805
transform 1 0 12777 0 1 -15718
box -10209 -388 10209 388
use ptap  ptap_312
timestamp 1624477805
transform 1 0 -9294 0 1 -15040
box 70 126 186 240
use ptap  ptap_313
timestamp 1624477805
transform 1 0 -8276 0 1 -15040
box 70 126 186 240
use ptap  ptap_314
timestamp 1624477805
transform 1 0 -7258 0 1 -15040
box 70 126 186 240
use ptap  ptap_315
timestamp 1624477805
transform 1 0 -6240 0 1 -15040
box 70 126 186 240
use ptap  ptap_316
timestamp 1624477805
transform 1 0 -5222 0 1 -15040
box 70 126 186 240
use ptap  ptap_317
timestamp 1624477805
transform 1 0 -4204 0 1 -15040
box 70 126 186 240
use ptap  ptap_318
timestamp 1624477805
transform 1 0 -3186 0 1 -15040
box 70 126 186 240
use ptap  ptap_319
timestamp 1624477805
transform 1 0 -2168 0 1 -15040
box 70 126 186 240
use ptap  ptap_320
timestamp 1624477805
transform 1 0 -1150 0 1 -15040
box 70 126 186 240
use ptap  ptap_321
timestamp 1624477805
transform 1 0 -132 0 1 -15040
box 70 126 186 240
use ptap  ptap_54
timestamp 1624477805
transform 1 0 2978 0 1 -15284
box 70 126 186 240
use ptap  ptap_55
timestamp 1624477805
transform 1 0 3996 0 1 -15284
box 70 126 186 240
use ptap  ptap_56
timestamp 1624477805
transform 1 0 5014 0 1 -15284
box 70 126 186 240
use ptap  ptap_57
timestamp 1624477805
transform 1 0 6032 0 1 -15284
box 70 126 186 240
use ptap  ptap_58
timestamp 1624477805
transform 1 0 7050 0 1 -15284
box 70 126 186 240
use ptap  ptap_59
timestamp 1624477805
transform 1 0 8068 0 1 -15284
box 70 126 186 240
use ptap  ptap_40
timestamp 1624477805
transform 1 0 9086 0 1 -15284
box 70 126 186 240
use ptap  ptap_41
timestamp 1624477805
transform 1 0 10104 0 1 -15284
box 70 126 186 240
use ptap  ptap_42
timestamp 1624477805
transform 1 0 11122 0 1 -15284
box 70 126 186 240
use ptap  ptap_43
timestamp 1624477805
transform 1 0 12140 0 1 -15284
box 70 126 186 240
use ptap  ptap_44
timestamp 1624477805
transform 1 0 13158 0 1 -15284
box 70 126 186 240
use ptap  ptap_45
timestamp 1624477805
transform 1 0 14176 0 1 -15284
box 70 126 186 240
use ptap  ptap_46
timestamp 1624477805
transform 1 0 15194 0 1 -15284
box 70 126 186 240
use ptap  ptap_47
timestamp 1624477805
transform 1 0 16212 0 1 -15284
box 70 126 186 240
use ptap  ptap_48
timestamp 1624477805
transform 1 0 17230 0 1 -15284
box 70 126 186 240
use ptap  ptap_49
timestamp 1624477805
transform 1 0 18248 0 1 -15284
box 70 126 186 240
use ptap  ptap_50
timestamp 1624477805
transform 1 0 19266 0 1 -15284
box 70 126 186 240
use ptap  ptap_51
timestamp 1624477805
transform 1 0 20284 0 1 -15284
box 70 126 186 240
use ptap  ptap_52
timestamp 1624477805
transform 1 0 21302 0 1 -15284
box 70 126 186 240
use ptap  ptap_53
timestamp 1624477805
transform 1 0 22320 0 1 -15284
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_8
timestamp 1624477805
transform 1 0 12779 0 1 -14484
box -10209 -388 10209 388
use ptap  ptap_302
timestamp 1624477805
transform 1 0 -9294 0 1 -14222
box 70 126 186 240
use ptap  ptap_303
timestamp 1624477805
transform 1 0 -8276 0 1 -14222
box 70 126 186 240
use ptap  ptap_304
timestamp 1624477805
transform 1 0 -7258 0 1 -14222
box 70 126 186 240
use ptap  ptap_305
timestamp 1624477805
transform 1 0 -6240 0 1 -14222
box 70 126 186 240
use ptap  ptap_306
timestamp 1624477805
transform 1 0 -5222 0 1 -14222
box 70 126 186 240
use ptap  ptap_307
timestamp 1624477805
transform 1 0 -4204 0 1 -14222
box 70 126 186 240
use ptap  ptap_308
timestamp 1624477805
transform 1 0 -3186 0 1 -14222
box 70 126 186 240
use ptap  ptap_309
timestamp 1624477805
transform 1 0 -2168 0 1 -14222
box 70 126 186 240
use ptap  ptap_310
timestamp 1624477805
transform 1 0 -1150 0 1 -14222
box 70 126 186 240
use ptap  ptap_311
timestamp 1624477805
transform 1 0 -132 0 1 -14222
box 70 126 186 240
use ptap  ptap_0
timestamp 1624477805
transform 1 0 2966 0 1 -14050
box 70 126 186 240
use ptap  ptap_2
timestamp 1624477805
transform 1 0 5002 0 1 -14050
box 70 126 186 240
use ptap  ptap_1
timestamp 1624477805
transform 1 0 3984 0 1 -14050
box 70 126 186 240
use ptap  ptap_4
timestamp 1624477805
transform 1 0 7038 0 1 -14050
box 70 126 186 240
use ptap  ptap_3
timestamp 1624477805
transform 1 0 6020 0 1 -14050
box 70 126 186 240
use ptap  ptap_5
timestamp 1624477805
transform 1 0 8056 0 1 -14050
box 70 126 186 240
use ptap  ptap_7
timestamp 1624477805
transform 1 0 10092 0 1 -14050
box 70 126 186 240
use ptap  ptap_6
timestamp 1624477805
transform 1 0 9074 0 1 -14050
box 70 126 186 240
use ptap  ptap_9
timestamp 1624477805
transform 1 0 12128 0 1 -14050
box 70 126 186 240
use ptap  ptap_8
timestamp 1624477805
transform 1 0 11110 0 1 -14050
box 70 126 186 240
use ptap  ptap_10
timestamp 1624477805
transform 1 0 13146 0 1 -14050
box 70 126 186 240
use ptap  ptap_12
timestamp 1624477805
transform 1 0 15182 0 1 -14050
box 70 126 186 240
use ptap  ptap_11
timestamp 1624477805
transform 1 0 14164 0 1 -14050
box 70 126 186 240
use ptap  ptap_14
timestamp 1624477805
transform 1 0 17218 0 1 -14050
box 70 126 186 240
use ptap  ptap_13
timestamp 1624477805
transform 1 0 16200 0 1 -14050
box 70 126 186 240
use ptap  ptap_16
timestamp 1624477805
transform 1 0 19254 0 1 -14050
box 70 126 186 240
use ptap  ptap_15
timestamp 1624477805
transform 1 0 18236 0 1 -14050
box 70 126 186 240
use ptap  ptap_17
timestamp 1624477805
transform 1 0 20272 0 1 -14050
box 70 126 186 240
use ptap  ptap_19
timestamp 1624477805
transform 1 0 22308 0 1 -14050
box 70 126 186 240
use ptap  ptap_18
timestamp 1624477805
transform 1 0 21290 0 1 -14050
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_7
timestamp 1624477805
transform 1 0 12779 0 1 -13252
box -10209 -388 10209 388
use ptap  ptap_293
timestamp 1624477805
transform 1 0 -9294 0 1 -13404
box 70 126 186 240
use ptap  ptap_292
timestamp 1624477805
transform 1 0 -8276 0 1 -13404
box 70 126 186 240
use ptap  ptap_295
timestamp 1624477805
transform 1 0 -6240 0 1 -13404
box 70 126 186 240
use ptap  ptap_294
timestamp 1624477805
transform 1 0 -7258 0 1 -13404
box 70 126 186 240
use ptap  ptap_297
timestamp 1624477805
transform 1 0 -4204 0 1 -13404
box 70 126 186 240
use ptap  ptap_296
timestamp 1624477805
transform 1 0 -5222 0 1 -13404
box 70 126 186 240
use ptap  ptap_299
timestamp 1624477805
transform 1 0 -2168 0 1 -13404
box 70 126 186 240
use ptap  ptap_298
timestamp 1624477805
transform 1 0 -3186 0 1 -13404
box 70 126 186 240
use ptap  ptap_301
timestamp 1624477805
transform 1 0 -132 0 1 -13404
box 70 126 186 240
use ptap  ptap_300
timestamp 1624477805
transform 1 0 -1150 0 1 -13404
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_lvt_XH9Q8F  sky130_fd_pr__nfet_01v8_lvt_XH9Q8F_0
timestamp 1624477805
transform 1 0 -4586 0 1 -14039
box -4610 -1615 4610 1615
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_3
timestamp 1624477805
transform 1 0 -11932 0 1 -10618
box -350 -300 349 300
use sky130_fd_pr__cap_mim_m3_1_P3BUE2  sky130_fd_pr__cap_mim_m3_1_P3BUE2_7
timestamp 1624477805
transform 1 0 -10134 0 1 -10619
box -1150 -300 1149 300
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_15
timestamp 1624477805
transform 1 0 -10133 0 1 -8921
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_3 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/sample_and_hold
timestamp 1624477805
transform 1 0 -11930 0 1 -8920
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_P3BUE2  sky130_fd_pr__cap_mim_m3_1_P3BUE2_6
timestamp 1624477805
transform 1 0 -7534 0 1 -10619
box -1150 -300 1149 300
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_14
timestamp 1624477805
transform 1 0 -7533 0 1 -8921
box -1150 -1100 1149 1100
use ptap  ptap_291
timestamp 1624477805
transform 1 0 -8756 0 1 -12422
box 70 126 186 240
use sky130_fd_pr__cap_mim_m3_1_P3BUE2  sky130_fd_pr__cap_mim_m3_1_P3BUE2_5
timestamp 1624477805
transform 1 0 -4934 0 1 -10619
box -1150 -300 1149 300
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_13
timestamp 1624477805
transform 1 0 -4933 0 1 -8921
box -1150 -1100 1149 1100
use ptap  ptap_290
timestamp 1624477805
transform 1 0 -7738 0 1 -12422
box 70 126 186 240
use ptap  ptap_289
timestamp 1624477805
transform 1 0 -6720 0 1 -12422
box 70 126 186 240
use ptap  ptap_288
timestamp 1624477805
transform 1 0 -5702 0 1 -12422
box 70 126 186 240
use sky130_fd_pr__cap_mim_m3_1_P3BUE2  sky130_fd_pr__cap_mim_m3_1_P3BUE2_4
timestamp 1624477805
transform 1 0 -2334 0 1 -10619
box -1150 -300 1149 300
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_12
timestamp 1624477805
transform 1 0 -2333 0 1 -8921
box -1150 -1100 1149 1100
use ptap  ptap_287
timestamp 1624477805
transform 1 0 -4684 0 1 -12422
box 70 126 186 240
use ptap  ptap_286
timestamp 1624477805
transform 1 0 -3666 0 1 -12422
box 70 126 186 240
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_2
timestamp 1624477805
transform 1 0 -534 0 1 -10618
box -350 -300 349 300
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_4
timestamp 1624477805
transform 1 0 -536 0 1 -8920
box -350 -1100 349 1100
use ptap  ptap_285
timestamp 1624477805
transform 1 0 -2648 0 1 -12422
box 70 126 186 240
use ptap  ptap_284
timestamp 1624477805
transform 1 0 -1630 0 1 -12422
box 70 126 186 240
use ptap  ptap_283
timestamp 1624477805
transform 1 0 -612 0 1 -12422
box 70 126 186 240
use ptap  ptap_34
timestamp 1624477805
transform 1 0 2978 0 1 -12814
box 70 126 186 240
use ptap  ptap_35
timestamp 1624477805
transform 1 0 3996 0 1 -12814
box 70 126 186 240
use ptap  ptap_36
timestamp 1624477805
transform 1 0 5014 0 1 -12814
box 70 126 186 240
use ptap  ptap_37
timestamp 1624477805
transform 1 0 6032 0 1 -12814
box 70 126 186 240
use ptap  ptap_38
timestamp 1624477805
transform 1 0 7050 0 1 -12814
box 70 126 186 240
use ptap  ptap_39
timestamp 1624477805
transform 1 0 8068 0 1 -12814
box 70 126 186 240
use ptap  ptap_20
timestamp 1624477805
transform 1 0 9086 0 1 -12814
box 70 126 186 240
use ptap  ptap_21
timestamp 1624477805
transform 1 0 10104 0 1 -12814
box 70 126 186 240
use ptap  ptap_22
timestamp 1624477805
transform 1 0 11122 0 1 -12814
box 70 126 186 240
use ptap  ptap_23
timestamp 1624477805
transform 1 0 12140 0 1 -12814
box 70 126 186 240
use ptap  ptap_24
timestamp 1624477805
transform 1 0 13158 0 1 -12814
box 70 126 186 240
use ptap  ptap_25
timestamp 1624477805
transform 1 0 14176 0 1 -12814
box 70 126 186 240
use ptap  ptap_26
timestamp 1624477805
transform 1 0 15194 0 1 -12814
box 70 126 186 240
use ptap  ptap_27
timestamp 1624477805
transform 1 0 16212 0 1 -12814
box 70 126 186 240
use ptap  ptap_28
timestamp 1624477805
transform 1 0 17230 0 1 -12814
box 70 126 186 240
use ptap  ptap_29
timestamp 1624477805
transform 1 0 18248 0 1 -12814
box 70 126 186 240
use ptap  ptap_30
timestamp 1624477805
transform 1 0 19266 0 1 -12814
box 70 126 186 240
use ptap  ptap_31
timestamp 1624477805
transform 1 0 20284 0 1 -12814
box 70 126 186 240
use ptap  ptap_32
timestamp 1624477805
transform 1 0 21302 0 1 -12814
box 70 126 186 240
use ptap  ptap_33
timestamp 1624477805
transform 1 0 22320 0 1 -12814
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_6
timestamp 1624477805
transform 1 0 12779 0 1 -12018
box -10209 -388 10209 388
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_5
timestamp 1624477805
transform 1 0 -536 0 1 -6420
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_2
timestamp 1624477805
transform 1 0 -11930 0 1 -6420
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_10
timestamp 1624477805
transform 1 0 -7533 0 1 -6421
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_9
timestamp 1624477805
transform 1 0 -4933 0 1 -6421
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_8
timestamp 1624477805
transform 1 0 -2333 0 1 -6421
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_11
timestamp 1624477805
transform 1 0 -10133 0 1 -6421
box -1150 -1100 1149 1100
use sky130_fd_pr__pfet_01v8_LEMKJU  sky130_fd_pr__pfet_01v8_LEMKJU_3
timestamp 1624477805
transform 1 0 4733 0 1 -7704
box -1155 -300 1155 300
use sky130_fd_pr__pfet_01v8_MSJKJ2  sky130_fd_pr__pfet_01v8_MSJKJ2_3 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/se_fold_casc_wide_swing_ota
timestamp 1624477805
transform 1 0 15126 0 1 -7674
box -7700 -400 7700 400
use sky130_fd_pr__pfet_01v8_LEMKJU  sky130_fd_pr__pfet_01v8_LEMKJU_2
timestamp 1624477805
transform 1 0 4733 0 1 -6766
box -1155 -300 1155 300
use ntap  ntap_73 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/ntap
timestamp 1624477805
transform 1 0 9664 0 1 -7356
box 250 218 480 436
use ntap  ntap_72
timestamp 1624477805
transform 1 0 8646 0 1 -7356
box 250 218 480 436
use ntap  ntap_71
timestamp 1624477805
transform 1 0 7628 0 1 -7356
box 250 218 480 436
use ntap  ntap_100
timestamp 1624477805
transform 1 0 5362 0 1 -7550
box 250 218 480 436
use ntap  ntap_101
timestamp 1624477805
transform 1 0 4344 0 1 -7550
box 250 218 480 436
use ntap  ntap_102
timestamp 1624477805
transform 1 0 3326 0 1 -7550
box 250 218 480 436
use ntap  ntap_66
timestamp 1624477805
transform 1 0 17808 0 1 -7356
box 250 218 480 436
use ntap  ntap_65
timestamp 1624477805
transform 1 0 16790 0 1 -7356
box 250 218 480 436
use ntap  ntap_63
timestamp 1624477805
transform 1 0 14754 0 1 -7356
box 250 218 480 436
use ntap  ntap_64
timestamp 1624477805
transform 1 0 15772 0 1 -7356
box 250 218 480 436
use ntap  ntap_62
timestamp 1624477805
transform 1 0 13736 0 1 -7356
box 250 218 480 436
use ntap  ntap_61
timestamp 1624477805
transform 1 0 12718 0 1 -7356
box 250 218 480 436
use ntap  ntap_74
timestamp 1624477805
transform 1 0 10682 0 1 -7356
box 250 218 480 436
use ntap  ntap_75
timestamp 1624477805
transform 1 0 11700 0 1 -7356
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_MSJKJ2  sky130_fd_pr__pfet_01v8_MSJKJ2_2
timestamp 1624477805
transform 1 0 15126 0 1 -6418
box -7700 -400 7700 400
use ntap  ntap_70
timestamp 1624477805
transform 1 0 21880 0 1 -7356
box 250 218 480 436
use ntap  ntap_69
timestamp 1624477805
transform 1 0 20862 0 1 -7356
box 250 218 480 436
use ntap  ntap_67
timestamp 1624477805
transform 1 0 18826 0 1 -7356
box 250 218 480 436
use ntap  ntap_68
timestamp 1624477805
transform 1 0 19844 0 1 -7356
box 250 218 480 436
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_6
timestamp 1624477805
transform 1 0 -536 0 1 -3920
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_1
timestamp 1624477805
transform 1 0 -11930 0 1 -3920
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_6
timestamp 1624477805
transform 1 0 -7533 0 1 -3921
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_5
timestamp 1624477805
transform 1 0 -4933 0 1 -3921
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_4
timestamp 1624477805
transform 1 0 -2333 0 1 -3921
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_7
timestamp 1624477805
transform 1 0 -10133 0 1 -3921
box -1150 -1100 1149 1100
use sky130_fd_pr__pfet_01v8_LEMKJU  sky130_fd_pr__pfet_01v8_LEMKJU_1
timestamp 1624477805
transform 1 0 4733 0 1 -5828
box -1155 -300 1155 300
use ntap  ntap_98
timestamp 1624477805
transform 1 0 4344 0 1 -6636
box 250 218 480 436
use ntap  ntap_99
timestamp 1624477805
transform 1 0 3326 0 1 -6636
box 250 218 480 436
use ntap  ntap_97
timestamp 1624477805
transform 1 0 5362 0 1 -6636
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_LEMKJU  sky130_fd_pr__pfet_01v8_LEMKJU_0
timestamp 1624477805
transform 1 0 4733 0 1 -4890
box -1155 -300 1155 300
use ntap  ntap_94
timestamp 1624477805
transform 1 0 5390 0 1 -5694
box 250 218 480 436
use ntap  ntap_95
timestamp 1624477805
transform 1 0 4372 0 1 -5694
box 250 218 480 436
use ntap  ntap_96
timestamp 1624477805
transform 1 0 3354 0 1 -5694
box 250 218 480 436
use ntap  ntap_56
timestamp 1624477805
transform 1 0 7628 0 1 -6118
box 250 218 480 436
use ntap  ntap_57
timestamp 1624477805
transform 1 0 8646 0 1 -6118
box 250 218 480 436
use ntap  ntap_58
timestamp 1624477805
transform 1 0 9664 0 1 -6118
box 250 218 480 436
use ntap  ntap_51
timestamp 1624477805
transform 1 0 17808 0 1 -6118
box 250 218 480 436
use ntap  ntap_50
timestamp 1624477805
transform 1 0 16790 0 1 -6118
box 250 218 480 436
use ntap  ntap_49
timestamp 1624477805
transform 1 0 15772 0 1 -6118
box 250 218 480 436
use ntap  ntap_48
timestamp 1624477805
transform 1 0 14754 0 1 -6118
box 250 218 480 436
use ntap  ntap_47
timestamp 1624477805
transform 1 0 13736 0 1 -6118
box 250 218 480 436
use ntap  ntap_46
timestamp 1624477805
transform 1 0 12718 0 1 -6118
box 250 218 480 436
use ntap  ntap_60
timestamp 1624477805
transform 1 0 11700 0 1 -6118
box 250 218 480 436
use ntap  ntap_59
timestamp 1624477805
transform 1 0 10682 0 1 -6118
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_MSJKJ2  sky130_fd_pr__pfet_01v8_MSJKJ2_0
timestamp 1624477805
transform 1 0 15126 0 1 -5162
box -7700 -400 7700 400
use ntap  ntap_93
timestamp 1624477805
transform 1 0 3396 0 1 -4610
box 250 218 480 436
use ntap  ntap_92
timestamp 1624477805
transform 1 0 4414 0 1 -4610
box 250 218 480 436
use ntap  ntap_91
timestamp 1624477805
transform 1 0 5432 0 1 -4610
box 250 218 480 436
use ntap  ntap_31
timestamp 1624477805
transform 1 0 7670 0 1 -4850
box 250 218 480 436
use ntap  ntap_32
timestamp 1624477805
transform 1 0 8688 0 1 -4850
box 250 218 480 436
use ntap  ntap_33
timestamp 1624477805
transform 1 0 9706 0 1 -4850
box 250 218 480 436
use ntap  ntap_34
timestamp 1624477805
transform 1 0 10724 0 1 -4850
box 250 218 480 436
use ntap  ntap_36
timestamp 1624477805
transform 1 0 12760 0 1 -4850
box 250 218 480 436
use ntap  ntap_35
timestamp 1624477805
transform 1 0 11742 0 1 -4850
box 250 218 480 436
use ntap  ntap_37
timestamp 1624477805
transform 1 0 13778 0 1 -4850
box 250 218 480 436
use ntap  ntap_38
timestamp 1624477805
transform 1 0 14796 0 1 -4850
box 250 218 480 436
use ntap  ntap_39
timestamp 1624477805
transform 1 0 15814 0 1 -4850
box 250 218 480 436
use ntap  ntap_40
timestamp 1624477805
transform 1 0 16832 0 1 -4850
box 250 218 480 436
use ntap  ntap_41
timestamp 1624477805
transform 1 0 17850 0 1 -4850
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_MSJKJ2  sky130_fd_pr__pfet_01v8_MSJKJ2_1
timestamp 1624477805
transform 1 0 15126 0 1 -3906
box -7700 -400 7700 400
use ntap  ntap_45
timestamp 1624477805
transform 1 0 21922 0 1 -4850
box 250 218 480 436
use ntap  ntap_44
timestamp 1624477805
transform 1 0 20904 0 1 -4850
box 250 218 480 436
use ntap  ntap_42
timestamp 1624477805
transform 1 0 18868 0 1 -4850
box 250 218 480 436
use ntap  ntap_43
timestamp 1624477805
transform 1 0 19886 0 1 -4850
box 250 218 480 436
use ntap  ntap_55
timestamp 1624477805
transform 1 0 21880 0 1 -6118
box 250 218 480 436
use ntap  ntap_54
timestamp 1624477805
transform 1 0 20862 0 1 -6118
box 250 218 480 436
use ntap  ntap_52
timestamp 1624477805
transform 1 0 18826 0 1 -6118
box 250 218 480 436
use ntap  ntap_53
timestamp 1624477805
transform 1 0 19844 0 1 -6118
box 250 218 480 436
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_7
timestamp 1624477805
transform 1 0 -536 0 1 -1420
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_0
timestamp 1624477805
transform 1 0 -11930 0 1 -1420
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_1
timestamp 1624477805
transform 1 0 -7533 0 1 -1420
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_2
timestamp 1624477805
transform 1 0 -4933 0 1 -1420
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_3
timestamp 1624477805
transform 1 0 -2333 0 1 -1420
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_0
timestamp 1624477805
transform 1 0 -10133 0 1 -1420
box -1150 -1100 1149 1100
use ntap  ntap_30
timestamp 1624477805
transform 1 0 7670 0 1 -3338
box 250 218 480 436
use ntap  ntap_29
timestamp 1624477805
transform 1 0 8688 0 1 -3338
box 250 218 480 436
use ntap  ntap_28
timestamp 1624477805
transform 1 0 9706 0 1 -3338
box 250 218 480 436
use ntap  ntap_27
timestamp 1624477805
transform 1 0 10724 0 1 -3338
box 250 218 480 436
use ntap  ntap_26
timestamp 1624477805
transform 1 0 11742 0 1 -3338
box 250 218 480 436
use ntap  ntap_24
timestamp 1624477805
transform 1 0 13778 0 1 -3338
box 250 218 480 436
use ntap  ntap_25
timestamp 1624477805
transform 1 0 12760 0 1 -3338
box 250 218 480 436
use ntap  ntap_23
timestamp 1624477805
transform 1 0 14796 0 1 -3338
box 250 218 480 436
use ntap  ntap_22
timestamp 1624477805
transform 1 0 15814 0 1 -3338
box 250 218 480 436
use ntap  ntap_21
timestamp 1624477805
transform 1 0 16832 0 1 -3338
box 250 218 480 436
use ntap  ntap_19
timestamp 1624477805
transform 1 0 18868 0 1 -3338
box 250 218 480 436
use ntap  ntap_20
timestamp 1624477805
transform 1 0 17850 0 1 -3338
box 250 218 480 436
use ntap  ntap_18
timestamp 1624477805
transform 1 0 19886 0 1 -3338
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_V2JKJ2  sky130_fd_pr__pfet_01v8_lvt_V2JKJ2_2 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/se_fold_casc_wide_swing_ota
timestamp 1624477805
transform 1 0 14649 0 1 -2132
box -8209 -400 8209 400
use ntap  ntap_0
timestamp 1624477805
transform 1 0 6652 0 1 -1894
box 250 218 480 436
use ntap  ntap_1
timestamp 1624477805
transform 1 0 7670 0 1 -1894
box 250 218 480 436
use ntap  ntap_3
timestamp 1624477805
transform 1 0 9706 0 1 -1894
box 250 218 480 436
use ntap  ntap_2
timestamp 1624477805
transform 1 0 8688 0 1 -1894
box 250 218 480 436
use ntap  ntap_4
timestamp 1624477805
transform 1 0 10724 0 1 -1894
box 250 218 480 436
use ntap  ntap_5
timestamp 1624477805
transform 1 0 11742 0 1 -1894
box 250 218 480 436
use ntap  ntap_6
timestamp 1624477805
transform 1 0 12760 0 1 -1894
box 250 218 480 436
use ntap  ntap_7
timestamp 1624477805
transform 1 0 13778 0 1 -1894
box 250 218 480 436
use ntap  ntap_8
timestamp 1624477805
transform 1 0 14796 0 1 -1894
box 250 218 480 436
use ntap  ntap_9
timestamp 1624477805
transform 1 0 15814 0 1 -1894
box 250 218 480 436
use ntap  ntap_10
timestamp 1624477805
transform 1 0 16832 0 1 -1894
box 250 218 480 436
use ntap  ntap_11
timestamp 1624477805
transform 1 0 17850 0 1 -1894
box 250 218 480 436
use ntap  ntap_12
timestamp 1624477805
transform 1 0 18868 0 1 -1894
box 250 218 480 436
use ntap  ntap_13
timestamp 1624477805
transform 1 0 19886 0 1 -1894
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_V2JKJ2  sky130_fd_pr__pfet_01v8_lvt_V2JKJ2_1
timestamp 1624477805
transform 1 0 14649 0 1 -996
box -8209 -400 8209 400
use ntap  ntap_86
timestamp 1624477805
transform 1 0 7670 0 1 -742
box 250 218 480 436
use ntap  ntap_87
timestamp 1624477805
transform 1 0 8688 0 1 -742
box 250 218 480 436
use ntap  ntap_88
timestamp 1624477805
transform 1 0 9706 0 1 -742
box 250 218 480 436
use ntap  ntap_89
timestamp 1624477805
transform 1 0 10724 0 1 -742
box 250 218 480 436
use ntap  ntap_90
timestamp 1624477805
transform 1 0 11742 0 1 -742
box 250 218 480 436
use ntap  ntap_77
timestamp 1624477805
transform 1 0 13778 0 1 -742
box 250 218 480 436
use ntap  ntap_76
timestamp 1624477805
transform 1 0 12760 0 1 -742
box 250 218 480 436
use ntap  ntap_78
timestamp 1624477805
transform 1 0 14796 0 1 -742
box 250 218 480 436
use ntap  ntap_79
timestamp 1624477805
transform 1 0 15814 0 1 -742
box 250 218 480 436
use ntap  ntap_80
timestamp 1624477805
transform 1 0 16832 0 1 -742
box 250 218 480 436
use ntap  ntap_82
timestamp 1624477805
transform 1 0 18868 0 1 -742
box 250 218 480 436
use ntap  ntap_81
timestamp 1624477805
transform 1 0 17850 0 1 -742
box 250 218 480 436
use ntap  ntap_83
timestamp 1624477805
transform 1 0 19886 0 1 -742
box 250 218 480 436
use ntap  ntap_84
timestamp 1624477805
transform 1 0 20904 0 1 -742
box 250 218 480 436
use ntap  ntap_85
timestamp 1624477805
transform 1 0 21922 0 1 -742
box 250 218 480 436
use ntap  ntap_15
timestamp 1624477805
transform 1 0 21922 0 1 -1894
box 250 218 480 436
use ntap  ntap_16
timestamp 1624477805
transform 1 0 21922 0 1 -3338
box 250 218 480 436
use ntap  ntap_14
timestamp 1624477805
transform 1 0 20904 0 1 -1894
box 250 218 480 436
use ntap  ntap_17
timestamp 1624477805
transform 1 0 20904 0 1 -3338
box 250 218 480 436
use sky130_fd_pr__cap_mim_m3_1_P3BUE2  sky130_fd_pr__cap_mim_m3_1_P3BUE2_0
timestamp 1624477805
transform 1 0 -10134 0 1 281
box -1150 -300 1149 300
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_0
timestamp 1624477805
transform 1 0 -11928 0 1 280
box -350 -300 349 300
use sky130_fd_pr__cap_mim_m3_1_P3BUE2  sky130_fd_pr__cap_mim_m3_1_P3BUE2_2
timestamp 1624477805
transform 1 0 -4934 0 1 281
box -1150 -300 1149 300
use sky130_fd_pr__cap_mim_m3_1_P3BUE2  sky130_fd_pr__cap_mim_m3_1_P3BUE2_1
timestamp 1624477805
transform 1 0 -7534 0 1 281
box -1150 -300 1149 300
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_1
timestamp 1624477805
transform 1 0 -534 0 1 280
box -350 -300 349 300
use sky130_fd_pr__cap_mim_m3_1_P3BUE2  sky130_fd_pr__cap_mim_m3_1_P3BUE2_3
timestamp 1624477805
transform 1 0 -2334 0 1 281
box -1150 -300 1149 300
use sky130_fd_pr__pfet_01v8_lvt_V2JKJ2  sky130_fd_pr__pfet_01v8_lvt_V2JKJ2_0
timestamp 1624477805
transform 1 0 14649 0 1 140
box -8209 -400 8209 400
<< labels >>
flabel metal2 9924 -2710 9924 -2710 1 FreeSans 480 0 0 0 vfoldm
flabel metal1 6356 -500 6356 -500 1 FreeSans 480 0 0 0 M1d
flabel metal1 7520 -2684 7520 -2684 1 FreeSans 480 0 0 0 M2d
flabel metal2 7798 -524 7798 -524 1 FreeSans 480 0 0 0 M6d
flabel metal1 7340 -3616 7340 -3616 1 FreeSans 480 0 0 0 M1d
flabel metal2 7618 -4582 7618 -4582 1 FreeSans 480 0 0 0 vbias1
flabel metal2 7514 -8154 7514 -8154 1 FreeSans 480 0 0 0 M2d
flabel metal2 16472 -5648 16472 -5648 1 FreeSans 480 0 0 0 M6d
flabel metal1 16668 -6000 16668 -6000 1 FreeSans 480 0 0 0 M13d
flabel metal2 11872 -8432 11872 -8432 1 FreeSans 480 0 0 0 M3d
flabel metal1 20726 -5618 20726 -5618 1 FreeSans 480 0 0 0 vfoldm
flabel metal2 20598 -6894 20598 -6894 1 FreeSans 480 0 0 0 vfoldp
flabel metal2 11830 716 11830 716 1 FreeSans 480 0 0 0 vfoldp
flabel metal2 3964 -6186 3964 -6186 1 FreeSans 480 0 0 0 vcmc_casc
flabel metal2 5800 -7134 5800 -7134 1 FreeSans 480 0 0 0 vcmcn_casc
flabel metal1 6080 -7670 6080 -7670 1 FreeSans 480 0 0 0 vcmcn2_casc
flabel metal1 3524 -7256 3524 -7256 1 FreeSans 480 0 0 0 vcmcn1_casc
flabel metal2 8324 850 8324 850 1 FreeSans 480 0 0 0 vbias1
flabel metal2 22386 -5742 22418 -5726 1 FreeSans 480 0 0 0 vom
port 16 n
flabel metal1 22574 -6900 22616 -6878 1 FreeSans 480 0 0 0 vop
port 17 n
flabel metal2 9302 588 9332 616 1 FreeSans 480 0 0 0 VDD
flabel metal2 -2498 -19392 -2424 -19358 1 FreeSans 480 0 0 0 vocm
port 15 n
flabel metal1 -6348 -21586 -6316 -21566 1 FreeSans 480 0 0 0 ibiasn
port 14 n
flabel metal1 2248 -17074 2270 -17046 1 FreeSans 480 0 0 0 vom
flabel metal2 12404 -15160 12436 -15142 1 FreeSans 480 0 0 0 vop
flabel metal1 23180 -18038 23204 -18008 1 FreeSans 480 0 0 0 VSS
flabel metal1 -5330 -24996 -5294 -24960 1 FreeSans 480 0 0 0 VSS
port 13 n
flabel metal1 23556 -17190 23556 -17190 1 FreeSans 480 0 0 0 vbias3
flabel metal1 2144 -12732 2144 -12732 1 FreeSans 480 0 0 0 vcmc_casc
flabel metal1 -2940 -20628 -2940 -20628 1 FreeSans 480 0 0 0 vcmn_casc_tail2
flabel metal2 -3068 -20216 -3068 -20216 1 FreeSans 480 0 0 0 vcmn_casc_tail1
flabel metal1 132 -19622 132 -19622 1 FreeSans 480 0 0 0 vcmcn2_casc
flabel metal1 -338 -20144 -338 -20144 1 FreeSans 480 0 0 0 vcmcn_casc
flabel metal1 18 -19488 18 -19488 1 FreeSans 480 0 0 0 vcmcn1_casc
flabel metal2 -1114 -21516 -1114 -21516 1 FreeSans 480 0 0 0 vfoldp
flabel metal1 -2656 -23502 -2622 -23470 1 FreeSans 480 0 0 0 vip
port 10 n
flabel metal1 1096 -23294 1122 -23264 1 FreeSans 480 0 0 0 vim
port 9 n
flabel metal1 4648 -16436 4648 -16436 1 FreeSans 480 0 0 0 vcascnp
flabel metal1 23300 -16984 23300 -16984 1 FreeSans 480 0 0 0 vcascnm
flabel metal1 23436 -21216 23436 -21216 1 FreeSans 480 0 0 0 vbias4
flabel metal1 2006 -14484 2006 -14484 1 FreeSans 480 0 0 0 vtail_casc
flabel metal1 23678 -12818 23678 -12814 1 FreeSans 480 0 0 0 M3d
flabel metal1 22954 -15336 22954 -15336 1 FreeSans 480 0 0 0 M13d
flabel metal1 592 -22748 592 -22748 1 FreeSans 480 0 0 0 vtail_casc
flabel metal1 -2092 -23816 -2092 -23816 1 FreeSans 480 0 0 0 vfoldm
flabel metal1 -9506 -22906 -9506 -22906 1 FreeSans 480 0 0 0 vcmn_casc_tail2
flabel metal1 -8364 -23636 -8364 -23636 1 FreeSans 480 0 0 0 vbias2
flabel metal1 -4292 -23864 -4292 -23864 1 FreeSans 480 0 0 0 vcmn_casc_tail1
flabel metal1 -8078 -12352 -8078 -12352 1 FreeSans 480 0 0 0 vbias1
flabel metal1 -6206 -19026 -6206 -19026 1 FreeSans 480 0 0 0 vbias2
flabel metal4 -1342 -5198 -1266 -5156 1 FreeSans 480 0 0 0 vom
flabel metal4 -10820 -2704 -10756 -2664 1 FreeSans 480 0 0 0 vop
flabel metal1 -2450 -19926 -2422 -19890 1 FreeSans 480 0 0 0 vom
flabel metal2 -768 -19990 -736 -19968 1 FreeSans 480 0 0 0 vop
flabel metal1 17510 -4394 17546 -4366 1 FreeSans 480 0 0 0 VDD
flabel metal4 -12400 1000 -12400 1800 3 FreeSans 3200 0 0 0 VDD
port 18 e
flabel metal4 -12400 -27200 -12400 -26400 3 FreeSans 3200 0 0 0 VSS
<< properties >>
string FIXED_BBOX -10872 -26372 24872 -10428
<< end >>
