magic
tech sky130A
magscale 1 2
timestamp 1623981089
<< nwell >>
rect -2622 123 3321 444
rect -2454 122 3321 123
rect -2622 -966 3320 -398
rect -2622 -2054 3320 -1486
rect -2622 -2896 3320 -2574
<< pwell >>
rect -2582 -342 3280 66
rect -2582 -1430 3280 -1022
rect -2582 -2518 3280 -2110
<< scnmos >>
rect -2163 -91 -2133 -7
rect -2079 -91 -2049 -7
rect -1891 -91 -1861 -7
rect -1779 -91 -1749 -19
rect -1680 -91 -1650 -19
rect -1581 -91 -1551 -7
rect -1462 -91 -1432 37
rect -1361 -91 -1331 -19
rect -1255 -91 -1225 -19
rect -1160 -91 -1130 -7
rect -970 -91 -940 39
rect -886 -91 -856 39
rect -698 -91 -668 -7
rect -603 -91 -573 39
rect -374 -91 -344 39
rect -129 -91 -99 39
rect -45 -91 -15 39
rect 39 -91 69 39
rect 123 -91 153 39
rect -2163 -269 -2133 -185
rect -2079 -269 -2049 -185
rect -1891 -269 -1861 -185
rect -1779 -257 -1749 -185
rect -1680 -257 -1650 -185
rect -1581 -269 -1551 -185
rect -1462 -313 -1432 -185
rect -1361 -257 -1331 -185
rect -1255 -257 -1225 -185
rect -1160 -269 -1130 -185
rect -970 -315 -940 -185
rect -886 -315 -856 -185
rect -698 -269 -668 -185
rect -603 -315 -573 -185
rect -374 -315 -344 -185
rect -129 -315 -99 -185
rect -45 -315 -15 -185
rect 39 -315 69 -185
rect 123 -315 153 -185
rect 535 -269 565 -185
rect 619 -269 649 -185
rect 807 -269 837 -185
rect 919 -257 949 -185
rect 1018 -257 1048 -185
rect 1117 -269 1147 -185
rect 1236 -313 1266 -185
rect 1337 -257 1367 -185
rect 1443 -257 1473 -185
rect 1538 -269 1568 -185
rect 1728 -315 1758 -185
rect 1812 -315 1842 -185
rect 2000 -269 2030 -185
rect 2095 -315 2125 -185
rect 2324 -315 2354 -185
rect 2569 -315 2599 -185
rect 2653 -315 2683 -185
rect 2737 -315 2767 -185
rect 2821 -315 2851 -185
rect -2163 -1179 -2133 -1095
rect -2079 -1179 -2049 -1095
rect -1891 -1179 -1861 -1095
rect -1779 -1179 -1749 -1107
rect -1680 -1179 -1650 -1107
rect -1581 -1179 -1551 -1095
rect -1462 -1179 -1432 -1051
rect -1361 -1179 -1331 -1107
rect -1255 -1179 -1225 -1107
rect -1160 -1179 -1130 -1095
rect -970 -1179 -940 -1049
rect -886 -1179 -856 -1049
rect -698 -1179 -668 -1095
rect -603 -1179 -573 -1049
rect -374 -1179 -344 -1049
rect -129 -1179 -99 -1049
rect -45 -1179 -15 -1049
rect 39 -1179 69 -1049
rect 123 -1179 153 -1049
rect 535 -1179 565 -1095
rect 619 -1179 649 -1095
rect 807 -1179 837 -1095
rect 919 -1179 949 -1107
rect 1018 -1179 1048 -1107
rect 1117 -1179 1147 -1095
rect 1236 -1179 1266 -1051
rect 1337 -1179 1367 -1107
rect 1443 -1179 1473 -1107
rect 1538 -1179 1568 -1095
rect 1728 -1179 1758 -1049
rect 1812 -1179 1842 -1049
rect 2000 -1179 2030 -1095
rect 2095 -1179 2125 -1049
rect 2324 -1179 2354 -1049
rect 2569 -1179 2599 -1049
rect 2653 -1179 2683 -1049
rect 2737 -1179 2767 -1049
rect 2821 -1179 2851 -1049
rect -2163 -1357 -2133 -1273
rect -2079 -1357 -2049 -1273
rect -1891 -1357 -1861 -1273
rect -1779 -1345 -1749 -1273
rect -1680 -1345 -1650 -1273
rect -1581 -1357 -1551 -1273
rect -1462 -1401 -1432 -1273
rect -1361 -1345 -1331 -1273
rect -1255 -1345 -1225 -1273
rect -1160 -1357 -1130 -1273
rect -970 -1403 -940 -1273
rect -886 -1403 -856 -1273
rect -698 -1357 -668 -1273
rect -603 -1403 -573 -1273
rect -374 -1403 -344 -1273
rect -129 -1403 -99 -1273
rect -45 -1403 -15 -1273
rect 39 -1403 69 -1273
rect 123 -1403 153 -1273
rect 535 -1357 565 -1273
rect 619 -1357 649 -1273
rect 807 -1357 837 -1273
rect 919 -1345 949 -1273
rect 1018 -1345 1048 -1273
rect 1117 -1357 1147 -1273
rect 1236 -1401 1266 -1273
rect 1337 -1345 1367 -1273
rect 1443 -1345 1473 -1273
rect 1538 -1357 1568 -1273
rect 1728 -1403 1758 -1273
rect 1812 -1403 1842 -1273
rect 2000 -1357 2030 -1273
rect 2095 -1403 2125 -1273
rect 2324 -1403 2354 -1273
rect 2569 -1403 2599 -1273
rect 2653 -1403 2683 -1273
rect 2737 -1403 2767 -1273
rect 2821 -1403 2851 -1273
rect -2163 -2267 -2133 -2183
rect -2079 -2267 -2049 -2183
rect -1891 -2267 -1861 -2183
rect -1779 -2267 -1749 -2195
rect -1680 -2267 -1650 -2195
rect -1581 -2267 -1551 -2183
rect -1462 -2267 -1432 -2139
rect -1361 -2267 -1331 -2195
rect -1255 -2267 -1225 -2195
rect -1160 -2267 -1130 -2183
rect -970 -2267 -940 -2137
rect -886 -2267 -856 -2137
rect -698 -2267 -668 -2183
rect -603 -2267 -573 -2137
rect -374 -2267 -344 -2137
rect -129 -2267 -99 -2137
rect -45 -2267 -15 -2137
rect 39 -2267 69 -2137
rect 123 -2267 153 -2137
rect 535 -2267 565 -2183
rect 619 -2267 649 -2183
rect 807 -2267 837 -2183
rect 919 -2267 949 -2195
rect 1018 -2267 1048 -2195
rect 1117 -2267 1147 -2183
rect 1236 -2267 1266 -2139
rect 1337 -2267 1367 -2195
rect 1443 -2267 1473 -2195
rect 1538 -2267 1568 -2183
rect 1728 -2267 1758 -2137
rect 1812 -2267 1842 -2137
rect 2000 -2267 2030 -2183
rect 2095 -2267 2125 -2137
rect 2324 -2267 2354 -2137
rect 2569 -2267 2599 -2137
rect 2653 -2267 2683 -2137
rect 2737 -2267 2767 -2137
rect 2821 -2267 2851 -2137
rect -2163 -2445 -2133 -2361
rect -2079 -2445 -2049 -2361
rect -1891 -2445 -1861 -2361
rect -1779 -2433 -1749 -2361
rect -1680 -2433 -1650 -2361
rect -1581 -2445 -1551 -2361
rect -1462 -2489 -1432 -2361
rect -1361 -2433 -1331 -2361
rect -1255 -2433 -1225 -2361
rect -1160 -2445 -1130 -2361
rect -970 -2491 -940 -2361
rect -886 -2491 -856 -2361
rect -698 -2445 -668 -2361
rect -603 -2491 -573 -2361
rect -374 -2491 -344 -2361
rect -129 -2491 -99 -2361
rect -45 -2491 -15 -2361
rect 39 -2491 69 -2361
rect 123 -2491 153 -2361
rect 535 -2445 565 -2361
rect 619 -2445 649 -2361
rect 807 -2445 837 -2361
rect 919 -2433 949 -2361
rect 1018 -2433 1048 -2361
rect 1117 -2445 1147 -2361
rect 1236 -2489 1266 -2361
rect 1337 -2433 1367 -2361
rect 1443 -2433 1473 -2361
rect 1538 -2445 1568 -2361
rect 1728 -2491 1758 -2361
rect 1812 -2491 1842 -2361
rect 2000 -2445 2030 -2361
rect 2095 -2491 2125 -2361
rect 2324 -2491 2354 -2361
rect 2569 -2491 2599 -2361
rect 2653 -2491 2683 -2361
rect 2737 -2491 2767 -2361
rect 2821 -2491 2851 -2361
<< scpmoshvt >>
rect -2163 225 -2133 353
rect -2079 225 -2049 353
rect -1891 275 -1861 359
rect -1806 275 -1776 359
rect -1711 275 -1681 359
rect -1608 275 -1578 359
rect -1476 209 -1446 359
rect -1381 275 -1351 359
rect -1297 275 -1267 359
rect -1183 275 -1153 359
rect -972 159 -942 359
rect -888 159 -858 359
rect -700 231 -670 359
rect -603 159 -573 359
rect -374 159 -344 359
rect -129 159 -99 359
rect -45 159 -15 359
rect 39 159 69 359
rect 123 159 153 359
rect -2163 -629 -2133 -501
rect -2079 -629 -2049 -501
rect -1891 -635 -1861 -551
rect -1806 -635 -1776 -551
rect -1711 -635 -1681 -551
rect -1608 -635 -1578 -551
rect -1476 -635 -1446 -485
rect -1381 -635 -1351 -551
rect -1297 -635 -1267 -551
rect -1183 -635 -1153 -551
rect -972 -635 -942 -435
rect -888 -635 -858 -435
rect -700 -635 -670 -507
rect -603 -635 -573 -435
rect -374 -635 -344 -435
rect -129 -635 -99 -435
rect -45 -635 -15 -435
rect 39 -635 69 -435
rect 123 -635 153 -435
rect 535 -629 565 -501
rect 619 -629 649 -501
rect 807 -635 837 -551
rect 892 -635 922 -551
rect 987 -635 1017 -551
rect 1090 -635 1120 -551
rect 1222 -635 1252 -485
rect 1317 -635 1347 -551
rect 1401 -635 1431 -551
rect 1515 -635 1545 -551
rect 1726 -635 1756 -435
rect 1810 -635 1840 -435
rect 1998 -635 2028 -507
rect 2095 -635 2125 -435
rect 2324 -635 2354 -435
rect 2569 -635 2599 -435
rect 2653 -635 2683 -435
rect 2737 -635 2767 -435
rect 2821 -635 2851 -435
rect -2163 -863 -2133 -735
rect -2079 -863 -2049 -735
rect -1891 -813 -1861 -729
rect -1806 -813 -1776 -729
rect -1711 -813 -1681 -729
rect -1608 -813 -1578 -729
rect -1476 -879 -1446 -729
rect -1381 -813 -1351 -729
rect -1297 -813 -1267 -729
rect -1183 -813 -1153 -729
rect -972 -929 -942 -729
rect -888 -929 -858 -729
rect -700 -857 -670 -729
rect -603 -929 -573 -729
rect -374 -929 -344 -729
rect -129 -929 -99 -729
rect -45 -929 -15 -729
rect 39 -929 69 -729
rect 123 -929 153 -729
rect 535 -863 565 -735
rect 619 -863 649 -735
rect 807 -813 837 -729
rect 892 -813 922 -729
rect 987 -813 1017 -729
rect 1090 -813 1120 -729
rect 1222 -879 1252 -729
rect 1317 -813 1347 -729
rect 1401 -813 1431 -729
rect 1515 -813 1545 -729
rect 1726 -929 1756 -729
rect 1810 -929 1840 -729
rect 1998 -857 2028 -729
rect 2095 -929 2125 -729
rect 2324 -929 2354 -729
rect 2569 -929 2599 -729
rect 2653 -929 2683 -729
rect 2737 -929 2767 -729
rect 2821 -929 2851 -729
rect -2163 -1717 -2133 -1589
rect -2079 -1717 -2049 -1589
rect -1891 -1723 -1861 -1639
rect -1806 -1723 -1776 -1639
rect -1711 -1723 -1681 -1639
rect -1608 -1723 -1578 -1639
rect -1476 -1723 -1446 -1573
rect -1381 -1723 -1351 -1639
rect -1297 -1723 -1267 -1639
rect -1183 -1723 -1153 -1639
rect -972 -1723 -942 -1523
rect -888 -1723 -858 -1523
rect -700 -1723 -670 -1595
rect -603 -1723 -573 -1523
rect -374 -1723 -344 -1523
rect -129 -1723 -99 -1523
rect -45 -1723 -15 -1523
rect 39 -1723 69 -1523
rect 123 -1723 153 -1523
rect 535 -1717 565 -1589
rect 619 -1717 649 -1589
rect 807 -1723 837 -1639
rect 892 -1723 922 -1639
rect 987 -1723 1017 -1639
rect 1090 -1723 1120 -1639
rect 1222 -1723 1252 -1573
rect 1317 -1723 1347 -1639
rect 1401 -1723 1431 -1639
rect 1515 -1723 1545 -1639
rect 1726 -1723 1756 -1523
rect 1810 -1723 1840 -1523
rect 1998 -1723 2028 -1595
rect 2095 -1723 2125 -1523
rect 2324 -1723 2354 -1523
rect 2569 -1723 2599 -1523
rect 2653 -1723 2683 -1523
rect 2737 -1723 2767 -1523
rect 2821 -1723 2851 -1523
rect -2163 -1951 -2133 -1823
rect -2079 -1951 -2049 -1823
rect -1891 -1901 -1861 -1817
rect -1806 -1901 -1776 -1817
rect -1711 -1901 -1681 -1817
rect -1608 -1901 -1578 -1817
rect -1476 -1967 -1446 -1817
rect -1381 -1901 -1351 -1817
rect -1297 -1901 -1267 -1817
rect -1183 -1901 -1153 -1817
rect -972 -2017 -942 -1817
rect -888 -2017 -858 -1817
rect -700 -1945 -670 -1817
rect -603 -2017 -573 -1817
rect -374 -2017 -344 -1817
rect -129 -2017 -99 -1817
rect -45 -2017 -15 -1817
rect 39 -2017 69 -1817
rect 123 -2017 153 -1817
rect 535 -1951 565 -1823
rect 619 -1951 649 -1823
rect 807 -1901 837 -1817
rect 892 -1901 922 -1817
rect 987 -1901 1017 -1817
rect 1090 -1901 1120 -1817
rect 1222 -1967 1252 -1817
rect 1317 -1901 1347 -1817
rect 1401 -1901 1431 -1817
rect 1515 -1901 1545 -1817
rect 1726 -2017 1756 -1817
rect 1810 -2017 1840 -1817
rect 1998 -1945 2028 -1817
rect 2095 -2017 2125 -1817
rect 2324 -2017 2354 -1817
rect 2569 -2017 2599 -1817
rect 2653 -2017 2683 -1817
rect 2737 -2017 2767 -1817
rect 2821 -2017 2851 -1817
rect -2163 -2805 -2133 -2677
rect -2079 -2805 -2049 -2677
rect -1891 -2811 -1861 -2727
rect -1806 -2811 -1776 -2727
rect -1711 -2811 -1681 -2727
rect -1608 -2811 -1578 -2727
rect -1476 -2811 -1446 -2661
rect -1381 -2811 -1351 -2727
rect -1297 -2811 -1267 -2727
rect -1183 -2811 -1153 -2727
rect -972 -2811 -942 -2611
rect -888 -2811 -858 -2611
rect -700 -2811 -670 -2683
rect -603 -2811 -573 -2611
rect -374 -2811 -344 -2611
rect -129 -2811 -99 -2611
rect -45 -2811 -15 -2611
rect 39 -2811 69 -2611
rect 123 -2811 153 -2611
rect 535 -2805 565 -2677
rect 619 -2805 649 -2677
rect 807 -2811 837 -2727
rect 892 -2811 922 -2727
rect 987 -2811 1017 -2727
rect 1090 -2811 1120 -2727
rect 1222 -2811 1252 -2661
rect 1317 -2811 1347 -2727
rect 1401 -2811 1431 -2727
rect 1515 -2811 1545 -2727
rect 1726 -2811 1756 -2611
rect 1810 -2811 1840 -2611
rect 1998 -2811 2028 -2683
rect 2095 -2811 2125 -2611
rect 2324 -2811 2354 -2611
rect 2569 -2811 2599 -2611
rect 2653 -2811 2683 -2611
rect 2737 -2811 2767 -2611
rect 2821 -2811 2851 -2611
<< ndiff >>
rect -2215 -19 -2163 -7
rect -2215 -53 -2207 -19
rect -2173 -53 -2163 -19
rect -2215 -91 -2163 -53
rect -2133 -45 -2079 -7
rect -2133 -79 -2123 -45
rect -2089 -79 -2079 -45
rect -2133 -91 -2079 -79
rect -2049 -19 -1997 -7
rect -2049 -53 -2039 -19
rect -2005 -53 -1997 -19
rect -2049 -91 -1997 -53
rect -1943 -45 -1891 -7
rect -1943 -79 -1935 -45
rect -1901 -79 -1891 -45
rect -1943 -91 -1891 -79
rect -1861 -19 -1811 -7
rect -1512 -7 -1462 37
rect -1631 -19 -1581 -7
rect -1861 -31 -1779 -19
rect -1861 -65 -1850 -31
rect -1816 -65 -1779 -31
rect -1861 -91 -1779 -65
rect -1749 -31 -1680 -19
rect -1749 -65 -1739 -31
rect -1705 -65 -1680 -31
rect -1749 -91 -1680 -65
rect -1650 -91 -1581 -19
rect -1551 -37 -1462 -7
rect -1551 -71 -1540 -37
rect -1506 -71 -1462 -37
rect -1551 -91 -1462 -71
rect -1432 -19 -1382 37
rect -1022 24 -970 39
rect -1210 -19 -1160 -7
rect -1432 -31 -1361 -19
rect -1432 -65 -1421 -31
rect -1387 -65 -1361 -31
rect -1432 -91 -1361 -65
rect -1331 -31 -1255 -19
rect -1331 -65 -1318 -31
rect -1284 -65 -1255 -31
rect -1331 -91 -1255 -65
rect -1225 -91 -1160 -19
rect -1130 -31 -1078 -7
rect -1130 -65 -1120 -31
rect -1086 -65 -1078 -31
rect -1130 -91 -1078 -65
rect -1022 -10 -1014 24
rect -980 -10 -970 24
rect -1022 -44 -970 -10
rect -1022 -78 -1014 -44
rect -980 -78 -970 -44
rect -1022 -91 -970 -78
rect -940 -15 -886 39
rect -940 -49 -930 -15
rect -896 -49 -886 -15
rect -940 -91 -886 -49
rect -856 26 -804 39
rect -856 -8 -846 26
rect -812 -8 -804 26
rect -653 -7 -603 39
rect -856 -42 -804 -8
rect -856 -76 -846 -42
rect -812 -76 -804 -42
rect -856 -91 -804 -76
rect -750 -19 -698 -7
rect -750 -53 -742 -19
rect -708 -53 -698 -19
rect -750 -91 -698 -53
rect -668 -45 -603 -7
rect -668 -79 -647 -45
rect -613 -79 -603 -45
rect -668 -91 -603 -79
rect -573 -7 -521 39
rect -573 -41 -563 -7
rect -529 -41 -521 -7
rect -573 -91 -521 -41
rect -426 27 -374 39
rect -426 -7 -418 27
rect -384 -7 -374 27
rect -426 -41 -374 -7
rect -426 -75 -418 -41
rect -384 -75 -374 -41
rect -426 -91 -374 -75
rect -344 27 -292 39
rect -344 -7 -334 27
rect -300 -7 -292 27
rect -344 -41 -292 -7
rect -344 -75 -334 -41
rect -300 -75 -292 -41
rect -344 -91 -292 -75
rect -181 -45 -129 39
rect -181 -79 -173 -45
rect -139 -79 -129 -45
rect -181 -91 -129 -79
rect -99 -37 -45 39
rect -99 -71 -89 -37
rect -55 -71 -45 -37
rect -99 -91 -45 -71
rect -15 -45 39 39
rect -15 -79 -5 -45
rect 29 -79 39 -45
rect -15 -91 39 -79
rect 69 -37 123 39
rect 69 -71 79 -37
rect 113 -71 123 -37
rect 69 -91 123 -71
rect 153 -44 205 39
rect 153 -78 163 -44
rect 197 -78 205 -44
rect 153 -91 205 -78
rect -2215 -223 -2163 -185
rect -2215 -257 -2207 -223
rect -2173 -257 -2163 -223
rect -2215 -269 -2163 -257
rect -2133 -197 -2079 -185
rect -2133 -231 -2123 -197
rect -2089 -231 -2079 -197
rect -2133 -269 -2079 -231
rect -2049 -223 -1997 -185
rect -2049 -257 -2039 -223
rect -2005 -257 -1997 -223
rect -2049 -269 -1997 -257
rect -1943 -197 -1891 -185
rect -1943 -231 -1935 -197
rect -1901 -231 -1891 -197
rect -1943 -269 -1891 -231
rect -1861 -211 -1779 -185
rect -1861 -245 -1850 -211
rect -1816 -245 -1779 -211
rect -1861 -257 -1779 -245
rect -1749 -211 -1680 -185
rect -1749 -245 -1739 -211
rect -1705 -245 -1680 -211
rect -1749 -257 -1680 -245
rect -1650 -257 -1581 -185
rect -1861 -269 -1811 -257
rect -1631 -269 -1581 -257
rect -1551 -205 -1462 -185
rect -1551 -239 -1540 -205
rect -1506 -239 -1462 -205
rect -1551 -269 -1462 -239
rect -1512 -313 -1462 -269
rect -1432 -211 -1361 -185
rect -1432 -245 -1421 -211
rect -1387 -245 -1361 -211
rect -1432 -257 -1361 -245
rect -1331 -211 -1255 -185
rect -1331 -245 -1318 -211
rect -1284 -245 -1255 -211
rect -1331 -257 -1255 -245
rect -1225 -257 -1160 -185
rect -1432 -313 -1382 -257
rect -1210 -269 -1160 -257
rect -1130 -211 -1078 -185
rect -1130 -245 -1120 -211
rect -1086 -245 -1078 -211
rect -1130 -269 -1078 -245
rect -1022 -198 -970 -185
rect -1022 -232 -1014 -198
rect -980 -232 -970 -198
rect -1022 -266 -970 -232
rect -1022 -300 -1014 -266
rect -980 -300 -970 -266
rect -1022 -315 -970 -300
rect -940 -227 -886 -185
rect -940 -261 -930 -227
rect -896 -261 -886 -227
rect -940 -315 -886 -261
rect -856 -200 -804 -185
rect -856 -234 -846 -200
rect -812 -234 -804 -200
rect -856 -268 -804 -234
rect -856 -302 -846 -268
rect -812 -302 -804 -268
rect -750 -223 -698 -185
rect -750 -257 -742 -223
rect -708 -257 -698 -223
rect -750 -269 -698 -257
rect -668 -197 -603 -185
rect -668 -231 -647 -197
rect -613 -231 -603 -197
rect -668 -269 -603 -231
rect -856 -315 -804 -302
rect -653 -315 -603 -269
rect -573 -235 -521 -185
rect -573 -269 -563 -235
rect -529 -269 -521 -235
rect -573 -315 -521 -269
rect -426 -201 -374 -185
rect -426 -235 -418 -201
rect -384 -235 -374 -201
rect -426 -269 -374 -235
rect -426 -303 -418 -269
rect -384 -303 -374 -269
rect -426 -315 -374 -303
rect -344 -201 -292 -185
rect -344 -235 -334 -201
rect -300 -235 -292 -201
rect -344 -269 -292 -235
rect -344 -303 -334 -269
rect -300 -303 -292 -269
rect -344 -315 -292 -303
rect -181 -197 -129 -185
rect -181 -231 -173 -197
rect -139 -231 -129 -197
rect -181 -315 -129 -231
rect -99 -205 -45 -185
rect -99 -239 -89 -205
rect -55 -239 -45 -205
rect -99 -315 -45 -239
rect -15 -197 39 -185
rect -15 -231 -5 -197
rect 29 -231 39 -197
rect -15 -315 39 -231
rect 69 -205 123 -185
rect 69 -239 79 -205
rect 113 -239 123 -205
rect 69 -315 123 -239
rect 153 -198 205 -185
rect 153 -232 163 -198
rect 197 -232 205 -198
rect 153 -315 205 -232
rect 483 -223 535 -185
rect 483 -257 491 -223
rect 525 -257 535 -223
rect 483 -269 535 -257
rect 565 -197 619 -185
rect 565 -231 575 -197
rect 609 -231 619 -197
rect 565 -269 619 -231
rect 649 -223 701 -185
rect 649 -257 659 -223
rect 693 -257 701 -223
rect 649 -269 701 -257
rect 755 -197 807 -185
rect 755 -231 763 -197
rect 797 -231 807 -197
rect 755 -269 807 -231
rect 837 -211 919 -185
rect 837 -245 848 -211
rect 882 -245 919 -211
rect 837 -257 919 -245
rect 949 -211 1018 -185
rect 949 -245 959 -211
rect 993 -245 1018 -211
rect 949 -257 1018 -245
rect 1048 -257 1117 -185
rect 837 -269 887 -257
rect 1067 -269 1117 -257
rect 1147 -205 1236 -185
rect 1147 -239 1158 -205
rect 1192 -239 1236 -205
rect 1147 -269 1236 -239
rect 1186 -313 1236 -269
rect 1266 -211 1337 -185
rect 1266 -245 1277 -211
rect 1311 -245 1337 -211
rect 1266 -257 1337 -245
rect 1367 -211 1443 -185
rect 1367 -245 1380 -211
rect 1414 -245 1443 -211
rect 1367 -257 1443 -245
rect 1473 -257 1538 -185
rect 1266 -313 1316 -257
rect 1488 -269 1538 -257
rect 1568 -211 1620 -185
rect 1568 -245 1578 -211
rect 1612 -245 1620 -211
rect 1568 -269 1620 -245
rect 1676 -198 1728 -185
rect 1676 -232 1684 -198
rect 1718 -232 1728 -198
rect 1676 -266 1728 -232
rect 1676 -300 1684 -266
rect 1718 -300 1728 -266
rect 1676 -315 1728 -300
rect 1758 -227 1812 -185
rect 1758 -261 1768 -227
rect 1802 -261 1812 -227
rect 1758 -315 1812 -261
rect 1842 -200 1894 -185
rect 1842 -234 1852 -200
rect 1886 -234 1894 -200
rect 1842 -268 1894 -234
rect 1842 -302 1852 -268
rect 1886 -302 1894 -268
rect 1948 -223 2000 -185
rect 1948 -257 1956 -223
rect 1990 -257 2000 -223
rect 1948 -269 2000 -257
rect 2030 -197 2095 -185
rect 2030 -231 2051 -197
rect 2085 -231 2095 -197
rect 2030 -269 2095 -231
rect 1842 -315 1894 -302
rect 2045 -315 2095 -269
rect 2125 -235 2177 -185
rect 2125 -269 2135 -235
rect 2169 -269 2177 -235
rect 2125 -315 2177 -269
rect 2272 -201 2324 -185
rect 2272 -235 2280 -201
rect 2314 -235 2324 -201
rect 2272 -269 2324 -235
rect 2272 -303 2280 -269
rect 2314 -303 2324 -269
rect 2272 -315 2324 -303
rect 2354 -201 2406 -185
rect 2354 -235 2364 -201
rect 2398 -235 2406 -201
rect 2354 -269 2406 -235
rect 2354 -303 2364 -269
rect 2398 -303 2406 -269
rect 2354 -315 2406 -303
rect 2517 -197 2569 -185
rect 2517 -231 2525 -197
rect 2559 -231 2569 -197
rect 2517 -315 2569 -231
rect 2599 -205 2653 -185
rect 2599 -239 2609 -205
rect 2643 -239 2653 -205
rect 2599 -315 2653 -239
rect 2683 -197 2737 -185
rect 2683 -231 2693 -197
rect 2727 -231 2737 -197
rect 2683 -315 2737 -231
rect 2767 -205 2821 -185
rect 2767 -239 2777 -205
rect 2811 -239 2821 -205
rect 2767 -315 2821 -239
rect 2851 -198 2903 -185
rect 2851 -232 2861 -198
rect 2895 -232 2903 -198
rect 2851 -315 2903 -232
rect -2215 -1107 -2163 -1095
rect -2215 -1141 -2207 -1107
rect -2173 -1141 -2163 -1107
rect -2215 -1179 -2163 -1141
rect -2133 -1133 -2079 -1095
rect -2133 -1167 -2123 -1133
rect -2089 -1167 -2079 -1133
rect -2133 -1179 -2079 -1167
rect -2049 -1107 -1997 -1095
rect -2049 -1141 -2039 -1107
rect -2005 -1141 -1997 -1107
rect -2049 -1179 -1997 -1141
rect -1943 -1133 -1891 -1095
rect -1943 -1167 -1935 -1133
rect -1901 -1167 -1891 -1133
rect -1943 -1179 -1891 -1167
rect -1861 -1107 -1811 -1095
rect -1512 -1095 -1462 -1051
rect -1631 -1107 -1581 -1095
rect -1861 -1119 -1779 -1107
rect -1861 -1153 -1850 -1119
rect -1816 -1153 -1779 -1119
rect -1861 -1179 -1779 -1153
rect -1749 -1119 -1680 -1107
rect -1749 -1153 -1739 -1119
rect -1705 -1153 -1680 -1119
rect -1749 -1179 -1680 -1153
rect -1650 -1179 -1581 -1107
rect -1551 -1125 -1462 -1095
rect -1551 -1159 -1540 -1125
rect -1506 -1159 -1462 -1125
rect -1551 -1179 -1462 -1159
rect -1432 -1107 -1382 -1051
rect -1022 -1064 -970 -1049
rect -1210 -1107 -1160 -1095
rect -1432 -1119 -1361 -1107
rect -1432 -1153 -1421 -1119
rect -1387 -1153 -1361 -1119
rect -1432 -1179 -1361 -1153
rect -1331 -1119 -1255 -1107
rect -1331 -1153 -1318 -1119
rect -1284 -1153 -1255 -1119
rect -1331 -1179 -1255 -1153
rect -1225 -1179 -1160 -1107
rect -1130 -1119 -1078 -1095
rect -1130 -1153 -1120 -1119
rect -1086 -1153 -1078 -1119
rect -1130 -1179 -1078 -1153
rect -1022 -1098 -1014 -1064
rect -980 -1098 -970 -1064
rect -1022 -1132 -970 -1098
rect -1022 -1166 -1014 -1132
rect -980 -1166 -970 -1132
rect -1022 -1179 -970 -1166
rect -940 -1103 -886 -1049
rect -940 -1137 -930 -1103
rect -896 -1137 -886 -1103
rect -940 -1179 -886 -1137
rect -856 -1062 -804 -1049
rect -856 -1096 -846 -1062
rect -812 -1096 -804 -1062
rect -653 -1095 -603 -1049
rect -856 -1130 -804 -1096
rect -856 -1164 -846 -1130
rect -812 -1164 -804 -1130
rect -856 -1179 -804 -1164
rect -750 -1107 -698 -1095
rect -750 -1141 -742 -1107
rect -708 -1141 -698 -1107
rect -750 -1179 -698 -1141
rect -668 -1133 -603 -1095
rect -668 -1167 -647 -1133
rect -613 -1167 -603 -1133
rect -668 -1179 -603 -1167
rect -573 -1095 -521 -1049
rect -573 -1129 -563 -1095
rect -529 -1129 -521 -1095
rect -573 -1179 -521 -1129
rect -426 -1061 -374 -1049
rect -426 -1095 -418 -1061
rect -384 -1095 -374 -1061
rect -426 -1129 -374 -1095
rect -426 -1163 -418 -1129
rect -384 -1163 -374 -1129
rect -426 -1179 -374 -1163
rect -344 -1061 -292 -1049
rect -344 -1095 -334 -1061
rect -300 -1095 -292 -1061
rect -344 -1129 -292 -1095
rect -344 -1163 -334 -1129
rect -300 -1163 -292 -1129
rect -344 -1179 -292 -1163
rect -181 -1133 -129 -1049
rect -181 -1167 -173 -1133
rect -139 -1167 -129 -1133
rect -181 -1179 -129 -1167
rect -99 -1125 -45 -1049
rect -99 -1159 -89 -1125
rect -55 -1159 -45 -1125
rect -99 -1179 -45 -1159
rect -15 -1133 39 -1049
rect -15 -1167 -5 -1133
rect 29 -1167 39 -1133
rect -15 -1179 39 -1167
rect 69 -1125 123 -1049
rect 69 -1159 79 -1125
rect 113 -1159 123 -1125
rect 69 -1179 123 -1159
rect 153 -1132 205 -1049
rect 153 -1166 163 -1132
rect 197 -1166 205 -1132
rect 153 -1179 205 -1166
rect 483 -1107 535 -1095
rect 483 -1141 491 -1107
rect 525 -1141 535 -1107
rect 483 -1179 535 -1141
rect 565 -1133 619 -1095
rect 565 -1167 575 -1133
rect 609 -1167 619 -1133
rect 565 -1179 619 -1167
rect 649 -1107 701 -1095
rect 649 -1141 659 -1107
rect 693 -1141 701 -1107
rect 649 -1179 701 -1141
rect 755 -1133 807 -1095
rect 755 -1167 763 -1133
rect 797 -1167 807 -1133
rect 755 -1179 807 -1167
rect 837 -1107 887 -1095
rect 1186 -1095 1236 -1051
rect 1067 -1107 1117 -1095
rect 837 -1119 919 -1107
rect 837 -1153 848 -1119
rect 882 -1153 919 -1119
rect 837 -1179 919 -1153
rect 949 -1119 1018 -1107
rect 949 -1153 959 -1119
rect 993 -1153 1018 -1119
rect 949 -1179 1018 -1153
rect 1048 -1179 1117 -1107
rect 1147 -1125 1236 -1095
rect 1147 -1159 1158 -1125
rect 1192 -1159 1236 -1125
rect 1147 -1179 1236 -1159
rect 1266 -1107 1316 -1051
rect 1676 -1064 1728 -1049
rect 1488 -1107 1538 -1095
rect 1266 -1119 1337 -1107
rect 1266 -1153 1277 -1119
rect 1311 -1153 1337 -1119
rect 1266 -1179 1337 -1153
rect 1367 -1119 1443 -1107
rect 1367 -1153 1380 -1119
rect 1414 -1153 1443 -1119
rect 1367 -1179 1443 -1153
rect 1473 -1179 1538 -1107
rect 1568 -1119 1620 -1095
rect 1568 -1153 1578 -1119
rect 1612 -1153 1620 -1119
rect 1568 -1179 1620 -1153
rect 1676 -1098 1684 -1064
rect 1718 -1098 1728 -1064
rect 1676 -1132 1728 -1098
rect 1676 -1166 1684 -1132
rect 1718 -1166 1728 -1132
rect 1676 -1179 1728 -1166
rect 1758 -1103 1812 -1049
rect 1758 -1137 1768 -1103
rect 1802 -1137 1812 -1103
rect 1758 -1179 1812 -1137
rect 1842 -1062 1894 -1049
rect 1842 -1096 1852 -1062
rect 1886 -1096 1894 -1062
rect 2045 -1095 2095 -1049
rect 1842 -1130 1894 -1096
rect 1842 -1164 1852 -1130
rect 1886 -1164 1894 -1130
rect 1842 -1179 1894 -1164
rect 1948 -1107 2000 -1095
rect 1948 -1141 1956 -1107
rect 1990 -1141 2000 -1107
rect 1948 -1179 2000 -1141
rect 2030 -1133 2095 -1095
rect 2030 -1167 2051 -1133
rect 2085 -1167 2095 -1133
rect 2030 -1179 2095 -1167
rect 2125 -1095 2177 -1049
rect 2125 -1129 2135 -1095
rect 2169 -1129 2177 -1095
rect 2125 -1179 2177 -1129
rect 2272 -1061 2324 -1049
rect 2272 -1095 2280 -1061
rect 2314 -1095 2324 -1061
rect 2272 -1129 2324 -1095
rect 2272 -1163 2280 -1129
rect 2314 -1163 2324 -1129
rect 2272 -1179 2324 -1163
rect 2354 -1061 2406 -1049
rect 2354 -1095 2364 -1061
rect 2398 -1095 2406 -1061
rect 2354 -1129 2406 -1095
rect 2354 -1163 2364 -1129
rect 2398 -1163 2406 -1129
rect 2354 -1179 2406 -1163
rect 2517 -1133 2569 -1049
rect 2517 -1167 2525 -1133
rect 2559 -1167 2569 -1133
rect 2517 -1179 2569 -1167
rect 2599 -1125 2653 -1049
rect 2599 -1159 2609 -1125
rect 2643 -1159 2653 -1125
rect 2599 -1179 2653 -1159
rect 2683 -1133 2737 -1049
rect 2683 -1167 2693 -1133
rect 2727 -1167 2737 -1133
rect 2683 -1179 2737 -1167
rect 2767 -1125 2821 -1049
rect 2767 -1159 2777 -1125
rect 2811 -1159 2821 -1125
rect 2767 -1179 2821 -1159
rect 2851 -1132 2903 -1049
rect 2851 -1166 2861 -1132
rect 2895 -1166 2903 -1132
rect 2851 -1179 2903 -1166
rect -2215 -1311 -2163 -1273
rect -2215 -1345 -2207 -1311
rect -2173 -1345 -2163 -1311
rect -2215 -1357 -2163 -1345
rect -2133 -1285 -2079 -1273
rect -2133 -1319 -2123 -1285
rect -2089 -1319 -2079 -1285
rect -2133 -1357 -2079 -1319
rect -2049 -1311 -1997 -1273
rect -2049 -1345 -2039 -1311
rect -2005 -1345 -1997 -1311
rect -2049 -1357 -1997 -1345
rect -1943 -1285 -1891 -1273
rect -1943 -1319 -1935 -1285
rect -1901 -1319 -1891 -1285
rect -1943 -1357 -1891 -1319
rect -1861 -1299 -1779 -1273
rect -1861 -1333 -1850 -1299
rect -1816 -1333 -1779 -1299
rect -1861 -1345 -1779 -1333
rect -1749 -1299 -1680 -1273
rect -1749 -1333 -1739 -1299
rect -1705 -1333 -1680 -1299
rect -1749 -1345 -1680 -1333
rect -1650 -1345 -1581 -1273
rect -1861 -1357 -1811 -1345
rect -1631 -1357 -1581 -1345
rect -1551 -1293 -1462 -1273
rect -1551 -1327 -1540 -1293
rect -1506 -1327 -1462 -1293
rect -1551 -1357 -1462 -1327
rect -1512 -1401 -1462 -1357
rect -1432 -1299 -1361 -1273
rect -1432 -1333 -1421 -1299
rect -1387 -1333 -1361 -1299
rect -1432 -1345 -1361 -1333
rect -1331 -1299 -1255 -1273
rect -1331 -1333 -1318 -1299
rect -1284 -1333 -1255 -1299
rect -1331 -1345 -1255 -1333
rect -1225 -1345 -1160 -1273
rect -1432 -1401 -1382 -1345
rect -1210 -1357 -1160 -1345
rect -1130 -1299 -1078 -1273
rect -1130 -1333 -1120 -1299
rect -1086 -1333 -1078 -1299
rect -1130 -1357 -1078 -1333
rect -1022 -1286 -970 -1273
rect -1022 -1320 -1014 -1286
rect -980 -1320 -970 -1286
rect -1022 -1354 -970 -1320
rect -1022 -1388 -1014 -1354
rect -980 -1388 -970 -1354
rect -1022 -1403 -970 -1388
rect -940 -1315 -886 -1273
rect -940 -1349 -930 -1315
rect -896 -1349 -886 -1315
rect -940 -1403 -886 -1349
rect -856 -1288 -804 -1273
rect -856 -1322 -846 -1288
rect -812 -1322 -804 -1288
rect -856 -1356 -804 -1322
rect -856 -1390 -846 -1356
rect -812 -1390 -804 -1356
rect -750 -1311 -698 -1273
rect -750 -1345 -742 -1311
rect -708 -1345 -698 -1311
rect -750 -1357 -698 -1345
rect -668 -1285 -603 -1273
rect -668 -1319 -647 -1285
rect -613 -1319 -603 -1285
rect -668 -1357 -603 -1319
rect -856 -1403 -804 -1390
rect -653 -1403 -603 -1357
rect -573 -1323 -521 -1273
rect -573 -1357 -563 -1323
rect -529 -1357 -521 -1323
rect -573 -1403 -521 -1357
rect -426 -1289 -374 -1273
rect -426 -1323 -418 -1289
rect -384 -1323 -374 -1289
rect -426 -1357 -374 -1323
rect -426 -1391 -418 -1357
rect -384 -1391 -374 -1357
rect -426 -1403 -374 -1391
rect -344 -1289 -292 -1273
rect -344 -1323 -334 -1289
rect -300 -1323 -292 -1289
rect -344 -1357 -292 -1323
rect -344 -1391 -334 -1357
rect -300 -1391 -292 -1357
rect -344 -1403 -292 -1391
rect -181 -1285 -129 -1273
rect -181 -1319 -173 -1285
rect -139 -1319 -129 -1285
rect -181 -1403 -129 -1319
rect -99 -1293 -45 -1273
rect -99 -1327 -89 -1293
rect -55 -1327 -45 -1293
rect -99 -1403 -45 -1327
rect -15 -1285 39 -1273
rect -15 -1319 -5 -1285
rect 29 -1319 39 -1285
rect -15 -1403 39 -1319
rect 69 -1293 123 -1273
rect 69 -1327 79 -1293
rect 113 -1327 123 -1293
rect 69 -1403 123 -1327
rect 153 -1286 205 -1273
rect 153 -1320 163 -1286
rect 197 -1320 205 -1286
rect 153 -1403 205 -1320
rect 483 -1311 535 -1273
rect 483 -1345 491 -1311
rect 525 -1345 535 -1311
rect 483 -1357 535 -1345
rect 565 -1285 619 -1273
rect 565 -1319 575 -1285
rect 609 -1319 619 -1285
rect 565 -1357 619 -1319
rect 649 -1311 701 -1273
rect 649 -1345 659 -1311
rect 693 -1345 701 -1311
rect 649 -1357 701 -1345
rect 755 -1285 807 -1273
rect 755 -1319 763 -1285
rect 797 -1319 807 -1285
rect 755 -1357 807 -1319
rect 837 -1299 919 -1273
rect 837 -1333 848 -1299
rect 882 -1333 919 -1299
rect 837 -1345 919 -1333
rect 949 -1299 1018 -1273
rect 949 -1333 959 -1299
rect 993 -1333 1018 -1299
rect 949 -1345 1018 -1333
rect 1048 -1345 1117 -1273
rect 837 -1357 887 -1345
rect 1067 -1357 1117 -1345
rect 1147 -1293 1236 -1273
rect 1147 -1327 1158 -1293
rect 1192 -1327 1236 -1293
rect 1147 -1357 1236 -1327
rect 1186 -1401 1236 -1357
rect 1266 -1299 1337 -1273
rect 1266 -1333 1277 -1299
rect 1311 -1333 1337 -1299
rect 1266 -1345 1337 -1333
rect 1367 -1299 1443 -1273
rect 1367 -1333 1380 -1299
rect 1414 -1333 1443 -1299
rect 1367 -1345 1443 -1333
rect 1473 -1345 1538 -1273
rect 1266 -1401 1316 -1345
rect 1488 -1357 1538 -1345
rect 1568 -1299 1620 -1273
rect 1568 -1333 1578 -1299
rect 1612 -1333 1620 -1299
rect 1568 -1357 1620 -1333
rect 1676 -1286 1728 -1273
rect 1676 -1320 1684 -1286
rect 1718 -1320 1728 -1286
rect 1676 -1354 1728 -1320
rect 1676 -1388 1684 -1354
rect 1718 -1388 1728 -1354
rect 1676 -1403 1728 -1388
rect 1758 -1315 1812 -1273
rect 1758 -1349 1768 -1315
rect 1802 -1349 1812 -1315
rect 1758 -1403 1812 -1349
rect 1842 -1288 1894 -1273
rect 1842 -1322 1852 -1288
rect 1886 -1322 1894 -1288
rect 1842 -1356 1894 -1322
rect 1842 -1390 1852 -1356
rect 1886 -1390 1894 -1356
rect 1948 -1311 2000 -1273
rect 1948 -1345 1956 -1311
rect 1990 -1345 2000 -1311
rect 1948 -1357 2000 -1345
rect 2030 -1285 2095 -1273
rect 2030 -1319 2051 -1285
rect 2085 -1319 2095 -1285
rect 2030 -1357 2095 -1319
rect 1842 -1403 1894 -1390
rect 2045 -1403 2095 -1357
rect 2125 -1323 2177 -1273
rect 2125 -1357 2135 -1323
rect 2169 -1357 2177 -1323
rect 2125 -1403 2177 -1357
rect 2272 -1289 2324 -1273
rect 2272 -1323 2280 -1289
rect 2314 -1323 2324 -1289
rect 2272 -1357 2324 -1323
rect 2272 -1391 2280 -1357
rect 2314 -1391 2324 -1357
rect 2272 -1403 2324 -1391
rect 2354 -1289 2406 -1273
rect 2354 -1323 2364 -1289
rect 2398 -1323 2406 -1289
rect 2354 -1357 2406 -1323
rect 2354 -1391 2364 -1357
rect 2398 -1391 2406 -1357
rect 2354 -1403 2406 -1391
rect 2517 -1285 2569 -1273
rect 2517 -1319 2525 -1285
rect 2559 -1319 2569 -1285
rect 2517 -1403 2569 -1319
rect 2599 -1293 2653 -1273
rect 2599 -1327 2609 -1293
rect 2643 -1327 2653 -1293
rect 2599 -1403 2653 -1327
rect 2683 -1285 2737 -1273
rect 2683 -1319 2693 -1285
rect 2727 -1319 2737 -1285
rect 2683 -1403 2737 -1319
rect 2767 -1293 2821 -1273
rect 2767 -1327 2777 -1293
rect 2811 -1327 2821 -1293
rect 2767 -1403 2821 -1327
rect 2851 -1286 2903 -1273
rect 2851 -1320 2861 -1286
rect 2895 -1320 2903 -1286
rect 2851 -1403 2903 -1320
rect -2215 -2195 -2163 -2183
rect -2215 -2229 -2207 -2195
rect -2173 -2229 -2163 -2195
rect -2215 -2267 -2163 -2229
rect -2133 -2221 -2079 -2183
rect -2133 -2255 -2123 -2221
rect -2089 -2255 -2079 -2221
rect -2133 -2267 -2079 -2255
rect -2049 -2195 -1997 -2183
rect -2049 -2229 -2039 -2195
rect -2005 -2229 -1997 -2195
rect -2049 -2267 -1997 -2229
rect -1943 -2221 -1891 -2183
rect -1943 -2255 -1935 -2221
rect -1901 -2255 -1891 -2221
rect -1943 -2267 -1891 -2255
rect -1861 -2195 -1811 -2183
rect -1512 -2183 -1462 -2139
rect -1631 -2195 -1581 -2183
rect -1861 -2207 -1779 -2195
rect -1861 -2241 -1850 -2207
rect -1816 -2241 -1779 -2207
rect -1861 -2267 -1779 -2241
rect -1749 -2207 -1680 -2195
rect -1749 -2241 -1739 -2207
rect -1705 -2241 -1680 -2207
rect -1749 -2267 -1680 -2241
rect -1650 -2267 -1581 -2195
rect -1551 -2213 -1462 -2183
rect -1551 -2247 -1540 -2213
rect -1506 -2247 -1462 -2213
rect -1551 -2267 -1462 -2247
rect -1432 -2195 -1382 -2139
rect -1022 -2152 -970 -2137
rect -1210 -2195 -1160 -2183
rect -1432 -2207 -1361 -2195
rect -1432 -2241 -1421 -2207
rect -1387 -2241 -1361 -2207
rect -1432 -2267 -1361 -2241
rect -1331 -2207 -1255 -2195
rect -1331 -2241 -1318 -2207
rect -1284 -2241 -1255 -2207
rect -1331 -2267 -1255 -2241
rect -1225 -2267 -1160 -2195
rect -1130 -2207 -1078 -2183
rect -1130 -2241 -1120 -2207
rect -1086 -2241 -1078 -2207
rect -1130 -2267 -1078 -2241
rect -1022 -2186 -1014 -2152
rect -980 -2186 -970 -2152
rect -1022 -2220 -970 -2186
rect -1022 -2254 -1014 -2220
rect -980 -2254 -970 -2220
rect -1022 -2267 -970 -2254
rect -940 -2191 -886 -2137
rect -940 -2225 -930 -2191
rect -896 -2225 -886 -2191
rect -940 -2267 -886 -2225
rect -856 -2150 -804 -2137
rect -856 -2184 -846 -2150
rect -812 -2184 -804 -2150
rect -653 -2183 -603 -2137
rect -856 -2218 -804 -2184
rect -856 -2252 -846 -2218
rect -812 -2252 -804 -2218
rect -856 -2267 -804 -2252
rect -750 -2195 -698 -2183
rect -750 -2229 -742 -2195
rect -708 -2229 -698 -2195
rect -750 -2267 -698 -2229
rect -668 -2221 -603 -2183
rect -668 -2255 -647 -2221
rect -613 -2255 -603 -2221
rect -668 -2267 -603 -2255
rect -573 -2183 -521 -2137
rect -573 -2217 -563 -2183
rect -529 -2217 -521 -2183
rect -573 -2267 -521 -2217
rect -426 -2149 -374 -2137
rect -426 -2183 -418 -2149
rect -384 -2183 -374 -2149
rect -426 -2217 -374 -2183
rect -426 -2251 -418 -2217
rect -384 -2251 -374 -2217
rect -426 -2267 -374 -2251
rect -344 -2149 -292 -2137
rect -344 -2183 -334 -2149
rect -300 -2183 -292 -2149
rect -344 -2217 -292 -2183
rect -344 -2251 -334 -2217
rect -300 -2251 -292 -2217
rect -344 -2267 -292 -2251
rect -181 -2221 -129 -2137
rect -181 -2255 -173 -2221
rect -139 -2255 -129 -2221
rect -181 -2267 -129 -2255
rect -99 -2213 -45 -2137
rect -99 -2247 -89 -2213
rect -55 -2247 -45 -2213
rect -99 -2267 -45 -2247
rect -15 -2221 39 -2137
rect -15 -2255 -5 -2221
rect 29 -2255 39 -2221
rect -15 -2267 39 -2255
rect 69 -2213 123 -2137
rect 69 -2247 79 -2213
rect 113 -2247 123 -2213
rect 69 -2267 123 -2247
rect 153 -2220 205 -2137
rect 153 -2254 163 -2220
rect 197 -2254 205 -2220
rect 153 -2267 205 -2254
rect 483 -2195 535 -2183
rect 483 -2229 491 -2195
rect 525 -2229 535 -2195
rect 483 -2267 535 -2229
rect 565 -2221 619 -2183
rect 565 -2255 575 -2221
rect 609 -2255 619 -2221
rect 565 -2267 619 -2255
rect 649 -2195 701 -2183
rect 649 -2229 659 -2195
rect 693 -2229 701 -2195
rect 649 -2267 701 -2229
rect 755 -2221 807 -2183
rect 755 -2255 763 -2221
rect 797 -2255 807 -2221
rect 755 -2267 807 -2255
rect 837 -2195 887 -2183
rect 1186 -2183 1236 -2139
rect 1067 -2195 1117 -2183
rect 837 -2207 919 -2195
rect 837 -2241 848 -2207
rect 882 -2241 919 -2207
rect 837 -2267 919 -2241
rect 949 -2207 1018 -2195
rect 949 -2241 959 -2207
rect 993 -2241 1018 -2207
rect 949 -2267 1018 -2241
rect 1048 -2267 1117 -2195
rect 1147 -2213 1236 -2183
rect 1147 -2247 1158 -2213
rect 1192 -2247 1236 -2213
rect 1147 -2267 1236 -2247
rect 1266 -2195 1316 -2139
rect 1676 -2152 1728 -2137
rect 1488 -2195 1538 -2183
rect 1266 -2207 1337 -2195
rect 1266 -2241 1277 -2207
rect 1311 -2241 1337 -2207
rect 1266 -2267 1337 -2241
rect 1367 -2207 1443 -2195
rect 1367 -2241 1380 -2207
rect 1414 -2241 1443 -2207
rect 1367 -2267 1443 -2241
rect 1473 -2267 1538 -2195
rect 1568 -2207 1620 -2183
rect 1568 -2241 1578 -2207
rect 1612 -2241 1620 -2207
rect 1568 -2267 1620 -2241
rect 1676 -2186 1684 -2152
rect 1718 -2186 1728 -2152
rect 1676 -2220 1728 -2186
rect 1676 -2254 1684 -2220
rect 1718 -2254 1728 -2220
rect 1676 -2267 1728 -2254
rect 1758 -2191 1812 -2137
rect 1758 -2225 1768 -2191
rect 1802 -2225 1812 -2191
rect 1758 -2267 1812 -2225
rect 1842 -2150 1894 -2137
rect 1842 -2184 1852 -2150
rect 1886 -2184 1894 -2150
rect 2045 -2183 2095 -2137
rect 1842 -2218 1894 -2184
rect 1842 -2252 1852 -2218
rect 1886 -2252 1894 -2218
rect 1842 -2267 1894 -2252
rect 1948 -2195 2000 -2183
rect 1948 -2229 1956 -2195
rect 1990 -2229 2000 -2195
rect 1948 -2267 2000 -2229
rect 2030 -2221 2095 -2183
rect 2030 -2255 2051 -2221
rect 2085 -2255 2095 -2221
rect 2030 -2267 2095 -2255
rect 2125 -2183 2177 -2137
rect 2125 -2217 2135 -2183
rect 2169 -2217 2177 -2183
rect 2125 -2267 2177 -2217
rect 2272 -2149 2324 -2137
rect 2272 -2183 2280 -2149
rect 2314 -2183 2324 -2149
rect 2272 -2217 2324 -2183
rect 2272 -2251 2280 -2217
rect 2314 -2251 2324 -2217
rect 2272 -2267 2324 -2251
rect 2354 -2149 2406 -2137
rect 2354 -2183 2364 -2149
rect 2398 -2183 2406 -2149
rect 2354 -2217 2406 -2183
rect 2354 -2251 2364 -2217
rect 2398 -2251 2406 -2217
rect 2354 -2267 2406 -2251
rect 2517 -2221 2569 -2137
rect 2517 -2255 2525 -2221
rect 2559 -2255 2569 -2221
rect 2517 -2267 2569 -2255
rect 2599 -2213 2653 -2137
rect 2599 -2247 2609 -2213
rect 2643 -2247 2653 -2213
rect 2599 -2267 2653 -2247
rect 2683 -2221 2737 -2137
rect 2683 -2255 2693 -2221
rect 2727 -2255 2737 -2221
rect 2683 -2267 2737 -2255
rect 2767 -2213 2821 -2137
rect 2767 -2247 2777 -2213
rect 2811 -2247 2821 -2213
rect 2767 -2267 2821 -2247
rect 2851 -2220 2903 -2137
rect 2851 -2254 2861 -2220
rect 2895 -2254 2903 -2220
rect 2851 -2267 2903 -2254
rect -2215 -2399 -2163 -2361
rect -2215 -2433 -2207 -2399
rect -2173 -2433 -2163 -2399
rect -2215 -2445 -2163 -2433
rect -2133 -2373 -2079 -2361
rect -2133 -2407 -2123 -2373
rect -2089 -2407 -2079 -2373
rect -2133 -2445 -2079 -2407
rect -2049 -2399 -1997 -2361
rect -2049 -2433 -2039 -2399
rect -2005 -2433 -1997 -2399
rect -2049 -2445 -1997 -2433
rect -1943 -2373 -1891 -2361
rect -1943 -2407 -1935 -2373
rect -1901 -2407 -1891 -2373
rect -1943 -2445 -1891 -2407
rect -1861 -2387 -1779 -2361
rect -1861 -2421 -1850 -2387
rect -1816 -2421 -1779 -2387
rect -1861 -2433 -1779 -2421
rect -1749 -2387 -1680 -2361
rect -1749 -2421 -1739 -2387
rect -1705 -2421 -1680 -2387
rect -1749 -2433 -1680 -2421
rect -1650 -2433 -1581 -2361
rect -1861 -2445 -1811 -2433
rect -1631 -2445 -1581 -2433
rect -1551 -2381 -1462 -2361
rect -1551 -2415 -1540 -2381
rect -1506 -2415 -1462 -2381
rect -1551 -2445 -1462 -2415
rect -1512 -2489 -1462 -2445
rect -1432 -2387 -1361 -2361
rect -1432 -2421 -1421 -2387
rect -1387 -2421 -1361 -2387
rect -1432 -2433 -1361 -2421
rect -1331 -2387 -1255 -2361
rect -1331 -2421 -1318 -2387
rect -1284 -2421 -1255 -2387
rect -1331 -2433 -1255 -2421
rect -1225 -2433 -1160 -2361
rect -1432 -2489 -1382 -2433
rect -1210 -2445 -1160 -2433
rect -1130 -2387 -1078 -2361
rect -1130 -2421 -1120 -2387
rect -1086 -2421 -1078 -2387
rect -1130 -2445 -1078 -2421
rect -1022 -2374 -970 -2361
rect -1022 -2408 -1014 -2374
rect -980 -2408 -970 -2374
rect -1022 -2442 -970 -2408
rect -1022 -2476 -1014 -2442
rect -980 -2476 -970 -2442
rect -1022 -2491 -970 -2476
rect -940 -2403 -886 -2361
rect -940 -2437 -930 -2403
rect -896 -2437 -886 -2403
rect -940 -2491 -886 -2437
rect -856 -2376 -804 -2361
rect -856 -2410 -846 -2376
rect -812 -2410 -804 -2376
rect -856 -2444 -804 -2410
rect -856 -2478 -846 -2444
rect -812 -2478 -804 -2444
rect -750 -2399 -698 -2361
rect -750 -2433 -742 -2399
rect -708 -2433 -698 -2399
rect -750 -2445 -698 -2433
rect -668 -2373 -603 -2361
rect -668 -2407 -647 -2373
rect -613 -2407 -603 -2373
rect -668 -2445 -603 -2407
rect -856 -2491 -804 -2478
rect -653 -2491 -603 -2445
rect -573 -2411 -521 -2361
rect -573 -2445 -563 -2411
rect -529 -2445 -521 -2411
rect -573 -2491 -521 -2445
rect -426 -2377 -374 -2361
rect -426 -2411 -418 -2377
rect -384 -2411 -374 -2377
rect -426 -2445 -374 -2411
rect -426 -2479 -418 -2445
rect -384 -2479 -374 -2445
rect -426 -2491 -374 -2479
rect -344 -2377 -292 -2361
rect -344 -2411 -334 -2377
rect -300 -2411 -292 -2377
rect -344 -2445 -292 -2411
rect -344 -2479 -334 -2445
rect -300 -2479 -292 -2445
rect -344 -2491 -292 -2479
rect -181 -2373 -129 -2361
rect -181 -2407 -173 -2373
rect -139 -2407 -129 -2373
rect -181 -2491 -129 -2407
rect -99 -2381 -45 -2361
rect -99 -2415 -89 -2381
rect -55 -2415 -45 -2381
rect -99 -2491 -45 -2415
rect -15 -2373 39 -2361
rect -15 -2407 -5 -2373
rect 29 -2407 39 -2373
rect -15 -2491 39 -2407
rect 69 -2381 123 -2361
rect 69 -2415 79 -2381
rect 113 -2415 123 -2381
rect 69 -2491 123 -2415
rect 153 -2374 205 -2361
rect 153 -2408 163 -2374
rect 197 -2408 205 -2374
rect 153 -2491 205 -2408
rect 483 -2399 535 -2361
rect 483 -2433 491 -2399
rect 525 -2433 535 -2399
rect 483 -2445 535 -2433
rect 565 -2373 619 -2361
rect 565 -2407 575 -2373
rect 609 -2407 619 -2373
rect 565 -2445 619 -2407
rect 649 -2399 701 -2361
rect 649 -2433 659 -2399
rect 693 -2433 701 -2399
rect 649 -2445 701 -2433
rect 755 -2373 807 -2361
rect 755 -2407 763 -2373
rect 797 -2407 807 -2373
rect 755 -2445 807 -2407
rect 837 -2387 919 -2361
rect 837 -2421 848 -2387
rect 882 -2421 919 -2387
rect 837 -2433 919 -2421
rect 949 -2387 1018 -2361
rect 949 -2421 959 -2387
rect 993 -2421 1018 -2387
rect 949 -2433 1018 -2421
rect 1048 -2433 1117 -2361
rect 837 -2445 887 -2433
rect 1067 -2445 1117 -2433
rect 1147 -2381 1236 -2361
rect 1147 -2415 1158 -2381
rect 1192 -2415 1236 -2381
rect 1147 -2445 1236 -2415
rect 1186 -2489 1236 -2445
rect 1266 -2387 1337 -2361
rect 1266 -2421 1277 -2387
rect 1311 -2421 1337 -2387
rect 1266 -2433 1337 -2421
rect 1367 -2387 1443 -2361
rect 1367 -2421 1380 -2387
rect 1414 -2421 1443 -2387
rect 1367 -2433 1443 -2421
rect 1473 -2433 1538 -2361
rect 1266 -2489 1316 -2433
rect 1488 -2445 1538 -2433
rect 1568 -2387 1620 -2361
rect 1568 -2421 1578 -2387
rect 1612 -2421 1620 -2387
rect 1568 -2445 1620 -2421
rect 1676 -2374 1728 -2361
rect 1676 -2408 1684 -2374
rect 1718 -2408 1728 -2374
rect 1676 -2442 1728 -2408
rect 1676 -2476 1684 -2442
rect 1718 -2476 1728 -2442
rect 1676 -2491 1728 -2476
rect 1758 -2403 1812 -2361
rect 1758 -2437 1768 -2403
rect 1802 -2437 1812 -2403
rect 1758 -2491 1812 -2437
rect 1842 -2376 1894 -2361
rect 1842 -2410 1852 -2376
rect 1886 -2410 1894 -2376
rect 1842 -2444 1894 -2410
rect 1842 -2478 1852 -2444
rect 1886 -2478 1894 -2444
rect 1948 -2399 2000 -2361
rect 1948 -2433 1956 -2399
rect 1990 -2433 2000 -2399
rect 1948 -2445 2000 -2433
rect 2030 -2373 2095 -2361
rect 2030 -2407 2051 -2373
rect 2085 -2407 2095 -2373
rect 2030 -2445 2095 -2407
rect 1842 -2491 1894 -2478
rect 2045 -2491 2095 -2445
rect 2125 -2411 2177 -2361
rect 2125 -2445 2135 -2411
rect 2169 -2445 2177 -2411
rect 2125 -2491 2177 -2445
rect 2272 -2377 2324 -2361
rect 2272 -2411 2280 -2377
rect 2314 -2411 2324 -2377
rect 2272 -2445 2324 -2411
rect 2272 -2479 2280 -2445
rect 2314 -2479 2324 -2445
rect 2272 -2491 2324 -2479
rect 2354 -2377 2406 -2361
rect 2354 -2411 2364 -2377
rect 2398 -2411 2406 -2377
rect 2354 -2445 2406 -2411
rect 2354 -2479 2364 -2445
rect 2398 -2479 2406 -2445
rect 2354 -2491 2406 -2479
rect 2517 -2373 2569 -2361
rect 2517 -2407 2525 -2373
rect 2559 -2407 2569 -2373
rect 2517 -2491 2569 -2407
rect 2599 -2381 2653 -2361
rect 2599 -2415 2609 -2381
rect 2643 -2415 2653 -2381
rect 2599 -2491 2653 -2415
rect 2683 -2373 2737 -2361
rect 2683 -2407 2693 -2373
rect 2727 -2407 2737 -2373
rect 2683 -2491 2737 -2407
rect 2767 -2381 2821 -2361
rect 2767 -2415 2777 -2381
rect 2811 -2415 2821 -2381
rect 2767 -2491 2821 -2415
rect 2851 -2374 2903 -2361
rect 2851 -2408 2861 -2374
rect 2895 -2408 2903 -2374
rect 2851 -2491 2903 -2408
<< pdiff >>
rect -2215 339 -2163 353
rect -2215 305 -2207 339
rect -2173 305 -2163 339
rect -2215 271 -2163 305
rect -2215 237 -2207 271
rect -2173 237 -2163 271
rect -2215 225 -2163 237
rect -2133 323 -2079 353
rect -2133 289 -2123 323
rect -2089 289 -2079 323
rect -2133 225 -2079 289
rect -2049 339 -1997 353
rect -2049 305 -2039 339
rect -2005 305 -1997 339
rect -2049 271 -1997 305
rect -1943 347 -1891 359
rect -1943 313 -1935 347
rect -1901 313 -1891 347
rect -1943 275 -1891 313
rect -1861 339 -1806 359
rect -1861 305 -1851 339
rect -1817 305 -1806 339
rect -1861 275 -1806 305
rect -1776 334 -1711 359
rect -1776 300 -1759 334
rect -1725 300 -1711 334
rect -1776 275 -1711 300
rect -1681 275 -1608 359
rect -1578 347 -1476 359
rect -1578 313 -1520 347
rect -1486 313 -1476 347
rect -1578 279 -1476 313
rect -1578 275 -1520 279
rect -2049 237 -2039 271
rect -2005 237 -1997 271
rect -2049 225 -1997 237
rect -1563 245 -1520 275
rect -1486 245 -1476 279
rect -1563 209 -1476 245
rect -1446 339 -1381 359
rect -1446 305 -1436 339
rect -1402 305 -1381 339
rect -1446 275 -1381 305
rect -1351 329 -1297 359
rect -1351 295 -1341 329
rect -1307 295 -1297 329
rect -1351 275 -1297 295
rect -1267 275 -1183 359
rect -1153 339 -1100 359
rect -1153 305 -1142 339
rect -1108 305 -1100 339
rect -1153 275 -1100 305
rect -1026 347 -972 359
rect -1026 313 -1018 347
rect -984 313 -972 347
rect -1026 276 -972 313
rect -1446 209 -1396 275
rect -1026 242 -1018 276
rect -984 242 -972 276
rect -1026 205 -972 242
rect -1026 171 -1018 205
rect -984 171 -972 205
rect -1026 159 -972 171
rect -942 317 -888 359
rect -942 283 -932 317
rect -898 283 -888 317
rect -942 237 -888 283
rect -942 203 -932 237
rect -898 203 -888 237
rect -942 159 -888 203
rect -858 341 -806 359
rect -858 307 -848 341
rect -814 307 -806 341
rect -858 273 -806 307
rect -858 239 -848 273
rect -814 239 -806 273
rect -858 205 -806 239
rect -752 347 -700 359
rect -752 313 -744 347
rect -710 313 -700 347
rect -752 279 -700 313
rect -752 245 -744 279
rect -710 245 -700 279
rect -752 231 -700 245
rect -670 347 -603 359
rect -670 313 -647 347
rect -613 313 -603 347
rect -670 279 -603 313
rect -670 245 -647 279
rect -613 245 -603 279
rect -670 231 -603 245
rect -858 171 -848 205
rect -814 171 -806 205
rect -858 159 -806 171
rect -655 211 -603 231
rect -655 177 -647 211
rect -613 177 -603 211
rect -655 159 -603 177
rect -573 347 -521 359
rect -573 313 -563 347
rect -529 313 -521 347
rect -573 276 -521 313
rect -573 242 -563 276
rect -529 242 -521 276
rect -573 205 -521 242
rect -573 171 -563 205
rect -529 171 -521 205
rect -573 159 -521 171
rect -426 347 -374 359
rect -426 313 -418 347
rect -384 313 -374 347
rect -426 279 -374 313
rect -426 245 -418 279
rect -384 245 -374 279
rect -426 211 -374 245
rect -426 177 -418 211
rect -384 177 -374 211
rect -426 159 -374 177
rect -344 347 -292 359
rect -344 313 -334 347
rect -300 313 -292 347
rect -344 279 -292 313
rect -344 245 -334 279
rect -300 245 -292 279
rect -344 211 -292 245
rect -344 177 -334 211
rect -300 177 -292 211
rect -344 159 -292 177
rect -181 347 -129 359
rect -181 313 -173 347
rect -139 313 -129 347
rect -181 279 -129 313
rect -181 245 -173 279
rect -139 245 -129 279
rect -181 211 -129 245
rect -181 177 -173 211
rect -139 177 -129 211
rect -181 159 -129 177
rect -99 347 -45 359
rect -99 313 -89 347
rect -55 313 -45 347
rect -99 279 -45 313
rect -99 245 -89 279
rect -55 245 -45 279
rect -99 211 -45 245
rect -99 177 -89 211
rect -55 177 -45 211
rect -99 159 -45 177
rect -15 347 39 359
rect -15 313 -5 347
rect 29 313 39 347
rect -15 279 39 313
rect -15 245 -5 279
rect 29 245 39 279
rect -15 159 39 245
rect 69 347 123 359
rect 69 313 79 347
rect 113 313 123 347
rect 69 279 123 313
rect 69 245 79 279
rect 113 245 123 279
rect 69 211 123 245
rect 69 177 79 211
rect 113 177 123 211
rect 69 159 123 177
rect 153 347 205 359
rect 153 313 163 347
rect 197 313 205 347
rect 153 159 205 313
rect -2215 -513 -2163 -501
rect -2215 -547 -2207 -513
rect -2173 -547 -2163 -513
rect -2215 -581 -2163 -547
rect -2215 -615 -2207 -581
rect -2173 -615 -2163 -581
rect -2215 -629 -2163 -615
rect -2133 -565 -2079 -501
rect -2133 -599 -2123 -565
rect -2089 -599 -2079 -565
rect -2133 -629 -2079 -599
rect -2049 -513 -1997 -501
rect -2049 -547 -2039 -513
rect -2005 -547 -1997 -513
rect -2049 -581 -1997 -547
rect -1026 -447 -972 -435
rect -1563 -521 -1476 -485
rect -1563 -551 -1520 -521
rect -2049 -615 -2039 -581
rect -2005 -615 -1997 -581
rect -2049 -629 -1997 -615
rect -1943 -589 -1891 -551
rect -1943 -623 -1935 -589
rect -1901 -623 -1891 -589
rect -1943 -635 -1891 -623
rect -1861 -581 -1806 -551
rect -1861 -615 -1851 -581
rect -1817 -615 -1806 -581
rect -1861 -635 -1806 -615
rect -1776 -576 -1711 -551
rect -1776 -610 -1759 -576
rect -1725 -610 -1711 -576
rect -1776 -635 -1711 -610
rect -1681 -635 -1608 -551
rect -1578 -555 -1520 -551
rect -1486 -555 -1476 -521
rect -1578 -589 -1476 -555
rect -1578 -623 -1520 -589
rect -1486 -623 -1476 -589
rect -1578 -635 -1476 -623
rect -1446 -551 -1396 -485
rect -1026 -481 -1018 -447
rect -984 -481 -972 -447
rect -1026 -518 -972 -481
rect -1446 -581 -1381 -551
rect -1446 -615 -1436 -581
rect -1402 -615 -1381 -581
rect -1446 -635 -1381 -615
rect -1351 -571 -1297 -551
rect -1351 -605 -1341 -571
rect -1307 -605 -1297 -571
rect -1351 -635 -1297 -605
rect -1267 -635 -1183 -551
rect -1153 -581 -1100 -551
rect -1153 -615 -1142 -581
rect -1108 -615 -1100 -581
rect -1153 -635 -1100 -615
rect -1026 -552 -1018 -518
rect -984 -552 -972 -518
rect -1026 -589 -972 -552
rect -1026 -623 -1018 -589
rect -984 -623 -972 -589
rect -1026 -635 -972 -623
rect -942 -479 -888 -435
rect -942 -513 -932 -479
rect -898 -513 -888 -479
rect -942 -559 -888 -513
rect -942 -593 -932 -559
rect -898 -593 -888 -559
rect -942 -635 -888 -593
rect -858 -447 -806 -435
rect -858 -481 -848 -447
rect -814 -481 -806 -447
rect -858 -515 -806 -481
rect -655 -453 -603 -435
rect -655 -487 -647 -453
rect -613 -487 -603 -453
rect -655 -507 -603 -487
rect -858 -549 -848 -515
rect -814 -549 -806 -515
rect -858 -583 -806 -549
rect -858 -617 -848 -583
rect -814 -617 -806 -583
rect -858 -635 -806 -617
rect -752 -521 -700 -507
rect -752 -555 -744 -521
rect -710 -555 -700 -521
rect -752 -589 -700 -555
rect -752 -623 -744 -589
rect -710 -623 -700 -589
rect -752 -635 -700 -623
rect -670 -521 -603 -507
rect -670 -555 -647 -521
rect -613 -555 -603 -521
rect -670 -589 -603 -555
rect -670 -623 -647 -589
rect -613 -623 -603 -589
rect -670 -635 -603 -623
rect -573 -447 -521 -435
rect -573 -481 -563 -447
rect -529 -481 -521 -447
rect -573 -518 -521 -481
rect -573 -552 -563 -518
rect -529 -552 -521 -518
rect -573 -589 -521 -552
rect -573 -623 -563 -589
rect -529 -623 -521 -589
rect -573 -635 -521 -623
rect -426 -453 -374 -435
rect -426 -487 -418 -453
rect -384 -487 -374 -453
rect -426 -521 -374 -487
rect -426 -555 -418 -521
rect -384 -555 -374 -521
rect -426 -589 -374 -555
rect -426 -623 -418 -589
rect -384 -623 -374 -589
rect -426 -635 -374 -623
rect -344 -453 -292 -435
rect -344 -487 -334 -453
rect -300 -487 -292 -453
rect -344 -521 -292 -487
rect -344 -555 -334 -521
rect -300 -555 -292 -521
rect -344 -589 -292 -555
rect -344 -623 -334 -589
rect -300 -623 -292 -589
rect -344 -635 -292 -623
rect -181 -453 -129 -435
rect -181 -487 -173 -453
rect -139 -487 -129 -453
rect -181 -521 -129 -487
rect -181 -555 -173 -521
rect -139 -555 -129 -521
rect -181 -589 -129 -555
rect -181 -623 -173 -589
rect -139 -623 -129 -589
rect -181 -635 -129 -623
rect -99 -453 -45 -435
rect -99 -487 -89 -453
rect -55 -487 -45 -453
rect -99 -521 -45 -487
rect -99 -555 -89 -521
rect -55 -555 -45 -521
rect -99 -589 -45 -555
rect -99 -623 -89 -589
rect -55 -623 -45 -589
rect -99 -635 -45 -623
rect -15 -521 39 -435
rect -15 -555 -5 -521
rect 29 -555 39 -521
rect -15 -589 39 -555
rect -15 -623 -5 -589
rect 29 -623 39 -589
rect -15 -635 39 -623
rect 69 -453 123 -435
rect 69 -487 79 -453
rect 113 -487 123 -453
rect 69 -521 123 -487
rect 69 -555 79 -521
rect 113 -555 123 -521
rect 69 -589 123 -555
rect 69 -623 79 -589
rect 113 -623 123 -589
rect 69 -635 123 -623
rect 153 -589 205 -435
rect 153 -623 163 -589
rect 197 -623 205 -589
rect 153 -635 205 -623
rect 483 -513 535 -501
rect 483 -547 491 -513
rect 525 -547 535 -513
rect 483 -581 535 -547
rect 483 -615 491 -581
rect 525 -615 535 -581
rect 483 -629 535 -615
rect 565 -565 619 -501
rect 565 -599 575 -565
rect 609 -599 619 -565
rect 565 -629 619 -599
rect 649 -513 701 -501
rect 649 -547 659 -513
rect 693 -547 701 -513
rect 649 -581 701 -547
rect 1672 -447 1726 -435
rect 1135 -521 1222 -485
rect 1135 -551 1178 -521
rect 649 -615 659 -581
rect 693 -615 701 -581
rect 649 -629 701 -615
rect 755 -589 807 -551
rect 755 -623 763 -589
rect 797 -623 807 -589
rect 755 -635 807 -623
rect 837 -581 892 -551
rect 837 -615 847 -581
rect 881 -615 892 -581
rect 837 -635 892 -615
rect 922 -576 987 -551
rect 922 -610 939 -576
rect 973 -610 987 -576
rect 922 -635 987 -610
rect 1017 -635 1090 -551
rect 1120 -555 1178 -551
rect 1212 -555 1222 -521
rect 1120 -589 1222 -555
rect 1120 -623 1178 -589
rect 1212 -623 1222 -589
rect 1120 -635 1222 -623
rect 1252 -551 1302 -485
rect 1672 -481 1680 -447
rect 1714 -481 1726 -447
rect 1672 -518 1726 -481
rect 1252 -581 1317 -551
rect 1252 -615 1262 -581
rect 1296 -615 1317 -581
rect 1252 -635 1317 -615
rect 1347 -571 1401 -551
rect 1347 -605 1357 -571
rect 1391 -605 1401 -571
rect 1347 -635 1401 -605
rect 1431 -635 1515 -551
rect 1545 -581 1598 -551
rect 1545 -615 1556 -581
rect 1590 -615 1598 -581
rect 1545 -635 1598 -615
rect 1672 -552 1680 -518
rect 1714 -552 1726 -518
rect 1672 -589 1726 -552
rect 1672 -623 1680 -589
rect 1714 -623 1726 -589
rect 1672 -635 1726 -623
rect 1756 -479 1810 -435
rect 1756 -513 1766 -479
rect 1800 -513 1810 -479
rect 1756 -559 1810 -513
rect 1756 -593 1766 -559
rect 1800 -593 1810 -559
rect 1756 -635 1810 -593
rect 1840 -447 1892 -435
rect 1840 -481 1850 -447
rect 1884 -481 1892 -447
rect 1840 -515 1892 -481
rect 2043 -453 2095 -435
rect 2043 -487 2051 -453
rect 2085 -487 2095 -453
rect 2043 -507 2095 -487
rect 1840 -549 1850 -515
rect 1884 -549 1892 -515
rect 1840 -583 1892 -549
rect 1840 -617 1850 -583
rect 1884 -617 1892 -583
rect 1840 -635 1892 -617
rect 1946 -521 1998 -507
rect 1946 -555 1954 -521
rect 1988 -555 1998 -521
rect 1946 -589 1998 -555
rect 1946 -623 1954 -589
rect 1988 -623 1998 -589
rect 1946 -635 1998 -623
rect 2028 -521 2095 -507
rect 2028 -555 2051 -521
rect 2085 -555 2095 -521
rect 2028 -589 2095 -555
rect 2028 -623 2051 -589
rect 2085 -623 2095 -589
rect 2028 -635 2095 -623
rect 2125 -447 2177 -435
rect 2125 -481 2135 -447
rect 2169 -481 2177 -447
rect 2125 -518 2177 -481
rect 2125 -552 2135 -518
rect 2169 -552 2177 -518
rect 2125 -589 2177 -552
rect 2125 -623 2135 -589
rect 2169 -623 2177 -589
rect 2125 -635 2177 -623
rect 2272 -453 2324 -435
rect 2272 -487 2280 -453
rect 2314 -487 2324 -453
rect 2272 -521 2324 -487
rect 2272 -555 2280 -521
rect 2314 -555 2324 -521
rect 2272 -589 2324 -555
rect 2272 -623 2280 -589
rect 2314 -623 2324 -589
rect 2272 -635 2324 -623
rect 2354 -453 2406 -435
rect 2354 -487 2364 -453
rect 2398 -487 2406 -453
rect 2354 -521 2406 -487
rect 2354 -555 2364 -521
rect 2398 -555 2406 -521
rect 2354 -589 2406 -555
rect 2354 -623 2364 -589
rect 2398 -623 2406 -589
rect 2354 -635 2406 -623
rect 2517 -453 2569 -435
rect 2517 -487 2525 -453
rect 2559 -487 2569 -453
rect 2517 -521 2569 -487
rect 2517 -555 2525 -521
rect 2559 -555 2569 -521
rect 2517 -589 2569 -555
rect 2517 -623 2525 -589
rect 2559 -623 2569 -589
rect 2517 -635 2569 -623
rect 2599 -453 2653 -435
rect 2599 -487 2609 -453
rect 2643 -487 2653 -453
rect 2599 -521 2653 -487
rect 2599 -555 2609 -521
rect 2643 -555 2653 -521
rect 2599 -589 2653 -555
rect 2599 -623 2609 -589
rect 2643 -623 2653 -589
rect 2599 -635 2653 -623
rect 2683 -521 2737 -435
rect 2683 -555 2693 -521
rect 2727 -555 2737 -521
rect 2683 -589 2737 -555
rect 2683 -623 2693 -589
rect 2727 -623 2737 -589
rect 2683 -635 2737 -623
rect 2767 -453 2821 -435
rect 2767 -487 2777 -453
rect 2811 -487 2821 -453
rect 2767 -521 2821 -487
rect 2767 -555 2777 -521
rect 2811 -555 2821 -521
rect 2767 -589 2821 -555
rect 2767 -623 2777 -589
rect 2811 -623 2821 -589
rect 2767 -635 2821 -623
rect 2851 -589 2903 -435
rect 2851 -623 2861 -589
rect 2895 -623 2903 -589
rect 2851 -635 2903 -623
rect -2215 -749 -2163 -735
rect -2215 -783 -2207 -749
rect -2173 -783 -2163 -749
rect -2215 -817 -2163 -783
rect -2215 -851 -2207 -817
rect -2173 -851 -2163 -817
rect -2215 -863 -2163 -851
rect -2133 -765 -2079 -735
rect -2133 -799 -2123 -765
rect -2089 -799 -2079 -765
rect -2133 -863 -2079 -799
rect -2049 -749 -1997 -735
rect -2049 -783 -2039 -749
rect -2005 -783 -1997 -749
rect -2049 -817 -1997 -783
rect -1943 -741 -1891 -729
rect -1943 -775 -1935 -741
rect -1901 -775 -1891 -741
rect -1943 -813 -1891 -775
rect -1861 -749 -1806 -729
rect -1861 -783 -1851 -749
rect -1817 -783 -1806 -749
rect -1861 -813 -1806 -783
rect -1776 -754 -1711 -729
rect -1776 -788 -1759 -754
rect -1725 -788 -1711 -754
rect -1776 -813 -1711 -788
rect -1681 -813 -1608 -729
rect -1578 -741 -1476 -729
rect -1578 -775 -1520 -741
rect -1486 -775 -1476 -741
rect -1578 -809 -1476 -775
rect -1578 -813 -1520 -809
rect -2049 -851 -2039 -817
rect -2005 -851 -1997 -817
rect -2049 -863 -1997 -851
rect -1563 -843 -1520 -813
rect -1486 -843 -1476 -809
rect -1563 -879 -1476 -843
rect -1446 -749 -1381 -729
rect -1446 -783 -1436 -749
rect -1402 -783 -1381 -749
rect -1446 -813 -1381 -783
rect -1351 -759 -1297 -729
rect -1351 -793 -1341 -759
rect -1307 -793 -1297 -759
rect -1351 -813 -1297 -793
rect -1267 -813 -1183 -729
rect -1153 -749 -1100 -729
rect -1153 -783 -1142 -749
rect -1108 -783 -1100 -749
rect -1153 -813 -1100 -783
rect -1026 -741 -972 -729
rect -1026 -775 -1018 -741
rect -984 -775 -972 -741
rect -1026 -812 -972 -775
rect -1446 -879 -1396 -813
rect -1026 -846 -1018 -812
rect -984 -846 -972 -812
rect -1026 -883 -972 -846
rect -1026 -917 -1018 -883
rect -984 -917 -972 -883
rect -1026 -929 -972 -917
rect -942 -771 -888 -729
rect -942 -805 -932 -771
rect -898 -805 -888 -771
rect -942 -851 -888 -805
rect -942 -885 -932 -851
rect -898 -885 -888 -851
rect -942 -929 -888 -885
rect -858 -747 -806 -729
rect -858 -781 -848 -747
rect -814 -781 -806 -747
rect -858 -815 -806 -781
rect -858 -849 -848 -815
rect -814 -849 -806 -815
rect -858 -883 -806 -849
rect -752 -741 -700 -729
rect -752 -775 -744 -741
rect -710 -775 -700 -741
rect -752 -809 -700 -775
rect -752 -843 -744 -809
rect -710 -843 -700 -809
rect -752 -857 -700 -843
rect -670 -741 -603 -729
rect -670 -775 -647 -741
rect -613 -775 -603 -741
rect -670 -809 -603 -775
rect -670 -843 -647 -809
rect -613 -843 -603 -809
rect -670 -857 -603 -843
rect -858 -917 -848 -883
rect -814 -917 -806 -883
rect -858 -929 -806 -917
rect -655 -877 -603 -857
rect -655 -911 -647 -877
rect -613 -911 -603 -877
rect -655 -929 -603 -911
rect -573 -741 -521 -729
rect -573 -775 -563 -741
rect -529 -775 -521 -741
rect -573 -812 -521 -775
rect -573 -846 -563 -812
rect -529 -846 -521 -812
rect -573 -883 -521 -846
rect -573 -917 -563 -883
rect -529 -917 -521 -883
rect -573 -929 -521 -917
rect -426 -741 -374 -729
rect -426 -775 -418 -741
rect -384 -775 -374 -741
rect -426 -809 -374 -775
rect -426 -843 -418 -809
rect -384 -843 -374 -809
rect -426 -877 -374 -843
rect -426 -911 -418 -877
rect -384 -911 -374 -877
rect -426 -929 -374 -911
rect -344 -741 -292 -729
rect -344 -775 -334 -741
rect -300 -775 -292 -741
rect -344 -809 -292 -775
rect -344 -843 -334 -809
rect -300 -843 -292 -809
rect -344 -877 -292 -843
rect -344 -911 -334 -877
rect -300 -911 -292 -877
rect -344 -929 -292 -911
rect -181 -741 -129 -729
rect -181 -775 -173 -741
rect -139 -775 -129 -741
rect -181 -809 -129 -775
rect -181 -843 -173 -809
rect -139 -843 -129 -809
rect -181 -877 -129 -843
rect -181 -911 -173 -877
rect -139 -911 -129 -877
rect -181 -929 -129 -911
rect -99 -741 -45 -729
rect -99 -775 -89 -741
rect -55 -775 -45 -741
rect -99 -809 -45 -775
rect -99 -843 -89 -809
rect -55 -843 -45 -809
rect -99 -877 -45 -843
rect -99 -911 -89 -877
rect -55 -911 -45 -877
rect -99 -929 -45 -911
rect -15 -741 39 -729
rect -15 -775 -5 -741
rect 29 -775 39 -741
rect -15 -809 39 -775
rect -15 -843 -5 -809
rect 29 -843 39 -809
rect -15 -929 39 -843
rect 69 -741 123 -729
rect 69 -775 79 -741
rect 113 -775 123 -741
rect 69 -809 123 -775
rect 69 -843 79 -809
rect 113 -843 123 -809
rect 69 -877 123 -843
rect 69 -911 79 -877
rect 113 -911 123 -877
rect 69 -929 123 -911
rect 153 -741 205 -729
rect 153 -775 163 -741
rect 197 -775 205 -741
rect 153 -929 205 -775
rect 483 -749 535 -735
rect 483 -783 491 -749
rect 525 -783 535 -749
rect 483 -817 535 -783
rect 483 -851 491 -817
rect 525 -851 535 -817
rect 483 -863 535 -851
rect 565 -765 619 -735
rect 565 -799 575 -765
rect 609 -799 619 -765
rect 565 -863 619 -799
rect 649 -749 701 -735
rect 649 -783 659 -749
rect 693 -783 701 -749
rect 649 -817 701 -783
rect 755 -741 807 -729
rect 755 -775 763 -741
rect 797 -775 807 -741
rect 755 -813 807 -775
rect 837 -749 892 -729
rect 837 -783 847 -749
rect 881 -783 892 -749
rect 837 -813 892 -783
rect 922 -754 987 -729
rect 922 -788 939 -754
rect 973 -788 987 -754
rect 922 -813 987 -788
rect 1017 -813 1090 -729
rect 1120 -741 1222 -729
rect 1120 -775 1178 -741
rect 1212 -775 1222 -741
rect 1120 -809 1222 -775
rect 1120 -813 1178 -809
rect 649 -851 659 -817
rect 693 -851 701 -817
rect 649 -863 701 -851
rect 1135 -843 1178 -813
rect 1212 -843 1222 -809
rect 1135 -879 1222 -843
rect 1252 -749 1317 -729
rect 1252 -783 1262 -749
rect 1296 -783 1317 -749
rect 1252 -813 1317 -783
rect 1347 -759 1401 -729
rect 1347 -793 1357 -759
rect 1391 -793 1401 -759
rect 1347 -813 1401 -793
rect 1431 -813 1515 -729
rect 1545 -749 1598 -729
rect 1545 -783 1556 -749
rect 1590 -783 1598 -749
rect 1545 -813 1598 -783
rect 1672 -741 1726 -729
rect 1672 -775 1680 -741
rect 1714 -775 1726 -741
rect 1672 -812 1726 -775
rect 1252 -879 1302 -813
rect 1672 -846 1680 -812
rect 1714 -846 1726 -812
rect 1672 -883 1726 -846
rect 1672 -917 1680 -883
rect 1714 -917 1726 -883
rect 1672 -929 1726 -917
rect 1756 -771 1810 -729
rect 1756 -805 1766 -771
rect 1800 -805 1810 -771
rect 1756 -851 1810 -805
rect 1756 -885 1766 -851
rect 1800 -885 1810 -851
rect 1756 -929 1810 -885
rect 1840 -747 1892 -729
rect 1840 -781 1850 -747
rect 1884 -781 1892 -747
rect 1840 -815 1892 -781
rect 1840 -849 1850 -815
rect 1884 -849 1892 -815
rect 1840 -883 1892 -849
rect 1946 -741 1998 -729
rect 1946 -775 1954 -741
rect 1988 -775 1998 -741
rect 1946 -809 1998 -775
rect 1946 -843 1954 -809
rect 1988 -843 1998 -809
rect 1946 -857 1998 -843
rect 2028 -741 2095 -729
rect 2028 -775 2051 -741
rect 2085 -775 2095 -741
rect 2028 -809 2095 -775
rect 2028 -843 2051 -809
rect 2085 -843 2095 -809
rect 2028 -857 2095 -843
rect 1840 -917 1850 -883
rect 1884 -917 1892 -883
rect 1840 -929 1892 -917
rect 2043 -877 2095 -857
rect 2043 -911 2051 -877
rect 2085 -911 2095 -877
rect 2043 -929 2095 -911
rect 2125 -741 2177 -729
rect 2125 -775 2135 -741
rect 2169 -775 2177 -741
rect 2125 -812 2177 -775
rect 2125 -846 2135 -812
rect 2169 -846 2177 -812
rect 2125 -883 2177 -846
rect 2125 -917 2135 -883
rect 2169 -917 2177 -883
rect 2125 -929 2177 -917
rect 2272 -741 2324 -729
rect 2272 -775 2280 -741
rect 2314 -775 2324 -741
rect 2272 -809 2324 -775
rect 2272 -843 2280 -809
rect 2314 -843 2324 -809
rect 2272 -877 2324 -843
rect 2272 -911 2280 -877
rect 2314 -911 2324 -877
rect 2272 -929 2324 -911
rect 2354 -741 2406 -729
rect 2354 -775 2364 -741
rect 2398 -775 2406 -741
rect 2354 -809 2406 -775
rect 2354 -843 2364 -809
rect 2398 -843 2406 -809
rect 2354 -877 2406 -843
rect 2354 -911 2364 -877
rect 2398 -911 2406 -877
rect 2354 -929 2406 -911
rect 2517 -741 2569 -729
rect 2517 -775 2525 -741
rect 2559 -775 2569 -741
rect 2517 -809 2569 -775
rect 2517 -843 2525 -809
rect 2559 -843 2569 -809
rect 2517 -877 2569 -843
rect 2517 -911 2525 -877
rect 2559 -911 2569 -877
rect 2517 -929 2569 -911
rect 2599 -741 2653 -729
rect 2599 -775 2609 -741
rect 2643 -775 2653 -741
rect 2599 -809 2653 -775
rect 2599 -843 2609 -809
rect 2643 -843 2653 -809
rect 2599 -877 2653 -843
rect 2599 -911 2609 -877
rect 2643 -911 2653 -877
rect 2599 -929 2653 -911
rect 2683 -741 2737 -729
rect 2683 -775 2693 -741
rect 2727 -775 2737 -741
rect 2683 -809 2737 -775
rect 2683 -843 2693 -809
rect 2727 -843 2737 -809
rect 2683 -929 2737 -843
rect 2767 -741 2821 -729
rect 2767 -775 2777 -741
rect 2811 -775 2821 -741
rect 2767 -809 2821 -775
rect 2767 -843 2777 -809
rect 2811 -843 2821 -809
rect 2767 -877 2821 -843
rect 2767 -911 2777 -877
rect 2811 -911 2821 -877
rect 2767 -929 2821 -911
rect 2851 -741 2903 -729
rect 2851 -775 2861 -741
rect 2895 -775 2903 -741
rect 2851 -929 2903 -775
rect -2215 -1601 -2163 -1589
rect -2215 -1635 -2207 -1601
rect -2173 -1635 -2163 -1601
rect -2215 -1669 -2163 -1635
rect -2215 -1703 -2207 -1669
rect -2173 -1703 -2163 -1669
rect -2215 -1717 -2163 -1703
rect -2133 -1653 -2079 -1589
rect -2133 -1687 -2123 -1653
rect -2089 -1687 -2079 -1653
rect -2133 -1717 -2079 -1687
rect -2049 -1601 -1997 -1589
rect -2049 -1635 -2039 -1601
rect -2005 -1635 -1997 -1601
rect -2049 -1669 -1997 -1635
rect -1026 -1535 -972 -1523
rect -1563 -1609 -1476 -1573
rect -1563 -1639 -1520 -1609
rect -2049 -1703 -2039 -1669
rect -2005 -1703 -1997 -1669
rect -2049 -1717 -1997 -1703
rect -1943 -1677 -1891 -1639
rect -1943 -1711 -1935 -1677
rect -1901 -1711 -1891 -1677
rect -1943 -1723 -1891 -1711
rect -1861 -1669 -1806 -1639
rect -1861 -1703 -1851 -1669
rect -1817 -1703 -1806 -1669
rect -1861 -1723 -1806 -1703
rect -1776 -1664 -1711 -1639
rect -1776 -1698 -1759 -1664
rect -1725 -1698 -1711 -1664
rect -1776 -1723 -1711 -1698
rect -1681 -1723 -1608 -1639
rect -1578 -1643 -1520 -1639
rect -1486 -1643 -1476 -1609
rect -1578 -1677 -1476 -1643
rect -1578 -1711 -1520 -1677
rect -1486 -1711 -1476 -1677
rect -1578 -1723 -1476 -1711
rect -1446 -1639 -1396 -1573
rect -1026 -1569 -1018 -1535
rect -984 -1569 -972 -1535
rect -1026 -1606 -972 -1569
rect -1446 -1669 -1381 -1639
rect -1446 -1703 -1436 -1669
rect -1402 -1703 -1381 -1669
rect -1446 -1723 -1381 -1703
rect -1351 -1659 -1297 -1639
rect -1351 -1693 -1341 -1659
rect -1307 -1693 -1297 -1659
rect -1351 -1723 -1297 -1693
rect -1267 -1723 -1183 -1639
rect -1153 -1669 -1100 -1639
rect -1153 -1703 -1142 -1669
rect -1108 -1703 -1100 -1669
rect -1153 -1723 -1100 -1703
rect -1026 -1640 -1018 -1606
rect -984 -1640 -972 -1606
rect -1026 -1677 -972 -1640
rect -1026 -1711 -1018 -1677
rect -984 -1711 -972 -1677
rect -1026 -1723 -972 -1711
rect -942 -1567 -888 -1523
rect -942 -1601 -932 -1567
rect -898 -1601 -888 -1567
rect -942 -1647 -888 -1601
rect -942 -1681 -932 -1647
rect -898 -1681 -888 -1647
rect -942 -1723 -888 -1681
rect -858 -1535 -806 -1523
rect -858 -1569 -848 -1535
rect -814 -1569 -806 -1535
rect -858 -1603 -806 -1569
rect -655 -1541 -603 -1523
rect -655 -1575 -647 -1541
rect -613 -1575 -603 -1541
rect -655 -1595 -603 -1575
rect -858 -1637 -848 -1603
rect -814 -1637 -806 -1603
rect -858 -1671 -806 -1637
rect -858 -1705 -848 -1671
rect -814 -1705 -806 -1671
rect -858 -1723 -806 -1705
rect -752 -1609 -700 -1595
rect -752 -1643 -744 -1609
rect -710 -1643 -700 -1609
rect -752 -1677 -700 -1643
rect -752 -1711 -744 -1677
rect -710 -1711 -700 -1677
rect -752 -1723 -700 -1711
rect -670 -1609 -603 -1595
rect -670 -1643 -647 -1609
rect -613 -1643 -603 -1609
rect -670 -1677 -603 -1643
rect -670 -1711 -647 -1677
rect -613 -1711 -603 -1677
rect -670 -1723 -603 -1711
rect -573 -1535 -521 -1523
rect -573 -1569 -563 -1535
rect -529 -1569 -521 -1535
rect -573 -1606 -521 -1569
rect -573 -1640 -563 -1606
rect -529 -1640 -521 -1606
rect -573 -1677 -521 -1640
rect -573 -1711 -563 -1677
rect -529 -1711 -521 -1677
rect -573 -1723 -521 -1711
rect -426 -1541 -374 -1523
rect -426 -1575 -418 -1541
rect -384 -1575 -374 -1541
rect -426 -1609 -374 -1575
rect -426 -1643 -418 -1609
rect -384 -1643 -374 -1609
rect -426 -1677 -374 -1643
rect -426 -1711 -418 -1677
rect -384 -1711 -374 -1677
rect -426 -1723 -374 -1711
rect -344 -1541 -292 -1523
rect -344 -1575 -334 -1541
rect -300 -1575 -292 -1541
rect -344 -1609 -292 -1575
rect -344 -1643 -334 -1609
rect -300 -1643 -292 -1609
rect -344 -1677 -292 -1643
rect -344 -1711 -334 -1677
rect -300 -1711 -292 -1677
rect -344 -1723 -292 -1711
rect -181 -1541 -129 -1523
rect -181 -1575 -173 -1541
rect -139 -1575 -129 -1541
rect -181 -1609 -129 -1575
rect -181 -1643 -173 -1609
rect -139 -1643 -129 -1609
rect -181 -1677 -129 -1643
rect -181 -1711 -173 -1677
rect -139 -1711 -129 -1677
rect -181 -1723 -129 -1711
rect -99 -1541 -45 -1523
rect -99 -1575 -89 -1541
rect -55 -1575 -45 -1541
rect -99 -1609 -45 -1575
rect -99 -1643 -89 -1609
rect -55 -1643 -45 -1609
rect -99 -1677 -45 -1643
rect -99 -1711 -89 -1677
rect -55 -1711 -45 -1677
rect -99 -1723 -45 -1711
rect -15 -1609 39 -1523
rect -15 -1643 -5 -1609
rect 29 -1643 39 -1609
rect -15 -1677 39 -1643
rect -15 -1711 -5 -1677
rect 29 -1711 39 -1677
rect -15 -1723 39 -1711
rect 69 -1541 123 -1523
rect 69 -1575 79 -1541
rect 113 -1575 123 -1541
rect 69 -1609 123 -1575
rect 69 -1643 79 -1609
rect 113 -1643 123 -1609
rect 69 -1677 123 -1643
rect 69 -1711 79 -1677
rect 113 -1711 123 -1677
rect 69 -1723 123 -1711
rect 153 -1677 205 -1523
rect 153 -1711 163 -1677
rect 197 -1711 205 -1677
rect 153 -1723 205 -1711
rect 483 -1601 535 -1589
rect 483 -1635 491 -1601
rect 525 -1635 535 -1601
rect 483 -1669 535 -1635
rect 483 -1703 491 -1669
rect 525 -1703 535 -1669
rect 483 -1717 535 -1703
rect 565 -1653 619 -1589
rect 565 -1687 575 -1653
rect 609 -1687 619 -1653
rect 565 -1717 619 -1687
rect 649 -1601 701 -1589
rect 649 -1635 659 -1601
rect 693 -1635 701 -1601
rect 649 -1669 701 -1635
rect 1672 -1535 1726 -1523
rect 1135 -1609 1222 -1573
rect 1135 -1639 1178 -1609
rect 649 -1703 659 -1669
rect 693 -1703 701 -1669
rect 649 -1717 701 -1703
rect 755 -1677 807 -1639
rect 755 -1711 763 -1677
rect 797 -1711 807 -1677
rect 755 -1723 807 -1711
rect 837 -1669 892 -1639
rect 837 -1703 847 -1669
rect 881 -1703 892 -1669
rect 837 -1723 892 -1703
rect 922 -1664 987 -1639
rect 922 -1698 939 -1664
rect 973 -1698 987 -1664
rect 922 -1723 987 -1698
rect 1017 -1723 1090 -1639
rect 1120 -1643 1178 -1639
rect 1212 -1643 1222 -1609
rect 1120 -1677 1222 -1643
rect 1120 -1711 1178 -1677
rect 1212 -1711 1222 -1677
rect 1120 -1723 1222 -1711
rect 1252 -1639 1302 -1573
rect 1672 -1569 1680 -1535
rect 1714 -1569 1726 -1535
rect 1672 -1606 1726 -1569
rect 1252 -1669 1317 -1639
rect 1252 -1703 1262 -1669
rect 1296 -1703 1317 -1669
rect 1252 -1723 1317 -1703
rect 1347 -1659 1401 -1639
rect 1347 -1693 1357 -1659
rect 1391 -1693 1401 -1659
rect 1347 -1723 1401 -1693
rect 1431 -1723 1515 -1639
rect 1545 -1669 1598 -1639
rect 1545 -1703 1556 -1669
rect 1590 -1703 1598 -1669
rect 1545 -1723 1598 -1703
rect 1672 -1640 1680 -1606
rect 1714 -1640 1726 -1606
rect 1672 -1677 1726 -1640
rect 1672 -1711 1680 -1677
rect 1714 -1711 1726 -1677
rect 1672 -1723 1726 -1711
rect 1756 -1567 1810 -1523
rect 1756 -1601 1766 -1567
rect 1800 -1601 1810 -1567
rect 1756 -1647 1810 -1601
rect 1756 -1681 1766 -1647
rect 1800 -1681 1810 -1647
rect 1756 -1723 1810 -1681
rect 1840 -1535 1892 -1523
rect 1840 -1569 1850 -1535
rect 1884 -1569 1892 -1535
rect 1840 -1603 1892 -1569
rect 2043 -1541 2095 -1523
rect 2043 -1575 2051 -1541
rect 2085 -1575 2095 -1541
rect 2043 -1595 2095 -1575
rect 1840 -1637 1850 -1603
rect 1884 -1637 1892 -1603
rect 1840 -1671 1892 -1637
rect 1840 -1705 1850 -1671
rect 1884 -1705 1892 -1671
rect 1840 -1723 1892 -1705
rect 1946 -1609 1998 -1595
rect 1946 -1643 1954 -1609
rect 1988 -1643 1998 -1609
rect 1946 -1677 1998 -1643
rect 1946 -1711 1954 -1677
rect 1988 -1711 1998 -1677
rect 1946 -1723 1998 -1711
rect 2028 -1609 2095 -1595
rect 2028 -1643 2051 -1609
rect 2085 -1643 2095 -1609
rect 2028 -1677 2095 -1643
rect 2028 -1711 2051 -1677
rect 2085 -1711 2095 -1677
rect 2028 -1723 2095 -1711
rect 2125 -1535 2177 -1523
rect 2125 -1569 2135 -1535
rect 2169 -1569 2177 -1535
rect 2125 -1606 2177 -1569
rect 2125 -1640 2135 -1606
rect 2169 -1640 2177 -1606
rect 2125 -1677 2177 -1640
rect 2125 -1711 2135 -1677
rect 2169 -1711 2177 -1677
rect 2125 -1723 2177 -1711
rect 2272 -1541 2324 -1523
rect 2272 -1575 2280 -1541
rect 2314 -1575 2324 -1541
rect 2272 -1609 2324 -1575
rect 2272 -1643 2280 -1609
rect 2314 -1643 2324 -1609
rect 2272 -1677 2324 -1643
rect 2272 -1711 2280 -1677
rect 2314 -1711 2324 -1677
rect 2272 -1723 2324 -1711
rect 2354 -1541 2406 -1523
rect 2354 -1575 2364 -1541
rect 2398 -1575 2406 -1541
rect 2354 -1609 2406 -1575
rect 2354 -1643 2364 -1609
rect 2398 -1643 2406 -1609
rect 2354 -1677 2406 -1643
rect 2354 -1711 2364 -1677
rect 2398 -1711 2406 -1677
rect 2354 -1723 2406 -1711
rect 2517 -1541 2569 -1523
rect 2517 -1575 2525 -1541
rect 2559 -1575 2569 -1541
rect 2517 -1609 2569 -1575
rect 2517 -1643 2525 -1609
rect 2559 -1643 2569 -1609
rect 2517 -1677 2569 -1643
rect 2517 -1711 2525 -1677
rect 2559 -1711 2569 -1677
rect 2517 -1723 2569 -1711
rect 2599 -1541 2653 -1523
rect 2599 -1575 2609 -1541
rect 2643 -1575 2653 -1541
rect 2599 -1609 2653 -1575
rect 2599 -1643 2609 -1609
rect 2643 -1643 2653 -1609
rect 2599 -1677 2653 -1643
rect 2599 -1711 2609 -1677
rect 2643 -1711 2653 -1677
rect 2599 -1723 2653 -1711
rect 2683 -1609 2737 -1523
rect 2683 -1643 2693 -1609
rect 2727 -1643 2737 -1609
rect 2683 -1677 2737 -1643
rect 2683 -1711 2693 -1677
rect 2727 -1711 2737 -1677
rect 2683 -1723 2737 -1711
rect 2767 -1541 2821 -1523
rect 2767 -1575 2777 -1541
rect 2811 -1575 2821 -1541
rect 2767 -1609 2821 -1575
rect 2767 -1643 2777 -1609
rect 2811 -1643 2821 -1609
rect 2767 -1677 2821 -1643
rect 2767 -1711 2777 -1677
rect 2811 -1711 2821 -1677
rect 2767 -1723 2821 -1711
rect 2851 -1677 2903 -1523
rect 2851 -1711 2861 -1677
rect 2895 -1711 2903 -1677
rect 2851 -1723 2903 -1711
rect -2215 -1837 -2163 -1823
rect -2215 -1871 -2207 -1837
rect -2173 -1871 -2163 -1837
rect -2215 -1905 -2163 -1871
rect -2215 -1939 -2207 -1905
rect -2173 -1939 -2163 -1905
rect -2215 -1951 -2163 -1939
rect -2133 -1853 -2079 -1823
rect -2133 -1887 -2123 -1853
rect -2089 -1887 -2079 -1853
rect -2133 -1951 -2079 -1887
rect -2049 -1837 -1997 -1823
rect -2049 -1871 -2039 -1837
rect -2005 -1871 -1997 -1837
rect -2049 -1905 -1997 -1871
rect -1943 -1829 -1891 -1817
rect -1943 -1863 -1935 -1829
rect -1901 -1863 -1891 -1829
rect -1943 -1901 -1891 -1863
rect -1861 -1837 -1806 -1817
rect -1861 -1871 -1851 -1837
rect -1817 -1871 -1806 -1837
rect -1861 -1901 -1806 -1871
rect -1776 -1842 -1711 -1817
rect -1776 -1876 -1759 -1842
rect -1725 -1876 -1711 -1842
rect -1776 -1901 -1711 -1876
rect -1681 -1901 -1608 -1817
rect -1578 -1829 -1476 -1817
rect -1578 -1863 -1520 -1829
rect -1486 -1863 -1476 -1829
rect -1578 -1897 -1476 -1863
rect -1578 -1901 -1520 -1897
rect -2049 -1939 -2039 -1905
rect -2005 -1939 -1997 -1905
rect -2049 -1951 -1997 -1939
rect -1563 -1931 -1520 -1901
rect -1486 -1931 -1476 -1897
rect -1563 -1967 -1476 -1931
rect -1446 -1837 -1381 -1817
rect -1446 -1871 -1436 -1837
rect -1402 -1871 -1381 -1837
rect -1446 -1901 -1381 -1871
rect -1351 -1847 -1297 -1817
rect -1351 -1881 -1341 -1847
rect -1307 -1881 -1297 -1847
rect -1351 -1901 -1297 -1881
rect -1267 -1901 -1183 -1817
rect -1153 -1837 -1100 -1817
rect -1153 -1871 -1142 -1837
rect -1108 -1871 -1100 -1837
rect -1153 -1901 -1100 -1871
rect -1026 -1829 -972 -1817
rect -1026 -1863 -1018 -1829
rect -984 -1863 -972 -1829
rect -1026 -1900 -972 -1863
rect -1446 -1967 -1396 -1901
rect -1026 -1934 -1018 -1900
rect -984 -1934 -972 -1900
rect -1026 -1971 -972 -1934
rect -1026 -2005 -1018 -1971
rect -984 -2005 -972 -1971
rect -1026 -2017 -972 -2005
rect -942 -1859 -888 -1817
rect -942 -1893 -932 -1859
rect -898 -1893 -888 -1859
rect -942 -1939 -888 -1893
rect -942 -1973 -932 -1939
rect -898 -1973 -888 -1939
rect -942 -2017 -888 -1973
rect -858 -1835 -806 -1817
rect -858 -1869 -848 -1835
rect -814 -1869 -806 -1835
rect -858 -1903 -806 -1869
rect -858 -1937 -848 -1903
rect -814 -1937 -806 -1903
rect -858 -1971 -806 -1937
rect -752 -1829 -700 -1817
rect -752 -1863 -744 -1829
rect -710 -1863 -700 -1829
rect -752 -1897 -700 -1863
rect -752 -1931 -744 -1897
rect -710 -1931 -700 -1897
rect -752 -1945 -700 -1931
rect -670 -1829 -603 -1817
rect -670 -1863 -647 -1829
rect -613 -1863 -603 -1829
rect -670 -1897 -603 -1863
rect -670 -1931 -647 -1897
rect -613 -1931 -603 -1897
rect -670 -1945 -603 -1931
rect -858 -2005 -848 -1971
rect -814 -2005 -806 -1971
rect -858 -2017 -806 -2005
rect -655 -1965 -603 -1945
rect -655 -1999 -647 -1965
rect -613 -1999 -603 -1965
rect -655 -2017 -603 -1999
rect -573 -1829 -521 -1817
rect -573 -1863 -563 -1829
rect -529 -1863 -521 -1829
rect -573 -1900 -521 -1863
rect -573 -1934 -563 -1900
rect -529 -1934 -521 -1900
rect -573 -1971 -521 -1934
rect -573 -2005 -563 -1971
rect -529 -2005 -521 -1971
rect -573 -2017 -521 -2005
rect -426 -1829 -374 -1817
rect -426 -1863 -418 -1829
rect -384 -1863 -374 -1829
rect -426 -1897 -374 -1863
rect -426 -1931 -418 -1897
rect -384 -1931 -374 -1897
rect -426 -1965 -374 -1931
rect -426 -1999 -418 -1965
rect -384 -1999 -374 -1965
rect -426 -2017 -374 -1999
rect -344 -1829 -292 -1817
rect -344 -1863 -334 -1829
rect -300 -1863 -292 -1829
rect -344 -1897 -292 -1863
rect -344 -1931 -334 -1897
rect -300 -1931 -292 -1897
rect -344 -1965 -292 -1931
rect -344 -1999 -334 -1965
rect -300 -1999 -292 -1965
rect -344 -2017 -292 -1999
rect -181 -1829 -129 -1817
rect -181 -1863 -173 -1829
rect -139 -1863 -129 -1829
rect -181 -1897 -129 -1863
rect -181 -1931 -173 -1897
rect -139 -1931 -129 -1897
rect -181 -1965 -129 -1931
rect -181 -1999 -173 -1965
rect -139 -1999 -129 -1965
rect -181 -2017 -129 -1999
rect -99 -1829 -45 -1817
rect -99 -1863 -89 -1829
rect -55 -1863 -45 -1829
rect -99 -1897 -45 -1863
rect -99 -1931 -89 -1897
rect -55 -1931 -45 -1897
rect -99 -1965 -45 -1931
rect -99 -1999 -89 -1965
rect -55 -1999 -45 -1965
rect -99 -2017 -45 -1999
rect -15 -1829 39 -1817
rect -15 -1863 -5 -1829
rect 29 -1863 39 -1829
rect -15 -1897 39 -1863
rect -15 -1931 -5 -1897
rect 29 -1931 39 -1897
rect -15 -2017 39 -1931
rect 69 -1829 123 -1817
rect 69 -1863 79 -1829
rect 113 -1863 123 -1829
rect 69 -1897 123 -1863
rect 69 -1931 79 -1897
rect 113 -1931 123 -1897
rect 69 -1965 123 -1931
rect 69 -1999 79 -1965
rect 113 -1999 123 -1965
rect 69 -2017 123 -1999
rect 153 -1829 205 -1817
rect 153 -1863 163 -1829
rect 197 -1863 205 -1829
rect 153 -2017 205 -1863
rect 483 -1837 535 -1823
rect 483 -1871 491 -1837
rect 525 -1871 535 -1837
rect 483 -1905 535 -1871
rect 483 -1939 491 -1905
rect 525 -1939 535 -1905
rect 483 -1951 535 -1939
rect 565 -1853 619 -1823
rect 565 -1887 575 -1853
rect 609 -1887 619 -1853
rect 565 -1951 619 -1887
rect 649 -1837 701 -1823
rect 649 -1871 659 -1837
rect 693 -1871 701 -1837
rect 649 -1905 701 -1871
rect 755 -1829 807 -1817
rect 755 -1863 763 -1829
rect 797 -1863 807 -1829
rect 755 -1901 807 -1863
rect 837 -1837 892 -1817
rect 837 -1871 847 -1837
rect 881 -1871 892 -1837
rect 837 -1901 892 -1871
rect 922 -1842 987 -1817
rect 922 -1876 939 -1842
rect 973 -1876 987 -1842
rect 922 -1901 987 -1876
rect 1017 -1901 1090 -1817
rect 1120 -1829 1222 -1817
rect 1120 -1863 1178 -1829
rect 1212 -1863 1222 -1829
rect 1120 -1897 1222 -1863
rect 1120 -1901 1178 -1897
rect 649 -1939 659 -1905
rect 693 -1939 701 -1905
rect 649 -1951 701 -1939
rect 1135 -1931 1178 -1901
rect 1212 -1931 1222 -1897
rect 1135 -1967 1222 -1931
rect 1252 -1837 1317 -1817
rect 1252 -1871 1262 -1837
rect 1296 -1871 1317 -1837
rect 1252 -1901 1317 -1871
rect 1347 -1847 1401 -1817
rect 1347 -1881 1357 -1847
rect 1391 -1881 1401 -1847
rect 1347 -1901 1401 -1881
rect 1431 -1901 1515 -1817
rect 1545 -1837 1598 -1817
rect 1545 -1871 1556 -1837
rect 1590 -1871 1598 -1837
rect 1545 -1901 1598 -1871
rect 1672 -1829 1726 -1817
rect 1672 -1863 1680 -1829
rect 1714 -1863 1726 -1829
rect 1672 -1900 1726 -1863
rect 1252 -1967 1302 -1901
rect 1672 -1934 1680 -1900
rect 1714 -1934 1726 -1900
rect 1672 -1971 1726 -1934
rect 1672 -2005 1680 -1971
rect 1714 -2005 1726 -1971
rect 1672 -2017 1726 -2005
rect 1756 -1859 1810 -1817
rect 1756 -1893 1766 -1859
rect 1800 -1893 1810 -1859
rect 1756 -1939 1810 -1893
rect 1756 -1973 1766 -1939
rect 1800 -1973 1810 -1939
rect 1756 -2017 1810 -1973
rect 1840 -1835 1892 -1817
rect 1840 -1869 1850 -1835
rect 1884 -1869 1892 -1835
rect 1840 -1903 1892 -1869
rect 1840 -1937 1850 -1903
rect 1884 -1937 1892 -1903
rect 1840 -1971 1892 -1937
rect 1946 -1829 1998 -1817
rect 1946 -1863 1954 -1829
rect 1988 -1863 1998 -1829
rect 1946 -1897 1998 -1863
rect 1946 -1931 1954 -1897
rect 1988 -1931 1998 -1897
rect 1946 -1945 1998 -1931
rect 2028 -1829 2095 -1817
rect 2028 -1863 2051 -1829
rect 2085 -1863 2095 -1829
rect 2028 -1897 2095 -1863
rect 2028 -1931 2051 -1897
rect 2085 -1931 2095 -1897
rect 2028 -1945 2095 -1931
rect 1840 -2005 1850 -1971
rect 1884 -2005 1892 -1971
rect 1840 -2017 1892 -2005
rect 2043 -1965 2095 -1945
rect 2043 -1999 2051 -1965
rect 2085 -1999 2095 -1965
rect 2043 -2017 2095 -1999
rect 2125 -1829 2177 -1817
rect 2125 -1863 2135 -1829
rect 2169 -1863 2177 -1829
rect 2125 -1900 2177 -1863
rect 2125 -1934 2135 -1900
rect 2169 -1934 2177 -1900
rect 2125 -1971 2177 -1934
rect 2125 -2005 2135 -1971
rect 2169 -2005 2177 -1971
rect 2125 -2017 2177 -2005
rect 2272 -1829 2324 -1817
rect 2272 -1863 2280 -1829
rect 2314 -1863 2324 -1829
rect 2272 -1897 2324 -1863
rect 2272 -1931 2280 -1897
rect 2314 -1931 2324 -1897
rect 2272 -1965 2324 -1931
rect 2272 -1999 2280 -1965
rect 2314 -1999 2324 -1965
rect 2272 -2017 2324 -1999
rect 2354 -1829 2406 -1817
rect 2354 -1863 2364 -1829
rect 2398 -1863 2406 -1829
rect 2354 -1897 2406 -1863
rect 2354 -1931 2364 -1897
rect 2398 -1931 2406 -1897
rect 2354 -1965 2406 -1931
rect 2354 -1999 2364 -1965
rect 2398 -1999 2406 -1965
rect 2354 -2017 2406 -1999
rect 2517 -1829 2569 -1817
rect 2517 -1863 2525 -1829
rect 2559 -1863 2569 -1829
rect 2517 -1897 2569 -1863
rect 2517 -1931 2525 -1897
rect 2559 -1931 2569 -1897
rect 2517 -1965 2569 -1931
rect 2517 -1999 2525 -1965
rect 2559 -1999 2569 -1965
rect 2517 -2017 2569 -1999
rect 2599 -1829 2653 -1817
rect 2599 -1863 2609 -1829
rect 2643 -1863 2653 -1829
rect 2599 -1897 2653 -1863
rect 2599 -1931 2609 -1897
rect 2643 -1931 2653 -1897
rect 2599 -1965 2653 -1931
rect 2599 -1999 2609 -1965
rect 2643 -1999 2653 -1965
rect 2599 -2017 2653 -1999
rect 2683 -1829 2737 -1817
rect 2683 -1863 2693 -1829
rect 2727 -1863 2737 -1829
rect 2683 -1897 2737 -1863
rect 2683 -1931 2693 -1897
rect 2727 -1931 2737 -1897
rect 2683 -2017 2737 -1931
rect 2767 -1829 2821 -1817
rect 2767 -1863 2777 -1829
rect 2811 -1863 2821 -1829
rect 2767 -1897 2821 -1863
rect 2767 -1931 2777 -1897
rect 2811 -1931 2821 -1897
rect 2767 -1965 2821 -1931
rect 2767 -1999 2777 -1965
rect 2811 -1999 2821 -1965
rect 2767 -2017 2821 -1999
rect 2851 -1829 2903 -1817
rect 2851 -1863 2861 -1829
rect 2895 -1863 2903 -1829
rect 2851 -2017 2903 -1863
rect -2215 -2689 -2163 -2677
rect -2215 -2723 -2207 -2689
rect -2173 -2723 -2163 -2689
rect -2215 -2757 -2163 -2723
rect -2215 -2791 -2207 -2757
rect -2173 -2791 -2163 -2757
rect -2215 -2805 -2163 -2791
rect -2133 -2741 -2079 -2677
rect -2133 -2775 -2123 -2741
rect -2089 -2775 -2079 -2741
rect -2133 -2805 -2079 -2775
rect -2049 -2689 -1997 -2677
rect -2049 -2723 -2039 -2689
rect -2005 -2723 -1997 -2689
rect -2049 -2757 -1997 -2723
rect -1026 -2623 -972 -2611
rect -1563 -2697 -1476 -2661
rect -1563 -2727 -1520 -2697
rect -2049 -2791 -2039 -2757
rect -2005 -2791 -1997 -2757
rect -2049 -2805 -1997 -2791
rect -1943 -2765 -1891 -2727
rect -1943 -2799 -1935 -2765
rect -1901 -2799 -1891 -2765
rect -1943 -2811 -1891 -2799
rect -1861 -2757 -1806 -2727
rect -1861 -2791 -1851 -2757
rect -1817 -2791 -1806 -2757
rect -1861 -2811 -1806 -2791
rect -1776 -2752 -1711 -2727
rect -1776 -2786 -1759 -2752
rect -1725 -2786 -1711 -2752
rect -1776 -2811 -1711 -2786
rect -1681 -2811 -1608 -2727
rect -1578 -2731 -1520 -2727
rect -1486 -2731 -1476 -2697
rect -1578 -2765 -1476 -2731
rect -1578 -2799 -1520 -2765
rect -1486 -2799 -1476 -2765
rect -1578 -2811 -1476 -2799
rect -1446 -2727 -1396 -2661
rect -1026 -2657 -1018 -2623
rect -984 -2657 -972 -2623
rect -1026 -2694 -972 -2657
rect -1446 -2757 -1381 -2727
rect -1446 -2791 -1436 -2757
rect -1402 -2791 -1381 -2757
rect -1446 -2811 -1381 -2791
rect -1351 -2747 -1297 -2727
rect -1351 -2781 -1341 -2747
rect -1307 -2781 -1297 -2747
rect -1351 -2811 -1297 -2781
rect -1267 -2811 -1183 -2727
rect -1153 -2757 -1100 -2727
rect -1153 -2791 -1142 -2757
rect -1108 -2791 -1100 -2757
rect -1153 -2811 -1100 -2791
rect -1026 -2728 -1018 -2694
rect -984 -2728 -972 -2694
rect -1026 -2765 -972 -2728
rect -1026 -2799 -1018 -2765
rect -984 -2799 -972 -2765
rect -1026 -2811 -972 -2799
rect -942 -2655 -888 -2611
rect -942 -2689 -932 -2655
rect -898 -2689 -888 -2655
rect -942 -2735 -888 -2689
rect -942 -2769 -932 -2735
rect -898 -2769 -888 -2735
rect -942 -2811 -888 -2769
rect -858 -2623 -806 -2611
rect -858 -2657 -848 -2623
rect -814 -2657 -806 -2623
rect -858 -2691 -806 -2657
rect -655 -2629 -603 -2611
rect -655 -2663 -647 -2629
rect -613 -2663 -603 -2629
rect -655 -2683 -603 -2663
rect -858 -2725 -848 -2691
rect -814 -2725 -806 -2691
rect -858 -2759 -806 -2725
rect -858 -2793 -848 -2759
rect -814 -2793 -806 -2759
rect -858 -2811 -806 -2793
rect -752 -2697 -700 -2683
rect -752 -2731 -744 -2697
rect -710 -2731 -700 -2697
rect -752 -2765 -700 -2731
rect -752 -2799 -744 -2765
rect -710 -2799 -700 -2765
rect -752 -2811 -700 -2799
rect -670 -2697 -603 -2683
rect -670 -2731 -647 -2697
rect -613 -2731 -603 -2697
rect -670 -2765 -603 -2731
rect -670 -2799 -647 -2765
rect -613 -2799 -603 -2765
rect -670 -2811 -603 -2799
rect -573 -2623 -521 -2611
rect -573 -2657 -563 -2623
rect -529 -2657 -521 -2623
rect -573 -2694 -521 -2657
rect -573 -2728 -563 -2694
rect -529 -2728 -521 -2694
rect -573 -2765 -521 -2728
rect -573 -2799 -563 -2765
rect -529 -2799 -521 -2765
rect -573 -2811 -521 -2799
rect -426 -2629 -374 -2611
rect -426 -2663 -418 -2629
rect -384 -2663 -374 -2629
rect -426 -2697 -374 -2663
rect -426 -2731 -418 -2697
rect -384 -2731 -374 -2697
rect -426 -2765 -374 -2731
rect -426 -2799 -418 -2765
rect -384 -2799 -374 -2765
rect -426 -2811 -374 -2799
rect -344 -2629 -292 -2611
rect -344 -2663 -334 -2629
rect -300 -2663 -292 -2629
rect -344 -2697 -292 -2663
rect -344 -2731 -334 -2697
rect -300 -2731 -292 -2697
rect -344 -2765 -292 -2731
rect -344 -2799 -334 -2765
rect -300 -2799 -292 -2765
rect -344 -2811 -292 -2799
rect -181 -2629 -129 -2611
rect -181 -2663 -173 -2629
rect -139 -2663 -129 -2629
rect -181 -2697 -129 -2663
rect -181 -2731 -173 -2697
rect -139 -2731 -129 -2697
rect -181 -2765 -129 -2731
rect -181 -2799 -173 -2765
rect -139 -2799 -129 -2765
rect -181 -2811 -129 -2799
rect -99 -2629 -45 -2611
rect -99 -2663 -89 -2629
rect -55 -2663 -45 -2629
rect -99 -2697 -45 -2663
rect -99 -2731 -89 -2697
rect -55 -2731 -45 -2697
rect -99 -2765 -45 -2731
rect -99 -2799 -89 -2765
rect -55 -2799 -45 -2765
rect -99 -2811 -45 -2799
rect -15 -2697 39 -2611
rect -15 -2731 -5 -2697
rect 29 -2731 39 -2697
rect -15 -2765 39 -2731
rect -15 -2799 -5 -2765
rect 29 -2799 39 -2765
rect -15 -2811 39 -2799
rect 69 -2629 123 -2611
rect 69 -2663 79 -2629
rect 113 -2663 123 -2629
rect 69 -2697 123 -2663
rect 69 -2731 79 -2697
rect 113 -2731 123 -2697
rect 69 -2765 123 -2731
rect 69 -2799 79 -2765
rect 113 -2799 123 -2765
rect 69 -2811 123 -2799
rect 153 -2765 205 -2611
rect 153 -2799 163 -2765
rect 197 -2799 205 -2765
rect 153 -2811 205 -2799
rect 483 -2689 535 -2677
rect 483 -2723 491 -2689
rect 525 -2723 535 -2689
rect 483 -2757 535 -2723
rect 483 -2791 491 -2757
rect 525 -2791 535 -2757
rect 483 -2805 535 -2791
rect 565 -2741 619 -2677
rect 565 -2775 575 -2741
rect 609 -2775 619 -2741
rect 565 -2805 619 -2775
rect 649 -2689 701 -2677
rect 649 -2723 659 -2689
rect 693 -2723 701 -2689
rect 649 -2757 701 -2723
rect 1672 -2623 1726 -2611
rect 1135 -2697 1222 -2661
rect 1135 -2727 1178 -2697
rect 649 -2791 659 -2757
rect 693 -2791 701 -2757
rect 649 -2805 701 -2791
rect 755 -2765 807 -2727
rect 755 -2799 763 -2765
rect 797 -2799 807 -2765
rect 755 -2811 807 -2799
rect 837 -2757 892 -2727
rect 837 -2791 847 -2757
rect 881 -2791 892 -2757
rect 837 -2811 892 -2791
rect 922 -2752 987 -2727
rect 922 -2786 939 -2752
rect 973 -2786 987 -2752
rect 922 -2811 987 -2786
rect 1017 -2811 1090 -2727
rect 1120 -2731 1178 -2727
rect 1212 -2731 1222 -2697
rect 1120 -2765 1222 -2731
rect 1120 -2799 1178 -2765
rect 1212 -2799 1222 -2765
rect 1120 -2811 1222 -2799
rect 1252 -2727 1302 -2661
rect 1672 -2657 1680 -2623
rect 1714 -2657 1726 -2623
rect 1672 -2694 1726 -2657
rect 1252 -2757 1317 -2727
rect 1252 -2791 1262 -2757
rect 1296 -2791 1317 -2757
rect 1252 -2811 1317 -2791
rect 1347 -2747 1401 -2727
rect 1347 -2781 1357 -2747
rect 1391 -2781 1401 -2747
rect 1347 -2811 1401 -2781
rect 1431 -2811 1515 -2727
rect 1545 -2757 1598 -2727
rect 1545 -2791 1556 -2757
rect 1590 -2791 1598 -2757
rect 1545 -2811 1598 -2791
rect 1672 -2728 1680 -2694
rect 1714 -2728 1726 -2694
rect 1672 -2765 1726 -2728
rect 1672 -2799 1680 -2765
rect 1714 -2799 1726 -2765
rect 1672 -2811 1726 -2799
rect 1756 -2655 1810 -2611
rect 1756 -2689 1766 -2655
rect 1800 -2689 1810 -2655
rect 1756 -2735 1810 -2689
rect 1756 -2769 1766 -2735
rect 1800 -2769 1810 -2735
rect 1756 -2811 1810 -2769
rect 1840 -2623 1892 -2611
rect 1840 -2657 1850 -2623
rect 1884 -2657 1892 -2623
rect 1840 -2691 1892 -2657
rect 2043 -2629 2095 -2611
rect 2043 -2663 2051 -2629
rect 2085 -2663 2095 -2629
rect 2043 -2683 2095 -2663
rect 1840 -2725 1850 -2691
rect 1884 -2725 1892 -2691
rect 1840 -2759 1892 -2725
rect 1840 -2793 1850 -2759
rect 1884 -2793 1892 -2759
rect 1840 -2811 1892 -2793
rect 1946 -2697 1998 -2683
rect 1946 -2731 1954 -2697
rect 1988 -2731 1998 -2697
rect 1946 -2765 1998 -2731
rect 1946 -2799 1954 -2765
rect 1988 -2799 1998 -2765
rect 1946 -2811 1998 -2799
rect 2028 -2697 2095 -2683
rect 2028 -2731 2051 -2697
rect 2085 -2731 2095 -2697
rect 2028 -2765 2095 -2731
rect 2028 -2799 2051 -2765
rect 2085 -2799 2095 -2765
rect 2028 -2811 2095 -2799
rect 2125 -2623 2177 -2611
rect 2125 -2657 2135 -2623
rect 2169 -2657 2177 -2623
rect 2125 -2694 2177 -2657
rect 2125 -2728 2135 -2694
rect 2169 -2728 2177 -2694
rect 2125 -2765 2177 -2728
rect 2125 -2799 2135 -2765
rect 2169 -2799 2177 -2765
rect 2125 -2811 2177 -2799
rect 2272 -2629 2324 -2611
rect 2272 -2663 2280 -2629
rect 2314 -2663 2324 -2629
rect 2272 -2697 2324 -2663
rect 2272 -2731 2280 -2697
rect 2314 -2731 2324 -2697
rect 2272 -2765 2324 -2731
rect 2272 -2799 2280 -2765
rect 2314 -2799 2324 -2765
rect 2272 -2811 2324 -2799
rect 2354 -2629 2406 -2611
rect 2354 -2663 2364 -2629
rect 2398 -2663 2406 -2629
rect 2354 -2697 2406 -2663
rect 2354 -2731 2364 -2697
rect 2398 -2731 2406 -2697
rect 2354 -2765 2406 -2731
rect 2354 -2799 2364 -2765
rect 2398 -2799 2406 -2765
rect 2354 -2811 2406 -2799
rect 2517 -2629 2569 -2611
rect 2517 -2663 2525 -2629
rect 2559 -2663 2569 -2629
rect 2517 -2697 2569 -2663
rect 2517 -2731 2525 -2697
rect 2559 -2731 2569 -2697
rect 2517 -2765 2569 -2731
rect 2517 -2799 2525 -2765
rect 2559 -2799 2569 -2765
rect 2517 -2811 2569 -2799
rect 2599 -2629 2653 -2611
rect 2599 -2663 2609 -2629
rect 2643 -2663 2653 -2629
rect 2599 -2697 2653 -2663
rect 2599 -2731 2609 -2697
rect 2643 -2731 2653 -2697
rect 2599 -2765 2653 -2731
rect 2599 -2799 2609 -2765
rect 2643 -2799 2653 -2765
rect 2599 -2811 2653 -2799
rect 2683 -2697 2737 -2611
rect 2683 -2731 2693 -2697
rect 2727 -2731 2737 -2697
rect 2683 -2765 2737 -2731
rect 2683 -2799 2693 -2765
rect 2727 -2799 2737 -2765
rect 2683 -2811 2737 -2799
rect 2767 -2629 2821 -2611
rect 2767 -2663 2777 -2629
rect 2811 -2663 2821 -2629
rect 2767 -2697 2821 -2663
rect 2767 -2731 2777 -2697
rect 2811 -2731 2821 -2697
rect 2767 -2765 2821 -2731
rect 2767 -2799 2777 -2765
rect 2811 -2799 2821 -2765
rect 2767 -2811 2821 -2799
rect 2851 -2765 2903 -2611
rect 2851 -2799 2861 -2765
rect 2895 -2799 2903 -2765
rect 2851 -2811 2903 -2799
<< ndiffc >>
rect -2207 -53 -2173 -19
rect -2123 -79 -2089 -45
rect -2039 -53 -2005 -19
rect -1935 -79 -1901 -45
rect -1850 -65 -1816 -31
rect -1739 -65 -1705 -31
rect -1540 -71 -1506 -37
rect -1421 -65 -1387 -31
rect -1318 -65 -1284 -31
rect -1120 -65 -1086 -31
rect -1014 -10 -980 24
rect -1014 -78 -980 -44
rect -930 -49 -896 -15
rect -846 -8 -812 26
rect -846 -76 -812 -42
rect -742 -53 -708 -19
rect -647 -79 -613 -45
rect -563 -41 -529 -7
rect -418 -7 -384 27
rect -418 -75 -384 -41
rect -334 -7 -300 27
rect -334 -75 -300 -41
rect -173 -79 -139 -45
rect -89 -71 -55 -37
rect -5 -79 29 -45
rect 79 -71 113 -37
rect 163 -78 197 -44
rect -2207 -257 -2173 -223
rect -2123 -231 -2089 -197
rect -2039 -257 -2005 -223
rect -1935 -231 -1901 -197
rect -1850 -245 -1816 -211
rect -1739 -245 -1705 -211
rect -1540 -239 -1506 -205
rect -1421 -245 -1387 -211
rect -1318 -245 -1284 -211
rect -1120 -245 -1086 -211
rect -1014 -232 -980 -198
rect -1014 -300 -980 -266
rect -930 -261 -896 -227
rect -846 -234 -812 -200
rect -846 -302 -812 -268
rect -742 -257 -708 -223
rect -647 -231 -613 -197
rect -563 -269 -529 -235
rect -418 -235 -384 -201
rect -418 -303 -384 -269
rect -334 -235 -300 -201
rect -334 -303 -300 -269
rect -173 -231 -139 -197
rect -89 -239 -55 -205
rect -5 -231 29 -197
rect 79 -239 113 -205
rect 163 -232 197 -198
rect 491 -257 525 -223
rect 575 -231 609 -197
rect 659 -257 693 -223
rect 763 -231 797 -197
rect 848 -245 882 -211
rect 959 -245 993 -211
rect 1158 -239 1192 -205
rect 1277 -245 1311 -211
rect 1380 -245 1414 -211
rect 1578 -245 1612 -211
rect 1684 -232 1718 -198
rect 1684 -300 1718 -266
rect 1768 -261 1802 -227
rect 1852 -234 1886 -200
rect 1852 -302 1886 -268
rect 1956 -257 1990 -223
rect 2051 -231 2085 -197
rect 2135 -269 2169 -235
rect 2280 -235 2314 -201
rect 2280 -303 2314 -269
rect 2364 -235 2398 -201
rect 2364 -303 2398 -269
rect 2525 -231 2559 -197
rect 2609 -239 2643 -205
rect 2693 -231 2727 -197
rect 2777 -239 2811 -205
rect 2861 -232 2895 -198
rect -2207 -1141 -2173 -1107
rect -2123 -1167 -2089 -1133
rect -2039 -1141 -2005 -1107
rect -1935 -1167 -1901 -1133
rect -1850 -1153 -1816 -1119
rect -1739 -1153 -1705 -1119
rect -1540 -1159 -1506 -1125
rect -1421 -1153 -1387 -1119
rect -1318 -1153 -1284 -1119
rect -1120 -1153 -1086 -1119
rect -1014 -1098 -980 -1064
rect -1014 -1166 -980 -1132
rect -930 -1137 -896 -1103
rect -846 -1096 -812 -1062
rect -846 -1164 -812 -1130
rect -742 -1141 -708 -1107
rect -647 -1167 -613 -1133
rect -563 -1129 -529 -1095
rect -418 -1095 -384 -1061
rect -418 -1163 -384 -1129
rect -334 -1095 -300 -1061
rect -334 -1163 -300 -1129
rect -173 -1167 -139 -1133
rect -89 -1159 -55 -1125
rect -5 -1167 29 -1133
rect 79 -1159 113 -1125
rect 163 -1166 197 -1132
rect 491 -1141 525 -1107
rect 575 -1167 609 -1133
rect 659 -1141 693 -1107
rect 763 -1167 797 -1133
rect 848 -1153 882 -1119
rect 959 -1153 993 -1119
rect 1158 -1159 1192 -1125
rect 1277 -1153 1311 -1119
rect 1380 -1153 1414 -1119
rect 1578 -1153 1612 -1119
rect 1684 -1098 1718 -1064
rect 1684 -1166 1718 -1132
rect 1768 -1137 1802 -1103
rect 1852 -1096 1886 -1062
rect 1852 -1164 1886 -1130
rect 1956 -1141 1990 -1107
rect 2051 -1167 2085 -1133
rect 2135 -1129 2169 -1095
rect 2280 -1095 2314 -1061
rect 2280 -1163 2314 -1129
rect 2364 -1095 2398 -1061
rect 2364 -1163 2398 -1129
rect 2525 -1167 2559 -1133
rect 2609 -1159 2643 -1125
rect 2693 -1167 2727 -1133
rect 2777 -1159 2811 -1125
rect 2861 -1166 2895 -1132
rect -2207 -1345 -2173 -1311
rect -2123 -1319 -2089 -1285
rect -2039 -1345 -2005 -1311
rect -1935 -1319 -1901 -1285
rect -1850 -1333 -1816 -1299
rect -1739 -1333 -1705 -1299
rect -1540 -1327 -1506 -1293
rect -1421 -1333 -1387 -1299
rect -1318 -1333 -1284 -1299
rect -1120 -1333 -1086 -1299
rect -1014 -1320 -980 -1286
rect -1014 -1388 -980 -1354
rect -930 -1349 -896 -1315
rect -846 -1322 -812 -1288
rect -846 -1390 -812 -1356
rect -742 -1345 -708 -1311
rect -647 -1319 -613 -1285
rect -563 -1357 -529 -1323
rect -418 -1323 -384 -1289
rect -418 -1391 -384 -1357
rect -334 -1323 -300 -1289
rect -334 -1391 -300 -1357
rect -173 -1319 -139 -1285
rect -89 -1327 -55 -1293
rect -5 -1319 29 -1285
rect 79 -1327 113 -1293
rect 163 -1320 197 -1286
rect 491 -1345 525 -1311
rect 575 -1319 609 -1285
rect 659 -1345 693 -1311
rect 763 -1319 797 -1285
rect 848 -1333 882 -1299
rect 959 -1333 993 -1299
rect 1158 -1327 1192 -1293
rect 1277 -1333 1311 -1299
rect 1380 -1333 1414 -1299
rect 1578 -1333 1612 -1299
rect 1684 -1320 1718 -1286
rect 1684 -1388 1718 -1354
rect 1768 -1349 1802 -1315
rect 1852 -1322 1886 -1288
rect 1852 -1390 1886 -1356
rect 1956 -1345 1990 -1311
rect 2051 -1319 2085 -1285
rect 2135 -1357 2169 -1323
rect 2280 -1323 2314 -1289
rect 2280 -1391 2314 -1357
rect 2364 -1323 2398 -1289
rect 2364 -1391 2398 -1357
rect 2525 -1319 2559 -1285
rect 2609 -1327 2643 -1293
rect 2693 -1319 2727 -1285
rect 2777 -1327 2811 -1293
rect 2861 -1320 2895 -1286
rect -2207 -2229 -2173 -2195
rect -2123 -2255 -2089 -2221
rect -2039 -2229 -2005 -2195
rect -1935 -2255 -1901 -2221
rect -1850 -2241 -1816 -2207
rect -1739 -2241 -1705 -2207
rect -1540 -2247 -1506 -2213
rect -1421 -2241 -1387 -2207
rect -1318 -2241 -1284 -2207
rect -1120 -2241 -1086 -2207
rect -1014 -2186 -980 -2152
rect -1014 -2254 -980 -2220
rect -930 -2225 -896 -2191
rect -846 -2184 -812 -2150
rect -846 -2252 -812 -2218
rect -742 -2229 -708 -2195
rect -647 -2255 -613 -2221
rect -563 -2217 -529 -2183
rect -418 -2183 -384 -2149
rect -418 -2251 -384 -2217
rect -334 -2183 -300 -2149
rect -334 -2251 -300 -2217
rect -173 -2255 -139 -2221
rect -89 -2247 -55 -2213
rect -5 -2255 29 -2221
rect 79 -2247 113 -2213
rect 163 -2254 197 -2220
rect 491 -2229 525 -2195
rect 575 -2255 609 -2221
rect 659 -2229 693 -2195
rect 763 -2255 797 -2221
rect 848 -2241 882 -2207
rect 959 -2241 993 -2207
rect 1158 -2247 1192 -2213
rect 1277 -2241 1311 -2207
rect 1380 -2241 1414 -2207
rect 1578 -2241 1612 -2207
rect 1684 -2186 1718 -2152
rect 1684 -2254 1718 -2220
rect 1768 -2225 1802 -2191
rect 1852 -2184 1886 -2150
rect 1852 -2252 1886 -2218
rect 1956 -2229 1990 -2195
rect 2051 -2255 2085 -2221
rect 2135 -2217 2169 -2183
rect 2280 -2183 2314 -2149
rect 2280 -2251 2314 -2217
rect 2364 -2183 2398 -2149
rect 2364 -2251 2398 -2217
rect 2525 -2255 2559 -2221
rect 2609 -2247 2643 -2213
rect 2693 -2255 2727 -2221
rect 2777 -2247 2811 -2213
rect 2861 -2254 2895 -2220
rect -2207 -2433 -2173 -2399
rect -2123 -2407 -2089 -2373
rect -2039 -2433 -2005 -2399
rect -1935 -2407 -1901 -2373
rect -1850 -2421 -1816 -2387
rect -1739 -2421 -1705 -2387
rect -1540 -2415 -1506 -2381
rect -1421 -2421 -1387 -2387
rect -1318 -2421 -1284 -2387
rect -1120 -2421 -1086 -2387
rect -1014 -2408 -980 -2374
rect -1014 -2476 -980 -2442
rect -930 -2437 -896 -2403
rect -846 -2410 -812 -2376
rect -846 -2478 -812 -2444
rect -742 -2433 -708 -2399
rect -647 -2407 -613 -2373
rect -563 -2445 -529 -2411
rect -418 -2411 -384 -2377
rect -418 -2479 -384 -2445
rect -334 -2411 -300 -2377
rect -334 -2479 -300 -2445
rect -173 -2407 -139 -2373
rect -89 -2415 -55 -2381
rect -5 -2407 29 -2373
rect 79 -2415 113 -2381
rect 163 -2408 197 -2374
rect 491 -2433 525 -2399
rect 575 -2407 609 -2373
rect 659 -2433 693 -2399
rect 763 -2407 797 -2373
rect 848 -2421 882 -2387
rect 959 -2421 993 -2387
rect 1158 -2415 1192 -2381
rect 1277 -2421 1311 -2387
rect 1380 -2421 1414 -2387
rect 1578 -2421 1612 -2387
rect 1684 -2408 1718 -2374
rect 1684 -2476 1718 -2442
rect 1768 -2437 1802 -2403
rect 1852 -2410 1886 -2376
rect 1852 -2478 1886 -2444
rect 1956 -2433 1990 -2399
rect 2051 -2407 2085 -2373
rect 2135 -2445 2169 -2411
rect 2280 -2411 2314 -2377
rect 2280 -2479 2314 -2445
rect 2364 -2411 2398 -2377
rect 2364 -2479 2398 -2445
rect 2525 -2407 2559 -2373
rect 2609 -2415 2643 -2381
rect 2693 -2407 2727 -2373
rect 2777 -2415 2811 -2381
rect 2861 -2408 2895 -2374
<< pdiffc >>
rect -2207 305 -2173 339
rect -2207 237 -2173 271
rect -2123 289 -2089 323
rect -2039 305 -2005 339
rect -1935 313 -1901 347
rect -1851 305 -1817 339
rect -1759 300 -1725 334
rect -1520 313 -1486 347
rect -2039 237 -2005 271
rect -1520 245 -1486 279
rect -1436 305 -1402 339
rect -1341 295 -1307 329
rect -1142 305 -1108 339
rect -1018 313 -984 347
rect -1018 242 -984 276
rect -1018 171 -984 205
rect -932 283 -898 317
rect -932 203 -898 237
rect -848 307 -814 341
rect -848 239 -814 273
rect -744 313 -710 347
rect -744 245 -710 279
rect -647 313 -613 347
rect -647 245 -613 279
rect -848 171 -814 205
rect -647 177 -613 211
rect -563 313 -529 347
rect -563 242 -529 276
rect -563 171 -529 205
rect -418 313 -384 347
rect -418 245 -384 279
rect -418 177 -384 211
rect -334 313 -300 347
rect -334 245 -300 279
rect -334 177 -300 211
rect -173 313 -139 347
rect -173 245 -139 279
rect -173 177 -139 211
rect -89 313 -55 347
rect -89 245 -55 279
rect -89 177 -55 211
rect -5 313 29 347
rect -5 245 29 279
rect 79 313 113 347
rect 79 245 113 279
rect 79 177 113 211
rect 163 313 197 347
rect -2207 -547 -2173 -513
rect -2207 -615 -2173 -581
rect -2123 -599 -2089 -565
rect -2039 -547 -2005 -513
rect -2039 -615 -2005 -581
rect -1935 -623 -1901 -589
rect -1851 -615 -1817 -581
rect -1759 -610 -1725 -576
rect -1520 -555 -1486 -521
rect -1520 -623 -1486 -589
rect -1018 -481 -984 -447
rect -1436 -615 -1402 -581
rect -1341 -605 -1307 -571
rect -1142 -615 -1108 -581
rect -1018 -552 -984 -518
rect -1018 -623 -984 -589
rect -932 -513 -898 -479
rect -932 -593 -898 -559
rect -848 -481 -814 -447
rect -647 -487 -613 -453
rect -848 -549 -814 -515
rect -848 -617 -814 -583
rect -744 -555 -710 -521
rect -744 -623 -710 -589
rect -647 -555 -613 -521
rect -647 -623 -613 -589
rect -563 -481 -529 -447
rect -563 -552 -529 -518
rect -563 -623 -529 -589
rect -418 -487 -384 -453
rect -418 -555 -384 -521
rect -418 -623 -384 -589
rect -334 -487 -300 -453
rect -334 -555 -300 -521
rect -334 -623 -300 -589
rect -173 -487 -139 -453
rect -173 -555 -139 -521
rect -173 -623 -139 -589
rect -89 -487 -55 -453
rect -89 -555 -55 -521
rect -89 -623 -55 -589
rect -5 -555 29 -521
rect -5 -623 29 -589
rect 79 -487 113 -453
rect 79 -555 113 -521
rect 79 -623 113 -589
rect 163 -623 197 -589
rect 491 -547 525 -513
rect 491 -615 525 -581
rect 575 -599 609 -565
rect 659 -547 693 -513
rect 659 -615 693 -581
rect 763 -623 797 -589
rect 847 -615 881 -581
rect 939 -610 973 -576
rect 1178 -555 1212 -521
rect 1178 -623 1212 -589
rect 1680 -481 1714 -447
rect 1262 -615 1296 -581
rect 1357 -605 1391 -571
rect 1556 -615 1590 -581
rect 1680 -552 1714 -518
rect 1680 -623 1714 -589
rect 1766 -513 1800 -479
rect 1766 -593 1800 -559
rect 1850 -481 1884 -447
rect 2051 -487 2085 -453
rect 1850 -549 1884 -515
rect 1850 -617 1884 -583
rect 1954 -555 1988 -521
rect 1954 -623 1988 -589
rect 2051 -555 2085 -521
rect 2051 -623 2085 -589
rect 2135 -481 2169 -447
rect 2135 -552 2169 -518
rect 2135 -623 2169 -589
rect 2280 -487 2314 -453
rect 2280 -555 2314 -521
rect 2280 -623 2314 -589
rect 2364 -487 2398 -453
rect 2364 -555 2398 -521
rect 2364 -623 2398 -589
rect 2525 -487 2559 -453
rect 2525 -555 2559 -521
rect 2525 -623 2559 -589
rect 2609 -487 2643 -453
rect 2609 -555 2643 -521
rect 2609 -623 2643 -589
rect 2693 -555 2727 -521
rect 2693 -623 2727 -589
rect 2777 -487 2811 -453
rect 2777 -555 2811 -521
rect 2777 -623 2811 -589
rect 2861 -623 2895 -589
rect -2207 -783 -2173 -749
rect -2207 -851 -2173 -817
rect -2123 -799 -2089 -765
rect -2039 -783 -2005 -749
rect -1935 -775 -1901 -741
rect -1851 -783 -1817 -749
rect -1759 -788 -1725 -754
rect -1520 -775 -1486 -741
rect -2039 -851 -2005 -817
rect -1520 -843 -1486 -809
rect -1436 -783 -1402 -749
rect -1341 -793 -1307 -759
rect -1142 -783 -1108 -749
rect -1018 -775 -984 -741
rect -1018 -846 -984 -812
rect -1018 -917 -984 -883
rect -932 -805 -898 -771
rect -932 -885 -898 -851
rect -848 -781 -814 -747
rect -848 -849 -814 -815
rect -744 -775 -710 -741
rect -744 -843 -710 -809
rect -647 -775 -613 -741
rect -647 -843 -613 -809
rect -848 -917 -814 -883
rect -647 -911 -613 -877
rect -563 -775 -529 -741
rect -563 -846 -529 -812
rect -563 -917 -529 -883
rect -418 -775 -384 -741
rect -418 -843 -384 -809
rect -418 -911 -384 -877
rect -334 -775 -300 -741
rect -334 -843 -300 -809
rect -334 -911 -300 -877
rect -173 -775 -139 -741
rect -173 -843 -139 -809
rect -173 -911 -139 -877
rect -89 -775 -55 -741
rect -89 -843 -55 -809
rect -89 -911 -55 -877
rect -5 -775 29 -741
rect -5 -843 29 -809
rect 79 -775 113 -741
rect 79 -843 113 -809
rect 79 -911 113 -877
rect 163 -775 197 -741
rect 491 -783 525 -749
rect 491 -851 525 -817
rect 575 -799 609 -765
rect 659 -783 693 -749
rect 763 -775 797 -741
rect 847 -783 881 -749
rect 939 -788 973 -754
rect 1178 -775 1212 -741
rect 659 -851 693 -817
rect 1178 -843 1212 -809
rect 1262 -783 1296 -749
rect 1357 -793 1391 -759
rect 1556 -783 1590 -749
rect 1680 -775 1714 -741
rect 1680 -846 1714 -812
rect 1680 -917 1714 -883
rect 1766 -805 1800 -771
rect 1766 -885 1800 -851
rect 1850 -781 1884 -747
rect 1850 -849 1884 -815
rect 1954 -775 1988 -741
rect 1954 -843 1988 -809
rect 2051 -775 2085 -741
rect 2051 -843 2085 -809
rect 1850 -917 1884 -883
rect 2051 -911 2085 -877
rect 2135 -775 2169 -741
rect 2135 -846 2169 -812
rect 2135 -917 2169 -883
rect 2280 -775 2314 -741
rect 2280 -843 2314 -809
rect 2280 -911 2314 -877
rect 2364 -775 2398 -741
rect 2364 -843 2398 -809
rect 2364 -911 2398 -877
rect 2525 -775 2559 -741
rect 2525 -843 2559 -809
rect 2525 -911 2559 -877
rect 2609 -775 2643 -741
rect 2609 -843 2643 -809
rect 2609 -911 2643 -877
rect 2693 -775 2727 -741
rect 2693 -843 2727 -809
rect 2777 -775 2811 -741
rect 2777 -843 2811 -809
rect 2777 -911 2811 -877
rect 2861 -775 2895 -741
rect -2207 -1635 -2173 -1601
rect -2207 -1703 -2173 -1669
rect -2123 -1687 -2089 -1653
rect -2039 -1635 -2005 -1601
rect -2039 -1703 -2005 -1669
rect -1935 -1711 -1901 -1677
rect -1851 -1703 -1817 -1669
rect -1759 -1698 -1725 -1664
rect -1520 -1643 -1486 -1609
rect -1520 -1711 -1486 -1677
rect -1018 -1569 -984 -1535
rect -1436 -1703 -1402 -1669
rect -1341 -1693 -1307 -1659
rect -1142 -1703 -1108 -1669
rect -1018 -1640 -984 -1606
rect -1018 -1711 -984 -1677
rect -932 -1601 -898 -1567
rect -932 -1681 -898 -1647
rect -848 -1569 -814 -1535
rect -647 -1575 -613 -1541
rect -848 -1637 -814 -1603
rect -848 -1705 -814 -1671
rect -744 -1643 -710 -1609
rect -744 -1711 -710 -1677
rect -647 -1643 -613 -1609
rect -647 -1711 -613 -1677
rect -563 -1569 -529 -1535
rect -563 -1640 -529 -1606
rect -563 -1711 -529 -1677
rect -418 -1575 -384 -1541
rect -418 -1643 -384 -1609
rect -418 -1711 -384 -1677
rect -334 -1575 -300 -1541
rect -334 -1643 -300 -1609
rect -334 -1711 -300 -1677
rect -173 -1575 -139 -1541
rect -173 -1643 -139 -1609
rect -173 -1711 -139 -1677
rect -89 -1575 -55 -1541
rect -89 -1643 -55 -1609
rect -89 -1711 -55 -1677
rect -5 -1643 29 -1609
rect -5 -1711 29 -1677
rect 79 -1575 113 -1541
rect 79 -1643 113 -1609
rect 79 -1711 113 -1677
rect 163 -1711 197 -1677
rect 491 -1635 525 -1601
rect 491 -1703 525 -1669
rect 575 -1687 609 -1653
rect 659 -1635 693 -1601
rect 659 -1703 693 -1669
rect 763 -1711 797 -1677
rect 847 -1703 881 -1669
rect 939 -1698 973 -1664
rect 1178 -1643 1212 -1609
rect 1178 -1711 1212 -1677
rect 1680 -1569 1714 -1535
rect 1262 -1703 1296 -1669
rect 1357 -1693 1391 -1659
rect 1556 -1703 1590 -1669
rect 1680 -1640 1714 -1606
rect 1680 -1711 1714 -1677
rect 1766 -1601 1800 -1567
rect 1766 -1681 1800 -1647
rect 1850 -1569 1884 -1535
rect 2051 -1575 2085 -1541
rect 1850 -1637 1884 -1603
rect 1850 -1705 1884 -1671
rect 1954 -1643 1988 -1609
rect 1954 -1711 1988 -1677
rect 2051 -1643 2085 -1609
rect 2051 -1711 2085 -1677
rect 2135 -1569 2169 -1535
rect 2135 -1640 2169 -1606
rect 2135 -1711 2169 -1677
rect 2280 -1575 2314 -1541
rect 2280 -1643 2314 -1609
rect 2280 -1711 2314 -1677
rect 2364 -1575 2398 -1541
rect 2364 -1643 2398 -1609
rect 2364 -1711 2398 -1677
rect 2525 -1575 2559 -1541
rect 2525 -1643 2559 -1609
rect 2525 -1711 2559 -1677
rect 2609 -1575 2643 -1541
rect 2609 -1643 2643 -1609
rect 2609 -1711 2643 -1677
rect 2693 -1643 2727 -1609
rect 2693 -1711 2727 -1677
rect 2777 -1575 2811 -1541
rect 2777 -1643 2811 -1609
rect 2777 -1711 2811 -1677
rect 2861 -1711 2895 -1677
rect -2207 -1871 -2173 -1837
rect -2207 -1939 -2173 -1905
rect -2123 -1887 -2089 -1853
rect -2039 -1871 -2005 -1837
rect -1935 -1863 -1901 -1829
rect -1851 -1871 -1817 -1837
rect -1759 -1876 -1725 -1842
rect -1520 -1863 -1486 -1829
rect -2039 -1939 -2005 -1905
rect -1520 -1931 -1486 -1897
rect -1436 -1871 -1402 -1837
rect -1341 -1881 -1307 -1847
rect -1142 -1871 -1108 -1837
rect -1018 -1863 -984 -1829
rect -1018 -1934 -984 -1900
rect -1018 -2005 -984 -1971
rect -932 -1893 -898 -1859
rect -932 -1973 -898 -1939
rect -848 -1869 -814 -1835
rect -848 -1937 -814 -1903
rect -744 -1863 -710 -1829
rect -744 -1931 -710 -1897
rect -647 -1863 -613 -1829
rect -647 -1931 -613 -1897
rect -848 -2005 -814 -1971
rect -647 -1999 -613 -1965
rect -563 -1863 -529 -1829
rect -563 -1934 -529 -1900
rect -563 -2005 -529 -1971
rect -418 -1863 -384 -1829
rect -418 -1931 -384 -1897
rect -418 -1999 -384 -1965
rect -334 -1863 -300 -1829
rect -334 -1931 -300 -1897
rect -334 -1999 -300 -1965
rect -173 -1863 -139 -1829
rect -173 -1931 -139 -1897
rect -173 -1999 -139 -1965
rect -89 -1863 -55 -1829
rect -89 -1931 -55 -1897
rect -89 -1999 -55 -1965
rect -5 -1863 29 -1829
rect -5 -1931 29 -1897
rect 79 -1863 113 -1829
rect 79 -1931 113 -1897
rect 79 -1999 113 -1965
rect 163 -1863 197 -1829
rect 491 -1871 525 -1837
rect 491 -1939 525 -1905
rect 575 -1887 609 -1853
rect 659 -1871 693 -1837
rect 763 -1863 797 -1829
rect 847 -1871 881 -1837
rect 939 -1876 973 -1842
rect 1178 -1863 1212 -1829
rect 659 -1939 693 -1905
rect 1178 -1931 1212 -1897
rect 1262 -1871 1296 -1837
rect 1357 -1881 1391 -1847
rect 1556 -1871 1590 -1837
rect 1680 -1863 1714 -1829
rect 1680 -1934 1714 -1900
rect 1680 -2005 1714 -1971
rect 1766 -1893 1800 -1859
rect 1766 -1973 1800 -1939
rect 1850 -1869 1884 -1835
rect 1850 -1937 1884 -1903
rect 1954 -1863 1988 -1829
rect 1954 -1931 1988 -1897
rect 2051 -1863 2085 -1829
rect 2051 -1931 2085 -1897
rect 1850 -2005 1884 -1971
rect 2051 -1999 2085 -1965
rect 2135 -1863 2169 -1829
rect 2135 -1934 2169 -1900
rect 2135 -2005 2169 -1971
rect 2280 -1863 2314 -1829
rect 2280 -1931 2314 -1897
rect 2280 -1999 2314 -1965
rect 2364 -1863 2398 -1829
rect 2364 -1931 2398 -1897
rect 2364 -1999 2398 -1965
rect 2525 -1863 2559 -1829
rect 2525 -1931 2559 -1897
rect 2525 -1999 2559 -1965
rect 2609 -1863 2643 -1829
rect 2609 -1931 2643 -1897
rect 2609 -1999 2643 -1965
rect 2693 -1863 2727 -1829
rect 2693 -1931 2727 -1897
rect 2777 -1863 2811 -1829
rect 2777 -1931 2811 -1897
rect 2777 -1999 2811 -1965
rect 2861 -1863 2895 -1829
rect -2207 -2723 -2173 -2689
rect -2207 -2791 -2173 -2757
rect -2123 -2775 -2089 -2741
rect -2039 -2723 -2005 -2689
rect -2039 -2791 -2005 -2757
rect -1935 -2799 -1901 -2765
rect -1851 -2791 -1817 -2757
rect -1759 -2786 -1725 -2752
rect -1520 -2731 -1486 -2697
rect -1520 -2799 -1486 -2765
rect -1018 -2657 -984 -2623
rect -1436 -2791 -1402 -2757
rect -1341 -2781 -1307 -2747
rect -1142 -2791 -1108 -2757
rect -1018 -2728 -984 -2694
rect -1018 -2799 -984 -2765
rect -932 -2689 -898 -2655
rect -932 -2769 -898 -2735
rect -848 -2657 -814 -2623
rect -647 -2663 -613 -2629
rect -848 -2725 -814 -2691
rect -848 -2793 -814 -2759
rect -744 -2731 -710 -2697
rect -744 -2799 -710 -2765
rect -647 -2731 -613 -2697
rect -647 -2799 -613 -2765
rect -563 -2657 -529 -2623
rect -563 -2728 -529 -2694
rect -563 -2799 -529 -2765
rect -418 -2663 -384 -2629
rect -418 -2731 -384 -2697
rect -418 -2799 -384 -2765
rect -334 -2663 -300 -2629
rect -334 -2731 -300 -2697
rect -334 -2799 -300 -2765
rect -173 -2663 -139 -2629
rect -173 -2731 -139 -2697
rect -173 -2799 -139 -2765
rect -89 -2663 -55 -2629
rect -89 -2731 -55 -2697
rect -89 -2799 -55 -2765
rect -5 -2731 29 -2697
rect -5 -2799 29 -2765
rect 79 -2663 113 -2629
rect 79 -2731 113 -2697
rect 79 -2799 113 -2765
rect 163 -2799 197 -2765
rect 491 -2723 525 -2689
rect 491 -2791 525 -2757
rect 575 -2775 609 -2741
rect 659 -2723 693 -2689
rect 659 -2791 693 -2757
rect 763 -2799 797 -2765
rect 847 -2791 881 -2757
rect 939 -2786 973 -2752
rect 1178 -2731 1212 -2697
rect 1178 -2799 1212 -2765
rect 1680 -2657 1714 -2623
rect 1262 -2791 1296 -2757
rect 1357 -2781 1391 -2747
rect 1556 -2791 1590 -2757
rect 1680 -2728 1714 -2694
rect 1680 -2799 1714 -2765
rect 1766 -2689 1800 -2655
rect 1766 -2769 1800 -2735
rect 1850 -2657 1884 -2623
rect 2051 -2663 2085 -2629
rect 1850 -2725 1884 -2691
rect 1850 -2793 1884 -2759
rect 1954 -2731 1988 -2697
rect 1954 -2799 1988 -2765
rect 2051 -2731 2085 -2697
rect 2051 -2799 2085 -2765
rect 2135 -2657 2169 -2623
rect 2135 -2728 2169 -2694
rect 2135 -2799 2169 -2765
rect 2280 -2663 2314 -2629
rect 2280 -2731 2314 -2697
rect 2280 -2799 2314 -2765
rect 2364 -2663 2398 -2629
rect 2364 -2731 2398 -2697
rect 2364 -2799 2398 -2765
rect 2525 -2663 2559 -2629
rect 2525 -2731 2559 -2697
rect 2525 -2799 2559 -2765
rect 2609 -2663 2643 -2629
rect 2609 -2731 2643 -2697
rect 2609 -2799 2643 -2765
rect 2693 -2731 2727 -2697
rect 2693 -2799 2727 -2765
rect 2777 -2663 2811 -2629
rect 2777 -2731 2811 -2697
rect 2777 -2799 2811 -2765
rect 2861 -2799 2895 -2765
<< psubdiff >>
rect -2555 7 -2521 31
rect -2555 -74 -2521 -27
rect 345 7 379 31
rect 345 -74 379 -27
rect 3219 7 3253 31
rect 3219 -74 3253 -27
rect -2555 -249 -2521 -202
rect -2555 -307 -2521 -283
rect 3219 -249 3253 -202
rect 3219 -307 3253 -283
rect -2555 -1081 -2521 -1057
rect -2555 -1162 -2521 -1115
rect 3219 -1081 3253 -1057
rect 3219 -1162 3253 -1115
rect -2555 -1337 -2521 -1290
rect -2555 -1395 -2521 -1371
rect 3219 -1337 3253 -1290
rect 3219 -1395 3253 -1371
rect -2555 -2169 -2521 -2145
rect -2555 -2250 -2521 -2203
rect 3219 -2169 3253 -2145
rect 3219 -2250 3253 -2203
rect -2555 -2425 -2521 -2378
rect -2555 -2483 -2521 -2459
rect 3219 -2425 3253 -2378
rect 3219 -2483 3253 -2459
<< nsubdiff >>
rect -2555 318 -2521 342
rect -2555 225 -2521 284
rect -2555 167 -2521 191
rect 345 318 379 342
rect 345 225 379 284
rect 345 167 379 191
rect 3219 318 3253 342
rect 3219 225 3253 284
rect 3219 167 3253 191
rect -2555 -467 -2521 -443
rect -2555 -560 -2521 -501
rect -2555 -618 -2521 -594
rect 3219 -467 3253 -443
rect 3219 -560 3253 -501
rect 3219 -618 3253 -594
rect -2555 -770 -2521 -746
rect -2555 -863 -2521 -804
rect -2555 -921 -2521 -897
rect 3219 -770 3253 -746
rect 3219 -863 3253 -804
rect 3219 -921 3253 -897
rect -2555 -1555 -2521 -1531
rect -2555 -1648 -2521 -1589
rect -2555 -1706 -2521 -1682
rect 3219 -1555 3253 -1531
rect 3219 -1648 3253 -1589
rect 3219 -1706 3253 -1682
rect -2555 -1858 -2521 -1834
rect -2555 -1951 -2521 -1892
rect -2555 -2009 -2521 -1985
rect 3219 -1858 3253 -1834
rect 3219 -1951 3253 -1892
rect 3219 -2009 3253 -1985
rect -2555 -2643 -2521 -2619
rect -2555 -2736 -2521 -2677
rect -2555 -2794 -2521 -2770
rect 3219 -2643 3253 -2619
rect 3219 -2736 3253 -2677
rect 3219 -2794 3253 -2770
<< psubdiffcont >>
rect -2555 -27 -2521 7
rect 345 -27 379 7
rect 3219 -27 3253 7
rect -2555 -283 -2521 -249
rect 3219 -283 3253 -249
rect -2555 -1115 -2521 -1081
rect 3219 -1115 3253 -1081
rect -2555 -1371 -2521 -1337
rect 3219 -1371 3253 -1337
rect -2555 -2203 -2521 -2169
rect 3219 -2203 3253 -2169
rect -2555 -2459 -2521 -2425
rect 3219 -2459 3253 -2425
<< nsubdiffcont >>
rect -2555 284 -2521 318
rect -2555 191 -2521 225
rect 345 284 379 318
rect 345 191 379 225
rect 3219 284 3253 318
rect 3219 191 3253 225
rect -2555 -501 -2521 -467
rect -2555 -594 -2521 -560
rect 3219 -501 3253 -467
rect 3219 -594 3253 -560
rect -2555 -804 -2521 -770
rect -2555 -897 -2521 -863
rect 3219 -804 3253 -770
rect 3219 -897 3253 -863
rect -2555 -1589 -2521 -1555
rect -2555 -1682 -2521 -1648
rect 3219 -1589 3253 -1555
rect 3219 -1682 3253 -1648
rect -2555 -1892 -2521 -1858
rect -2555 -1985 -2521 -1951
rect 3219 -1892 3253 -1858
rect 3219 -1985 3253 -1951
rect -2555 -2677 -2521 -2643
rect -2555 -2770 -2521 -2736
rect 3219 -2677 3253 -2643
rect 3219 -2770 3253 -2736
<< poly >>
rect -2163 353 -2133 379
rect -2079 353 -2049 379
rect -1891 359 -1861 385
rect -1806 359 -1776 385
rect -1711 359 -1681 385
rect -1608 359 -1578 385
rect -1476 359 -1446 385
rect -1381 359 -1351 385
rect -1297 359 -1267 385
rect -1183 359 -1153 385
rect -972 359 -942 385
rect -888 359 -858 385
rect -700 359 -670 385
rect -603 359 -573 385
rect -374 359 -344 385
rect -129 359 -99 385
rect -45 359 -15 385
rect 39 359 69 385
rect 123 359 153 385
rect -2163 210 -2133 225
rect -2196 180 -2133 210
rect -2196 127 -2166 180
rect -2079 136 -2049 225
rect -1891 195 -1861 275
rect -2220 111 -2166 127
rect -2220 77 -2210 111
rect -2176 77 -2166 111
rect -2124 126 -2049 136
rect -1956 179 -1861 195
rect -1956 145 -1946 179
rect -1912 145 -1861 179
rect -1806 159 -1776 275
rect -1711 243 -1681 275
rect -1711 227 -1650 243
rect -1711 193 -1694 227
rect -1660 193 -1650 227
rect -1711 177 -1650 193
rect -1956 129 -1861 145
rect -2124 92 -2108 126
rect -2074 92 -2049 126
rect -2124 82 -2049 92
rect -2220 61 -2166 77
rect -2196 38 -2166 61
rect -2196 8 -2133 38
rect -2163 -7 -2133 8
rect -2079 -7 -2049 82
rect -1891 -7 -1861 129
rect -1819 149 -1753 159
rect -1819 115 -1803 149
rect -1769 135 -1753 149
rect -1769 115 -1650 135
rect -1819 105 -1650 115
rect -1799 53 -1733 63
rect -1799 19 -1783 53
rect -1749 19 -1733 53
rect -1799 9 -1733 19
rect -1779 -19 -1749 9
rect -1680 -19 -1650 105
rect -1608 75 -1578 275
rect -1476 171 -1446 209
rect -1381 177 -1351 275
rect -1297 237 -1267 275
rect -1183 243 -1153 275
rect -1298 227 -1232 237
rect -1298 193 -1282 227
rect -1248 193 -1232 227
rect -1298 183 -1232 193
rect -1183 227 -1102 243
rect -1183 193 -1146 227
rect -1112 193 -1102 227
rect -1183 177 -1102 193
rect -1536 161 -1446 171
rect -1536 127 -1520 161
rect -1486 127 -1446 161
rect -1536 117 -1446 127
rect -1476 82 -1446 117
rect -1394 161 -1340 177
rect -1394 127 -1384 161
rect -1350 141 -1340 161
rect -1350 127 -1225 141
rect -1394 111 -1225 127
rect -1608 65 -1534 75
rect -1608 31 -1584 65
rect -1550 31 -1534 65
rect -1476 52 -1432 82
rect -1462 37 -1432 52
rect -1361 53 -1297 69
rect -1608 21 -1534 31
rect -1581 -7 -1551 21
rect -1361 19 -1341 53
rect -1307 19 -1297 53
rect -1361 3 -1297 19
rect -1361 -19 -1331 3
rect -1255 -19 -1225 111
rect -1160 -7 -1130 177
rect -700 195 -670 231
rect -709 165 -670 195
rect -972 127 -942 159
rect -888 127 -858 159
rect -709 127 -679 165
rect -603 127 -573 159
rect -374 127 -344 159
rect -129 127 -99 159
rect -45 127 -15 159
rect 39 127 69 159
rect 123 127 153 159
rect -1082 111 -940 127
rect -1082 77 -1072 111
rect -1038 77 -940 111
rect -1082 61 -940 77
rect -898 111 -679 127
rect -898 77 -888 111
rect -854 77 -679 111
rect -898 61 -679 77
rect -637 111 -573 127
rect -637 77 -627 111
rect -593 77 -573 111
rect -637 61 -573 77
rect -430 111 -344 127
rect -430 77 -414 111
rect -380 77 -344 111
rect -430 61 -344 77
rect -197 111 153 127
rect -197 77 -181 111
rect -147 77 -89 111
rect -55 77 -5 111
rect 29 77 79 111
rect 113 77 153 111
rect -197 61 153 77
rect -970 39 -940 61
rect -886 39 -856 61
rect -709 32 -679 61
rect -603 39 -573 61
rect -374 39 -344 61
rect -129 39 -99 61
rect -45 39 -15 61
rect 39 39 69 61
rect 123 39 153 61
rect -709 8 -668 32
rect -698 -7 -668 8
rect -2163 -117 -2133 -91
rect -2079 -117 -2049 -91
rect -1891 -117 -1861 -91
rect -1779 -117 -1749 -91
rect -1680 -117 -1650 -91
rect -1581 -117 -1551 -91
rect -1462 -117 -1432 -91
rect -1361 -117 -1331 -91
rect -1255 -117 -1225 -91
rect -1160 -117 -1130 -91
rect -970 -117 -940 -91
rect -886 -117 -856 -91
rect -698 -117 -668 -91
rect -603 -117 -573 -91
rect -374 -117 -344 -91
rect -129 -117 -99 -91
rect -45 -117 -15 -91
rect 39 -117 69 -91
rect 123 -117 153 -91
rect -2163 -185 -2133 -159
rect -2079 -185 -2049 -159
rect -1891 -185 -1861 -159
rect -1779 -185 -1749 -159
rect -1680 -185 -1650 -159
rect -1581 -185 -1551 -159
rect -1462 -185 -1432 -159
rect -1361 -185 -1331 -159
rect -1255 -185 -1225 -159
rect -1160 -185 -1130 -159
rect -970 -185 -940 -159
rect -886 -185 -856 -159
rect -698 -185 -668 -159
rect -603 -185 -573 -159
rect -374 -185 -344 -159
rect -129 -185 -99 -159
rect -45 -185 -15 -159
rect 39 -185 69 -159
rect 123 -185 153 -159
rect 535 -185 565 -159
rect 619 -185 649 -159
rect 807 -185 837 -159
rect 919 -185 949 -159
rect 1018 -185 1048 -159
rect 1117 -185 1147 -159
rect 1236 -185 1266 -159
rect 1337 -185 1367 -159
rect 1443 -185 1473 -159
rect 1538 -185 1568 -159
rect 1728 -185 1758 -159
rect 1812 -185 1842 -159
rect 2000 -185 2030 -159
rect 2095 -185 2125 -159
rect 2324 -185 2354 -159
rect 2569 -185 2599 -159
rect 2653 -185 2683 -159
rect 2737 -185 2767 -159
rect 2821 -185 2851 -159
rect -2163 -284 -2133 -269
rect -2196 -314 -2133 -284
rect -2196 -337 -2166 -314
rect -2220 -353 -2166 -337
rect -2220 -387 -2210 -353
rect -2176 -387 -2166 -353
rect -2079 -358 -2049 -269
rect -2220 -403 -2166 -387
rect -2196 -456 -2166 -403
rect -2124 -368 -2049 -358
rect -2124 -402 -2108 -368
rect -2074 -402 -2049 -368
rect -2124 -412 -2049 -402
rect -1891 -405 -1861 -269
rect -1779 -285 -1749 -257
rect -1799 -295 -1733 -285
rect -1799 -329 -1783 -295
rect -1749 -329 -1733 -295
rect -1799 -339 -1733 -329
rect -1680 -381 -1650 -257
rect -1581 -297 -1551 -269
rect -2196 -486 -2133 -456
rect -2163 -501 -2133 -486
rect -2079 -501 -2049 -412
rect -1956 -421 -1861 -405
rect -1956 -455 -1946 -421
rect -1912 -455 -1861 -421
rect -1819 -391 -1650 -381
rect -1819 -425 -1803 -391
rect -1769 -411 -1650 -391
rect -1608 -307 -1534 -297
rect -1608 -341 -1584 -307
rect -1550 -341 -1534 -307
rect -1361 -279 -1331 -257
rect -1361 -295 -1297 -279
rect -1462 -328 -1432 -313
rect -1608 -351 -1534 -341
rect -1769 -425 -1753 -411
rect -1819 -435 -1753 -425
rect -1956 -471 -1861 -455
rect -1891 -551 -1861 -471
rect -1806 -551 -1776 -435
rect -1711 -469 -1650 -453
rect -1711 -503 -1694 -469
rect -1660 -503 -1650 -469
rect -1711 -519 -1650 -503
rect -1711 -551 -1681 -519
rect -1608 -551 -1578 -351
rect -1476 -358 -1432 -328
rect -1361 -329 -1341 -295
rect -1307 -329 -1297 -295
rect -1361 -345 -1297 -329
rect -1476 -393 -1446 -358
rect -1255 -387 -1225 -257
rect -1536 -403 -1446 -393
rect -1536 -437 -1520 -403
rect -1486 -437 -1446 -403
rect -1536 -447 -1446 -437
rect -1476 -485 -1446 -447
rect -1394 -403 -1225 -387
rect -1394 -437 -1384 -403
rect -1350 -417 -1225 -403
rect -1350 -437 -1340 -417
rect -1394 -453 -1340 -437
rect -1160 -453 -1130 -269
rect -698 -284 -668 -269
rect -709 -308 -668 -284
rect -970 -337 -940 -315
rect -886 -337 -856 -315
rect -709 -337 -679 -308
rect 535 -284 565 -269
rect 502 -314 565 -284
rect -603 -337 -573 -315
rect -374 -337 -344 -315
rect -129 -337 -99 -315
rect -45 -337 -15 -315
rect 39 -337 69 -315
rect 123 -337 153 -315
rect 502 -337 532 -314
rect -1082 -353 -940 -337
rect -1082 -387 -1072 -353
rect -1038 -387 -940 -353
rect -1082 -403 -940 -387
rect -898 -353 -679 -337
rect -898 -387 -888 -353
rect -854 -387 -679 -353
rect -898 -403 -679 -387
rect -637 -353 -573 -337
rect -637 -387 -627 -353
rect -593 -387 -573 -353
rect -637 -403 -573 -387
rect -430 -353 -344 -337
rect -430 -387 -414 -353
rect -380 -387 -344 -353
rect -430 -403 -344 -387
rect -197 -353 153 -337
rect -197 -387 -181 -353
rect -147 -387 -89 -353
rect -55 -387 -5 -353
rect 29 -387 79 -353
rect 113 -387 153 -353
rect -197 -403 153 -387
rect 478 -353 532 -337
rect 478 -387 488 -353
rect 522 -387 532 -353
rect 619 -358 649 -269
rect 478 -403 532 -387
rect -972 -435 -942 -403
rect -888 -435 -858 -403
rect -2163 -655 -2133 -629
rect -2079 -655 -2049 -629
rect -1381 -551 -1351 -453
rect -1298 -469 -1232 -459
rect -1298 -503 -1282 -469
rect -1248 -503 -1232 -469
rect -1298 -513 -1232 -503
rect -1183 -469 -1102 -453
rect -1183 -503 -1146 -469
rect -1112 -503 -1102 -469
rect -1297 -551 -1267 -513
rect -1183 -519 -1102 -503
rect -1183 -551 -1153 -519
rect -709 -441 -679 -403
rect -603 -435 -573 -403
rect -374 -435 -344 -403
rect -129 -435 -99 -403
rect -45 -435 -15 -403
rect 39 -435 69 -403
rect 123 -435 153 -403
rect -709 -471 -670 -441
rect -700 -507 -670 -471
rect 502 -456 532 -403
rect 574 -368 649 -358
rect 574 -402 590 -368
rect 624 -402 649 -368
rect 574 -412 649 -402
rect 807 -405 837 -269
rect 919 -285 949 -257
rect 899 -295 965 -285
rect 899 -329 915 -295
rect 949 -329 965 -295
rect 899 -339 965 -329
rect 1018 -381 1048 -257
rect 1117 -297 1147 -269
rect 502 -486 565 -456
rect 535 -501 565 -486
rect 619 -501 649 -412
rect 742 -421 837 -405
rect 742 -455 752 -421
rect 786 -455 837 -421
rect 879 -391 1048 -381
rect 879 -425 895 -391
rect 929 -411 1048 -391
rect 1090 -307 1164 -297
rect 1090 -341 1114 -307
rect 1148 -341 1164 -307
rect 1337 -279 1367 -257
rect 1337 -295 1401 -279
rect 1236 -328 1266 -313
rect 1090 -351 1164 -341
rect 929 -425 945 -411
rect 879 -435 945 -425
rect 742 -471 837 -455
rect 807 -551 837 -471
rect 892 -551 922 -435
rect 987 -469 1048 -453
rect 987 -503 1004 -469
rect 1038 -503 1048 -469
rect 987 -519 1048 -503
rect 987 -551 1017 -519
rect 1090 -551 1120 -351
rect 1222 -358 1266 -328
rect 1337 -329 1357 -295
rect 1391 -329 1401 -295
rect 1337 -345 1401 -329
rect 1222 -393 1252 -358
rect 1443 -387 1473 -257
rect 1162 -403 1252 -393
rect 1162 -437 1178 -403
rect 1212 -437 1252 -403
rect 1162 -447 1252 -437
rect 1222 -485 1252 -447
rect 1304 -403 1473 -387
rect 1304 -437 1314 -403
rect 1348 -417 1473 -403
rect 1348 -437 1358 -417
rect 1304 -453 1358 -437
rect 1538 -453 1568 -269
rect 2000 -284 2030 -269
rect 1989 -308 2030 -284
rect 1728 -337 1758 -315
rect 1812 -337 1842 -315
rect 1989 -337 2019 -308
rect 2095 -337 2125 -315
rect 2324 -337 2354 -315
rect 2569 -337 2599 -315
rect 2653 -337 2683 -315
rect 2737 -337 2767 -315
rect 2821 -337 2851 -315
rect 1616 -353 1758 -337
rect 1616 -387 1626 -353
rect 1660 -387 1758 -353
rect 1616 -403 1758 -387
rect 1800 -353 2019 -337
rect 1800 -387 1810 -353
rect 1844 -387 2019 -353
rect 1800 -403 2019 -387
rect 2061 -353 2125 -337
rect 2061 -387 2071 -353
rect 2105 -387 2125 -353
rect 2061 -403 2125 -387
rect 2268 -353 2354 -337
rect 2268 -387 2284 -353
rect 2318 -387 2354 -353
rect 2268 -403 2354 -387
rect 2501 -353 2851 -337
rect 2501 -387 2517 -353
rect 2551 -387 2609 -353
rect 2643 -387 2693 -353
rect 2727 -387 2777 -353
rect 2811 -387 2851 -353
rect 2501 -403 2851 -387
rect 1726 -435 1756 -403
rect 1810 -435 1840 -403
rect -1891 -661 -1861 -635
rect -1806 -661 -1776 -635
rect -1711 -661 -1681 -635
rect -1608 -661 -1578 -635
rect -1476 -661 -1446 -635
rect -1381 -661 -1351 -635
rect -1297 -661 -1267 -635
rect -1183 -661 -1153 -635
rect -972 -661 -942 -635
rect -888 -661 -858 -635
rect -700 -661 -670 -635
rect -603 -661 -573 -635
rect -374 -661 -344 -635
rect -129 -661 -99 -635
rect -45 -661 -15 -635
rect 39 -661 69 -635
rect 123 -661 153 -635
rect 535 -655 565 -629
rect 619 -655 649 -629
rect 1317 -551 1347 -453
rect 1400 -469 1466 -459
rect 1400 -503 1416 -469
rect 1450 -503 1466 -469
rect 1400 -513 1466 -503
rect 1515 -469 1596 -453
rect 1515 -503 1552 -469
rect 1586 -503 1596 -469
rect 1401 -551 1431 -513
rect 1515 -519 1596 -503
rect 1515 -551 1545 -519
rect 1989 -441 2019 -403
rect 2095 -435 2125 -403
rect 2324 -435 2354 -403
rect 2569 -435 2599 -403
rect 2653 -435 2683 -403
rect 2737 -435 2767 -403
rect 2821 -435 2851 -403
rect 1989 -471 2028 -441
rect 1998 -507 2028 -471
rect 807 -661 837 -635
rect 892 -661 922 -635
rect 987 -661 1017 -635
rect 1090 -661 1120 -635
rect 1222 -661 1252 -635
rect 1317 -661 1347 -635
rect 1401 -661 1431 -635
rect 1515 -661 1545 -635
rect 1726 -661 1756 -635
rect 1810 -661 1840 -635
rect 1998 -661 2028 -635
rect 2095 -661 2125 -635
rect 2324 -661 2354 -635
rect 2569 -661 2599 -635
rect 2653 -661 2683 -635
rect 2737 -661 2767 -635
rect 2821 -661 2851 -635
rect -2163 -735 -2133 -709
rect -2079 -735 -2049 -709
rect -1891 -729 -1861 -703
rect -1806 -729 -1776 -703
rect -1711 -729 -1681 -703
rect -1608 -729 -1578 -703
rect -1476 -729 -1446 -703
rect -1381 -729 -1351 -703
rect -1297 -729 -1267 -703
rect -1183 -729 -1153 -703
rect -972 -729 -942 -703
rect -888 -729 -858 -703
rect -700 -729 -670 -703
rect -603 -729 -573 -703
rect -374 -729 -344 -703
rect -129 -729 -99 -703
rect -45 -729 -15 -703
rect 39 -729 69 -703
rect 123 -729 153 -703
rect -2163 -878 -2133 -863
rect -2196 -908 -2133 -878
rect -2196 -961 -2166 -908
rect -2079 -952 -2049 -863
rect -1891 -893 -1861 -813
rect -2220 -977 -2166 -961
rect -2220 -1011 -2210 -977
rect -2176 -1011 -2166 -977
rect -2124 -962 -2049 -952
rect -1956 -909 -1861 -893
rect -1956 -943 -1946 -909
rect -1912 -943 -1861 -909
rect -1806 -929 -1776 -813
rect -1711 -845 -1681 -813
rect -1711 -861 -1650 -845
rect -1711 -895 -1694 -861
rect -1660 -895 -1650 -861
rect -1711 -911 -1650 -895
rect -1956 -959 -1861 -943
rect -2124 -996 -2108 -962
rect -2074 -996 -2049 -962
rect -2124 -1006 -2049 -996
rect -2220 -1027 -2166 -1011
rect -2196 -1050 -2166 -1027
rect -2196 -1080 -2133 -1050
rect -2163 -1095 -2133 -1080
rect -2079 -1095 -2049 -1006
rect -1891 -1095 -1861 -959
rect -1819 -939 -1753 -929
rect -1819 -973 -1803 -939
rect -1769 -953 -1753 -939
rect -1769 -973 -1650 -953
rect -1819 -983 -1650 -973
rect -1799 -1035 -1733 -1025
rect -1799 -1069 -1783 -1035
rect -1749 -1069 -1733 -1035
rect -1799 -1079 -1733 -1069
rect -1779 -1107 -1749 -1079
rect -1680 -1107 -1650 -983
rect -1608 -1013 -1578 -813
rect -1476 -917 -1446 -879
rect -1381 -911 -1351 -813
rect -1297 -851 -1267 -813
rect -1183 -845 -1153 -813
rect -1298 -861 -1232 -851
rect -1298 -895 -1282 -861
rect -1248 -895 -1232 -861
rect -1298 -905 -1232 -895
rect -1183 -861 -1102 -845
rect -1183 -895 -1146 -861
rect -1112 -895 -1102 -861
rect -1183 -911 -1102 -895
rect -1536 -927 -1446 -917
rect -1536 -961 -1520 -927
rect -1486 -961 -1446 -927
rect -1536 -971 -1446 -961
rect -1476 -1006 -1446 -971
rect -1394 -927 -1340 -911
rect -1394 -961 -1384 -927
rect -1350 -947 -1340 -927
rect -1350 -961 -1225 -947
rect -1394 -977 -1225 -961
rect -1608 -1023 -1534 -1013
rect -1608 -1057 -1584 -1023
rect -1550 -1057 -1534 -1023
rect -1476 -1036 -1432 -1006
rect -1462 -1051 -1432 -1036
rect -1361 -1035 -1297 -1019
rect -1608 -1067 -1534 -1057
rect -1581 -1095 -1551 -1067
rect -1361 -1069 -1341 -1035
rect -1307 -1069 -1297 -1035
rect -1361 -1085 -1297 -1069
rect -1361 -1107 -1331 -1085
rect -1255 -1107 -1225 -977
rect -1160 -1095 -1130 -911
rect -700 -893 -670 -857
rect -709 -923 -670 -893
rect -972 -961 -942 -929
rect -888 -961 -858 -929
rect -709 -961 -679 -923
rect 535 -735 565 -709
rect 619 -735 649 -709
rect 807 -729 837 -703
rect 892 -729 922 -703
rect 987 -729 1017 -703
rect 1090 -729 1120 -703
rect 1222 -729 1252 -703
rect 1317 -729 1347 -703
rect 1401 -729 1431 -703
rect 1515 -729 1545 -703
rect 1726 -729 1756 -703
rect 1810 -729 1840 -703
rect 1998 -729 2028 -703
rect 2095 -729 2125 -703
rect 2324 -729 2354 -703
rect 2569 -729 2599 -703
rect 2653 -729 2683 -703
rect 2737 -729 2767 -703
rect 2821 -729 2851 -703
rect 535 -878 565 -863
rect 502 -908 565 -878
rect -603 -961 -573 -929
rect -374 -961 -344 -929
rect -129 -961 -99 -929
rect -45 -961 -15 -929
rect 39 -961 69 -929
rect 123 -961 153 -929
rect 502 -961 532 -908
rect 619 -952 649 -863
rect 807 -893 837 -813
rect -1082 -977 -940 -961
rect -1082 -1011 -1072 -977
rect -1038 -1011 -940 -977
rect -1082 -1027 -940 -1011
rect -898 -977 -679 -961
rect -898 -1011 -888 -977
rect -854 -1011 -679 -977
rect -898 -1027 -679 -1011
rect -637 -977 -573 -961
rect -637 -1011 -627 -977
rect -593 -1011 -573 -977
rect -637 -1027 -573 -1011
rect -430 -977 -344 -961
rect -430 -1011 -414 -977
rect -380 -1011 -344 -977
rect -430 -1027 -344 -1011
rect -197 -977 153 -961
rect -197 -1011 -181 -977
rect -147 -1011 -89 -977
rect -55 -1011 -5 -977
rect 29 -1011 79 -977
rect 113 -1011 153 -977
rect -197 -1027 153 -1011
rect 478 -977 532 -961
rect 478 -1011 488 -977
rect 522 -1011 532 -977
rect 574 -962 649 -952
rect 742 -909 837 -893
rect 742 -943 752 -909
rect 786 -943 837 -909
rect 892 -929 922 -813
rect 987 -845 1017 -813
rect 987 -861 1048 -845
rect 987 -895 1004 -861
rect 1038 -895 1048 -861
rect 987 -911 1048 -895
rect 742 -959 837 -943
rect 574 -996 590 -962
rect 624 -996 649 -962
rect 574 -1006 649 -996
rect 478 -1027 532 -1011
rect -970 -1049 -940 -1027
rect -886 -1049 -856 -1027
rect -709 -1056 -679 -1027
rect -603 -1049 -573 -1027
rect -374 -1049 -344 -1027
rect -129 -1049 -99 -1027
rect -45 -1049 -15 -1027
rect 39 -1049 69 -1027
rect 123 -1049 153 -1027
rect -709 -1080 -668 -1056
rect -698 -1095 -668 -1080
rect 502 -1050 532 -1027
rect 502 -1080 565 -1050
rect 535 -1095 565 -1080
rect 619 -1095 649 -1006
rect 807 -1095 837 -959
rect 879 -939 945 -929
rect 879 -973 895 -939
rect 929 -953 945 -939
rect 929 -973 1048 -953
rect 879 -983 1048 -973
rect 899 -1035 965 -1025
rect 899 -1069 915 -1035
rect 949 -1069 965 -1035
rect 899 -1079 965 -1069
rect 919 -1107 949 -1079
rect 1018 -1107 1048 -983
rect 1090 -1013 1120 -813
rect 1222 -917 1252 -879
rect 1317 -911 1347 -813
rect 1401 -851 1431 -813
rect 1515 -845 1545 -813
rect 1400 -861 1466 -851
rect 1400 -895 1416 -861
rect 1450 -895 1466 -861
rect 1400 -905 1466 -895
rect 1515 -861 1596 -845
rect 1515 -895 1552 -861
rect 1586 -895 1596 -861
rect 1515 -911 1596 -895
rect 1162 -927 1252 -917
rect 1162 -961 1178 -927
rect 1212 -961 1252 -927
rect 1162 -971 1252 -961
rect 1222 -1006 1252 -971
rect 1304 -927 1358 -911
rect 1304 -961 1314 -927
rect 1348 -947 1358 -927
rect 1348 -961 1473 -947
rect 1304 -977 1473 -961
rect 1090 -1023 1164 -1013
rect 1090 -1057 1114 -1023
rect 1148 -1057 1164 -1023
rect 1222 -1036 1266 -1006
rect 1236 -1051 1266 -1036
rect 1337 -1035 1401 -1019
rect 1090 -1067 1164 -1057
rect 1117 -1095 1147 -1067
rect 1337 -1069 1357 -1035
rect 1391 -1069 1401 -1035
rect 1337 -1085 1401 -1069
rect 1337 -1107 1367 -1085
rect 1443 -1107 1473 -977
rect 1538 -1095 1568 -911
rect 1998 -893 2028 -857
rect 1989 -923 2028 -893
rect 1726 -961 1756 -929
rect 1810 -961 1840 -929
rect 1989 -961 2019 -923
rect 2095 -961 2125 -929
rect 2324 -961 2354 -929
rect 2569 -961 2599 -929
rect 2653 -961 2683 -929
rect 2737 -961 2767 -929
rect 2821 -961 2851 -929
rect 1616 -977 1758 -961
rect 1616 -1011 1626 -977
rect 1660 -1011 1758 -977
rect 1616 -1027 1758 -1011
rect 1800 -977 2019 -961
rect 1800 -1011 1810 -977
rect 1844 -1011 2019 -977
rect 1800 -1027 2019 -1011
rect 2061 -977 2125 -961
rect 2061 -1011 2071 -977
rect 2105 -1011 2125 -977
rect 2061 -1027 2125 -1011
rect 2268 -977 2354 -961
rect 2268 -1011 2284 -977
rect 2318 -1011 2354 -977
rect 2268 -1027 2354 -1011
rect 2501 -977 2851 -961
rect 2501 -1011 2517 -977
rect 2551 -1011 2609 -977
rect 2643 -1011 2693 -977
rect 2727 -1011 2777 -977
rect 2811 -1011 2851 -977
rect 2501 -1027 2851 -1011
rect 1728 -1049 1758 -1027
rect 1812 -1049 1842 -1027
rect 1989 -1056 2019 -1027
rect 2095 -1049 2125 -1027
rect 2324 -1049 2354 -1027
rect 2569 -1049 2599 -1027
rect 2653 -1049 2683 -1027
rect 2737 -1049 2767 -1027
rect 2821 -1049 2851 -1027
rect 1989 -1080 2030 -1056
rect 2000 -1095 2030 -1080
rect -2163 -1205 -2133 -1179
rect -2079 -1205 -2049 -1179
rect -1891 -1205 -1861 -1179
rect -1779 -1205 -1749 -1179
rect -1680 -1205 -1650 -1179
rect -1581 -1205 -1551 -1179
rect -1462 -1205 -1432 -1179
rect -1361 -1205 -1331 -1179
rect -1255 -1205 -1225 -1179
rect -1160 -1205 -1130 -1179
rect -970 -1205 -940 -1179
rect -886 -1205 -856 -1179
rect -698 -1205 -668 -1179
rect -603 -1205 -573 -1179
rect -374 -1205 -344 -1179
rect -129 -1205 -99 -1179
rect -45 -1205 -15 -1179
rect 39 -1205 69 -1179
rect 123 -1205 153 -1179
rect 535 -1205 565 -1179
rect 619 -1205 649 -1179
rect 807 -1205 837 -1179
rect 919 -1205 949 -1179
rect 1018 -1205 1048 -1179
rect 1117 -1205 1147 -1179
rect 1236 -1205 1266 -1179
rect 1337 -1205 1367 -1179
rect 1443 -1205 1473 -1179
rect 1538 -1205 1568 -1179
rect 1728 -1205 1758 -1179
rect 1812 -1205 1842 -1179
rect 2000 -1205 2030 -1179
rect 2095 -1205 2125 -1179
rect 2324 -1205 2354 -1179
rect 2569 -1205 2599 -1179
rect 2653 -1205 2683 -1179
rect 2737 -1205 2767 -1179
rect 2821 -1205 2851 -1179
rect -2163 -1273 -2133 -1247
rect -2079 -1273 -2049 -1247
rect -1891 -1273 -1861 -1247
rect -1779 -1273 -1749 -1247
rect -1680 -1273 -1650 -1247
rect -1581 -1273 -1551 -1247
rect -1462 -1273 -1432 -1247
rect -1361 -1273 -1331 -1247
rect -1255 -1273 -1225 -1247
rect -1160 -1273 -1130 -1247
rect -970 -1273 -940 -1247
rect -886 -1273 -856 -1247
rect -698 -1273 -668 -1247
rect -603 -1273 -573 -1247
rect -374 -1273 -344 -1247
rect -129 -1273 -99 -1247
rect -45 -1273 -15 -1247
rect 39 -1273 69 -1247
rect 123 -1273 153 -1247
rect 535 -1273 565 -1247
rect 619 -1273 649 -1247
rect 807 -1273 837 -1247
rect 919 -1273 949 -1247
rect 1018 -1273 1048 -1247
rect 1117 -1273 1147 -1247
rect 1236 -1273 1266 -1247
rect 1337 -1273 1367 -1247
rect 1443 -1273 1473 -1247
rect 1538 -1273 1568 -1247
rect 1728 -1273 1758 -1247
rect 1812 -1273 1842 -1247
rect 2000 -1273 2030 -1247
rect 2095 -1273 2125 -1247
rect 2324 -1273 2354 -1247
rect 2569 -1273 2599 -1247
rect 2653 -1273 2683 -1247
rect 2737 -1273 2767 -1247
rect 2821 -1273 2851 -1247
rect -2163 -1372 -2133 -1357
rect -2196 -1402 -2133 -1372
rect -2196 -1425 -2166 -1402
rect -2220 -1441 -2166 -1425
rect -2220 -1475 -2210 -1441
rect -2176 -1475 -2166 -1441
rect -2079 -1446 -2049 -1357
rect -2220 -1491 -2166 -1475
rect -2196 -1544 -2166 -1491
rect -2124 -1456 -2049 -1446
rect -2124 -1490 -2108 -1456
rect -2074 -1490 -2049 -1456
rect -2124 -1500 -2049 -1490
rect -1891 -1493 -1861 -1357
rect -1779 -1373 -1749 -1345
rect -1799 -1383 -1733 -1373
rect -1799 -1417 -1783 -1383
rect -1749 -1417 -1733 -1383
rect -1799 -1427 -1733 -1417
rect -1680 -1469 -1650 -1345
rect -1581 -1385 -1551 -1357
rect -2196 -1574 -2133 -1544
rect -2163 -1589 -2133 -1574
rect -2079 -1589 -2049 -1500
rect -1956 -1509 -1861 -1493
rect -1956 -1543 -1946 -1509
rect -1912 -1543 -1861 -1509
rect -1819 -1479 -1650 -1469
rect -1819 -1513 -1803 -1479
rect -1769 -1499 -1650 -1479
rect -1608 -1395 -1534 -1385
rect -1608 -1429 -1584 -1395
rect -1550 -1429 -1534 -1395
rect -1361 -1367 -1331 -1345
rect -1361 -1383 -1297 -1367
rect -1462 -1416 -1432 -1401
rect -1608 -1439 -1534 -1429
rect -1769 -1513 -1753 -1499
rect -1819 -1523 -1753 -1513
rect -1956 -1559 -1861 -1543
rect -1891 -1639 -1861 -1559
rect -1806 -1639 -1776 -1523
rect -1711 -1557 -1650 -1541
rect -1711 -1591 -1694 -1557
rect -1660 -1591 -1650 -1557
rect -1711 -1607 -1650 -1591
rect -1711 -1639 -1681 -1607
rect -1608 -1639 -1578 -1439
rect -1476 -1446 -1432 -1416
rect -1361 -1417 -1341 -1383
rect -1307 -1417 -1297 -1383
rect -1361 -1433 -1297 -1417
rect -1476 -1481 -1446 -1446
rect -1255 -1475 -1225 -1345
rect -1536 -1491 -1446 -1481
rect -1536 -1525 -1520 -1491
rect -1486 -1525 -1446 -1491
rect -1536 -1535 -1446 -1525
rect -1476 -1573 -1446 -1535
rect -1394 -1491 -1225 -1475
rect -1394 -1525 -1384 -1491
rect -1350 -1505 -1225 -1491
rect -1350 -1525 -1340 -1505
rect -1394 -1541 -1340 -1525
rect -1160 -1541 -1130 -1357
rect -698 -1372 -668 -1357
rect -709 -1396 -668 -1372
rect -970 -1425 -940 -1403
rect -886 -1425 -856 -1403
rect -709 -1425 -679 -1396
rect 535 -1372 565 -1357
rect 502 -1402 565 -1372
rect -603 -1425 -573 -1403
rect -374 -1425 -344 -1403
rect -129 -1425 -99 -1403
rect -45 -1425 -15 -1403
rect 39 -1425 69 -1403
rect 123 -1425 153 -1403
rect 502 -1425 532 -1402
rect -1082 -1441 -940 -1425
rect -1082 -1475 -1072 -1441
rect -1038 -1475 -940 -1441
rect -1082 -1491 -940 -1475
rect -898 -1441 -679 -1425
rect -898 -1475 -888 -1441
rect -854 -1475 -679 -1441
rect -898 -1491 -679 -1475
rect -637 -1441 -573 -1425
rect -637 -1475 -627 -1441
rect -593 -1475 -573 -1441
rect -637 -1491 -573 -1475
rect -430 -1441 -344 -1425
rect -430 -1475 -414 -1441
rect -380 -1475 -344 -1441
rect -430 -1491 -344 -1475
rect -197 -1441 153 -1425
rect -197 -1475 -181 -1441
rect -147 -1475 -89 -1441
rect -55 -1475 -5 -1441
rect 29 -1475 79 -1441
rect 113 -1475 153 -1441
rect -197 -1491 153 -1475
rect 478 -1441 532 -1425
rect 478 -1475 488 -1441
rect 522 -1475 532 -1441
rect 619 -1446 649 -1357
rect 478 -1491 532 -1475
rect -972 -1523 -942 -1491
rect -888 -1523 -858 -1491
rect -2163 -1743 -2133 -1717
rect -2079 -1743 -2049 -1717
rect -1381 -1639 -1351 -1541
rect -1298 -1557 -1232 -1547
rect -1298 -1591 -1282 -1557
rect -1248 -1591 -1232 -1557
rect -1298 -1601 -1232 -1591
rect -1183 -1557 -1102 -1541
rect -1183 -1591 -1146 -1557
rect -1112 -1591 -1102 -1557
rect -1297 -1639 -1267 -1601
rect -1183 -1607 -1102 -1591
rect -1183 -1639 -1153 -1607
rect -709 -1529 -679 -1491
rect -603 -1523 -573 -1491
rect -374 -1523 -344 -1491
rect -129 -1523 -99 -1491
rect -45 -1523 -15 -1491
rect 39 -1523 69 -1491
rect 123 -1523 153 -1491
rect -709 -1559 -670 -1529
rect -700 -1595 -670 -1559
rect 502 -1544 532 -1491
rect 574 -1456 649 -1446
rect 574 -1490 590 -1456
rect 624 -1490 649 -1456
rect 574 -1500 649 -1490
rect 807 -1493 837 -1357
rect 919 -1373 949 -1345
rect 899 -1383 965 -1373
rect 899 -1417 915 -1383
rect 949 -1417 965 -1383
rect 899 -1427 965 -1417
rect 1018 -1469 1048 -1345
rect 1117 -1385 1147 -1357
rect 502 -1574 565 -1544
rect 535 -1589 565 -1574
rect 619 -1589 649 -1500
rect 742 -1509 837 -1493
rect 742 -1543 752 -1509
rect 786 -1543 837 -1509
rect 879 -1479 1048 -1469
rect 879 -1513 895 -1479
rect 929 -1499 1048 -1479
rect 1090 -1395 1164 -1385
rect 1090 -1429 1114 -1395
rect 1148 -1429 1164 -1395
rect 1337 -1367 1367 -1345
rect 1337 -1383 1401 -1367
rect 1236 -1416 1266 -1401
rect 1090 -1439 1164 -1429
rect 929 -1513 945 -1499
rect 879 -1523 945 -1513
rect 742 -1559 837 -1543
rect 807 -1639 837 -1559
rect 892 -1639 922 -1523
rect 987 -1557 1048 -1541
rect 987 -1591 1004 -1557
rect 1038 -1591 1048 -1557
rect 987 -1607 1048 -1591
rect 987 -1639 1017 -1607
rect 1090 -1639 1120 -1439
rect 1222 -1446 1266 -1416
rect 1337 -1417 1357 -1383
rect 1391 -1417 1401 -1383
rect 1337 -1433 1401 -1417
rect 1222 -1481 1252 -1446
rect 1443 -1475 1473 -1345
rect 1162 -1491 1252 -1481
rect 1162 -1525 1178 -1491
rect 1212 -1525 1252 -1491
rect 1162 -1535 1252 -1525
rect 1222 -1573 1252 -1535
rect 1304 -1491 1473 -1475
rect 1304 -1525 1314 -1491
rect 1348 -1505 1473 -1491
rect 1348 -1525 1358 -1505
rect 1304 -1541 1358 -1525
rect 1538 -1541 1568 -1357
rect 2000 -1372 2030 -1357
rect 1989 -1396 2030 -1372
rect 1728 -1425 1758 -1403
rect 1812 -1425 1842 -1403
rect 1989 -1425 2019 -1396
rect 2095 -1425 2125 -1403
rect 2324 -1425 2354 -1403
rect 2569 -1425 2599 -1403
rect 2653 -1425 2683 -1403
rect 2737 -1425 2767 -1403
rect 2821 -1425 2851 -1403
rect 1616 -1441 1758 -1425
rect 1616 -1475 1626 -1441
rect 1660 -1475 1758 -1441
rect 1616 -1491 1758 -1475
rect 1800 -1441 2019 -1425
rect 1800 -1475 1810 -1441
rect 1844 -1475 2019 -1441
rect 1800 -1491 2019 -1475
rect 2061 -1441 2125 -1425
rect 2061 -1475 2071 -1441
rect 2105 -1475 2125 -1441
rect 2061 -1491 2125 -1475
rect 2268 -1441 2354 -1425
rect 2268 -1475 2284 -1441
rect 2318 -1475 2354 -1441
rect 2268 -1491 2354 -1475
rect 2501 -1441 2851 -1425
rect 2501 -1475 2517 -1441
rect 2551 -1475 2609 -1441
rect 2643 -1475 2693 -1441
rect 2727 -1475 2777 -1441
rect 2811 -1475 2851 -1441
rect 2501 -1491 2851 -1475
rect 1726 -1523 1756 -1491
rect 1810 -1523 1840 -1491
rect -1891 -1749 -1861 -1723
rect -1806 -1749 -1776 -1723
rect -1711 -1749 -1681 -1723
rect -1608 -1749 -1578 -1723
rect -1476 -1749 -1446 -1723
rect -1381 -1749 -1351 -1723
rect -1297 -1749 -1267 -1723
rect -1183 -1749 -1153 -1723
rect -972 -1749 -942 -1723
rect -888 -1749 -858 -1723
rect -700 -1749 -670 -1723
rect -603 -1749 -573 -1723
rect -374 -1749 -344 -1723
rect -129 -1749 -99 -1723
rect -45 -1749 -15 -1723
rect 39 -1749 69 -1723
rect 123 -1749 153 -1723
rect 535 -1743 565 -1717
rect 619 -1743 649 -1717
rect 1317 -1639 1347 -1541
rect 1400 -1557 1466 -1547
rect 1400 -1591 1416 -1557
rect 1450 -1591 1466 -1557
rect 1400 -1601 1466 -1591
rect 1515 -1557 1596 -1541
rect 1515 -1591 1552 -1557
rect 1586 -1591 1596 -1557
rect 1401 -1639 1431 -1601
rect 1515 -1607 1596 -1591
rect 1515 -1639 1545 -1607
rect 1989 -1529 2019 -1491
rect 2095 -1523 2125 -1491
rect 2324 -1523 2354 -1491
rect 2569 -1523 2599 -1491
rect 2653 -1523 2683 -1491
rect 2737 -1523 2767 -1491
rect 2821 -1523 2851 -1491
rect 1989 -1559 2028 -1529
rect 1998 -1595 2028 -1559
rect 807 -1749 837 -1723
rect 892 -1749 922 -1723
rect 987 -1749 1017 -1723
rect 1090 -1749 1120 -1723
rect 1222 -1749 1252 -1723
rect 1317 -1749 1347 -1723
rect 1401 -1749 1431 -1723
rect 1515 -1749 1545 -1723
rect 1726 -1749 1756 -1723
rect 1810 -1749 1840 -1723
rect 1998 -1749 2028 -1723
rect 2095 -1749 2125 -1723
rect 2324 -1749 2354 -1723
rect 2569 -1749 2599 -1723
rect 2653 -1749 2683 -1723
rect 2737 -1749 2767 -1723
rect 2821 -1749 2851 -1723
rect -2163 -1823 -2133 -1797
rect -2079 -1823 -2049 -1797
rect -1891 -1817 -1861 -1791
rect -1806 -1817 -1776 -1791
rect -1711 -1817 -1681 -1791
rect -1608 -1817 -1578 -1791
rect -1476 -1817 -1446 -1791
rect -1381 -1817 -1351 -1791
rect -1297 -1817 -1267 -1791
rect -1183 -1817 -1153 -1791
rect -972 -1817 -942 -1791
rect -888 -1817 -858 -1791
rect -700 -1817 -670 -1791
rect -603 -1817 -573 -1791
rect -374 -1817 -344 -1791
rect -129 -1817 -99 -1791
rect -45 -1817 -15 -1791
rect 39 -1817 69 -1791
rect 123 -1817 153 -1791
rect -2163 -1966 -2133 -1951
rect -2196 -1996 -2133 -1966
rect -2196 -2049 -2166 -1996
rect -2079 -2040 -2049 -1951
rect -1891 -1981 -1861 -1901
rect -2220 -2065 -2166 -2049
rect -2220 -2099 -2210 -2065
rect -2176 -2099 -2166 -2065
rect -2124 -2050 -2049 -2040
rect -1956 -1997 -1861 -1981
rect -1956 -2031 -1946 -1997
rect -1912 -2031 -1861 -1997
rect -1806 -2017 -1776 -1901
rect -1711 -1933 -1681 -1901
rect -1711 -1949 -1650 -1933
rect -1711 -1983 -1694 -1949
rect -1660 -1983 -1650 -1949
rect -1711 -1999 -1650 -1983
rect -1956 -2047 -1861 -2031
rect -2124 -2084 -2108 -2050
rect -2074 -2084 -2049 -2050
rect -2124 -2094 -2049 -2084
rect -2220 -2115 -2166 -2099
rect -2196 -2138 -2166 -2115
rect -2196 -2168 -2133 -2138
rect -2163 -2183 -2133 -2168
rect -2079 -2183 -2049 -2094
rect -1891 -2183 -1861 -2047
rect -1819 -2027 -1753 -2017
rect -1819 -2061 -1803 -2027
rect -1769 -2041 -1753 -2027
rect -1769 -2061 -1650 -2041
rect -1819 -2071 -1650 -2061
rect -1799 -2123 -1733 -2113
rect -1799 -2157 -1783 -2123
rect -1749 -2157 -1733 -2123
rect -1799 -2167 -1733 -2157
rect -1779 -2195 -1749 -2167
rect -1680 -2195 -1650 -2071
rect -1608 -2101 -1578 -1901
rect -1476 -2005 -1446 -1967
rect -1381 -1999 -1351 -1901
rect -1297 -1939 -1267 -1901
rect -1183 -1933 -1153 -1901
rect -1298 -1949 -1232 -1939
rect -1298 -1983 -1282 -1949
rect -1248 -1983 -1232 -1949
rect -1298 -1993 -1232 -1983
rect -1183 -1949 -1102 -1933
rect -1183 -1983 -1146 -1949
rect -1112 -1983 -1102 -1949
rect -1183 -1999 -1102 -1983
rect -1536 -2015 -1446 -2005
rect -1536 -2049 -1520 -2015
rect -1486 -2049 -1446 -2015
rect -1536 -2059 -1446 -2049
rect -1476 -2094 -1446 -2059
rect -1394 -2015 -1340 -1999
rect -1394 -2049 -1384 -2015
rect -1350 -2035 -1340 -2015
rect -1350 -2049 -1225 -2035
rect -1394 -2065 -1225 -2049
rect -1608 -2111 -1534 -2101
rect -1608 -2145 -1584 -2111
rect -1550 -2145 -1534 -2111
rect -1476 -2124 -1432 -2094
rect -1462 -2139 -1432 -2124
rect -1361 -2123 -1297 -2107
rect -1608 -2155 -1534 -2145
rect -1581 -2183 -1551 -2155
rect -1361 -2157 -1341 -2123
rect -1307 -2157 -1297 -2123
rect -1361 -2173 -1297 -2157
rect -1361 -2195 -1331 -2173
rect -1255 -2195 -1225 -2065
rect -1160 -2183 -1130 -1999
rect -700 -1981 -670 -1945
rect -709 -2011 -670 -1981
rect -972 -2049 -942 -2017
rect -888 -2049 -858 -2017
rect -709 -2049 -679 -2011
rect 535 -1823 565 -1797
rect 619 -1823 649 -1797
rect 807 -1817 837 -1791
rect 892 -1817 922 -1791
rect 987 -1817 1017 -1791
rect 1090 -1817 1120 -1791
rect 1222 -1817 1252 -1791
rect 1317 -1817 1347 -1791
rect 1401 -1817 1431 -1791
rect 1515 -1817 1545 -1791
rect 1726 -1817 1756 -1791
rect 1810 -1817 1840 -1791
rect 1998 -1817 2028 -1791
rect 2095 -1817 2125 -1791
rect 2324 -1817 2354 -1791
rect 2569 -1817 2599 -1791
rect 2653 -1817 2683 -1791
rect 2737 -1817 2767 -1791
rect 2821 -1817 2851 -1791
rect 535 -1966 565 -1951
rect 502 -1996 565 -1966
rect -603 -2049 -573 -2017
rect -374 -2049 -344 -2017
rect -129 -2049 -99 -2017
rect -45 -2049 -15 -2017
rect 39 -2049 69 -2017
rect 123 -2049 153 -2017
rect 502 -2049 532 -1996
rect 619 -2040 649 -1951
rect 807 -1981 837 -1901
rect -1082 -2065 -940 -2049
rect -1082 -2099 -1072 -2065
rect -1038 -2099 -940 -2065
rect -1082 -2115 -940 -2099
rect -898 -2065 -679 -2049
rect -898 -2099 -888 -2065
rect -854 -2099 -679 -2065
rect -898 -2115 -679 -2099
rect -637 -2065 -573 -2049
rect -637 -2099 -627 -2065
rect -593 -2099 -573 -2065
rect -637 -2115 -573 -2099
rect -430 -2065 -344 -2049
rect -430 -2099 -414 -2065
rect -380 -2099 -344 -2065
rect -430 -2115 -344 -2099
rect -197 -2065 153 -2049
rect -197 -2099 -181 -2065
rect -147 -2099 -89 -2065
rect -55 -2099 -5 -2065
rect 29 -2099 79 -2065
rect 113 -2099 153 -2065
rect -197 -2115 153 -2099
rect 478 -2065 532 -2049
rect 478 -2099 488 -2065
rect 522 -2099 532 -2065
rect 574 -2050 649 -2040
rect 742 -1997 837 -1981
rect 742 -2031 752 -1997
rect 786 -2031 837 -1997
rect 892 -2017 922 -1901
rect 987 -1933 1017 -1901
rect 987 -1949 1048 -1933
rect 987 -1983 1004 -1949
rect 1038 -1983 1048 -1949
rect 987 -1999 1048 -1983
rect 742 -2047 837 -2031
rect 574 -2084 590 -2050
rect 624 -2084 649 -2050
rect 574 -2094 649 -2084
rect 478 -2115 532 -2099
rect -970 -2137 -940 -2115
rect -886 -2137 -856 -2115
rect -709 -2144 -679 -2115
rect -603 -2137 -573 -2115
rect -374 -2137 -344 -2115
rect -129 -2137 -99 -2115
rect -45 -2137 -15 -2115
rect 39 -2137 69 -2115
rect 123 -2137 153 -2115
rect -709 -2168 -668 -2144
rect -698 -2183 -668 -2168
rect 502 -2138 532 -2115
rect 502 -2168 565 -2138
rect 535 -2183 565 -2168
rect 619 -2183 649 -2094
rect 807 -2183 837 -2047
rect 879 -2027 945 -2017
rect 879 -2061 895 -2027
rect 929 -2041 945 -2027
rect 929 -2061 1048 -2041
rect 879 -2071 1048 -2061
rect 899 -2123 965 -2113
rect 899 -2157 915 -2123
rect 949 -2157 965 -2123
rect 899 -2167 965 -2157
rect 919 -2195 949 -2167
rect 1018 -2195 1048 -2071
rect 1090 -2101 1120 -1901
rect 1222 -2005 1252 -1967
rect 1317 -1999 1347 -1901
rect 1401 -1939 1431 -1901
rect 1515 -1933 1545 -1901
rect 1400 -1949 1466 -1939
rect 1400 -1983 1416 -1949
rect 1450 -1983 1466 -1949
rect 1400 -1993 1466 -1983
rect 1515 -1949 1596 -1933
rect 1515 -1983 1552 -1949
rect 1586 -1983 1596 -1949
rect 1515 -1999 1596 -1983
rect 1162 -2015 1252 -2005
rect 1162 -2049 1178 -2015
rect 1212 -2049 1252 -2015
rect 1162 -2059 1252 -2049
rect 1222 -2094 1252 -2059
rect 1304 -2015 1358 -1999
rect 1304 -2049 1314 -2015
rect 1348 -2035 1358 -2015
rect 1348 -2049 1473 -2035
rect 1304 -2065 1473 -2049
rect 1090 -2111 1164 -2101
rect 1090 -2145 1114 -2111
rect 1148 -2145 1164 -2111
rect 1222 -2124 1266 -2094
rect 1236 -2139 1266 -2124
rect 1337 -2123 1401 -2107
rect 1090 -2155 1164 -2145
rect 1117 -2183 1147 -2155
rect 1337 -2157 1357 -2123
rect 1391 -2157 1401 -2123
rect 1337 -2173 1401 -2157
rect 1337 -2195 1367 -2173
rect 1443 -2195 1473 -2065
rect 1538 -2183 1568 -1999
rect 1998 -1981 2028 -1945
rect 1989 -2011 2028 -1981
rect 1726 -2049 1756 -2017
rect 1810 -2049 1840 -2017
rect 1989 -2049 2019 -2011
rect 2095 -2049 2125 -2017
rect 2324 -2049 2354 -2017
rect 2569 -2049 2599 -2017
rect 2653 -2049 2683 -2017
rect 2737 -2049 2767 -2017
rect 2821 -2049 2851 -2017
rect 1616 -2065 1758 -2049
rect 1616 -2099 1626 -2065
rect 1660 -2099 1758 -2065
rect 1616 -2115 1758 -2099
rect 1800 -2065 2019 -2049
rect 1800 -2099 1810 -2065
rect 1844 -2099 2019 -2065
rect 1800 -2115 2019 -2099
rect 2061 -2065 2125 -2049
rect 2061 -2099 2071 -2065
rect 2105 -2099 2125 -2065
rect 2061 -2115 2125 -2099
rect 2268 -2065 2354 -2049
rect 2268 -2099 2284 -2065
rect 2318 -2099 2354 -2065
rect 2268 -2115 2354 -2099
rect 2501 -2065 2851 -2049
rect 2501 -2099 2517 -2065
rect 2551 -2099 2609 -2065
rect 2643 -2099 2693 -2065
rect 2727 -2099 2777 -2065
rect 2811 -2099 2851 -2065
rect 2501 -2115 2851 -2099
rect 1728 -2137 1758 -2115
rect 1812 -2137 1842 -2115
rect 1989 -2144 2019 -2115
rect 2095 -2137 2125 -2115
rect 2324 -2137 2354 -2115
rect 2569 -2137 2599 -2115
rect 2653 -2137 2683 -2115
rect 2737 -2137 2767 -2115
rect 2821 -2137 2851 -2115
rect 1989 -2168 2030 -2144
rect 2000 -2183 2030 -2168
rect -2163 -2293 -2133 -2267
rect -2079 -2293 -2049 -2267
rect -1891 -2293 -1861 -2267
rect -1779 -2293 -1749 -2267
rect -1680 -2293 -1650 -2267
rect -1581 -2293 -1551 -2267
rect -1462 -2293 -1432 -2267
rect -1361 -2293 -1331 -2267
rect -1255 -2293 -1225 -2267
rect -1160 -2293 -1130 -2267
rect -970 -2293 -940 -2267
rect -886 -2293 -856 -2267
rect -698 -2293 -668 -2267
rect -603 -2293 -573 -2267
rect -374 -2293 -344 -2267
rect -129 -2293 -99 -2267
rect -45 -2293 -15 -2267
rect 39 -2293 69 -2267
rect 123 -2293 153 -2267
rect 535 -2293 565 -2267
rect 619 -2293 649 -2267
rect 807 -2293 837 -2267
rect 919 -2293 949 -2267
rect 1018 -2293 1048 -2267
rect 1117 -2293 1147 -2267
rect 1236 -2293 1266 -2267
rect 1337 -2293 1367 -2267
rect 1443 -2293 1473 -2267
rect 1538 -2293 1568 -2267
rect 1728 -2293 1758 -2267
rect 1812 -2293 1842 -2267
rect 2000 -2293 2030 -2267
rect 2095 -2293 2125 -2267
rect 2324 -2293 2354 -2267
rect 2569 -2293 2599 -2267
rect 2653 -2293 2683 -2267
rect 2737 -2293 2767 -2267
rect 2821 -2293 2851 -2267
rect -2163 -2361 -2133 -2335
rect -2079 -2361 -2049 -2335
rect -1891 -2361 -1861 -2335
rect -1779 -2361 -1749 -2335
rect -1680 -2361 -1650 -2335
rect -1581 -2361 -1551 -2335
rect -1462 -2361 -1432 -2335
rect -1361 -2361 -1331 -2335
rect -1255 -2361 -1225 -2335
rect -1160 -2361 -1130 -2335
rect -970 -2361 -940 -2335
rect -886 -2361 -856 -2335
rect -698 -2361 -668 -2335
rect -603 -2361 -573 -2335
rect -374 -2361 -344 -2335
rect -129 -2361 -99 -2335
rect -45 -2361 -15 -2335
rect 39 -2361 69 -2335
rect 123 -2361 153 -2335
rect 535 -2361 565 -2335
rect 619 -2361 649 -2335
rect 807 -2361 837 -2335
rect 919 -2361 949 -2335
rect 1018 -2361 1048 -2335
rect 1117 -2361 1147 -2335
rect 1236 -2361 1266 -2335
rect 1337 -2361 1367 -2335
rect 1443 -2361 1473 -2335
rect 1538 -2361 1568 -2335
rect 1728 -2361 1758 -2335
rect 1812 -2361 1842 -2335
rect 2000 -2361 2030 -2335
rect 2095 -2361 2125 -2335
rect 2324 -2361 2354 -2335
rect 2569 -2361 2599 -2335
rect 2653 -2361 2683 -2335
rect 2737 -2361 2767 -2335
rect 2821 -2361 2851 -2335
rect -2163 -2460 -2133 -2445
rect -2196 -2490 -2133 -2460
rect -2196 -2513 -2166 -2490
rect -2220 -2529 -2166 -2513
rect -2220 -2563 -2210 -2529
rect -2176 -2563 -2166 -2529
rect -2079 -2534 -2049 -2445
rect -2220 -2579 -2166 -2563
rect -2196 -2632 -2166 -2579
rect -2124 -2544 -2049 -2534
rect -2124 -2578 -2108 -2544
rect -2074 -2578 -2049 -2544
rect -2124 -2588 -2049 -2578
rect -1891 -2581 -1861 -2445
rect -1779 -2461 -1749 -2433
rect -1799 -2471 -1733 -2461
rect -1799 -2505 -1783 -2471
rect -1749 -2505 -1733 -2471
rect -1799 -2515 -1733 -2505
rect -1680 -2557 -1650 -2433
rect -1581 -2473 -1551 -2445
rect -2196 -2662 -2133 -2632
rect -2163 -2677 -2133 -2662
rect -2079 -2677 -2049 -2588
rect -1956 -2597 -1861 -2581
rect -1956 -2631 -1946 -2597
rect -1912 -2631 -1861 -2597
rect -1819 -2567 -1650 -2557
rect -1819 -2601 -1803 -2567
rect -1769 -2587 -1650 -2567
rect -1608 -2483 -1534 -2473
rect -1608 -2517 -1584 -2483
rect -1550 -2517 -1534 -2483
rect -1361 -2455 -1331 -2433
rect -1361 -2471 -1297 -2455
rect -1462 -2504 -1432 -2489
rect -1608 -2527 -1534 -2517
rect -1769 -2601 -1753 -2587
rect -1819 -2611 -1753 -2601
rect -1956 -2647 -1861 -2631
rect -1891 -2727 -1861 -2647
rect -1806 -2727 -1776 -2611
rect -1711 -2645 -1650 -2629
rect -1711 -2679 -1694 -2645
rect -1660 -2679 -1650 -2645
rect -1711 -2695 -1650 -2679
rect -1711 -2727 -1681 -2695
rect -1608 -2727 -1578 -2527
rect -1476 -2534 -1432 -2504
rect -1361 -2505 -1341 -2471
rect -1307 -2505 -1297 -2471
rect -1361 -2521 -1297 -2505
rect -1476 -2569 -1446 -2534
rect -1255 -2563 -1225 -2433
rect -1536 -2579 -1446 -2569
rect -1536 -2613 -1520 -2579
rect -1486 -2613 -1446 -2579
rect -1536 -2623 -1446 -2613
rect -1476 -2661 -1446 -2623
rect -1394 -2579 -1225 -2563
rect -1394 -2613 -1384 -2579
rect -1350 -2593 -1225 -2579
rect -1350 -2613 -1340 -2593
rect -1394 -2629 -1340 -2613
rect -1160 -2629 -1130 -2445
rect -698 -2460 -668 -2445
rect -709 -2484 -668 -2460
rect -970 -2513 -940 -2491
rect -886 -2513 -856 -2491
rect -709 -2513 -679 -2484
rect 535 -2460 565 -2445
rect 502 -2490 565 -2460
rect -603 -2513 -573 -2491
rect -374 -2513 -344 -2491
rect -129 -2513 -99 -2491
rect -45 -2513 -15 -2491
rect 39 -2513 69 -2491
rect 123 -2513 153 -2491
rect 502 -2513 532 -2490
rect -1082 -2529 -940 -2513
rect -1082 -2563 -1072 -2529
rect -1038 -2563 -940 -2529
rect -1082 -2579 -940 -2563
rect -898 -2529 -679 -2513
rect -898 -2563 -888 -2529
rect -854 -2563 -679 -2529
rect -898 -2579 -679 -2563
rect -637 -2529 -573 -2513
rect -637 -2563 -627 -2529
rect -593 -2563 -573 -2529
rect -637 -2579 -573 -2563
rect -430 -2529 -344 -2513
rect -430 -2563 -414 -2529
rect -380 -2563 -344 -2529
rect -430 -2579 -344 -2563
rect -197 -2529 153 -2513
rect -197 -2563 -181 -2529
rect -147 -2563 -89 -2529
rect -55 -2563 -5 -2529
rect 29 -2563 79 -2529
rect 113 -2563 153 -2529
rect -197 -2579 153 -2563
rect 478 -2529 532 -2513
rect 478 -2563 488 -2529
rect 522 -2563 532 -2529
rect 619 -2534 649 -2445
rect 478 -2579 532 -2563
rect -972 -2611 -942 -2579
rect -888 -2611 -858 -2579
rect -2163 -2831 -2133 -2805
rect -2079 -2831 -2049 -2805
rect -1381 -2727 -1351 -2629
rect -1298 -2645 -1232 -2635
rect -1298 -2679 -1282 -2645
rect -1248 -2679 -1232 -2645
rect -1298 -2689 -1232 -2679
rect -1183 -2645 -1102 -2629
rect -1183 -2679 -1146 -2645
rect -1112 -2679 -1102 -2645
rect -1297 -2727 -1267 -2689
rect -1183 -2695 -1102 -2679
rect -1183 -2727 -1153 -2695
rect -709 -2617 -679 -2579
rect -603 -2611 -573 -2579
rect -374 -2611 -344 -2579
rect -129 -2611 -99 -2579
rect -45 -2611 -15 -2579
rect 39 -2611 69 -2579
rect 123 -2611 153 -2579
rect -709 -2647 -670 -2617
rect -700 -2683 -670 -2647
rect 502 -2632 532 -2579
rect 574 -2544 649 -2534
rect 574 -2578 590 -2544
rect 624 -2578 649 -2544
rect 574 -2588 649 -2578
rect 807 -2581 837 -2445
rect 919 -2461 949 -2433
rect 899 -2471 965 -2461
rect 899 -2505 915 -2471
rect 949 -2505 965 -2471
rect 899 -2515 965 -2505
rect 1018 -2557 1048 -2433
rect 1117 -2473 1147 -2445
rect 502 -2662 565 -2632
rect 535 -2677 565 -2662
rect 619 -2677 649 -2588
rect 742 -2597 837 -2581
rect 742 -2631 752 -2597
rect 786 -2631 837 -2597
rect 879 -2567 1048 -2557
rect 879 -2601 895 -2567
rect 929 -2587 1048 -2567
rect 1090 -2483 1164 -2473
rect 1090 -2517 1114 -2483
rect 1148 -2517 1164 -2483
rect 1337 -2455 1367 -2433
rect 1337 -2471 1401 -2455
rect 1236 -2504 1266 -2489
rect 1090 -2527 1164 -2517
rect 929 -2601 945 -2587
rect 879 -2611 945 -2601
rect 742 -2647 837 -2631
rect 807 -2727 837 -2647
rect 892 -2727 922 -2611
rect 987 -2645 1048 -2629
rect 987 -2679 1004 -2645
rect 1038 -2679 1048 -2645
rect 987 -2695 1048 -2679
rect 987 -2727 1017 -2695
rect 1090 -2727 1120 -2527
rect 1222 -2534 1266 -2504
rect 1337 -2505 1357 -2471
rect 1391 -2505 1401 -2471
rect 1337 -2521 1401 -2505
rect 1222 -2569 1252 -2534
rect 1443 -2563 1473 -2433
rect 1162 -2579 1252 -2569
rect 1162 -2613 1178 -2579
rect 1212 -2613 1252 -2579
rect 1162 -2623 1252 -2613
rect 1222 -2661 1252 -2623
rect 1304 -2579 1473 -2563
rect 1304 -2613 1314 -2579
rect 1348 -2593 1473 -2579
rect 1348 -2613 1358 -2593
rect 1304 -2629 1358 -2613
rect 1538 -2629 1568 -2445
rect 2000 -2460 2030 -2445
rect 1989 -2484 2030 -2460
rect 1728 -2513 1758 -2491
rect 1812 -2513 1842 -2491
rect 1989 -2513 2019 -2484
rect 2095 -2513 2125 -2491
rect 2324 -2513 2354 -2491
rect 2569 -2513 2599 -2491
rect 2653 -2513 2683 -2491
rect 2737 -2513 2767 -2491
rect 2821 -2513 2851 -2491
rect 1616 -2529 1758 -2513
rect 1616 -2563 1626 -2529
rect 1660 -2563 1758 -2529
rect 1616 -2579 1758 -2563
rect 1800 -2529 2019 -2513
rect 1800 -2563 1810 -2529
rect 1844 -2563 2019 -2529
rect 1800 -2579 2019 -2563
rect 2061 -2529 2125 -2513
rect 2061 -2563 2071 -2529
rect 2105 -2563 2125 -2529
rect 2061 -2579 2125 -2563
rect 2268 -2529 2354 -2513
rect 2268 -2563 2284 -2529
rect 2318 -2563 2354 -2529
rect 2268 -2579 2354 -2563
rect 2501 -2529 2851 -2513
rect 2501 -2563 2517 -2529
rect 2551 -2563 2609 -2529
rect 2643 -2563 2693 -2529
rect 2727 -2563 2777 -2529
rect 2811 -2563 2851 -2529
rect 2501 -2579 2851 -2563
rect 1726 -2611 1756 -2579
rect 1810 -2611 1840 -2579
rect -1891 -2837 -1861 -2811
rect -1806 -2837 -1776 -2811
rect -1711 -2837 -1681 -2811
rect -1608 -2837 -1578 -2811
rect -1476 -2837 -1446 -2811
rect -1381 -2837 -1351 -2811
rect -1297 -2837 -1267 -2811
rect -1183 -2837 -1153 -2811
rect -972 -2837 -942 -2811
rect -888 -2837 -858 -2811
rect -700 -2837 -670 -2811
rect -603 -2837 -573 -2811
rect -374 -2837 -344 -2811
rect -129 -2837 -99 -2811
rect -45 -2837 -15 -2811
rect 39 -2837 69 -2811
rect 123 -2837 153 -2811
rect 535 -2831 565 -2805
rect 619 -2831 649 -2805
rect 1317 -2727 1347 -2629
rect 1400 -2645 1466 -2635
rect 1400 -2679 1416 -2645
rect 1450 -2679 1466 -2645
rect 1400 -2689 1466 -2679
rect 1515 -2645 1596 -2629
rect 1515 -2679 1552 -2645
rect 1586 -2679 1596 -2645
rect 1401 -2727 1431 -2689
rect 1515 -2695 1596 -2679
rect 1515 -2727 1545 -2695
rect 1989 -2617 2019 -2579
rect 2095 -2611 2125 -2579
rect 2324 -2611 2354 -2579
rect 2569 -2611 2599 -2579
rect 2653 -2611 2683 -2579
rect 2737 -2611 2767 -2579
rect 2821 -2611 2851 -2579
rect 1989 -2647 2028 -2617
rect 1998 -2683 2028 -2647
rect 807 -2837 837 -2811
rect 892 -2837 922 -2811
rect 987 -2837 1017 -2811
rect 1090 -2837 1120 -2811
rect 1222 -2837 1252 -2811
rect 1317 -2837 1347 -2811
rect 1401 -2837 1431 -2811
rect 1515 -2837 1545 -2811
rect 1726 -2837 1756 -2811
rect 1810 -2837 1840 -2811
rect 1998 -2837 2028 -2811
rect 2095 -2837 2125 -2811
rect 2324 -2837 2354 -2811
rect 2569 -2837 2599 -2811
rect 2653 -2837 2683 -2811
rect 2737 -2837 2767 -2811
rect 2821 -2837 2851 -2811
<< polycont >>
rect -2210 77 -2176 111
rect -1946 145 -1912 179
rect -1694 193 -1660 227
rect -2108 92 -2074 126
rect -1803 115 -1769 149
rect -1783 19 -1749 53
rect -1282 193 -1248 227
rect -1146 193 -1112 227
rect -1520 127 -1486 161
rect -1384 127 -1350 161
rect -1584 31 -1550 65
rect -1341 19 -1307 53
rect -1072 77 -1038 111
rect -888 77 -854 111
rect -627 77 -593 111
rect -414 77 -380 111
rect -181 77 -147 111
rect -89 77 -55 111
rect -5 77 29 111
rect 79 77 113 111
rect -2210 -387 -2176 -353
rect -2108 -402 -2074 -368
rect -1783 -329 -1749 -295
rect -1946 -455 -1912 -421
rect -1803 -425 -1769 -391
rect -1584 -341 -1550 -307
rect -1694 -503 -1660 -469
rect -1341 -329 -1307 -295
rect -1520 -437 -1486 -403
rect -1384 -437 -1350 -403
rect -1072 -387 -1038 -353
rect -888 -387 -854 -353
rect -627 -387 -593 -353
rect -414 -387 -380 -353
rect -181 -387 -147 -353
rect -89 -387 -55 -353
rect -5 -387 29 -353
rect 79 -387 113 -353
rect 488 -387 522 -353
rect -1282 -503 -1248 -469
rect -1146 -503 -1112 -469
rect 590 -402 624 -368
rect 915 -329 949 -295
rect 752 -455 786 -421
rect 895 -425 929 -391
rect 1114 -341 1148 -307
rect 1004 -503 1038 -469
rect 1357 -329 1391 -295
rect 1178 -437 1212 -403
rect 1314 -437 1348 -403
rect 1626 -387 1660 -353
rect 1810 -387 1844 -353
rect 2071 -387 2105 -353
rect 2284 -387 2318 -353
rect 2517 -387 2551 -353
rect 2609 -387 2643 -353
rect 2693 -387 2727 -353
rect 2777 -387 2811 -353
rect 1416 -503 1450 -469
rect 1552 -503 1586 -469
rect -2210 -1011 -2176 -977
rect -1946 -943 -1912 -909
rect -1694 -895 -1660 -861
rect -2108 -996 -2074 -962
rect -1803 -973 -1769 -939
rect -1783 -1069 -1749 -1035
rect -1282 -895 -1248 -861
rect -1146 -895 -1112 -861
rect -1520 -961 -1486 -927
rect -1384 -961 -1350 -927
rect -1584 -1057 -1550 -1023
rect -1341 -1069 -1307 -1035
rect -1072 -1011 -1038 -977
rect -888 -1011 -854 -977
rect -627 -1011 -593 -977
rect -414 -1011 -380 -977
rect -181 -1011 -147 -977
rect -89 -1011 -55 -977
rect -5 -1011 29 -977
rect 79 -1011 113 -977
rect 488 -1011 522 -977
rect 752 -943 786 -909
rect 1004 -895 1038 -861
rect 590 -996 624 -962
rect 895 -973 929 -939
rect 915 -1069 949 -1035
rect 1416 -895 1450 -861
rect 1552 -895 1586 -861
rect 1178 -961 1212 -927
rect 1314 -961 1348 -927
rect 1114 -1057 1148 -1023
rect 1357 -1069 1391 -1035
rect 1626 -1011 1660 -977
rect 1810 -1011 1844 -977
rect 2071 -1011 2105 -977
rect 2284 -1011 2318 -977
rect 2517 -1011 2551 -977
rect 2609 -1011 2643 -977
rect 2693 -1011 2727 -977
rect 2777 -1011 2811 -977
rect -2210 -1475 -2176 -1441
rect -2108 -1490 -2074 -1456
rect -1783 -1417 -1749 -1383
rect -1946 -1543 -1912 -1509
rect -1803 -1513 -1769 -1479
rect -1584 -1429 -1550 -1395
rect -1694 -1591 -1660 -1557
rect -1341 -1417 -1307 -1383
rect -1520 -1525 -1486 -1491
rect -1384 -1525 -1350 -1491
rect -1072 -1475 -1038 -1441
rect -888 -1475 -854 -1441
rect -627 -1475 -593 -1441
rect -414 -1475 -380 -1441
rect -181 -1475 -147 -1441
rect -89 -1475 -55 -1441
rect -5 -1475 29 -1441
rect 79 -1475 113 -1441
rect 488 -1475 522 -1441
rect -1282 -1591 -1248 -1557
rect -1146 -1591 -1112 -1557
rect 590 -1490 624 -1456
rect 915 -1417 949 -1383
rect 752 -1543 786 -1509
rect 895 -1513 929 -1479
rect 1114 -1429 1148 -1395
rect 1004 -1591 1038 -1557
rect 1357 -1417 1391 -1383
rect 1178 -1525 1212 -1491
rect 1314 -1525 1348 -1491
rect 1626 -1475 1660 -1441
rect 1810 -1475 1844 -1441
rect 2071 -1475 2105 -1441
rect 2284 -1475 2318 -1441
rect 2517 -1475 2551 -1441
rect 2609 -1475 2643 -1441
rect 2693 -1475 2727 -1441
rect 2777 -1475 2811 -1441
rect 1416 -1591 1450 -1557
rect 1552 -1591 1586 -1557
rect -2210 -2099 -2176 -2065
rect -1946 -2031 -1912 -1997
rect -1694 -1983 -1660 -1949
rect -2108 -2084 -2074 -2050
rect -1803 -2061 -1769 -2027
rect -1783 -2157 -1749 -2123
rect -1282 -1983 -1248 -1949
rect -1146 -1983 -1112 -1949
rect -1520 -2049 -1486 -2015
rect -1384 -2049 -1350 -2015
rect -1584 -2145 -1550 -2111
rect -1341 -2157 -1307 -2123
rect -1072 -2099 -1038 -2065
rect -888 -2099 -854 -2065
rect -627 -2099 -593 -2065
rect -414 -2099 -380 -2065
rect -181 -2099 -147 -2065
rect -89 -2099 -55 -2065
rect -5 -2099 29 -2065
rect 79 -2099 113 -2065
rect 488 -2099 522 -2065
rect 752 -2031 786 -1997
rect 1004 -1983 1038 -1949
rect 590 -2084 624 -2050
rect 895 -2061 929 -2027
rect 915 -2157 949 -2123
rect 1416 -1983 1450 -1949
rect 1552 -1983 1586 -1949
rect 1178 -2049 1212 -2015
rect 1314 -2049 1348 -2015
rect 1114 -2145 1148 -2111
rect 1357 -2157 1391 -2123
rect 1626 -2099 1660 -2065
rect 1810 -2099 1844 -2065
rect 2071 -2099 2105 -2065
rect 2284 -2099 2318 -2065
rect 2517 -2099 2551 -2065
rect 2609 -2099 2643 -2065
rect 2693 -2099 2727 -2065
rect 2777 -2099 2811 -2065
rect -2210 -2563 -2176 -2529
rect -2108 -2578 -2074 -2544
rect -1783 -2505 -1749 -2471
rect -1946 -2631 -1912 -2597
rect -1803 -2601 -1769 -2567
rect -1584 -2517 -1550 -2483
rect -1694 -2679 -1660 -2645
rect -1341 -2505 -1307 -2471
rect -1520 -2613 -1486 -2579
rect -1384 -2613 -1350 -2579
rect -1072 -2563 -1038 -2529
rect -888 -2563 -854 -2529
rect -627 -2563 -593 -2529
rect -414 -2563 -380 -2529
rect -181 -2563 -147 -2529
rect -89 -2563 -55 -2529
rect -5 -2563 29 -2529
rect 79 -2563 113 -2529
rect 488 -2563 522 -2529
rect -1282 -2679 -1248 -2645
rect -1146 -2679 -1112 -2645
rect 590 -2578 624 -2544
rect 915 -2505 949 -2471
rect 752 -2631 786 -2597
rect 895 -2601 929 -2567
rect 1114 -2517 1148 -2483
rect 1004 -2679 1038 -2645
rect 1357 -2505 1391 -2471
rect 1178 -2613 1212 -2579
rect 1314 -2613 1348 -2579
rect 1626 -2563 1660 -2529
rect 1810 -2563 1844 -2529
rect 2071 -2563 2105 -2529
rect 2284 -2563 2318 -2529
rect 2517 -2563 2551 -2529
rect 2609 -2563 2643 -2529
rect 2693 -2563 2727 -2529
rect 2777 -2563 2811 -2529
rect 1416 -2679 1450 -2645
rect 1552 -2679 1586 -2645
<< locali >>
rect -2584 389 -2555 423
rect -2521 389 -2492 423
rect -2242 389 -2213 423
rect -2179 389 -2121 423
rect -2087 389 -2029 423
rect -1995 389 -1937 423
rect -1903 389 -1845 423
rect -1811 389 -1753 423
rect -1719 389 -1661 423
rect -1627 389 -1569 423
rect -1535 389 -1477 423
rect -1443 389 -1385 423
rect -1351 389 -1293 423
rect -1259 389 -1201 423
rect -1167 389 -1109 423
rect -1075 389 -1017 423
rect -983 389 -925 423
rect -891 389 -833 423
rect -799 389 -741 423
rect -707 389 -649 423
rect -615 389 -557 423
rect -523 389 -465 423
rect -431 389 -373 423
rect -339 389 -281 423
rect -247 389 -189 423
rect -155 389 -97 423
rect -63 389 -5 423
rect 29 389 87 423
rect 121 389 179 423
rect 213 389 242 423
rect 316 389 345 423
rect 379 389 408 423
rect 3190 389 3219 423
rect 3253 389 3282 423
rect -2567 318 -2509 389
rect -2567 284 -2555 318
rect -2521 284 -2509 318
rect -2567 225 -2509 284
rect -2567 191 -2555 225
rect -2521 191 -2509 225
rect -2207 339 -2173 355
rect -2207 271 -2173 305
rect -2139 323 -2073 389
rect -2139 289 -2123 323
rect -2089 289 -2073 323
rect -2039 339 -2002 355
rect -2005 305 -2002 339
rect -2039 271 -2002 305
rect -1954 347 -1901 389
rect -1954 313 -1935 347
rect -1954 297 -1901 313
rect -1867 339 -1817 355
rect -1867 305 -1851 339
rect -1520 347 -1486 389
rect -2173 253 -2074 255
rect -2173 237 -2116 253
rect -2207 221 -2116 237
rect -2567 156 -2509 191
rect -2120 219 -2116 221
rect -2082 219 -2074 253
rect -2224 146 -2154 187
rect -2224 98 -2214 146
rect -2166 98 -2154 146
rect -2224 77 -2210 98
rect -2176 77 -2154 98
rect -2224 57 -2154 77
rect -2120 126 -2074 219
rect -2120 92 -2108 126
rect -2567 7 -2509 24
rect -2120 23 -2074 92
rect -2567 -27 -2555 7
rect -2521 -27 -2509 7
rect -2567 -121 -2509 -27
rect -2207 -11 -2074 23
rect -2005 237 -2002 271
rect -1867 270 -1817 305
rect -1775 300 -1759 334
rect -1725 300 -1554 334
rect -2039 185 -2002 237
rect -1878 244 -1817 270
rect -1728 253 -1622 266
rect -2039 151 -2037 185
rect -2003 151 -2002 185
rect -2207 -19 -2173 -11
rect -2039 -19 -2002 151
rect -1968 179 -1912 195
rect -1968 145 -1946 179
rect -1968 88 -1912 145
rect -1968 40 -1962 88
rect -1914 40 -1912 88
rect -1968 5 -1912 40
rect -1878 23 -1844 244
rect -1728 219 -1696 253
rect -1662 227 -1622 253
rect -1810 185 -1762 206
rect -1810 151 -1799 185
rect -1765 151 -1762 185
rect -1810 149 -1762 151
rect -1810 115 -1803 149
rect -1769 115 -1762 149
rect -1810 87 -1762 115
rect -1728 53 -1694 219
rect -1660 193 -1622 227
rect -1588 177 -1554 300
rect -1520 279 -1486 313
rect -1520 229 -1486 245
rect -1452 339 -1402 355
rect -1452 305 -1436 339
rect -1144 339 -1081 389
rect -1452 289 -1402 305
rect -1357 295 -1341 329
rect -1307 295 -1180 329
rect -1588 161 -1486 177
rect -1588 159 -1520 161
rect -1878 -3 -1833 23
rect -1799 19 -1783 53
rect -1749 19 -1694 53
rect -1799 9 -1694 19
rect -1660 127 -1520 159
rect -1660 125 -1486 127
rect -2207 -69 -2173 -53
rect -2139 -79 -2123 -45
rect -2089 -79 -2073 -45
rect -2005 -53 -2002 -19
rect -2039 -69 -2002 -53
rect -1951 -45 -1901 -29
rect -2139 -121 -2073 -79
rect -1951 -79 -1935 -45
rect -1867 -31 -1833 -3
rect -1660 -31 -1626 125
rect -1520 111 -1486 125
rect -1584 75 -1544 81
rect -1452 75 -1418 289
rect -1384 253 -1346 255
rect -1384 219 -1382 253
rect -1348 219 -1346 253
rect -1384 161 -1346 219
rect -1350 127 -1346 161
rect -1384 111 -1346 127
rect -1312 227 -1248 261
rect -1312 193 -1282 227
rect -1312 185 -1248 193
rect -1312 151 -1295 185
rect -1261 151 -1248 185
rect -1584 65 -1418 75
rect -1312 69 -1248 151
rect -1550 31 -1418 65
rect -1584 15 -1418 31
rect -1867 -65 -1850 -31
rect -1816 -65 -1800 -31
rect -1761 -65 -1739 -31
rect -1705 -65 -1626 -31
rect -1562 -37 -1488 -21
rect -1951 -121 -1901 -79
rect -1562 -71 -1540 -37
rect -1506 -71 -1488 -37
rect -1452 -31 -1418 15
rect -1341 53 -1248 69
rect -1307 19 -1248 53
rect -1341 3 -1248 19
rect -1214 127 -1180 295
rect -1144 305 -1142 339
rect -1108 305 -1081 339
rect -1144 289 -1081 305
rect -1034 347 -966 355
rect -1034 313 -1018 347
rect -984 313 -966 347
rect -1034 276 -966 313
rect -1034 243 -1018 276
rect -1146 242 -1018 243
rect -984 242 -966 276
rect -1146 227 -966 242
rect -1112 205 -966 227
rect -1112 193 -1018 205
rect -1146 171 -1018 193
rect -984 171 -966 205
rect -932 317 -898 389
rect -760 347 -694 351
rect -932 237 -898 283
rect -932 187 -898 203
rect -864 341 -798 346
rect -864 307 -848 341
rect -814 307 -798 341
rect -864 273 -798 307
rect -864 239 -848 273
rect -814 239 -798 273
rect -864 205 -798 239
rect -760 313 -744 347
rect -710 313 -694 347
rect -760 279 -694 313
rect -760 245 -744 279
rect -710 245 -694 279
rect -760 205 -694 245
rect -1146 168 -966 171
rect -1004 127 -966 168
rect -864 171 -848 205
rect -814 177 -798 205
rect -814 171 -782 177
rect -864 161 -782 171
rect -829 151 -782 161
rect -1214 111 -1038 127
rect -1214 77 -1072 111
rect -1214 61 -1038 77
rect -1004 111 -854 127
rect -1004 77 -888 111
rect -1004 61 -854 77
rect -1214 -31 -1180 61
rect -1004 27 -964 61
rect -820 35 -782 151
rect -831 27 -782 35
rect -1030 24 -964 27
rect -1030 -10 -1014 24
rect -980 -10 -964 24
rect -862 26 -782 27
rect -862 8 -846 26
rect -812 10 -782 26
rect -748 127 -694 205
rect -656 347 -613 389
rect -656 313 -647 347
rect -656 279 -613 313
rect -656 245 -647 279
rect -656 211 -613 245
rect -656 177 -647 211
rect -656 161 -613 177
rect -579 347 -512 355
rect -579 313 -563 347
rect -529 313 -512 347
rect -579 276 -512 313
rect -579 242 -563 276
rect -529 242 -512 276
rect -579 205 -512 242
rect -579 171 -563 205
rect -529 171 -512 205
rect -579 158 -512 171
rect -426 347 -384 389
rect -426 313 -418 347
rect -426 279 -384 313
rect -426 245 -418 279
rect -426 211 -384 245
rect -426 177 -418 211
rect -426 161 -384 177
rect -350 347 -284 355
rect -350 313 -334 347
rect -300 313 -284 347
rect -350 279 -284 313
rect -350 245 -334 279
rect -300 245 -284 279
rect -350 211 -284 245
rect -350 177 -334 211
rect -300 177 -284 211
rect -350 159 -284 177
rect -192 347 -139 389
rect -192 313 -173 347
rect -192 279 -139 313
rect -192 245 -173 279
rect -192 211 -139 245
rect -192 177 -173 211
rect -192 161 -139 177
rect -105 347 -39 355
rect -105 313 -89 347
rect -55 313 -39 347
rect -105 279 -39 313
rect -105 245 -89 279
rect -55 245 -39 279
rect -105 211 -39 245
rect -5 347 29 389
rect -5 279 29 313
rect -5 229 29 245
rect 63 347 129 355
rect 63 313 79 347
rect 113 313 129 347
rect 63 279 129 313
rect 163 347 205 389
rect 197 313 205 347
rect 163 297 205 313
rect 333 318 391 389
rect 63 245 79 279
rect 113 245 129 279
rect -105 177 -89 211
rect -55 195 -39 211
rect 63 211 129 245
rect 63 195 79 211
rect -55 177 79 195
rect 113 199 129 211
rect 333 284 345 318
rect 379 284 391 318
rect 333 225 391 284
rect 113 177 216 199
rect -105 161 216 177
rect -748 111 -593 127
rect -748 77 -627 111
rect -748 61 -593 77
rect -559 126 -512 158
rect -330 126 -284 159
rect -197 126 129 127
rect -559 78 -552 126
rect -388 111 -364 125
rect -812 8 -796 10
rect -1452 -65 -1421 -31
rect -1387 -65 -1371 -31
rect -1337 -65 -1318 -31
rect -1284 -65 -1180 -31
rect -1125 -31 -1083 -15
rect -1125 -65 -1120 -31
rect -1086 -65 -1083 -31
rect -1562 -121 -1488 -71
rect -1125 -121 -1083 -65
rect -1030 -44 -964 -10
rect -1030 -78 -1014 -44
rect -980 -78 -964 -44
rect -930 -15 -896 1
rect -930 -121 -896 -49
rect -862 -40 -858 8
rect -810 -40 -796 8
rect -748 -15 -708 61
rect -559 44 -512 78
rect -430 77 -414 78
rect -380 77 -364 111
rect -330 78 -324 126
rect -197 78 -192 126
rect -144 111 -82 126
rect -34 111 34 126
rect 82 111 129 126
rect -144 78 -89 111
rect -34 78 -5 111
rect -862 -42 -796 -40
rect -862 -76 -846 -42
rect -812 -76 -796 -42
rect -758 -19 -708 -15
rect -758 -53 -742 -19
rect -563 -7 -512 44
rect -758 -69 -708 -53
rect -661 -45 -597 -29
rect -862 -77 -796 -76
rect -661 -79 -647 -45
rect -613 -79 -597 -45
rect -661 -121 -597 -79
rect -529 -41 -512 -7
rect -563 -87 -512 -41
rect -430 27 -384 43
rect -330 39 -284 78
rect -197 77 -181 78
rect -147 77 -89 78
rect -55 77 -5 78
rect 29 78 34 111
rect 29 77 79 78
rect 113 77 129 111
rect 163 124 216 161
rect 333 191 345 225
rect 379 191 391 225
rect 333 156 391 191
rect 3207 318 3265 389
rect 3207 284 3219 318
rect 3253 284 3265 318
rect 3207 225 3265 284
rect 3207 191 3219 225
rect 3253 191 3265 225
rect 3207 156 3265 191
rect 163 76 166 124
rect 214 76 216 124
rect 163 43 216 76
rect -430 -7 -418 27
rect -430 -41 -384 -7
rect -430 -75 -418 -41
rect -430 -121 -384 -75
rect -350 27 -284 39
rect -350 -7 -334 27
rect -300 -7 -284 27
rect -350 -41 -284 -7
rect -105 7 216 43
rect 333 7 391 24
rect -350 -75 -334 -41
rect -300 -75 -284 -41
rect -350 -87 -284 -75
rect -192 -45 -139 -29
rect -192 -79 -173 -45
rect -192 -121 -139 -79
rect -105 -37 -39 7
rect -105 -71 -89 -37
rect -55 -71 -39 -37
rect -105 -87 -39 -71
rect -5 -45 29 -29
rect -5 -121 29 -79
rect 63 -37 129 7
rect 333 -27 345 7
rect 379 -27 391 7
rect 63 -71 79 -37
rect 113 -71 129 -37
rect 63 -87 129 -71
rect 163 -44 213 -28
rect 197 -78 213 -44
rect 163 -121 213 -78
rect 333 -121 391 -27
rect 3207 7 3265 24
rect 3207 -27 3219 7
rect 3253 -27 3265 7
rect 3207 -121 3265 -27
rect -2584 -155 -2555 -121
rect -2521 -155 -2492 -121
rect -2242 -155 -2213 -121
rect -2179 -155 -2121 -121
rect -2087 -155 -2029 -121
rect -1995 -155 -1937 -121
rect -1903 -155 -1845 -121
rect -1811 -155 -1753 -121
rect -1719 -155 -1661 -121
rect -1627 -155 -1569 -121
rect -1535 -155 -1477 -121
rect -1443 -155 -1385 -121
rect -1351 -155 -1293 -121
rect -1259 -155 -1201 -121
rect -1167 -155 -1109 -121
rect -1075 -155 -1017 -121
rect -983 -155 -925 -121
rect -891 -155 -833 -121
rect -799 -155 -741 -121
rect -707 -155 -649 -121
rect -615 -155 -557 -121
rect -523 -155 -465 -121
rect -431 -155 -373 -121
rect -339 -155 -281 -121
rect -247 -155 -189 -121
rect -155 -155 -97 -121
rect -63 -155 -5 -121
rect 29 -155 87 -121
rect 121 -155 179 -121
rect 213 -155 242 -121
rect 316 -155 345 -121
rect 379 -155 408 -121
rect 456 -155 485 -121
rect 519 -155 577 -121
rect 611 -155 669 -121
rect 703 -155 761 -121
rect 795 -155 853 -121
rect 887 -155 945 -121
rect 979 -155 1037 -121
rect 1071 -155 1129 -121
rect 1163 -155 1221 -121
rect 1255 -155 1313 -121
rect 1347 -155 1405 -121
rect 1439 -155 1497 -121
rect 1531 -155 1589 -121
rect 1623 -155 1681 -121
rect 1715 -155 1773 -121
rect 1807 -155 1865 -121
rect 1899 -155 1957 -121
rect 1991 -155 2049 -121
rect 2083 -155 2141 -121
rect 2175 -155 2233 -121
rect 2267 -155 2325 -121
rect 2359 -155 2417 -121
rect 2451 -155 2509 -121
rect 2543 -155 2601 -121
rect 2635 -155 2693 -121
rect 2727 -155 2785 -121
rect 2819 -155 2877 -121
rect 2911 -155 2940 -121
rect 3190 -155 3219 -121
rect 3253 -155 3282 -121
rect -2567 -249 -2509 -155
rect -2139 -197 -2073 -155
rect -2567 -283 -2555 -249
rect -2521 -283 -2509 -249
rect -2567 -300 -2509 -283
rect -2207 -223 -2173 -207
rect -2139 -231 -2123 -197
rect -2089 -231 -2073 -197
rect -1951 -197 -1901 -155
rect -2039 -223 -2002 -207
rect -2207 -265 -2173 -257
rect -2005 -257 -2002 -223
rect -1951 -231 -1935 -197
rect -1562 -205 -1488 -155
rect -1951 -247 -1901 -231
rect -1867 -245 -1850 -211
rect -1816 -245 -1800 -211
rect -1761 -245 -1739 -211
rect -1705 -245 -1626 -211
rect -2207 -299 -2074 -265
rect -2224 -353 -2154 -333
rect -2224 -364 -2210 -353
rect -2176 -364 -2154 -353
rect -2224 -412 -2218 -364
rect -2170 -412 -2154 -364
rect -2567 -467 -2509 -432
rect -2224 -463 -2154 -412
rect -2120 -368 -2074 -299
rect -2120 -402 -2108 -368
rect -2567 -501 -2555 -467
rect -2521 -501 -2509 -467
rect -2120 -495 -2074 -402
rect -2120 -497 -2116 -495
rect -2567 -560 -2509 -501
rect -2567 -594 -2555 -560
rect -2521 -594 -2509 -560
rect -2567 -665 -2509 -594
rect -2207 -513 -2116 -497
rect -2173 -529 -2116 -513
rect -2082 -529 -2074 -495
rect -2173 -531 -2074 -529
rect -2039 -427 -2002 -257
rect -1867 -273 -1833 -245
rect -2039 -461 -2037 -427
rect -2003 -461 -2002 -427
rect -2039 -513 -2002 -461
rect -1968 -316 -1912 -281
rect -1968 -364 -1962 -316
rect -1914 -364 -1912 -316
rect -1968 -421 -1912 -364
rect -1968 -455 -1946 -421
rect -1968 -471 -1912 -455
rect -1878 -299 -1833 -273
rect -1799 -295 -1694 -285
rect -2207 -581 -2173 -547
rect -2005 -547 -2002 -513
rect -1878 -520 -1844 -299
rect -1799 -329 -1783 -295
rect -1749 -329 -1694 -295
rect -1810 -391 -1762 -363
rect -1810 -425 -1803 -391
rect -1769 -425 -1762 -391
rect -1810 -427 -1762 -425
rect -1810 -461 -1799 -427
rect -1765 -461 -1762 -427
rect -1810 -482 -1762 -461
rect -1728 -495 -1694 -329
rect -1660 -401 -1626 -245
rect -1562 -239 -1540 -205
rect -1506 -239 -1488 -205
rect -1125 -211 -1083 -155
rect -1562 -255 -1488 -239
rect -1452 -245 -1421 -211
rect -1387 -245 -1371 -211
rect -1337 -245 -1318 -211
rect -1284 -245 -1180 -211
rect -1452 -291 -1418 -245
rect -1584 -307 -1418 -291
rect -1550 -341 -1418 -307
rect -1584 -351 -1418 -341
rect -1341 -295 -1248 -279
rect -1307 -329 -1248 -295
rect -1341 -345 -1248 -329
rect -1584 -357 -1544 -351
rect -1520 -401 -1486 -387
rect -1660 -403 -1486 -401
rect -1660 -435 -1520 -403
rect -1588 -437 -1520 -435
rect -1588 -453 -1486 -437
rect -1878 -546 -1817 -520
rect -1728 -529 -1696 -495
rect -1660 -503 -1622 -469
rect -1662 -529 -1622 -503
rect -1728 -542 -1622 -529
rect -2207 -631 -2173 -615
rect -2139 -599 -2123 -565
rect -2089 -599 -2073 -565
rect -2139 -665 -2073 -599
rect -2039 -581 -2002 -547
rect -2005 -615 -2002 -581
rect -2039 -631 -2002 -615
rect -1954 -589 -1901 -573
rect -1954 -623 -1935 -589
rect -1954 -665 -1901 -623
rect -1867 -581 -1817 -546
rect -1588 -576 -1554 -453
rect -1867 -615 -1851 -581
rect -1775 -610 -1759 -576
rect -1725 -610 -1554 -576
rect -1520 -521 -1486 -505
rect -1520 -589 -1486 -555
rect -1867 -631 -1817 -615
rect -1520 -665 -1486 -623
rect -1452 -565 -1418 -351
rect -1384 -403 -1346 -387
rect -1350 -437 -1346 -403
rect -1384 -495 -1346 -437
rect -1384 -529 -1382 -495
rect -1348 -529 -1346 -495
rect -1384 -531 -1346 -529
rect -1312 -427 -1248 -345
rect -1312 -461 -1295 -427
rect -1261 -461 -1248 -427
rect -1312 -469 -1248 -461
rect -1312 -503 -1282 -469
rect -1312 -537 -1248 -503
rect -1214 -337 -1180 -245
rect -1125 -245 -1120 -211
rect -1086 -245 -1083 -211
rect -1125 -261 -1083 -245
rect -1030 -232 -1014 -198
rect -980 -232 -964 -198
rect -1030 -266 -964 -232
rect -1030 -300 -1014 -266
rect -980 -300 -964 -266
rect -930 -227 -896 -155
rect -661 -197 -597 -155
rect -930 -277 -896 -261
rect -862 -200 -796 -199
rect -862 -234 -846 -200
rect -812 -234 -796 -200
rect -862 -268 -796 -234
rect -758 -223 -708 -207
rect -758 -257 -742 -223
rect -661 -231 -647 -197
rect -613 -231 -597 -197
rect -661 -247 -597 -231
rect -563 -235 -512 -189
rect -758 -261 -708 -257
rect -1030 -303 -964 -300
rect -862 -302 -846 -268
rect -812 -286 -796 -268
rect -812 -302 -782 -286
rect -862 -303 -782 -302
rect -1004 -337 -964 -303
rect -831 -311 -782 -303
rect -1214 -353 -1038 -337
rect -1214 -387 -1072 -353
rect -1214 -403 -1038 -387
rect -1004 -353 -854 -337
rect -1004 -387 -888 -353
rect -1004 -403 -854 -387
rect -1452 -581 -1402 -565
rect -1214 -571 -1180 -403
rect -1004 -444 -966 -403
rect -820 -427 -782 -311
rect -829 -437 -782 -427
rect -1146 -447 -966 -444
rect -1146 -469 -1018 -447
rect -1112 -481 -1018 -469
rect -984 -481 -966 -447
rect -864 -447 -782 -437
rect -1112 -503 -966 -481
rect -1146 -518 -966 -503
rect -1146 -519 -1018 -518
rect -1034 -552 -1018 -519
rect -984 -552 -966 -518
rect -1452 -615 -1436 -581
rect -1357 -605 -1341 -571
rect -1307 -605 -1180 -571
rect -1144 -581 -1081 -565
rect -1452 -631 -1402 -615
rect -1144 -615 -1142 -581
rect -1108 -615 -1081 -581
rect -1144 -665 -1081 -615
rect -1034 -589 -966 -552
rect -1034 -623 -1018 -589
rect -984 -623 -966 -589
rect -1034 -631 -966 -623
rect -932 -479 -898 -463
rect -932 -559 -898 -513
rect -932 -665 -898 -593
rect -864 -481 -848 -447
rect -814 -453 -782 -447
rect -748 -337 -708 -261
rect -529 -269 -512 -235
rect -563 -320 -512 -269
rect -430 -201 -384 -155
rect -430 -235 -418 -201
rect -430 -269 -384 -235
rect -430 -303 -418 -269
rect -430 -319 -384 -303
rect -350 -201 -284 -189
rect -350 -235 -334 -201
rect -300 -235 -284 -201
rect -350 -269 -284 -235
rect -192 -197 -139 -155
rect -192 -231 -173 -197
rect -192 -247 -139 -231
rect -105 -205 -39 -189
rect -105 -239 -89 -205
rect -55 -239 -39 -205
rect -350 -303 -334 -269
rect -300 -303 -284 -269
rect -350 -315 -284 -303
rect -748 -353 -593 -337
rect -748 -387 -627 -353
rect -748 -403 -593 -387
rect -559 -354 -512 -320
rect -430 -354 -414 -353
rect -559 -402 -552 -354
rect -380 -387 -364 -353
rect -388 -401 -364 -387
rect -330 -354 -284 -315
rect -105 -283 -39 -239
rect -5 -197 29 -155
rect -5 -247 29 -231
rect 63 -205 129 -189
rect 63 -239 79 -205
rect 113 -239 129 -205
rect 63 -283 129 -239
rect 163 -198 213 -155
rect 197 -232 213 -198
rect 559 -197 625 -155
rect 163 -248 213 -232
rect 491 -223 525 -207
rect 559 -231 575 -197
rect 609 -231 625 -197
rect 747 -197 797 -155
rect 659 -223 696 -207
rect 491 -265 525 -257
rect 693 -257 696 -223
rect 747 -231 763 -197
rect 1136 -205 1210 -155
rect 747 -247 797 -231
rect 831 -245 848 -211
rect 882 -245 898 -211
rect 937 -245 959 -211
rect 993 -245 1072 -211
rect -105 -319 216 -283
rect 491 -299 624 -265
rect 163 -352 216 -319
rect -197 -354 -181 -353
rect -147 -354 -89 -353
rect -55 -354 -5 -353
rect -330 -402 -324 -354
rect -197 -402 -192 -354
rect -144 -387 -89 -354
rect -34 -387 -5 -354
rect 29 -354 79 -353
rect 29 -387 34 -354
rect 113 -387 129 -353
rect -144 -402 -82 -387
rect -34 -402 34 -387
rect 82 -402 129 -387
rect -814 -481 -798 -453
rect -748 -481 -694 -403
rect -559 -434 -512 -402
rect -864 -515 -798 -481
rect -864 -538 -848 -515
rect -814 -538 -798 -515
rect -864 -586 -858 -538
rect -810 -586 -798 -538
rect -864 -617 -848 -586
rect -814 -617 -798 -586
rect -864 -622 -798 -617
rect -760 -521 -694 -481
rect -760 -555 -744 -521
rect -710 -555 -694 -521
rect -760 -589 -694 -555
rect -760 -623 -744 -589
rect -710 -623 -694 -589
rect -760 -627 -694 -623
rect -656 -453 -613 -437
rect -656 -487 -647 -453
rect -656 -521 -613 -487
rect -656 -555 -647 -521
rect -656 -589 -613 -555
rect -656 -623 -647 -589
rect -656 -665 -613 -623
rect -579 -447 -512 -434
rect -330 -435 -284 -402
rect -197 -403 129 -402
rect 163 -400 170 -352
rect 474 -353 544 -333
rect 474 -387 488 -353
rect 522 -387 544 -353
rect -579 -481 -563 -447
rect -529 -481 -512 -447
rect -579 -518 -512 -481
rect -579 -552 -563 -518
rect -529 -552 -512 -518
rect -579 -589 -512 -552
rect -579 -623 -563 -589
rect -529 -623 -512 -589
rect -579 -631 -512 -623
rect -426 -453 -384 -437
rect -426 -487 -418 -453
rect -426 -521 -384 -487
rect -426 -555 -418 -521
rect -426 -589 -384 -555
rect -426 -623 -418 -589
rect -426 -665 -384 -623
rect -350 -453 -284 -435
rect 163 -437 216 -400
rect -350 -487 -334 -453
rect -300 -487 -284 -453
rect -350 -521 -284 -487
rect -350 -555 -334 -521
rect -300 -555 -284 -521
rect -350 -589 -284 -555
rect -350 -623 -334 -589
rect -300 -623 -284 -589
rect -350 -631 -284 -623
rect -192 -453 -139 -437
rect -192 -487 -173 -453
rect -192 -521 -139 -487
rect -192 -555 -173 -521
rect -192 -589 -139 -555
rect -192 -623 -173 -589
rect -192 -665 -139 -623
rect -105 -453 216 -437
rect -105 -487 -89 -453
rect -55 -471 79 -453
rect -55 -487 -39 -471
rect -105 -521 -39 -487
rect 63 -487 79 -471
rect 113 -475 216 -453
rect 474 -406 544 -387
rect 474 -454 480 -406
rect 528 -454 544 -406
rect 474 -463 544 -454
rect 578 -368 624 -299
rect 578 -402 590 -368
rect 113 -487 129 -475
rect -105 -555 -89 -521
rect -55 -555 -39 -521
rect -105 -589 -39 -555
rect -105 -623 -89 -589
rect -55 -623 -39 -589
rect -105 -631 -39 -623
rect -5 -521 29 -505
rect -5 -589 29 -555
rect -5 -665 29 -623
rect 63 -521 129 -487
rect 578 -495 624 -402
rect 578 -497 582 -495
rect 63 -555 79 -521
rect 113 -555 129 -521
rect 63 -589 129 -555
rect 491 -513 582 -497
rect 525 -529 582 -513
rect 616 -529 624 -495
rect 525 -531 624 -529
rect 659 -427 696 -257
rect 831 -273 865 -245
rect 659 -461 661 -427
rect 695 -461 696 -427
rect 659 -513 696 -461
rect 730 -316 786 -281
rect 730 -364 736 -316
rect 784 -364 786 -316
rect 730 -421 786 -364
rect 730 -455 752 -421
rect 730 -471 786 -455
rect 820 -299 865 -273
rect 899 -295 1004 -285
rect 63 -623 79 -589
rect 113 -623 129 -589
rect 63 -631 129 -623
rect 163 -589 205 -573
rect 197 -623 205 -589
rect 163 -665 205 -623
rect 491 -581 525 -547
rect 693 -547 696 -513
rect 820 -520 854 -299
rect 899 -329 915 -295
rect 949 -329 1004 -295
rect 888 -391 936 -363
rect 888 -425 895 -391
rect 929 -425 936 -391
rect 888 -427 936 -425
rect 888 -461 899 -427
rect 933 -461 936 -427
rect 888 -482 936 -461
rect 970 -495 1004 -329
rect 1038 -401 1072 -245
rect 1136 -239 1158 -205
rect 1192 -239 1210 -205
rect 1573 -211 1615 -155
rect 1136 -255 1210 -239
rect 1246 -245 1277 -211
rect 1311 -245 1327 -211
rect 1361 -245 1380 -211
rect 1414 -245 1518 -211
rect 1246 -291 1280 -245
rect 1114 -307 1280 -291
rect 1148 -341 1280 -307
rect 1114 -351 1280 -341
rect 1357 -295 1450 -279
rect 1391 -329 1450 -295
rect 1357 -345 1450 -329
rect 1114 -357 1154 -351
rect 1178 -401 1212 -387
rect 1038 -403 1212 -401
rect 1038 -435 1178 -403
rect 1110 -437 1178 -435
rect 1110 -453 1212 -437
rect 820 -546 881 -520
rect 970 -529 1002 -495
rect 1038 -503 1076 -469
rect 1036 -529 1076 -503
rect 970 -542 1076 -529
rect 491 -631 525 -615
rect 559 -599 575 -565
rect 609 -599 625 -565
rect 559 -665 625 -599
rect 659 -581 696 -547
rect 693 -615 696 -581
rect 659 -631 696 -615
rect 744 -589 797 -573
rect 744 -623 763 -589
rect 744 -665 797 -623
rect 831 -581 881 -546
rect 1110 -576 1144 -453
rect 831 -615 847 -581
rect 923 -610 939 -576
rect 973 -610 1144 -576
rect 1178 -521 1212 -505
rect 1178 -589 1212 -555
rect 831 -631 881 -615
rect 1178 -665 1212 -623
rect 1246 -565 1280 -351
rect 1314 -403 1352 -387
rect 1348 -437 1352 -403
rect 1314 -495 1352 -437
rect 1314 -529 1316 -495
rect 1350 -529 1352 -495
rect 1314 -531 1352 -529
rect 1386 -427 1450 -345
rect 1386 -461 1403 -427
rect 1437 -461 1450 -427
rect 1386 -469 1450 -461
rect 1386 -503 1416 -469
rect 1386 -537 1450 -503
rect 1484 -337 1518 -245
rect 1573 -245 1578 -211
rect 1612 -245 1615 -211
rect 1573 -261 1615 -245
rect 1668 -232 1684 -198
rect 1718 -232 1734 -198
rect 1668 -266 1734 -232
rect 1668 -300 1684 -266
rect 1718 -300 1734 -266
rect 1768 -227 1802 -155
rect 2037 -197 2101 -155
rect 1768 -277 1802 -261
rect 1836 -200 1902 -199
rect 1836 -234 1852 -200
rect 1886 -234 1902 -200
rect 1836 -240 1902 -234
rect 1668 -303 1734 -300
rect 1836 -288 1842 -240
rect 1890 -286 1902 -240
rect 1940 -223 1990 -207
rect 1940 -257 1956 -223
rect 2037 -231 2051 -197
rect 2085 -231 2101 -197
rect 2037 -247 2101 -231
rect 2135 -235 2186 -189
rect 1940 -261 1990 -257
rect 1890 -288 1916 -286
rect 1836 -302 1852 -288
rect 1886 -302 1916 -288
rect 1836 -303 1916 -302
rect 1694 -337 1734 -303
rect 1867 -311 1916 -303
rect 1484 -353 1660 -337
rect 1484 -387 1626 -353
rect 1484 -403 1660 -387
rect 1694 -353 1844 -337
rect 1694 -387 1810 -353
rect 1694 -403 1844 -387
rect 1246 -581 1296 -565
rect 1484 -571 1518 -403
rect 1694 -444 1732 -403
rect 1878 -427 1916 -311
rect 1869 -437 1916 -427
rect 1552 -447 1732 -444
rect 1552 -469 1680 -447
rect 1586 -481 1680 -469
rect 1714 -481 1732 -447
rect 1834 -447 1916 -437
rect 1586 -503 1732 -481
rect 1552 -518 1732 -503
rect 1552 -519 1680 -518
rect 1664 -552 1680 -519
rect 1714 -552 1732 -518
rect 1246 -615 1262 -581
rect 1341 -605 1357 -571
rect 1391 -605 1518 -571
rect 1554 -581 1617 -565
rect 1246 -631 1296 -615
rect 1554 -615 1556 -581
rect 1590 -615 1617 -581
rect 1554 -665 1617 -615
rect 1664 -589 1732 -552
rect 1664 -623 1680 -589
rect 1714 -623 1732 -589
rect 1664 -631 1732 -623
rect 1766 -479 1800 -463
rect 1766 -559 1800 -513
rect 1766 -665 1800 -593
rect 1834 -481 1850 -447
rect 1884 -453 1916 -447
rect 1950 -337 1990 -261
rect 2169 -269 2186 -235
rect 2135 -320 2186 -269
rect 2268 -201 2314 -155
rect 2268 -235 2280 -201
rect 2268 -269 2314 -235
rect 2268 -303 2280 -269
rect 2268 -319 2314 -303
rect 2348 -201 2414 -189
rect 2348 -235 2364 -201
rect 2398 -235 2414 -201
rect 2348 -269 2414 -235
rect 2506 -197 2559 -155
rect 2506 -231 2525 -197
rect 2506 -247 2559 -231
rect 2593 -205 2659 -189
rect 2593 -239 2609 -205
rect 2643 -239 2659 -205
rect 2348 -303 2364 -269
rect 2398 -303 2414 -269
rect 2348 -315 2414 -303
rect 1950 -353 2105 -337
rect 1950 -387 2071 -353
rect 1950 -403 2105 -387
rect 2139 -354 2186 -320
rect 2268 -354 2284 -353
rect 2139 -402 2146 -354
rect 2318 -387 2334 -353
rect 2310 -401 2334 -387
rect 2368 -354 2414 -315
rect 2593 -283 2659 -239
rect 2693 -197 2727 -155
rect 2693 -247 2727 -231
rect 2761 -205 2827 -189
rect 2761 -239 2777 -205
rect 2811 -239 2827 -205
rect 2761 -283 2827 -239
rect 2861 -198 2911 -155
rect 2895 -232 2911 -198
rect 2861 -248 2911 -232
rect 3207 -249 3265 -155
rect 3207 -283 3219 -249
rect 3253 -283 3265 -249
rect 2593 -319 2914 -283
rect 3207 -300 3265 -283
rect 2861 -352 2914 -319
rect 2501 -354 2517 -353
rect 2551 -354 2609 -353
rect 2643 -354 2693 -353
rect 2368 -402 2374 -354
rect 2501 -402 2506 -354
rect 2554 -387 2609 -354
rect 2664 -387 2693 -354
rect 2727 -354 2777 -353
rect 2727 -387 2732 -354
rect 2811 -387 2827 -353
rect 2554 -402 2616 -387
rect 2664 -402 2732 -387
rect 2780 -402 2827 -387
rect 1884 -481 1900 -453
rect 1950 -481 2004 -403
rect 2139 -434 2186 -402
rect 1834 -515 1900 -481
rect 1834 -549 1850 -515
rect 1884 -549 1900 -515
rect 1834 -583 1900 -549
rect 1834 -617 1850 -583
rect 1884 -617 1900 -583
rect 1834 -622 1900 -617
rect 1938 -521 2004 -481
rect 1938 -555 1954 -521
rect 1988 -555 2004 -521
rect 1938 -589 2004 -555
rect 1938 -623 1954 -589
rect 1988 -623 2004 -589
rect 1938 -627 2004 -623
rect 2042 -453 2085 -437
rect 2042 -487 2051 -453
rect 2042 -521 2085 -487
rect 2042 -555 2051 -521
rect 2042 -589 2085 -555
rect 2042 -623 2051 -589
rect 2042 -665 2085 -623
rect 2119 -447 2186 -434
rect 2368 -435 2414 -402
rect 2501 -403 2827 -402
rect 2861 -400 2864 -352
rect 2912 -400 2914 -352
rect 2119 -481 2135 -447
rect 2169 -481 2186 -447
rect 2119 -518 2186 -481
rect 2119 -552 2135 -518
rect 2169 -552 2186 -518
rect 2119 -589 2186 -552
rect 2119 -623 2135 -589
rect 2169 -623 2186 -589
rect 2119 -631 2186 -623
rect 2272 -453 2314 -437
rect 2272 -487 2280 -453
rect 2272 -521 2314 -487
rect 2272 -555 2280 -521
rect 2272 -589 2314 -555
rect 2272 -623 2280 -589
rect 2272 -665 2314 -623
rect 2348 -453 2414 -435
rect 2861 -437 2914 -400
rect 2348 -487 2364 -453
rect 2398 -487 2414 -453
rect 2348 -521 2414 -487
rect 2348 -555 2364 -521
rect 2398 -555 2414 -521
rect 2348 -589 2414 -555
rect 2348 -623 2364 -589
rect 2398 -623 2414 -589
rect 2348 -631 2414 -623
rect 2506 -453 2559 -437
rect 2506 -487 2525 -453
rect 2506 -521 2559 -487
rect 2506 -555 2525 -521
rect 2506 -589 2559 -555
rect 2506 -623 2525 -589
rect 2506 -665 2559 -623
rect 2593 -453 2914 -437
rect 2593 -487 2609 -453
rect 2643 -471 2777 -453
rect 2643 -487 2659 -471
rect 2593 -521 2659 -487
rect 2761 -487 2777 -471
rect 2811 -475 2914 -453
rect 3207 -467 3265 -432
rect 2811 -487 2827 -475
rect 2593 -555 2609 -521
rect 2643 -555 2659 -521
rect 2593 -589 2659 -555
rect 2593 -623 2609 -589
rect 2643 -623 2659 -589
rect 2593 -631 2659 -623
rect 2693 -521 2727 -505
rect 2693 -589 2727 -555
rect 2693 -665 2727 -623
rect 2761 -521 2827 -487
rect 2761 -555 2777 -521
rect 2811 -555 2827 -521
rect 2761 -589 2827 -555
rect 3207 -501 3219 -467
rect 3253 -501 3265 -467
rect 3207 -560 3265 -501
rect 2761 -623 2777 -589
rect 2811 -623 2827 -589
rect 2761 -631 2827 -623
rect 2861 -589 2903 -573
rect 2895 -623 2903 -589
rect 2861 -665 2903 -623
rect 3207 -594 3219 -560
rect 3253 -594 3265 -560
rect 3207 -665 3265 -594
rect -2584 -699 -2555 -665
rect -2521 -699 -2492 -665
rect -2242 -699 -2213 -665
rect -2179 -699 -2121 -665
rect -2087 -699 -2029 -665
rect -1995 -699 -1937 -665
rect -1903 -699 -1845 -665
rect -1811 -699 -1753 -665
rect -1719 -699 -1661 -665
rect -1627 -699 -1569 -665
rect -1535 -699 -1477 -665
rect -1443 -699 -1385 -665
rect -1351 -699 -1293 -665
rect -1259 -699 -1201 -665
rect -1167 -699 -1109 -665
rect -1075 -699 -1017 -665
rect -983 -699 -925 -665
rect -891 -699 -833 -665
rect -799 -699 -741 -665
rect -707 -699 -649 -665
rect -615 -699 -557 -665
rect -523 -699 -465 -665
rect -431 -699 -373 -665
rect -339 -699 -281 -665
rect -247 -699 -189 -665
rect -155 -699 -97 -665
rect -63 -699 -5 -665
rect 29 -699 87 -665
rect 121 -699 179 -665
rect 213 -699 242 -665
rect 456 -699 485 -665
rect 519 -699 577 -665
rect 611 -699 669 -665
rect 703 -699 761 -665
rect 795 -699 853 -665
rect 887 -699 945 -665
rect 979 -699 1037 -665
rect 1071 -699 1129 -665
rect 1163 -699 1221 -665
rect 1255 -699 1313 -665
rect 1347 -699 1405 -665
rect 1439 -699 1497 -665
rect 1531 -699 1589 -665
rect 1623 -699 1681 -665
rect 1715 -699 1773 -665
rect 1807 -699 1865 -665
rect 1899 -699 1957 -665
rect 1991 -699 2049 -665
rect 2083 -699 2141 -665
rect 2175 -699 2233 -665
rect 2267 -699 2325 -665
rect 2359 -699 2417 -665
rect 2451 -699 2509 -665
rect 2543 -699 2601 -665
rect 2635 -699 2693 -665
rect 2727 -699 2785 -665
rect 2819 -699 2877 -665
rect 2911 -699 2940 -665
rect 3190 -699 3219 -665
rect 3253 -699 3282 -665
rect -2567 -770 -2509 -699
rect -2567 -804 -2555 -770
rect -2521 -804 -2509 -770
rect -2567 -863 -2509 -804
rect -2567 -897 -2555 -863
rect -2521 -897 -2509 -863
rect -2207 -749 -2173 -733
rect -2207 -817 -2173 -783
rect -2139 -765 -2073 -699
rect -2139 -799 -2123 -765
rect -2089 -799 -2073 -765
rect -2039 -749 -2002 -733
rect -2005 -783 -2002 -749
rect -2039 -817 -2002 -783
rect -1954 -741 -1901 -699
rect -1954 -775 -1935 -741
rect -1954 -791 -1901 -775
rect -1867 -749 -1817 -733
rect -1867 -783 -1851 -749
rect -1520 -741 -1486 -699
rect -2173 -835 -2074 -833
rect -2173 -851 -2116 -835
rect -2207 -867 -2116 -851
rect -2567 -932 -2509 -897
rect -2120 -869 -2116 -867
rect -2082 -869 -2074 -835
rect -2224 -910 -2154 -901
rect -2224 -958 -2218 -910
rect -2170 -958 -2154 -910
rect -2224 -977 -2154 -958
rect -2224 -1011 -2210 -977
rect -2176 -1011 -2154 -977
rect -2224 -1031 -2154 -1011
rect -2120 -962 -2074 -869
rect -2120 -996 -2108 -962
rect -2567 -1081 -2509 -1064
rect -2120 -1065 -2074 -996
rect -2567 -1115 -2555 -1081
rect -2521 -1115 -2509 -1081
rect -2567 -1209 -2509 -1115
rect -2207 -1099 -2074 -1065
rect -2005 -851 -2002 -817
rect -1867 -818 -1817 -783
rect -1775 -788 -1759 -754
rect -1725 -788 -1554 -754
rect -2039 -903 -2002 -851
rect -1878 -844 -1817 -818
rect -1728 -835 -1622 -822
rect -2039 -937 -2037 -903
rect -2003 -937 -2002 -903
rect -2207 -1107 -2173 -1099
rect -2039 -1107 -2002 -937
rect -1968 -909 -1912 -893
rect -1968 -943 -1946 -909
rect -1968 -1000 -1912 -943
rect -1968 -1048 -1962 -1000
rect -1914 -1048 -1912 -1000
rect -1968 -1083 -1912 -1048
rect -1878 -1065 -1844 -844
rect -1728 -869 -1696 -835
rect -1662 -861 -1622 -835
rect -1810 -903 -1762 -882
rect -1810 -937 -1799 -903
rect -1765 -937 -1762 -903
rect -1810 -939 -1762 -937
rect -1810 -973 -1803 -939
rect -1769 -973 -1762 -939
rect -1810 -1001 -1762 -973
rect -1728 -1035 -1694 -869
rect -1660 -895 -1622 -861
rect -1588 -911 -1554 -788
rect -1520 -809 -1486 -775
rect -1520 -859 -1486 -843
rect -1452 -749 -1402 -733
rect -1452 -783 -1436 -749
rect -1144 -749 -1081 -699
rect -1452 -799 -1402 -783
rect -1357 -793 -1341 -759
rect -1307 -793 -1180 -759
rect -1588 -927 -1486 -911
rect -1588 -929 -1520 -927
rect -1878 -1091 -1833 -1065
rect -1799 -1069 -1783 -1035
rect -1749 -1069 -1694 -1035
rect -1799 -1079 -1694 -1069
rect -1660 -961 -1520 -929
rect -1660 -963 -1486 -961
rect -2207 -1157 -2173 -1141
rect -2139 -1167 -2123 -1133
rect -2089 -1167 -2073 -1133
rect -2005 -1141 -2002 -1107
rect -2039 -1157 -2002 -1141
rect -1951 -1133 -1901 -1117
rect -2139 -1209 -2073 -1167
rect -1951 -1167 -1935 -1133
rect -1867 -1119 -1833 -1091
rect -1660 -1119 -1626 -963
rect -1520 -977 -1486 -963
rect -1584 -1013 -1544 -1007
rect -1452 -1013 -1418 -799
rect -1384 -835 -1346 -833
rect -1384 -869 -1382 -835
rect -1348 -869 -1346 -835
rect -1384 -927 -1346 -869
rect -1350 -961 -1346 -927
rect -1384 -977 -1346 -961
rect -1312 -861 -1248 -827
rect -1312 -895 -1282 -861
rect -1312 -903 -1248 -895
rect -1312 -937 -1295 -903
rect -1261 -937 -1248 -903
rect -1584 -1023 -1418 -1013
rect -1312 -1019 -1248 -937
rect -1550 -1057 -1418 -1023
rect -1584 -1073 -1418 -1057
rect -1867 -1153 -1850 -1119
rect -1816 -1153 -1800 -1119
rect -1761 -1153 -1739 -1119
rect -1705 -1153 -1626 -1119
rect -1562 -1125 -1488 -1109
rect -1951 -1209 -1901 -1167
rect -1562 -1159 -1540 -1125
rect -1506 -1159 -1488 -1125
rect -1452 -1119 -1418 -1073
rect -1341 -1035 -1248 -1019
rect -1307 -1069 -1248 -1035
rect -1341 -1085 -1248 -1069
rect -1214 -961 -1180 -793
rect -1144 -783 -1142 -749
rect -1108 -783 -1081 -749
rect -1144 -799 -1081 -783
rect -1034 -741 -966 -733
rect -1034 -775 -1018 -741
rect -984 -775 -966 -741
rect -1034 -812 -966 -775
rect -1034 -845 -1018 -812
rect -1146 -846 -1018 -845
rect -984 -846 -966 -812
rect -1146 -861 -966 -846
rect -1112 -883 -966 -861
rect -1112 -895 -1018 -883
rect -1146 -917 -1018 -895
rect -984 -917 -966 -883
rect -932 -771 -898 -699
rect -760 -741 -694 -737
rect -932 -851 -898 -805
rect -932 -901 -898 -885
rect -864 -747 -798 -742
rect -864 -781 -848 -747
rect -814 -781 -798 -747
rect -864 -815 -798 -781
rect -864 -849 -848 -815
rect -814 -849 -798 -815
rect -864 -883 -798 -849
rect -760 -775 -744 -741
rect -710 -775 -694 -741
rect -760 -809 -694 -775
rect -760 -843 -744 -809
rect -710 -843 -694 -809
rect -760 -883 -694 -843
rect -1146 -920 -966 -917
rect -1004 -961 -966 -920
rect -864 -917 -848 -883
rect -814 -911 -798 -883
rect -814 -917 -782 -911
rect -864 -927 -782 -917
rect -829 -937 -782 -927
rect -1214 -977 -1038 -961
rect -1214 -1011 -1072 -977
rect -1214 -1027 -1038 -1011
rect -1004 -977 -854 -961
rect -1004 -1011 -888 -977
rect -1004 -1027 -854 -1011
rect -1214 -1119 -1180 -1027
rect -1004 -1061 -964 -1027
rect -820 -1053 -782 -937
rect -831 -1061 -782 -1053
rect -1030 -1064 -964 -1061
rect -1030 -1098 -1014 -1064
rect -980 -1098 -964 -1064
rect -862 -1062 -782 -1061
rect -862 -1082 -846 -1062
rect -812 -1078 -782 -1062
rect -748 -961 -694 -883
rect -656 -741 -613 -699
rect -656 -775 -647 -741
rect -656 -809 -613 -775
rect -656 -843 -647 -809
rect -656 -877 -613 -843
rect -656 -911 -647 -877
rect -656 -927 -613 -911
rect -579 -741 -512 -733
rect -579 -775 -563 -741
rect -529 -775 -512 -741
rect -579 -812 -512 -775
rect -579 -846 -563 -812
rect -529 -846 -512 -812
rect -579 -883 -512 -846
rect -579 -917 -563 -883
rect -529 -917 -512 -883
rect -579 -930 -512 -917
rect -426 -741 -384 -699
rect -426 -775 -418 -741
rect -426 -809 -384 -775
rect -426 -843 -418 -809
rect -426 -877 -384 -843
rect -426 -911 -418 -877
rect -426 -927 -384 -911
rect -350 -741 -284 -733
rect -350 -775 -334 -741
rect -300 -775 -284 -741
rect -350 -809 -284 -775
rect -350 -843 -334 -809
rect -300 -843 -284 -809
rect -350 -877 -284 -843
rect -350 -911 -334 -877
rect -300 -911 -284 -877
rect -350 -929 -284 -911
rect -192 -741 -139 -699
rect -192 -775 -173 -741
rect -192 -809 -139 -775
rect -192 -843 -173 -809
rect -192 -877 -139 -843
rect -192 -911 -173 -877
rect -192 -927 -139 -911
rect -105 -741 -39 -733
rect -105 -775 -89 -741
rect -55 -775 -39 -741
rect -105 -809 -39 -775
rect -105 -843 -89 -809
rect -55 -843 -39 -809
rect -105 -877 -39 -843
rect -5 -741 29 -699
rect -5 -809 29 -775
rect -5 -859 29 -843
rect 63 -741 129 -733
rect 63 -775 79 -741
rect 113 -775 129 -741
rect 63 -809 129 -775
rect 163 -741 205 -699
rect 197 -775 205 -741
rect 163 -791 205 -775
rect 491 -749 525 -733
rect 63 -843 79 -809
rect 113 -843 129 -809
rect -105 -911 -89 -877
rect -55 -893 -39 -877
rect 63 -877 129 -843
rect 491 -817 525 -783
rect 559 -765 625 -699
rect 559 -799 575 -765
rect 609 -799 625 -765
rect 659 -749 696 -733
rect 693 -783 696 -749
rect 659 -817 696 -783
rect 744 -741 797 -699
rect 744 -775 763 -741
rect 744 -791 797 -775
rect 831 -749 881 -733
rect 831 -783 847 -749
rect 1178 -741 1212 -699
rect 525 -835 624 -833
rect 525 -851 582 -835
rect 491 -867 582 -851
rect 63 -893 79 -877
rect -55 -911 79 -893
rect 113 -889 129 -877
rect 578 -869 582 -867
rect 616 -869 624 -835
rect 113 -911 216 -889
rect -105 -927 216 -911
rect -748 -977 -593 -961
rect -748 -1011 -627 -977
rect -748 -1027 -593 -1011
rect -559 -962 -512 -930
rect -330 -962 -284 -929
rect -197 -962 129 -961
rect -559 -1010 -552 -962
rect -388 -977 -364 -963
rect -812 -1082 -796 -1078
rect -1452 -1153 -1421 -1119
rect -1387 -1153 -1371 -1119
rect -1337 -1153 -1318 -1119
rect -1284 -1153 -1180 -1119
rect -1125 -1119 -1083 -1103
rect -1125 -1153 -1120 -1119
rect -1086 -1153 -1083 -1119
rect -1562 -1209 -1488 -1159
rect -1125 -1209 -1083 -1153
rect -1030 -1132 -964 -1098
rect -1030 -1166 -1014 -1132
rect -980 -1166 -964 -1132
rect -930 -1103 -896 -1087
rect -930 -1209 -896 -1137
rect -862 -1130 -858 -1082
rect -810 -1130 -796 -1082
rect -748 -1103 -708 -1027
rect -559 -1044 -512 -1010
rect -430 -1011 -414 -1010
rect -380 -1011 -364 -977
rect -330 -1010 -324 -962
rect -197 -1010 -192 -962
rect -144 -977 -82 -962
rect -34 -977 34 -962
rect 82 -977 129 -962
rect -144 -1010 -89 -977
rect -34 -1010 -5 -977
rect -862 -1164 -846 -1130
rect -812 -1164 -796 -1130
rect -758 -1107 -708 -1103
rect -758 -1141 -742 -1107
rect -563 -1095 -512 -1044
rect -758 -1157 -708 -1141
rect -661 -1133 -597 -1117
rect -862 -1165 -796 -1164
rect -661 -1167 -647 -1133
rect -613 -1167 -597 -1133
rect -661 -1209 -597 -1167
rect -529 -1129 -512 -1095
rect -563 -1175 -512 -1129
rect -430 -1061 -384 -1045
rect -330 -1049 -284 -1010
rect -197 -1011 -181 -1010
rect -147 -1011 -89 -1010
rect -55 -1011 -5 -1010
rect 29 -1010 34 -977
rect 29 -1011 79 -1010
rect 113 -1011 129 -977
rect 163 -964 216 -927
rect 474 -950 544 -901
rect 163 -1012 166 -964
rect 474 -998 480 -950
rect 528 -998 544 -950
rect 474 -1011 488 -998
rect 522 -1011 544 -998
rect 163 -1045 216 -1012
rect 474 -1031 544 -1011
rect 578 -962 624 -869
rect 578 -996 590 -962
rect -430 -1095 -418 -1061
rect -430 -1129 -384 -1095
rect -430 -1163 -418 -1129
rect -430 -1209 -384 -1163
rect -350 -1061 -284 -1049
rect -350 -1095 -334 -1061
rect -300 -1095 -284 -1061
rect -350 -1129 -284 -1095
rect -105 -1081 216 -1045
rect 578 -1065 624 -996
rect -350 -1163 -334 -1129
rect -300 -1163 -284 -1129
rect -350 -1175 -284 -1163
rect -192 -1133 -139 -1117
rect -192 -1167 -173 -1133
rect -192 -1209 -139 -1167
rect -105 -1125 -39 -1081
rect -105 -1159 -89 -1125
rect -55 -1159 -39 -1125
rect -105 -1175 -39 -1159
rect -5 -1133 29 -1117
rect -5 -1209 29 -1167
rect 63 -1125 129 -1081
rect 491 -1099 624 -1065
rect 693 -851 696 -817
rect 831 -818 881 -783
rect 923 -788 939 -754
rect 973 -788 1144 -754
rect 659 -903 696 -851
rect 820 -844 881 -818
rect 970 -835 1076 -822
rect 659 -937 661 -903
rect 695 -937 696 -903
rect 491 -1107 525 -1099
rect 63 -1159 79 -1125
rect 113 -1159 129 -1125
rect 63 -1175 129 -1159
rect 163 -1132 213 -1116
rect 197 -1166 213 -1132
rect 659 -1107 696 -937
rect 730 -909 786 -893
rect 730 -943 752 -909
rect 730 -1000 786 -943
rect 730 -1048 736 -1000
rect 784 -1048 786 -1000
rect 730 -1083 786 -1048
rect 820 -1065 854 -844
rect 970 -869 1002 -835
rect 1036 -861 1076 -835
rect 888 -903 936 -882
rect 888 -937 899 -903
rect 933 -937 936 -903
rect 888 -939 936 -937
rect 888 -973 895 -939
rect 929 -973 936 -939
rect 888 -1001 936 -973
rect 970 -1035 1004 -869
rect 1038 -895 1076 -861
rect 1110 -911 1144 -788
rect 1178 -809 1212 -775
rect 1178 -859 1212 -843
rect 1246 -749 1296 -733
rect 1246 -783 1262 -749
rect 1554 -749 1617 -699
rect 1246 -799 1296 -783
rect 1341 -793 1357 -759
rect 1391 -793 1518 -759
rect 1110 -927 1212 -911
rect 1110 -929 1178 -927
rect 820 -1091 865 -1065
rect 899 -1069 915 -1035
rect 949 -1069 1004 -1035
rect 899 -1079 1004 -1069
rect 1038 -961 1178 -929
rect 1038 -963 1212 -961
rect 491 -1157 525 -1141
rect 163 -1209 213 -1166
rect 559 -1167 575 -1133
rect 609 -1167 625 -1133
rect 693 -1141 696 -1107
rect 659 -1157 696 -1141
rect 747 -1133 797 -1117
rect 559 -1209 625 -1167
rect 747 -1167 763 -1133
rect 831 -1119 865 -1091
rect 1038 -1119 1072 -963
rect 1178 -977 1212 -963
rect 1114 -1013 1154 -1007
rect 1246 -1013 1280 -799
rect 1314 -835 1352 -833
rect 1314 -869 1316 -835
rect 1350 -869 1352 -835
rect 1314 -927 1352 -869
rect 1348 -961 1352 -927
rect 1314 -977 1352 -961
rect 1386 -861 1450 -827
rect 1386 -895 1416 -861
rect 1386 -903 1450 -895
rect 1386 -937 1403 -903
rect 1437 -937 1450 -903
rect 1114 -1023 1280 -1013
rect 1386 -1019 1450 -937
rect 1148 -1057 1280 -1023
rect 1114 -1073 1280 -1057
rect 831 -1153 848 -1119
rect 882 -1153 898 -1119
rect 937 -1153 959 -1119
rect 993 -1153 1072 -1119
rect 1136 -1125 1210 -1109
rect 747 -1209 797 -1167
rect 1136 -1159 1158 -1125
rect 1192 -1159 1210 -1125
rect 1246 -1119 1280 -1073
rect 1357 -1035 1450 -1019
rect 1391 -1069 1450 -1035
rect 1357 -1085 1450 -1069
rect 1484 -961 1518 -793
rect 1554 -783 1556 -749
rect 1590 -783 1617 -749
rect 1554 -799 1617 -783
rect 1664 -741 1732 -733
rect 1664 -775 1680 -741
rect 1714 -775 1732 -741
rect 1664 -812 1732 -775
rect 1664 -845 1680 -812
rect 1552 -846 1680 -845
rect 1714 -846 1732 -812
rect 1552 -861 1732 -846
rect 1586 -883 1732 -861
rect 1586 -895 1680 -883
rect 1552 -917 1680 -895
rect 1714 -917 1732 -883
rect 1766 -771 1800 -699
rect 1938 -741 2004 -737
rect 1766 -851 1800 -805
rect 1766 -901 1800 -885
rect 1834 -747 1900 -742
rect 1834 -778 1850 -747
rect 1884 -778 1900 -747
rect 1834 -826 1840 -778
rect 1888 -826 1900 -778
rect 1834 -849 1850 -826
rect 1884 -849 1900 -826
rect 1834 -883 1900 -849
rect 1938 -775 1954 -741
rect 1988 -775 2004 -741
rect 1938 -809 2004 -775
rect 1938 -843 1954 -809
rect 1988 -843 2004 -809
rect 1938 -883 2004 -843
rect 1552 -920 1732 -917
rect 1694 -961 1732 -920
rect 1834 -917 1850 -883
rect 1884 -911 1900 -883
rect 1884 -917 1916 -911
rect 1834 -927 1916 -917
rect 1869 -937 1916 -927
rect 1484 -977 1660 -961
rect 1484 -1011 1626 -977
rect 1484 -1027 1660 -1011
rect 1694 -977 1844 -961
rect 1694 -1011 1810 -977
rect 1694 -1027 1844 -1011
rect 1484 -1119 1518 -1027
rect 1694 -1061 1734 -1027
rect 1878 -1053 1916 -937
rect 1867 -1061 1916 -1053
rect 1668 -1064 1734 -1061
rect 1668 -1098 1684 -1064
rect 1718 -1098 1734 -1064
rect 1836 -1062 1916 -1061
rect 1246 -1153 1277 -1119
rect 1311 -1153 1327 -1119
rect 1361 -1153 1380 -1119
rect 1414 -1153 1518 -1119
rect 1573 -1119 1615 -1103
rect 1573 -1153 1578 -1119
rect 1612 -1153 1615 -1119
rect 1136 -1209 1210 -1159
rect 1573 -1209 1615 -1153
rect 1668 -1132 1734 -1098
rect 1668 -1166 1684 -1132
rect 1718 -1166 1734 -1132
rect 1768 -1103 1802 -1087
rect 1768 -1209 1802 -1137
rect 1836 -1096 1852 -1062
rect 1886 -1078 1916 -1062
rect 1950 -961 2004 -883
rect 2042 -741 2085 -699
rect 2042 -775 2051 -741
rect 2042 -809 2085 -775
rect 2042 -843 2051 -809
rect 2042 -877 2085 -843
rect 2042 -911 2051 -877
rect 2042 -927 2085 -911
rect 2119 -741 2186 -733
rect 2119 -775 2135 -741
rect 2169 -775 2186 -741
rect 2119 -812 2186 -775
rect 2119 -846 2135 -812
rect 2169 -846 2186 -812
rect 2119 -883 2186 -846
rect 2119 -917 2135 -883
rect 2169 -917 2186 -883
rect 2119 -930 2186 -917
rect 2272 -741 2314 -699
rect 2272 -775 2280 -741
rect 2272 -809 2314 -775
rect 2272 -843 2280 -809
rect 2272 -877 2314 -843
rect 2272 -911 2280 -877
rect 2272 -927 2314 -911
rect 2348 -741 2414 -733
rect 2348 -775 2364 -741
rect 2398 -775 2414 -741
rect 2348 -809 2414 -775
rect 2348 -843 2364 -809
rect 2398 -843 2414 -809
rect 2348 -877 2414 -843
rect 2348 -911 2364 -877
rect 2398 -911 2414 -877
rect 2348 -929 2414 -911
rect 2506 -741 2559 -699
rect 2506 -775 2525 -741
rect 2506 -809 2559 -775
rect 2506 -843 2525 -809
rect 2506 -877 2559 -843
rect 2506 -911 2525 -877
rect 2506 -927 2559 -911
rect 2593 -741 2659 -733
rect 2593 -775 2609 -741
rect 2643 -775 2659 -741
rect 2593 -809 2659 -775
rect 2593 -843 2609 -809
rect 2643 -843 2659 -809
rect 2593 -877 2659 -843
rect 2693 -741 2727 -699
rect 2693 -809 2727 -775
rect 2693 -859 2727 -843
rect 2761 -741 2827 -733
rect 2761 -775 2777 -741
rect 2811 -775 2827 -741
rect 2761 -809 2827 -775
rect 2861 -741 2903 -699
rect 2895 -775 2903 -741
rect 2861 -791 2903 -775
rect 3207 -770 3265 -699
rect 2761 -843 2777 -809
rect 2811 -843 2827 -809
rect 2593 -911 2609 -877
rect 2643 -893 2659 -877
rect 2761 -877 2827 -843
rect 2761 -893 2777 -877
rect 2643 -911 2777 -893
rect 2811 -889 2827 -877
rect 3207 -804 3219 -770
rect 3253 -804 3265 -770
rect 3207 -863 3265 -804
rect 2811 -911 2914 -889
rect 2593 -927 2914 -911
rect 1950 -977 2105 -961
rect 1950 -1011 2071 -977
rect 1950 -1027 2105 -1011
rect 2139 -962 2186 -930
rect 2368 -962 2414 -929
rect 2501 -962 2827 -961
rect 2139 -1010 2146 -962
rect 2310 -977 2334 -963
rect 1886 -1096 1902 -1078
rect 1836 -1130 1902 -1096
rect 1950 -1103 1990 -1027
rect 2139 -1044 2186 -1010
rect 2268 -1011 2284 -1010
rect 2318 -1011 2334 -977
rect 2368 -1010 2374 -962
rect 2501 -1010 2506 -962
rect 2554 -977 2616 -962
rect 2664 -977 2732 -962
rect 2780 -977 2827 -962
rect 2554 -1010 2609 -977
rect 2664 -1010 2693 -977
rect 1836 -1164 1852 -1130
rect 1886 -1164 1902 -1130
rect 1940 -1107 1990 -1103
rect 1940 -1141 1956 -1107
rect 2135 -1095 2186 -1044
rect 1940 -1157 1990 -1141
rect 2037 -1133 2101 -1117
rect 1836 -1165 1902 -1164
rect 2037 -1167 2051 -1133
rect 2085 -1167 2101 -1133
rect 2037 -1209 2101 -1167
rect 2169 -1129 2186 -1095
rect 2135 -1175 2186 -1129
rect 2268 -1061 2314 -1045
rect 2368 -1049 2414 -1010
rect 2501 -1011 2517 -1010
rect 2551 -1011 2609 -1010
rect 2643 -1011 2693 -1010
rect 2727 -1010 2732 -977
rect 2727 -1011 2777 -1010
rect 2811 -1011 2827 -977
rect 2861 -964 2914 -927
rect 3207 -897 3219 -863
rect 3253 -897 3265 -863
rect 3207 -932 3265 -897
rect 2861 -1012 2864 -964
rect 2912 -1012 2914 -964
rect 2861 -1045 2914 -1012
rect 2268 -1095 2280 -1061
rect 2268 -1129 2314 -1095
rect 2268 -1163 2280 -1129
rect 2268 -1209 2314 -1163
rect 2348 -1061 2414 -1049
rect 2348 -1095 2364 -1061
rect 2398 -1095 2414 -1061
rect 2348 -1129 2414 -1095
rect 2593 -1081 2914 -1045
rect 3207 -1081 3265 -1064
rect 2348 -1163 2364 -1129
rect 2398 -1163 2414 -1129
rect 2348 -1175 2414 -1163
rect 2506 -1133 2559 -1117
rect 2506 -1167 2525 -1133
rect 2506 -1209 2559 -1167
rect 2593 -1125 2659 -1081
rect 2593 -1159 2609 -1125
rect 2643 -1159 2659 -1125
rect 2593 -1175 2659 -1159
rect 2693 -1133 2727 -1117
rect 2693 -1209 2727 -1167
rect 2761 -1125 2827 -1081
rect 3207 -1115 3219 -1081
rect 3253 -1115 3265 -1081
rect 2761 -1159 2777 -1125
rect 2811 -1159 2827 -1125
rect 2761 -1175 2827 -1159
rect 2861 -1132 2911 -1116
rect 2895 -1166 2911 -1132
rect 2861 -1209 2911 -1166
rect 3207 -1209 3265 -1115
rect -2584 -1243 -2555 -1209
rect -2521 -1243 -2492 -1209
rect -2242 -1243 -2213 -1209
rect -2179 -1243 -2121 -1209
rect -2087 -1243 -2029 -1209
rect -1995 -1243 -1937 -1209
rect -1903 -1243 -1845 -1209
rect -1811 -1243 -1753 -1209
rect -1719 -1243 -1661 -1209
rect -1627 -1243 -1569 -1209
rect -1535 -1243 -1477 -1209
rect -1443 -1243 -1385 -1209
rect -1351 -1243 -1293 -1209
rect -1259 -1243 -1201 -1209
rect -1167 -1243 -1109 -1209
rect -1075 -1243 -1017 -1209
rect -983 -1243 -925 -1209
rect -891 -1243 -833 -1209
rect -799 -1243 -741 -1209
rect -707 -1243 -649 -1209
rect -615 -1243 -557 -1209
rect -523 -1243 -465 -1209
rect -431 -1243 -373 -1209
rect -339 -1243 -281 -1209
rect -247 -1243 -189 -1209
rect -155 -1243 -97 -1209
rect -63 -1243 -5 -1209
rect 29 -1243 87 -1209
rect 121 -1243 179 -1209
rect 213 -1243 242 -1209
rect 456 -1243 485 -1209
rect 519 -1243 577 -1209
rect 611 -1243 669 -1209
rect 703 -1243 761 -1209
rect 795 -1243 853 -1209
rect 887 -1243 945 -1209
rect 979 -1243 1037 -1209
rect 1071 -1243 1129 -1209
rect 1163 -1243 1221 -1209
rect 1255 -1243 1313 -1209
rect 1347 -1243 1405 -1209
rect 1439 -1243 1497 -1209
rect 1531 -1243 1589 -1209
rect 1623 -1243 1681 -1209
rect 1715 -1243 1773 -1209
rect 1807 -1243 1865 -1209
rect 1899 -1243 1957 -1209
rect 1991 -1243 2049 -1209
rect 2083 -1243 2141 -1209
rect 2175 -1243 2233 -1209
rect 2267 -1243 2325 -1209
rect 2359 -1243 2417 -1209
rect 2451 -1243 2509 -1209
rect 2543 -1243 2601 -1209
rect 2635 -1243 2693 -1209
rect 2727 -1243 2785 -1209
rect 2819 -1243 2877 -1209
rect 2911 -1243 2940 -1209
rect 3190 -1243 3219 -1209
rect 3253 -1243 3282 -1209
rect -2567 -1337 -2509 -1243
rect -2139 -1285 -2073 -1243
rect -2567 -1371 -2555 -1337
rect -2521 -1371 -2509 -1337
rect -2567 -1388 -2509 -1371
rect -2207 -1311 -2173 -1295
rect -2139 -1319 -2123 -1285
rect -2089 -1319 -2073 -1285
rect -1951 -1285 -1901 -1243
rect -2039 -1311 -2002 -1295
rect -2207 -1353 -2173 -1345
rect -2005 -1345 -2002 -1311
rect -1951 -1319 -1935 -1285
rect -1562 -1293 -1488 -1243
rect -1951 -1335 -1901 -1319
rect -1867 -1333 -1850 -1299
rect -1816 -1333 -1800 -1299
rect -1761 -1333 -1739 -1299
rect -1705 -1333 -1626 -1299
rect -2207 -1387 -2074 -1353
rect -2224 -1441 -2154 -1421
rect -2224 -1454 -2210 -1441
rect -2176 -1454 -2154 -1441
rect -2224 -1502 -2218 -1454
rect -2170 -1502 -2154 -1454
rect -2567 -1555 -2509 -1520
rect -2224 -1551 -2154 -1502
rect -2120 -1456 -2074 -1387
rect -2120 -1490 -2108 -1456
rect -2567 -1589 -2555 -1555
rect -2521 -1589 -2509 -1555
rect -2120 -1583 -2074 -1490
rect -2120 -1585 -2116 -1583
rect -2567 -1648 -2509 -1589
rect -2567 -1682 -2555 -1648
rect -2521 -1682 -2509 -1648
rect -2567 -1753 -2509 -1682
rect -2207 -1601 -2116 -1585
rect -2173 -1617 -2116 -1601
rect -2082 -1617 -2074 -1583
rect -2173 -1619 -2074 -1617
rect -2039 -1515 -2002 -1345
rect -1867 -1361 -1833 -1333
rect -2039 -1549 -2037 -1515
rect -2003 -1549 -2002 -1515
rect -2039 -1601 -2002 -1549
rect -1968 -1404 -1912 -1369
rect -1968 -1452 -1962 -1404
rect -1914 -1452 -1912 -1404
rect -1968 -1509 -1912 -1452
rect -1968 -1543 -1946 -1509
rect -1968 -1559 -1912 -1543
rect -1878 -1387 -1833 -1361
rect -1799 -1383 -1694 -1373
rect -2207 -1669 -2173 -1635
rect -2005 -1635 -2002 -1601
rect -1878 -1608 -1844 -1387
rect -1799 -1417 -1783 -1383
rect -1749 -1417 -1694 -1383
rect -1810 -1479 -1762 -1451
rect -1810 -1513 -1803 -1479
rect -1769 -1513 -1762 -1479
rect -1810 -1515 -1762 -1513
rect -1810 -1549 -1799 -1515
rect -1765 -1549 -1762 -1515
rect -1810 -1570 -1762 -1549
rect -1728 -1583 -1694 -1417
rect -1660 -1489 -1626 -1333
rect -1562 -1327 -1540 -1293
rect -1506 -1327 -1488 -1293
rect -1125 -1299 -1083 -1243
rect -1562 -1343 -1488 -1327
rect -1452 -1333 -1421 -1299
rect -1387 -1333 -1371 -1299
rect -1337 -1333 -1318 -1299
rect -1284 -1333 -1180 -1299
rect -1452 -1379 -1418 -1333
rect -1584 -1395 -1418 -1379
rect -1550 -1429 -1418 -1395
rect -1584 -1439 -1418 -1429
rect -1341 -1383 -1248 -1367
rect -1307 -1417 -1248 -1383
rect -1341 -1433 -1248 -1417
rect -1584 -1445 -1544 -1439
rect -1520 -1489 -1486 -1475
rect -1660 -1491 -1486 -1489
rect -1660 -1523 -1520 -1491
rect -1588 -1525 -1520 -1523
rect -1588 -1541 -1486 -1525
rect -1878 -1634 -1817 -1608
rect -1728 -1617 -1696 -1583
rect -1660 -1591 -1622 -1557
rect -1662 -1617 -1622 -1591
rect -1728 -1630 -1622 -1617
rect -2207 -1719 -2173 -1703
rect -2139 -1687 -2123 -1653
rect -2089 -1687 -2073 -1653
rect -2139 -1753 -2073 -1687
rect -2039 -1669 -2002 -1635
rect -2005 -1703 -2002 -1669
rect -2039 -1719 -2002 -1703
rect -1954 -1677 -1901 -1661
rect -1954 -1711 -1935 -1677
rect -1954 -1753 -1901 -1711
rect -1867 -1669 -1817 -1634
rect -1588 -1664 -1554 -1541
rect -1867 -1703 -1851 -1669
rect -1775 -1698 -1759 -1664
rect -1725 -1698 -1554 -1664
rect -1520 -1609 -1486 -1593
rect -1520 -1677 -1486 -1643
rect -1867 -1719 -1817 -1703
rect -1520 -1753 -1486 -1711
rect -1452 -1653 -1418 -1439
rect -1384 -1491 -1346 -1475
rect -1350 -1525 -1346 -1491
rect -1384 -1583 -1346 -1525
rect -1384 -1617 -1382 -1583
rect -1348 -1617 -1346 -1583
rect -1384 -1619 -1346 -1617
rect -1312 -1515 -1248 -1433
rect -1312 -1549 -1295 -1515
rect -1261 -1549 -1248 -1515
rect -1312 -1557 -1248 -1549
rect -1312 -1591 -1282 -1557
rect -1312 -1625 -1248 -1591
rect -1214 -1425 -1180 -1333
rect -1125 -1333 -1120 -1299
rect -1086 -1333 -1083 -1299
rect -1125 -1349 -1083 -1333
rect -1030 -1320 -1014 -1286
rect -980 -1320 -964 -1286
rect -1030 -1354 -964 -1320
rect -1030 -1388 -1014 -1354
rect -980 -1388 -964 -1354
rect -930 -1315 -896 -1243
rect -661 -1285 -597 -1243
rect -930 -1365 -896 -1349
rect -862 -1288 -796 -1287
rect -862 -1322 -846 -1288
rect -812 -1322 -796 -1288
rect -862 -1356 -796 -1322
rect -758 -1311 -708 -1295
rect -758 -1345 -742 -1311
rect -661 -1319 -647 -1285
rect -613 -1319 -597 -1285
rect -661 -1335 -597 -1319
rect -563 -1323 -512 -1277
rect -758 -1349 -708 -1345
rect -1030 -1391 -964 -1388
rect -862 -1390 -846 -1356
rect -812 -1374 -796 -1356
rect -812 -1390 -782 -1374
rect -862 -1391 -782 -1390
rect -1004 -1425 -964 -1391
rect -831 -1399 -782 -1391
rect -1214 -1441 -1038 -1425
rect -1214 -1475 -1072 -1441
rect -1214 -1491 -1038 -1475
rect -1004 -1441 -854 -1425
rect -1004 -1475 -888 -1441
rect -1004 -1491 -854 -1475
rect -1452 -1669 -1402 -1653
rect -1214 -1659 -1180 -1491
rect -1004 -1532 -966 -1491
rect -820 -1515 -782 -1399
rect -829 -1525 -782 -1515
rect -1146 -1535 -966 -1532
rect -1146 -1557 -1018 -1535
rect -1112 -1569 -1018 -1557
rect -984 -1569 -966 -1535
rect -864 -1535 -782 -1525
rect -1112 -1591 -966 -1569
rect -1146 -1606 -966 -1591
rect -1146 -1607 -1018 -1606
rect -1034 -1640 -1018 -1607
rect -984 -1640 -966 -1606
rect -1452 -1703 -1436 -1669
rect -1357 -1693 -1341 -1659
rect -1307 -1693 -1180 -1659
rect -1144 -1669 -1081 -1653
rect -1452 -1719 -1402 -1703
rect -1144 -1703 -1142 -1669
rect -1108 -1703 -1081 -1669
rect -1144 -1753 -1081 -1703
rect -1034 -1677 -966 -1640
rect -1034 -1711 -1018 -1677
rect -984 -1711 -966 -1677
rect -1034 -1719 -966 -1711
rect -932 -1567 -898 -1551
rect -932 -1647 -898 -1601
rect -932 -1753 -898 -1681
rect -864 -1569 -848 -1535
rect -814 -1541 -782 -1535
rect -748 -1425 -708 -1349
rect -529 -1357 -512 -1323
rect -563 -1408 -512 -1357
rect -430 -1289 -384 -1243
rect -430 -1323 -418 -1289
rect -430 -1357 -384 -1323
rect -430 -1391 -418 -1357
rect -430 -1407 -384 -1391
rect -350 -1289 -284 -1277
rect -350 -1323 -334 -1289
rect -300 -1323 -284 -1289
rect -350 -1357 -284 -1323
rect -192 -1285 -139 -1243
rect -192 -1319 -173 -1285
rect -192 -1335 -139 -1319
rect -105 -1293 -39 -1277
rect -105 -1327 -89 -1293
rect -55 -1327 -39 -1293
rect -350 -1391 -334 -1357
rect -300 -1391 -284 -1357
rect -350 -1403 -284 -1391
rect -748 -1441 -593 -1425
rect -748 -1475 -627 -1441
rect -748 -1491 -593 -1475
rect -559 -1442 -512 -1408
rect -430 -1442 -414 -1441
rect -559 -1490 -552 -1442
rect -380 -1475 -364 -1441
rect -388 -1489 -364 -1475
rect -330 -1442 -284 -1403
rect -105 -1371 -39 -1327
rect -5 -1285 29 -1243
rect -5 -1335 29 -1319
rect 63 -1293 129 -1277
rect 63 -1327 79 -1293
rect 113 -1327 129 -1293
rect 63 -1371 129 -1327
rect 163 -1286 213 -1243
rect 197 -1320 213 -1286
rect 559 -1285 625 -1243
rect 163 -1336 213 -1320
rect 491 -1311 525 -1295
rect 559 -1319 575 -1285
rect 609 -1319 625 -1285
rect 747 -1285 797 -1243
rect 659 -1311 696 -1295
rect 491 -1353 525 -1345
rect 693 -1345 696 -1311
rect 747 -1319 763 -1285
rect 1136 -1293 1210 -1243
rect 747 -1335 797 -1319
rect 831 -1333 848 -1299
rect 882 -1333 898 -1299
rect 937 -1333 959 -1299
rect 993 -1333 1072 -1299
rect -105 -1407 216 -1371
rect 491 -1387 624 -1353
rect 163 -1440 216 -1407
rect -197 -1442 -181 -1441
rect -147 -1442 -89 -1441
rect -55 -1442 -5 -1441
rect -330 -1490 -324 -1442
rect -197 -1490 -192 -1442
rect -144 -1475 -89 -1442
rect -34 -1475 -5 -1442
rect 29 -1442 79 -1441
rect 29 -1475 34 -1442
rect 113 -1475 129 -1441
rect -144 -1490 -82 -1475
rect -34 -1490 34 -1475
rect 82 -1490 129 -1475
rect -814 -1569 -798 -1541
rect -748 -1569 -694 -1491
rect -559 -1522 -512 -1490
rect -864 -1603 -798 -1569
rect -864 -1626 -848 -1603
rect -814 -1626 -798 -1603
rect -864 -1674 -858 -1626
rect -810 -1674 -798 -1626
rect -864 -1705 -848 -1674
rect -814 -1705 -798 -1674
rect -864 -1710 -798 -1705
rect -760 -1609 -694 -1569
rect -760 -1643 -744 -1609
rect -710 -1643 -694 -1609
rect -760 -1677 -694 -1643
rect -760 -1711 -744 -1677
rect -710 -1711 -694 -1677
rect -760 -1715 -694 -1711
rect -656 -1541 -613 -1525
rect -656 -1575 -647 -1541
rect -656 -1609 -613 -1575
rect -656 -1643 -647 -1609
rect -656 -1677 -613 -1643
rect -656 -1711 -647 -1677
rect -656 -1753 -613 -1711
rect -579 -1535 -512 -1522
rect -330 -1523 -284 -1490
rect -197 -1491 129 -1490
rect 163 -1488 166 -1440
rect 214 -1488 216 -1440
rect -579 -1569 -563 -1535
rect -529 -1569 -512 -1535
rect -579 -1606 -512 -1569
rect -579 -1640 -563 -1606
rect -529 -1640 -512 -1606
rect -579 -1677 -512 -1640
rect -579 -1711 -563 -1677
rect -529 -1711 -512 -1677
rect -579 -1719 -512 -1711
rect -426 -1541 -384 -1525
rect -426 -1575 -418 -1541
rect -426 -1609 -384 -1575
rect -426 -1643 -418 -1609
rect -426 -1677 -384 -1643
rect -426 -1711 -418 -1677
rect -426 -1753 -384 -1711
rect -350 -1541 -284 -1523
rect 163 -1525 216 -1488
rect -350 -1575 -334 -1541
rect -300 -1575 -284 -1541
rect -350 -1609 -284 -1575
rect -350 -1643 -334 -1609
rect -300 -1643 -284 -1609
rect -350 -1677 -284 -1643
rect -350 -1711 -334 -1677
rect -300 -1711 -284 -1677
rect -350 -1719 -284 -1711
rect -192 -1541 -139 -1525
rect -192 -1575 -173 -1541
rect -192 -1609 -139 -1575
rect -192 -1643 -173 -1609
rect -192 -1677 -139 -1643
rect -192 -1711 -173 -1677
rect -192 -1753 -139 -1711
rect -105 -1541 216 -1525
rect -105 -1575 -89 -1541
rect -55 -1559 79 -1541
rect -55 -1575 -39 -1559
rect -105 -1609 -39 -1575
rect 63 -1575 79 -1559
rect 113 -1563 216 -1541
rect 474 -1441 544 -1421
rect 474 -1475 488 -1441
rect 522 -1475 544 -1441
rect 474 -1494 544 -1475
rect 474 -1542 480 -1494
rect 528 -1542 544 -1494
rect 474 -1551 544 -1542
rect 578 -1456 624 -1387
rect 578 -1490 590 -1456
rect 113 -1575 129 -1563
rect -105 -1643 -89 -1609
rect -55 -1643 -39 -1609
rect -105 -1677 -39 -1643
rect -105 -1711 -89 -1677
rect -55 -1711 -39 -1677
rect -105 -1719 -39 -1711
rect -5 -1609 29 -1593
rect -5 -1677 29 -1643
rect -5 -1753 29 -1711
rect 63 -1609 129 -1575
rect 578 -1583 624 -1490
rect 578 -1585 582 -1583
rect 63 -1643 79 -1609
rect 113 -1643 129 -1609
rect 63 -1677 129 -1643
rect 491 -1601 582 -1585
rect 525 -1617 582 -1601
rect 616 -1617 624 -1583
rect 525 -1619 624 -1617
rect 659 -1515 696 -1345
rect 831 -1361 865 -1333
rect 659 -1549 661 -1515
rect 695 -1549 696 -1515
rect 659 -1601 696 -1549
rect 730 -1404 786 -1369
rect 730 -1452 736 -1404
rect 784 -1452 786 -1404
rect 730 -1509 786 -1452
rect 730 -1543 752 -1509
rect 730 -1559 786 -1543
rect 820 -1387 865 -1361
rect 899 -1383 1004 -1373
rect 63 -1711 79 -1677
rect 113 -1711 129 -1677
rect 63 -1719 129 -1711
rect 163 -1677 205 -1661
rect 197 -1711 205 -1677
rect 163 -1753 205 -1711
rect 491 -1669 525 -1635
rect 693 -1635 696 -1601
rect 820 -1608 854 -1387
rect 899 -1417 915 -1383
rect 949 -1417 1004 -1383
rect 888 -1479 936 -1451
rect 888 -1513 895 -1479
rect 929 -1513 936 -1479
rect 888 -1515 936 -1513
rect 888 -1549 899 -1515
rect 933 -1549 936 -1515
rect 888 -1570 936 -1549
rect 970 -1583 1004 -1417
rect 1038 -1489 1072 -1333
rect 1136 -1327 1158 -1293
rect 1192 -1327 1210 -1293
rect 1573 -1299 1615 -1243
rect 1136 -1343 1210 -1327
rect 1246 -1333 1277 -1299
rect 1311 -1333 1327 -1299
rect 1361 -1333 1380 -1299
rect 1414 -1333 1518 -1299
rect 1246 -1379 1280 -1333
rect 1114 -1395 1280 -1379
rect 1148 -1429 1280 -1395
rect 1114 -1439 1280 -1429
rect 1357 -1383 1450 -1367
rect 1391 -1417 1450 -1383
rect 1357 -1433 1450 -1417
rect 1114 -1445 1154 -1439
rect 1178 -1489 1212 -1475
rect 1038 -1491 1212 -1489
rect 1038 -1523 1178 -1491
rect 1110 -1525 1178 -1523
rect 1110 -1541 1212 -1525
rect 820 -1634 881 -1608
rect 970 -1617 1002 -1583
rect 1038 -1591 1076 -1557
rect 1036 -1617 1076 -1591
rect 970 -1630 1076 -1617
rect 491 -1719 525 -1703
rect 559 -1687 575 -1653
rect 609 -1687 625 -1653
rect 559 -1753 625 -1687
rect 659 -1669 696 -1635
rect 693 -1703 696 -1669
rect 659 -1719 696 -1703
rect 744 -1677 797 -1661
rect 744 -1711 763 -1677
rect 744 -1753 797 -1711
rect 831 -1669 881 -1634
rect 1110 -1664 1144 -1541
rect 831 -1703 847 -1669
rect 923 -1698 939 -1664
rect 973 -1698 1144 -1664
rect 1178 -1609 1212 -1593
rect 1178 -1677 1212 -1643
rect 831 -1719 881 -1703
rect 1178 -1753 1212 -1711
rect 1246 -1653 1280 -1439
rect 1314 -1491 1352 -1475
rect 1348 -1525 1352 -1491
rect 1314 -1583 1352 -1525
rect 1314 -1617 1316 -1583
rect 1350 -1617 1352 -1583
rect 1314 -1619 1352 -1617
rect 1386 -1515 1450 -1433
rect 1386 -1549 1403 -1515
rect 1437 -1549 1450 -1515
rect 1386 -1557 1450 -1549
rect 1386 -1591 1416 -1557
rect 1386 -1625 1450 -1591
rect 1484 -1425 1518 -1333
rect 1573 -1333 1578 -1299
rect 1612 -1333 1615 -1299
rect 1573 -1349 1615 -1333
rect 1668 -1320 1684 -1286
rect 1718 -1320 1734 -1286
rect 1668 -1354 1734 -1320
rect 1668 -1388 1684 -1354
rect 1718 -1388 1734 -1354
rect 1768 -1315 1802 -1243
rect 2037 -1285 2101 -1243
rect 1768 -1365 1802 -1349
rect 1836 -1288 1902 -1287
rect 1836 -1322 1852 -1288
rect 1886 -1322 1902 -1288
rect 1668 -1391 1734 -1388
rect 1836 -1370 1840 -1322
rect 1888 -1370 1902 -1322
rect 1940 -1311 1990 -1295
rect 1940 -1345 1956 -1311
rect 2037 -1319 2051 -1285
rect 2085 -1319 2101 -1285
rect 2037 -1335 2101 -1319
rect 2135 -1323 2186 -1277
rect 1940 -1349 1990 -1345
rect 1836 -1390 1852 -1370
rect 1886 -1374 1902 -1370
rect 1886 -1390 1916 -1374
rect 1836 -1391 1916 -1390
rect 1694 -1425 1734 -1391
rect 1867 -1399 1916 -1391
rect 1484 -1441 1660 -1425
rect 1484 -1475 1626 -1441
rect 1484 -1491 1660 -1475
rect 1694 -1441 1844 -1425
rect 1694 -1475 1810 -1441
rect 1694 -1491 1844 -1475
rect 1246 -1669 1296 -1653
rect 1484 -1659 1518 -1491
rect 1694 -1532 1732 -1491
rect 1878 -1515 1916 -1399
rect 1869 -1525 1916 -1515
rect 1552 -1535 1732 -1532
rect 1552 -1557 1680 -1535
rect 1586 -1569 1680 -1557
rect 1714 -1569 1732 -1535
rect 1834 -1535 1916 -1525
rect 1586 -1591 1732 -1569
rect 1552 -1606 1732 -1591
rect 1552 -1607 1680 -1606
rect 1664 -1640 1680 -1607
rect 1714 -1640 1732 -1606
rect 1246 -1703 1262 -1669
rect 1341 -1693 1357 -1659
rect 1391 -1693 1518 -1659
rect 1554 -1669 1617 -1653
rect 1246 -1719 1296 -1703
rect 1554 -1703 1556 -1669
rect 1590 -1703 1617 -1669
rect 1554 -1753 1617 -1703
rect 1664 -1677 1732 -1640
rect 1664 -1711 1680 -1677
rect 1714 -1711 1732 -1677
rect 1664 -1719 1732 -1711
rect 1766 -1567 1800 -1551
rect 1766 -1647 1800 -1601
rect 1766 -1753 1800 -1681
rect 1834 -1569 1850 -1535
rect 1884 -1541 1916 -1535
rect 1950 -1425 1990 -1349
rect 2169 -1357 2186 -1323
rect 2135 -1408 2186 -1357
rect 2268 -1289 2314 -1243
rect 2268 -1323 2280 -1289
rect 2268 -1357 2314 -1323
rect 2268 -1391 2280 -1357
rect 2268 -1407 2314 -1391
rect 2348 -1289 2414 -1277
rect 2348 -1323 2364 -1289
rect 2398 -1323 2414 -1289
rect 2348 -1357 2414 -1323
rect 2506 -1285 2559 -1243
rect 2506 -1319 2525 -1285
rect 2506 -1335 2559 -1319
rect 2593 -1293 2659 -1277
rect 2593 -1327 2609 -1293
rect 2643 -1327 2659 -1293
rect 2348 -1391 2364 -1357
rect 2398 -1391 2414 -1357
rect 2348 -1403 2414 -1391
rect 1950 -1441 2105 -1425
rect 1950 -1475 2071 -1441
rect 1950 -1491 2105 -1475
rect 2139 -1442 2186 -1408
rect 2268 -1442 2284 -1441
rect 2139 -1490 2146 -1442
rect 2318 -1475 2334 -1441
rect 2310 -1489 2334 -1475
rect 2368 -1442 2414 -1403
rect 2593 -1371 2659 -1327
rect 2693 -1285 2727 -1243
rect 2693 -1335 2727 -1319
rect 2761 -1293 2827 -1277
rect 2761 -1327 2777 -1293
rect 2811 -1327 2827 -1293
rect 2761 -1371 2827 -1327
rect 2861 -1286 2911 -1243
rect 2895 -1320 2911 -1286
rect 2861 -1336 2911 -1320
rect 3207 -1337 3265 -1243
rect 3207 -1371 3219 -1337
rect 3253 -1371 3265 -1337
rect 2593 -1407 2914 -1371
rect 3207 -1388 3265 -1371
rect 2861 -1440 2914 -1407
rect 2501 -1442 2517 -1441
rect 2551 -1442 2609 -1441
rect 2643 -1442 2693 -1441
rect 2368 -1490 2374 -1442
rect 2501 -1490 2506 -1442
rect 2554 -1475 2609 -1442
rect 2664 -1475 2693 -1442
rect 2727 -1442 2777 -1441
rect 2727 -1475 2732 -1442
rect 2811 -1475 2827 -1441
rect 2554 -1490 2616 -1475
rect 2664 -1490 2732 -1475
rect 2780 -1490 2827 -1475
rect 1884 -1569 1900 -1541
rect 1950 -1569 2004 -1491
rect 2139 -1522 2186 -1490
rect 1834 -1603 1900 -1569
rect 1834 -1637 1850 -1603
rect 1884 -1637 1900 -1603
rect 1834 -1671 1900 -1637
rect 1834 -1705 1850 -1671
rect 1884 -1705 1900 -1671
rect 1834 -1710 1900 -1705
rect 1938 -1609 2004 -1569
rect 1938 -1643 1954 -1609
rect 1988 -1643 2004 -1609
rect 1938 -1677 2004 -1643
rect 1938 -1711 1954 -1677
rect 1988 -1711 2004 -1677
rect 1938 -1715 2004 -1711
rect 2042 -1541 2085 -1525
rect 2042 -1575 2051 -1541
rect 2042 -1609 2085 -1575
rect 2042 -1643 2051 -1609
rect 2042 -1677 2085 -1643
rect 2042 -1711 2051 -1677
rect 2042 -1753 2085 -1711
rect 2119 -1535 2186 -1522
rect 2368 -1523 2414 -1490
rect 2501 -1491 2827 -1490
rect 2861 -1488 2864 -1440
rect 2119 -1569 2135 -1535
rect 2169 -1569 2186 -1535
rect 2119 -1606 2186 -1569
rect 2119 -1640 2135 -1606
rect 2169 -1640 2186 -1606
rect 2119 -1677 2186 -1640
rect 2119 -1711 2135 -1677
rect 2169 -1711 2186 -1677
rect 2119 -1719 2186 -1711
rect 2272 -1541 2314 -1525
rect 2272 -1575 2280 -1541
rect 2272 -1609 2314 -1575
rect 2272 -1643 2280 -1609
rect 2272 -1677 2314 -1643
rect 2272 -1711 2280 -1677
rect 2272 -1753 2314 -1711
rect 2348 -1541 2414 -1523
rect 2861 -1525 2914 -1488
rect 2348 -1575 2364 -1541
rect 2398 -1575 2414 -1541
rect 2348 -1609 2414 -1575
rect 2348 -1643 2364 -1609
rect 2398 -1643 2414 -1609
rect 2348 -1677 2414 -1643
rect 2348 -1711 2364 -1677
rect 2398 -1711 2414 -1677
rect 2348 -1719 2414 -1711
rect 2506 -1541 2559 -1525
rect 2506 -1575 2525 -1541
rect 2506 -1609 2559 -1575
rect 2506 -1643 2525 -1609
rect 2506 -1677 2559 -1643
rect 2506 -1711 2525 -1677
rect 2506 -1753 2559 -1711
rect 2593 -1541 2914 -1525
rect 2593 -1575 2609 -1541
rect 2643 -1559 2777 -1541
rect 2643 -1575 2659 -1559
rect 2593 -1609 2659 -1575
rect 2761 -1575 2777 -1559
rect 2811 -1563 2914 -1541
rect 3207 -1555 3265 -1520
rect 2811 -1575 2827 -1563
rect 2593 -1643 2609 -1609
rect 2643 -1643 2659 -1609
rect 2593 -1677 2659 -1643
rect 2593 -1711 2609 -1677
rect 2643 -1711 2659 -1677
rect 2593 -1719 2659 -1711
rect 2693 -1609 2727 -1593
rect 2693 -1677 2727 -1643
rect 2693 -1753 2727 -1711
rect 2761 -1609 2827 -1575
rect 2761 -1643 2777 -1609
rect 2811 -1643 2827 -1609
rect 2761 -1677 2827 -1643
rect 3207 -1589 3219 -1555
rect 3253 -1589 3265 -1555
rect 3207 -1648 3265 -1589
rect 2761 -1711 2777 -1677
rect 2811 -1711 2827 -1677
rect 2761 -1719 2827 -1711
rect 2861 -1677 2903 -1661
rect 2895 -1711 2903 -1677
rect 2861 -1753 2903 -1711
rect 3207 -1682 3219 -1648
rect 3253 -1682 3265 -1648
rect 3207 -1753 3265 -1682
rect -2584 -1787 -2555 -1753
rect -2521 -1787 -2492 -1753
rect -2242 -1787 -2213 -1753
rect -2179 -1787 -2121 -1753
rect -2087 -1787 -2029 -1753
rect -1995 -1787 -1937 -1753
rect -1903 -1787 -1845 -1753
rect -1811 -1787 -1753 -1753
rect -1719 -1787 -1661 -1753
rect -1627 -1787 -1569 -1753
rect -1535 -1787 -1477 -1753
rect -1443 -1787 -1385 -1753
rect -1351 -1787 -1293 -1753
rect -1259 -1787 -1201 -1753
rect -1167 -1787 -1109 -1753
rect -1075 -1787 -1017 -1753
rect -983 -1787 -925 -1753
rect -891 -1787 -833 -1753
rect -799 -1787 -741 -1753
rect -707 -1787 -649 -1753
rect -615 -1787 -557 -1753
rect -523 -1787 -465 -1753
rect -431 -1787 -373 -1753
rect -339 -1787 -281 -1753
rect -247 -1787 -189 -1753
rect -155 -1787 -97 -1753
rect -63 -1787 -5 -1753
rect 29 -1787 87 -1753
rect 121 -1787 179 -1753
rect 213 -1787 242 -1753
rect 456 -1787 485 -1753
rect 519 -1787 577 -1753
rect 611 -1787 669 -1753
rect 703 -1787 761 -1753
rect 795 -1787 853 -1753
rect 887 -1787 945 -1753
rect 979 -1787 1037 -1753
rect 1071 -1787 1129 -1753
rect 1163 -1787 1221 -1753
rect 1255 -1787 1313 -1753
rect 1347 -1787 1405 -1753
rect 1439 -1787 1497 -1753
rect 1531 -1787 1589 -1753
rect 1623 -1787 1681 -1753
rect 1715 -1787 1773 -1753
rect 1807 -1787 1865 -1753
rect 1899 -1787 1957 -1753
rect 1991 -1787 2049 -1753
rect 2083 -1787 2141 -1753
rect 2175 -1787 2233 -1753
rect 2267 -1787 2325 -1753
rect 2359 -1787 2417 -1753
rect 2451 -1787 2509 -1753
rect 2543 -1787 2601 -1753
rect 2635 -1787 2693 -1753
rect 2727 -1787 2785 -1753
rect 2819 -1787 2877 -1753
rect 2911 -1787 2940 -1753
rect 3190 -1787 3219 -1753
rect 3253 -1787 3282 -1753
rect -2567 -1858 -2509 -1787
rect -2567 -1892 -2555 -1858
rect -2521 -1892 -2509 -1858
rect -2567 -1951 -2509 -1892
rect -2567 -1985 -2555 -1951
rect -2521 -1985 -2509 -1951
rect -2207 -1837 -2173 -1821
rect -2207 -1905 -2173 -1871
rect -2139 -1853 -2073 -1787
rect -2139 -1887 -2123 -1853
rect -2089 -1887 -2073 -1853
rect -2039 -1837 -2002 -1821
rect -2005 -1871 -2002 -1837
rect -2039 -1905 -2002 -1871
rect -1954 -1829 -1901 -1787
rect -1954 -1863 -1935 -1829
rect -1954 -1879 -1901 -1863
rect -1867 -1837 -1817 -1821
rect -1867 -1871 -1851 -1837
rect -1520 -1829 -1486 -1787
rect -2173 -1923 -2074 -1921
rect -2173 -1939 -2116 -1923
rect -2207 -1955 -2116 -1939
rect -2567 -2020 -2509 -1985
rect -2120 -1957 -2116 -1955
rect -2082 -1957 -2074 -1923
rect -2224 -1998 -2154 -1989
rect -2224 -2046 -2218 -1998
rect -2170 -2046 -2154 -1998
rect -2224 -2065 -2154 -2046
rect -2224 -2099 -2210 -2065
rect -2176 -2099 -2154 -2065
rect -2224 -2119 -2154 -2099
rect -2120 -2050 -2074 -1957
rect -2120 -2084 -2108 -2050
rect -2567 -2169 -2509 -2152
rect -2120 -2153 -2074 -2084
rect -2567 -2203 -2555 -2169
rect -2521 -2203 -2509 -2169
rect -2567 -2297 -2509 -2203
rect -2207 -2187 -2074 -2153
rect -2005 -1939 -2002 -1905
rect -1867 -1906 -1817 -1871
rect -1775 -1876 -1759 -1842
rect -1725 -1876 -1554 -1842
rect -2039 -1991 -2002 -1939
rect -1878 -1932 -1817 -1906
rect -1728 -1923 -1622 -1910
rect -2039 -2025 -2037 -1991
rect -2003 -2025 -2002 -1991
rect -2207 -2195 -2173 -2187
rect -2039 -2195 -2002 -2025
rect -1968 -1997 -1912 -1981
rect -1968 -2031 -1946 -1997
rect -1968 -2088 -1912 -2031
rect -1968 -2136 -1962 -2088
rect -1914 -2136 -1912 -2088
rect -1968 -2171 -1912 -2136
rect -1878 -2153 -1844 -1932
rect -1728 -1957 -1696 -1923
rect -1662 -1949 -1622 -1923
rect -1810 -1991 -1762 -1970
rect -1810 -2025 -1799 -1991
rect -1765 -2025 -1762 -1991
rect -1810 -2027 -1762 -2025
rect -1810 -2061 -1803 -2027
rect -1769 -2061 -1762 -2027
rect -1810 -2089 -1762 -2061
rect -1728 -2123 -1694 -1957
rect -1660 -1983 -1622 -1949
rect -1588 -1999 -1554 -1876
rect -1520 -1897 -1486 -1863
rect -1520 -1947 -1486 -1931
rect -1452 -1837 -1402 -1821
rect -1452 -1871 -1436 -1837
rect -1144 -1837 -1081 -1787
rect -1452 -1887 -1402 -1871
rect -1357 -1881 -1341 -1847
rect -1307 -1881 -1180 -1847
rect -1588 -2015 -1486 -1999
rect -1588 -2017 -1520 -2015
rect -1878 -2179 -1833 -2153
rect -1799 -2157 -1783 -2123
rect -1749 -2157 -1694 -2123
rect -1799 -2167 -1694 -2157
rect -1660 -2049 -1520 -2017
rect -1660 -2051 -1486 -2049
rect -2207 -2245 -2173 -2229
rect -2139 -2255 -2123 -2221
rect -2089 -2255 -2073 -2221
rect -2005 -2229 -2002 -2195
rect -2039 -2245 -2002 -2229
rect -1951 -2221 -1901 -2205
rect -2139 -2297 -2073 -2255
rect -1951 -2255 -1935 -2221
rect -1867 -2207 -1833 -2179
rect -1660 -2207 -1626 -2051
rect -1520 -2065 -1486 -2051
rect -1584 -2101 -1544 -2095
rect -1452 -2101 -1418 -1887
rect -1384 -1923 -1346 -1921
rect -1384 -1957 -1382 -1923
rect -1348 -1957 -1346 -1923
rect -1384 -2015 -1346 -1957
rect -1350 -2049 -1346 -2015
rect -1384 -2065 -1346 -2049
rect -1312 -1949 -1248 -1915
rect -1312 -1983 -1282 -1949
rect -1312 -1991 -1248 -1983
rect -1312 -2025 -1295 -1991
rect -1261 -2025 -1248 -1991
rect -1584 -2111 -1418 -2101
rect -1312 -2107 -1248 -2025
rect -1550 -2145 -1418 -2111
rect -1584 -2161 -1418 -2145
rect -1867 -2241 -1850 -2207
rect -1816 -2241 -1800 -2207
rect -1761 -2241 -1739 -2207
rect -1705 -2241 -1626 -2207
rect -1562 -2213 -1488 -2197
rect -1951 -2297 -1901 -2255
rect -1562 -2247 -1540 -2213
rect -1506 -2247 -1488 -2213
rect -1452 -2207 -1418 -2161
rect -1341 -2123 -1248 -2107
rect -1307 -2157 -1248 -2123
rect -1341 -2173 -1248 -2157
rect -1214 -2049 -1180 -1881
rect -1144 -1871 -1142 -1837
rect -1108 -1871 -1081 -1837
rect -1144 -1887 -1081 -1871
rect -1034 -1829 -966 -1821
rect -1034 -1863 -1018 -1829
rect -984 -1863 -966 -1829
rect -1034 -1900 -966 -1863
rect -1034 -1933 -1018 -1900
rect -1146 -1934 -1018 -1933
rect -984 -1934 -966 -1900
rect -1146 -1949 -966 -1934
rect -1112 -1971 -966 -1949
rect -1112 -1983 -1018 -1971
rect -1146 -2005 -1018 -1983
rect -984 -2005 -966 -1971
rect -932 -1859 -898 -1787
rect -760 -1829 -694 -1825
rect -932 -1939 -898 -1893
rect -932 -1989 -898 -1973
rect -864 -1835 -798 -1830
rect -864 -1869 -848 -1835
rect -814 -1869 -798 -1835
rect -864 -1903 -798 -1869
rect -864 -1937 -848 -1903
rect -814 -1937 -798 -1903
rect -864 -1971 -798 -1937
rect -760 -1863 -744 -1829
rect -710 -1863 -694 -1829
rect -760 -1897 -694 -1863
rect -760 -1931 -744 -1897
rect -710 -1931 -694 -1897
rect -760 -1971 -694 -1931
rect -1146 -2008 -966 -2005
rect -1004 -2049 -966 -2008
rect -864 -2005 -848 -1971
rect -814 -1999 -798 -1971
rect -814 -2005 -782 -1999
rect -864 -2015 -782 -2005
rect -829 -2025 -782 -2015
rect -1214 -2065 -1038 -2049
rect -1214 -2099 -1072 -2065
rect -1214 -2115 -1038 -2099
rect -1004 -2065 -854 -2049
rect -1004 -2099 -888 -2065
rect -1004 -2115 -854 -2099
rect -1214 -2207 -1180 -2115
rect -1004 -2149 -964 -2115
rect -820 -2141 -782 -2025
rect -831 -2149 -782 -2141
rect -1030 -2152 -964 -2149
rect -1030 -2186 -1014 -2152
rect -980 -2186 -964 -2152
rect -862 -2150 -782 -2149
rect -862 -2168 -846 -2150
rect -812 -2166 -782 -2150
rect -748 -2049 -694 -1971
rect -656 -1829 -613 -1787
rect -656 -1863 -647 -1829
rect -656 -1897 -613 -1863
rect -656 -1931 -647 -1897
rect -656 -1965 -613 -1931
rect -656 -1999 -647 -1965
rect -656 -2015 -613 -1999
rect -579 -1829 -512 -1821
rect -579 -1863 -563 -1829
rect -529 -1863 -512 -1829
rect -579 -1900 -512 -1863
rect -579 -1934 -563 -1900
rect -529 -1934 -512 -1900
rect -579 -1971 -512 -1934
rect -579 -2005 -563 -1971
rect -529 -2005 -512 -1971
rect -579 -2018 -512 -2005
rect -426 -1829 -384 -1787
rect -426 -1863 -418 -1829
rect -426 -1897 -384 -1863
rect -426 -1931 -418 -1897
rect -426 -1965 -384 -1931
rect -426 -1999 -418 -1965
rect -426 -2015 -384 -1999
rect -350 -1829 -284 -1821
rect -350 -1863 -334 -1829
rect -300 -1863 -284 -1829
rect -350 -1897 -284 -1863
rect -350 -1931 -334 -1897
rect -300 -1931 -284 -1897
rect -350 -1965 -284 -1931
rect -350 -1999 -334 -1965
rect -300 -1999 -284 -1965
rect -350 -2017 -284 -1999
rect -192 -1829 -139 -1787
rect -192 -1863 -173 -1829
rect -192 -1897 -139 -1863
rect -192 -1931 -173 -1897
rect -192 -1965 -139 -1931
rect -192 -1999 -173 -1965
rect -192 -2015 -139 -1999
rect -105 -1829 -39 -1821
rect -105 -1863 -89 -1829
rect -55 -1863 -39 -1829
rect -105 -1897 -39 -1863
rect -105 -1931 -89 -1897
rect -55 -1931 -39 -1897
rect -105 -1965 -39 -1931
rect -5 -1829 29 -1787
rect -5 -1897 29 -1863
rect -5 -1947 29 -1931
rect 63 -1829 129 -1821
rect 63 -1863 79 -1829
rect 113 -1863 129 -1829
rect 63 -1897 129 -1863
rect 163 -1829 205 -1787
rect 197 -1863 205 -1829
rect 163 -1879 205 -1863
rect 491 -1837 525 -1821
rect 63 -1931 79 -1897
rect 113 -1931 129 -1897
rect -105 -1999 -89 -1965
rect -55 -1981 -39 -1965
rect 63 -1965 129 -1931
rect 491 -1905 525 -1871
rect 559 -1853 625 -1787
rect 559 -1887 575 -1853
rect 609 -1887 625 -1853
rect 659 -1837 696 -1821
rect 693 -1871 696 -1837
rect 659 -1905 696 -1871
rect 744 -1829 797 -1787
rect 744 -1863 763 -1829
rect 744 -1879 797 -1863
rect 831 -1837 881 -1821
rect 831 -1871 847 -1837
rect 1178 -1829 1212 -1787
rect 525 -1923 624 -1921
rect 525 -1939 582 -1923
rect 491 -1955 582 -1939
rect 63 -1981 79 -1965
rect -55 -1999 79 -1981
rect 113 -1977 129 -1965
rect 578 -1957 582 -1955
rect 616 -1957 624 -1923
rect 113 -1999 216 -1977
rect -105 -2015 216 -1999
rect -748 -2065 -593 -2049
rect -748 -2099 -627 -2065
rect -748 -2115 -593 -2099
rect -559 -2050 -512 -2018
rect -330 -2050 -284 -2017
rect -197 -2050 129 -2049
rect -559 -2098 -552 -2050
rect -388 -2065 -364 -2051
rect -812 -2168 -796 -2166
rect -1452 -2241 -1421 -2207
rect -1387 -2241 -1371 -2207
rect -1337 -2241 -1318 -2207
rect -1284 -2241 -1180 -2207
rect -1125 -2207 -1083 -2191
rect -1125 -2241 -1120 -2207
rect -1086 -2241 -1083 -2207
rect -1562 -2297 -1488 -2247
rect -1125 -2297 -1083 -2241
rect -1030 -2220 -964 -2186
rect -1030 -2254 -1014 -2220
rect -980 -2254 -964 -2220
rect -930 -2191 -896 -2175
rect -930 -2297 -896 -2225
rect -862 -2216 -858 -2168
rect -810 -2216 -796 -2168
rect -748 -2191 -708 -2115
rect -559 -2132 -512 -2098
rect -430 -2099 -414 -2098
rect -380 -2099 -364 -2065
rect -330 -2098 -324 -2050
rect -197 -2098 -192 -2050
rect -144 -2065 -82 -2050
rect -34 -2065 34 -2050
rect 82 -2065 129 -2050
rect -144 -2098 -89 -2065
rect -34 -2098 -5 -2065
rect -862 -2218 -796 -2216
rect -862 -2252 -846 -2218
rect -812 -2252 -796 -2218
rect -758 -2195 -708 -2191
rect -758 -2229 -742 -2195
rect -563 -2183 -512 -2132
rect -758 -2245 -708 -2229
rect -661 -2221 -597 -2205
rect -862 -2253 -796 -2252
rect -661 -2255 -647 -2221
rect -613 -2255 -597 -2221
rect -661 -2297 -597 -2255
rect -529 -2217 -512 -2183
rect -563 -2263 -512 -2217
rect -430 -2149 -384 -2133
rect -330 -2137 -284 -2098
rect -197 -2099 -181 -2098
rect -147 -2099 -89 -2098
rect -55 -2099 -5 -2098
rect 29 -2098 34 -2065
rect 29 -2099 79 -2098
rect 113 -2099 129 -2065
rect 163 -2052 216 -2015
rect 163 -2100 166 -2052
rect 214 -2100 216 -2052
rect 163 -2133 216 -2100
rect 474 -2040 544 -1989
rect 474 -2088 480 -2040
rect 528 -2088 544 -2040
rect 474 -2099 488 -2088
rect 522 -2099 544 -2088
rect 474 -2119 544 -2099
rect 578 -2050 624 -1957
rect 578 -2084 590 -2050
rect -430 -2183 -418 -2149
rect -430 -2217 -384 -2183
rect -430 -2251 -418 -2217
rect -430 -2297 -384 -2251
rect -350 -2149 -284 -2137
rect -350 -2183 -334 -2149
rect -300 -2183 -284 -2149
rect -350 -2217 -284 -2183
rect -105 -2169 216 -2133
rect 578 -2153 624 -2084
rect -350 -2251 -334 -2217
rect -300 -2251 -284 -2217
rect -350 -2263 -284 -2251
rect -192 -2221 -139 -2205
rect -192 -2255 -173 -2221
rect -192 -2297 -139 -2255
rect -105 -2213 -39 -2169
rect -105 -2247 -89 -2213
rect -55 -2247 -39 -2213
rect -105 -2263 -39 -2247
rect -5 -2221 29 -2205
rect -5 -2297 29 -2255
rect 63 -2213 129 -2169
rect 491 -2187 624 -2153
rect 693 -1939 696 -1905
rect 831 -1906 881 -1871
rect 923 -1876 939 -1842
rect 973 -1876 1144 -1842
rect 659 -1991 696 -1939
rect 820 -1932 881 -1906
rect 970 -1923 1076 -1910
rect 659 -2025 661 -1991
rect 695 -2025 696 -1991
rect 491 -2195 525 -2187
rect 63 -2247 79 -2213
rect 113 -2247 129 -2213
rect 63 -2263 129 -2247
rect 163 -2220 213 -2204
rect 197 -2254 213 -2220
rect 659 -2195 696 -2025
rect 730 -1997 786 -1981
rect 730 -2031 752 -1997
rect 730 -2088 786 -2031
rect 730 -2136 736 -2088
rect 784 -2136 786 -2088
rect 730 -2171 786 -2136
rect 820 -2153 854 -1932
rect 970 -1957 1002 -1923
rect 1036 -1949 1076 -1923
rect 888 -1991 936 -1970
rect 888 -2025 899 -1991
rect 933 -2025 936 -1991
rect 888 -2027 936 -2025
rect 888 -2061 895 -2027
rect 929 -2061 936 -2027
rect 888 -2089 936 -2061
rect 970 -2123 1004 -1957
rect 1038 -1983 1076 -1949
rect 1110 -1999 1144 -1876
rect 1178 -1897 1212 -1863
rect 1178 -1947 1212 -1931
rect 1246 -1837 1296 -1821
rect 1246 -1871 1262 -1837
rect 1554 -1837 1617 -1787
rect 1246 -1887 1296 -1871
rect 1341 -1881 1357 -1847
rect 1391 -1881 1518 -1847
rect 1110 -2015 1212 -1999
rect 1110 -2017 1178 -2015
rect 820 -2179 865 -2153
rect 899 -2157 915 -2123
rect 949 -2157 1004 -2123
rect 899 -2167 1004 -2157
rect 1038 -2049 1178 -2017
rect 1038 -2051 1212 -2049
rect 491 -2245 525 -2229
rect 163 -2297 213 -2254
rect 559 -2255 575 -2221
rect 609 -2255 625 -2221
rect 693 -2229 696 -2195
rect 659 -2245 696 -2229
rect 747 -2221 797 -2205
rect 559 -2297 625 -2255
rect 747 -2255 763 -2221
rect 831 -2207 865 -2179
rect 1038 -2207 1072 -2051
rect 1178 -2065 1212 -2051
rect 1114 -2101 1154 -2095
rect 1246 -2101 1280 -1887
rect 1314 -1923 1352 -1921
rect 1314 -1957 1316 -1923
rect 1350 -1957 1352 -1923
rect 1314 -2015 1352 -1957
rect 1348 -2049 1352 -2015
rect 1314 -2065 1352 -2049
rect 1386 -1949 1450 -1915
rect 1386 -1983 1416 -1949
rect 1386 -1991 1450 -1983
rect 1386 -2025 1403 -1991
rect 1437 -2025 1450 -1991
rect 1114 -2111 1280 -2101
rect 1386 -2107 1450 -2025
rect 1148 -2145 1280 -2111
rect 1114 -2161 1280 -2145
rect 831 -2241 848 -2207
rect 882 -2241 898 -2207
rect 937 -2241 959 -2207
rect 993 -2241 1072 -2207
rect 1136 -2213 1210 -2197
rect 747 -2297 797 -2255
rect 1136 -2247 1158 -2213
rect 1192 -2247 1210 -2213
rect 1246 -2207 1280 -2161
rect 1357 -2123 1450 -2107
rect 1391 -2157 1450 -2123
rect 1357 -2173 1450 -2157
rect 1484 -2049 1518 -1881
rect 1554 -1871 1556 -1837
rect 1590 -1871 1617 -1837
rect 1554 -1887 1617 -1871
rect 1664 -1829 1732 -1821
rect 1664 -1863 1680 -1829
rect 1714 -1863 1732 -1829
rect 1664 -1900 1732 -1863
rect 1664 -1933 1680 -1900
rect 1552 -1934 1680 -1933
rect 1714 -1934 1732 -1900
rect 1552 -1949 1732 -1934
rect 1586 -1971 1732 -1949
rect 1586 -1983 1680 -1971
rect 1552 -2005 1680 -1983
rect 1714 -2005 1732 -1971
rect 1766 -1859 1800 -1787
rect 1938 -1829 2004 -1825
rect 1766 -1939 1800 -1893
rect 1766 -1989 1800 -1973
rect 1834 -1835 1900 -1830
rect 1834 -1866 1850 -1835
rect 1884 -1866 1900 -1835
rect 1834 -1914 1840 -1866
rect 1888 -1914 1900 -1866
rect 1834 -1937 1850 -1914
rect 1884 -1937 1900 -1914
rect 1834 -1971 1900 -1937
rect 1938 -1863 1954 -1829
rect 1988 -1863 2004 -1829
rect 1938 -1897 2004 -1863
rect 1938 -1931 1954 -1897
rect 1988 -1931 2004 -1897
rect 1938 -1971 2004 -1931
rect 1552 -2008 1732 -2005
rect 1694 -2049 1732 -2008
rect 1834 -2005 1850 -1971
rect 1884 -1999 1900 -1971
rect 1884 -2005 1916 -1999
rect 1834 -2015 1916 -2005
rect 1869 -2025 1916 -2015
rect 1484 -2065 1660 -2049
rect 1484 -2099 1626 -2065
rect 1484 -2115 1660 -2099
rect 1694 -2065 1844 -2049
rect 1694 -2099 1810 -2065
rect 1694 -2115 1844 -2099
rect 1484 -2207 1518 -2115
rect 1694 -2149 1734 -2115
rect 1878 -2141 1916 -2025
rect 1867 -2149 1916 -2141
rect 1668 -2152 1734 -2149
rect 1668 -2186 1684 -2152
rect 1718 -2186 1734 -2152
rect 1836 -2150 1916 -2149
rect 1246 -2241 1277 -2207
rect 1311 -2241 1327 -2207
rect 1361 -2241 1380 -2207
rect 1414 -2241 1518 -2207
rect 1573 -2207 1615 -2191
rect 1573 -2241 1578 -2207
rect 1612 -2241 1615 -2207
rect 1136 -2297 1210 -2247
rect 1573 -2297 1615 -2241
rect 1668 -2220 1734 -2186
rect 1668 -2254 1684 -2220
rect 1718 -2254 1734 -2220
rect 1768 -2191 1802 -2175
rect 1768 -2297 1802 -2225
rect 1836 -2184 1852 -2150
rect 1886 -2166 1916 -2150
rect 1950 -2049 2004 -1971
rect 2042 -1829 2085 -1787
rect 2042 -1863 2051 -1829
rect 2042 -1897 2085 -1863
rect 2042 -1931 2051 -1897
rect 2042 -1965 2085 -1931
rect 2042 -1999 2051 -1965
rect 2042 -2015 2085 -1999
rect 2119 -1829 2186 -1821
rect 2119 -1863 2135 -1829
rect 2169 -1863 2186 -1829
rect 2119 -1900 2186 -1863
rect 2119 -1934 2135 -1900
rect 2169 -1934 2186 -1900
rect 2119 -1971 2186 -1934
rect 2119 -2005 2135 -1971
rect 2169 -2005 2186 -1971
rect 2119 -2018 2186 -2005
rect 2272 -1829 2314 -1787
rect 2272 -1863 2280 -1829
rect 2272 -1897 2314 -1863
rect 2272 -1931 2280 -1897
rect 2272 -1965 2314 -1931
rect 2272 -1999 2280 -1965
rect 2272 -2015 2314 -1999
rect 2348 -1829 2414 -1821
rect 2348 -1863 2364 -1829
rect 2398 -1863 2414 -1829
rect 2348 -1897 2414 -1863
rect 2348 -1931 2364 -1897
rect 2398 -1931 2414 -1897
rect 2348 -1965 2414 -1931
rect 2348 -1999 2364 -1965
rect 2398 -1999 2414 -1965
rect 2348 -2017 2414 -1999
rect 2506 -1829 2559 -1787
rect 2506 -1863 2525 -1829
rect 2506 -1897 2559 -1863
rect 2506 -1931 2525 -1897
rect 2506 -1965 2559 -1931
rect 2506 -1999 2525 -1965
rect 2506 -2015 2559 -1999
rect 2593 -1829 2659 -1821
rect 2593 -1863 2609 -1829
rect 2643 -1863 2659 -1829
rect 2593 -1897 2659 -1863
rect 2593 -1931 2609 -1897
rect 2643 -1931 2659 -1897
rect 2593 -1965 2659 -1931
rect 2693 -1829 2727 -1787
rect 2693 -1897 2727 -1863
rect 2693 -1947 2727 -1931
rect 2761 -1829 2827 -1821
rect 2761 -1863 2777 -1829
rect 2811 -1863 2827 -1829
rect 2761 -1897 2827 -1863
rect 2861 -1829 2903 -1787
rect 2895 -1863 2903 -1829
rect 2861 -1879 2903 -1863
rect 3207 -1858 3265 -1787
rect 2761 -1931 2777 -1897
rect 2811 -1931 2827 -1897
rect 2593 -1999 2609 -1965
rect 2643 -1981 2659 -1965
rect 2761 -1965 2827 -1931
rect 2761 -1981 2777 -1965
rect 2643 -1999 2777 -1981
rect 2811 -1977 2827 -1965
rect 3207 -1892 3219 -1858
rect 3253 -1892 3265 -1858
rect 3207 -1951 3265 -1892
rect 2811 -1999 2914 -1977
rect 2593 -2015 2914 -1999
rect 1950 -2065 2105 -2049
rect 1950 -2099 2071 -2065
rect 1950 -2115 2105 -2099
rect 2139 -2050 2186 -2018
rect 2368 -2050 2414 -2017
rect 2501 -2050 2827 -2049
rect 2139 -2098 2146 -2050
rect 2310 -2065 2334 -2051
rect 1886 -2184 1902 -2166
rect 1836 -2218 1902 -2184
rect 1950 -2191 1990 -2115
rect 2139 -2132 2186 -2098
rect 2268 -2099 2284 -2098
rect 2318 -2099 2334 -2065
rect 2368 -2098 2374 -2050
rect 2501 -2098 2506 -2050
rect 2554 -2065 2616 -2050
rect 2664 -2065 2732 -2050
rect 2780 -2065 2827 -2050
rect 2554 -2098 2609 -2065
rect 2664 -2098 2693 -2065
rect 1836 -2252 1852 -2218
rect 1886 -2252 1902 -2218
rect 1940 -2195 1990 -2191
rect 1940 -2229 1956 -2195
rect 2135 -2183 2186 -2132
rect 1940 -2245 1990 -2229
rect 2037 -2221 2101 -2205
rect 1836 -2253 1902 -2252
rect 2037 -2255 2051 -2221
rect 2085 -2255 2101 -2221
rect 2037 -2297 2101 -2255
rect 2169 -2217 2186 -2183
rect 2135 -2263 2186 -2217
rect 2268 -2149 2314 -2133
rect 2368 -2137 2414 -2098
rect 2501 -2099 2517 -2098
rect 2551 -2099 2609 -2098
rect 2643 -2099 2693 -2098
rect 2727 -2098 2732 -2065
rect 2727 -2099 2777 -2098
rect 2811 -2099 2827 -2065
rect 2861 -2052 2914 -2015
rect 3207 -1985 3219 -1951
rect 3253 -1985 3265 -1951
rect 3207 -2020 3265 -1985
rect 2861 -2100 2868 -2052
rect 2861 -2133 2914 -2100
rect 2268 -2183 2280 -2149
rect 2268 -2217 2314 -2183
rect 2268 -2251 2280 -2217
rect 2268 -2297 2314 -2251
rect 2348 -2149 2414 -2137
rect 2348 -2183 2364 -2149
rect 2398 -2183 2414 -2149
rect 2348 -2217 2414 -2183
rect 2593 -2169 2914 -2133
rect 3207 -2169 3265 -2152
rect 2348 -2251 2364 -2217
rect 2398 -2251 2414 -2217
rect 2348 -2263 2414 -2251
rect 2506 -2221 2559 -2205
rect 2506 -2255 2525 -2221
rect 2506 -2297 2559 -2255
rect 2593 -2213 2659 -2169
rect 2593 -2247 2609 -2213
rect 2643 -2247 2659 -2213
rect 2593 -2263 2659 -2247
rect 2693 -2221 2727 -2205
rect 2693 -2297 2727 -2255
rect 2761 -2213 2827 -2169
rect 3207 -2203 3219 -2169
rect 3253 -2203 3265 -2169
rect 2761 -2247 2777 -2213
rect 2811 -2247 2827 -2213
rect 2761 -2263 2827 -2247
rect 2861 -2220 2911 -2204
rect 2895 -2254 2911 -2220
rect 2861 -2297 2911 -2254
rect 3207 -2297 3265 -2203
rect -2584 -2331 -2555 -2297
rect -2521 -2331 -2492 -2297
rect -2242 -2331 -2213 -2297
rect -2179 -2331 -2121 -2297
rect -2087 -2331 -2029 -2297
rect -1995 -2331 -1937 -2297
rect -1903 -2331 -1845 -2297
rect -1811 -2331 -1753 -2297
rect -1719 -2331 -1661 -2297
rect -1627 -2331 -1569 -2297
rect -1535 -2331 -1477 -2297
rect -1443 -2331 -1385 -2297
rect -1351 -2331 -1293 -2297
rect -1259 -2331 -1201 -2297
rect -1167 -2331 -1109 -2297
rect -1075 -2331 -1017 -2297
rect -983 -2331 -925 -2297
rect -891 -2331 -833 -2297
rect -799 -2331 -741 -2297
rect -707 -2331 -649 -2297
rect -615 -2331 -557 -2297
rect -523 -2331 -465 -2297
rect -431 -2331 -373 -2297
rect -339 -2331 -281 -2297
rect -247 -2331 -189 -2297
rect -155 -2331 -97 -2297
rect -63 -2331 -5 -2297
rect 29 -2331 87 -2297
rect 121 -2331 179 -2297
rect 213 -2331 242 -2297
rect 456 -2331 485 -2297
rect 519 -2331 577 -2297
rect 611 -2331 669 -2297
rect 703 -2331 761 -2297
rect 795 -2331 853 -2297
rect 887 -2331 945 -2297
rect 979 -2331 1037 -2297
rect 1071 -2331 1129 -2297
rect 1163 -2331 1221 -2297
rect 1255 -2331 1313 -2297
rect 1347 -2331 1405 -2297
rect 1439 -2331 1497 -2297
rect 1531 -2331 1589 -2297
rect 1623 -2331 1681 -2297
rect 1715 -2331 1773 -2297
rect 1807 -2331 1865 -2297
rect 1899 -2331 1957 -2297
rect 1991 -2331 2049 -2297
rect 2083 -2331 2141 -2297
rect 2175 -2331 2233 -2297
rect 2267 -2331 2325 -2297
rect 2359 -2331 2417 -2297
rect 2451 -2331 2509 -2297
rect 2543 -2331 2601 -2297
rect 2635 -2331 2693 -2297
rect 2727 -2331 2785 -2297
rect 2819 -2331 2877 -2297
rect 2911 -2331 2940 -2297
rect 3190 -2331 3219 -2297
rect 3253 -2331 3282 -2297
rect -2567 -2425 -2509 -2331
rect -2139 -2373 -2073 -2331
rect -2567 -2459 -2555 -2425
rect -2521 -2459 -2509 -2425
rect -2567 -2476 -2509 -2459
rect -2207 -2399 -2173 -2383
rect -2139 -2407 -2123 -2373
rect -2089 -2407 -2073 -2373
rect -1951 -2373 -1901 -2331
rect -2039 -2399 -2002 -2383
rect -2207 -2441 -2173 -2433
rect -2005 -2433 -2002 -2399
rect -1951 -2407 -1935 -2373
rect -1562 -2381 -1488 -2331
rect -1951 -2423 -1901 -2407
rect -1867 -2421 -1850 -2387
rect -1816 -2421 -1800 -2387
rect -1761 -2421 -1739 -2387
rect -1705 -2421 -1626 -2387
rect -2207 -2475 -2074 -2441
rect -2224 -2529 -2154 -2509
rect -2224 -2540 -2210 -2529
rect -2176 -2540 -2154 -2529
rect -2224 -2588 -2218 -2540
rect -2170 -2588 -2154 -2540
rect -2567 -2643 -2509 -2608
rect -2224 -2639 -2154 -2588
rect -2120 -2544 -2074 -2475
rect -2120 -2578 -2108 -2544
rect -2567 -2677 -2555 -2643
rect -2521 -2677 -2509 -2643
rect -2120 -2671 -2074 -2578
rect -2120 -2673 -2116 -2671
rect -2567 -2736 -2509 -2677
rect -2567 -2770 -2555 -2736
rect -2521 -2770 -2509 -2736
rect -2567 -2841 -2509 -2770
rect -2207 -2689 -2116 -2673
rect -2173 -2705 -2116 -2689
rect -2082 -2705 -2074 -2671
rect -2173 -2707 -2074 -2705
rect -2039 -2603 -2002 -2433
rect -1867 -2449 -1833 -2421
rect -2039 -2637 -2037 -2603
rect -2003 -2637 -2002 -2603
rect -2039 -2689 -2002 -2637
rect -1968 -2492 -1912 -2457
rect -1968 -2540 -1962 -2492
rect -1914 -2540 -1912 -2492
rect -1968 -2597 -1912 -2540
rect -1968 -2631 -1946 -2597
rect -1968 -2647 -1912 -2631
rect -1878 -2475 -1833 -2449
rect -1799 -2471 -1694 -2461
rect -2207 -2757 -2173 -2723
rect -2005 -2723 -2002 -2689
rect -1878 -2696 -1844 -2475
rect -1799 -2505 -1783 -2471
rect -1749 -2505 -1694 -2471
rect -1810 -2567 -1762 -2539
rect -1810 -2601 -1803 -2567
rect -1769 -2601 -1762 -2567
rect -1810 -2603 -1762 -2601
rect -1810 -2637 -1799 -2603
rect -1765 -2637 -1762 -2603
rect -1810 -2658 -1762 -2637
rect -1728 -2671 -1694 -2505
rect -1660 -2577 -1626 -2421
rect -1562 -2415 -1540 -2381
rect -1506 -2415 -1488 -2381
rect -1125 -2387 -1083 -2331
rect -1562 -2431 -1488 -2415
rect -1452 -2421 -1421 -2387
rect -1387 -2421 -1371 -2387
rect -1337 -2421 -1318 -2387
rect -1284 -2421 -1180 -2387
rect -1452 -2467 -1418 -2421
rect -1584 -2483 -1418 -2467
rect -1550 -2517 -1418 -2483
rect -1584 -2527 -1418 -2517
rect -1341 -2471 -1248 -2455
rect -1307 -2505 -1248 -2471
rect -1341 -2521 -1248 -2505
rect -1584 -2533 -1544 -2527
rect -1520 -2577 -1486 -2563
rect -1660 -2579 -1486 -2577
rect -1660 -2611 -1520 -2579
rect -1588 -2613 -1520 -2611
rect -1588 -2629 -1486 -2613
rect -1878 -2722 -1817 -2696
rect -1728 -2705 -1696 -2671
rect -1660 -2679 -1622 -2645
rect -1662 -2705 -1622 -2679
rect -1728 -2718 -1622 -2705
rect -2207 -2807 -2173 -2791
rect -2139 -2775 -2123 -2741
rect -2089 -2775 -2073 -2741
rect -2139 -2841 -2073 -2775
rect -2039 -2757 -2002 -2723
rect -2005 -2791 -2002 -2757
rect -2039 -2807 -2002 -2791
rect -1954 -2765 -1901 -2749
rect -1954 -2799 -1935 -2765
rect -1954 -2841 -1901 -2799
rect -1867 -2757 -1817 -2722
rect -1588 -2752 -1554 -2629
rect -1867 -2791 -1851 -2757
rect -1775 -2786 -1759 -2752
rect -1725 -2786 -1554 -2752
rect -1520 -2697 -1486 -2681
rect -1520 -2765 -1486 -2731
rect -1867 -2807 -1817 -2791
rect -1520 -2841 -1486 -2799
rect -1452 -2741 -1418 -2527
rect -1384 -2579 -1346 -2563
rect -1350 -2613 -1346 -2579
rect -1384 -2671 -1346 -2613
rect -1384 -2705 -1382 -2671
rect -1348 -2705 -1346 -2671
rect -1384 -2707 -1346 -2705
rect -1312 -2603 -1248 -2521
rect -1312 -2637 -1295 -2603
rect -1261 -2637 -1248 -2603
rect -1312 -2645 -1248 -2637
rect -1312 -2679 -1282 -2645
rect -1312 -2713 -1248 -2679
rect -1214 -2513 -1180 -2421
rect -1125 -2421 -1120 -2387
rect -1086 -2421 -1083 -2387
rect -1125 -2437 -1083 -2421
rect -1030 -2408 -1014 -2374
rect -980 -2408 -964 -2374
rect -1030 -2442 -964 -2408
rect -1030 -2476 -1014 -2442
rect -980 -2476 -964 -2442
rect -930 -2403 -896 -2331
rect -661 -2373 -597 -2331
rect -930 -2453 -896 -2437
rect -862 -2376 -796 -2375
rect -862 -2410 -846 -2376
rect -812 -2410 -796 -2376
rect -862 -2444 -796 -2410
rect -758 -2399 -708 -2383
rect -758 -2433 -742 -2399
rect -661 -2407 -647 -2373
rect -613 -2407 -597 -2373
rect -661 -2423 -597 -2407
rect -563 -2411 -512 -2365
rect -758 -2437 -708 -2433
rect -1030 -2479 -964 -2476
rect -862 -2478 -846 -2444
rect -812 -2462 -796 -2444
rect -812 -2478 -782 -2462
rect -862 -2479 -782 -2478
rect -1004 -2513 -964 -2479
rect -831 -2487 -782 -2479
rect -1214 -2529 -1038 -2513
rect -1214 -2563 -1072 -2529
rect -1214 -2579 -1038 -2563
rect -1004 -2529 -854 -2513
rect -1004 -2563 -888 -2529
rect -1004 -2579 -854 -2563
rect -1452 -2757 -1402 -2741
rect -1214 -2747 -1180 -2579
rect -1004 -2620 -966 -2579
rect -820 -2603 -782 -2487
rect -829 -2613 -782 -2603
rect -1146 -2623 -966 -2620
rect -1146 -2645 -1018 -2623
rect -1112 -2657 -1018 -2645
rect -984 -2657 -966 -2623
rect -864 -2623 -782 -2613
rect -1112 -2679 -966 -2657
rect -1146 -2694 -966 -2679
rect -1146 -2695 -1018 -2694
rect -1034 -2728 -1018 -2695
rect -984 -2728 -966 -2694
rect -1452 -2791 -1436 -2757
rect -1357 -2781 -1341 -2747
rect -1307 -2781 -1180 -2747
rect -1144 -2757 -1081 -2741
rect -1452 -2807 -1402 -2791
rect -1144 -2791 -1142 -2757
rect -1108 -2791 -1081 -2757
rect -1144 -2841 -1081 -2791
rect -1034 -2765 -966 -2728
rect -1034 -2799 -1018 -2765
rect -984 -2799 -966 -2765
rect -1034 -2807 -966 -2799
rect -932 -2655 -898 -2639
rect -932 -2735 -898 -2689
rect -932 -2841 -898 -2769
rect -864 -2657 -848 -2623
rect -814 -2629 -782 -2623
rect -748 -2513 -708 -2437
rect -529 -2445 -512 -2411
rect -563 -2496 -512 -2445
rect -430 -2377 -384 -2331
rect -430 -2411 -418 -2377
rect -430 -2445 -384 -2411
rect -430 -2479 -418 -2445
rect -430 -2495 -384 -2479
rect -350 -2377 -284 -2365
rect -350 -2411 -334 -2377
rect -300 -2411 -284 -2377
rect -350 -2445 -284 -2411
rect -192 -2373 -139 -2331
rect -192 -2407 -173 -2373
rect -192 -2423 -139 -2407
rect -105 -2381 -39 -2365
rect -105 -2415 -89 -2381
rect -55 -2415 -39 -2381
rect -350 -2479 -334 -2445
rect -300 -2479 -284 -2445
rect -350 -2491 -284 -2479
rect -748 -2529 -593 -2513
rect -748 -2563 -627 -2529
rect -748 -2579 -593 -2563
rect -559 -2530 -512 -2496
rect -430 -2530 -414 -2529
rect -559 -2578 -552 -2530
rect -380 -2563 -364 -2529
rect -388 -2577 -364 -2563
rect -330 -2530 -284 -2491
rect -105 -2459 -39 -2415
rect -5 -2373 29 -2331
rect -5 -2423 29 -2407
rect 63 -2381 129 -2365
rect 63 -2415 79 -2381
rect 113 -2415 129 -2381
rect 63 -2459 129 -2415
rect 163 -2374 213 -2331
rect 197 -2408 213 -2374
rect 559 -2373 625 -2331
rect 163 -2424 213 -2408
rect 491 -2399 525 -2383
rect 559 -2407 575 -2373
rect 609 -2407 625 -2373
rect 747 -2373 797 -2331
rect 659 -2399 696 -2383
rect 491 -2441 525 -2433
rect 693 -2433 696 -2399
rect 747 -2407 763 -2373
rect 1136 -2381 1210 -2331
rect 747 -2423 797 -2407
rect 831 -2421 848 -2387
rect 882 -2421 898 -2387
rect 937 -2421 959 -2387
rect 993 -2421 1072 -2387
rect -105 -2495 216 -2459
rect 491 -2475 624 -2441
rect 163 -2528 216 -2495
rect 474 -2522 544 -2509
rect -197 -2530 -181 -2529
rect -147 -2530 -89 -2529
rect -55 -2530 -5 -2529
rect -330 -2578 -324 -2530
rect -197 -2578 -192 -2530
rect -144 -2563 -89 -2530
rect -34 -2563 -5 -2530
rect 29 -2530 79 -2529
rect 29 -2563 34 -2530
rect 113 -2563 129 -2529
rect -144 -2578 -82 -2563
rect -34 -2578 34 -2563
rect 82 -2578 129 -2563
rect -814 -2657 -798 -2629
rect -748 -2657 -694 -2579
rect -559 -2610 -512 -2578
rect -864 -2691 -798 -2657
rect -864 -2712 -848 -2691
rect -814 -2712 -798 -2691
rect -864 -2760 -858 -2712
rect -810 -2760 -798 -2712
rect -864 -2793 -848 -2760
rect -814 -2793 -798 -2760
rect -864 -2798 -798 -2793
rect -760 -2697 -694 -2657
rect -760 -2731 -744 -2697
rect -710 -2731 -694 -2697
rect -760 -2765 -694 -2731
rect -760 -2799 -744 -2765
rect -710 -2799 -694 -2765
rect -760 -2803 -694 -2799
rect -656 -2629 -613 -2613
rect -656 -2663 -647 -2629
rect -656 -2697 -613 -2663
rect -656 -2731 -647 -2697
rect -656 -2765 -613 -2731
rect -656 -2799 -647 -2765
rect -656 -2841 -613 -2799
rect -579 -2623 -512 -2610
rect -330 -2611 -284 -2578
rect -197 -2579 129 -2578
rect 163 -2576 166 -2528
rect 474 -2570 488 -2522
rect 536 -2570 544 -2522
rect -579 -2657 -563 -2623
rect -529 -2657 -512 -2623
rect -579 -2694 -512 -2657
rect -579 -2728 -563 -2694
rect -529 -2728 -512 -2694
rect -579 -2765 -512 -2728
rect -579 -2799 -563 -2765
rect -529 -2799 -512 -2765
rect -579 -2807 -512 -2799
rect -426 -2629 -384 -2613
rect -426 -2663 -418 -2629
rect -426 -2697 -384 -2663
rect -426 -2731 -418 -2697
rect -426 -2765 -384 -2731
rect -426 -2799 -418 -2765
rect -426 -2841 -384 -2799
rect -350 -2629 -284 -2611
rect 163 -2613 216 -2576
rect -350 -2663 -334 -2629
rect -300 -2663 -284 -2629
rect -350 -2697 -284 -2663
rect -350 -2731 -334 -2697
rect -300 -2731 -284 -2697
rect -350 -2765 -284 -2731
rect -350 -2799 -334 -2765
rect -300 -2799 -284 -2765
rect -350 -2807 -284 -2799
rect -192 -2629 -139 -2613
rect -192 -2663 -173 -2629
rect -192 -2697 -139 -2663
rect -192 -2731 -173 -2697
rect -192 -2765 -139 -2731
rect -192 -2799 -173 -2765
rect -192 -2841 -139 -2799
rect -105 -2629 216 -2613
rect -105 -2663 -89 -2629
rect -55 -2647 79 -2629
rect -55 -2663 -39 -2647
rect -105 -2697 -39 -2663
rect 63 -2663 79 -2647
rect 113 -2651 216 -2629
rect 474 -2639 544 -2570
rect 578 -2544 624 -2475
rect 578 -2578 590 -2544
rect 113 -2663 129 -2651
rect -105 -2731 -89 -2697
rect -55 -2731 -39 -2697
rect -105 -2765 -39 -2731
rect -105 -2799 -89 -2765
rect -55 -2799 -39 -2765
rect -105 -2807 -39 -2799
rect -5 -2697 29 -2681
rect -5 -2765 29 -2731
rect -5 -2841 29 -2799
rect 63 -2697 129 -2663
rect 578 -2671 624 -2578
rect 578 -2673 582 -2671
rect 63 -2731 79 -2697
rect 113 -2731 129 -2697
rect 63 -2765 129 -2731
rect 491 -2689 582 -2673
rect 525 -2705 582 -2689
rect 616 -2705 624 -2671
rect 525 -2707 624 -2705
rect 659 -2603 696 -2433
rect 831 -2449 865 -2421
rect 659 -2637 661 -2603
rect 695 -2637 696 -2603
rect 659 -2689 696 -2637
rect 730 -2492 786 -2457
rect 730 -2540 736 -2492
rect 784 -2540 786 -2492
rect 730 -2597 786 -2540
rect 730 -2631 752 -2597
rect 730 -2647 786 -2631
rect 820 -2475 865 -2449
rect 899 -2471 1004 -2461
rect 63 -2799 79 -2765
rect 113 -2799 129 -2765
rect 63 -2807 129 -2799
rect 163 -2765 205 -2749
rect 197 -2799 205 -2765
rect 163 -2841 205 -2799
rect 491 -2757 525 -2723
rect 693 -2723 696 -2689
rect 820 -2696 854 -2475
rect 899 -2505 915 -2471
rect 949 -2505 1004 -2471
rect 888 -2567 936 -2539
rect 888 -2601 895 -2567
rect 929 -2601 936 -2567
rect 888 -2603 936 -2601
rect 888 -2637 899 -2603
rect 933 -2637 936 -2603
rect 888 -2658 936 -2637
rect 970 -2671 1004 -2505
rect 1038 -2577 1072 -2421
rect 1136 -2415 1158 -2381
rect 1192 -2415 1210 -2381
rect 1573 -2387 1615 -2331
rect 1136 -2431 1210 -2415
rect 1246 -2421 1277 -2387
rect 1311 -2421 1327 -2387
rect 1361 -2421 1380 -2387
rect 1414 -2421 1518 -2387
rect 1246 -2467 1280 -2421
rect 1114 -2483 1280 -2467
rect 1148 -2517 1280 -2483
rect 1114 -2527 1280 -2517
rect 1357 -2471 1450 -2455
rect 1391 -2505 1450 -2471
rect 1357 -2521 1450 -2505
rect 1114 -2533 1154 -2527
rect 1178 -2577 1212 -2563
rect 1038 -2579 1212 -2577
rect 1038 -2611 1178 -2579
rect 1110 -2613 1178 -2611
rect 1110 -2629 1212 -2613
rect 820 -2722 881 -2696
rect 970 -2705 1002 -2671
rect 1038 -2679 1076 -2645
rect 1036 -2705 1076 -2679
rect 970 -2718 1076 -2705
rect 491 -2807 525 -2791
rect 559 -2775 575 -2741
rect 609 -2775 625 -2741
rect 559 -2841 625 -2775
rect 659 -2757 696 -2723
rect 693 -2791 696 -2757
rect 659 -2807 696 -2791
rect 744 -2765 797 -2749
rect 744 -2799 763 -2765
rect 744 -2841 797 -2799
rect 831 -2757 881 -2722
rect 1110 -2752 1144 -2629
rect 831 -2791 847 -2757
rect 923 -2786 939 -2752
rect 973 -2786 1144 -2752
rect 1178 -2697 1212 -2681
rect 1178 -2765 1212 -2731
rect 831 -2807 881 -2791
rect 1178 -2841 1212 -2799
rect 1246 -2741 1280 -2527
rect 1314 -2579 1352 -2563
rect 1348 -2613 1352 -2579
rect 1314 -2671 1352 -2613
rect 1314 -2705 1316 -2671
rect 1350 -2705 1352 -2671
rect 1314 -2707 1352 -2705
rect 1386 -2603 1450 -2521
rect 1386 -2637 1403 -2603
rect 1437 -2637 1450 -2603
rect 1386 -2645 1450 -2637
rect 1386 -2679 1416 -2645
rect 1386 -2713 1450 -2679
rect 1484 -2513 1518 -2421
rect 1573 -2421 1578 -2387
rect 1612 -2421 1615 -2387
rect 1573 -2437 1615 -2421
rect 1668 -2408 1684 -2374
rect 1718 -2408 1734 -2374
rect 1668 -2442 1734 -2408
rect 1668 -2476 1684 -2442
rect 1718 -2476 1734 -2442
rect 1768 -2403 1802 -2331
rect 2037 -2373 2101 -2331
rect 1768 -2453 1802 -2437
rect 1836 -2376 1902 -2375
rect 1836 -2410 1852 -2376
rect 1886 -2410 1902 -2376
rect 1836 -2412 1902 -2410
rect 1668 -2479 1734 -2476
rect 1836 -2460 1840 -2412
rect 1888 -2460 1902 -2412
rect 1940 -2399 1990 -2383
rect 1940 -2433 1956 -2399
rect 2037 -2407 2051 -2373
rect 2085 -2407 2101 -2373
rect 2037 -2423 2101 -2407
rect 2135 -2411 2186 -2365
rect 1940 -2437 1990 -2433
rect 1836 -2478 1852 -2460
rect 1886 -2462 1902 -2460
rect 1886 -2478 1916 -2462
rect 1836 -2479 1916 -2478
rect 1694 -2513 1734 -2479
rect 1867 -2487 1916 -2479
rect 1484 -2529 1660 -2513
rect 1484 -2563 1626 -2529
rect 1484 -2579 1660 -2563
rect 1694 -2529 1844 -2513
rect 1694 -2563 1810 -2529
rect 1694 -2579 1844 -2563
rect 1246 -2757 1296 -2741
rect 1484 -2747 1518 -2579
rect 1694 -2620 1732 -2579
rect 1878 -2603 1916 -2487
rect 1869 -2613 1916 -2603
rect 1552 -2623 1732 -2620
rect 1552 -2645 1680 -2623
rect 1586 -2657 1680 -2645
rect 1714 -2657 1732 -2623
rect 1834 -2623 1916 -2613
rect 1586 -2679 1732 -2657
rect 1552 -2694 1732 -2679
rect 1552 -2695 1680 -2694
rect 1664 -2728 1680 -2695
rect 1714 -2728 1732 -2694
rect 1246 -2791 1262 -2757
rect 1341 -2781 1357 -2747
rect 1391 -2781 1518 -2747
rect 1554 -2757 1617 -2741
rect 1246 -2807 1296 -2791
rect 1554 -2791 1556 -2757
rect 1590 -2791 1617 -2757
rect 1554 -2841 1617 -2791
rect 1664 -2765 1732 -2728
rect 1664 -2799 1680 -2765
rect 1714 -2799 1732 -2765
rect 1664 -2807 1732 -2799
rect 1766 -2655 1800 -2639
rect 1766 -2735 1800 -2689
rect 1766 -2841 1800 -2769
rect 1834 -2657 1850 -2623
rect 1884 -2629 1916 -2623
rect 1950 -2513 1990 -2437
rect 2169 -2445 2186 -2411
rect 2135 -2496 2186 -2445
rect 2268 -2377 2314 -2331
rect 2268 -2411 2280 -2377
rect 2268 -2445 2314 -2411
rect 2268 -2479 2280 -2445
rect 2268 -2495 2314 -2479
rect 2348 -2377 2414 -2365
rect 2348 -2411 2364 -2377
rect 2398 -2411 2414 -2377
rect 2348 -2445 2414 -2411
rect 2506 -2373 2559 -2331
rect 2506 -2407 2525 -2373
rect 2506 -2423 2559 -2407
rect 2593 -2381 2659 -2365
rect 2593 -2415 2609 -2381
rect 2643 -2415 2659 -2381
rect 2348 -2479 2364 -2445
rect 2398 -2479 2414 -2445
rect 2348 -2491 2414 -2479
rect 1950 -2529 2105 -2513
rect 1950 -2563 2071 -2529
rect 1950 -2579 2105 -2563
rect 2139 -2530 2186 -2496
rect 2268 -2530 2284 -2529
rect 2139 -2578 2146 -2530
rect 2318 -2563 2334 -2529
rect 2310 -2577 2334 -2563
rect 2368 -2530 2414 -2491
rect 2593 -2459 2659 -2415
rect 2693 -2373 2727 -2331
rect 2693 -2423 2727 -2407
rect 2761 -2381 2827 -2365
rect 2761 -2415 2777 -2381
rect 2811 -2415 2827 -2381
rect 2761 -2459 2827 -2415
rect 2861 -2374 2911 -2331
rect 2895 -2408 2911 -2374
rect 2861 -2424 2911 -2408
rect 3207 -2425 3265 -2331
rect 3207 -2459 3219 -2425
rect 3253 -2459 3265 -2425
rect 2593 -2495 2914 -2459
rect 3207 -2476 3265 -2459
rect 2861 -2528 2914 -2495
rect 2501 -2530 2517 -2529
rect 2551 -2530 2609 -2529
rect 2643 -2530 2693 -2529
rect 2368 -2578 2374 -2530
rect 2501 -2578 2506 -2530
rect 2554 -2563 2609 -2530
rect 2664 -2563 2693 -2530
rect 2727 -2530 2777 -2529
rect 2727 -2563 2732 -2530
rect 2811 -2563 2827 -2529
rect 2554 -2578 2616 -2563
rect 2664 -2578 2732 -2563
rect 2780 -2578 2827 -2563
rect 1884 -2657 1900 -2629
rect 1950 -2657 2004 -2579
rect 2139 -2610 2186 -2578
rect 1834 -2691 1900 -2657
rect 1834 -2725 1850 -2691
rect 1884 -2725 1900 -2691
rect 1834 -2759 1900 -2725
rect 1834 -2793 1850 -2759
rect 1884 -2793 1900 -2759
rect 1834 -2798 1900 -2793
rect 1938 -2697 2004 -2657
rect 1938 -2731 1954 -2697
rect 1988 -2731 2004 -2697
rect 1938 -2765 2004 -2731
rect 1938 -2799 1954 -2765
rect 1988 -2799 2004 -2765
rect 1938 -2803 2004 -2799
rect 2042 -2629 2085 -2613
rect 2042 -2663 2051 -2629
rect 2042 -2697 2085 -2663
rect 2042 -2731 2051 -2697
rect 2042 -2765 2085 -2731
rect 2042 -2799 2051 -2765
rect 2042 -2841 2085 -2799
rect 2119 -2623 2186 -2610
rect 2368 -2611 2414 -2578
rect 2501 -2579 2827 -2578
rect 2861 -2576 2864 -2528
rect 2912 -2576 2914 -2528
rect 2119 -2657 2135 -2623
rect 2169 -2657 2186 -2623
rect 2119 -2694 2186 -2657
rect 2119 -2728 2135 -2694
rect 2169 -2728 2186 -2694
rect 2119 -2765 2186 -2728
rect 2119 -2799 2135 -2765
rect 2169 -2799 2186 -2765
rect 2119 -2807 2186 -2799
rect 2272 -2629 2314 -2613
rect 2272 -2663 2280 -2629
rect 2272 -2697 2314 -2663
rect 2272 -2731 2280 -2697
rect 2272 -2765 2314 -2731
rect 2272 -2799 2280 -2765
rect 2272 -2841 2314 -2799
rect 2348 -2629 2414 -2611
rect 2861 -2613 2914 -2576
rect 2348 -2663 2364 -2629
rect 2398 -2663 2414 -2629
rect 2348 -2697 2414 -2663
rect 2348 -2731 2364 -2697
rect 2398 -2731 2414 -2697
rect 2348 -2765 2414 -2731
rect 2348 -2799 2364 -2765
rect 2398 -2799 2414 -2765
rect 2348 -2807 2414 -2799
rect 2506 -2629 2559 -2613
rect 2506 -2663 2525 -2629
rect 2506 -2697 2559 -2663
rect 2506 -2731 2525 -2697
rect 2506 -2765 2559 -2731
rect 2506 -2799 2525 -2765
rect 2506 -2841 2559 -2799
rect 2593 -2629 2914 -2613
rect 2593 -2663 2609 -2629
rect 2643 -2647 2777 -2629
rect 2643 -2663 2659 -2647
rect 2593 -2697 2659 -2663
rect 2761 -2663 2777 -2647
rect 2811 -2651 2914 -2629
rect 3207 -2643 3265 -2608
rect 2811 -2663 2827 -2651
rect 2593 -2731 2609 -2697
rect 2643 -2731 2659 -2697
rect 2593 -2765 2659 -2731
rect 2593 -2799 2609 -2765
rect 2643 -2799 2659 -2765
rect 2593 -2807 2659 -2799
rect 2693 -2697 2727 -2681
rect 2693 -2765 2727 -2731
rect 2693 -2841 2727 -2799
rect 2761 -2697 2827 -2663
rect 2761 -2731 2777 -2697
rect 2811 -2731 2827 -2697
rect 2761 -2765 2827 -2731
rect 3207 -2677 3219 -2643
rect 3253 -2677 3265 -2643
rect 3207 -2736 3265 -2677
rect 2761 -2799 2777 -2765
rect 2811 -2799 2827 -2765
rect 2761 -2807 2827 -2799
rect 2861 -2765 2903 -2749
rect 2895 -2799 2903 -2765
rect 2861 -2841 2903 -2799
rect 3207 -2770 3219 -2736
rect 3253 -2770 3265 -2736
rect 3207 -2841 3265 -2770
rect -2584 -2875 -2555 -2841
rect -2521 -2875 -2492 -2841
rect -2242 -2875 -2213 -2841
rect -2179 -2875 -2121 -2841
rect -2087 -2875 -2029 -2841
rect -1995 -2875 -1937 -2841
rect -1903 -2875 -1845 -2841
rect -1811 -2875 -1753 -2841
rect -1719 -2875 -1661 -2841
rect -1627 -2875 -1569 -2841
rect -1535 -2875 -1477 -2841
rect -1443 -2875 -1385 -2841
rect -1351 -2875 -1293 -2841
rect -1259 -2875 -1201 -2841
rect -1167 -2875 -1109 -2841
rect -1075 -2875 -1017 -2841
rect -983 -2875 -925 -2841
rect -891 -2875 -833 -2841
rect -799 -2875 -741 -2841
rect -707 -2875 -649 -2841
rect -615 -2875 -557 -2841
rect -523 -2875 -465 -2841
rect -431 -2875 -373 -2841
rect -339 -2875 -281 -2841
rect -247 -2875 -189 -2841
rect -155 -2875 -97 -2841
rect -63 -2875 -5 -2841
rect 29 -2875 87 -2841
rect 121 -2875 179 -2841
rect 213 -2875 242 -2841
rect 456 -2875 485 -2841
rect 519 -2875 577 -2841
rect 611 -2875 669 -2841
rect 703 -2875 761 -2841
rect 795 -2875 853 -2841
rect 887 -2875 945 -2841
rect 979 -2875 1037 -2841
rect 1071 -2875 1129 -2841
rect 1163 -2875 1221 -2841
rect 1255 -2875 1313 -2841
rect 1347 -2875 1405 -2841
rect 1439 -2875 1497 -2841
rect 1531 -2875 1589 -2841
rect 1623 -2875 1681 -2841
rect 1715 -2875 1773 -2841
rect 1807 -2875 1865 -2841
rect 1899 -2875 1957 -2841
rect 1991 -2875 2049 -2841
rect 2083 -2875 2141 -2841
rect 2175 -2875 2233 -2841
rect 2267 -2875 2325 -2841
rect 2359 -2875 2417 -2841
rect 2451 -2875 2509 -2841
rect 2543 -2875 2601 -2841
rect 2635 -2875 2693 -2841
rect 2727 -2875 2785 -2841
rect 2819 -2875 2877 -2841
rect 2911 -2875 2940 -2841
rect 3190 -2875 3219 -2841
rect 3253 -2875 3282 -2841
<< viali >>
rect -2555 389 -2521 423
rect -2213 389 -2179 423
rect -2121 389 -2087 423
rect -2029 389 -1995 423
rect -1937 389 -1903 423
rect -1845 389 -1811 423
rect -1753 389 -1719 423
rect -1661 389 -1627 423
rect -1569 389 -1535 423
rect -1477 389 -1443 423
rect -1385 389 -1351 423
rect -1293 389 -1259 423
rect -1201 389 -1167 423
rect -1109 389 -1075 423
rect -1017 389 -983 423
rect -925 389 -891 423
rect -833 389 -799 423
rect -741 389 -707 423
rect -649 389 -615 423
rect -557 389 -523 423
rect -465 389 -431 423
rect -373 389 -339 423
rect -281 389 -247 423
rect -189 389 -155 423
rect -97 389 -63 423
rect -5 389 29 423
rect 87 389 121 423
rect 179 389 213 423
rect 345 389 379 423
rect 3219 389 3253 423
rect -2116 219 -2082 253
rect -2214 111 -2166 146
rect -2214 98 -2210 111
rect -2210 98 -2176 111
rect -2176 98 -2166 111
rect -2037 151 -2003 185
rect -1962 40 -1914 88
rect -1696 227 -1662 253
rect -1696 219 -1694 227
rect -1694 219 -1662 227
rect -1799 151 -1765 185
rect -1382 219 -1348 253
rect -1295 151 -1261 185
rect -552 78 -504 126
rect -436 111 -388 126
rect -436 78 -414 111
rect -414 78 -388 111
rect -858 -8 -846 8
rect -846 -8 -812 8
rect -812 -8 -810 8
rect -858 -40 -810 -8
rect -324 78 -276 126
rect -192 111 -144 126
rect -82 111 -34 126
rect 34 111 82 126
rect -192 78 -181 111
rect -181 78 -147 111
rect -147 78 -144 111
rect -82 78 -55 111
rect -55 78 -34 111
rect 34 78 79 111
rect 79 78 82 111
rect 166 76 214 124
rect -2555 -155 -2521 -121
rect -2213 -155 -2179 -121
rect -2121 -155 -2087 -121
rect -2029 -155 -1995 -121
rect -1937 -155 -1903 -121
rect -1845 -155 -1811 -121
rect -1753 -155 -1719 -121
rect -1661 -155 -1627 -121
rect -1569 -155 -1535 -121
rect -1477 -155 -1443 -121
rect -1385 -155 -1351 -121
rect -1293 -155 -1259 -121
rect -1201 -155 -1167 -121
rect -1109 -155 -1075 -121
rect -1017 -155 -983 -121
rect -925 -155 -891 -121
rect -833 -155 -799 -121
rect -741 -155 -707 -121
rect -649 -155 -615 -121
rect -557 -155 -523 -121
rect -465 -155 -431 -121
rect -373 -155 -339 -121
rect -281 -155 -247 -121
rect -189 -155 -155 -121
rect -97 -155 -63 -121
rect -5 -155 29 -121
rect 87 -155 121 -121
rect 179 -155 213 -121
rect 345 -155 379 -121
rect 485 -155 519 -121
rect 577 -155 611 -121
rect 669 -155 703 -121
rect 761 -155 795 -121
rect 853 -155 887 -121
rect 945 -155 979 -121
rect 1037 -155 1071 -121
rect 1129 -155 1163 -121
rect 1221 -155 1255 -121
rect 1313 -155 1347 -121
rect 1405 -155 1439 -121
rect 1497 -155 1531 -121
rect 1589 -155 1623 -121
rect 1681 -155 1715 -121
rect 1773 -155 1807 -121
rect 1865 -155 1899 -121
rect 1957 -155 1991 -121
rect 2049 -155 2083 -121
rect 2141 -155 2175 -121
rect 2233 -155 2267 -121
rect 2325 -155 2359 -121
rect 2417 -155 2451 -121
rect 2509 -155 2543 -121
rect 2601 -155 2635 -121
rect 2693 -155 2727 -121
rect 2785 -155 2819 -121
rect 2877 -155 2911 -121
rect 3219 -155 3253 -121
rect -2218 -387 -2210 -364
rect -2210 -387 -2176 -364
rect -2176 -387 -2170 -364
rect -2218 -412 -2170 -387
rect -2116 -529 -2082 -495
rect -2037 -461 -2003 -427
rect -1962 -364 -1914 -316
rect -1799 -461 -1765 -427
rect -1696 -503 -1694 -495
rect -1694 -503 -1662 -495
rect -1696 -529 -1662 -503
rect -1382 -529 -1348 -495
rect -1295 -461 -1261 -427
rect -552 -402 -504 -354
rect -436 -387 -414 -354
rect -414 -387 -388 -354
rect -436 -402 -388 -387
rect -324 -402 -276 -354
rect -192 -387 -181 -354
rect -181 -387 -147 -354
rect -147 -387 -144 -354
rect -82 -387 -55 -354
rect -55 -387 -34 -354
rect 34 -387 79 -354
rect 79 -387 82 -354
rect -192 -402 -144 -387
rect -82 -402 -34 -387
rect 34 -402 82 -387
rect -858 -549 -848 -538
rect -848 -549 -814 -538
rect -814 -549 -810 -538
rect -858 -583 -810 -549
rect -858 -586 -848 -583
rect -848 -586 -814 -583
rect -814 -586 -810 -583
rect 170 -400 218 -352
rect 480 -454 528 -406
rect 582 -529 616 -495
rect 661 -461 695 -427
rect 736 -364 784 -316
rect 899 -461 933 -427
rect 1002 -503 1004 -495
rect 1004 -503 1036 -495
rect 1002 -529 1036 -503
rect 1316 -529 1350 -495
rect 1403 -461 1437 -427
rect 1842 -268 1890 -240
rect 1842 -288 1852 -268
rect 1852 -288 1886 -268
rect 1886 -288 1890 -268
rect 2146 -402 2194 -354
rect 2262 -387 2284 -354
rect 2284 -387 2310 -354
rect 2262 -402 2310 -387
rect 2374 -402 2422 -354
rect 2506 -387 2517 -354
rect 2517 -387 2551 -354
rect 2551 -387 2554 -354
rect 2616 -387 2643 -354
rect 2643 -387 2664 -354
rect 2732 -387 2777 -354
rect 2777 -387 2780 -354
rect 2506 -402 2554 -387
rect 2616 -402 2664 -387
rect 2732 -402 2780 -387
rect 2864 -400 2912 -352
rect -2555 -699 -2521 -665
rect -2213 -699 -2179 -665
rect -2121 -699 -2087 -665
rect -2029 -699 -1995 -665
rect -1937 -699 -1903 -665
rect -1845 -699 -1811 -665
rect -1753 -699 -1719 -665
rect -1661 -699 -1627 -665
rect -1569 -699 -1535 -665
rect -1477 -699 -1443 -665
rect -1385 -699 -1351 -665
rect -1293 -699 -1259 -665
rect -1201 -699 -1167 -665
rect -1109 -699 -1075 -665
rect -1017 -699 -983 -665
rect -925 -699 -891 -665
rect -833 -699 -799 -665
rect -741 -699 -707 -665
rect -649 -699 -615 -665
rect -557 -699 -523 -665
rect -465 -699 -431 -665
rect -373 -699 -339 -665
rect -281 -699 -247 -665
rect -189 -699 -155 -665
rect -97 -699 -63 -665
rect -5 -699 29 -665
rect 87 -699 121 -665
rect 179 -699 213 -665
rect 485 -699 519 -665
rect 577 -699 611 -665
rect 669 -699 703 -665
rect 761 -699 795 -665
rect 853 -699 887 -665
rect 945 -699 979 -665
rect 1037 -699 1071 -665
rect 1129 -699 1163 -665
rect 1221 -699 1255 -665
rect 1313 -699 1347 -665
rect 1405 -699 1439 -665
rect 1497 -699 1531 -665
rect 1589 -699 1623 -665
rect 1681 -699 1715 -665
rect 1773 -699 1807 -665
rect 1865 -699 1899 -665
rect 1957 -699 1991 -665
rect 2049 -699 2083 -665
rect 2141 -699 2175 -665
rect 2233 -699 2267 -665
rect 2325 -699 2359 -665
rect 2417 -699 2451 -665
rect 2509 -699 2543 -665
rect 2601 -699 2635 -665
rect 2693 -699 2727 -665
rect 2785 -699 2819 -665
rect 2877 -699 2911 -665
rect 3219 -699 3253 -665
rect -2116 -869 -2082 -835
rect -2218 -958 -2170 -910
rect -2037 -937 -2003 -903
rect -1962 -1048 -1914 -1000
rect -1696 -861 -1662 -835
rect -1696 -869 -1694 -861
rect -1694 -869 -1662 -861
rect -1799 -937 -1765 -903
rect -1382 -869 -1348 -835
rect -1295 -937 -1261 -903
rect 582 -869 616 -835
rect -552 -1010 -504 -962
rect -436 -977 -388 -962
rect -436 -1010 -414 -977
rect -414 -1010 -388 -977
rect -858 -1096 -846 -1082
rect -846 -1096 -812 -1082
rect -812 -1096 -810 -1082
rect -858 -1130 -810 -1096
rect -324 -1010 -276 -962
rect -192 -977 -144 -962
rect -82 -977 -34 -962
rect 34 -977 82 -962
rect -192 -1010 -181 -977
rect -181 -1010 -147 -977
rect -147 -1010 -144 -977
rect -82 -1010 -55 -977
rect -55 -1010 -34 -977
rect 34 -1010 79 -977
rect 79 -1010 82 -977
rect 166 -1012 218 -964
rect 480 -977 528 -950
rect 480 -998 488 -977
rect 488 -998 522 -977
rect 522 -998 528 -977
rect 661 -937 695 -903
rect 736 -1048 784 -1000
rect 1002 -861 1036 -835
rect 1002 -869 1004 -861
rect 1004 -869 1036 -861
rect 899 -937 933 -903
rect 1316 -869 1350 -835
rect 1403 -937 1437 -903
rect 1840 -781 1850 -778
rect 1850 -781 1884 -778
rect 1884 -781 1888 -778
rect 1840 -815 1888 -781
rect 1840 -826 1850 -815
rect 1850 -826 1884 -815
rect 1884 -826 1888 -815
rect 2146 -1010 2194 -962
rect 2262 -977 2310 -962
rect 2262 -1010 2284 -977
rect 2284 -1010 2310 -977
rect 2374 -1010 2422 -962
rect 2506 -977 2554 -962
rect 2616 -977 2664 -962
rect 2732 -977 2780 -962
rect 2506 -1010 2517 -977
rect 2517 -1010 2551 -977
rect 2551 -1010 2554 -977
rect 2616 -1010 2643 -977
rect 2643 -1010 2664 -977
rect 2732 -1010 2777 -977
rect 2777 -1010 2780 -977
rect 2864 -1012 2912 -964
rect -2555 -1243 -2521 -1209
rect -2213 -1243 -2179 -1209
rect -2121 -1243 -2087 -1209
rect -2029 -1243 -1995 -1209
rect -1937 -1243 -1903 -1209
rect -1845 -1243 -1811 -1209
rect -1753 -1243 -1719 -1209
rect -1661 -1243 -1627 -1209
rect -1569 -1243 -1535 -1209
rect -1477 -1243 -1443 -1209
rect -1385 -1243 -1351 -1209
rect -1293 -1243 -1259 -1209
rect -1201 -1243 -1167 -1209
rect -1109 -1243 -1075 -1209
rect -1017 -1243 -983 -1209
rect -925 -1243 -891 -1209
rect -833 -1243 -799 -1209
rect -741 -1243 -707 -1209
rect -649 -1243 -615 -1209
rect -557 -1243 -523 -1209
rect -465 -1243 -431 -1209
rect -373 -1243 -339 -1209
rect -281 -1243 -247 -1209
rect -189 -1243 -155 -1209
rect -97 -1243 -63 -1209
rect -5 -1243 29 -1209
rect 87 -1243 121 -1209
rect 179 -1243 213 -1209
rect 485 -1243 519 -1209
rect 577 -1243 611 -1209
rect 669 -1243 703 -1209
rect 761 -1243 795 -1209
rect 853 -1243 887 -1209
rect 945 -1243 979 -1209
rect 1037 -1243 1071 -1209
rect 1129 -1243 1163 -1209
rect 1221 -1243 1255 -1209
rect 1313 -1243 1347 -1209
rect 1405 -1243 1439 -1209
rect 1497 -1243 1531 -1209
rect 1589 -1243 1623 -1209
rect 1681 -1243 1715 -1209
rect 1773 -1243 1807 -1209
rect 1865 -1243 1899 -1209
rect 1957 -1243 1991 -1209
rect 2049 -1243 2083 -1209
rect 2141 -1243 2175 -1209
rect 2233 -1243 2267 -1209
rect 2325 -1243 2359 -1209
rect 2417 -1243 2451 -1209
rect 2509 -1243 2543 -1209
rect 2601 -1243 2635 -1209
rect 2693 -1243 2727 -1209
rect 2785 -1243 2819 -1209
rect 2877 -1243 2911 -1209
rect 3219 -1243 3253 -1209
rect -2218 -1475 -2210 -1454
rect -2210 -1475 -2176 -1454
rect -2176 -1475 -2170 -1454
rect -2218 -1502 -2170 -1475
rect -2116 -1617 -2082 -1583
rect -2037 -1549 -2003 -1515
rect -1962 -1452 -1914 -1404
rect -1799 -1549 -1765 -1515
rect -1696 -1591 -1694 -1583
rect -1694 -1591 -1662 -1583
rect -1696 -1617 -1662 -1591
rect -1382 -1617 -1348 -1583
rect -1295 -1549 -1261 -1515
rect -552 -1490 -504 -1442
rect -436 -1475 -414 -1442
rect -414 -1475 -388 -1442
rect -436 -1490 -388 -1475
rect -324 -1490 -276 -1442
rect -192 -1475 -181 -1442
rect -181 -1475 -147 -1442
rect -147 -1475 -144 -1442
rect -82 -1475 -55 -1442
rect -55 -1475 -34 -1442
rect 34 -1475 79 -1442
rect 79 -1475 82 -1442
rect -192 -1490 -144 -1475
rect -82 -1490 -34 -1475
rect 34 -1490 82 -1475
rect -858 -1637 -848 -1626
rect -848 -1637 -814 -1626
rect -814 -1637 -810 -1626
rect -858 -1671 -810 -1637
rect -858 -1674 -848 -1671
rect -848 -1674 -814 -1671
rect -814 -1674 -810 -1671
rect 166 -1488 214 -1440
rect 480 -1542 528 -1494
rect 582 -1617 616 -1583
rect 661 -1549 695 -1515
rect 736 -1452 784 -1404
rect 899 -1549 933 -1515
rect 1002 -1591 1004 -1583
rect 1004 -1591 1036 -1583
rect 1002 -1617 1036 -1591
rect 1316 -1617 1350 -1583
rect 1403 -1549 1437 -1515
rect 1840 -1356 1888 -1322
rect 1840 -1370 1852 -1356
rect 1852 -1370 1886 -1356
rect 1886 -1370 1888 -1356
rect 2146 -1490 2194 -1442
rect 2262 -1475 2284 -1442
rect 2284 -1475 2310 -1442
rect 2262 -1490 2310 -1475
rect 2374 -1490 2422 -1442
rect 2506 -1475 2517 -1442
rect 2517 -1475 2551 -1442
rect 2551 -1475 2554 -1442
rect 2616 -1475 2643 -1442
rect 2643 -1475 2664 -1442
rect 2732 -1475 2777 -1442
rect 2777 -1475 2780 -1442
rect 2506 -1490 2554 -1475
rect 2616 -1490 2664 -1475
rect 2732 -1490 2780 -1475
rect 2864 -1488 2916 -1440
rect -2555 -1787 -2521 -1753
rect -2213 -1787 -2179 -1753
rect -2121 -1787 -2087 -1753
rect -2029 -1787 -1995 -1753
rect -1937 -1787 -1903 -1753
rect -1845 -1787 -1811 -1753
rect -1753 -1787 -1719 -1753
rect -1661 -1787 -1627 -1753
rect -1569 -1787 -1535 -1753
rect -1477 -1787 -1443 -1753
rect -1385 -1787 -1351 -1753
rect -1293 -1787 -1259 -1753
rect -1201 -1787 -1167 -1753
rect -1109 -1787 -1075 -1753
rect -1017 -1787 -983 -1753
rect -925 -1787 -891 -1753
rect -833 -1787 -799 -1753
rect -741 -1787 -707 -1753
rect -649 -1787 -615 -1753
rect -557 -1787 -523 -1753
rect -465 -1787 -431 -1753
rect -373 -1787 -339 -1753
rect -281 -1787 -247 -1753
rect -189 -1787 -155 -1753
rect -97 -1787 -63 -1753
rect -5 -1787 29 -1753
rect 87 -1787 121 -1753
rect 179 -1787 213 -1753
rect 485 -1787 519 -1753
rect 577 -1787 611 -1753
rect 669 -1787 703 -1753
rect 761 -1787 795 -1753
rect 853 -1787 887 -1753
rect 945 -1787 979 -1753
rect 1037 -1787 1071 -1753
rect 1129 -1787 1163 -1753
rect 1221 -1787 1255 -1753
rect 1313 -1787 1347 -1753
rect 1405 -1787 1439 -1753
rect 1497 -1787 1531 -1753
rect 1589 -1787 1623 -1753
rect 1681 -1787 1715 -1753
rect 1773 -1787 1807 -1753
rect 1865 -1787 1899 -1753
rect 1957 -1787 1991 -1753
rect 2049 -1787 2083 -1753
rect 2141 -1787 2175 -1753
rect 2233 -1787 2267 -1753
rect 2325 -1787 2359 -1753
rect 2417 -1787 2451 -1753
rect 2509 -1787 2543 -1753
rect 2601 -1787 2635 -1753
rect 2693 -1787 2727 -1753
rect 2785 -1787 2819 -1753
rect 2877 -1787 2911 -1753
rect 3219 -1787 3253 -1753
rect -2116 -1957 -2082 -1923
rect -2218 -2046 -2170 -1998
rect -2037 -2025 -2003 -1991
rect -1962 -2136 -1914 -2088
rect -1696 -1949 -1662 -1923
rect -1696 -1957 -1694 -1949
rect -1694 -1957 -1662 -1949
rect -1799 -2025 -1765 -1991
rect -1382 -1957 -1348 -1923
rect -1295 -2025 -1261 -1991
rect 582 -1957 616 -1923
rect -552 -2098 -504 -2050
rect -436 -2065 -388 -2050
rect -436 -2098 -414 -2065
rect -414 -2098 -388 -2065
rect -858 -2184 -846 -2168
rect -846 -2184 -812 -2168
rect -812 -2184 -810 -2168
rect -858 -2216 -810 -2184
rect -324 -2098 -276 -2050
rect -192 -2065 -144 -2050
rect -82 -2065 -34 -2050
rect 34 -2065 82 -2050
rect -192 -2098 -181 -2065
rect -181 -2098 -147 -2065
rect -147 -2098 -144 -2065
rect -82 -2098 -55 -2065
rect -55 -2098 -34 -2065
rect 34 -2098 79 -2065
rect 79 -2098 82 -2065
rect 166 -2100 214 -2052
rect 480 -2065 528 -2040
rect 480 -2088 488 -2065
rect 488 -2088 522 -2065
rect 522 -2088 528 -2065
rect 661 -2025 695 -1991
rect 736 -2136 784 -2088
rect 1002 -1949 1036 -1923
rect 1002 -1957 1004 -1949
rect 1004 -1957 1036 -1949
rect 899 -2025 933 -1991
rect 1316 -1957 1350 -1923
rect 1403 -2025 1437 -1991
rect 1840 -1869 1850 -1866
rect 1850 -1869 1884 -1866
rect 1884 -1869 1888 -1866
rect 1840 -1903 1888 -1869
rect 1840 -1914 1850 -1903
rect 1850 -1914 1884 -1903
rect 1884 -1914 1888 -1903
rect 2146 -2098 2194 -2050
rect 2262 -2065 2310 -2050
rect 2262 -2098 2284 -2065
rect 2284 -2098 2310 -2065
rect 2374 -2098 2422 -2050
rect 2506 -2065 2554 -2050
rect 2616 -2065 2664 -2050
rect 2732 -2065 2780 -2050
rect 2506 -2098 2517 -2065
rect 2517 -2098 2551 -2065
rect 2551 -2098 2554 -2065
rect 2616 -2098 2643 -2065
rect 2643 -2098 2664 -2065
rect 2732 -2098 2777 -2065
rect 2777 -2098 2780 -2065
rect 2868 -2100 2916 -2052
rect -2555 -2331 -2521 -2297
rect -2213 -2331 -2179 -2297
rect -2121 -2331 -2087 -2297
rect -2029 -2331 -1995 -2297
rect -1937 -2331 -1903 -2297
rect -1845 -2331 -1811 -2297
rect -1753 -2331 -1719 -2297
rect -1661 -2331 -1627 -2297
rect -1569 -2331 -1535 -2297
rect -1477 -2331 -1443 -2297
rect -1385 -2331 -1351 -2297
rect -1293 -2331 -1259 -2297
rect -1201 -2331 -1167 -2297
rect -1109 -2331 -1075 -2297
rect -1017 -2331 -983 -2297
rect -925 -2331 -891 -2297
rect -833 -2331 -799 -2297
rect -741 -2331 -707 -2297
rect -649 -2331 -615 -2297
rect -557 -2331 -523 -2297
rect -465 -2331 -431 -2297
rect -373 -2331 -339 -2297
rect -281 -2331 -247 -2297
rect -189 -2331 -155 -2297
rect -97 -2331 -63 -2297
rect -5 -2331 29 -2297
rect 87 -2331 121 -2297
rect 179 -2331 213 -2297
rect 485 -2331 519 -2297
rect 577 -2331 611 -2297
rect 669 -2331 703 -2297
rect 761 -2331 795 -2297
rect 853 -2331 887 -2297
rect 945 -2331 979 -2297
rect 1037 -2331 1071 -2297
rect 1129 -2331 1163 -2297
rect 1221 -2331 1255 -2297
rect 1313 -2331 1347 -2297
rect 1405 -2331 1439 -2297
rect 1497 -2331 1531 -2297
rect 1589 -2331 1623 -2297
rect 1681 -2331 1715 -2297
rect 1773 -2331 1807 -2297
rect 1865 -2331 1899 -2297
rect 1957 -2331 1991 -2297
rect 2049 -2331 2083 -2297
rect 2141 -2331 2175 -2297
rect 2233 -2331 2267 -2297
rect 2325 -2331 2359 -2297
rect 2417 -2331 2451 -2297
rect 2509 -2331 2543 -2297
rect 2601 -2331 2635 -2297
rect 2693 -2331 2727 -2297
rect 2785 -2331 2819 -2297
rect 2877 -2331 2911 -2297
rect 3219 -2331 3253 -2297
rect -2218 -2563 -2210 -2540
rect -2210 -2563 -2176 -2540
rect -2176 -2563 -2170 -2540
rect -2218 -2588 -2170 -2563
rect -2116 -2705 -2082 -2671
rect -2037 -2637 -2003 -2603
rect -1962 -2540 -1914 -2492
rect -1799 -2637 -1765 -2603
rect -1696 -2679 -1694 -2671
rect -1694 -2679 -1662 -2671
rect -1696 -2705 -1662 -2679
rect -1382 -2705 -1348 -2671
rect -1295 -2637 -1261 -2603
rect -552 -2578 -504 -2530
rect -436 -2563 -414 -2530
rect -414 -2563 -388 -2530
rect -436 -2578 -388 -2563
rect -324 -2578 -276 -2530
rect -192 -2563 -181 -2530
rect -181 -2563 -147 -2530
rect -147 -2563 -144 -2530
rect -82 -2563 -55 -2530
rect -55 -2563 -34 -2530
rect 34 -2563 79 -2530
rect 79 -2563 82 -2530
rect -192 -2578 -144 -2563
rect -82 -2578 -34 -2563
rect 34 -2578 82 -2563
rect -858 -2725 -848 -2712
rect -848 -2725 -814 -2712
rect -814 -2725 -810 -2712
rect -858 -2759 -810 -2725
rect -858 -2760 -848 -2759
rect -848 -2760 -814 -2759
rect -814 -2760 -810 -2759
rect 166 -2576 218 -2528
rect 488 -2529 536 -2522
rect 488 -2563 522 -2529
rect 522 -2563 536 -2529
rect 488 -2570 536 -2563
rect 582 -2705 616 -2671
rect 661 -2637 695 -2603
rect 736 -2540 784 -2492
rect 899 -2637 933 -2603
rect 1002 -2679 1004 -2671
rect 1004 -2679 1036 -2671
rect 1002 -2705 1036 -2679
rect 1316 -2705 1350 -2671
rect 1403 -2637 1437 -2603
rect 1840 -2444 1888 -2412
rect 1840 -2460 1852 -2444
rect 1852 -2460 1886 -2444
rect 1886 -2460 1888 -2444
rect 2146 -2578 2194 -2530
rect 2262 -2563 2284 -2530
rect 2284 -2563 2310 -2530
rect 2262 -2578 2310 -2563
rect 2374 -2578 2422 -2530
rect 2506 -2563 2517 -2530
rect 2517 -2563 2551 -2530
rect 2551 -2563 2554 -2530
rect 2616 -2563 2643 -2530
rect 2643 -2563 2664 -2530
rect 2732 -2563 2777 -2530
rect 2777 -2563 2780 -2530
rect 2506 -2578 2554 -2563
rect 2616 -2578 2664 -2563
rect 2732 -2578 2780 -2563
rect 2864 -2576 2912 -2528
rect -2555 -2875 -2521 -2841
rect -2213 -2875 -2179 -2841
rect -2121 -2875 -2087 -2841
rect -2029 -2875 -1995 -2841
rect -1937 -2875 -1903 -2841
rect -1845 -2875 -1811 -2841
rect -1753 -2875 -1719 -2841
rect -1661 -2875 -1627 -2841
rect -1569 -2875 -1535 -2841
rect -1477 -2875 -1443 -2841
rect -1385 -2875 -1351 -2841
rect -1293 -2875 -1259 -2841
rect -1201 -2875 -1167 -2841
rect -1109 -2875 -1075 -2841
rect -1017 -2875 -983 -2841
rect -925 -2875 -891 -2841
rect -833 -2875 -799 -2841
rect -741 -2875 -707 -2841
rect -649 -2875 -615 -2841
rect -557 -2875 -523 -2841
rect -465 -2875 -431 -2841
rect -373 -2875 -339 -2841
rect -281 -2875 -247 -2841
rect -189 -2875 -155 -2841
rect -97 -2875 -63 -2841
rect -5 -2875 29 -2841
rect 87 -2875 121 -2841
rect 179 -2875 213 -2841
rect 485 -2875 519 -2841
rect 577 -2875 611 -2841
rect 669 -2875 703 -2841
rect 761 -2875 795 -2841
rect 853 -2875 887 -2841
rect 945 -2875 979 -2841
rect 1037 -2875 1071 -2841
rect 1129 -2875 1163 -2841
rect 1221 -2875 1255 -2841
rect 1313 -2875 1347 -2841
rect 1405 -2875 1439 -2841
rect 1497 -2875 1531 -2841
rect 1589 -2875 1623 -2841
rect 1681 -2875 1715 -2841
rect 1773 -2875 1807 -2841
rect 1865 -2875 1899 -2841
rect 1957 -2875 1991 -2841
rect 2049 -2875 2083 -2841
rect 2141 -2875 2175 -2841
rect 2233 -2875 2267 -2841
rect 2325 -2875 2359 -2841
rect 2417 -2875 2451 -2841
rect 2509 -2875 2543 -2841
rect 2601 -2875 2635 -2841
rect 2693 -2875 2727 -2841
rect 2785 -2875 2819 -2841
rect 2877 -2875 2911 -2841
rect 3219 -2875 3253 -2841
<< metal1 >>
rect -2584 442 3282 454
rect -2584 423 292 442
rect 388 423 3282 442
rect -2584 389 -2555 423
rect -2521 389 -2213 423
rect -2179 389 -2121 423
rect -2087 389 -2029 423
rect -1995 389 -1937 423
rect -1903 389 -1845 423
rect -1811 389 -1753 423
rect -1719 389 -1661 423
rect -1627 389 -1569 423
rect -1535 389 -1477 423
rect -1443 389 -1385 423
rect -1351 389 -1293 423
rect -1259 389 -1201 423
rect -1167 389 -1109 423
rect -1075 389 -1017 423
rect -983 389 -925 423
rect -891 389 -833 423
rect -799 389 -741 423
rect -707 389 -649 423
rect -615 389 -557 423
rect -523 389 -465 423
rect -431 389 -373 423
rect -339 389 -281 423
rect -247 389 -189 423
rect -155 389 -97 423
rect -63 389 -5 423
rect 29 389 87 423
rect 121 389 179 423
rect 213 389 292 423
rect 388 389 3219 423
rect 3253 389 3282 423
rect -2584 370 292 389
rect 388 370 3282 389
rect -2584 358 3282 370
rect -2128 253 -2070 259
rect -2128 219 -2116 253
rect -2082 250 -2070 253
rect -1708 253 -1650 259
rect -1708 250 -1696 253
rect -2082 222 -1696 250
rect -2082 219 -2070 222
rect -2128 213 -2070 219
rect -1708 219 -1696 222
rect -1662 250 -1650 253
rect -1394 253 -1336 259
rect -1394 250 -1382 253
rect -1662 222 -1382 250
rect -1662 219 -1650 222
rect -1708 213 -1650 219
rect -1394 219 -1382 222
rect -1348 219 -1336 253
rect -1394 213 -1336 219
rect -2049 185 -1991 191
rect -2674 146 -2154 152
rect -2674 98 -2214 146
rect -2166 98 -2154 146
rect -2049 151 -2037 185
rect -2003 182 -1991 185
rect -1811 185 -1753 191
rect -1811 182 -1799 185
rect -2003 154 -1799 182
rect -2003 151 -1991 154
rect -2049 145 -1991 151
rect -1811 151 -1799 154
rect -1765 182 -1753 185
rect -1307 185 -1249 191
rect -1307 182 -1295 185
rect -1765 154 -1295 182
rect -1765 151 -1753 154
rect -1811 145 -1753 151
rect -1307 151 -1295 154
rect -1261 151 -1249 185
rect -1307 145 -1249 151
rect -564 126 -376 132
rect -2674 92 -2154 98
rect -1968 94 -1908 100
rect -1974 34 -1968 94
rect -1908 34 -1902 94
rect -564 78 -552 126
rect -504 78 -436 126
rect -388 78 -376 126
rect -564 72 -376 78
rect -336 126 94 132
rect 160 130 220 136
rect -336 78 -324 126
rect -276 78 -192 126
rect -144 78 -82 126
rect -34 78 34 126
rect 82 78 94 126
rect -336 72 94 78
rect 154 70 160 130
rect 220 70 226 130
rect 160 64 220 70
rect -1968 28 -1908 34
rect -864 14 -804 20
rect -870 -46 -864 14
rect -804 -46 -798 14
rect -864 -52 -804 -46
rect -2584 -102 3282 -90
rect -2584 -121 -2388 -102
rect -2584 -155 -2555 -121
rect -2521 -155 -2388 -121
rect -2584 -174 -2388 -155
rect -2292 -121 2990 -102
rect -2292 -155 -2213 -121
rect -2179 -155 -2121 -121
rect -2087 -155 -2029 -121
rect -1995 -155 -1937 -121
rect -1903 -155 -1845 -121
rect -1811 -155 -1753 -121
rect -1719 -155 -1661 -121
rect -1627 -155 -1569 -121
rect -1535 -155 -1477 -121
rect -1443 -155 -1385 -121
rect -1351 -155 -1293 -121
rect -1259 -155 -1201 -121
rect -1167 -155 -1109 -121
rect -1075 -155 -1017 -121
rect -983 -155 -925 -121
rect -891 -155 -833 -121
rect -799 -155 -741 -121
rect -707 -155 -649 -121
rect -615 -155 -557 -121
rect -523 -155 -465 -121
rect -431 -155 -373 -121
rect -339 -155 -281 -121
rect -247 -155 -189 -121
rect -155 -155 -97 -121
rect -63 -155 -5 -121
rect 29 -155 87 -121
rect 121 -155 179 -121
rect 213 -155 345 -121
rect 379 -155 485 -121
rect 519 -155 577 -121
rect 611 -155 669 -121
rect 703 -155 761 -121
rect 795 -155 853 -121
rect 887 -155 945 -121
rect 979 -155 1037 -121
rect 1071 -155 1129 -121
rect 1163 -155 1221 -121
rect 1255 -155 1313 -121
rect 1347 -155 1405 -121
rect 1439 -155 1497 -121
rect 1531 -155 1589 -121
rect 1623 -155 1681 -121
rect 1715 -155 1773 -121
rect 1807 -155 1865 -121
rect 1899 -155 1957 -121
rect 1991 -155 2049 -121
rect 2083 -155 2141 -121
rect 2175 -155 2233 -121
rect 2267 -155 2325 -121
rect 2359 -155 2417 -121
rect 2451 -155 2509 -121
rect 2543 -155 2601 -121
rect 2635 -155 2693 -121
rect 2727 -155 2785 -121
rect 2819 -155 2877 -121
rect 2911 -155 2990 -121
rect -2292 -174 2990 -155
rect 3086 -121 3282 -102
rect 3086 -155 3219 -121
rect 3253 -155 3282 -121
rect 3086 -174 3282 -155
rect -2584 -186 3282 -174
rect 1836 -234 1896 -228
rect 1830 -294 1836 -234
rect 1896 -294 1902 -234
rect 1836 -300 1896 -294
rect -1968 -310 -1908 -304
rect 730 -310 790 -304
rect -2224 -358 -2164 -352
rect -2230 -418 -2224 -358
rect -2164 -418 -2158 -358
rect -1974 -370 -1968 -310
rect -1908 -370 -1902 -310
rect -564 -354 -376 -348
rect -1968 -376 -1908 -370
rect -564 -402 -552 -354
rect -504 -402 -436 -354
rect -388 -402 -376 -354
rect -564 -408 -376 -402
rect -336 -354 94 -348
rect -336 -402 -324 -354
rect -276 -402 -192 -354
rect -144 -402 -82 -354
rect -34 -402 34 -354
rect 82 -402 94 -354
rect -336 -408 94 -402
rect 152 -406 158 -346
rect 218 -406 230 -346
rect 724 -370 730 -310
rect 790 -370 796 -310
rect 2858 -346 2918 -340
rect 2134 -354 2322 -348
rect 730 -376 790 -370
rect 474 -400 534 -394
rect -2224 -424 -2164 -418
rect -2049 -427 -1991 -421
rect -2049 -461 -2037 -427
rect -2003 -430 -1991 -427
rect -1811 -427 -1753 -421
rect -1811 -430 -1799 -427
rect -2003 -458 -1799 -430
rect -2003 -461 -1991 -458
rect -2049 -467 -1991 -461
rect -1811 -461 -1799 -458
rect -1765 -430 -1753 -427
rect -1307 -427 -1249 -421
rect -1307 -430 -1295 -427
rect -1765 -458 -1295 -430
rect -1765 -461 -1753 -458
rect -1811 -467 -1753 -461
rect -1307 -461 -1295 -458
rect -1261 -461 -1249 -427
rect 468 -460 474 -400
rect 534 -460 540 -400
rect 2134 -402 2146 -354
rect 2194 -402 2262 -354
rect 2310 -402 2322 -354
rect 2134 -408 2322 -402
rect 2362 -354 2792 -348
rect 2362 -402 2374 -354
rect 2422 -402 2506 -354
rect 2554 -402 2616 -354
rect 2664 -402 2732 -354
rect 2780 -402 2792 -354
rect 2362 -408 2792 -402
rect 2852 -406 2858 -346
rect 2918 -406 2924 -346
rect 2858 -412 2918 -406
rect 649 -427 707 -421
rect -1307 -467 -1249 -461
rect 474 -466 534 -460
rect 649 -461 661 -427
rect 695 -430 707 -427
rect 887 -427 945 -421
rect 887 -430 899 -427
rect 695 -458 899 -430
rect 695 -461 707 -458
rect 649 -467 707 -461
rect 887 -461 899 -458
rect 933 -430 945 -427
rect 1391 -427 1449 -421
rect 1391 -430 1403 -427
rect 933 -458 1403 -430
rect 933 -461 945 -458
rect 887 -467 945 -461
rect 1391 -461 1403 -458
rect 1437 -461 1449 -427
rect 1391 -467 1449 -461
rect -2128 -495 -2070 -489
rect -2128 -529 -2116 -495
rect -2082 -498 -2070 -495
rect -1708 -495 -1650 -489
rect -1708 -498 -1696 -495
rect -2082 -526 -1696 -498
rect -2082 -529 -2070 -526
rect -2128 -535 -2070 -529
rect -1708 -529 -1696 -526
rect -1662 -498 -1650 -495
rect -1394 -495 -1336 -489
rect -1394 -498 -1382 -495
rect -1662 -526 -1382 -498
rect -1662 -529 -1650 -526
rect -1708 -535 -1650 -529
rect -1394 -529 -1382 -526
rect -1348 -529 -1336 -495
rect 570 -495 628 -489
rect -1394 -535 -1336 -529
rect -864 -532 -804 -526
rect 570 -529 582 -495
rect 616 -498 628 -495
rect 990 -495 1048 -489
rect 990 -498 1002 -495
rect 616 -526 1002 -498
rect 616 -529 628 -526
rect -870 -592 -864 -532
rect -804 -592 -798 -532
rect 570 -535 628 -529
rect 990 -529 1002 -526
rect 1036 -498 1048 -495
rect 1304 -495 1362 -489
rect 1304 -498 1316 -495
rect 1036 -526 1316 -498
rect 1036 -529 1048 -526
rect 990 -535 1048 -529
rect 1304 -529 1316 -526
rect 1350 -529 1362 -495
rect 1304 -535 1362 -529
rect -864 -598 -804 -592
rect -2584 -646 3282 -634
rect -2584 -665 292 -646
rect -2584 -699 -2555 -665
rect -2521 -699 -2213 -665
rect -2179 -699 -2121 -665
rect -2087 -699 -2029 -665
rect -1995 -699 -1937 -665
rect -1903 -699 -1845 -665
rect -1811 -699 -1753 -665
rect -1719 -699 -1661 -665
rect -1627 -699 -1569 -665
rect -1535 -699 -1477 -665
rect -1443 -699 -1385 -665
rect -1351 -699 -1293 -665
rect -1259 -699 -1201 -665
rect -1167 -699 -1109 -665
rect -1075 -699 -1017 -665
rect -983 -699 -925 -665
rect -891 -699 -833 -665
rect -799 -699 -741 -665
rect -707 -699 -649 -665
rect -615 -699 -557 -665
rect -523 -699 -465 -665
rect -431 -699 -373 -665
rect -339 -699 -281 -665
rect -247 -699 -189 -665
rect -155 -699 -97 -665
rect -63 -699 -5 -665
rect 29 -699 87 -665
rect 121 -699 179 -665
rect 213 -699 292 -665
rect -2584 -718 292 -699
rect 388 -665 3282 -646
rect 388 -699 485 -665
rect 519 -699 577 -665
rect 611 -699 669 -665
rect 703 -699 761 -665
rect 795 -699 853 -665
rect 887 -699 945 -665
rect 979 -699 1037 -665
rect 1071 -699 1129 -665
rect 1163 -699 1221 -665
rect 1255 -699 1313 -665
rect 1347 -699 1405 -665
rect 1439 -699 1497 -665
rect 1531 -699 1589 -665
rect 1623 -699 1681 -665
rect 1715 -699 1773 -665
rect 1807 -699 1865 -665
rect 1899 -699 1957 -665
rect 1991 -699 2049 -665
rect 2083 -699 2141 -665
rect 2175 -699 2233 -665
rect 2267 -699 2325 -665
rect 2359 -699 2417 -665
rect 2451 -699 2509 -665
rect 2543 -699 2601 -665
rect 2635 -699 2693 -665
rect 2727 -699 2785 -665
rect 2819 -699 2877 -665
rect 2911 -699 3219 -665
rect 3253 -699 3282 -665
rect 388 -718 3282 -699
rect -2584 -730 3282 -718
rect 1834 -772 1894 -766
rect -2128 -835 -2070 -829
rect -2128 -869 -2116 -835
rect -2082 -838 -2070 -835
rect -1708 -835 -1650 -829
rect -1708 -838 -1696 -835
rect -2082 -866 -1696 -838
rect -2082 -869 -2070 -866
rect -2128 -875 -2070 -869
rect -1708 -869 -1696 -866
rect -1662 -838 -1650 -835
rect -1394 -835 -1336 -829
rect -1394 -838 -1382 -835
rect -1662 -866 -1382 -838
rect -1662 -869 -1650 -866
rect -1708 -875 -1650 -869
rect -1394 -869 -1382 -866
rect -1348 -869 -1336 -835
rect -1394 -875 -1336 -869
rect 570 -835 628 -829
rect 570 -869 582 -835
rect 616 -838 628 -835
rect 990 -835 1048 -829
rect 990 -838 1002 -835
rect 616 -866 1002 -838
rect 616 -869 628 -866
rect 570 -875 628 -869
rect 990 -869 1002 -866
rect 1036 -838 1048 -835
rect 1304 -835 1362 -829
rect 1828 -832 1834 -772
rect 1894 -832 1900 -772
rect 1304 -838 1316 -835
rect 1036 -866 1316 -838
rect 1036 -869 1048 -866
rect 990 -875 1048 -869
rect 1304 -869 1316 -866
rect 1350 -869 1362 -835
rect 1834 -838 1894 -832
rect 1304 -875 1362 -869
rect -2224 -904 -2164 -898
rect -2049 -903 -1991 -897
rect -2230 -964 -2224 -904
rect -2164 -964 -2158 -904
rect -2049 -937 -2037 -903
rect -2003 -906 -1991 -903
rect -1811 -903 -1753 -897
rect -1811 -906 -1799 -903
rect -2003 -934 -1799 -906
rect -2003 -937 -1991 -934
rect -2049 -943 -1991 -937
rect -1811 -937 -1799 -934
rect -1765 -906 -1753 -903
rect -1307 -903 -1249 -897
rect -1307 -906 -1295 -903
rect -1765 -934 -1295 -906
rect -1765 -937 -1753 -934
rect -1811 -943 -1753 -937
rect -1307 -937 -1295 -934
rect -1261 -937 -1249 -903
rect -1307 -943 -1249 -937
rect 649 -903 707 -897
rect 649 -937 661 -903
rect 695 -906 707 -903
rect 887 -903 945 -897
rect 887 -906 899 -903
rect 695 -934 899 -906
rect 695 -937 707 -934
rect 474 -944 534 -938
rect 649 -943 707 -937
rect 887 -937 899 -934
rect 933 -906 945 -903
rect 1391 -903 1449 -897
rect 1391 -906 1403 -903
rect 933 -934 1403 -906
rect 933 -937 945 -934
rect 887 -943 945 -937
rect 1391 -937 1403 -934
rect 1437 -937 1449 -903
rect 1391 -943 1449 -937
rect -564 -962 -376 -956
rect -2224 -970 -2164 -964
rect -1968 -994 -1908 -988
rect -1974 -1054 -1968 -994
rect -1908 -1054 -1902 -994
rect -564 -1010 -552 -962
rect -504 -1010 -436 -962
rect -388 -1010 -376 -962
rect -564 -1016 -376 -1010
rect -336 -962 94 -956
rect 160 -958 220 -952
rect -336 -1010 -324 -962
rect -276 -1010 -192 -962
rect -144 -1010 -82 -962
rect -34 -1010 34 -962
rect 82 -1010 94 -962
rect -336 -1016 94 -1010
rect 154 -1018 160 -958
rect 220 -1018 226 -958
rect 468 -1004 474 -944
rect 534 -1004 540 -944
rect 2134 -962 2322 -956
rect 730 -994 790 -988
rect 474 -1010 534 -1004
rect 160 -1024 220 -1018
rect 724 -1054 730 -994
rect 790 -1054 796 -994
rect 2134 -1010 2146 -962
rect 2194 -1010 2262 -962
rect 2310 -1010 2322 -962
rect 2134 -1016 2322 -1010
rect 2362 -962 2792 -956
rect 2858 -958 2918 -952
rect 2362 -1010 2374 -962
rect 2422 -1010 2506 -962
rect 2554 -1010 2616 -962
rect 2664 -1010 2732 -962
rect 2780 -1010 2792 -962
rect 2362 -1016 2792 -1010
rect 2852 -1018 2858 -958
rect 2918 -1018 2924 -958
rect 2858 -1024 2918 -1018
rect -1968 -1060 -1908 -1054
rect 730 -1060 790 -1054
rect -864 -1076 -804 -1070
rect -870 -1136 -864 -1076
rect -804 -1136 -798 -1076
rect -864 -1142 -804 -1136
rect -2584 -1190 3282 -1178
rect -2584 -1209 -2388 -1190
rect -2584 -1243 -2555 -1209
rect -2521 -1243 -2388 -1209
rect -2584 -1262 -2388 -1243
rect -2292 -1209 2990 -1190
rect -2292 -1243 -2213 -1209
rect -2179 -1243 -2121 -1209
rect -2087 -1243 -2029 -1209
rect -1995 -1243 -1937 -1209
rect -1903 -1243 -1845 -1209
rect -1811 -1243 -1753 -1209
rect -1719 -1243 -1661 -1209
rect -1627 -1243 -1569 -1209
rect -1535 -1243 -1477 -1209
rect -1443 -1243 -1385 -1209
rect -1351 -1243 -1293 -1209
rect -1259 -1243 -1201 -1209
rect -1167 -1243 -1109 -1209
rect -1075 -1243 -1017 -1209
rect -983 -1243 -925 -1209
rect -891 -1243 -833 -1209
rect -799 -1243 -741 -1209
rect -707 -1243 -649 -1209
rect -615 -1243 -557 -1209
rect -523 -1243 -465 -1209
rect -431 -1243 -373 -1209
rect -339 -1243 -281 -1209
rect -247 -1243 -189 -1209
rect -155 -1243 -97 -1209
rect -63 -1243 -5 -1209
rect 29 -1243 87 -1209
rect 121 -1243 179 -1209
rect 213 -1243 485 -1209
rect 519 -1243 577 -1209
rect 611 -1243 669 -1209
rect 703 -1243 761 -1209
rect 795 -1243 853 -1209
rect 887 -1243 945 -1209
rect 979 -1243 1037 -1209
rect 1071 -1243 1129 -1209
rect 1163 -1243 1221 -1209
rect 1255 -1243 1313 -1209
rect 1347 -1243 1405 -1209
rect 1439 -1243 1497 -1209
rect 1531 -1243 1589 -1209
rect 1623 -1243 1681 -1209
rect 1715 -1243 1773 -1209
rect 1807 -1243 1865 -1209
rect 1899 -1243 1957 -1209
rect 1991 -1243 2049 -1209
rect 2083 -1243 2141 -1209
rect 2175 -1243 2233 -1209
rect 2267 -1243 2325 -1209
rect 2359 -1243 2417 -1209
rect 2451 -1243 2509 -1209
rect 2543 -1243 2601 -1209
rect 2635 -1243 2693 -1209
rect 2727 -1243 2785 -1209
rect 2819 -1243 2877 -1209
rect 2911 -1243 2990 -1209
rect -2292 -1262 2990 -1243
rect 3086 -1209 3282 -1190
rect 3086 -1243 3219 -1209
rect 3253 -1243 3282 -1209
rect 3086 -1262 3282 -1243
rect -2584 -1274 3282 -1262
rect 1834 -1316 1894 -1310
rect 1828 -1376 1834 -1316
rect 1894 -1376 1900 -1316
rect 1834 -1382 1894 -1376
rect -1968 -1398 -1908 -1392
rect 730 -1398 790 -1392
rect -2224 -1448 -2164 -1442
rect -2230 -1508 -2224 -1448
rect -2164 -1508 -2158 -1448
rect -1974 -1458 -1968 -1398
rect -1908 -1458 -1902 -1398
rect 160 -1434 220 -1428
rect -564 -1442 -376 -1436
rect -1968 -1464 -1908 -1458
rect -564 -1490 -552 -1442
rect -504 -1490 -436 -1442
rect -388 -1490 -376 -1442
rect -564 -1496 -376 -1490
rect -336 -1442 94 -1436
rect -336 -1490 -324 -1442
rect -276 -1490 -192 -1442
rect -144 -1490 -82 -1442
rect -34 -1490 34 -1442
rect 82 -1490 94 -1442
rect -336 -1496 94 -1490
rect 154 -1494 160 -1434
rect 220 -1494 226 -1434
rect 724 -1458 730 -1398
rect 790 -1458 796 -1398
rect 2858 -1434 2918 -1428
rect 2134 -1442 2322 -1436
rect 730 -1464 790 -1458
rect 474 -1488 534 -1482
rect 160 -1500 220 -1494
rect -2224 -1514 -2164 -1508
rect -2049 -1515 -1991 -1509
rect -2049 -1549 -2037 -1515
rect -2003 -1518 -1991 -1515
rect -1811 -1515 -1753 -1509
rect -1811 -1518 -1799 -1515
rect -2003 -1546 -1799 -1518
rect -2003 -1549 -1991 -1546
rect -2049 -1555 -1991 -1549
rect -1811 -1549 -1799 -1546
rect -1765 -1518 -1753 -1515
rect -1307 -1515 -1249 -1509
rect -1307 -1518 -1295 -1515
rect -1765 -1546 -1295 -1518
rect -1765 -1549 -1753 -1546
rect -1811 -1555 -1753 -1549
rect -1307 -1549 -1295 -1546
rect -1261 -1549 -1249 -1515
rect 468 -1548 474 -1488
rect 534 -1548 540 -1488
rect 2134 -1490 2146 -1442
rect 2194 -1490 2262 -1442
rect 2310 -1490 2322 -1442
rect 2134 -1496 2322 -1490
rect 2362 -1442 2792 -1436
rect 2362 -1490 2374 -1442
rect 2422 -1490 2506 -1442
rect 2554 -1490 2616 -1442
rect 2664 -1490 2732 -1442
rect 2780 -1490 2792 -1442
rect 2362 -1496 2792 -1490
rect 2852 -1494 2858 -1434
rect 2918 -1494 2924 -1434
rect 2858 -1500 2918 -1494
rect 649 -1515 707 -1509
rect -1307 -1555 -1249 -1549
rect 474 -1554 534 -1548
rect 649 -1549 661 -1515
rect 695 -1518 707 -1515
rect 887 -1515 945 -1509
rect 887 -1518 899 -1515
rect 695 -1546 899 -1518
rect 695 -1549 707 -1546
rect 649 -1555 707 -1549
rect 887 -1549 899 -1546
rect 933 -1518 945 -1515
rect 1391 -1515 1449 -1509
rect 1391 -1518 1403 -1515
rect 933 -1546 1403 -1518
rect 933 -1549 945 -1546
rect 887 -1555 945 -1549
rect 1391 -1549 1403 -1546
rect 1437 -1549 1449 -1515
rect 1391 -1555 1449 -1549
rect -2128 -1583 -2070 -1577
rect -2128 -1617 -2116 -1583
rect -2082 -1586 -2070 -1583
rect -1708 -1583 -1650 -1577
rect -1708 -1586 -1696 -1583
rect -2082 -1614 -1696 -1586
rect -2082 -1617 -2070 -1614
rect -2128 -1623 -2070 -1617
rect -1708 -1617 -1696 -1614
rect -1662 -1586 -1650 -1583
rect -1394 -1583 -1336 -1577
rect -1394 -1586 -1382 -1583
rect -1662 -1614 -1382 -1586
rect -1662 -1617 -1650 -1614
rect -1708 -1623 -1650 -1617
rect -1394 -1617 -1382 -1614
rect -1348 -1617 -1336 -1583
rect 570 -1583 628 -1577
rect -1394 -1623 -1336 -1617
rect -864 -1620 -804 -1614
rect 570 -1617 582 -1583
rect 616 -1586 628 -1583
rect 990 -1583 1048 -1577
rect 990 -1586 1002 -1583
rect 616 -1614 1002 -1586
rect 616 -1617 628 -1614
rect -870 -1680 -864 -1620
rect -804 -1680 -798 -1620
rect 570 -1623 628 -1617
rect 990 -1617 1002 -1614
rect 1036 -1586 1048 -1583
rect 1304 -1583 1362 -1577
rect 1304 -1586 1316 -1583
rect 1036 -1614 1316 -1586
rect 1036 -1617 1048 -1614
rect 990 -1623 1048 -1617
rect 1304 -1617 1316 -1614
rect 1350 -1617 1362 -1583
rect 1304 -1623 1362 -1617
rect -864 -1686 -804 -1680
rect -2584 -1734 3282 -1722
rect -2584 -1753 292 -1734
rect -2584 -1787 -2555 -1753
rect -2521 -1787 -2213 -1753
rect -2179 -1787 -2121 -1753
rect -2087 -1787 -2029 -1753
rect -1995 -1787 -1937 -1753
rect -1903 -1787 -1845 -1753
rect -1811 -1787 -1753 -1753
rect -1719 -1787 -1661 -1753
rect -1627 -1787 -1569 -1753
rect -1535 -1787 -1477 -1753
rect -1443 -1787 -1385 -1753
rect -1351 -1787 -1293 -1753
rect -1259 -1787 -1201 -1753
rect -1167 -1787 -1109 -1753
rect -1075 -1787 -1017 -1753
rect -983 -1787 -925 -1753
rect -891 -1787 -833 -1753
rect -799 -1787 -741 -1753
rect -707 -1787 -649 -1753
rect -615 -1787 -557 -1753
rect -523 -1787 -465 -1753
rect -431 -1787 -373 -1753
rect -339 -1787 -281 -1753
rect -247 -1787 -189 -1753
rect -155 -1787 -97 -1753
rect -63 -1787 -5 -1753
rect 29 -1787 87 -1753
rect 121 -1787 179 -1753
rect 213 -1787 292 -1753
rect -2584 -1806 292 -1787
rect 388 -1753 3282 -1734
rect 388 -1787 485 -1753
rect 519 -1787 577 -1753
rect 611 -1787 669 -1753
rect 703 -1787 761 -1753
rect 795 -1787 853 -1753
rect 887 -1787 945 -1753
rect 979 -1787 1037 -1753
rect 1071 -1787 1129 -1753
rect 1163 -1787 1221 -1753
rect 1255 -1787 1313 -1753
rect 1347 -1787 1405 -1753
rect 1439 -1787 1497 -1753
rect 1531 -1787 1589 -1753
rect 1623 -1787 1681 -1753
rect 1715 -1787 1773 -1753
rect 1807 -1787 1865 -1753
rect 1899 -1787 1957 -1753
rect 1991 -1787 2049 -1753
rect 2083 -1787 2141 -1753
rect 2175 -1787 2233 -1753
rect 2267 -1787 2325 -1753
rect 2359 -1787 2417 -1753
rect 2451 -1787 2509 -1753
rect 2543 -1787 2601 -1753
rect 2635 -1787 2693 -1753
rect 2727 -1787 2785 -1753
rect 2819 -1787 2877 -1753
rect 2911 -1787 3219 -1753
rect 3253 -1787 3282 -1753
rect 388 -1806 3282 -1787
rect -2584 -1818 3282 -1806
rect 1834 -1860 1894 -1854
rect -2128 -1923 -2070 -1917
rect -2128 -1957 -2116 -1923
rect -2082 -1926 -2070 -1923
rect -1708 -1923 -1650 -1917
rect -1708 -1926 -1696 -1923
rect -2082 -1954 -1696 -1926
rect -2082 -1957 -2070 -1954
rect -2128 -1963 -2070 -1957
rect -1708 -1957 -1696 -1954
rect -1662 -1926 -1650 -1923
rect -1394 -1923 -1336 -1917
rect -1394 -1926 -1382 -1923
rect -1662 -1954 -1382 -1926
rect -1662 -1957 -1650 -1954
rect -1708 -1963 -1650 -1957
rect -1394 -1957 -1382 -1954
rect -1348 -1957 -1336 -1923
rect -1394 -1963 -1336 -1957
rect 570 -1923 628 -1917
rect 570 -1957 582 -1923
rect 616 -1926 628 -1923
rect 990 -1923 1048 -1917
rect 990 -1926 1002 -1923
rect 616 -1954 1002 -1926
rect 616 -1957 628 -1954
rect 570 -1963 628 -1957
rect 990 -1957 1002 -1954
rect 1036 -1926 1048 -1923
rect 1304 -1923 1362 -1917
rect 1828 -1920 1834 -1860
rect 1894 -1920 1900 -1860
rect 1304 -1926 1316 -1923
rect 1036 -1954 1316 -1926
rect 1036 -1957 1048 -1954
rect 990 -1963 1048 -1957
rect 1304 -1957 1316 -1954
rect 1350 -1957 1362 -1923
rect 1834 -1926 1894 -1920
rect 1304 -1963 1362 -1957
rect -2224 -1992 -2164 -1986
rect -2049 -1991 -1991 -1985
rect -2230 -2052 -2224 -1992
rect -2164 -2052 -2158 -1992
rect -2049 -2025 -2037 -1991
rect -2003 -1994 -1991 -1991
rect -1811 -1991 -1753 -1985
rect -1811 -1994 -1799 -1991
rect -2003 -2022 -1799 -1994
rect -2003 -2025 -1991 -2022
rect -2049 -2031 -1991 -2025
rect -1811 -2025 -1799 -2022
rect -1765 -1994 -1753 -1991
rect -1307 -1991 -1249 -1985
rect -1307 -1994 -1295 -1991
rect -1765 -2022 -1295 -1994
rect -1765 -2025 -1753 -2022
rect -1811 -2031 -1753 -2025
rect -1307 -2025 -1295 -2022
rect -1261 -2025 -1249 -1991
rect -1307 -2031 -1249 -2025
rect 649 -1991 707 -1985
rect 649 -2025 661 -1991
rect 695 -1994 707 -1991
rect 887 -1991 945 -1985
rect 887 -1994 899 -1991
rect 695 -2022 899 -1994
rect 695 -2025 707 -2022
rect 474 -2034 534 -2028
rect 649 -2031 707 -2025
rect 887 -2025 899 -2022
rect 933 -1994 945 -1991
rect 1391 -1991 1449 -1985
rect 1391 -1994 1403 -1991
rect 933 -2022 1403 -1994
rect 933 -2025 945 -2022
rect 887 -2031 945 -2025
rect 1391 -2025 1403 -2022
rect 1437 -2025 1449 -1991
rect 1391 -2031 1449 -2025
rect -564 -2050 -376 -2044
rect -2224 -2058 -2164 -2052
rect -1968 -2082 -1908 -2076
rect -1974 -2142 -1968 -2082
rect -1908 -2142 -1902 -2082
rect -564 -2098 -552 -2050
rect -504 -2098 -436 -2050
rect -388 -2098 -376 -2050
rect -564 -2104 -376 -2098
rect -336 -2050 94 -2044
rect 160 -2046 220 -2040
rect -336 -2098 -324 -2050
rect -276 -2098 -192 -2050
rect -144 -2098 -82 -2050
rect -34 -2098 34 -2050
rect 82 -2098 94 -2050
rect -336 -2104 94 -2098
rect 154 -2106 160 -2046
rect 220 -2106 226 -2046
rect 468 -2094 474 -2034
rect 534 -2094 540 -2034
rect 2134 -2050 2322 -2044
rect 730 -2082 790 -2076
rect 474 -2100 534 -2094
rect 160 -2112 220 -2106
rect 724 -2142 730 -2082
rect 790 -2142 796 -2082
rect 2134 -2098 2146 -2050
rect 2194 -2098 2262 -2050
rect 2310 -2098 2322 -2050
rect 2134 -2104 2322 -2098
rect 2362 -2050 2792 -2044
rect 2362 -2098 2374 -2050
rect 2422 -2098 2506 -2050
rect 2554 -2098 2616 -2050
rect 2664 -2098 2732 -2050
rect 2780 -2098 2792 -2050
rect 2362 -2104 2792 -2098
rect 2850 -2106 2856 -2046
rect 2916 -2106 2928 -2046
rect -1968 -2148 -1908 -2142
rect 730 -2148 790 -2142
rect -864 -2162 -804 -2156
rect -870 -2222 -864 -2162
rect -804 -2222 -798 -2162
rect -864 -2228 -804 -2222
rect -2584 -2278 3282 -2266
rect -2584 -2297 -2388 -2278
rect -2584 -2331 -2555 -2297
rect -2521 -2331 -2388 -2297
rect -2584 -2350 -2388 -2331
rect -2292 -2297 2990 -2278
rect -2292 -2331 -2213 -2297
rect -2179 -2331 -2121 -2297
rect -2087 -2331 -2029 -2297
rect -1995 -2331 -1937 -2297
rect -1903 -2331 -1845 -2297
rect -1811 -2331 -1753 -2297
rect -1719 -2331 -1661 -2297
rect -1627 -2331 -1569 -2297
rect -1535 -2331 -1477 -2297
rect -1443 -2331 -1385 -2297
rect -1351 -2331 -1293 -2297
rect -1259 -2331 -1201 -2297
rect -1167 -2331 -1109 -2297
rect -1075 -2331 -1017 -2297
rect -983 -2331 -925 -2297
rect -891 -2331 -833 -2297
rect -799 -2331 -741 -2297
rect -707 -2331 -649 -2297
rect -615 -2331 -557 -2297
rect -523 -2331 -465 -2297
rect -431 -2331 -373 -2297
rect -339 -2331 -281 -2297
rect -247 -2331 -189 -2297
rect -155 -2331 -97 -2297
rect -63 -2331 -5 -2297
rect 29 -2331 87 -2297
rect 121 -2331 179 -2297
rect 213 -2331 485 -2297
rect 519 -2331 577 -2297
rect 611 -2331 669 -2297
rect 703 -2331 761 -2297
rect 795 -2331 853 -2297
rect 887 -2331 945 -2297
rect 979 -2331 1037 -2297
rect 1071 -2331 1129 -2297
rect 1163 -2331 1221 -2297
rect 1255 -2331 1313 -2297
rect 1347 -2331 1405 -2297
rect 1439 -2331 1497 -2297
rect 1531 -2331 1589 -2297
rect 1623 -2331 1681 -2297
rect 1715 -2331 1773 -2297
rect 1807 -2331 1865 -2297
rect 1899 -2331 1957 -2297
rect 1991 -2331 2049 -2297
rect 2083 -2331 2141 -2297
rect 2175 -2331 2233 -2297
rect 2267 -2331 2325 -2297
rect 2359 -2331 2417 -2297
rect 2451 -2331 2509 -2297
rect 2543 -2331 2601 -2297
rect 2635 -2331 2693 -2297
rect 2727 -2331 2785 -2297
rect 2819 -2331 2877 -2297
rect 2911 -2331 2990 -2297
rect -2292 -2350 2990 -2331
rect 3086 -2297 3282 -2278
rect 3086 -2331 3219 -2297
rect 3253 -2331 3282 -2297
rect 3086 -2350 3282 -2331
rect -2584 -2362 3282 -2350
rect 1834 -2406 1894 -2400
rect 1828 -2466 1834 -2406
rect 1894 -2466 1900 -2406
rect 1834 -2472 1894 -2466
rect -1968 -2486 -1908 -2480
rect 730 -2486 790 -2480
rect -2224 -2534 -2164 -2528
rect -2230 -2594 -2224 -2534
rect -2164 -2594 -2158 -2534
rect -1974 -2546 -1968 -2486
rect -1908 -2546 -1902 -2486
rect 482 -2516 542 -2510
rect 160 -2522 220 -2516
rect -564 -2530 -376 -2524
rect -1968 -2552 -1908 -2546
rect -564 -2578 -552 -2530
rect -504 -2578 -436 -2530
rect -388 -2578 -376 -2530
rect -564 -2584 -376 -2578
rect -336 -2530 94 -2524
rect -336 -2578 -324 -2530
rect -276 -2578 -192 -2530
rect -144 -2578 -82 -2530
rect -34 -2578 34 -2530
rect 82 -2578 94 -2530
rect -336 -2584 94 -2578
rect 154 -2582 160 -2522
rect 220 -2582 226 -2522
rect 476 -2576 482 -2516
rect 542 -2576 548 -2516
rect 724 -2546 730 -2486
rect 790 -2546 796 -2486
rect 2858 -2522 2918 -2516
rect 2134 -2530 2322 -2524
rect 730 -2552 790 -2546
rect 482 -2582 542 -2576
rect 2134 -2578 2146 -2530
rect 2194 -2578 2262 -2530
rect 2310 -2578 2322 -2530
rect 160 -2588 220 -2582
rect 2134 -2584 2322 -2578
rect 2362 -2530 2792 -2524
rect 2362 -2578 2374 -2530
rect 2422 -2578 2506 -2530
rect 2554 -2578 2616 -2530
rect 2664 -2578 2732 -2530
rect 2780 -2578 2792 -2530
rect 2362 -2584 2792 -2578
rect 2852 -2582 2858 -2522
rect 2918 -2582 2924 -2522
rect 2858 -2588 2918 -2582
rect -2224 -2600 -2164 -2594
rect -2049 -2603 -1991 -2597
rect -2049 -2637 -2037 -2603
rect -2003 -2606 -1991 -2603
rect -1811 -2603 -1753 -2597
rect -1811 -2606 -1799 -2603
rect -2003 -2634 -1799 -2606
rect -2003 -2637 -1991 -2634
rect -2049 -2643 -1991 -2637
rect -1811 -2637 -1799 -2634
rect -1765 -2606 -1753 -2603
rect -1307 -2603 -1249 -2597
rect -1307 -2606 -1295 -2603
rect -1765 -2634 -1295 -2606
rect -1765 -2637 -1753 -2634
rect -1811 -2643 -1753 -2637
rect -1307 -2637 -1295 -2634
rect -1261 -2637 -1249 -2603
rect -1307 -2643 -1249 -2637
rect 649 -2603 707 -2597
rect 649 -2637 661 -2603
rect 695 -2606 707 -2603
rect 887 -2603 945 -2597
rect 887 -2606 899 -2603
rect 695 -2634 899 -2606
rect 695 -2637 707 -2634
rect 649 -2643 707 -2637
rect 887 -2637 899 -2634
rect 933 -2606 945 -2603
rect 1391 -2603 1449 -2597
rect 1391 -2606 1403 -2603
rect 933 -2634 1403 -2606
rect 933 -2637 945 -2634
rect 887 -2643 945 -2637
rect 1391 -2637 1403 -2634
rect 1437 -2637 1449 -2603
rect 1391 -2643 1449 -2637
rect -2128 -2671 -2070 -2665
rect -2128 -2705 -2116 -2671
rect -2082 -2674 -2070 -2671
rect -1708 -2671 -1650 -2665
rect -1708 -2674 -1696 -2671
rect -2082 -2702 -1696 -2674
rect -2082 -2705 -2070 -2702
rect -2128 -2711 -2070 -2705
rect -1708 -2705 -1696 -2702
rect -1662 -2674 -1650 -2671
rect -1394 -2671 -1336 -2665
rect -1394 -2674 -1382 -2671
rect -1662 -2702 -1382 -2674
rect -1662 -2705 -1650 -2702
rect -1708 -2711 -1650 -2705
rect -1394 -2705 -1382 -2702
rect -1348 -2705 -1336 -2671
rect 570 -2671 628 -2665
rect -1394 -2711 -1336 -2705
rect -864 -2706 -804 -2700
rect 570 -2705 582 -2671
rect 616 -2674 628 -2671
rect 990 -2671 1048 -2665
rect 990 -2674 1002 -2671
rect 616 -2702 1002 -2674
rect 616 -2705 628 -2702
rect -870 -2766 -864 -2706
rect -804 -2766 -798 -2706
rect 570 -2711 628 -2705
rect 990 -2705 1002 -2702
rect 1036 -2674 1048 -2671
rect 1304 -2671 1362 -2665
rect 1304 -2674 1316 -2671
rect 1036 -2702 1316 -2674
rect 1036 -2705 1048 -2702
rect 990 -2711 1048 -2705
rect 1304 -2705 1316 -2702
rect 1350 -2705 1362 -2671
rect 1304 -2711 1362 -2705
rect -864 -2772 -804 -2766
rect -2584 -2822 3282 -2810
rect -2584 -2841 292 -2822
rect -2584 -2875 -2555 -2841
rect -2521 -2875 -2213 -2841
rect -2179 -2875 -2121 -2841
rect -2087 -2875 -2029 -2841
rect -1995 -2875 -1937 -2841
rect -1903 -2875 -1845 -2841
rect -1811 -2875 -1753 -2841
rect -1719 -2875 -1661 -2841
rect -1627 -2875 -1569 -2841
rect -1535 -2875 -1477 -2841
rect -1443 -2875 -1385 -2841
rect -1351 -2875 -1293 -2841
rect -1259 -2875 -1201 -2841
rect -1167 -2875 -1109 -2841
rect -1075 -2875 -1017 -2841
rect -983 -2875 -925 -2841
rect -891 -2875 -833 -2841
rect -799 -2875 -741 -2841
rect -707 -2875 -649 -2841
rect -615 -2875 -557 -2841
rect -523 -2875 -465 -2841
rect -431 -2875 -373 -2841
rect -339 -2875 -281 -2841
rect -247 -2875 -189 -2841
rect -155 -2875 -97 -2841
rect -63 -2875 -5 -2841
rect 29 -2875 87 -2841
rect 121 -2875 179 -2841
rect 213 -2875 292 -2841
rect -2584 -2894 292 -2875
rect 388 -2841 3282 -2822
rect 388 -2875 485 -2841
rect 519 -2875 577 -2841
rect 611 -2875 669 -2841
rect 703 -2875 761 -2841
rect 795 -2875 853 -2841
rect 887 -2875 945 -2841
rect 979 -2875 1037 -2841
rect 1071 -2875 1129 -2841
rect 1163 -2875 1221 -2841
rect 1255 -2875 1313 -2841
rect 1347 -2875 1405 -2841
rect 1439 -2875 1497 -2841
rect 1531 -2875 1589 -2841
rect 1623 -2875 1681 -2841
rect 1715 -2875 1773 -2841
rect 1807 -2875 1865 -2841
rect 1899 -2875 1957 -2841
rect 1991 -2875 2049 -2841
rect 2083 -2875 2141 -2841
rect 2175 -2875 2233 -2841
rect 2267 -2875 2325 -2841
rect 2359 -2875 2417 -2841
rect 2451 -2875 2509 -2841
rect 2543 -2875 2601 -2841
rect 2635 -2875 2693 -2841
rect 2727 -2875 2785 -2841
rect 2819 -2875 2877 -2841
rect 2911 -2875 3219 -2841
rect 3253 -2875 3282 -2841
rect 388 -2894 3282 -2875
rect -2584 -2906 3282 -2894
<< via1 >>
rect 292 423 388 442
rect 292 389 345 423
rect 345 389 379 423
rect 379 389 388 423
rect 292 370 388 389
rect -1968 88 -1908 94
rect -1968 40 -1962 88
rect -1962 40 -1914 88
rect -1914 40 -1908 88
rect -1968 34 -1908 40
rect 160 124 220 130
rect 160 76 166 124
rect 166 76 214 124
rect 214 76 220 124
rect 160 70 220 76
rect -864 8 -804 14
rect -864 -40 -858 8
rect -858 -40 -810 8
rect -810 -40 -804 8
rect -864 -46 -804 -40
rect -2388 -174 -2292 -102
rect 2990 -174 3086 -102
rect 1836 -240 1896 -234
rect 1836 -288 1842 -240
rect 1842 -288 1890 -240
rect 1890 -288 1896 -240
rect 1836 -294 1896 -288
rect -2224 -364 -2164 -358
rect -2224 -412 -2218 -364
rect -2218 -412 -2170 -364
rect -2170 -412 -2164 -364
rect -2224 -418 -2164 -412
rect -1968 -316 -1908 -310
rect -1968 -364 -1962 -316
rect -1962 -364 -1914 -316
rect -1914 -364 -1908 -316
rect -1968 -370 -1908 -364
rect 158 -352 218 -346
rect 158 -400 170 -352
rect 170 -400 218 -352
rect 158 -406 218 -400
rect 730 -316 790 -310
rect 730 -364 736 -316
rect 736 -364 784 -316
rect 784 -364 790 -316
rect 730 -370 790 -364
rect 474 -406 534 -400
rect 474 -454 480 -406
rect 480 -454 528 -406
rect 528 -454 534 -406
rect 474 -460 534 -454
rect 2858 -352 2918 -346
rect 2858 -400 2864 -352
rect 2864 -400 2912 -352
rect 2912 -400 2918 -352
rect 2858 -406 2918 -400
rect -864 -538 -804 -532
rect -864 -586 -858 -538
rect -858 -586 -810 -538
rect -810 -586 -804 -538
rect -864 -592 -804 -586
rect 292 -718 388 -646
rect 1834 -778 1894 -772
rect 1834 -826 1840 -778
rect 1840 -826 1888 -778
rect 1888 -826 1894 -778
rect 1834 -832 1894 -826
rect -2224 -910 -2164 -904
rect -2224 -958 -2218 -910
rect -2218 -958 -2170 -910
rect -2170 -958 -2164 -910
rect -2224 -964 -2164 -958
rect -1968 -1000 -1908 -994
rect -1968 -1048 -1962 -1000
rect -1962 -1048 -1914 -1000
rect -1914 -1048 -1908 -1000
rect -1968 -1054 -1908 -1048
rect 160 -964 220 -958
rect 160 -1012 166 -964
rect 166 -1012 218 -964
rect 218 -1012 220 -964
rect 160 -1018 220 -1012
rect 474 -950 534 -944
rect 474 -998 480 -950
rect 480 -998 528 -950
rect 528 -998 534 -950
rect 474 -1004 534 -998
rect 730 -1000 790 -994
rect 730 -1048 736 -1000
rect 736 -1048 784 -1000
rect 784 -1048 790 -1000
rect 730 -1054 790 -1048
rect 2858 -964 2918 -958
rect 2858 -1012 2864 -964
rect 2864 -1012 2912 -964
rect 2912 -1012 2918 -964
rect 2858 -1018 2918 -1012
rect -864 -1082 -804 -1076
rect -864 -1130 -858 -1082
rect -858 -1130 -810 -1082
rect -810 -1130 -804 -1082
rect -864 -1136 -804 -1130
rect -2388 -1262 -2292 -1190
rect 2990 -1262 3086 -1190
rect 1834 -1322 1894 -1316
rect 1834 -1370 1840 -1322
rect 1840 -1370 1888 -1322
rect 1888 -1370 1894 -1322
rect 1834 -1376 1894 -1370
rect -2224 -1454 -2164 -1448
rect -2224 -1502 -2218 -1454
rect -2218 -1502 -2170 -1454
rect -2170 -1502 -2164 -1454
rect -2224 -1508 -2164 -1502
rect -1968 -1404 -1908 -1398
rect -1968 -1452 -1962 -1404
rect -1962 -1452 -1914 -1404
rect -1914 -1452 -1908 -1404
rect -1968 -1458 -1908 -1452
rect 160 -1440 220 -1434
rect 160 -1488 166 -1440
rect 166 -1488 214 -1440
rect 214 -1488 220 -1440
rect 160 -1494 220 -1488
rect 730 -1404 790 -1398
rect 730 -1452 736 -1404
rect 736 -1452 784 -1404
rect 784 -1452 790 -1404
rect 730 -1458 790 -1452
rect 474 -1494 534 -1488
rect 474 -1542 480 -1494
rect 480 -1542 528 -1494
rect 528 -1542 534 -1494
rect 474 -1548 534 -1542
rect 2858 -1440 2918 -1434
rect 2858 -1488 2864 -1440
rect 2864 -1488 2916 -1440
rect 2916 -1488 2918 -1440
rect 2858 -1494 2918 -1488
rect -864 -1626 -804 -1620
rect -864 -1674 -858 -1626
rect -858 -1674 -810 -1626
rect -810 -1674 -804 -1626
rect -864 -1680 -804 -1674
rect 292 -1806 388 -1734
rect 1834 -1866 1894 -1860
rect 1834 -1914 1840 -1866
rect 1840 -1914 1888 -1866
rect 1888 -1914 1894 -1866
rect 1834 -1920 1894 -1914
rect -2224 -1998 -2164 -1992
rect -2224 -2046 -2218 -1998
rect -2218 -2046 -2170 -1998
rect -2170 -2046 -2164 -1998
rect -2224 -2052 -2164 -2046
rect -1968 -2088 -1908 -2082
rect -1968 -2136 -1962 -2088
rect -1962 -2136 -1914 -2088
rect -1914 -2136 -1908 -2088
rect -1968 -2142 -1908 -2136
rect 160 -2052 220 -2046
rect 160 -2100 166 -2052
rect 166 -2100 214 -2052
rect 214 -2100 220 -2052
rect 160 -2106 220 -2100
rect 474 -2040 534 -2034
rect 474 -2088 480 -2040
rect 480 -2088 528 -2040
rect 528 -2088 534 -2040
rect 474 -2094 534 -2088
rect 730 -2088 790 -2082
rect 730 -2136 736 -2088
rect 736 -2136 784 -2088
rect 784 -2136 790 -2088
rect 730 -2142 790 -2136
rect 2856 -2052 2916 -2046
rect 2856 -2100 2868 -2052
rect 2868 -2100 2916 -2052
rect 2856 -2106 2916 -2100
rect -864 -2168 -804 -2162
rect -864 -2216 -858 -2168
rect -858 -2216 -810 -2168
rect -810 -2216 -804 -2168
rect -864 -2222 -804 -2216
rect -2388 -2350 -2292 -2278
rect 2990 -2350 3086 -2278
rect 1834 -2412 1894 -2406
rect 1834 -2460 1840 -2412
rect 1840 -2460 1888 -2412
rect 1888 -2460 1894 -2412
rect 1834 -2466 1894 -2460
rect -2224 -2540 -2164 -2534
rect -2224 -2588 -2218 -2540
rect -2218 -2588 -2170 -2540
rect -2170 -2588 -2164 -2540
rect -2224 -2594 -2164 -2588
rect -1968 -2492 -1908 -2486
rect -1968 -2540 -1962 -2492
rect -1962 -2540 -1914 -2492
rect -1914 -2540 -1908 -2492
rect -1968 -2546 -1908 -2540
rect 160 -2528 220 -2522
rect 160 -2576 166 -2528
rect 166 -2576 218 -2528
rect 218 -2576 220 -2528
rect 160 -2582 220 -2576
rect 482 -2522 542 -2516
rect 482 -2570 488 -2522
rect 488 -2570 536 -2522
rect 536 -2570 542 -2522
rect 482 -2576 542 -2570
rect 730 -2492 790 -2486
rect 730 -2540 736 -2492
rect 736 -2540 784 -2492
rect 784 -2540 790 -2492
rect 730 -2546 790 -2540
rect 2858 -2528 2918 -2522
rect 2858 -2576 2864 -2528
rect 2864 -2576 2912 -2528
rect 2912 -2576 2918 -2528
rect 2858 -2582 2918 -2576
rect -864 -2712 -804 -2706
rect -864 -2760 -858 -2712
rect -858 -2760 -810 -2712
rect -810 -2760 -804 -2712
rect -864 -2766 -804 -2760
rect 292 -2894 388 -2822
<< metal2 >>
rect 280 442 400 454
rect 280 370 292 442
rect 388 370 400 442
rect 280 358 400 370
rect -1968 94 160 130
rect -1908 70 160 94
rect 220 70 226 130
rect -1968 28 -1908 34
rect -864 14 -804 20
rect -2400 -102 -2280 -90
rect -2400 -174 -2388 -102
rect -2292 -174 -2280 -102
rect -864 -106 -804 -46
rect -2400 -186 -2280 -174
rect -2224 -166 -804 -106
rect -2224 -358 -2164 -166
rect 1836 -234 1896 104
rect 2978 -102 3098 -90
rect 2978 -174 2990 -102
rect 3086 -174 3098 -102
rect 2978 -186 3098 -174
rect 1830 -294 1836 -234
rect 1896 -294 1902 -234
rect -1968 -310 -1908 -304
rect 730 -310 790 -304
rect 158 -346 224 -340
rect -1908 -370 158 -346
rect -1968 -406 158 -370
rect 218 -406 224 -346
rect 790 -370 2858 -346
rect 158 -412 224 -406
rect 474 -400 534 -394
rect -2224 -424 -2164 -418
rect 730 -406 2858 -370
rect 2918 -406 2924 -346
rect -864 -532 -804 -526
rect -864 -652 -804 -592
rect -2224 -712 -804 -652
rect 280 -646 400 -634
rect -2224 -904 -2164 -712
rect 280 -718 292 -646
rect 388 -718 400 -646
rect 474 -652 534 -460
rect 474 -712 1894 -652
rect 280 -730 400 -718
rect 1834 -772 1894 -712
rect 1834 -838 1894 -832
rect 474 -944 534 -938
rect -2224 -970 -2164 -964
rect -1968 -994 160 -958
rect -1908 -1018 160 -994
rect 220 -1018 226 -958
rect -1968 -1060 -1908 -1054
rect -864 -1076 -804 -1070
rect -2400 -1190 -2280 -1178
rect -2400 -1262 -2388 -1190
rect -2292 -1262 -2280 -1190
rect -864 -1196 -804 -1136
rect -2400 -1274 -2280 -1262
rect -2224 -1256 -804 -1196
rect 474 -1196 534 -1004
rect 730 -994 2858 -958
rect 790 -1018 2858 -994
rect 2918 -1018 2924 -958
rect 730 -1060 790 -1054
rect 2978 -1190 3098 -1178
rect 474 -1256 1894 -1196
rect -2224 -1448 -2164 -1256
rect 1834 -1316 1894 -1256
rect 2978 -1262 2990 -1190
rect 3086 -1262 3098 -1190
rect 2978 -1274 3098 -1262
rect 1834 -1382 1894 -1376
rect -1968 -1398 -1908 -1392
rect 730 -1398 790 -1392
rect -1908 -1458 160 -1434
rect -1968 -1494 160 -1458
rect 220 -1494 226 -1434
rect 790 -1458 2858 -1434
rect 474 -1488 534 -1482
rect -2224 -1514 -2164 -1508
rect 730 -1494 2858 -1458
rect 2918 -1494 2924 -1434
rect -864 -1620 -804 -1614
rect -864 -1740 -804 -1680
rect -2224 -1800 -804 -1740
rect 280 -1734 400 -1722
rect -2224 -1992 -2164 -1800
rect 280 -1806 292 -1734
rect 388 -1806 400 -1734
rect 474 -1740 534 -1548
rect 474 -1800 1894 -1740
rect 280 -1818 400 -1806
rect 1834 -1860 1894 -1800
rect 1834 -1926 1894 -1920
rect 474 -2034 534 -2028
rect -2224 -2058 -2164 -2052
rect -1968 -2082 160 -2046
rect -1908 -2106 160 -2082
rect 220 -2106 226 -2046
rect 2856 -2046 2922 -2040
rect -1968 -2148 -1908 -2142
rect -864 -2162 -804 -2156
rect -2400 -2278 -2280 -2266
rect -2400 -2350 -2388 -2278
rect -2292 -2350 -2280 -2278
rect -864 -2282 -804 -2222
rect -2400 -2362 -2280 -2350
rect -2224 -2342 -804 -2282
rect 474 -2286 534 -2094
rect 730 -2082 2856 -2046
rect 790 -2106 2856 -2082
rect 2916 -2106 2922 -2046
rect 2856 -2112 2922 -2106
rect 730 -2148 790 -2142
rect 2978 -2278 3098 -2266
rect -2224 -2534 -2164 -2342
rect 474 -2346 1894 -2286
rect 1834 -2406 1894 -2346
rect 2978 -2350 2990 -2278
rect 3086 -2350 3098 -2278
rect 2978 -2362 3098 -2350
rect 1834 -2472 1894 -2466
rect -1968 -2486 -1908 -2480
rect 730 -2486 790 -2480
rect 482 -2516 542 -2510
rect -1908 -2546 160 -2522
rect -1968 -2582 160 -2546
rect 220 -2582 226 -2522
rect 376 -2576 482 -2516
rect -2224 -2600 -2164 -2594
rect -864 -2706 -804 -2700
rect 376 -2706 436 -2576
rect 482 -2582 542 -2576
rect 790 -2546 2858 -2522
rect 730 -2582 2858 -2546
rect 2918 -2582 2924 -2522
rect -804 -2766 436 -2706
rect -864 -2772 -804 -2766
rect 280 -2822 400 -2810
rect 280 -2894 292 -2822
rect 388 -2894 400 -2822
rect 280 -2906 400 -2894
<< via2 >>
rect 292 370 388 442
rect -2388 -174 -2292 -102
rect 2990 -174 3086 -102
rect 292 -718 388 -646
rect -2388 -1262 -2292 -1190
rect 2990 -1262 3086 -1190
rect 292 -1806 388 -1734
rect -2388 -2350 -2292 -2278
rect 2990 -2350 3086 -2278
rect 292 -2894 388 -2822
<< metal3 >>
rect 280 442 400 454
rect 280 370 292 442
rect 388 370 400 442
rect 280 358 400 370
rect -2400 -102 -2280 -90
rect -2400 -174 -2388 -102
rect -2292 -174 -2280 -102
rect -2400 -186 -2280 -174
rect 2978 -102 3098 -90
rect 2978 -174 2990 -102
rect 3086 -174 3098 -102
rect 2978 -186 3098 -174
rect 280 -646 400 -634
rect 280 -718 292 -646
rect 388 -718 400 -646
rect 280 -730 400 -718
rect -2400 -1190 -2280 -1178
rect -2400 -1262 -2388 -1190
rect -2292 -1262 -2280 -1190
rect -2400 -1274 -2280 -1262
rect 2978 -1190 3098 -1178
rect 2978 -1262 2990 -1190
rect 3086 -1262 3098 -1190
rect 2978 -1274 3098 -1262
rect 280 -1734 400 -1722
rect 280 -1806 292 -1734
rect 388 -1806 400 -1734
rect 280 -1818 400 -1806
rect -2400 -2278 -2280 -2266
rect -2400 -2350 -2388 -2278
rect -2292 -2350 -2280 -2278
rect -2400 -2362 -2280 -2350
rect 2978 -2278 3098 -2266
rect 2978 -2350 2990 -2278
rect 3086 -2350 3098 -2278
rect 2978 -2362 3098 -2350
rect 280 -2822 400 -2810
rect 280 -2894 292 -2822
rect 388 -2894 400 -2822
rect 280 -2906 400 -2894
<< via3 >>
rect 292 370 388 442
rect -2388 -174 -2292 -102
rect 2990 -174 3086 -102
rect 292 -718 388 -646
rect -2388 -1262 -2292 -1190
rect 2990 -1262 3086 -1190
rect 292 -1806 388 -1734
rect -2388 -2350 -2292 -2278
rect 2990 -2350 3086 -2278
rect 292 -2894 388 -2822
<< metal4 >>
rect -2400 -102 -2280 454
rect -2400 -174 -2388 -102
rect -2292 -174 -2280 -102
rect -2400 -1190 -2280 -174
rect -2400 -1262 -2388 -1190
rect -2292 -1262 -2280 -1190
rect -2400 -2278 -2280 -1262
rect -2400 -2350 -2388 -2278
rect -2292 -2350 -2280 -2278
rect -2400 -2906 -2280 -2350
rect 280 442 400 454
rect 280 370 292 442
rect 388 370 400 442
rect 280 -646 400 370
rect 280 -718 292 -646
rect 388 -718 400 -646
rect 280 -1734 400 -718
rect 280 -1806 292 -1734
rect 388 -1806 400 -1734
rect 280 -2822 400 -1806
rect 280 -2894 292 -2822
rect 388 -2894 400 -2822
rect 280 -2906 400 -2894
rect 2978 -102 3098 454
rect 2978 -174 2990 -102
rect 3086 -174 3098 -102
rect 2978 -1190 3098 -174
rect 2978 -1262 2990 -1190
rect 3086 -1262 3098 -1190
rect 2978 -2278 3098 -1262
rect 2978 -2350 2990 -2278
rect 3086 -2350 3098 -2278
rect 2978 -2906 3098 -2350
<< labels >>
rlabel comment s -2242 -1226 -2242 -1226 4 dfxbp_1
rlabel comment s -2242 -2314 -2242 -2314 4 dfxbp_1
flabel metal1 s -2562 -691 -2509 -662 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel comment s -2584 -138 -2584 -138 2 tapvpwrvgnd_1
flabel metal1 s -2562 -702 -2509 -673 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s -2562 -1779 -2509 -1750 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel comment s -2584 -1226 -2584 -1226 2 tapvpwrvgnd_1
flabel metal1 s -2562 -1790 -2509 -1761 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s -2562 -2867 -2509 -2838 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel comment s -2584 -2314 -2584 -2314 2 tapvpwrvgnd_1
rlabel comment s 3282 -2314 3282 -2314 8 tapvpwrvgnd_1
flabel metal1 s 3207 -2867 3260 -2838 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 3207 -1790 3260 -1761 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel comment s 3282 -1226 3282 -1226 8 tapvpwrvgnd_1
flabel metal1 s 3207 -1779 3260 -1750 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 3207 -702 3260 -673 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel comment s 3282 -138 3282 -138 8 tapvpwrvgnd_1
flabel metal1 s 3207 -691 3260 -662 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 -2660 116 -2654 122 1 FreeSans 480 0 0 0 vin
port 1 n
flabel metal1 s 3210 -1244 3261 -1206 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 3210 -1246 3261 -1208 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 3210 -2332 3261 -2294 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 3210 -2334 3261 -2296 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s -2563 -2334 -2512 -2296 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s -2563 -2332 -2512 -2294 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s -2563 -1246 -2512 -1208 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s -2563 -1244 -2512 -1206 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s -2563 -158 -2512 -120 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 3210 -158 3261 -120 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal4 -2348 -374 -2344 -370 1 FreeSans 480 0 0 0 VSS
port 4 n ground bidirectional
flabel metal4 332 -378 342 -370 1 FreeSans 480 0 0 0 VDD
port 3 n power bidirectional
flabel metal2 1856 80 1866 88 1 FreeSans 480 0 0 0 vout
port 2 n
flabel metal1 -2213 -2331 -2179 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_5/VGND
flabel metal1 -2213 -2875 -2179 -2841 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_5/VPWR
flabel locali -557 -2652 -523 -2618 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_5/Q_N
flabel locali -1953 -2569 -1919 -2535 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_5/D
flabel locali -2213 -2569 -2179 -2535 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_5/CLK
flabel locali -852 -2433 -818 -2399 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_5/Q
flabel pwell -2213 -2331 -2179 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_5/VNB
flabel pwell -2196 -2314 -2196 -2314 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_5/VNB
flabel nwell -2213 -2875 -2179 -2841 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_5/VPB
flabel nwell -2196 -2858 -2196 -2858 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_5/VPB
rlabel comment -2242 -2314 -2242 -2314 2 sky130_fd_sc_hd__dfxbp_1_5/dfxbp_1
flabel metal1 -2213 -2331 -2179 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_4/VGND
flabel metal1 -2213 -1787 -2179 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_4/VPWR
flabel locali -557 -2010 -523 -1976 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_4/Q_N
flabel locali -1953 -2093 -1919 -2059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_4/D
flabel locali -2213 -2093 -2179 -2059 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_4/CLK
flabel locali -852 -2229 -818 -2195 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_4/Q
flabel pwell -2213 -2331 -2179 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_4/VNB
flabel pwell -2196 -2314 -2196 -2314 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_4/VNB
flabel nwell -2213 -1787 -2179 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_4/VPB
flabel nwell -2196 -1770 -2196 -1770 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_4/VPB
rlabel comment -2242 -2314 -2242 -2314 4 sky130_fd_sc_hd__dfxbp_1_4/dfxbp_1
flabel metal1 -2562 -2867 -2509 -2838 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_6/VPWR
flabel metal1 -2563 -2334 -2512 -2296 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_6/VGND
rlabel comment -2584 -2314 -2584 -2314 2 sky130_fd_sc_hd__tapvpwrvgnd_1_6/tapvpwrvgnd_1
flabel metal1 -2562 -1790 -2509 -1761 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_5/VPWR
flabel metal1 -2563 -2332 -2512 -2294 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_5/VGND
rlabel comment -2584 -2314 -2584 -2314 4 sky130_fd_sc_hd__tapvpwrvgnd_1_5/tapvpwrvgnd_1
flabel locali 179 -2501 213 -2467 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_5/Y
flabel locali 179 -2569 213 -2535 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_5/Y
flabel locali 179 -2637 213 -2603 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_5/Y
flabel locali -189 -2569 -155 -2535 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_5/A
flabel locali -97 -2569 -63 -2535 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_5/A
flabel locali -5 -2569 29 -2535 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_5/A
flabel locali 87 -2569 121 -2535 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_5/A
flabel nwell -189 -2875 -155 -2841 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_5/VPB
flabel pwell -189 -2331 -155 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_5/VNB
flabel metal1 -189 -2875 -155 -2841 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_5/VPWR
flabel metal1 -189 -2331 -155 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_5/VGND
rlabel comment -218 -2314 -218 -2314 2 sky130_fd_sc_hd__inv_4_5/inv_4
flabel locali 179 -2161 213 -2127 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_4/Y
flabel locali 179 -2093 213 -2059 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_4/Y
flabel locali 179 -2025 213 -1991 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_4/Y
flabel locali -189 -2093 -155 -2059 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_4/A
flabel locali -97 -2093 -63 -2059 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_4/A
flabel locali -5 -2093 29 -2059 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_4/A
flabel locali 87 -2093 121 -2059 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_4/A
flabel nwell -189 -1787 -155 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_4/VPB
flabel pwell -189 -2331 -155 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_4/VNB
flabel metal1 -189 -1787 -155 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_4/VPWR
flabel metal1 -189 -2331 -155 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_4/VGND
rlabel comment -218 -2314 -218 -2314 4 sky130_fd_sc_hd__inv_4_4/inv_4
flabel locali -330 -2637 -296 -2603 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_5/Y
flabel locali -330 -2569 -296 -2535 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_5/Y
flabel locali -422 -2569 -388 -2535 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_5/A
flabel nwell -465 -2875 -431 -2841 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_5/VPB
flabel pwell -465 -2331 -431 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_5/VNB
flabel metal1 -465 -2331 -431 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_5/VGND
flabel metal1 -465 -2875 -431 -2841 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_5/VPWR
rlabel comment -494 -2314 -494 -2314 2 sky130_fd_sc_hd__inv_1_5/inv_1
flabel locali -330 -2025 -296 -1991 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_4/Y
flabel locali -330 -2093 -296 -2059 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_4/Y
flabel locali -422 -2093 -388 -2059 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_4/A
flabel nwell -465 -1787 -431 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_4/VPB
flabel pwell -465 -2331 -431 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_4/VNB
flabel metal1 -465 -2331 -431 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_4/VGND
flabel metal1 -465 -1787 -431 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_4/VPWR
rlabel comment -494 -2314 -494 -2314 4 sky130_fd_sc_hd__inv_1_4/inv_1
flabel metal1 485 -2331 519 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_10/VGND
flabel metal1 485 -2875 519 -2841 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_10/VPWR
flabel locali 2141 -2652 2175 -2618 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_10/Q_N
flabel locali 745 -2569 779 -2535 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_10/D
flabel locali 485 -2569 519 -2535 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_10/CLK
flabel locali 1846 -2433 1880 -2399 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_10/Q
flabel pwell 485 -2331 519 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_10/VNB
flabel pwell 502 -2314 502 -2314 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_10/VNB
flabel nwell 485 -2875 519 -2841 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_10/VPB
flabel nwell 502 -2858 502 -2858 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_10/VPB
rlabel comment 456 -2314 456 -2314 2 sky130_fd_sc_hd__dfxbp_1_10/dfxbp_1
flabel metal1 485 -2331 519 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_9/VGND
flabel metal1 485 -1787 519 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_9/VPWR
flabel locali 2141 -2010 2175 -1976 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_9/Q_N
flabel locali 745 -2093 779 -2059 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_9/D
flabel locali 485 -2093 519 -2059 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_9/CLK
flabel locali 1846 -2229 1880 -2195 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_9/Q
flabel pwell 485 -2331 519 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_9/VNB
flabel pwell 502 -2314 502 -2314 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_9/VNB
flabel nwell 485 -1787 519 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_9/VPB
flabel nwell 502 -1770 502 -1770 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_9/VPB
rlabel comment 456 -2314 456 -2314 4 sky130_fd_sc_hd__dfxbp_1_9/dfxbp_1
flabel locali 2877 -2501 2911 -2467 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_10/Y
flabel locali 2877 -2569 2911 -2535 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_10/Y
flabel locali 2877 -2637 2911 -2603 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_10/Y
flabel locali 2509 -2569 2543 -2535 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_10/A
flabel locali 2601 -2569 2635 -2535 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_10/A
flabel locali 2693 -2569 2727 -2535 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_10/A
flabel locali 2785 -2569 2819 -2535 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_10/A
flabel nwell 2509 -2875 2543 -2841 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_10/VPB
flabel pwell 2509 -2331 2543 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_10/VNB
flabel metal1 2509 -2875 2543 -2841 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_10/VPWR
flabel metal1 2509 -2331 2543 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_10/VGND
rlabel comment 2480 -2314 2480 -2314 2 sky130_fd_sc_hd__inv_4_10/inv_4
flabel locali 2877 -2161 2911 -2127 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_9/Y
flabel locali 2877 -2093 2911 -2059 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_9/Y
flabel locali 2877 -2025 2911 -1991 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_9/Y
flabel locali 2509 -2093 2543 -2059 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_9/A
flabel locali 2601 -2093 2635 -2059 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_9/A
flabel locali 2693 -2093 2727 -2059 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_9/A
flabel locali 2785 -2093 2819 -2059 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_9/A
flabel nwell 2509 -1787 2543 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_9/VPB
flabel pwell 2509 -2331 2543 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_9/VNB
flabel metal1 2509 -1787 2543 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_9/VPWR
flabel metal1 2509 -2331 2543 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_9/VGND
rlabel comment 2480 -2314 2480 -2314 4 sky130_fd_sc_hd__inv_4_9/inv_4
flabel locali 2368 -2637 2402 -2603 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_10/Y
flabel locali 2368 -2569 2402 -2535 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_10/Y
flabel locali 2276 -2569 2310 -2535 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_10/A
flabel nwell 2233 -2875 2267 -2841 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_10/VPB
flabel pwell 2233 -2331 2267 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_10/VNB
flabel metal1 2233 -2331 2267 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_10/VGND
flabel metal1 2233 -2875 2267 -2841 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_10/VPWR
rlabel comment 2204 -2314 2204 -2314 2 sky130_fd_sc_hd__inv_1_10/inv_1
flabel locali 2368 -2025 2402 -1991 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_9/Y
flabel locali 2368 -2093 2402 -2059 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_9/Y
flabel locali 2276 -2093 2310 -2059 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_9/A
flabel nwell 2233 -1787 2267 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_9/VPB
flabel pwell 2233 -2331 2267 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_9/VNB
flabel metal1 2233 -2331 2267 -2297 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_9/VGND
flabel metal1 2233 -1787 2267 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_9/VPWR
rlabel comment 2204 -2314 2204 -2314 4 sky130_fd_sc_hd__inv_1_9/inv_1
flabel metal1 3207 -2867 3260 -2838 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_7/VPWR
flabel metal1 3210 -2334 3261 -2296 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_7/VGND
rlabel comment 3282 -2314 3282 -2314 8 sky130_fd_sc_hd__tapvpwrvgnd_1_7/tapvpwrvgnd_1
flabel metal1 3207 -1790 3260 -1761 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_8/VPWR
flabel metal1 3210 -2332 3261 -2294 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_8/VGND
rlabel comment 3282 -2314 3282 -2314 6 sky130_fd_sc_hd__tapvpwrvgnd_1_8/tapvpwrvgnd_1
flabel metal1 -2213 -1243 -2179 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/VGND
flabel metal1 -2213 -1787 -2179 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/VPWR
flabel locali -557 -1564 -523 -1530 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/Q_N
flabel locali -1953 -1481 -1919 -1447 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/D
flabel locali -2213 -1481 -2179 -1447 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/CLK
flabel locali -852 -1345 -818 -1311 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/Q
flabel pwell -2213 -1243 -2179 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/VNB
flabel pwell -2196 -1226 -2196 -1226 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/VNB
flabel nwell -2213 -1787 -2179 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/VPB
flabel nwell -2196 -1770 -2196 -1770 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2/VPB
rlabel comment -2242 -1226 -2242 -1226 2 sky130_fd_sc_hd__dfxbp_1_2/dfxbp_1
flabel metal1 -2562 -1779 -2509 -1750 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_4/VPWR
flabel metal1 -2563 -1246 -2512 -1208 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_4/VGND
rlabel comment -2584 -1226 -2584 -1226 2 sky130_fd_sc_hd__tapvpwrvgnd_1_4/tapvpwrvgnd_1
flabel locali 179 -1413 213 -1379 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_2/Y
flabel locali 179 -1481 213 -1447 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_2/Y
flabel locali 179 -1549 213 -1515 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_2/Y
flabel locali -189 -1481 -155 -1447 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_2/A
flabel locali -97 -1481 -63 -1447 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_2/A
flabel locali -5 -1481 29 -1447 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_2/A
flabel locali 87 -1481 121 -1447 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_2/A
flabel nwell -189 -1787 -155 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_2/VPB
flabel pwell -189 -1243 -155 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_2/VNB
flabel metal1 -189 -1787 -155 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_2/VPWR
flabel metal1 -189 -1243 -155 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_2/VGND
rlabel comment -218 -1226 -218 -1226 2 sky130_fd_sc_hd__inv_4_2/inv_4
flabel locali -330 -1549 -296 -1515 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_2/Y
flabel locali -330 -1481 -296 -1447 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_2/Y
flabel locali -422 -1481 -388 -1447 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_2/A
flabel nwell -465 -1787 -431 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_2/VPB
flabel pwell -465 -1243 -431 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_2/VNB
flabel metal1 -465 -1243 -431 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_2/VGND
flabel metal1 -465 -1787 -431 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_2/VPWR
rlabel comment -494 -1226 -494 -1226 2 sky130_fd_sc_hd__inv_1_2/inv_1
flabel metal1 485 -1243 519 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_8/VGND
flabel metal1 485 -1787 519 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_8/VPWR
flabel locali 2141 -1564 2175 -1530 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_8/Q_N
flabel locali 745 -1481 779 -1447 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_8/D
flabel locali 485 -1481 519 -1447 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_8/CLK
flabel locali 1846 -1345 1880 -1311 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_8/Q
flabel pwell 485 -1243 519 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_8/VNB
flabel pwell 502 -1226 502 -1226 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_8/VNB
flabel nwell 485 -1787 519 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_8/VPB
flabel nwell 502 -1770 502 -1770 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_8/VPB
rlabel comment 456 -1226 456 -1226 2 sky130_fd_sc_hd__dfxbp_1_8/dfxbp_1
flabel locali 2877 -1413 2911 -1379 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_8/Y
flabel locali 2877 -1481 2911 -1447 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_8/Y
flabel locali 2877 -1549 2911 -1515 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_8/Y
flabel locali 2509 -1481 2543 -1447 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_8/A
flabel locali 2601 -1481 2635 -1447 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_8/A
flabel locali 2693 -1481 2727 -1447 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_8/A
flabel locali 2785 -1481 2819 -1447 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_8/A
flabel nwell 2509 -1787 2543 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_8/VPB
flabel pwell 2509 -1243 2543 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_8/VNB
flabel metal1 2509 -1787 2543 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_8/VPWR
flabel metal1 2509 -1243 2543 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_8/VGND
rlabel comment 2480 -1226 2480 -1226 2 sky130_fd_sc_hd__inv_4_8/inv_4
flabel locali 2368 -1549 2402 -1515 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_8/Y
flabel locali 2368 -1481 2402 -1447 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_8/Y
flabel locali 2276 -1481 2310 -1447 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_8/A
flabel nwell 2233 -1787 2267 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_8/VPB
flabel pwell 2233 -1243 2267 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_8/VNB
flabel metal1 2233 -1243 2267 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_8/VGND
flabel metal1 2233 -1787 2267 -1753 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_8/VPWR
rlabel comment 2204 -1226 2204 -1226 2 sky130_fd_sc_hd__inv_1_8/inv_1
flabel metal1 3207 -1779 3260 -1750 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_9/VPWR
flabel metal1 3210 -1246 3261 -1208 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_9/VGND
rlabel comment 3282 -1226 3282 -1226 8 sky130_fd_sc_hd__tapvpwrvgnd_1_9/tapvpwrvgnd_1
flabel metal1 -2213 -1243 -2179 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/VGND
flabel metal1 -2213 -699 -2179 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/VPWR
flabel locali -557 -922 -523 -888 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/Q_N
flabel locali -1953 -1005 -1919 -971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/D
flabel locali -2213 -1005 -2179 -971 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/CLK
flabel locali -852 -1141 -818 -1107 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/Q
flabel pwell -2213 -1243 -2179 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/VNB
flabel pwell -2196 -1226 -2196 -1226 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/VNB
flabel nwell -2213 -699 -2179 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/VPB
flabel nwell -2196 -682 -2196 -682 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3/VPB
rlabel comment -2242 -1226 -2242 -1226 4 sky130_fd_sc_hd__dfxbp_1_3/dfxbp_1
flabel metal1 -2562 -702 -2509 -673 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_3/VPWR
flabel metal1 -2563 -1244 -2512 -1206 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_3/VGND
rlabel comment -2584 -1226 -2584 -1226 4 sky130_fd_sc_hd__tapvpwrvgnd_1_3/tapvpwrvgnd_1
flabel locali 179 -1073 213 -1039 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_3/Y
flabel locali 179 -1005 213 -971 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_3/Y
flabel locali 179 -937 213 -903 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_3/Y
flabel locali -189 -1005 -155 -971 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_3/A
flabel locali -97 -1005 -63 -971 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_3/A
flabel locali -5 -1005 29 -971 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_3/A
flabel locali 87 -1005 121 -971 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_3/A
flabel nwell -189 -699 -155 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_3/VPB
flabel pwell -189 -1243 -155 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_3/VNB
flabel metal1 -189 -699 -155 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_3/VPWR
flabel metal1 -189 -1243 -155 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_3/VGND
rlabel comment -218 -1226 -218 -1226 4 sky130_fd_sc_hd__inv_4_3/inv_4
flabel locali -330 -937 -296 -903 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_3/Y
flabel locali -330 -1005 -296 -971 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_3/Y
flabel locali -422 -1005 -388 -971 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_3/A
flabel nwell -465 -699 -431 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_3/VPB
flabel pwell -465 -1243 -431 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_3/VNB
flabel metal1 -465 -1243 -431 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_3/VGND
flabel metal1 -465 -699 -431 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_3/VPWR
rlabel comment -494 -1226 -494 -1226 4 sky130_fd_sc_hd__inv_1_3/inv_1
flabel metal1 485 -1243 519 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_7/VGND
flabel metal1 485 -699 519 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_7/VPWR
flabel locali 2141 -922 2175 -888 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_7/Q_N
flabel locali 745 -1005 779 -971 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_7/D
flabel locali 485 -1005 519 -971 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_7/CLK
flabel locali 1846 -1141 1880 -1107 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_7/Q
flabel pwell 485 -1243 519 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_7/VNB
flabel pwell 502 -1226 502 -1226 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_7/VNB
flabel nwell 485 -699 519 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_7/VPB
flabel nwell 502 -682 502 -682 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_7/VPB
rlabel comment 456 -1226 456 -1226 4 sky130_fd_sc_hd__dfxbp_1_7/dfxbp_1
flabel locali 2877 -1073 2911 -1039 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_7/Y
flabel locali 2877 -1005 2911 -971 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_7/Y
flabel locali 2877 -937 2911 -903 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_7/Y
flabel locali 2509 -1005 2543 -971 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_7/A
flabel locali 2601 -1005 2635 -971 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_7/A
flabel locali 2693 -1005 2727 -971 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_7/A
flabel locali 2785 -1005 2819 -971 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_7/A
flabel nwell 2509 -699 2543 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_7/VPB
flabel pwell 2509 -1243 2543 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_7/VNB
flabel metal1 2509 -699 2543 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_7/VPWR
flabel metal1 2509 -1243 2543 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_7/VGND
rlabel comment 2480 -1226 2480 -1226 4 sky130_fd_sc_hd__inv_4_7/inv_4
flabel locali 2368 -937 2402 -903 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_7/Y
flabel locali 2368 -1005 2402 -971 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_7/Y
flabel locali 2276 -1005 2310 -971 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_7/A
flabel nwell 2233 -699 2267 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_7/VPB
flabel pwell 2233 -1243 2267 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_7/VNB
flabel metal1 2233 -1243 2267 -1209 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_7/VGND
flabel metal1 2233 -699 2267 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_7/VPWR
rlabel comment 2204 -1226 2204 -1226 4 sky130_fd_sc_hd__inv_1_7/inv_1
flabel metal1 3207 -702 3260 -673 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_10/VPWR
flabel metal1 3210 -1244 3261 -1206 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_10/VGND
rlabel comment 3282 -1226 3282 -1226 6 sky130_fd_sc_hd__tapvpwrvgnd_1_10/tapvpwrvgnd_1
flabel metal1 -2213 -155 -2179 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VGND
flabel metal1 -2213 -699 -2179 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VPWR
flabel locali -557 -476 -523 -442 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/Q_N
flabel locali -1953 -393 -1919 -359 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/D
flabel locali -2213 -393 -2179 -359 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/CLK
flabel locali -852 -257 -818 -223 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/Q
flabel pwell -2213 -155 -2179 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VNB
flabel pwell -2196 -138 -2196 -138 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VNB
flabel nwell -2213 -699 -2179 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VPB
flabel nwell -2196 -682 -2196 -682 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1/VPB
rlabel comment -2242 -138 -2242 -138 2 sky130_fd_sc_hd__dfxbp_1_1/dfxbp_1
flabel metal1 -2562 -691 -2509 -662 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_2/VPWR
flabel metal1 -2563 -158 -2512 -120 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_2/VGND
rlabel comment -2584 -138 -2584 -138 2 sky130_fd_sc_hd__tapvpwrvgnd_1_2/tapvpwrvgnd_1
flabel locali 179 -325 213 -291 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_1/Y
flabel locali 179 -393 213 -359 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_1/Y
flabel locali 179 -461 213 -427 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_1/Y
flabel locali -189 -393 -155 -359 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_1/A
flabel locali -97 -393 -63 -359 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_1/A
flabel locali -5 -393 29 -359 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_1/A
flabel locali 87 -393 121 -359 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_1/A
flabel nwell -189 -699 -155 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_1/VPB
flabel pwell -189 -155 -155 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_1/VNB
flabel metal1 -189 -699 -155 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_1/VPWR
flabel metal1 -189 -155 -155 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_1/VGND
rlabel comment -218 -138 -218 -138 2 sky130_fd_sc_hd__inv_4_1/inv_4
flabel locali -330 -461 -296 -427 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/Y
flabel locali -330 -393 -296 -359 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/Y
flabel locali -422 -393 -388 -359 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/A
flabel nwell -465 -699 -431 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VPB
flabel pwell -465 -155 -431 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VNB
flabel metal1 -465 -155 -431 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VGND
flabel metal1 -465 -699 -431 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VPWR
rlabel comment -494 -138 -494 -138 2 sky130_fd_sc_hd__inv_1_1/inv_1
flabel metal1 485 -155 519 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_6/VGND
flabel metal1 485 -699 519 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_6/VPWR
flabel locali 2141 -476 2175 -442 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_6/Q_N
flabel locali 745 -393 779 -359 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_6/D
flabel locali 485 -393 519 -359 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_6/CLK
flabel locali 1846 -257 1880 -223 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_6/Q
flabel pwell 485 -155 519 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_6/VNB
flabel pwell 502 -138 502 -138 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_6/VNB
flabel nwell 485 -699 519 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_6/VPB
flabel nwell 502 -682 502 -682 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_6/VPB
rlabel comment 456 -138 456 -138 2 sky130_fd_sc_hd__dfxbp_1_6/dfxbp_1
flabel locali 2877 -325 2911 -291 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_6/Y
flabel locali 2877 -393 2911 -359 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_6/Y
flabel locali 2877 -461 2911 -427 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_6/Y
flabel locali 2509 -393 2543 -359 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_6/A
flabel locali 2601 -393 2635 -359 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_6/A
flabel locali 2693 -393 2727 -359 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_6/A
flabel locali 2785 -393 2819 -359 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_6/A
flabel nwell 2509 -699 2543 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_6/VPB
flabel pwell 2509 -155 2543 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_6/VNB
flabel metal1 2509 -699 2543 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_6/VPWR
flabel metal1 2509 -155 2543 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_6/VGND
rlabel comment 2480 -138 2480 -138 2 sky130_fd_sc_hd__inv_4_6/inv_4
flabel locali 2368 -461 2402 -427 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_6/Y
flabel locali 2368 -393 2402 -359 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_6/Y
flabel locali 2276 -393 2310 -359 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_6/A
flabel nwell 2233 -699 2267 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_6/VPB
flabel pwell 2233 -155 2267 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_6/VNB
flabel metal1 2233 -155 2267 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_6/VGND
flabel metal1 2233 -699 2267 -665 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_6/VPWR
rlabel comment 2204 -138 2204 -138 2 sky130_fd_sc_hd__inv_1_6/inv_1
flabel metal1 3207 -691 3260 -662 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_11/VPWR
flabel metal1 3210 -158 3261 -120 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_11/VGND
rlabel comment 3282 -138 3282 -138 8 sky130_fd_sc_hd__tapvpwrvgnd_1_11/tapvpwrvgnd_1
flabel metal1 -2213 -155 -2179 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VGND
flabel metal1 -2213 389 -2179 423 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VPWR
flabel locali -557 166 -523 200 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/Q_N
flabel locali -1953 83 -1919 117 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/D
flabel locali -2213 83 -2179 117 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/CLK
flabel locali -852 -53 -818 -19 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/Q
flabel pwell -2213 -155 -2179 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VNB
flabel pwell -2196 -138 -2196 -138 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VNB
flabel nwell -2213 389 -2179 423 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VPB
flabel nwell -2196 406 -2196 406 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0/VPB
rlabel comment -2242 -138 -2242 -138 4 sky130_fd_sc_hd__dfxbp_1_0/dfxbp_1
flabel metal1 -2562 386 -2509 415 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VPWR
flabel metal1 -2563 -156 -2512 -118 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VGND
rlabel comment -2584 -138 -2584 -138 4 sky130_fd_sc_hd__tapvpwrvgnd_1_1/tapvpwrvgnd_1
flabel locali 179 15 213 49 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/Y
flabel locali 179 83 213 117 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/Y
flabel locali 179 151 213 185 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/Y
flabel locali -189 83 -155 117 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/A
flabel locali -97 83 -63 117 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/A
flabel locali -5 83 29 117 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/A
flabel locali 87 83 121 117 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/A
flabel nwell -189 389 -155 423 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0/VPB
flabel pwell -189 -155 -155 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0/VNB
flabel metal1 -189 389 -155 423 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0/VPWR
flabel metal1 -189 -155 -155 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0/VGND
rlabel comment -218 -138 -218 -138 4 sky130_fd_sc_hd__inv_4_0/inv_4
flabel locali -330 151 -296 185 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali -330 83 -296 117 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali -422 83 -388 117 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/A
flabel nwell -465 389 -431 423 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -465 -155 -431 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -465 -155 -431 -121 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -465 389 -431 423 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -494 -138 -494 -138 4 sky130_fd_sc_hd__inv_1_0/inv_1
flabel metal1 338 386 391 415 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VPWR
flabel metal1 337 -156 388 -118 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VGND
rlabel comment 316 -138 316 -138 4 sky130_fd_sc_hd__tapvpwrvgnd_1_0/tapvpwrvgnd_1
flabel metal1 3207 386 3260 415 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_12/VPWR
flabel metal1 3210 -156 3261 -118 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_12/VGND
rlabel comment 3282 -138 3282 -138 6 sky130_fd_sc_hd__tapvpwrvgnd_1_12/tapvpwrvgnd_1
<< end >>
