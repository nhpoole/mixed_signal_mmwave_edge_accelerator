magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -2699 -1460 2699 1460
<< nwell >>
rect -1439 -200 1439 200
<< pmos >>
rect -1345 -100 -945 100
rect -887 -100 -487 100
rect -429 -100 -29 100
rect 29 -100 429 100
rect 487 -100 887 100
rect 945 -100 1345 100
<< pdiff >>
rect -1403 85 -1345 100
rect -1403 51 -1391 85
rect -1357 51 -1345 85
rect -1403 17 -1345 51
rect -1403 -17 -1391 17
rect -1357 -17 -1345 17
rect -1403 -51 -1345 -17
rect -1403 -85 -1391 -51
rect -1357 -85 -1345 -51
rect -1403 -100 -1345 -85
rect -945 85 -887 100
rect -945 51 -933 85
rect -899 51 -887 85
rect -945 17 -887 51
rect -945 -17 -933 17
rect -899 -17 -887 17
rect -945 -51 -887 -17
rect -945 -85 -933 -51
rect -899 -85 -887 -51
rect -945 -100 -887 -85
rect -487 85 -429 100
rect -487 51 -475 85
rect -441 51 -429 85
rect -487 17 -429 51
rect -487 -17 -475 17
rect -441 -17 -429 17
rect -487 -51 -429 -17
rect -487 -85 -475 -51
rect -441 -85 -429 -51
rect -487 -100 -429 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 429 85 487 100
rect 429 51 441 85
rect 475 51 487 85
rect 429 17 487 51
rect 429 -17 441 17
rect 475 -17 487 17
rect 429 -51 487 -17
rect 429 -85 441 -51
rect 475 -85 487 -51
rect 429 -100 487 -85
rect 887 85 945 100
rect 887 51 899 85
rect 933 51 945 85
rect 887 17 945 51
rect 887 -17 899 17
rect 933 -17 945 17
rect 887 -51 945 -17
rect 887 -85 899 -51
rect 933 -85 945 -51
rect 887 -100 945 -85
rect 1345 85 1403 100
rect 1345 51 1357 85
rect 1391 51 1403 85
rect 1345 17 1403 51
rect 1345 -17 1357 17
rect 1391 -17 1403 17
rect 1345 -51 1403 -17
rect 1345 -85 1357 -51
rect 1391 -85 1403 -51
rect 1345 -100 1403 -85
<< pdiffc >>
rect -1391 51 -1357 85
rect -1391 -17 -1357 17
rect -1391 -85 -1357 -51
rect -933 51 -899 85
rect -933 -17 -899 17
rect -933 -85 -899 -51
rect -475 51 -441 85
rect -475 -17 -441 17
rect -475 -85 -441 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 441 51 475 85
rect 441 -17 475 17
rect 441 -85 475 -51
rect 899 51 933 85
rect 899 -17 933 17
rect 899 -85 933 -51
rect 1357 51 1391 85
rect 1357 -17 1391 17
rect 1357 -85 1391 -51
<< poly >>
rect -1271 181 -1019 197
rect -1271 164 -1230 181
rect -1345 147 -1230 164
rect -1196 147 -1162 181
rect -1128 147 -1094 181
rect -1060 164 -1019 181
rect -813 181 -561 197
rect -813 164 -772 181
rect -1060 147 -945 164
rect -1345 100 -945 147
rect -887 147 -772 164
rect -738 147 -704 181
rect -670 147 -636 181
rect -602 164 -561 181
rect -355 181 -103 197
rect -355 164 -314 181
rect -602 147 -487 164
rect -887 100 -487 147
rect -429 147 -314 164
rect -280 147 -246 181
rect -212 147 -178 181
rect -144 164 -103 181
rect 103 181 355 197
rect 103 164 144 181
rect -144 147 -29 164
rect -429 100 -29 147
rect 29 147 144 164
rect 178 147 212 181
rect 246 147 280 181
rect 314 164 355 181
rect 561 181 813 197
rect 561 164 602 181
rect 314 147 429 164
rect 29 100 429 147
rect 487 147 602 164
rect 636 147 670 181
rect 704 147 738 181
rect 772 164 813 181
rect 1019 181 1271 197
rect 1019 164 1060 181
rect 772 147 887 164
rect 487 100 887 147
rect 945 147 1060 164
rect 1094 147 1128 181
rect 1162 147 1196 181
rect 1230 164 1271 181
rect 1230 147 1345 164
rect 945 100 1345 147
rect -1345 -147 -945 -100
rect -1345 -164 -1230 -147
rect -1271 -181 -1230 -164
rect -1196 -181 -1162 -147
rect -1128 -181 -1094 -147
rect -1060 -164 -945 -147
rect -887 -147 -487 -100
rect -887 -164 -772 -147
rect -1060 -181 -1019 -164
rect -1271 -197 -1019 -181
rect -813 -181 -772 -164
rect -738 -181 -704 -147
rect -670 -181 -636 -147
rect -602 -164 -487 -147
rect -429 -147 -29 -100
rect -429 -164 -314 -147
rect -602 -181 -561 -164
rect -813 -197 -561 -181
rect -355 -181 -314 -164
rect -280 -181 -246 -147
rect -212 -181 -178 -147
rect -144 -164 -29 -147
rect 29 -147 429 -100
rect 29 -164 144 -147
rect -144 -181 -103 -164
rect -355 -197 -103 -181
rect 103 -181 144 -164
rect 178 -181 212 -147
rect 246 -181 280 -147
rect 314 -164 429 -147
rect 487 -147 887 -100
rect 487 -164 602 -147
rect 314 -181 355 -164
rect 103 -197 355 -181
rect 561 -181 602 -164
rect 636 -181 670 -147
rect 704 -181 738 -147
rect 772 -164 887 -147
rect 945 -147 1345 -100
rect 945 -164 1060 -147
rect 772 -181 813 -164
rect 561 -197 813 -181
rect 1019 -181 1060 -164
rect 1094 -181 1128 -147
rect 1162 -181 1196 -147
rect 1230 -164 1345 -147
rect 1230 -181 1271 -164
rect 1019 -197 1271 -181
<< polycont >>
rect -1230 147 -1196 181
rect -1162 147 -1128 181
rect -1094 147 -1060 181
rect -772 147 -738 181
rect -704 147 -670 181
rect -636 147 -602 181
rect -314 147 -280 181
rect -246 147 -212 181
rect -178 147 -144 181
rect 144 147 178 181
rect 212 147 246 181
rect 280 147 314 181
rect 602 147 636 181
rect 670 147 704 181
rect 738 147 772 181
rect 1060 147 1094 181
rect 1128 147 1162 181
rect 1196 147 1230 181
rect -1230 -181 -1196 -147
rect -1162 -181 -1128 -147
rect -1094 -181 -1060 -147
rect -772 -181 -738 -147
rect -704 -181 -670 -147
rect -636 -181 -602 -147
rect -314 -181 -280 -147
rect -246 -181 -212 -147
rect -178 -181 -144 -147
rect 144 -181 178 -147
rect 212 -181 246 -147
rect 280 -181 314 -147
rect 602 -181 636 -147
rect 670 -181 704 -147
rect 738 -181 772 -147
rect 1060 -181 1094 -147
rect 1128 -181 1162 -147
rect 1196 -181 1230 -147
<< locali >>
rect -1271 147 -1234 181
rect -1196 147 -1162 181
rect -1128 147 -1094 181
rect -1056 147 -1019 181
rect -813 147 -776 181
rect -738 147 -704 181
rect -670 147 -636 181
rect -598 147 -561 181
rect -355 147 -318 181
rect -280 147 -246 181
rect -212 147 -178 181
rect -140 147 -103 181
rect 103 147 140 181
rect 178 147 212 181
rect 246 147 280 181
rect 318 147 355 181
rect 561 147 598 181
rect 636 147 670 181
rect 704 147 738 181
rect 776 147 813 181
rect 1019 147 1056 181
rect 1094 147 1128 181
rect 1162 147 1196 181
rect 1234 147 1271 181
rect -1391 85 -1357 104
rect -1391 17 -1357 19
rect -1391 -19 -1357 -17
rect -1391 -104 -1357 -85
rect -933 85 -899 104
rect -933 17 -899 19
rect -933 -19 -899 -17
rect -933 -104 -899 -85
rect -475 85 -441 104
rect -475 17 -441 19
rect -475 -19 -441 -17
rect -475 -104 -441 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 441 85 475 104
rect 441 17 475 19
rect 441 -19 475 -17
rect 441 -104 475 -85
rect 899 85 933 104
rect 899 17 933 19
rect 899 -19 933 -17
rect 899 -104 933 -85
rect 1357 85 1391 104
rect 1357 17 1391 19
rect 1357 -19 1391 -17
rect 1357 -104 1391 -85
rect -1271 -181 -1234 -147
rect -1196 -181 -1162 -147
rect -1128 -181 -1094 -147
rect -1056 -181 -1019 -147
rect -813 -181 -776 -147
rect -738 -181 -704 -147
rect -670 -181 -636 -147
rect -598 -181 -561 -147
rect -355 -181 -318 -147
rect -280 -181 -246 -147
rect -212 -181 -178 -147
rect -140 -181 -103 -147
rect 103 -181 140 -147
rect 178 -181 212 -147
rect 246 -181 280 -147
rect 318 -181 355 -147
rect 561 -181 598 -147
rect 636 -181 670 -147
rect 704 -181 738 -147
rect 776 -181 813 -147
rect 1019 -181 1056 -147
rect 1094 -181 1128 -147
rect 1162 -181 1196 -147
rect 1234 -181 1271 -147
<< viali >>
rect -1234 147 -1230 181
rect -1230 147 -1200 181
rect -1162 147 -1128 181
rect -1090 147 -1060 181
rect -1060 147 -1056 181
rect -776 147 -772 181
rect -772 147 -742 181
rect -704 147 -670 181
rect -632 147 -602 181
rect -602 147 -598 181
rect -318 147 -314 181
rect -314 147 -284 181
rect -246 147 -212 181
rect -174 147 -144 181
rect -144 147 -140 181
rect 140 147 144 181
rect 144 147 174 181
rect 212 147 246 181
rect 284 147 314 181
rect 314 147 318 181
rect 598 147 602 181
rect 602 147 632 181
rect 670 147 704 181
rect 742 147 772 181
rect 772 147 776 181
rect 1056 147 1060 181
rect 1060 147 1090 181
rect 1128 147 1162 181
rect 1200 147 1230 181
rect 1230 147 1234 181
rect -1391 51 -1357 53
rect -1391 19 -1357 51
rect -1391 -51 -1357 -19
rect -1391 -53 -1357 -51
rect -933 51 -899 53
rect -933 19 -899 51
rect -933 -51 -899 -19
rect -933 -53 -899 -51
rect -475 51 -441 53
rect -475 19 -441 51
rect -475 -51 -441 -19
rect -475 -53 -441 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 441 51 475 53
rect 441 19 475 51
rect 441 -51 475 -19
rect 441 -53 475 -51
rect 899 51 933 53
rect 899 19 933 51
rect 899 -51 933 -19
rect 899 -53 933 -51
rect 1357 51 1391 53
rect 1357 19 1391 51
rect 1357 -51 1391 -19
rect 1357 -53 1391 -51
rect -1234 -181 -1230 -147
rect -1230 -181 -1200 -147
rect -1162 -181 -1128 -147
rect -1090 -181 -1060 -147
rect -1060 -181 -1056 -147
rect -776 -181 -772 -147
rect -772 -181 -742 -147
rect -704 -181 -670 -147
rect -632 -181 -602 -147
rect -602 -181 -598 -147
rect -318 -181 -314 -147
rect -314 -181 -284 -147
rect -246 -181 -212 -147
rect -174 -181 -144 -147
rect -144 -181 -140 -147
rect 140 -181 144 -147
rect 144 -181 174 -147
rect 212 -181 246 -147
rect 284 -181 314 -147
rect 314 -181 318 -147
rect 598 -181 602 -147
rect 602 -181 632 -147
rect 670 -181 704 -147
rect 742 -181 772 -147
rect 772 -181 776 -147
rect 1056 -181 1060 -147
rect 1060 -181 1090 -147
rect 1128 -181 1162 -147
rect 1200 -181 1230 -147
rect 1230 -181 1234 -147
<< metal1 >>
rect -1249 181 -1041 187
rect -1249 147 -1234 181
rect -1200 147 -1162 181
rect -1128 147 -1090 181
rect -1056 147 -1041 181
rect -1249 141 -1041 147
rect -791 181 -583 187
rect -791 147 -776 181
rect -742 147 -704 181
rect -670 147 -632 181
rect -598 147 -583 181
rect -791 141 -583 147
rect -333 181 -125 187
rect -333 147 -318 181
rect -284 147 -246 181
rect -212 147 -174 181
rect -140 147 -125 181
rect -333 141 -125 147
rect 125 181 333 187
rect 125 147 140 181
rect 174 147 212 181
rect 246 147 284 181
rect 318 147 333 181
rect 125 141 333 147
rect 583 181 791 187
rect 583 147 598 181
rect 632 147 670 181
rect 704 147 742 181
rect 776 147 791 181
rect 583 141 791 147
rect 1041 181 1249 187
rect 1041 147 1056 181
rect 1090 147 1128 181
rect 1162 147 1200 181
rect 1234 147 1249 181
rect 1041 141 1249 147
rect -1397 53 -1351 100
rect -1397 19 -1391 53
rect -1357 19 -1351 53
rect -1397 -19 -1351 19
rect -1397 -53 -1391 -19
rect -1357 -53 -1351 -19
rect -1397 -100 -1351 -53
rect -939 53 -893 100
rect -939 19 -933 53
rect -899 19 -893 53
rect -939 -19 -893 19
rect -939 -53 -933 -19
rect -899 -53 -893 -19
rect -939 -100 -893 -53
rect -481 53 -435 100
rect -481 19 -475 53
rect -441 19 -435 53
rect -481 -19 -435 19
rect -481 -53 -475 -19
rect -441 -53 -435 -19
rect -481 -100 -435 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 435 53 481 100
rect 435 19 441 53
rect 475 19 481 53
rect 435 -19 481 19
rect 435 -53 441 -19
rect 475 -53 481 -19
rect 435 -100 481 -53
rect 893 53 939 100
rect 893 19 899 53
rect 933 19 939 53
rect 893 -19 939 19
rect 893 -53 899 -19
rect 933 -53 939 -19
rect 893 -100 939 -53
rect 1351 53 1397 100
rect 1351 19 1357 53
rect 1391 19 1397 53
rect 1351 -19 1397 19
rect 1351 -53 1357 -19
rect 1391 -53 1397 -19
rect 1351 -100 1397 -53
rect -1249 -147 -1041 -141
rect -1249 -181 -1234 -147
rect -1200 -181 -1162 -147
rect -1128 -181 -1090 -147
rect -1056 -181 -1041 -147
rect -1249 -187 -1041 -181
rect -791 -147 -583 -141
rect -791 -181 -776 -147
rect -742 -181 -704 -147
rect -670 -181 -632 -147
rect -598 -181 -583 -147
rect -791 -187 -583 -181
rect -333 -147 -125 -141
rect -333 -181 -318 -147
rect -284 -181 -246 -147
rect -212 -181 -174 -147
rect -140 -181 -125 -147
rect -333 -187 -125 -181
rect 125 -147 333 -141
rect 125 -181 140 -147
rect 174 -181 212 -147
rect 246 -181 284 -147
rect 318 -181 333 -147
rect 125 -187 333 -181
rect 583 -147 791 -141
rect 583 -181 598 -147
rect 632 -181 670 -147
rect 704 -181 742 -147
rect 776 -181 791 -147
rect 583 -187 791 -181
rect 1041 -147 1249 -141
rect 1041 -181 1056 -147
rect 1090 -181 1128 -147
rect 1162 -181 1200 -147
rect 1234 -181 1249 -147
rect 1041 -187 1249 -181
<< end >>
