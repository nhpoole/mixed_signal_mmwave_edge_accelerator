magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1296 -1309 2464 11211
<< metal1 >>
rect 552 9872 616 9924
rect 552 8458 616 8510
rect 552 7044 616 7096
rect 552 5630 616 5682
rect 552 4216 616 4268
rect 552 2802 616 2854
rect 552 1388 616 1440
rect 552 -26 616 26
<< metal2 >>
rect 137 9022 203 9074
rect 137 7894 203 7946
rect 137 6194 203 6246
rect 137 5066 203 5118
rect 137 3366 203 3418
rect 137 2238 203 2290
rect 137 538 203 590
rect 369 0 397 9898
rect 556 9874 612 9922
rect 1082 9093 1148 9145
rect 556 8460 612 8508
rect 1082 7823 1148 7875
rect 556 7046 612 7094
rect 1082 6265 1148 6317
rect 556 5632 612 5680
rect 1082 4995 1148 5047
rect 556 4218 612 4266
rect 1082 3437 1148 3489
rect 556 2804 612 2852
rect 1082 2167 1148 2219
rect 556 1390 612 1438
rect 1082 609 1148 661
rect 556 -24 612 24
<< metal3 >>
rect 535 9849 633 9947
rect 535 8435 633 8533
rect 535 7021 633 7119
rect 535 5607 633 5705
rect 535 4193 633 4291
rect 535 2779 633 2877
rect 535 1365 633 1463
rect 0 278 1168 338
rect 535 -49 633 49
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_6
timestamp 1626065694
transform 1 0 0 0 1 0
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_5
timestamp 1626065694
transform 1 0 0 0 -1 2828
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_4
timestamp 1626065694
transform 1 0 0 0 1 2828
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_3
timestamp 1626065694
transform 1 0 0 0 -1 5656
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_2
timestamp 1626065694
transform 1 0 0 0 1 5656
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_1
timestamp 1626065694
transform 1 0 0 0 -1 8484
box -36 -43 1204 1467
use sky130_fd_bd_sram__openram_dff  sky130_fd_bd_sram__openram_dff_0
timestamp 1626065694
transform 1 0 0 0 1 8484
box -36 -43 1204 1467
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1626065694
transform 1 0 363 0 1 271
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1626065694
transform 1 0 551 0 1 8447
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1626065694
transform 1 0 552 0 1 8452
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_0
timestamp 1626065694
transform 1 0 555 0 1 8451
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_2
timestamp 1626065694
transform 1 0 551 0 1 9861
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1626065694
transform 1 0 552 0 1 9866
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1
timestamp 1626065694
transform 1 0 555 0 1 9865
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_3
timestamp 1626065694
transform 1 0 551 0 1 8447
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1626065694
transform 1 0 552 0 1 8452
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_2
timestamp 1626065694
transform 1 0 555 0 1 8451
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_4
timestamp 1626065694
transform 1 0 551 0 1 7033
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_3
timestamp 1626065694
transform 1 0 552 0 1 7038
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_3
timestamp 1626065694
transform 1 0 555 0 1 7037
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_5
timestamp 1626065694
transform 1 0 551 0 1 5619
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_4
timestamp 1626065694
transform 1 0 552 0 1 5624
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_4
timestamp 1626065694
transform 1 0 555 0 1 5623
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_6
timestamp 1626065694
transform 1 0 551 0 1 7033
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_5
timestamp 1626065694
transform 1 0 552 0 1 7038
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_5
timestamp 1626065694
transform 1 0 555 0 1 7037
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_7
timestamp 1626065694
transform 1 0 551 0 1 5619
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_6
timestamp 1626065694
transform 1 0 552 0 1 5624
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_6
timestamp 1626065694
transform 1 0 555 0 1 5623
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_8
timestamp 1626065694
transform 1 0 551 0 1 4205
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_7
timestamp 1626065694
transform 1 0 552 0 1 4210
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_7
timestamp 1626065694
transform 1 0 555 0 1 4209
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_9
timestamp 1626065694
transform 1 0 551 0 1 2791
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_8
timestamp 1626065694
transform 1 0 552 0 1 2796
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_8
timestamp 1626065694
transform 1 0 555 0 1 2795
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_10
timestamp 1626065694
transform 1 0 551 0 1 4205
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_9
timestamp 1626065694
transform 1 0 552 0 1 4210
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_9
timestamp 1626065694
transform 1 0 555 0 1 4209
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_11
timestamp 1626065694
transform 1 0 551 0 1 2791
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_10
timestamp 1626065694
transform 1 0 552 0 1 2796
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_10
timestamp 1626065694
transform 1 0 555 0 1 2795
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_12
timestamp 1626065694
transform 1 0 551 0 1 1377
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_11
timestamp 1626065694
transform 1 0 552 0 1 1382
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_11
timestamp 1626065694
transform 1 0 555 0 1 1381
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_13
timestamp 1626065694
transform 1 0 551 0 1 -37
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_12
timestamp 1626065694
transform 1 0 552 0 1 -32
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_12
timestamp 1626065694
transform 1 0 555 0 1 -33
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_14
timestamp 1626065694
transform 1 0 551 0 1 1377
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_13
timestamp 1626065694
transform 1 0 552 0 1 1382
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_13
timestamp 1626065694
transform 1 0 555 0 1 1381
box 0 0 58 66
<< labels >>
rlabel metal3 s 535 7021 633 7119 4 vdd
rlabel metal3 s 535 1365 633 1463 4 vdd
rlabel metal3 s 535 4193 633 4291 4 vdd
rlabel metal3 s 535 9849 633 9947 4 vdd
rlabel metal3 s 535 2779 633 2877 4 gnd
rlabel metal3 s 535 -49 633 49 4 gnd
rlabel metal3 s 535 8435 633 8533 4 gnd
rlabel metal3 s 535 5607 633 5705 4 gnd
rlabel metal3 s 0 278 1168 338 4 clk
rlabel metal2 s 137 538 203 590 4 din_0
rlabel metal2 s 1082 609 1148 661 4 dout_0
rlabel metal2 s 137 2238 203 2290 4 din_1
rlabel metal2 s 1082 2167 1148 2219 4 dout_1
rlabel metal2 s 137 3366 203 3418 4 din_2
rlabel metal2 s 1082 3437 1148 3489 4 dout_2
rlabel metal2 s 137 5066 203 5118 4 din_3
rlabel metal2 s 1082 4995 1148 5047 4 dout_3
rlabel metal2 s 137 6194 203 6246 4 din_4
rlabel metal2 s 1082 6265 1148 6317 4 dout_4
rlabel metal2 s 137 7894 203 7946 4 din_5
rlabel metal2 s 1082 7823 1148 7875 4 dout_5
rlabel metal2 s 137 9022 203 9074 4 din_6
rlabel metal2 s 1082 9093 1148 9145 4 dout_6
<< properties >>
string FIXED_BBOX 0 0 1168 9898
<< end >>
