../../0-lvs_setup/outputs/design_extracted.spice