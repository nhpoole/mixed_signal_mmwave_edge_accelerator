magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -3026 -3428 43300 30798
<< pwell >>
rect -228 816 4428 968
rect -228 -1916 -76 816
rect 4276 -1916 4428 816
rect -228 -2068 4428 -1916
<< psubdiff >>
rect -202 909 4402 942
rect -202 875 -25 909
rect 9 875 43 909
rect 77 875 111 909
rect 145 875 179 909
rect 213 875 247 909
rect 281 875 315 909
rect 349 875 383 909
rect 417 875 451 909
rect 485 875 519 909
rect 553 875 587 909
rect 621 875 655 909
rect 689 875 723 909
rect 757 875 791 909
rect 825 875 859 909
rect 893 875 927 909
rect 961 875 995 909
rect 1029 875 1063 909
rect 1097 875 1131 909
rect 1165 875 1199 909
rect 1233 875 1267 909
rect 1301 875 1335 909
rect 1369 875 1403 909
rect 1437 875 1471 909
rect 1505 875 1539 909
rect 1573 875 1607 909
rect 1641 875 1675 909
rect 1709 875 1743 909
rect 1777 875 1811 909
rect 1845 875 1879 909
rect 1913 875 1947 909
rect 1981 875 2015 909
rect 2049 875 2083 909
rect 2117 875 2151 909
rect 2185 875 2219 909
rect 2253 875 2287 909
rect 2321 875 2355 909
rect 2389 875 2423 909
rect 2457 875 2491 909
rect 2525 875 2559 909
rect 2593 875 2627 909
rect 2661 875 2695 909
rect 2729 875 2763 909
rect 2797 875 2831 909
rect 2865 875 2899 909
rect 2933 875 2967 909
rect 3001 875 3035 909
rect 3069 875 3103 909
rect 3137 875 3171 909
rect 3205 875 3239 909
rect 3273 875 3307 909
rect 3341 875 3375 909
rect 3409 875 3443 909
rect 3477 875 3511 909
rect 3545 875 3579 909
rect 3613 875 3647 909
rect 3681 875 3715 909
rect 3749 875 3783 909
rect 3817 875 3851 909
rect 3885 875 3919 909
rect 3953 875 3987 909
rect 4021 875 4055 909
rect 4089 875 4123 909
rect 4157 875 4191 909
rect 4225 875 4402 909
rect -202 842 4402 875
rect -202 759 -102 842
rect -202 725 -169 759
rect -135 725 -102 759
rect -202 691 -102 725
rect -202 657 -169 691
rect -135 657 -102 691
rect -202 623 -102 657
rect -202 589 -169 623
rect -135 589 -102 623
rect -202 555 -102 589
rect -202 521 -169 555
rect -135 521 -102 555
rect -202 487 -102 521
rect -202 453 -169 487
rect -135 453 -102 487
rect -202 419 -102 453
rect -202 385 -169 419
rect -135 385 -102 419
rect -202 351 -102 385
rect -202 317 -169 351
rect -135 317 -102 351
rect -202 283 -102 317
rect -202 249 -169 283
rect -135 249 -102 283
rect -202 215 -102 249
rect -202 181 -169 215
rect -135 181 -102 215
rect -202 147 -102 181
rect -202 113 -169 147
rect -135 113 -102 147
rect -202 79 -102 113
rect -202 45 -169 79
rect -135 45 -102 79
rect -202 11 -102 45
rect -202 -23 -169 11
rect -135 -23 -102 11
rect -202 -57 -102 -23
rect -202 -91 -169 -57
rect -135 -91 -102 -57
rect -202 -125 -102 -91
rect -202 -159 -169 -125
rect -135 -159 -102 -125
rect -202 -193 -102 -159
rect -202 -227 -169 -193
rect -135 -227 -102 -193
rect -202 -261 -102 -227
rect -202 -295 -169 -261
rect -135 -295 -102 -261
rect -202 -329 -102 -295
rect -202 -363 -169 -329
rect -135 -363 -102 -329
rect -202 -397 -102 -363
rect -202 -431 -169 -397
rect -135 -431 -102 -397
rect -202 -465 -102 -431
rect -202 -499 -169 -465
rect -135 -499 -102 -465
rect -202 -533 -102 -499
rect -202 -567 -169 -533
rect -135 -567 -102 -533
rect -202 -601 -102 -567
rect -202 -635 -169 -601
rect -135 -635 -102 -601
rect -202 -669 -102 -635
rect -202 -703 -169 -669
rect -135 -703 -102 -669
rect -202 -737 -102 -703
rect -202 -771 -169 -737
rect -135 -771 -102 -737
rect -202 -805 -102 -771
rect -202 -839 -169 -805
rect -135 -839 -102 -805
rect -202 -873 -102 -839
rect -202 -907 -169 -873
rect -135 -907 -102 -873
rect -202 -941 -102 -907
rect -202 -975 -169 -941
rect -135 -975 -102 -941
rect -202 -1009 -102 -975
rect -202 -1043 -169 -1009
rect -135 -1043 -102 -1009
rect -202 -1077 -102 -1043
rect -202 -1111 -169 -1077
rect -135 -1111 -102 -1077
rect -202 -1145 -102 -1111
rect -202 -1179 -169 -1145
rect -135 -1179 -102 -1145
rect -202 -1213 -102 -1179
rect -202 -1247 -169 -1213
rect -135 -1247 -102 -1213
rect -202 -1281 -102 -1247
rect -202 -1315 -169 -1281
rect -135 -1315 -102 -1281
rect -202 -1349 -102 -1315
rect -202 -1383 -169 -1349
rect -135 -1383 -102 -1349
rect -202 -1417 -102 -1383
rect -202 -1451 -169 -1417
rect -135 -1451 -102 -1417
rect -202 -1485 -102 -1451
rect -202 -1519 -169 -1485
rect -135 -1519 -102 -1485
rect -202 -1553 -102 -1519
rect -202 -1587 -169 -1553
rect -135 -1587 -102 -1553
rect -202 -1621 -102 -1587
rect -202 -1655 -169 -1621
rect -135 -1655 -102 -1621
rect -202 -1689 -102 -1655
rect -202 -1723 -169 -1689
rect -135 -1723 -102 -1689
rect -202 -1757 -102 -1723
rect -202 -1791 -169 -1757
rect -135 -1791 -102 -1757
rect -202 -1825 -102 -1791
rect -202 -1859 -169 -1825
rect -135 -1859 -102 -1825
rect -202 -1942 -102 -1859
rect 4302 759 4402 842
rect 4302 725 4335 759
rect 4369 725 4402 759
rect 4302 691 4402 725
rect 4302 657 4335 691
rect 4369 657 4402 691
rect 4302 623 4402 657
rect 4302 589 4335 623
rect 4369 589 4402 623
rect 4302 555 4402 589
rect 4302 521 4335 555
rect 4369 521 4402 555
rect 4302 487 4402 521
rect 4302 453 4335 487
rect 4369 453 4402 487
rect 4302 419 4402 453
rect 4302 385 4335 419
rect 4369 385 4402 419
rect 4302 351 4402 385
rect 4302 317 4335 351
rect 4369 317 4402 351
rect 4302 283 4402 317
rect 4302 249 4335 283
rect 4369 249 4402 283
rect 4302 215 4402 249
rect 4302 181 4335 215
rect 4369 181 4402 215
rect 4302 147 4402 181
rect 4302 113 4335 147
rect 4369 113 4402 147
rect 4302 79 4402 113
rect 4302 45 4335 79
rect 4369 45 4402 79
rect 4302 11 4402 45
rect 4302 -23 4335 11
rect 4369 -23 4402 11
rect 4302 -57 4402 -23
rect 4302 -91 4335 -57
rect 4369 -91 4402 -57
rect 4302 -125 4402 -91
rect 4302 -159 4335 -125
rect 4369 -159 4402 -125
rect 4302 -193 4402 -159
rect 4302 -227 4335 -193
rect 4369 -227 4402 -193
rect 4302 -261 4402 -227
rect 4302 -295 4335 -261
rect 4369 -295 4402 -261
rect 4302 -329 4402 -295
rect 4302 -363 4335 -329
rect 4369 -363 4402 -329
rect 4302 -397 4402 -363
rect 4302 -431 4335 -397
rect 4369 -431 4402 -397
rect 4302 -465 4402 -431
rect 4302 -499 4335 -465
rect 4369 -499 4402 -465
rect 4302 -533 4402 -499
rect 4302 -567 4335 -533
rect 4369 -567 4402 -533
rect 4302 -601 4402 -567
rect 4302 -635 4335 -601
rect 4369 -635 4402 -601
rect 4302 -669 4402 -635
rect 4302 -703 4335 -669
rect 4369 -703 4402 -669
rect 4302 -737 4402 -703
rect 4302 -771 4335 -737
rect 4369 -771 4402 -737
rect 4302 -805 4402 -771
rect 4302 -839 4335 -805
rect 4369 -839 4402 -805
rect 4302 -873 4402 -839
rect 4302 -907 4335 -873
rect 4369 -907 4402 -873
rect 4302 -941 4402 -907
rect 4302 -975 4335 -941
rect 4369 -975 4402 -941
rect 4302 -1009 4402 -975
rect 4302 -1043 4335 -1009
rect 4369 -1043 4402 -1009
rect 4302 -1077 4402 -1043
rect 4302 -1111 4335 -1077
rect 4369 -1111 4402 -1077
rect 4302 -1145 4402 -1111
rect 4302 -1179 4335 -1145
rect 4369 -1179 4402 -1145
rect 4302 -1213 4402 -1179
rect 4302 -1247 4335 -1213
rect 4369 -1247 4402 -1213
rect 4302 -1281 4402 -1247
rect 4302 -1315 4335 -1281
rect 4369 -1315 4402 -1281
rect 4302 -1349 4402 -1315
rect 4302 -1383 4335 -1349
rect 4369 -1383 4402 -1349
rect 4302 -1417 4402 -1383
rect 4302 -1451 4335 -1417
rect 4369 -1451 4402 -1417
rect 4302 -1485 4402 -1451
rect 4302 -1519 4335 -1485
rect 4369 -1519 4402 -1485
rect 4302 -1553 4402 -1519
rect 4302 -1587 4335 -1553
rect 4369 -1587 4402 -1553
rect 4302 -1621 4402 -1587
rect 4302 -1655 4335 -1621
rect 4369 -1655 4402 -1621
rect 4302 -1689 4402 -1655
rect 4302 -1723 4335 -1689
rect 4369 -1723 4402 -1689
rect 4302 -1757 4402 -1723
rect 4302 -1791 4335 -1757
rect 4369 -1791 4402 -1757
rect 4302 -1825 4402 -1791
rect 4302 -1859 4335 -1825
rect 4369 -1859 4402 -1825
rect 4302 -1942 4402 -1859
rect -202 -1975 4402 -1942
rect -202 -2009 -25 -1975
rect 9 -2009 43 -1975
rect 77 -2009 111 -1975
rect 145 -2009 179 -1975
rect 213 -2009 247 -1975
rect 281 -2009 315 -1975
rect 349 -2009 383 -1975
rect 417 -2009 451 -1975
rect 485 -2009 519 -1975
rect 553 -2009 587 -1975
rect 621 -2009 655 -1975
rect 689 -2009 723 -1975
rect 757 -2009 791 -1975
rect 825 -2009 859 -1975
rect 893 -2009 927 -1975
rect 961 -2009 995 -1975
rect 1029 -2009 1063 -1975
rect 1097 -2009 1131 -1975
rect 1165 -2009 1199 -1975
rect 1233 -2009 1267 -1975
rect 1301 -2009 1335 -1975
rect 1369 -2009 1403 -1975
rect 1437 -2009 1471 -1975
rect 1505 -2009 1539 -1975
rect 1573 -2009 1607 -1975
rect 1641 -2009 1675 -1975
rect 1709 -2009 1743 -1975
rect 1777 -2009 1811 -1975
rect 1845 -2009 1879 -1975
rect 1913 -2009 1947 -1975
rect 1981 -2009 2015 -1975
rect 2049 -2009 2083 -1975
rect 2117 -2009 2151 -1975
rect 2185 -2009 2219 -1975
rect 2253 -2009 2287 -1975
rect 2321 -2009 2355 -1975
rect 2389 -2009 2423 -1975
rect 2457 -2009 2491 -1975
rect 2525 -2009 2559 -1975
rect 2593 -2009 2627 -1975
rect 2661 -2009 2695 -1975
rect 2729 -2009 2763 -1975
rect 2797 -2009 2831 -1975
rect 2865 -2009 2899 -1975
rect 2933 -2009 2967 -1975
rect 3001 -2009 3035 -1975
rect 3069 -2009 3103 -1975
rect 3137 -2009 3171 -1975
rect 3205 -2009 3239 -1975
rect 3273 -2009 3307 -1975
rect 3341 -2009 3375 -1975
rect 3409 -2009 3443 -1975
rect 3477 -2009 3511 -1975
rect 3545 -2009 3579 -1975
rect 3613 -2009 3647 -1975
rect 3681 -2009 3715 -1975
rect 3749 -2009 3783 -1975
rect 3817 -2009 3851 -1975
rect 3885 -2009 3919 -1975
rect 3953 -2009 3987 -1975
rect 4021 -2009 4055 -1975
rect 4089 -2009 4123 -1975
rect 4157 -2009 4191 -1975
rect 4225 -2009 4402 -1975
rect -202 -2042 4402 -2009
<< psubdiffcont >>
rect -25 875 9 909
rect 43 875 77 909
rect 111 875 145 909
rect 179 875 213 909
rect 247 875 281 909
rect 315 875 349 909
rect 383 875 417 909
rect 451 875 485 909
rect 519 875 553 909
rect 587 875 621 909
rect 655 875 689 909
rect 723 875 757 909
rect 791 875 825 909
rect 859 875 893 909
rect 927 875 961 909
rect 995 875 1029 909
rect 1063 875 1097 909
rect 1131 875 1165 909
rect 1199 875 1233 909
rect 1267 875 1301 909
rect 1335 875 1369 909
rect 1403 875 1437 909
rect 1471 875 1505 909
rect 1539 875 1573 909
rect 1607 875 1641 909
rect 1675 875 1709 909
rect 1743 875 1777 909
rect 1811 875 1845 909
rect 1879 875 1913 909
rect 1947 875 1981 909
rect 2015 875 2049 909
rect 2083 875 2117 909
rect 2151 875 2185 909
rect 2219 875 2253 909
rect 2287 875 2321 909
rect 2355 875 2389 909
rect 2423 875 2457 909
rect 2491 875 2525 909
rect 2559 875 2593 909
rect 2627 875 2661 909
rect 2695 875 2729 909
rect 2763 875 2797 909
rect 2831 875 2865 909
rect 2899 875 2933 909
rect 2967 875 3001 909
rect 3035 875 3069 909
rect 3103 875 3137 909
rect 3171 875 3205 909
rect 3239 875 3273 909
rect 3307 875 3341 909
rect 3375 875 3409 909
rect 3443 875 3477 909
rect 3511 875 3545 909
rect 3579 875 3613 909
rect 3647 875 3681 909
rect 3715 875 3749 909
rect 3783 875 3817 909
rect 3851 875 3885 909
rect 3919 875 3953 909
rect 3987 875 4021 909
rect 4055 875 4089 909
rect 4123 875 4157 909
rect 4191 875 4225 909
rect -169 725 -135 759
rect -169 657 -135 691
rect -169 589 -135 623
rect -169 521 -135 555
rect -169 453 -135 487
rect -169 385 -135 419
rect -169 317 -135 351
rect -169 249 -135 283
rect -169 181 -135 215
rect -169 113 -135 147
rect -169 45 -135 79
rect -169 -23 -135 11
rect -169 -91 -135 -57
rect -169 -159 -135 -125
rect -169 -227 -135 -193
rect -169 -295 -135 -261
rect -169 -363 -135 -329
rect -169 -431 -135 -397
rect -169 -499 -135 -465
rect -169 -567 -135 -533
rect -169 -635 -135 -601
rect -169 -703 -135 -669
rect -169 -771 -135 -737
rect -169 -839 -135 -805
rect -169 -907 -135 -873
rect -169 -975 -135 -941
rect -169 -1043 -135 -1009
rect -169 -1111 -135 -1077
rect -169 -1179 -135 -1145
rect -169 -1247 -135 -1213
rect -169 -1315 -135 -1281
rect -169 -1383 -135 -1349
rect -169 -1451 -135 -1417
rect -169 -1519 -135 -1485
rect -169 -1587 -135 -1553
rect -169 -1655 -135 -1621
rect -169 -1723 -135 -1689
rect -169 -1791 -135 -1757
rect -169 -1859 -135 -1825
rect 4335 725 4369 759
rect 4335 657 4369 691
rect 4335 589 4369 623
rect 4335 521 4369 555
rect 4335 453 4369 487
rect 4335 385 4369 419
rect 4335 317 4369 351
rect 4335 249 4369 283
rect 4335 181 4369 215
rect 4335 113 4369 147
rect 4335 45 4369 79
rect 4335 -23 4369 11
rect 4335 -91 4369 -57
rect 4335 -159 4369 -125
rect 4335 -227 4369 -193
rect 4335 -295 4369 -261
rect 4335 -363 4369 -329
rect 4335 -431 4369 -397
rect 4335 -499 4369 -465
rect 4335 -567 4369 -533
rect 4335 -635 4369 -601
rect 4335 -703 4369 -669
rect 4335 -771 4369 -737
rect 4335 -839 4369 -805
rect 4335 -907 4369 -873
rect 4335 -975 4369 -941
rect 4335 -1043 4369 -1009
rect 4335 -1111 4369 -1077
rect 4335 -1179 4369 -1145
rect 4335 -1247 4369 -1213
rect 4335 -1315 4369 -1281
rect 4335 -1383 4369 -1349
rect 4335 -1451 4369 -1417
rect 4335 -1519 4369 -1485
rect 4335 -1587 4369 -1553
rect 4335 -1655 4369 -1621
rect 4335 -1723 4369 -1689
rect 4335 -1791 4369 -1757
rect 4335 -1859 4369 -1825
rect -25 -2009 9 -1975
rect 43 -2009 77 -1975
rect 111 -2009 145 -1975
rect 179 -2009 213 -1975
rect 247 -2009 281 -1975
rect 315 -2009 349 -1975
rect 383 -2009 417 -1975
rect 451 -2009 485 -1975
rect 519 -2009 553 -1975
rect 587 -2009 621 -1975
rect 655 -2009 689 -1975
rect 723 -2009 757 -1975
rect 791 -2009 825 -1975
rect 859 -2009 893 -1975
rect 927 -2009 961 -1975
rect 995 -2009 1029 -1975
rect 1063 -2009 1097 -1975
rect 1131 -2009 1165 -1975
rect 1199 -2009 1233 -1975
rect 1267 -2009 1301 -1975
rect 1335 -2009 1369 -1975
rect 1403 -2009 1437 -1975
rect 1471 -2009 1505 -1975
rect 1539 -2009 1573 -1975
rect 1607 -2009 1641 -1975
rect 1675 -2009 1709 -1975
rect 1743 -2009 1777 -1975
rect 1811 -2009 1845 -1975
rect 1879 -2009 1913 -1975
rect 1947 -2009 1981 -1975
rect 2015 -2009 2049 -1975
rect 2083 -2009 2117 -1975
rect 2151 -2009 2185 -1975
rect 2219 -2009 2253 -1975
rect 2287 -2009 2321 -1975
rect 2355 -2009 2389 -1975
rect 2423 -2009 2457 -1975
rect 2491 -2009 2525 -1975
rect 2559 -2009 2593 -1975
rect 2627 -2009 2661 -1975
rect 2695 -2009 2729 -1975
rect 2763 -2009 2797 -1975
rect 2831 -2009 2865 -1975
rect 2899 -2009 2933 -1975
rect 2967 -2009 3001 -1975
rect 3035 -2009 3069 -1975
rect 3103 -2009 3137 -1975
rect 3171 -2009 3205 -1975
rect 3239 -2009 3273 -1975
rect 3307 -2009 3341 -1975
rect 3375 -2009 3409 -1975
rect 3443 -2009 3477 -1975
rect 3511 -2009 3545 -1975
rect 3579 -2009 3613 -1975
rect 3647 -2009 3681 -1975
rect 3715 -2009 3749 -1975
rect 3783 -2009 3817 -1975
rect 3851 -2009 3885 -1975
rect 3919 -2009 3953 -1975
rect 3987 -2009 4021 -1975
rect 4055 -2009 4089 -1975
rect 4123 -2009 4157 -1975
rect 4191 -2009 4225 -1975
<< locali >>
rect -202 909 4402 942
rect -202 875 -77 909
rect -43 875 -25 909
rect 29 875 43 909
rect 101 875 111 909
rect 173 875 179 909
rect 245 875 247 909
rect 281 875 283 909
rect 349 875 355 909
rect 417 875 427 909
rect 485 875 499 909
rect 553 875 571 909
rect 621 875 643 909
rect 689 875 715 909
rect 757 875 787 909
rect 825 875 859 909
rect 893 875 927 909
rect 965 875 995 909
rect 1037 875 1063 909
rect 1109 875 1131 909
rect 1181 875 1199 909
rect 1253 875 1267 909
rect 1325 875 1335 909
rect 1397 875 1403 909
rect 1469 875 1471 909
rect 1505 875 1507 909
rect 1573 875 1579 909
rect 1641 875 1651 909
rect 1709 875 1723 909
rect 1777 875 1795 909
rect 1845 875 1867 909
rect 1913 875 1939 909
rect 1981 875 2011 909
rect 2049 875 2083 909
rect 2117 875 2151 909
rect 2189 875 2219 909
rect 2261 875 2287 909
rect 2333 875 2355 909
rect 2405 875 2423 909
rect 2477 875 2491 909
rect 2549 875 2559 909
rect 2621 875 2627 909
rect 2693 875 2695 909
rect 2729 875 2731 909
rect 2797 875 2803 909
rect 2865 875 2875 909
rect 2933 875 2947 909
rect 3001 875 3019 909
rect 3069 875 3091 909
rect 3137 875 3163 909
rect 3205 875 3235 909
rect 3273 875 3307 909
rect 3341 875 3375 909
rect 3413 875 3443 909
rect 3485 875 3511 909
rect 3557 875 3579 909
rect 3629 875 3647 909
rect 3701 875 3715 909
rect 3773 875 3783 909
rect 3845 875 3851 909
rect 3917 875 3919 909
rect 3953 875 3955 909
rect 4021 875 4027 909
rect 4089 875 4099 909
rect 4157 875 4171 909
rect 4225 875 4243 909
rect 4277 875 4402 909
rect -202 842 4402 875
rect -202 759 -102 842
rect -202 725 -169 759
rect -135 725 -102 759
rect -202 691 -102 725
rect -202 657 -169 691
rect -135 657 -102 691
rect -202 655 -102 657
rect -202 589 -169 655
rect -135 589 -102 655
rect -202 583 -102 589
rect -202 521 -169 583
rect -135 521 -102 583
rect -202 511 -102 521
rect -202 453 -169 511
rect -135 453 -102 511
rect -202 439 -102 453
rect -202 385 -169 439
rect -135 385 -102 439
rect -202 367 -102 385
rect -202 317 -169 367
rect -135 317 -102 367
rect -202 295 -102 317
rect -202 249 -169 295
rect -135 249 -102 295
rect -202 223 -102 249
rect -202 181 -169 223
rect -135 181 -102 223
rect -202 151 -102 181
rect -202 113 -169 151
rect -135 113 -102 151
rect -202 79 -102 113
rect -202 45 -169 79
rect -135 45 -102 79
rect -202 11 -102 45
rect -202 -27 -169 11
rect -135 -27 -102 11
rect -202 -57 -102 -27
rect -202 -99 -169 -57
rect -135 -99 -102 -57
rect -202 -125 -102 -99
rect -202 -171 -169 -125
rect -135 -171 -102 -125
rect -202 -193 -102 -171
rect -202 -243 -169 -193
rect -135 -243 -102 -193
rect -202 -261 -102 -243
rect -202 -315 -169 -261
rect -135 -315 -102 -261
rect -202 -329 -102 -315
rect -202 -387 -169 -329
rect -135 -387 -102 -329
rect -202 -397 -102 -387
rect -202 -459 -169 -397
rect -135 -459 -102 -397
rect -202 -465 -102 -459
rect -202 -531 -169 -465
rect -135 -531 -102 -465
rect -202 -533 -102 -531
rect -202 -567 -169 -533
rect -135 -567 -102 -533
rect -202 -569 -102 -567
rect -202 -635 -169 -569
rect -135 -635 -102 -569
rect -202 -641 -102 -635
rect -202 -703 -169 -641
rect -135 -703 -102 -641
rect -202 -713 -102 -703
rect -202 -771 -169 -713
rect -135 -771 -102 -713
rect -202 -785 -102 -771
rect -202 -839 -169 -785
rect -135 -839 -102 -785
rect -202 -857 -102 -839
rect -202 -907 -169 -857
rect -135 -907 -102 -857
rect -202 -929 -102 -907
rect -202 -975 -169 -929
rect -135 -975 -102 -929
rect -202 -1001 -102 -975
rect -202 -1043 -169 -1001
rect -135 -1043 -102 -1001
rect -202 -1073 -102 -1043
rect -202 -1111 -169 -1073
rect -135 -1111 -102 -1073
rect -202 -1145 -102 -1111
rect -202 -1179 -169 -1145
rect -135 -1179 -102 -1145
rect -202 -1213 -102 -1179
rect -202 -1251 -169 -1213
rect -135 -1251 -102 -1213
rect -202 -1281 -102 -1251
rect -202 -1323 -169 -1281
rect -135 -1323 -102 -1281
rect -202 -1349 -102 -1323
rect -202 -1395 -169 -1349
rect -135 -1395 -102 -1349
rect -202 -1417 -102 -1395
rect -202 -1467 -169 -1417
rect -135 -1467 -102 -1417
rect -202 -1485 -102 -1467
rect -202 -1539 -169 -1485
rect -135 -1539 -102 -1485
rect -202 -1553 -102 -1539
rect -202 -1611 -169 -1553
rect -135 -1611 -102 -1553
rect -202 -1621 -102 -1611
rect -202 -1683 -169 -1621
rect -135 -1683 -102 -1621
rect -202 -1689 -102 -1683
rect -202 -1755 -169 -1689
rect -135 -1755 -102 -1689
rect -202 -1757 -102 -1755
rect -202 -1791 -169 -1757
rect -135 -1791 -102 -1757
rect -202 -1825 -102 -1791
rect -202 -1859 -169 -1825
rect -135 -1859 -102 -1825
rect -202 -1942 -102 -1859
rect 4302 759 4402 842
rect 4302 725 4335 759
rect 4369 725 4402 759
rect 4302 691 4402 725
rect 4302 657 4335 691
rect 4369 657 4402 691
rect 4302 655 4402 657
rect 4302 589 4335 655
rect 4369 589 4402 655
rect 4302 583 4402 589
rect 4302 521 4335 583
rect 4369 521 4402 583
rect 4302 511 4402 521
rect 4302 453 4335 511
rect 4369 453 4402 511
rect 4302 439 4402 453
rect 4302 385 4335 439
rect 4369 385 4402 439
rect 4302 367 4402 385
rect 4302 317 4335 367
rect 4369 317 4402 367
rect 4302 295 4402 317
rect 4302 249 4335 295
rect 4369 249 4402 295
rect 4302 223 4402 249
rect 4302 181 4335 223
rect 4369 181 4402 223
rect 4302 151 4402 181
rect 4302 113 4335 151
rect 4369 113 4402 151
rect 4302 79 4402 113
rect 4302 45 4335 79
rect 4369 45 4402 79
rect 4302 11 4402 45
rect 4302 -27 4335 11
rect 4369 -27 4402 11
rect 4302 -57 4402 -27
rect 4302 -99 4335 -57
rect 4369 -99 4402 -57
rect 4302 -125 4402 -99
rect 4302 -171 4335 -125
rect 4369 -171 4402 -125
rect 4302 -193 4402 -171
rect 4302 -243 4335 -193
rect 4369 -243 4402 -193
rect 4302 -261 4402 -243
rect 4302 -315 4335 -261
rect 4369 -315 4402 -261
rect 4302 -329 4402 -315
rect 4302 -387 4335 -329
rect 4369 -387 4402 -329
rect 4302 -397 4402 -387
rect 4302 -459 4335 -397
rect 4369 -459 4402 -397
rect 4302 -465 4402 -459
rect 4302 -531 4335 -465
rect 4369 -531 4402 -465
rect 4302 -533 4402 -531
rect 4302 -567 4335 -533
rect 4369 -567 4402 -533
rect 4302 -569 4402 -567
rect 4302 -635 4335 -569
rect 4369 -635 4402 -569
rect 4302 -641 4402 -635
rect 4302 -703 4335 -641
rect 4369 -703 4402 -641
rect 4302 -713 4402 -703
rect 4302 -771 4335 -713
rect 4369 -771 4402 -713
rect 4302 -785 4402 -771
rect 4302 -839 4335 -785
rect 4369 -839 4402 -785
rect 4302 -857 4402 -839
rect 4302 -907 4335 -857
rect 4369 -907 4402 -857
rect 4302 -929 4402 -907
rect 4302 -975 4335 -929
rect 4369 -975 4402 -929
rect 4302 -1001 4402 -975
rect 4302 -1043 4335 -1001
rect 4369 -1043 4402 -1001
rect 4302 -1073 4402 -1043
rect 4302 -1111 4335 -1073
rect 4369 -1111 4402 -1073
rect 4302 -1145 4402 -1111
rect 4302 -1179 4335 -1145
rect 4369 -1179 4402 -1145
rect 4302 -1213 4402 -1179
rect 4302 -1251 4335 -1213
rect 4369 -1251 4402 -1213
rect 4302 -1281 4402 -1251
rect 4302 -1323 4335 -1281
rect 4369 -1323 4402 -1281
rect 4302 -1349 4402 -1323
rect 4302 -1395 4335 -1349
rect 4369 -1395 4402 -1349
rect 4302 -1417 4402 -1395
rect 4302 -1467 4335 -1417
rect 4369 -1467 4402 -1417
rect 4302 -1485 4402 -1467
rect 4302 -1539 4335 -1485
rect 4369 -1539 4402 -1485
rect 4302 -1553 4402 -1539
rect 4302 -1611 4335 -1553
rect 4369 -1611 4402 -1553
rect 4302 -1621 4402 -1611
rect 4302 -1683 4335 -1621
rect 4369 -1683 4402 -1621
rect 4302 -1689 4402 -1683
rect 4302 -1755 4335 -1689
rect 4369 -1755 4402 -1689
rect 4302 -1757 4402 -1755
rect 4302 -1791 4335 -1757
rect 4369 -1791 4402 -1757
rect 4302 -1825 4402 -1791
rect 4302 -1859 4335 -1825
rect 4369 -1859 4402 -1825
rect 4302 -1942 4402 -1859
rect -202 -1975 4402 -1942
rect -202 -2009 -77 -1975
rect -43 -2009 -25 -1975
rect 29 -2009 43 -1975
rect 101 -2009 111 -1975
rect 173 -2009 179 -1975
rect 245 -2009 247 -1975
rect 281 -2009 283 -1975
rect 349 -2009 355 -1975
rect 417 -2009 427 -1975
rect 485 -2009 499 -1975
rect 553 -2009 571 -1975
rect 621 -2009 643 -1975
rect 689 -2009 715 -1975
rect 757 -2009 787 -1975
rect 825 -2009 859 -1975
rect 893 -2009 927 -1975
rect 965 -2009 995 -1975
rect 1037 -2009 1063 -1975
rect 1109 -2009 1131 -1975
rect 1181 -2009 1199 -1975
rect 1253 -2009 1267 -1975
rect 1325 -2009 1335 -1975
rect 1397 -2009 1403 -1975
rect 1469 -2009 1471 -1975
rect 1505 -2009 1507 -1975
rect 1573 -2009 1579 -1975
rect 1641 -2009 1651 -1975
rect 1709 -2009 1723 -1975
rect 1777 -2009 1795 -1975
rect 1845 -2009 1867 -1975
rect 1913 -2009 1939 -1975
rect 1981 -2009 2011 -1975
rect 2049 -2009 2083 -1975
rect 2117 -2009 2151 -1975
rect 2189 -2009 2219 -1975
rect 2261 -2009 2287 -1975
rect 2333 -2009 2355 -1975
rect 2405 -2009 2423 -1975
rect 2477 -2009 2491 -1975
rect 2549 -2009 2559 -1975
rect 2621 -2009 2627 -1975
rect 2693 -2009 2695 -1975
rect 2729 -2009 2731 -1975
rect 2797 -2009 2803 -1975
rect 2865 -2009 2875 -1975
rect 2933 -2009 2947 -1975
rect 3001 -2009 3019 -1975
rect 3069 -2009 3091 -1975
rect 3137 -2009 3163 -1975
rect 3205 -2009 3235 -1975
rect 3273 -2009 3307 -1975
rect 3341 -2009 3375 -1975
rect 3413 -2009 3443 -1975
rect 3485 -2009 3511 -1975
rect 3557 -2009 3579 -1975
rect 3629 -2009 3647 -1975
rect 3701 -2009 3715 -1975
rect 3773 -2009 3783 -1975
rect 3845 -2009 3851 -1975
rect 3917 -2009 3919 -1975
rect 3953 -2009 3955 -1975
rect 4021 -2009 4027 -1975
rect 4089 -2009 4099 -1975
rect 4157 -2009 4171 -1975
rect 4225 -2009 4243 -1975
rect 4277 -2009 4402 -1975
rect -202 -2042 4402 -2009
<< viali >>
rect -77 875 -43 909
rect -5 875 9 909
rect 9 875 29 909
rect 67 875 77 909
rect 77 875 101 909
rect 139 875 145 909
rect 145 875 173 909
rect 211 875 213 909
rect 213 875 245 909
rect 283 875 315 909
rect 315 875 317 909
rect 355 875 383 909
rect 383 875 389 909
rect 427 875 451 909
rect 451 875 461 909
rect 499 875 519 909
rect 519 875 533 909
rect 571 875 587 909
rect 587 875 605 909
rect 643 875 655 909
rect 655 875 677 909
rect 715 875 723 909
rect 723 875 749 909
rect 787 875 791 909
rect 791 875 821 909
rect 859 875 893 909
rect 931 875 961 909
rect 961 875 965 909
rect 1003 875 1029 909
rect 1029 875 1037 909
rect 1075 875 1097 909
rect 1097 875 1109 909
rect 1147 875 1165 909
rect 1165 875 1181 909
rect 1219 875 1233 909
rect 1233 875 1253 909
rect 1291 875 1301 909
rect 1301 875 1325 909
rect 1363 875 1369 909
rect 1369 875 1397 909
rect 1435 875 1437 909
rect 1437 875 1469 909
rect 1507 875 1539 909
rect 1539 875 1541 909
rect 1579 875 1607 909
rect 1607 875 1613 909
rect 1651 875 1675 909
rect 1675 875 1685 909
rect 1723 875 1743 909
rect 1743 875 1757 909
rect 1795 875 1811 909
rect 1811 875 1829 909
rect 1867 875 1879 909
rect 1879 875 1901 909
rect 1939 875 1947 909
rect 1947 875 1973 909
rect 2011 875 2015 909
rect 2015 875 2045 909
rect 2083 875 2117 909
rect 2155 875 2185 909
rect 2185 875 2189 909
rect 2227 875 2253 909
rect 2253 875 2261 909
rect 2299 875 2321 909
rect 2321 875 2333 909
rect 2371 875 2389 909
rect 2389 875 2405 909
rect 2443 875 2457 909
rect 2457 875 2477 909
rect 2515 875 2525 909
rect 2525 875 2549 909
rect 2587 875 2593 909
rect 2593 875 2621 909
rect 2659 875 2661 909
rect 2661 875 2693 909
rect 2731 875 2763 909
rect 2763 875 2765 909
rect 2803 875 2831 909
rect 2831 875 2837 909
rect 2875 875 2899 909
rect 2899 875 2909 909
rect 2947 875 2967 909
rect 2967 875 2981 909
rect 3019 875 3035 909
rect 3035 875 3053 909
rect 3091 875 3103 909
rect 3103 875 3125 909
rect 3163 875 3171 909
rect 3171 875 3197 909
rect 3235 875 3239 909
rect 3239 875 3269 909
rect 3307 875 3341 909
rect 3379 875 3409 909
rect 3409 875 3413 909
rect 3451 875 3477 909
rect 3477 875 3485 909
rect 3523 875 3545 909
rect 3545 875 3557 909
rect 3595 875 3613 909
rect 3613 875 3629 909
rect 3667 875 3681 909
rect 3681 875 3701 909
rect 3739 875 3749 909
rect 3749 875 3773 909
rect 3811 875 3817 909
rect 3817 875 3845 909
rect 3883 875 3885 909
rect 3885 875 3917 909
rect 3955 875 3987 909
rect 3987 875 3989 909
rect 4027 875 4055 909
rect 4055 875 4061 909
rect 4099 875 4123 909
rect 4123 875 4133 909
rect 4171 875 4191 909
rect 4191 875 4205 909
rect 4243 875 4277 909
rect -169 623 -135 655
rect -169 621 -135 623
rect -169 555 -135 583
rect -169 549 -135 555
rect -169 487 -135 511
rect -169 477 -135 487
rect -169 419 -135 439
rect -169 405 -135 419
rect -169 351 -135 367
rect -169 333 -135 351
rect -169 283 -135 295
rect -169 261 -135 283
rect -169 215 -135 223
rect -169 189 -135 215
rect -169 147 -135 151
rect -169 117 -135 147
rect -169 45 -135 79
rect -169 -23 -135 7
rect -169 -27 -135 -23
rect -169 -91 -135 -65
rect -169 -99 -135 -91
rect -169 -159 -135 -137
rect -169 -171 -135 -159
rect -169 -227 -135 -209
rect -169 -243 -135 -227
rect -169 -295 -135 -281
rect -169 -315 -135 -295
rect -169 -363 -135 -353
rect -169 -387 -135 -363
rect -169 -431 -135 -425
rect -169 -459 -135 -431
rect -169 -499 -135 -497
rect -169 -531 -135 -499
rect -169 -601 -135 -569
rect -169 -603 -135 -601
rect -169 -669 -135 -641
rect -169 -675 -135 -669
rect -169 -737 -135 -713
rect -169 -747 -135 -737
rect -169 -805 -135 -785
rect -169 -819 -135 -805
rect -169 -873 -135 -857
rect -169 -891 -135 -873
rect -169 -941 -135 -929
rect -169 -963 -135 -941
rect -169 -1009 -135 -1001
rect -169 -1035 -135 -1009
rect -169 -1077 -135 -1073
rect -169 -1107 -135 -1077
rect -169 -1179 -135 -1145
rect -169 -1247 -135 -1217
rect -169 -1251 -135 -1247
rect -169 -1315 -135 -1289
rect -169 -1323 -135 -1315
rect -169 -1383 -135 -1361
rect -169 -1395 -135 -1383
rect -169 -1451 -135 -1433
rect -169 -1467 -135 -1451
rect -169 -1519 -135 -1505
rect -169 -1539 -135 -1519
rect -169 -1587 -135 -1577
rect -169 -1611 -135 -1587
rect -169 -1655 -135 -1649
rect -169 -1683 -135 -1655
rect -169 -1723 -135 -1721
rect -169 -1755 -135 -1723
rect 4335 623 4369 655
rect 4335 621 4369 623
rect 4335 555 4369 583
rect 4335 549 4369 555
rect 4335 487 4369 511
rect 4335 477 4369 487
rect 4335 419 4369 439
rect 4335 405 4369 419
rect 4335 351 4369 367
rect 4335 333 4369 351
rect 4335 283 4369 295
rect 4335 261 4369 283
rect 4335 215 4369 223
rect 4335 189 4369 215
rect 4335 147 4369 151
rect 4335 117 4369 147
rect 4335 45 4369 79
rect 4335 -23 4369 7
rect 4335 -27 4369 -23
rect 4335 -91 4369 -65
rect 4335 -99 4369 -91
rect 4335 -159 4369 -137
rect 4335 -171 4369 -159
rect 4335 -227 4369 -209
rect 4335 -243 4369 -227
rect 4335 -295 4369 -281
rect 4335 -315 4369 -295
rect 4335 -363 4369 -353
rect 4335 -387 4369 -363
rect 4335 -431 4369 -425
rect 4335 -459 4369 -431
rect 4335 -499 4369 -497
rect 4335 -531 4369 -499
rect 4335 -601 4369 -569
rect 4335 -603 4369 -601
rect 4335 -669 4369 -641
rect 4335 -675 4369 -669
rect 4335 -737 4369 -713
rect 4335 -747 4369 -737
rect 4335 -805 4369 -785
rect 4335 -819 4369 -805
rect 4335 -873 4369 -857
rect 4335 -891 4369 -873
rect 4335 -941 4369 -929
rect 4335 -963 4369 -941
rect 4335 -1009 4369 -1001
rect 4335 -1035 4369 -1009
rect 4335 -1077 4369 -1073
rect 4335 -1107 4369 -1077
rect 4335 -1179 4369 -1145
rect 4335 -1247 4369 -1217
rect 4335 -1251 4369 -1247
rect 4335 -1315 4369 -1289
rect 4335 -1323 4369 -1315
rect 4335 -1383 4369 -1361
rect 4335 -1395 4369 -1383
rect 4335 -1451 4369 -1433
rect 4335 -1467 4369 -1451
rect 4335 -1519 4369 -1505
rect 4335 -1539 4369 -1519
rect 4335 -1587 4369 -1577
rect 4335 -1611 4369 -1587
rect 4335 -1655 4369 -1649
rect 4335 -1683 4369 -1655
rect 4335 -1723 4369 -1721
rect 4335 -1755 4369 -1723
rect -77 -2009 -43 -1975
rect -5 -2009 9 -1975
rect 9 -2009 29 -1975
rect 67 -2009 77 -1975
rect 77 -2009 101 -1975
rect 139 -2009 145 -1975
rect 145 -2009 173 -1975
rect 211 -2009 213 -1975
rect 213 -2009 245 -1975
rect 283 -2009 315 -1975
rect 315 -2009 317 -1975
rect 355 -2009 383 -1975
rect 383 -2009 389 -1975
rect 427 -2009 451 -1975
rect 451 -2009 461 -1975
rect 499 -2009 519 -1975
rect 519 -2009 533 -1975
rect 571 -2009 587 -1975
rect 587 -2009 605 -1975
rect 643 -2009 655 -1975
rect 655 -2009 677 -1975
rect 715 -2009 723 -1975
rect 723 -2009 749 -1975
rect 787 -2009 791 -1975
rect 791 -2009 821 -1975
rect 859 -2009 893 -1975
rect 931 -2009 961 -1975
rect 961 -2009 965 -1975
rect 1003 -2009 1029 -1975
rect 1029 -2009 1037 -1975
rect 1075 -2009 1097 -1975
rect 1097 -2009 1109 -1975
rect 1147 -2009 1165 -1975
rect 1165 -2009 1181 -1975
rect 1219 -2009 1233 -1975
rect 1233 -2009 1253 -1975
rect 1291 -2009 1301 -1975
rect 1301 -2009 1325 -1975
rect 1363 -2009 1369 -1975
rect 1369 -2009 1397 -1975
rect 1435 -2009 1437 -1975
rect 1437 -2009 1469 -1975
rect 1507 -2009 1539 -1975
rect 1539 -2009 1541 -1975
rect 1579 -2009 1607 -1975
rect 1607 -2009 1613 -1975
rect 1651 -2009 1675 -1975
rect 1675 -2009 1685 -1975
rect 1723 -2009 1743 -1975
rect 1743 -2009 1757 -1975
rect 1795 -2009 1811 -1975
rect 1811 -2009 1829 -1975
rect 1867 -2009 1879 -1975
rect 1879 -2009 1901 -1975
rect 1939 -2009 1947 -1975
rect 1947 -2009 1973 -1975
rect 2011 -2009 2015 -1975
rect 2015 -2009 2045 -1975
rect 2083 -2009 2117 -1975
rect 2155 -2009 2185 -1975
rect 2185 -2009 2189 -1975
rect 2227 -2009 2253 -1975
rect 2253 -2009 2261 -1975
rect 2299 -2009 2321 -1975
rect 2321 -2009 2333 -1975
rect 2371 -2009 2389 -1975
rect 2389 -2009 2405 -1975
rect 2443 -2009 2457 -1975
rect 2457 -2009 2477 -1975
rect 2515 -2009 2525 -1975
rect 2525 -2009 2549 -1975
rect 2587 -2009 2593 -1975
rect 2593 -2009 2621 -1975
rect 2659 -2009 2661 -1975
rect 2661 -2009 2693 -1975
rect 2731 -2009 2763 -1975
rect 2763 -2009 2765 -1975
rect 2803 -2009 2831 -1975
rect 2831 -2009 2837 -1975
rect 2875 -2009 2899 -1975
rect 2899 -2009 2909 -1975
rect 2947 -2009 2967 -1975
rect 2967 -2009 2981 -1975
rect 3019 -2009 3035 -1975
rect 3035 -2009 3053 -1975
rect 3091 -2009 3103 -1975
rect 3103 -2009 3125 -1975
rect 3163 -2009 3171 -1975
rect 3171 -2009 3197 -1975
rect 3235 -2009 3239 -1975
rect 3239 -2009 3269 -1975
rect 3307 -2009 3341 -1975
rect 3379 -2009 3409 -1975
rect 3409 -2009 3413 -1975
rect 3451 -2009 3477 -1975
rect 3477 -2009 3485 -1975
rect 3523 -2009 3545 -1975
rect 3545 -2009 3557 -1975
rect 3595 -2009 3613 -1975
rect 3613 -2009 3629 -1975
rect 3667 -2009 3681 -1975
rect 3681 -2009 3701 -1975
rect 3739 -2009 3749 -1975
rect 3749 -2009 3773 -1975
rect 3811 -2009 3817 -1975
rect 3817 -2009 3845 -1975
rect 3883 -2009 3885 -1975
rect 3885 -2009 3917 -1975
rect 3955 -2009 3987 -1975
rect 3987 -2009 3989 -1975
rect 4027 -2009 4055 -1975
rect 4055 -2009 4061 -1975
rect 4099 -2009 4123 -1975
rect 4123 -2009 4133 -1975
rect 4171 -2009 4191 -1975
rect 4191 -2009 4205 -1975
rect 4243 -2009 4277 -1975
<< metal1 >>
rect 4662 12780 5100 12860
rect 4662 1208 4711 12780
rect 4955 1208 5100 12780
rect 4662 1148 5100 1208
rect -210 967 4968 1022
rect -210 915 -138 967
rect -86 915 -74 967
rect -22 915 -10 967
rect 42 915 54 967
rect 106 915 118 967
rect 170 915 182 967
rect 234 915 246 967
rect 298 915 310 967
rect 362 915 374 967
rect 426 915 438 967
rect 490 915 502 967
rect 554 915 566 967
rect 618 915 630 967
rect 682 915 694 967
rect 746 915 758 967
rect 810 915 822 967
rect 874 915 886 967
rect 938 915 950 967
rect 1002 915 1014 967
rect 1066 915 1078 967
rect 1130 915 1142 967
rect 1194 915 1206 967
rect 1258 915 1270 967
rect 1322 915 1334 967
rect 1386 915 1398 967
rect 1450 915 1462 967
rect 1514 915 1526 967
rect 1578 915 1590 967
rect 1642 915 1654 967
rect 1706 915 1718 967
rect 1770 915 1782 967
rect 1834 915 1846 967
rect 1898 915 1910 967
rect 1962 915 1974 967
rect 2026 915 2038 967
rect 2090 915 2102 967
rect 2154 915 2166 967
rect 2218 915 2230 967
rect 2282 915 2294 967
rect 2346 915 2358 967
rect 2410 915 2422 967
rect 2474 915 2486 967
rect 2538 915 2550 967
rect 2602 915 2614 967
rect 2666 915 2678 967
rect 2730 915 2742 967
rect 2794 915 2806 967
rect 2858 915 2870 967
rect 2922 915 2934 967
rect 2986 915 2998 967
rect 3050 915 3062 967
rect 3114 915 3126 967
rect 3178 915 3190 967
rect 3242 915 3254 967
rect 3306 915 3318 967
rect 3370 915 3382 967
rect 3434 915 3446 967
rect 3498 915 3510 967
rect 3562 915 3574 967
rect 3626 915 3638 967
rect 3690 915 3702 967
rect 3754 915 3766 967
rect 3818 915 3830 967
rect 3882 915 3894 967
rect 3946 915 3958 967
rect 4010 915 4022 967
rect 4074 915 4086 967
rect 4138 915 4150 967
rect 4202 915 4214 967
rect 4266 915 4278 967
rect 4330 915 4342 967
rect 4394 915 4406 967
rect 4458 915 4470 967
rect 4522 915 4534 967
rect 4586 915 4598 967
rect 4650 915 4662 967
rect 4714 915 4726 967
rect 4778 915 4790 967
rect 4842 915 4854 967
rect 4906 915 4968 967
rect -210 909 4968 915
rect -210 875 -77 909
rect -43 875 -5 909
rect 29 875 67 909
rect 101 875 139 909
rect 173 875 211 909
rect 245 875 283 909
rect 317 875 355 909
rect 389 875 427 909
rect 461 875 499 909
rect 533 875 571 909
rect 605 875 643 909
rect 677 875 715 909
rect 749 875 787 909
rect 821 875 859 909
rect 893 875 931 909
rect 965 875 1003 909
rect 1037 875 1075 909
rect 1109 875 1147 909
rect 1181 875 1219 909
rect 1253 875 1291 909
rect 1325 875 1363 909
rect 1397 875 1435 909
rect 1469 875 1507 909
rect 1541 875 1579 909
rect 1613 875 1651 909
rect 1685 875 1723 909
rect 1757 875 1795 909
rect 1829 875 1867 909
rect 1901 875 1939 909
rect 1973 875 2011 909
rect 2045 875 2083 909
rect 2117 875 2155 909
rect 2189 875 2227 909
rect 2261 875 2299 909
rect 2333 875 2371 909
rect 2405 875 2443 909
rect 2477 875 2515 909
rect 2549 875 2587 909
rect 2621 875 2659 909
rect 2693 875 2731 909
rect 2765 875 2803 909
rect 2837 875 2875 909
rect 2909 875 2947 909
rect 2981 875 3019 909
rect 3053 875 3091 909
rect 3125 875 3163 909
rect 3197 875 3235 909
rect 3269 875 3307 909
rect 3341 875 3379 909
rect 3413 875 3451 909
rect 3485 875 3523 909
rect 3557 875 3595 909
rect 3629 875 3667 909
rect 3701 875 3739 909
rect 3773 875 3811 909
rect 3845 875 3883 909
rect 3917 875 3955 909
rect 3989 875 4027 909
rect 4061 875 4099 909
rect 4133 875 4171 909
rect 4205 875 4243 909
rect 4277 875 4968 909
rect -210 838 4968 875
rect -208 836 4408 838
rect -208 655 -96 836
rect -8 744 64 748
rect -8 692 2 744
rect 54 692 64 744
rect -8 688 64 692
rect -208 621 -169 655
rect -135 621 -96 655
rect -208 583 -96 621
rect -208 549 -169 583
rect -135 549 -96 583
rect -208 511 -96 549
rect -208 477 -169 511
rect -135 477 -96 511
rect -208 439 -96 477
rect -208 405 -169 439
rect -135 405 -96 439
rect -208 367 -96 405
rect -208 333 -169 367
rect -135 333 -96 367
rect -208 295 -96 333
rect -208 261 -169 295
rect -135 261 -96 295
rect -208 223 -96 261
rect -208 189 -169 223
rect -135 189 -96 223
rect -208 151 -96 189
rect -208 117 -169 151
rect -135 117 -96 151
rect -208 79 -96 117
rect -208 45 -169 79
rect -135 45 -96 79
rect -208 7 -96 45
rect -208 -27 -169 7
rect -135 -27 -96 7
rect -208 -65 -96 -27
rect -208 -99 -169 -65
rect -135 -99 -96 -65
rect -208 -137 -96 -99
rect -208 -171 -169 -137
rect -135 -171 -96 -137
rect -208 -209 -96 -171
rect -208 -243 -169 -209
rect -135 -243 -96 -209
rect -208 -281 -96 -243
rect -208 -315 -169 -281
rect -135 -315 -96 -281
rect -208 -353 -96 -315
rect -208 -387 -169 -353
rect -135 -387 -96 -353
rect -208 -425 -96 -387
rect -208 -459 -169 -425
rect -135 -459 -96 -425
rect -208 -497 -96 -459
rect -208 -531 -169 -497
rect -135 -531 -96 -497
rect -208 -569 -96 -531
rect -208 -603 -169 -569
rect -135 -603 -96 -569
rect -208 -641 -96 -603
rect -208 -675 -169 -641
rect -135 -675 -96 -641
rect -208 -713 -96 -675
rect -208 -747 -169 -713
rect -135 -747 -96 -713
rect -208 -785 -96 -747
rect -208 -819 -169 -785
rect -135 -819 -96 -785
rect -208 -857 -96 -819
rect -208 -891 -169 -857
rect -135 -891 -96 -857
rect -208 -929 -96 -891
rect -208 -963 -169 -929
rect -135 -963 -96 -929
rect -208 -1001 -96 -963
rect -208 -1035 -169 -1001
rect -135 -1035 -96 -1001
rect -208 -1073 -96 -1035
rect -208 -1107 -169 -1073
rect -135 -1107 -96 -1073
rect -208 -1145 -96 -1107
rect -208 -1179 -169 -1145
rect -135 -1179 -96 -1145
rect -208 -1217 -96 -1179
rect -208 -1251 -169 -1217
rect -135 -1251 -96 -1217
rect -2 -1218 58 688
rect 136 620 208 624
rect 136 568 146 620
rect 198 568 208 620
rect 136 564 208 568
rect 272 620 332 836
rect 404 620 464 836
rect 784 744 856 748
rect 784 692 794 744
rect 846 692 856 744
rect 784 688 856 692
rect 142 -1092 202 564
rect 272 560 464 620
rect 272 -244 332 560
rect 404 478 464 560
rect 790 382 850 688
rect 1172 624 1232 836
rect 1304 624 1364 836
rect 1432 624 1492 836
rect 1172 564 1492 624
rect 1812 620 1884 624
rect 1812 568 1822 620
rect 1874 568 1884 620
rect 1812 564 1884 568
rect 2332 620 2404 624
rect 2332 568 2342 620
rect 2394 568 2404 620
rect 2332 564 2404 568
rect 2724 622 2784 836
rect 2856 622 2916 836
rect 2984 622 3044 836
rect 3360 744 3432 748
rect 3360 692 3370 744
rect 3422 692 3432 744
rect 3360 688 3432 692
rect 1172 480 1232 564
rect 1304 562 1492 564
rect 404 -244 464 6
rect 272 -304 464 -244
rect 272 -1090 332 -304
rect 404 -520 464 -304
rect 532 -358 592 80
rect 662 -110 722 4
rect 920 -108 980 0
rect 656 -114 728 -110
rect 656 -166 666 -114
rect 718 -166 728 -114
rect 656 -170 728 -166
rect 914 -112 986 -108
rect 914 -164 924 -112
rect 976 -164 986 -112
rect 914 -168 986 -164
rect 526 -362 598 -358
rect 526 -414 536 -362
rect 588 -414 598 -362
rect 526 -418 598 -414
rect 662 -520 722 -170
rect 784 -244 856 -240
rect 784 -296 794 -244
rect 846 -296 856 -244
rect 784 -300 856 -296
rect 790 -620 850 -300
rect 920 -518 980 -168
rect 1050 -358 1110 102
rect 1172 -242 1232 6
rect 1304 -242 1364 562
rect 1432 482 1492 562
rect 1818 386 1878 564
rect 2338 390 2398 564
rect 2724 562 3044 622
rect 2724 478 2784 562
rect 2856 560 3044 562
rect 1172 -244 1364 -242
rect 1434 -244 1494 6
rect 1564 -240 1624 104
rect 1692 -110 1752 2
rect 1952 -110 2012 4
rect 1686 -114 1758 -110
rect 1686 -166 1696 -114
rect 1748 -166 1758 -114
rect 1686 -170 1758 -166
rect 1946 -114 2018 -110
rect 1946 -166 1956 -114
rect 2008 -166 2018 -114
rect 1946 -170 2018 -166
rect 1172 -302 1494 -244
rect 1558 -244 1630 -240
rect 1558 -296 1568 -244
rect 1620 -296 1630 -244
rect 1558 -300 1630 -296
rect 1044 -362 1116 -358
rect 1044 -414 1054 -362
rect 1106 -414 1116 -362
rect 1044 -418 1116 -414
rect 1172 -518 1232 -302
rect 1304 -304 1494 -302
rect 398 -1090 458 -994
rect 136 -1096 208 -1092
rect 136 -1148 146 -1096
rect 198 -1148 208 -1096
rect 136 -1152 208 -1148
rect 272 -1150 458 -1090
rect 532 -1092 592 -902
rect 1048 -1092 1108 -910
rect 1170 -1092 1230 -992
rect 1304 -1092 1364 -304
rect 1434 -516 1494 -304
rect 1692 -522 1752 -170
rect 1816 -362 1888 -358
rect 1816 -414 1826 -362
rect 1878 -414 1888 -362
rect 1816 -418 1888 -414
rect 1822 -616 1882 -418
rect 1952 -522 2012 -170
rect 2080 -240 2140 110
rect 2208 -110 2268 8
rect 2466 -110 2526 10
rect 2202 -114 2274 -110
rect 2202 -166 2212 -114
rect 2264 -166 2274 -114
rect 2202 -170 2274 -166
rect 2460 -114 2532 -110
rect 2460 -166 2470 -114
rect 2522 -166 2532 -114
rect 2460 -170 2532 -166
rect 2074 -244 2146 -240
rect 2074 -296 2084 -244
rect 2136 -296 2146 -244
rect 2074 -300 2146 -296
rect 2208 -522 2268 -170
rect 2330 -362 2402 -358
rect 2330 -414 2340 -362
rect 2392 -414 2402 -362
rect 2330 -418 2402 -414
rect 2336 -616 2396 -418
rect 2466 -522 2526 -170
rect 2598 -240 2658 120
rect 2592 -244 2664 -240
rect 2592 -296 2602 -244
rect 2654 -296 2664 -244
rect 2592 -300 2664 -296
rect 2724 -244 2784 4
rect 2856 -244 2916 560
rect 2984 480 3044 560
rect 3366 370 3426 688
rect 3758 624 3818 836
rect 3882 624 3942 836
rect 4128 744 4200 748
rect 4128 692 4138 744
rect 4190 692 4200 744
rect 4128 688 4200 692
rect 3758 564 3942 624
rect 3992 620 4064 624
rect 3992 568 4002 620
rect 4054 568 4064 620
rect 3992 564 4064 568
rect 3758 480 3818 564
rect 2724 -246 2916 -244
rect 2986 -246 3046 4
rect 2724 -304 3046 -246
rect 2724 -520 2784 -304
rect 2856 -306 3046 -304
rect 1432 -1092 1492 -992
rect -208 -1289 -96 -1251
rect -8 -1222 64 -1218
rect -8 -1274 2 -1222
rect 54 -1274 64 -1222
rect -8 -1278 64 -1274
rect -208 -1323 -169 -1289
rect -135 -1323 -96 -1289
rect -208 -1361 -96 -1323
rect 272 -1352 332 -1150
rect 398 -1352 458 -1150
rect 526 -1096 598 -1092
rect 526 -1148 536 -1096
rect 588 -1148 598 -1096
rect 526 -1152 598 -1148
rect 1042 -1096 1114 -1092
rect 1042 -1148 1052 -1096
rect 1104 -1148 1114 -1096
rect 1042 -1152 1114 -1148
rect 1170 -1152 1492 -1092
rect 1170 -1352 1230 -1152
rect 1304 -1352 1364 -1152
rect 1432 -1352 1492 -1152
rect 1560 -1218 1620 -888
rect 2082 -1218 2142 -894
rect 2596 -1218 2656 -890
rect 2722 -1094 2782 -994
rect 2856 -1094 2916 -306
rect 2986 -518 3046 -306
rect 3112 -358 3172 126
rect 3242 -110 3302 -2
rect 3502 -110 3562 4
rect 3236 -114 3308 -110
rect 3236 -166 3246 -114
rect 3298 -166 3308 -114
rect 3236 -170 3308 -166
rect 3496 -114 3568 -110
rect 3496 -166 3506 -114
rect 3558 -166 3568 -114
rect 3496 -170 3568 -166
rect 3106 -362 3178 -358
rect 3106 -414 3116 -362
rect 3168 -414 3178 -362
rect 3106 -418 3178 -414
rect 3242 -520 3302 -170
rect 3362 -244 3434 -240
rect 3362 -296 3372 -244
rect 3424 -296 3434 -244
rect 3362 -300 3434 -296
rect 3368 -632 3428 -300
rect 3502 -520 3562 -170
rect 3626 -358 3686 102
rect 3754 -240 3814 4
rect 3882 -240 3942 564
rect 3754 -300 3942 -240
rect 3620 -362 3692 -358
rect 3620 -414 3630 -362
rect 3682 -414 3692 -362
rect 3620 -418 3692 -414
rect 3754 -518 3814 -300
rect 2984 -1094 3044 -994
rect 3112 -1092 3172 -902
rect 3626 -1092 3686 -906
rect 3752 -1092 3812 -992
rect 3882 -1092 3942 -300
rect 3998 -1092 4058 564
rect 2722 -1154 3044 -1094
rect 3106 -1096 3178 -1092
rect 3106 -1148 3116 -1096
rect 3168 -1148 3178 -1096
rect 3106 -1152 3178 -1148
rect 3620 -1096 3692 -1092
rect 3620 -1148 3630 -1096
rect 3682 -1148 3692 -1096
rect 3620 -1152 3692 -1148
rect 3752 -1152 3942 -1092
rect 3992 -1096 4064 -1092
rect 3992 -1148 4002 -1096
rect 4054 -1148 4064 -1096
rect 3992 -1152 4064 -1148
rect 1554 -1222 1626 -1218
rect 1554 -1274 1564 -1222
rect 1616 -1274 1626 -1222
rect 1554 -1278 1626 -1274
rect 2076 -1222 2148 -1218
rect 2076 -1274 2086 -1222
rect 2138 -1274 2148 -1222
rect 2076 -1278 2148 -1274
rect 2590 -1222 2662 -1218
rect 2590 -1274 2600 -1222
rect 2652 -1274 2662 -1222
rect 2590 -1278 2662 -1274
rect 2722 -1352 2782 -1154
rect 2856 -1352 2916 -1154
rect 2984 -1352 3044 -1154
rect 3752 -1352 3812 -1152
rect 3882 -1352 3942 -1152
rect 4134 -1218 4194 688
rect 4296 655 4408 836
rect 4296 621 4335 655
rect 4369 621 4408 655
rect 4296 583 4408 621
rect 4296 549 4335 583
rect 4369 549 4408 583
rect 4296 511 4408 549
rect 4296 477 4335 511
rect 4369 477 4408 511
rect 4296 439 4408 477
rect 4296 405 4335 439
rect 4369 405 4408 439
rect 4296 367 4408 405
rect 4296 333 4335 367
rect 4369 333 4408 367
rect 4296 295 4408 333
rect 4296 261 4335 295
rect 4369 261 4408 295
rect 4296 223 4408 261
rect 4296 189 4335 223
rect 4369 189 4408 223
rect 4296 151 4408 189
rect 4296 117 4335 151
rect 4369 117 4408 151
rect 4296 79 4408 117
rect 6942 104 7222 164
rect 4296 45 4335 79
rect 4369 45 4408 79
rect 4296 7 4408 45
rect 4296 -27 4335 7
rect 4369 -27 4408 7
rect 4296 -65 4408 -27
rect 4296 -99 4335 -65
rect 4369 -99 4408 -65
rect 4296 -137 4408 -99
rect 4296 -171 4335 -137
rect 4369 -171 4408 -137
rect 4296 -209 4408 -171
rect 4296 -243 4335 -209
rect 4369 -243 4408 -209
rect 4296 -281 4408 -243
rect 4296 -315 4335 -281
rect 4369 -315 4408 -281
rect 4296 -353 4408 -315
rect 4296 -387 4335 -353
rect 4369 -387 4408 -353
rect 4296 -425 4408 -387
rect 4296 -459 4335 -425
rect 4369 -459 4408 -425
rect 4296 -497 4408 -459
rect 4296 -531 4335 -497
rect 4369 -531 4408 -497
rect 4296 -569 4408 -531
rect 4296 -603 4335 -569
rect 4369 -603 4408 -569
rect 4296 -641 4408 -603
rect 4296 -675 4335 -641
rect 4369 -675 4408 -641
rect 4296 -713 4408 -675
rect 4296 -747 4335 -713
rect 4369 -747 4408 -713
rect 4296 -785 4408 -747
rect 4296 -819 4335 -785
rect 4369 -819 4408 -785
rect 4296 -857 4408 -819
rect 4296 -891 4335 -857
rect 4369 -891 4408 -857
rect 4296 -929 4408 -891
rect 4296 -963 4335 -929
rect 4369 -963 4408 -929
rect 4296 -1001 4408 -963
rect 4296 -1035 4335 -1001
rect 4369 -1035 4408 -1001
rect 4296 -1073 4408 -1035
rect 4296 -1107 4335 -1073
rect 4369 -1107 4408 -1073
rect 4296 -1145 4408 -1107
rect 4296 -1179 4335 -1145
rect 4369 -1179 4408 -1145
rect 4296 -1217 4408 -1179
rect 4128 -1222 4200 -1218
rect 4128 -1274 4138 -1222
rect 4190 -1274 4200 -1222
rect 4128 -1278 4200 -1274
rect 4296 -1251 4335 -1217
rect 4369 -1251 4408 -1217
rect 4296 -1289 4408 -1251
rect 4296 -1323 4335 -1289
rect 4369 -1323 4408 -1289
rect -208 -1395 -169 -1361
rect -135 -1395 -96 -1361
rect -208 -1433 -96 -1395
rect -208 -1467 -169 -1433
rect -135 -1467 -96 -1433
rect -208 -1505 -96 -1467
rect -208 -1539 -169 -1505
rect -135 -1539 -96 -1505
rect -208 -1577 -96 -1539
rect 204 -1428 3996 -1352
rect 204 -1480 286 -1428
rect 338 -1480 350 -1428
rect 402 -1480 414 -1428
rect 466 -1480 478 -1428
rect 530 -1480 542 -1428
rect 594 -1480 606 -1428
rect 658 -1480 670 -1428
rect 722 -1480 734 -1428
rect 786 -1480 798 -1428
rect 850 -1480 862 -1428
rect 914 -1480 926 -1428
rect 978 -1480 990 -1428
rect 1042 -1480 1054 -1428
rect 1106 -1480 1118 -1428
rect 1170 -1480 1182 -1428
rect 1234 -1480 1246 -1428
rect 1298 -1480 1310 -1428
rect 1362 -1480 1374 -1428
rect 1426 -1480 1438 -1428
rect 1490 -1480 1502 -1428
rect 1554 -1480 1566 -1428
rect 1618 -1480 1630 -1428
rect 1682 -1480 1694 -1428
rect 1746 -1480 1758 -1428
rect 1810 -1480 1822 -1428
rect 1874 -1480 1886 -1428
rect 1938 -1480 1950 -1428
rect 2002 -1480 2014 -1428
rect 2066 -1480 2078 -1428
rect 2130 -1480 2142 -1428
rect 2194 -1480 2206 -1428
rect 2258 -1480 2270 -1428
rect 2322 -1480 2334 -1428
rect 2386 -1480 2398 -1428
rect 2450 -1480 2462 -1428
rect 2514 -1480 2526 -1428
rect 2578 -1480 2590 -1428
rect 2642 -1480 2654 -1428
rect 2706 -1480 2718 -1428
rect 2770 -1480 2782 -1428
rect 2834 -1480 2846 -1428
rect 2898 -1480 2910 -1428
rect 2962 -1480 2974 -1428
rect 3026 -1480 3038 -1428
rect 3090 -1480 3102 -1428
rect 3154 -1480 3166 -1428
rect 3218 -1480 3230 -1428
rect 3282 -1480 3294 -1428
rect 3346 -1480 3358 -1428
rect 3410 -1480 3422 -1428
rect 3474 -1480 3486 -1428
rect 3538 -1480 3550 -1428
rect 3602 -1480 3614 -1428
rect 3666 -1480 3678 -1428
rect 3730 -1480 3742 -1428
rect 3794 -1480 3806 -1428
rect 3858 -1480 3870 -1428
rect 3922 -1480 3996 -1428
rect 204 -1550 3996 -1480
rect 4296 -1361 4408 -1323
rect 4296 -1395 4335 -1361
rect 4369 -1395 4408 -1361
rect 4296 -1433 4408 -1395
rect 4296 -1467 4335 -1433
rect 4369 -1467 4408 -1433
rect 4296 -1505 4408 -1467
rect 4296 -1539 4335 -1505
rect 4369 -1539 4408 -1505
rect -208 -1611 -169 -1577
rect -135 -1611 -96 -1577
rect -208 -1636 -96 -1611
rect 4296 -1577 4408 -1539
rect 4296 -1611 4335 -1577
rect 4369 -1611 4408 -1577
rect 4296 -1636 4408 -1611
rect -208 -1649 514 -1636
rect -208 -1683 -169 -1649
rect -135 -1664 514 -1649
rect -135 -1683 -78 -1664
rect -208 -1721 -78 -1683
rect -208 -1755 -169 -1721
rect -135 -1755 -78 -1721
rect -208 -1908 -78 -1755
rect 486 -1908 514 -1664
rect -208 -1936 514 -1908
rect 3686 -1649 4408 -1636
rect 3686 -1664 4335 -1649
rect 3686 -1908 3714 -1664
rect 4278 -1683 4335 -1664
rect 4369 -1683 4408 -1649
rect 4278 -1721 4408 -1683
rect 4278 -1755 4335 -1721
rect 4369 -1755 4408 -1721
rect 4278 -1908 4408 -1755
rect 3686 -1936 4408 -1908
rect -208 -1975 4408 -1936
rect -208 -2009 -77 -1975
rect -43 -2009 -5 -1975
rect 29 -2009 67 -1975
rect 101 -2009 139 -1975
rect 173 -2009 211 -1975
rect 245 -2009 283 -1975
rect 317 -2009 355 -1975
rect 389 -2009 427 -1975
rect 461 -2009 499 -1975
rect 533 -2009 571 -1975
rect 605 -2009 643 -1975
rect 677 -2009 715 -1975
rect 749 -2009 787 -1975
rect 821 -2009 859 -1975
rect 893 -2009 931 -1975
rect 965 -2009 1003 -1975
rect 1037 -2009 1075 -1975
rect 1109 -2009 1147 -1975
rect 1181 -2009 1219 -1975
rect 1253 -2009 1291 -1975
rect 1325 -2009 1363 -1975
rect 1397 -2009 1435 -1975
rect 1469 -2009 1507 -1975
rect 1541 -2009 1579 -1975
rect 1613 -2009 1651 -1975
rect 1685 -2009 1723 -1975
rect 1757 -2009 1795 -1975
rect 1829 -2009 1867 -1975
rect 1901 -2009 1939 -1975
rect 1973 -2009 2011 -1975
rect 2045 -2009 2083 -1975
rect 2117 -2009 2155 -1975
rect 2189 -2009 2227 -1975
rect 2261 -2009 2299 -1975
rect 2333 -2009 2371 -1975
rect 2405 -2009 2443 -1975
rect 2477 -2009 2515 -1975
rect 2549 -2009 2587 -1975
rect 2621 -2009 2659 -1975
rect 2693 -2009 2731 -1975
rect 2765 -2009 2803 -1975
rect 2837 -2009 2875 -1975
rect 2909 -2009 2947 -1975
rect 2981 -2009 3019 -1975
rect 3053 -2009 3091 -1975
rect 3125 -2009 3163 -1975
rect 3197 -2009 3235 -1975
rect 3269 -2009 3307 -1975
rect 3341 -2009 3379 -1975
rect 3413 -2009 3451 -1975
rect 3485 -2009 3523 -1975
rect 3557 -2009 3595 -1975
rect 3629 -2009 3667 -1975
rect 3701 -2009 3739 -1975
rect 3773 -2009 3811 -1975
rect 3845 -2009 3883 -1975
rect 3917 -2009 3955 -1975
rect 3989 -2009 4027 -1975
rect 4061 -2009 4099 -1975
rect 4133 -2009 4171 -1975
rect 4205 -2009 4243 -1975
rect 4277 -2009 4408 -1975
rect -208 -2048 4408 -2009
<< via1 >>
rect 4711 1208 4955 12780
rect -138 915 -86 967
rect -74 915 -22 967
rect -10 915 42 967
rect 54 915 106 967
rect 118 915 170 967
rect 182 915 234 967
rect 246 915 298 967
rect 310 915 362 967
rect 374 915 426 967
rect 438 915 490 967
rect 502 915 554 967
rect 566 915 618 967
rect 630 915 682 967
rect 694 915 746 967
rect 758 915 810 967
rect 822 915 874 967
rect 886 915 938 967
rect 950 915 1002 967
rect 1014 915 1066 967
rect 1078 915 1130 967
rect 1142 915 1194 967
rect 1206 915 1258 967
rect 1270 915 1322 967
rect 1334 915 1386 967
rect 1398 915 1450 967
rect 1462 915 1514 967
rect 1526 915 1578 967
rect 1590 915 1642 967
rect 1654 915 1706 967
rect 1718 915 1770 967
rect 1782 915 1834 967
rect 1846 915 1898 967
rect 1910 915 1962 967
rect 1974 915 2026 967
rect 2038 915 2090 967
rect 2102 915 2154 967
rect 2166 915 2218 967
rect 2230 915 2282 967
rect 2294 915 2346 967
rect 2358 915 2410 967
rect 2422 915 2474 967
rect 2486 915 2538 967
rect 2550 915 2602 967
rect 2614 915 2666 967
rect 2678 915 2730 967
rect 2742 915 2794 967
rect 2806 915 2858 967
rect 2870 915 2922 967
rect 2934 915 2986 967
rect 2998 915 3050 967
rect 3062 915 3114 967
rect 3126 915 3178 967
rect 3190 915 3242 967
rect 3254 915 3306 967
rect 3318 915 3370 967
rect 3382 915 3434 967
rect 3446 915 3498 967
rect 3510 915 3562 967
rect 3574 915 3626 967
rect 3638 915 3690 967
rect 3702 915 3754 967
rect 3766 915 3818 967
rect 3830 915 3882 967
rect 3894 915 3946 967
rect 3958 915 4010 967
rect 4022 915 4074 967
rect 4086 915 4138 967
rect 4150 915 4202 967
rect 4214 915 4266 967
rect 4278 915 4330 967
rect 4342 915 4394 967
rect 4406 915 4458 967
rect 4470 915 4522 967
rect 4534 915 4586 967
rect 4598 915 4650 967
rect 4662 915 4714 967
rect 4726 915 4778 967
rect 4790 915 4842 967
rect 4854 915 4906 967
rect 2 692 54 744
rect 146 568 198 620
rect 794 692 846 744
rect 1822 568 1874 620
rect 2342 568 2394 620
rect 3370 692 3422 744
rect 666 -166 718 -114
rect 924 -164 976 -112
rect 536 -414 588 -362
rect 794 -296 846 -244
rect 1696 -166 1748 -114
rect 1956 -166 2008 -114
rect 1568 -296 1620 -244
rect 1054 -414 1106 -362
rect 146 -1148 198 -1096
rect 1826 -414 1878 -362
rect 2212 -166 2264 -114
rect 2470 -166 2522 -114
rect 2084 -296 2136 -244
rect 2340 -414 2392 -362
rect 2602 -296 2654 -244
rect 4138 692 4190 744
rect 4002 568 4054 620
rect 2 -1274 54 -1222
rect 536 -1148 588 -1096
rect 1052 -1148 1104 -1096
rect 3246 -166 3298 -114
rect 3506 -166 3558 -114
rect 3116 -414 3168 -362
rect 3372 -296 3424 -244
rect 3630 -414 3682 -362
rect 3116 -1148 3168 -1096
rect 3630 -1148 3682 -1096
rect 4002 -1148 4054 -1096
rect 1564 -1274 1616 -1222
rect 2086 -1274 2138 -1222
rect 2600 -1274 2652 -1222
rect 4138 -1274 4190 -1222
rect 286 -1480 338 -1428
rect 350 -1480 402 -1428
rect 414 -1480 466 -1428
rect 478 -1480 530 -1428
rect 542 -1480 594 -1428
rect 606 -1480 658 -1428
rect 670 -1480 722 -1428
rect 734 -1480 786 -1428
rect 798 -1480 850 -1428
rect 862 -1480 914 -1428
rect 926 -1480 978 -1428
rect 990 -1480 1042 -1428
rect 1054 -1480 1106 -1428
rect 1118 -1480 1170 -1428
rect 1182 -1480 1234 -1428
rect 1246 -1480 1298 -1428
rect 1310 -1480 1362 -1428
rect 1374 -1480 1426 -1428
rect 1438 -1480 1490 -1428
rect 1502 -1480 1554 -1428
rect 1566 -1480 1618 -1428
rect 1630 -1480 1682 -1428
rect 1694 -1480 1746 -1428
rect 1758 -1480 1810 -1428
rect 1822 -1480 1874 -1428
rect 1886 -1480 1938 -1428
rect 1950 -1480 2002 -1428
rect 2014 -1480 2066 -1428
rect 2078 -1480 2130 -1428
rect 2142 -1480 2194 -1428
rect 2206 -1480 2258 -1428
rect 2270 -1480 2322 -1428
rect 2334 -1480 2386 -1428
rect 2398 -1480 2450 -1428
rect 2462 -1480 2514 -1428
rect 2526 -1480 2578 -1428
rect 2590 -1480 2642 -1428
rect 2654 -1480 2706 -1428
rect 2718 -1480 2770 -1428
rect 2782 -1480 2834 -1428
rect 2846 -1480 2898 -1428
rect 2910 -1480 2962 -1428
rect 2974 -1480 3026 -1428
rect 3038 -1480 3090 -1428
rect 3102 -1480 3154 -1428
rect 3166 -1480 3218 -1428
rect 3230 -1480 3282 -1428
rect 3294 -1480 3346 -1428
rect 3358 -1480 3410 -1428
rect 3422 -1480 3474 -1428
rect 3486 -1480 3538 -1428
rect 3550 -1480 3602 -1428
rect 3614 -1480 3666 -1428
rect 3678 -1480 3730 -1428
rect 3742 -1480 3794 -1428
rect 3806 -1480 3858 -1428
rect 3870 -1480 3922 -1428
rect -78 -1908 486 -1664
rect 3714 -1908 4278 -1664
<< metal2 >>
rect 4216 12972 5348 13072
rect 1875 12090 1965 12094
rect 4216 12090 4316 12972
rect 1870 12068 4316 12090
rect 1870 12012 1892 12068
rect 1948 12012 4316 12068
rect 1870 11990 4316 12012
rect 4636 12782 5024 12860
rect 4636 12780 4725 12782
rect 4941 12780 5024 12782
rect 1875 11986 1965 11990
rect 1574 9681 1676 9686
rect 1570 9663 1680 9681
rect 1570 9607 1597 9663
rect 1653 9607 1680 9663
rect 1570 9589 1680 9607
rect 1574 9539 1676 9589
rect 919 9437 1676 9539
rect 919 9364 1021 9437
rect 919 9308 942 9364
rect 998 9308 1021 9364
rect 919 9276 1021 9308
rect 1286 4681 1390 4686
rect 1282 4662 1394 4681
rect 1282 4606 1310 4662
rect 1366 4606 1394 4662
rect 1282 4587 1394 4606
rect 1286 4532 1390 4587
rect 1286 4428 1746 4532
rect 1642 4342 1746 4428
rect 1642 4286 1666 4342
rect 1722 4286 1746 4342
rect 1642 4253 1746 4286
rect 4636 1208 4711 12780
rect 4955 1208 5024 12780
rect 5248 12762 5348 12972
rect 5248 12706 5270 12762
rect 5326 12706 5348 12762
rect 5248 12675 5348 12706
rect 4636 1206 4725 1208
rect 4941 1206 5024 1208
rect 4636 1148 5024 1206
rect 5564 1602 8252 1662
rect -202 969 4964 1026
rect -202 967 -124 969
rect -68 967 -44 969
rect 12 967 36 969
rect 92 967 116 969
rect 172 967 196 969
rect 252 967 276 969
rect 332 967 356 969
rect 412 967 436 969
rect 492 967 516 969
rect 572 967 596 969
rect 652 967 676 969
rect 732 967 756 969
rect 812 967 836 969
rect 892 967 916 969
rect 972 967 996 969
rect 1052 967 1076 969
rect 1132 967 1156 969
rect 1212 967 1236 969
rect 1292 967 1316 969
rect 1372 967 1396 969
rect 1452 967 1476 969
rect 1532 967 1556 969
rect 1612 967 1636 969
rect 1692 967 1716 969
rect 1772 967 1796 969
rect 1852 967 1876 969
rect 1932 967 1956 969
rect 2012 967 2036 969
rect 2092 967 2116 969
rect 2172 967 2196 969
rect 2252 967 2276 969
rect 2332 967 2356 969
rect 2412 967 2436 969
rect 2492 967 2516 969
rect 2572 967 2596 969
rect 2652 967 2676 969
rect 2732 967 2756 969
rect 2812 967 2836 969
rect 2892 967 2916 969
rect 2972 967 2996 969
rect 3052 967 3076 969
rect 3132 967 3156 969
rect 3212 967 3236 969
rect 3292 967 3316 969
rect 3372 967 3396 969
rect 3452 967 3476 969
rect 3532 967 3556 969
rect 3612 967 3636 969
rect 3692 967 3716 969
rect 3772 967 3796 969
rect 3852 967 3876 969
rect 3932 967 3956 969
rect 4012 967 4036 969
rect 4092 967 4116 969
rect 4172 967 4196 969
rect 4252 967 4276 969
rect 4332 967 4356 969
rect 4412 967 4436 969
rect 4492 967 4516 969
rect 4572 967 4596 969
rect 4652 967 4676 969
rect 4732 967 4756 969
rect 4812 967 4836 969
rect 4892 967 4964 969
rect -202 915 -138 967
rect 106 915 116 967
rect 172 915 182 967
rect 426 915 436 967
rect 492 915 502 967
rect 746 915 756 967
rect 812 915 822 967
rect 1066 915 1076 967
rect 1132 915 1142 967
rect 1386 915 1396 967
rect 1452 915 1462 967
rect 1706 915 1716 967
rect 1772 915 1782 967
rect 2026 915 2036 967
rect 2092 915 2102 967
rect 2346 915 2356 967
rect 2412 915 2422 967
rect 2666 915 2676 967
rect 2732 915 2742 967
rect 2986 915 2996 967
rect 3052 915 3062 967
rect 3306 915 3316 967
rect 3372 915 3382 967
rect 3626 915 3636 967
rect 3692 915 3702 967
rect 3946 915 3956 967
rect 4012 915 4022 967
rect 4266 915 4276 967
rect 4332 915 4342 967
rect 4586 915 4596 967
rect 4652 915 4662 967
rect 4906 915 4964 967
rect -202 913 -124 915
rect -68 913 -44 915
rect 12 913 36 915
rect 92 913 116 915
rect 172 913 196 915
rect 252 913 276 915
rect 332 913 356 915
rect 412 913 436 915
rect 492 913 516 915
rect 572 913 596 915
rect 652 913 676 915
rect 732 913 756 915
rect 812 913 836 915
rect 892 913 916 915
rect 972 913 996 915
rect 1052 913 1076 915
rect 1132 913 1156 915
rect 1212 913 1236 915
rect 1292 913 1316 915
rect 1372 913 1396 915
rect 1452 913 1476 915
rect 1532 913 1556 915
rect 1612 913 1636 915
rect 1692 913 1716 915
rect 1772 913 1796 915
rect 1852 913 1876 915
rect 1932 913 1956 915
rect 2012 913 2036 915
rect 2092 913 2116 915
rect 2172 913 2196 915
rect 2252 913 2276 915
rect 2332 913 2356 915
rect 2412 913 2436 915
rect 2492 913 2516 915
rect 2572 913 2596 915
rect 2652 913 2676 915
rect 2732 913 2756 915
rect 2812 913 2836 915
rect 2892 913 2916 915
rect 2972 913 2996 915
rect 3052 913 3076 915
rect 3132 913 3156 915
rect 3212 913 3236 915
rect 3292 913 3316 915
rect 3372 913 3396 915
rect 3452 913 3476 915
rect 3532 913 3556 915
rect 3612 913 3636 915
rect 3692 913 3716 915
rect 3772 913 3796 915
rect 3852 913 3876 915
rect 3932 913 3956 915
rect 4012 913 4036 915
rect 4092 913 4116 915
rect 4172 913 4196 915
rect 4252 913 4276 915
rect 4332 913 4356 915
rect 4412 913 4436 915
rect 4492 913 4516 915
rect 4572 913 4596 915
rect 4652 913 4676 915
rect 4732 913 4756 915
rect 4812 913 4836 915
rect 4892 913 4964 915
rect -202 846 4964 913
rect -2 748 58 754
rect 790 748 850 754
rect 3366 748 3426 754
rect 4134 748 4194 754
rect -2 744 4194 748
rect -2 692 2 744
rect 54 692 794 744
rect 846 692 3370 744
rect 3422 692 4138 744
rect 4190 692 4194 744
rect -2 688 4194 692
rect -2 682 58 688
rect 790 682 850 688
rect 3366 682 3426 688
rect 4134 682 4194 688
rect 142 624 202 630
rect 1033 624 1123 648
rect 1818 624 1878 630
rect 2338 624 2398 630
rect 3998 624 4058 630
rect 5564 624 5624 1602
rect 6398 640 6596 700
rect 6391 634 6508 640
rect 142 622 5624 624
rect 142 620 1050 622
rect 142 568 146 620
rect 198 568 1050 620
rect 142 566 1050 568
rect 1106 620 5624 622
rect 1106 568 1822 620
rect 1874 568 2342 620
rect 2394 568 4002 620
rect 4054 568 5624 620
rect 1106 566 5624 568
rect 142 564 5624 566
rect 142 558 202 564
rect 1033 540 1123 564
rect 1818 558 1878 564
rect 2338 558 2398 564
rect 3998 558 4058 564
rect 662 -110 722 -104
rect 920 -110 980 -102
rect 1692 -110 1752 -104
rect 1952 -110 2012 -104
rect 2208 -110 2268 -104
rect 2466 -110 2526 -104
rect 3242 -110 3302 -104
rect 3502 -110 3562 -104
rect 662 -112 3562 -110
rect 662 -114 924 -112
rect 662 -166 666 -114
rect 718 -164 924 -114
rect 976 -114 3562 -112
rect 976 -164 1696 -114
rect 718 -166 1696 -164
rect 1748 -166 1956 -114
rect 2008 -166 2212 -114
rect 2264 -166 2470 -114
rect 2522 -166 3246 -114
rect 3298 -166 3506 -114
rect 3558 -166 3562 -114
rect 662 -170 3562 -166
rect 662 -176 722 -170
rect 920 -174 980 -170
rect 1692 -176 1752 -170
rect 1952 -176 2012 -170
rect 2208 -176 2268 -170
rect 2466 -176 2526 -170
rect 3242 -176 3302 -170
rect 3502 -176 3562 -170
rect 790 -240 850 -234
rect 1564 -240 1624 -234
rect 2080 -240 2140 -234
rect 2598 -240 2658 -234
rect 3368 -240 3428 -234
rect 790 -242 5181 -240
rect 790 -244 5114 -242
rect 790 -296 794 -244
rect 846 -296 1568 -244
rect 1620 -296 2084 -244
rect 2136 -296 2602 -244
rect 2654 -296 3372 -244
rect 3424 -296 5114 -244
rect 790 -298 5114 -296
rect 5170 -298 5181 -242
rect 790 -300 5181 -298
rect 790 -306 850 -300
rect 1564 -306 1624 -300
rect 2080 -306 2140 -300
rect 2598 -306 2658 -300
rect 3368 -306 3428 -300
rect 532 -358 592 -352
rect 1050 -358 1110 -352
rect 1822 -358 1882 -352
rect 2336 -358 2396 -352
rect 3112 -358 3172 -352
rect 3607 -358 3697 -332
rect 6448 -358 6508 634
rect 532 -362 3624 -358
rect 3680 -362 6508 -358
rect 532 -414 536 -362
rect 588 -414 1054 -362
rect 1106 -414 1826 -362
rect 1878 -414 2340 -362
rect 2392 -414 3116 -362
rect 3168 -414 3624 -362
rect 3682 -414 6508 -362
rect 532 -418 6508 -414
rect 532 -424 592 -418
rect 1050 -424 1110 -418
rect 1822 -424 1882 -418
rect 2336 -424 2396 -418
rect 3112 -424 3172 -418
rect 3607 -440 3697 -418
rect 142 -1092 202 -1086
rect 532 -1092 592 -1086
rect 1048 -1092 1108 -1086
rect 3112 -1092 3172 -1086
rect 3626 -1092 3686 -1086
rect 3998 -1092 4058 -1086
rect 142 -1096 4058 -1092
rect 142 -1148 146 -1096
rect 198 -1148 536 -1096
rect 588 -1148 1052 -1096
rect 1104 -1148 3116 -1096
rect 3168 -1148 3630 -1096
rect 3682 -1148 4002 -1096
rect 4054 -1148 4058 -1096
rect 142 -1152 4058 -1148
rect 142 -1158 202 -1152
rect 532 -1158 592 -1152
rect 1048 -1158 1108 -1152
rect 3112 -1158 3172 -1152
rect 3626 -1158 3686 -1152
rect 3998 -1158 4058 -1152
rect -2 -1218 58 -1212
rect 1560 -1218 1620 -1212
rect 2082 -1218 2142 -1212
rect 2596 -1218 2656 -1212
rect 4134 -1218 4194 -1212
rect -2 -1222 4194 -1218
rect -2 -1274 2 -1222
rect 54 -1274 1564 -1222
rect 1616 -1274 2086 -1222
rect 2138 -1274 2600 -1222
rect 2652 -1274 4138 -1222
rect 4190 -1274 4194 -1222
rect -2 -1278 4194 -1274
rect -2 -1284 58 -1278
rect 1560 -1284 1620 -1278
rect 2082 -1284 2142 -1278
rect 2596 -1284 2656 -1278
rect 4134 -1284 4194 -1278
rect 204 -1426 3996 -1352
rect 204 -1482 276 -1426
rect 332 -1428 356 -1426
rect 412 -1428 436 -1426
rect 492 -1428 516 -1426
rect 572 -1428 596 -1426
rect 652 -1428 676 -1426
rect 732 -1428 756 -1426
rect 812 -1428 836 -1426
rect 892 -1428 916 -1426
rect 972 -1428 996 -1426
rect 1052 -1428 1076 -1426
rect 1132 -1428 1156 -1426
rect 1212 -1428 1236 -1426
rect 1292 -1428 1316 -1426
rect 1372 -1428 1396 -1426
rect 1452 -1428 1476 -1426
rect 1532 -1428 1556 -1426
rect 1612 -1428 1636 -1426
rect 1692 -1428 1716 -1426
rect 1772 -1428 1796 -1426
rect 1852 -1428 1876 -1426
rect 1932 -1428 1956 -1426
rect 2012 -1428 2036 -1426
rect 2092 -1428 2116 -1426
rect 2172 -1428 2196 -1426
rect 2252 -1428 2276 -1426
rect 2332 -1428 2356 -1426
rect 2412 -1428 2436 -1426
rect 2492 -1428 2516 -1426
rect 2572 -1428 2596 -1426
rect 2652 -1428 2676 -1426
rect 2732 -1428 2756 -1426
rect 2812 -1428 2836 -1426
rect 2892 -1428 2916 -1426
rect 2972 -1428 2996 -1426
rect 3052 -1428 3076 -1426
rect 3132 -1428 3156 -1426
rect 3212 -1428 3236 -1426
rect 3292 -1428 3316 -1426
rect 3372 -1428 3396 -1426
rect 3452 -1428 3476 -1426
rect 3532 -1428 3556 -1426
rect 3612 -1428 3636 -1426
rect 3692 -1428 3716 -1426
rect 3772 -1428 3796 -1426
rect 3852 -1428 3876 -1426
rect 338 -1480 350 -1428
rect 412 -1480 414 -1428
rect 594 -1480 596 -1428
rect 658 -1480 670 -1428
rect 732 -1480 734 -1428
rect 914 -1480 916 -1428
rect 978 -1480 990 -1428
rect 1052 -1480 1054 -1428
rect 1234 -1480 1236 -1428
rect 1298 -1480 1310 -1428
rect 1372 -1480 1374 -1428
rect 1554 -1480 1556 -1428
rect 1618 -1480 1630 -1428
rect 1692 -1480 1694 -1428
rect 1874 -1480 1876 -1428
rect 1938 -1480 1950 -1428
rect 2012 -1480 2014 -1428
rect 2194 -1480 2196 -1428
rect 2258 -1480 2270 -1428
rect 2332 -1480 2334 -1428
rect 2514 -1480 2516 -1428
rect 2578 -1480 2590 -1428
rect 2652 -1480 2654 -1428
rect 2834 -1480 2836 -1428
rect 2898 -1480 2910 -1428
rect 2972 -1480 2974 -1428
rect 3154 -1480 3156 -1428
rect 3218 -1480 3230 -1428
rect 3292 -1480 3294 -1428
rect 3474 -1480 3476 -1428
rect 3538 -1480 3550 -1428
rect 3612 -1480 3614 -1428
rect 3794 -1480 3796 -1428
rect 3858 -1480 3870 -1428
rect 332 -1482 356 -1480
rect 412 -1482 436 -1480
rect 492 -1482 516 -1480
rect 572 -1482 596 -1480
rect 652 -1482 676 -1480
rect 732 -1482 756 -1480
rect 812 -1482 836 -1480
rect 892 -1482 916 -1480
rect 972 -1482 996 -1480
rect 1052 -1482 1076 -1480
rect 1132 -1482 1156 -1480
rect 1212 -1482 1236 -1480
rect 1292 -1482 1316 -1480
rect 1372 -1482 1396 -1480
rect 1452 -1482 1476 -1480
rect 1532 -1482 1556 -1480
rect 1612 -1482 1636 -1480
rect 1692 -1482 1716 -1480
rect 1772 -1482 1796 -1480
rect 1852 -1482 1876 -1480
rect 1932 -1482 1956 -1480
rect 2012 -1482 2036 -1480
rect 2092 -1482 2116 -1480
rect 2172 -1482 2196 -1480
rect 2252 -1482 2276 -1480
rect 2332 -1482 2356 -1480
rect 2412 -1482 2436 -1480
rect 2492 -1482 2516 -1480
rect 2572 -1482 2596 -1480
rect 2652 -1482 2676 -1480
rect 2732 -1482 2756 -1480
rect 2812 -1482 2836 -1480
rect 2892 -1482 2916 -1480
rect 2972 -1482 2996 -1480
rect 3052 -1482 3076 -1480
rect 3132 -1482 3156 -1480
rect 3212 -1482 3236 -1480
rect 3292 -1482 3316 -1480
rect 3372 -1482 3396 -1480
rect 3452 -1482 3476 -1480
rect 3532 -1482 3556 -1480
rect 3612 -1482 3636 -1480
rect 3692 -1482 3716 -1480
rect 3772 -1482 3796 -1480
rect 3852 -1482 3876 -1480
rect 3932 -1482 3996 -1426
rect 204 -1550 3996 -1482
rect -96 -1638 504 -1626
rect -96 -1664 -64 -1638
rect 472 -1664 504 -1638
rect -96 -1908 -78 -1664
rect 486 -1908 504 -1664
rect -96 -1934 -64 -1908
rect 472 -1934 504 -1908
rect -96 -1946 504 -1934
rect 3696 -1638 4296 -1626
rect 3696 -1664 3728 -1638
rect 4264 -1664 4296 -1638
rect 3696 -1908 3714 -1664
rect 4278 -1908 4296 -1664
rect 3696 -1934 3728 -1908
rect 4264 -1934 4296 -1908
rect 3696 -1946 4296 -1934
<< via2 >>
rect 1892 12012 1948 12068
rect 4725 12780 4941 12782
rect 1597 9607 1653 9663
rect 942 9308 998 9364
rect 1310 4606 1366 4662
rect 1666 4286 1722 4342
rect 4725 1208 4941 12780
rect 5270 12706 5326 12762
rect 4725 1206 4941 1208
rect -124 967 -68 969
rect -44 967 12 969
rect 36 967 92 969
rect 116 967 172 969
rect 196 967 252 969
rect 276 967 332 969
rect 356 967 412 969
rect 436 967 492 969
rect 516 967 572 969
rect 596 967 652 969
rect 676 967 732 969
rect 756 967 812 969
rect 836 967 892 969
rect 916 967 972 969
rect 996 967 1052 969
rect 1076 967 1132 969
rect 1156 967 1212 969
rect 1236 967 1292 969
rect 1316 967 1372 969
rect 1396 967 1452 969
rect 1476 967 1532 969
rect 1556 967 1612 969
rect 1636 967 1692 969
rect 1716 967 1772 969
rect 1796 967 1852 969
rect 1876 967 1932 969
rect 1956 967 2012 969
rect 2036 967 2092 969
rect 2116 967 2172 969
rect 2196 967 2252 969
rect 2276 967 2332 969
rect 2356 967 2412 969
rect 2436 967 2492 969
rect 2516 967 2572 969
rect 2596 967 2652 969
rect 2676 967 2732 969
rect 2756 967 2812 969
rect 2836 967 2892 969
rect 2916 967 2972 969
rect 2996 967 3052 969
rect 3076 967 3132 969
rect 3156 967 3212 969
rect 3236 967 3292 969
rect 3316 967 3372 969
rect 3396 967 3452 969
rect 3476 967 3532 969
rect 3556 967 3612 969
rect 3636 967 3692 969
rect 3716 967 3772 969
rect 3796 967 3852 969
rect 3876 967 3932 969
rect 3956 967 4012 969
rect 4036 967 4092 969
rect 4116 967 4172 969
rect 4196 967 4252 969
rect 4276 967 4332 969
rect 4356 967 4412 969
rect 4436 967 4492 969
rect 4516 967 4572 969
rect 4596 967 4652 969
rect 4676 967 4732 969
rect 4756 967 4812 969
rect 4836 967 4892 969
rect -124 915 -86 967
rect -86 915 -74 967
rect -74 915 -68 967
rect -44 915 -22 967
rect -22 915 -10 967
rect -10 915 12 967
rect 36 915 42 967
rect 42 915 54 967
rect 54 915 92 967
rect 116 915 118 967
rect 118 915 170 967
rect 170 915 172 967
rect 196 915 234 967
rect 234 915 246 967
rect 246 915 252 967
rect 276 915 298 967
rect 298 915 310 967
rect 310 915 332 967
rect 356 915 362 967
rect 362 915 374 967
rect 374 915 412 967
rect 436 915 438 967
rect 438 915 490 967
rect 490 915 492 967
rect 516 915 554 967
rect 554 915 566 967
rect 566 915 572 967
rect 596 915 618 967
rect 618 915 630 967
rect 630 915 652 967
rect 676 915 682 967
rect 682 915 694 967
rect 694 915 732 967
rect 756 915 758 967
rect 758 915 810 967
rect 810 915 812 967
rect 836 915 874 967
rect 874 915 886 967
rect 886 915 892 967
rect 916 915 938 967
rect 938 915 950 967
rect 950 915 972 967
rect 996 915 1002 967
rect 1002 915 1014 967
rect 1014 915 1052 967
rect 1076 915 1078 967
rect 1078 915 1130 967
rect 1130 915 1132 967
rect 1156 915 1194 967
rect 1194 915 1206 967
rect 1206 915 1212 967
rect 1236 915 1258 967
rect 1258 915 1270 967
rect 1270 915 1292 967
rect 1316 915 1322 967
rect 1322 915 1334 967
rect 1334 915 1372 967
rect 1396 915 1398 967
rect 1398 915 1450 967
rect 1450 915 1452 967
rect 1476 915 1514 967
rect 1514 915 1526 967
rect 1526 915 1532 967
rect 1556 915 1578 967
rect 1578 915 1590 967
rect 1590 915 1612 967
rect 1636 915 1642 967
rect 1642 915 1654 967
rect 1654 915 1692 967
rect 1716 915 1718 967
rect 1718 915 1770 967
rect 1770 915 1772 967
rect 1796 915 1834 967
rect 1834 915 1846 967
rect 1846 915 1852 967
rect 1876 915 1898 967
rect 1898 915 1910 967
rect 1910 915 1932 967
rect 1956 915 1962 967
rect 1962 915 1974 967
rect 1974 915 2012 967
rect 2036 915 2038 967
rect 2038 915 2090 967
rect 2090 915 2092 967
rect 2116 915 2154 967
rect 2154 915 2166 967
rect 2166 915 2172 967
rect 2196 915 2218 967
rect 2218 915 2230 967
rect 2230 915 2252 967
rect 2276 915 2282 967
rect 2282 915 2294 967
rect 2294 915 2332 967
rect 2356 915 2358 967
rect 2358 915 2410 967
rect 2410 915 2412 967
rect 2436 915 2474 967
rect 2474 915 2486 967
rect 2486 915 2492 967
rect 2516 915 2538 967
rect 2538 915 2550 967
rect 2550 915 2572 967
rect 2596 915 2602 967
rect 2602 915 2614 967
rect 2614 915 2652 967
rect 2676 915 2678 967
rect 2678 915 2730 967
rect 2730 915 2732 967
rect 2756 915 2794 967
rect 2794 915 2806 967
rect 2806 915 2812 967
rect 2836 915 2858 967
rect 2858 915 2870 967
rect 2870 915 2892 967
rect 2916 915 2922 967
rect 2922 915 2934 967
rect 2934 915 2972 967
rect 2996 915 2998 967
rect 2998 915 3050 967
rect 3050 915 3052 967
rect 3076 915 3114 967
rect 3114 915 3126 967
rect 3126 915 3132 967
rect 3156 915 3178 967
rect 3178 915 3190 967
rect 3190 915 3212 967
rect 3236 915 3242 967
rect 3242 915 3254 967
rect 3254 915 3292 967
rect 3316 915 3318 967
rect 3318 915 3370 967
rect 3370 915 3372 967
rect 3396 915 3434 967
rect 3434 915 3446 967
rect 3446 915 3452 967
rect 3476 915 3498 967
rect 3498 915 3510 967
rect 3510 915 3532 967
rect 3556 915 3562 967
rect 3562 915 3574 967
rect 3574 915 3612 967
rect 3636 915 3638 967
rect 3638 915 3690 967
rect 3690 915 3692 967
rect 3716 915 3754 967
rect 3754 915 3766 967
rect 3766 915 3772 967
rect 3796 915 3818 967
rect 3818 915 3830 967
rect 3830 915 3852 967
rect 3876 915 3882 967
rect 3882 915 3894 967
rect 3894 915 3932 967
rect 3956 915 3958 967
rect 3958 915 4010 967
rect 4010 915 4012 967
rect 4036 915 4074 967
rect 4074 915 4086 967
rect 4086 915 4092 967
rect 4116 915 4138 967
rect 4138 915 4150 967
rect 4150 915 4172 967
rect 4196 915 4202 967
rect 4202 915 4214 967
rect 4214 915 4252 967
rect 4276 915 4278 967
rect 4278 915 4330 967
rect 4330 915 4332 967
rect 4356 915 4394 967
rect 4394 915 4406 967
rect 4406 915 4412 967
rect 4436 915 4458 967
rect 4458 915 4470 967
rect 4470 915 4492 967
rect 4516 915 4522 967
rect 4522 915 4534 967
rect 4534 915 4572 967
rect 4596 915 4598 967
rect 4598 915 4650 967
rect 4650 915 4652 967
rect 4676 915 4714 967
rect 4714 915 4726 967
rect 4726 915 4732 967
rect 4756 915 4778 967
rect 4778 915 4790 967
rect 4790 915 4812 967
rect 4836 915 4842 967
rect 4842 915 4854 967
rect 4854 915 4892 967
rect -124 913 -68 915
rect -44 913 12 915
rect 36 913 92 915
rect 116 913 172 915
rect 196 913 252 915
rect 276 913 332 915
rect 356 913 412 915
rect 436 913 492 915
rect 516 913 572 915
rect 596 913 652 915
rect 676 913 732 915
rect 756 913 812 915
rect 836 913 892 915
rect 916 913 972 915
rect 996 913 1052 915
rect 1076 913 1132 915
rect 1156 913 1212 915
rect 1236 913 1292 915
rect 1316 913 1372 915
rect 1396 913 1452 915
rect 1476 913 1532 915
rect 1556 913 1612 915
rect 1636 913 1692 915
rect 1716 913 1772 915
rect 1796 913 1852 915
rect 1876 913 1932 915
rect 1956 913 2012 915
rect 2036 913 2092 915
rect 2116 913 2172 915
rect 2196 913 2252 915
rect 2276 913 2332 915
rect 2356 913 2412 915
rect 2436 913 2492 915
rect 2516 913 2572 915
rect 2596 913 2652 915
rect 2676 913 2732 915
rect 2756 913 2812 915
rect 2836 913 2892 915
rect 2916 913 2972 915
rect 2996 913 3052 915
rect 3076 913 3132 915
rect 3156 913 3212 915
rect 3236 913 3292 915
rect 3316 913 3372 915
rect 3396 913 3452 915
rect 3476 913 3532 915
rect 3556 913 3612 915
rect 3636 913 3692 915
rect 3716 913 3772 915
rect 3796 913 3852 915
rect 3876 913 3932 915
rect 3956 913 4012 915
rect 4036 913 4092 915
rect 4116 913 4172 915
rect 4196 913 4252 915
rect 4276 913 4332 915
rect 4356 913 4412 915
rect 4436 913 4492 915
rect 4516 913 4572 915
rect 4596 913 4652 915
rect 4676 913 4732 915
rect 4756 913 4812 915
rect 4836 913 4892 915
rect 1050 566 1106 622
rect 5114 -298 5170 -242
rect 3624 -362 3680 -358
rect 3624 -414 3630 -362
rect 3630 -414 3680 -362
rect 276 -1428 332 -1426
rect 356 -1428 412 -1426
rect 436 -1428 492 -1426
rect 516 -1428 572 -1426
rect 596 -1428 652 -1426
rect 676 -1428 732 -1426
rect 756 -1428 812 -1426
rect 836 -1428 892 -1426
rect 916 -1428 972 -1426
rect 996 -1428 1052 -1426
rect 1076 -1428 1132 -1426
rect 1156 -1428 1212 -1426
rect 1236 -1428 1292 -1426
rect 1316 -1428 1372 -1426
rect 1396 -1428 1452 -1426
rect 1476 -1428 1532 -1426
rect 1556 -1428 1612 -1426
rect 1636 -1428 1692 -1426
rect 1716 -1428 1772 -1426
rect 1796 -1428 1852 -1426
rect 1876 -1428 1932 -1426
rect 1956 -1428 2012 -1426
rect 2036 -1428 2092 -1426
rect 2116 -1428 2172 -1426
rect 2196 -1428 2252 -1426
rect 2276 -1428 2332 -1426
rect 2356 -1428 2412 -1426
rect 2436 -1428 2492 -1426
rect 2516 -1428 2572 -1426
rect 2596 -1428 2652 -1426
rect 2676 -1428 2732 -1426
rect 2756 -1428 2812 -1426
rect 2836 -1428 2892 -1426
rect 2916 -1428 2972 -1426
rect 2996 -1428 3052 -1426
rect 3076 -1428 3132 -1426
rect 3156 -1428 3212 -1426
rect 3236 -1428 3292 -1426
rect 3316 -1428 3372 -1426
rect 3396 -1428 3452 -1426
rect 3476 -1428 3532 -1426
rect 3556 -1428 3612 -1426
rect 3636 -1428 3692 -1426
rect 3716 -1428 3772 -1426
rect 3796 -1428 3852 -1426
rect 3876 -1428 3932 -1426
rect 276 -1480 286 -1428
rect 286 -1480 332 -1428
rect 356 -1480 402 -1428
rect 402 -1480 412 -1428
rect 436 -1480 466 -1428
rect 466 -1480 478 -1428
rect 478 -1480 492 -1428
rect 516 -1480 530 -1428
rect 530 -1480 542 -1428
rect 542 -1480 572 -1428
rect 596 -1480 606 -1428
rect 606 -1480 652 -1428
rect 676 -1480 722 -1428
rect 722 -1480 732 -1428
rect 756 -1480 786 -1428
rect 786 -1480 798 -1428
rect 798 -1480 812 -1428
rect 836 -1480 850 -1428
rect 850 -1480 862 -1428
rect 862 -1480 892 -1428
rect 916 -1480 926 -1428
rect 926 -1480 972 -1428
rect 996 -1480 1042 -1428
rect 1042 -1480 1052 -1428
rect 1076 -1480 1106 -1428
rect 1106 -1480 1118 -1428
rect 1118 -1480 1132 -1428
rect 1156 -1480 1170 -1428
rect 1170 -1480 1182 -1428
rect 1182 -1480 1212 -1428
rect 1236 -1480 1246 -1428
rect 1246 -1480 1292 -1428
rect 1316 -1480 1362 -1428
rect 1362 -1480 1372 -1428
rect 1396 -1480 1426 -1428
rect 1426 -1480 1438 -1428
rect 1438 -1480 1452 -1428
rect 1476 -1480 1490 -1428
rect 1490 -1480 1502 -1428
rect 1502 -1480 1532 -1428
rect 1556 -1480 1566 -1428
rect 1566 -1480 1612 -1428
rect 1636 -1480 1682 -1428
rect 1682 -1480 1692 -1428
rect 1716 -1480 1746 -1428
rect 1746 -1480 1758 -1428
rect 1758 -1480 1772 -1428
rect 1796 -1480 1810 -1428
rect 1810 -1480 1822 -1428
rect 1822 -1480 1852 -1428
rect 1876 -1480 1886 -1428
rect 1886 -1480 1932 -1428
rect 1956 -1480 2002 -1428
rect 2002 -1480 2012 -1428
rect 2036 -1480 2066 -1428
rect 2066 -1480 2078 -1428
rect 2078 -1480 2092 -1428
rect 2116 -1480 2130 -1428
rect 2130 -1480 2142 -1428
rect 2142 -1480 2172 -1428
rect 2196 -1480 2206 -1428
rect 2206 -1480 2252 -1428
rect 2276 -1480 2322 -1428
rect 2322 -1480 2332 -1428
rect 2356 -1480 2386 -1428
rect 2386 -1480 2398 -1428
rect 2398 -1480 2412 -1428
rect 2436 -1480 2450 -1428
rect 2450 -1480 2462 -1428
rect 2462 -1480 2492 -1428
rect 2516 -1480 2526 -1428
rect 2526 -1480 2572 -1428
rect 2596 -1480 2642 -1428
rect 2642 -1480 2652 -1428
rect 2676 -1480 2706 -1428
rect 2706 -1480 2718 -1428
rect 2718 -1480 2732 -1428
rect 2756 -1480 2770 -1428
rect 2770 -1480 2782 -1428
rect 2782 -1480 2812 -1428
rect 2836 -1480 2846 -1428
rect 2846 -1480 2892 -1428
rect 2916 -1480 2962 -1428
rect 2962 -1480 2972 -1428
rect 2996 -1480 3026 -1428
rect 3026 -1480 3038 -1428
rect 3038 -1480 3052 -1428
rect 3076 -1480 3090 -1428
rect 3090 -1480 3102 -1428
rect 3102 -1480 3132 -1428
rect 3156 -1480 3166 -1428
rect 3166 -1480 3212 -1428
rect 3236 -1480 3282 -1428
rect 3282 -1480 3292 -1428
rect 3316 -1480 3346 -1428
rect 3346 -1480 3358 -1428
rect 3358 -1480 3372 -1428
rect 3396 -1480 3410 -1428
rect 3410 -1480 3422 -1428
rect 3422 -1480 3452 -1428
rect 3476 -1480 3486 -1428
rect 3486 -1480 3532 -1428
rect 3556 -1480 3602 -1428
rect 3602 -1480 3612 -1428
rect 3636 -1480 3666 -1428
rect 3666 -1480 3678 -1428
rect 3678 -1480 3692 -1428
rect 3716 -1480 3730 -1428
rect 3730 -1480 3742 -1428
rect 3742 -1480 3772 -1428
rect 3796 -1480 3806 -1428
rect 3806 -1480 3852 -1428
rect 3876 -1480 3922 -1428
rect 3922 -1480 3932 -1428
rect 276 -1482 332 -1480
rect 356 -1482 412 -1480
rect 436 -1482 492 -1480
rect 516 -1482 572 -1480
rect 596 -1482 652 -1480
rect 676 -1482 732 -1480
rect 756 -1482 812 -1480
rect 836 -1482 892 -1480
rect 916 -1482 972 -1480
rect 996 -1482 1052 -1480
rect 1076 -1482 1132 -1480
rect 1156 -1482 1212 -1480
rect 1236 -1482 1292 -1480
rect 1316 -1482 1372 -1480
rect 1396 -1482 1452 -1480
rect 1476 -1482 1532 -1480
rect 1556 -1482 1612 -1480
rect 1636 -1482 1692 -1480
rect 1716 -1482 1772 -1480
rect 1796 -1482 1852 -1480
rect 1876 -1482 1932 -1480
rect 1956 -1482 2012 -1480
rect 2036 -1482 2092 -1480
rect 2116 -1482 2172 -1480
rect 2196 -1482 2252 -1480
rect 2276 -1482 2332 -1480
rect 2356 -1482 2412 -1480
rect 2436 -1482 2492 -1480
rect 2516 -1482 2572 -1480
rect 2596 -1482 2652 -1480
rect 2676 -1482 2732 -1480
rect 2756 -1482 2812 -1480
rect 2836 -1482 2892 -1480
rect 2916 -1482 2972 -1480
rect 2996 -1482 3052 -1480
rect 3076 -1482 3132 -1480
rect 3156 -1482 3212 -1480
rect 3236 -1482 3292 -1480
rect 3316 -1482 3372 -1480
rect 3396 -1482 3452 -1480
rect 3476 -1482 3532 -1480
rect 3556 -1482 3612 -1480
rect 3636 -1482 3692 -1480
rect 3716 -1482 3772 -1480
rect 3796 -1482 3852 -1480
rect 3876 -1482 3932 -1480
rect -64 -1664 472 -1638
rect -64 -1908 472 -1664
rect -64 -1934 472 -1908
rect 3728 -1664 4264 -1638
rect 3728 -1908 4264 -1664
rect 3728 -1934 4264 -1908
<< metal3 >>
rect 1944 13222 5056 13468
rect 1872 12944 5056 13222
rect -1766 12782 5056 12944
rect -1766 12340 4725 12782
rect -1766 11834 -1052 12340
rect 3922 12198 4725 12340
rect 1870 12068 1970 12090
rect -841 12038 -743 12043
rect 1627 12038 1725 12043
rect -844 12020 1726 12038
rect -844 11956 -824 12020
rect -760 11956 1644 12020
rect 1708 11956 1726 12020
rect -844 11938 1726 11956
rect 1870 12012 1892 12068
rect 1948 12012 1970 12068
rect -841 11933 -743 11938
rect 1627 11933 1725 11938
rect 1870 11834 1970 12012
rect -1766 11818 -734 11834
rect -1766 9672 -736 11818
rect 1890 11744 1970 11834
rect 522 9691 634 9912
rect 517 9672 639 9691
rect -1766 9668 639 9672
rect -1766 9634 546 9668
rect -1766 4336 -1052 9634
rect 517 9604 546 9634
rect 610 9604 639 9668
rect 756 9634 1166 9672
rect 1574 9663 1676 9812
rect 517 9581 639 9604
rect 1574 9607 1597 9663
rect 1653 9607 1676 9663
rect 1574 9584 1676 9607
rect 522 9580 634 9581
rect 914 9364 1026 9392
rect 2088 9387 2200 9388
rect 914 9334 942 9364
rect -804 9308 942 9334
rect 998 9336 1026 9364
rect 2083 9364 2205 9387
rect 998 9334 1298 9336
rect 2083 9334 2112 9364
rect 998 9308 1396 9334
rect -804 4876 1396 9308
rect 1992 9300 2112 9334
rect 2176 9334 2205 9364
rect 3928 9334 4725 12198
rect 2176 9300 4725 9334
rect 1992 7200 4725 9300
rect 1734 6802 4725 7200
rect 1992 5096 4725 6802
rect -804 4844 1224 4876
rect 1286 4844 1396 4876
rect 1286 4662 1390 4844
rect 2112 4665 2204 4880
rect 1286 4606 1310 4662
rect 1366 4606 1390 4662
rect 1286 4582 1390 4606
rect 2107 4652 2209 4665
rect 2107 4588 2126 4652
rect 2190 4588 2209 4652
rect 2358 4643 4725 5096
rect 2107 4575 2209 4588
rect 2112 4574 2204 4575
rect 3922 4404 4725 4643
rect 834 4366 938 4380
rect -1766 2134 -478 4336
rect 834 4302 854 4366
rect 918 4302 938 4366
rect 834 4288 938 4302
rect 1637 4342 1751 4371
rect 840 4180 932 4288
rect 1637 4286 1666 4342
rect 1722 4286 1751 4342
rect 1637 4257 1751 4286
rect 1642 4150 1746 4257
rect -1766 1726 -1052 2134
rect 1291 2030 1389 2035
rect 1290 2029 1796 2030
rect 1290 2012 1801 2029
rect 1290 1948 1308 2012
rect 1372 1948 1714 2012
rect 1778 1948 1801 2012
rect 1290 1931 1801 1948
rect 1290 1930 1796 1931
rect 1291 1925 1389 1930
rect 3928 1810 4725 4404
rect 3922 1726 4725 1810
rect -1766 1206 4725 1726
rect 4941 1206 5056 12782
rect 5243 12762 5353 12789
rect 5243 12761 5270 12762
rect 5326 12761 5353 12762
rect 5243 12697 5266 12761
rect 5330 12697 5353 12761
rect 5243 12673 5353 12697
rect -1766 1126 5056 1206
rect -242 1124 5056 1126
rect -242 969 5054 1124
rect -242 913 -124 969
rect -68 913 -44 969
rect 12 913 36 969
rect 92 913 116 969
rect 172 913 196 969
rect 252 913 276 969
rect 332 913 356 969
rect 412 913 436 969
rect 492 913 516 969
rect 572 913 596 969
rect 652 913 676 969
rect 732 913 756 969
rect 812 913 836 969
rect 892 913 916 969
rect 972 913 996 969
rect 1052 913 1076 969
rect 1132 913 1156 969
rect 1212 913 1236 969
rect 1292 913 1316 969
rect 1372 913 1396 969
rect 1452 913 1476 969
rect 1532 913 1556 969
rect 1612 913 1636 969
rect 1692 913 1716 969
rect 1772 913 1796 969
rect 1852 913 1876 969
rect 1932 913 1956 969
rect 2012 913 2036 969
rect 2092 913 2116 969
rect 2172 913 2196 969
rect 2252 913 2276 969
rect 2332 913 2356 969
rect 2412 913 2436 969
rect 2492 913 2516 969
rect 2572 913 2596 969
rect 2652 913 2676 969
rect 2732 913 2756 969
rect 2812 913 2836 969
rect 2892 913 2916 969
rect 2972 913 2996 969
rect 3052 913 3076 969
rect 3132 913 3156 969
rect 3212 913 3236 969
rect 3292 913 3316 969
rect 3372 913 3396 969
rect 3452 913 3476 969
rect 3532 913 3556 969
rect 3612 913 3636 969
rect 3692 913 3716 969
rect 3772 913 3796 969
rect 3852 913 3876 969
rect 3932 913 3956 969
rect 4012 913 4036 969
rect 4092 913 4116 969
rect 4172 913 4196 969
rect 4252 913 4276 969
rect 4332 913 4356 969
rect 4412 913 4436 969
rect 4492 913 4516 969
rect 4572 913 4596 969
rect 4652 913 4676 969
rect 4732 913 4756 969
rect 4812 913 4836 969
rect 4892 913 5054 969
rect -242 818 5054 913
rect 1291 644 1389 649
rect 1028 626 1390 644
rect 1028 622 1308 626
rect 1028 566 1050 622
rect 1106 566 1308 622
rect 1028 562 1308 566
rect 1372 562 1390 626
rect 1028 544 1390 562
rect 1291 539 1389 544
rect 5247 -220 5345 -215
rect 5094 -238 5346 -220
rect 5094 -242 5264 -238
rect 5094 -298 5114 -242
rect 5170 -298 5264 -242
rect 5094 -302 5264 -298
rect 5328 -302 5346 -238
rect 5094 -320 5346 -302
rect 5247 -325 5345 -320
rect 4043 -336 4141 -331
rect 3602 -354 4142 -336
rect 3602 -358 4060 -354
rect 3602 -414 3624 -358
rect 3680 -414 4060 -358
rect 3602 -418 4060 -414
rect 4124 -418 4142 -354
rect 3602 -436 4142 -418
rect 4043 -441 4141 -436
rect 204 -1422 3996 -1352
rect 204 -1486 272 -1422
rect 336 -1486 352 -1422
rect 416 -1486 432 -1422
rect 496 -1486 512 -1422
rect 576 -1486 592 -1422
rect 656 -1486 672 -1422
rect 736 -1486 752 -1422
rect 816 -1486 832 -1422
rect 896 -1486 912 -1422
rect 976 -1486 992 -1422
rect 1056 -1486 1072 -1422
rect 1136 -1486 1152 -1422
rect 1216 -1486 1232 -1422
rect 1296 -1486 1312 -1422
rect 1376 -1486 1392 -1422
rect 1456 -1486 1472 -1422
rect 1536 -1486 1552 -1422
rect 1616 -1486 1632 -1422
rect 1696 -1486 1712 -1422
rect 1776 -1486 1792 -1422
rect 1856 -1486 1872 -1422
rect 1936 -1486 1952 -1422
rect 2016 -1486 2032 -1422
rect 2096 -1486 2112 -1422
rect 2176 -1486 2192 -1422
rect 2256 -1486 2272 -1422
rect 2336 -1486 2352 -1422
rect 2416 -1486 2432 -1422
rect 2496 -1486 2512 -1422
rect 2576 -1486 2592 -1422
rect 2656 -1486 2672 -1422
rect 2736 -1486 2752 -1422
rect 2816 -1486 2832 -1422
rect 2896 -1486 2912 -1422
rect 2976 -1486 2992 -1422
rect 3056 -1486 3072 -1422
rect 3136 -1486 3152 -1422
rect 3216 -1486 3232 -1422
rect 3296 -1486 3312 -1422
rect 3376 -1486 3392 -1422
rect 3456 -1486 3472 -1422
rect 3536 -1486 3552 -1422
rect 3616 -1486 3632 -1422
rect 3696 -1486 3712 -1422
rect 3776 -1486 3792 -1422
rect 3856 -1486 3872 -1422
rect 3936 -1486 3996 -1422
rect 204 -1550 3996 -1486
rect -106 -1638 514 -1631
rect -106 -1674 -64 -1638
rect 472 -1674 514 -1638
rect -106 -1898 -68 -1674
rect 476 -1898 514 -1674
rect -106 -1934 -64 -1898
rect 472 -1934 514 -1898
rect -106 -1941 514 -1934
rect 3686 -1638 4306 -1631
rect 3686 -1674 3728 -1638
rect 4264 -1674 4306 -1638
rect 3686 -1898 3724 -1674
rect 4268 -1898 4306 -1674
rect 3686 -1934 3728 -1898
rect 4264 -1934 4306 -1898
rect 3686 -1941 4306 -1934
<< via3 >>
rect -824 11956 -760 12020
rect 1644 11956 1708 12020
rect 546 9604 610 9668
rect 2112 9300 2176 9364
rect 2126 4588 2190 4652
rect 854 4302 918 4366
rect 1308 1948 1372 2012
rect 1714 1948 1778 2012
rect 5266 12706 5270 12761
rect 5270 12706 5326 12761
rect 5326 12706 5330 12761
rect 5266 12697 5330 12706
rect 1308 562 1372 626
rect 5264 -302 5328 -238
rect 4060 -418 4124 -354
rect 272 -1426 336 -1422
rect 272 -1482 276 -1426
rect 276 -1482 332 -1426
rect 332 -1482 336 -1426
rect 272 -1486 336 -1482
rect 352 -1426 416 -1422
rect 352 -1482 356 -1426
rect 356 -1482 412 -1426
rect 412 -1482 416 -1426
rect 352 -1486 416 -1482
rect 432 -1426 496 -1422
rect 432 -1482 436 -1426
rect 436 -1482 492 -1426
rect 492 -1482 496 -1426
rect 432 -1486 496 -1482
rect 512 -1426 576 -1422
rect 512 -1482 516 -1426
rect 516 -1482 572 -1426
rect 572 -1482 576 -1426
rect 512 -1486 576 -1482
rect 592 -1426 656 -1422
rect 592 -1482 596 -1426
rect 596 -1482 652 -1426
rect 652 -1482 656 -1426
rect 592 -1486 656 -1482
rect 672 -1426 736 -1422
rect 672 -1482 676 -1426
rect 676 -1482 732 -1426
rect 732 -1482 736 -1426
rect 672 -1486 736 -1482
rect 752 -1426 816 -1422
rect 752 -1482 756 -1426
rect 756 -1482 812 -1426
rect 812 -1482 816 -1426
rect 752 -1486 816 -1482
rect 832 -1426 896 -1422
rect 832 -1482 836 -1426
rect 836 -1482 892 -1426
rect 892 -1482 896 -1426
rect 832 -1486 896 -1482
rect 912 -1426 976 -1422
rect 912 -1482 916 -1426
rect 916 -1482 972 -1426
rect 972 -1482 976 -1426
rect 912 -1486 976 -1482
rect 992 -1426 1056 -1422
rect 992 -1482 996 -1426
rect 996 -1482 1052 -1426
rect 1052 -1482 1056 -1426
rect 992 -1486 1056 -1482
rect 1072 -1426 1136 -1422
rect 1072 -1482 1076 -1426
rect 1076 -1482 1132 -1426
rect 1132 -1482 1136 -1426
rect 1072 -1486 1136 -1482
rect 1152 -1426 1216 -1422
rect 1152 -1482 1156 -1426
rect 1156 -1482 1212 -1426
rect 1212 -1482 1216 -1426
rect 1152 -1486 1216 -1482
rect 1232 -1426 1296 -1422
rect 1232 -1482 1236 -1426
rect 1236 -1482 1292 -1426
rect 1292 -1482 1296 -1426
rect 1232 -1486 1296 -1482
rect 1312 -1426 1376 -1422
rect 1312 -1482 1316 -1426
rect 1316 -1482 1372 -1426
rect 1372 -1482 1376 -1426
rect 1312 -1486 1376 -1482
rect 1392 -1426 1456 -1422
rect 1392 -1482 1396 -1426
rect 1396 -1482 1452 -1426
rect 1452 -1482 1456 -1426
rect 1392 -1486 1456 -1482
rect 1472 -1426 1536 -1422
rect 1472 -1482 1476 -1426
rect 1476 -1482 1532 -1426
rect 1532 -1482 1536 -1426
rect 1472 -1486 1536 -1482
rect 1552 -1426 1616 -1422
rect 1552 -1482 1556 -1426
rect 1556 -1482 1612 -1426
rect 1612 -1482 1616 -1426
rect 1552 -1486 1616 -1482
rect 1632 -1426 1696 -1422
rect 1632 -1482 1636 -1426
rect 1636 -1482 1692 -1426
rect 1692 -1482 1696 -1426
rect 1632 -1486 1696 -1482
rect 1712 -1426 1776 -1422
rect 1712 -1482 1716 -1426
rect 1716 -1482 1772 -1426
rect 1772 -1482 1776 -1426
rect 1712 -1486 1776 -1482
rect 1792 -1426 1856 -1422
rect 1792 -1482 1796 -1426
rect 1796 -1482 1852 -1426
rect 1852 -1482 1856 -1426
rect 1792 -1486 1856 -1482
rect 1872 -1426 1936 -1422
rect 1872 -1482 1876 -1426
rect 1876 -1482 1932 -1426
rect 1932 -1482 1936 -1426
rect 1872 -1486 1936 -1482
rect 1952 -1426 2016 -1422
rect 1952 -1482 1956 -1426
rect 1956 -1482 2012 -1426
rect 2012 -1482 2016 -1426
rect 1952 -1486 2016 -1482
rect 2032 -1426 2096 -1422
rect 2032 -1482 2036 -1426
rect 2036 -1482 2092 -1426
rect 2092 -1482 2096 -1426
rect 2032 -1486 2096 -1482
rect 2112 -1426 2176 -1422
rect 2112 -1482 2116 -1426
rect 2116 -1482 2172 -1426
rect 2172 -1482 2176 -1426
rect 2112 -1486 2176 -1482
rect 2192 -1426 2256 -1422
rect 2192 -1482 2196 -1426
rect 2196 -1482 2252 -1426
rect 2252 -1482 2256 -1426
rect 2192 -1486 2256 -1482
rect 2272 -1426 2336 -1422
rect 2272 -1482 2276 -1426
rect 2276 -1482 2332 -1426
rect 2332 -1482 2336 -1426
rect 2272 -1486 2336 -1482
rect 2352 -1426 2416 -1422
rect 2352 -1482 2356 -1426
rect 2356 -1482 2412 -1426
rect 2412 -1482 2416 -1426
rect 2352 -1486 2416 -1482
rect 2432 -1426 2496 -1422
rect 2432 -1482 2436 -1426
rect 2436 -1482 2492 -1426
rect 2492 -1482 2496 -1426
rect 2432 -1486 2496 -1482
rect 2512 -1426 2576 -1422
rect 2512 -1482 2516 -1426
rect 2516 -1482 2572 -1426
rect 2572 -1482 2576 -1426
rect 2512 -1486 2576 -1482
rect 2592 -1426 2656 -1422
rect 2592 -1482 2596 -1426
rect 2596 -1482 2652 -1426
rect 2652 -1482 2656 -1426
rect 2592 -1486 2656 -1482
rect 2672 -1426 2736 -1422
rect 2672 -1482 2676 -1426
rect 2676 -1482 2732 -1426
rect 2732 -1482 2736 -1426
rect 2672 -1486 2736 -1482
rect 2752 -1426 2816 -1422
rect 2752 -1482 2756 -1426
rect 2756 -1482 2812 -1426
rect 2812 -1482 2816 -1426
rect 2752 -1486 2816 -1482
rect 2832 -1426 2896 -1422
rect 2832 -1482 2836 -1426
rect 2836 -1482 2892 -1426
rect 2892 -1482 2896 -1426
rect 2832 -1486 2896 -1482
rect 2912 -1426 2976 -1422
rect 2912 -1482 2916 -1426
rect 2916 -1482 2972 -1426
rect 2972 -1482 2976 -1426
rect 2912 -1486 2976 -1482
rect 2992 -1426 3056 -1422
rect 2992 -1482 2996 -1426
rect 2996 -1482 3052 -1426
rect 3052 -1482 3056 -1426
rect 2992 -1486 3056 -1482
rect 3072 -1426 3136 -1422
rect 3072 -1482 3076 -1426
rect 3076 -1482 3132 -1426
rect 3132 -1482 3136 -1426
rect 3072 -1486 3136 -1482
rect 3152 -1426 3216 -1422
rect 3152 -1482 3156 -1426
rect 3156 -1482 3212 -1426
rect 3212 -1482 3216 -1426
rect 3152 -1486 3216 -1482
rect 3232 -1426 3296 -1422
rect 3232 -1482 3236 -1426
rect 3236 -1482 3292 -1426
rect 3292 -1482 3296 -1426
rect 3232 -1486 3296 -1482
rect 3312 -1426 3376 -1422
rect 3312 -1482 3316 -1426
rect 3316 -1482 3372 -1426
rect 3372 -1482 3376 -1426
rect 3312 -1486 3376 -1482
rect 3392 -1426 3456 -1422
rect 3392 -1482 3396 -1426
rect 3396 -1482 3452 -1426
rect 3452 -1482 3456 -1426
rect 3392 -1486 3456 -1482
rect 3472 -1426 3536 -1422
rect 3472 -1482 3476 -1426
rect 3476 -1482 3532 -1426
rect 3532 -1482 3536 -1426
rect 3472 -1486 3536 -1482
rect 3552 -1426 3616 -1422
rect 3552 -1482 3556 -1426
rect 3556 -1482 3612 -1426
rect 3612 -1482 3616 -1426
rect 3552 -1486 3616 -1482
rect 3632 -1426 3696 -1422
rect 3632 -1482 3636 -1426
rect 3636 -1482 3692 -1426
rect 3692 -1482 3696 -1426
rect 3632 -1486 3696 -1482
rect 3712 -1426 3776 -1422
rect 3712 -1482 3716 -1426
rect 3716 -1482 3772 -1426
rect 3772 -1482 3776 -1426
rect 3712 -1486 3776 -1482
rect 3792 -1426 3856 -1422
rect 3792 -1482 3796 -1426
rect 3796 -1482 3852 -1426
rect 3852 -1482 3856 -1426
rect 3792 -1486 3856 -1482
rect 3872 -1426 3936 -1422
rect 3872 -1482 3876 -1426
rect 3876 -1482 3932 -1426
rect 3932 -1482 3936 -1426
rect 3872 -1486 3936 -1482
rect -68 -1898 -64 -1674
rect -64 -1898 472 -1674
rect 472 -1898 476 -1674
rect 3724 -1898 3728 -1674
rect 3728 -1898 4264 -1674
rect 4264 -1898 4268 -1674
<< metal4 >>
rect 1944 28680 2742 29480
rect 17174 13068 17274 13680
rect 15670 12968 17274 13068
rect 15670 12784 15770 12968
rect 5246 12780 15770 12784
rect 5242 12761 15770 12780
rect -1744 12706 -1644 12734
rect -1750 12606 1212 12706
rect 1654 12606 4620 12706
rect 5242 12697 5266 12761
rect 5330 12697 15770 12761
rect 5242 12684 15770 12697
rect 5242 12678 5354 12684
rect -1744 10950 -1644 12606
rect 1238 12182 3888 12282
rect -1110 12020 -742 12038
rect -1110 11956 -824 12020
rect -760 11956 -742 12020
rect -1110 11938 -742 11956
rect -1744 10850 -1318 10950
rect -1744 8336 -1644 10850
rect -1110 9134 -1010 11938
rect 1238 11660 1338 12182
rect 884 11560 1338 11660
rect 1626 12020 1726 12038
rect 1626 11956 1644 12020
rect 1708 11956 1726 12020
rect 1626 11086 1726 11956
rect 522 9668 2200 9692
rect 522 9604 546 9668
rect 610 9604 2200 9668
rect 522 9580 2200 9604
rect 2088 9364 2200 9580
rect 2088 9300 2112 9364
rect 2176 9300 2200 9364
rect 2088 9276 2200 9300
rect 3788 9134 3888 12182
rect 4520 10936 4620 12606
rect 4162 10828 4620 10936
rect -1110 9034 -434 9134
rect 3246 9034 3888 9134
rect 4520 8336 4620 10828
rect -1752 8228 -1294 8336
rect 4162 8228 4620 8336
rect -1744 5836 -1644 8228
rect 246 6546 346 7417
rect 2522 6546 2622 7417
rect -1752 5728 -1294 5836
rect 4520 5736 4620 8228
rect -1744 3236 -1644 5728
rect 4162 5628 4620 5736
rect -1108 4782 -358 4882
rect 3020 4786 3891 4886
rect -1752 3128 -1264 3236
rect -1744 1478 -1644 3128
rect -1108 2030 -1008 4782
rect 2112 4652 2204 4666
rect 2112 4588 2126 4652
rect 2190 4588 2204 4652
rect 839 4380 933 4381
rect 2112 4380 2204 4588
rect 839 4366 2204 4380
rect 839 4302 854 4366
rect 918 4302 2204 4366
rect 839 4288 2204 4302
rect 839 4287 933 4288
rect 890 2196 1018 2414
rect 890 2096 1590 2196
rect -1108 2012 1390 2030
rect -1108 1948 1308 2012
rect 1372 1948 1390 2012
rect -1108 1930 1390 1948
rect -1744 1378 1206 1478
rect 1290 626 1390 1930
rect 1490 1840 1590 2096
rect 1696 2012 1796 2654
rect 1696 1948 1714 2012
rect 1778 1948 1796 2012
rect 1696 1930 1796 1948
rect 3791 1840 3891 4786
rect 4520 3236 4620 5628
rect 4162 3128 4620 3236
rect 1490 1740 3891 1840
rect 1490 1140 1590 1740
rect 4520 1478 4620 3128
rect 1658 1378 4620 1478
rect 1490 1040 4142 1140
rect 1290 562 1308 626
rect 1372 562 1390 626
rect 1290 544 1390 562
rect 4042 -354 4142 1040
rect 5246 -238 5346 12678
rect 5246 -302 5264 -238
rect 5328 -302 5346 -238
rect 5246 -320 5346 -302
rect 4042 -418 4060 -354
rect 4124 -418 4142 -354
rect 4042 -436 4142 -418
rect -280 -1422 4480 -1320
rect -280 -1486 272 -1422
rect 336 -1486 352 -1422
rect 416 -1486 432 -1422
rect 496 -1486 512 -1422
rect 576 -1486 592 -1422
rect 656 -1486 672 -1422
rect 736 -1486 752 -1422
rect 816 -1486 832 -1422
rect 896 -1486 912 -1422
rect 976 -1486 992 -1422
rect 1056 -1486 1072 -1422
rect 1136 -1486 1152 -1422
rect 1216 -1486 1232 -1422
rect 1296 -1486 1312 -1422
rect 1376 -1486 1392 -1422
rect 1456 -1486 1472 -1422
rect 1536 -1486 1552 -1422
rect 1616 -1486 1632 -1422
rect 1696 -1486 1712 -1422
rect 1776 -1486 1792 -1422
rect 1856 -1486 1872 -1422
rect 1936 -1486 1952 -1422
rect 2016 -1486 2032 -1422
rect 2096 -1486 2112 -1422
rect 2176 -1486 2192 -1422
rect 2256 -1486 2272 -1422
rect 2336 -1486 2352 -1422
rect 2416 -1486 2432 -1422
rect 2496 -1486 2512 -1422
rect 2576 -1486 2592 -1422
rect 2656 -1486 2672 -1422
rect 2736 -1486 2752 -1422
rect 2816 -1486 2832 -1422
rect 2896 -1486 2912 -1422
rect 2976 -1486 2992 -1422
rect 3056 -1486 3072 -1422
rect 3136 -1486 3152 -1422
rect 3216 -1486 3232 -1422
rect 3296 -1486 3312 -1422
rect 3376 -1486 3392 -1422
rect 3456 -1486 3472 -1422
rect 3536 -1486 3552 -1422
rect 3616 -1486 3632 -1422
rect 3696 -1486 3712 -1422
rect 3776 -1486 3792 -1422
rect 3856 -1486 3872 -1422
rect 3936 -1486 4480 -1422
rect -280 -1674 4480 -1486
rect -280 -1898 -68 -1674
rect 476 -1898 3724 -1674
rect 4268 -1898 4480 -1674
rect -280 -2120 4480 -1898
use sky130_fd_pr__cap_mim_m3_1_KBZ9JD  sky130_fd_pr__cap_mim_m3_1_KBZ9JD_7
timestamp 1626486988
transform 1 0 106 0 1 3234
box -1150 -1100 1050 1100
use sky130_fd_pr__cap_mim_m3_1_KBZ9JD  sky130_fd_pr__cap_mim_m3_1_KBZ9JD_6
timestamp 1626486988
transform 1 0 2628 0 1 3234
box -1150 -1100 1050 1100
use sky130_fd_pr__nfet_01v8_USKJ3F  sky130_fd_pr__nfet_01v8_USKJ3F_1
timestamp 1626486988
transform 1 0 2109 0 1 242
box -1861 -288 1861 288
use sky130_fd_pr__nfet_01v8_USKJ3F  sky130_fd_pr__nfet_01v8_USKJ3F_0
timestamp 1626486988
transform 1 0 2109 0 1 -758
box -1861 -288 1861 288
use sky130_fd_pr__cap_mim_m3_1_XQCLDR  sky130_fd_pr__cap_mim_m3_1_XQCLDR_3
timestamp 1626486988
transform -1 0 -1407 0 -1 3106
box -350 -1300 349 1300
use sky130_fd_pr__cap_mim_m3_1_5E2G4H  sky130_fd_pr__cap_mim_m3_1_5E2G4H_3
timestamp 1626486988
transform 1 0 3068 0 -1 1426
box -1550 -300 1549 300
use sky130_fd_pr__cap_mim_m3_1_5E2G4H  sky130_fd_pr__cap_mim_m3_1_5E2G4H_2
timestamp 1626486988
transform -1 0 -203 0 -1 1426
box -1550 -300 1549 300
use sky130_fd_pr__cap_mim_m3_1_XQCLDR  sky130_fd_pr__cap_mim_m3_1_XQCLDR_2
timestamp 1626486988
transform 1 0 4272 0 -1 3106
box -350 -1300 349 1300
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_3
timestamp 1626486988
transform -1 0 -1407 0 -1 8250
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_2
timestamp 1626486988
transform -1 0 -1407 0 1 5756
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_KBZ9JD  sky130_fd_pr__cap_mim_m3_1_KBZ9JD_5
timestamp 1626486988
transform 1 0 346 0 1 5734
box -1150 -1100 1050 1100
use sky130_fd_pr__cap_mim_m3_1_KBZ9JD  sky130_fd_pr__cap_mim_m3_1_KBZ9JD_4
timestamp 1626486988
transform 1 0 346 0 1 8234
box -1150 -1100 1050 1100
use sky130_fd_pr__cap_mim_m3_1_KBZ9JD  sky130_fd_pr__cap_mim_m3_1_KBZ9JD_3
timestamp 1626486988
transform 1 0 2884 0 1 8234
box -1150 -1100 1050 1100
use sky130_fd_pr__cap_mim_m3_1_KBZ9JD  sky130_fd_pr__cap_mim_m3_1_KBZ9JD_2
timestamp 1626486988
transform 1 0 2884 0 1 5734
box -1150 -1100 1050 1100
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_1
timestamp 1626486988
transform 1 0 4272 0 1 5756
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_0
timestamp 1626486988
transform 1 0 4272 0 -1 8250
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_KBZ9JD  sky130_fd_pr__cap_mim_m3_1_KBZ9JD_1
timestamp 1626486988
transform 1 0 116 0 1 10734
box -1150 -1100 1050 1100
use sky130_fd_pr__cap_mim_m3_1_KBZ9JD  sky130_fd_pr__cap_mim_m3_1_KBZ9JD_0
timestamp 1626486988
transform 1 0 2626 0 1 10734
box -1150 -1100 1050 1100
use sky130_fd_pr__cap_mim_m3_1_XQCLDR  sky130_fd_pr__cap_mim_m3_1_XQCLDR_1
timestamp 1626486988
transform -1 0 -1407 0 1 10900
box -350 -1300 349 1300
use sky130_fd_pr__cap_mim_m3_1_5E2G4H  sky130_fd_pr__cap_mim_m3_1_5E2G4H_1
timestamp 1626486988
transform 1 0 3068 0 1 12640
box -1550 -300 1549 300
use sky130_fd_pr__cap_mim_m3_1_5E2G4H  sky130_fd_pr__cap_mim_m3_1_5E2G4H_0
timestamp 1626486988
transform -1 0 -203 0 1 12640
box -1550 -300 1549 300
use sky130_fd_pr__cap_mim_m3_1_XQCLDR  sky130_fd_pr__cap_mim_m3_1_XQCLDR_0
timestamp 1626486988
transform 1 0 4272 0 1 10900
box -350 -1300 349 1300
use se_fold_casc_wide_swing_ota  se_fold_casc_wide_swing_ota_0
timestamp 1626486988
transform 1 0 17040 0 1 25080
box -15168 -27248 25000 4400
<< labels >>
flabel metal2 s 2362 -152 2380 -136 1 FreeSans 600 0 0 0 clk
flabel metal2 s 2348 -280 2366 -264 1 FreeSans 600 0 0 0 vout
flabel metal1 s 18 -178 30 -162 1 FreeSans 600 0 0 0 vin
flabel metal2 s 1848 -1132 1870 -1116 1 FreeSans 600 0 0 0 vholdm
flabel metal2 s 2620 -404 2638 -386 1 FreeSans 600 0 0 0 vhold
flabel metal4 s 3836 11340 3852 11354 1 FreeSans 600 0 0 0 vhold
flabel metal1 s 6974 124 6984 136 1 FreeSans 600 0 0 0 ibiasn
flabel metal4 s 2134 29128 2186 29174 1 FreeSans 600 0 0 0 VDD
flabel metal4 s -1076 11268 -1050 11288 1 FreeSans 600 0 0 0 vholdm
flabel metal3 s 1324 6968 1358 6998 1 FreeSans 600 0 0 0 vout
flabel metal4 s -266 -1346 -260 -1342 1 FreeSans 600 0 0 0 VSS
<< properties >>
string FIXED_BBOX -152 -1992 4352 1492
<< end >>
