magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< locali >>
rect 94 3062 1942 3096
rect 3259 3023 3836 3057
rect 174 2950 1832 2984
rect 254 2860 1942 2894
rect 1636 2636 1942 2670
rect 1556 2546 1832 2580
rect 3259 2473 3836 2507
rect 1236 2434 1942 2468
rect 1476 2272 1942 2306
rect 3259 2233 3836 2267
rect 1316 2160 1832 2194
rect 1636 2070 1942 2104
rect 1636 1846 1942 1880
rect 1316 1756 1832 1790
rect 3259 1683 3836 1717
rect 1236 1644 1942 1678
rect 1476 1482 1942 1516
rect 3259 1443 3836 1477
rect 1556 1370 1832 1404
rect 1396 1280 1942 1314
rect 1396 1056 1942 1090
rect 254 943 494 977
rect 1556 966 1832 1000
rect 3259 893 3836 927
rect 1236 854 1942 888
rect 1476 692 1942 726
rect 3259 653 3836 687
rect 174 603 494 637
rect 1316 580 1832 614
rect 1396 490 1942 524
rect 1396 266 1942 300
rect 94 153 494 187
rect 1316 176 1832 210
rect 3259 103 3836 137
rect 1236 64 1942 98
<< metal1 >>
rect 80 199 108 3080
rect 160 649 188 3080
rect 240 989 268 3080
rect 231 931 277 989
rect 151 591 197 649
rect 71 141 117 199
rect 80 80 108 141
rect 160 80 188 591
rect 240 80 268 931
rect 584 80 612 1185
rect 980 80 1008 1185
rect 1110 884 1174 936
rect 1110 644 1174 696
rect 1110 94 1174 146
rect 1222 80 1250 3080
rect 1302 80 1330 3080
rect 1382 80 1410 3080
rect 1462 80 1490 3080
rect 1542 80 1570 3080
rect 1622 80 1650 3080
rect 2030 80 2076 3204
rect 2454 80 2502 3146
rect 2886 80 2934 3146
rect 3278 80 3306 3160
rect 3674 80 3702 3160
<< metal2 >>
rect 2025 2764 2081 2812
rect 2450 2764 2506 2812
rect 2882 2764 2938 2812
rect 3264 2741 3320 2789
rect 3660 2741 3716 2789
rect 2025 1974 2081 2022
rect 2450 1974 2506 2022
rect 2882 1974 2938 2022
rect 3264 1951 3320 1999
rect 3660 1951 3716 1999
rect 2025 1184 2081 1232
rect 2450 1184 2506 1232
rect 2882 1184 2938 1232
rect 3264 1161 3320 1209
rect 3660 1161 3716 1209
rect 1128 1087 1396 1115
rect 1128 910 1156 1087
rect 1128 692 1316 720
rect 1128 670 1156 692
rect 570 371 626 419
rect 966 371 1022 419
rect 2025 394 2081 442
rect 2450 394 2506 442
rect 2882 394 2938 442
rect 3264 371 3320 419
rect 3660 371 3716 419
rect 1128 297 1236 325
rect 1128 120 1156 297
<< metal3 >>
rect 2004 2739 2102 2837
rect 2429 2739 2527 2837
rect 2861 2739 2959 2837
rect 3243 2716 3341 2814
rect 3639 2716 3737 2814
rect 2004 1949 2102 2047
rect 2429 1949 2527 2047
rect 2861 1949 2959 2047
rect 3243 1926 3341 2024
rect 3639 1926 3737 2024
rect 2004 1159 2102 1257
rect 2429 1159 2527 1257
rect 2861 1159 2959 1257
rect 3243 1136 3341 1234
rect 3639 1136 3737 1234
rect 549 346 647 444
rect 945 346 1043 444
rect 2004 369 2102 467
rect 2429 369 2527 467
rect 2861 369 2959 467
rect 3243 346 3341 444
rect 3639 346 3737 444
use contact_16  contact_16_26
timestamp 1624494425
transform 1 0 61 0 1 141
box 0 0 66 58
use contact_8  contact_8_8
timestamp 1624494425
transform 1 0 566 0 1 363
box 0 0 64 64
use contact_9  contact_9_8
timestamp 1624494425
transform 1 0 565 0 1 358
box 0 0 66 74
use pinv_dec  pinv_dec_1
timestamp 1624494425
transform 1 0 400 0 -1 790
box 44 0 760 490
use pinv_dec  pinv_dec_2
timestamp 1624494425
transform 1 0 400 0 1 0
box 44 0 760 490
use contact_7  contact_7_8
timestamp 1624494425
transform 1 0 1113 0 1 87
box 0 0 58 66
use contact_8  contact_8_24
timestamp 1624494425
transform 1 0 1110 0 1 88
box 0 0 64 64
use contact_17  contact_17_2
timestamp 1624494425
transform 1 0 1204 0 1 279
box 0 0 64 64
use contact_16  contact_16_23
timestamp 1624494425
transform 1 0 1203 0 1 52
box 0 0 66 58
use contact_16  contact_16_22
timestamp 1624494425
transform 1 0 1283 0 1 164
box 0 0 66 58
use contact_16  contact_16_21
timestamp 1624494425
transform 1 0 1363 0 1 254
box 0 0 66 58
use contact_16  contact_16_18
timestamp 1624494425
transform 1 0 1363 0 1 478
box 0 0 66 58
use contact_8  contact_8_21
timestamp 1624494425
transform 1 0 962 0 1 363
box 0 0 64 64
use contact_9  contact_9_21
timestamp 1624494425
transform 1 0 961 0 1 358
box 0 0 66 74
use contact_8  contact_8_7
timestamp 1624494425
transform 1 0 2021 0 1 386
box 0 0 64 64
use contact_9  contact_9_7
timestamp 1624494425
transform 1 0 2020 0 1 381
box 0 0 66 74
use contact_8  contact_8_19
timestamp 1624494425
transform 1 0 2446 0 1 386
box 0 0 64 64
use contact_9  contact_9_19
timestamp 1624494425
transform 1 0 2445 0 1 381
box 0 0 66 74
use contact_8  contact_8_20
timestamp 1624494425
transform 1 0 2878 0 1 386
box 0 0 64 64
use contact_9  contact_9_20
timestamp 1624494425
transform 1 0 2877 0 1 381
box 0 0 66 74
use contact_8  contact_8_6
timestamp 1624494425
transform 1 0 3260 0 1 363
box 0 0 64 64
use contact_9  contact_9_6
timestamp 1624494425
transform 1 0 3259 0 1 358
box 0 0 66 74
use contact_8  contact_8_18
timestamp 1624494425
transform 1 0 3656 0 1 363
box 0 0 64 64
use contact_9  contact_9_18
timestamp 1624494425
transform 1 0 3655 0 1 358
box 0 0 66 74
use and3_dec  and3_dec_7
timestamp 1624494425
transform 1 0 1782 0 1 0
box 0 -60 2072 490
use and3_dec  and3_dec_6
timestamp 1624494425
transform 1 0 1782 0 -1 790
box 0 -60 2072 490
use contact_16  contact_16_25
timestamp 1624494425
transform 1 0 141 0 1 591
box 0 0 66 58
use contact_16  contact_16_24
timestamp 1624494425
transform 1 0 221 0 1 931
box 0 0 66 58
use pinv_dec  pinv_dec_0
timestamp 1624494425
transform 1 0 400 0 1 790
box 44 0 760 490
use contact_7  contact_7_7
timestamp 1624494425
transform 1 0 1113 0 1 637
box 0 0 58 66
use contact_8  contact_8_23
timestamp 1624494425
transform 1 0 1110 0 1 638
box 0 0 64 64
use contact_17  contact_17_1
timestamp 1624494425
transform 1 0 1284 0 1 674
box 0 0 64 64
use contact_7  contact_7_6
timestamp 1624494425
transform 1 0 1113 0 1 877
box 0 0 58 66
use contact_8  contact_8_22
timestamp 1624494425
transform 1 0 1110 0 1 878
box 0 0 64 64
use contact_16  contact_16_20
timestamp 1624494425
transform 1 0 1443 0 1 680
box 0 0 66 58
use contact_16  contact_16_19
timestamp 1624494425
transform 1 0 1283 0 1 568
box 0 0 66 58
use contact_16  contact_16_17
timestamp 1624494425
transform 1 0 1203 0 1 842
box 0 0 66 58
use contact_16  contact_16_16
timestamp 1624494425
transform 1 0 1523 0 1 954
box 0 0 66 58
use and3_dec  and3_dec_5
timestamp 1624494425
transform 1 0 1782 0 1 790
box 0 -60 2072 490
use contact_17  contact_17_0
timestamp 1624494425
transform 1 0 1364 0 1 1069
box 0 0 64 64
use contact_16  contact_16_15
timestamp 1624494425
transform 1 0 1363 0 1 1044
box 0 0 66 58
use contact_16  contact_16_12
timestamp 1624494425
transform 1 0 1363 0 1 1268
box 0 0 66 58
use contact_8  contact_8_5
timestamp 1624494425
transform 1 0 2021 0 1 1176
box 0 0 64 64
use contact_9  contact_9_5
timestamp 1624494425
transform 1 0 2020 0 1 1171
box 0 0 66 74
use contact_8  contact_8_16
timestamp 1624494425
transform 1 0 2446 0 1 1176
box 0 0 64 64
use contact_9  contact_9_16
timestamp 1624494425
transform 1 0 2445 0 1 1171
box 0 0 66 74
use contact_8  contact_8_17
timestamp 1624494425
transform 1 0 2878 0 1 1176
box 0 0 64 64
use contact_9  contact_9_17
timestamp 1624494425
transform 1 0 2877 0 1 1171
box 0 0 66 74
use contact_8  contact_8_4
timestamp 1624494425
transform 1 0 3260 0 1 1153
box 0 0 64 64
use contact_9  contact_9_4
timestamp 1624494425
transform 1 0 3259 0 1 1148
box 0 0 66 74
use contact_8  contact_8_15
timestamp 1624494425
transform 1 0 3656 0 1 1153
box 0 0 64 64
use contact_9  contact_9_15
timestamp 1624494425
transform 1 0 3655 0 1 1148
box 0 0 66 74
use contact_16  contact_16_13
timestamp 1624494425
transform 1 0 1523 0 1 1358
box 0 0 66 58
use contact_16  contact_16_14
timestamp 1624494425
transform 1 0 1443 0 1 1470
box 0 0 66 58
use and3_dec  and3_dec_4
timestamp 1624494425
transform 1 0 1782 0 -1 1580
box 0 -60 2072 490
use and3_dec  and3_dec_3
timestamp 1624494425
transform 1 0 1782 0 1 1580
box 0 -60 2072 490
use contact_16  contact_16_9
timestamp 1624494425
transform 1 0 1603 0 1 1834
box 0 0 66 58
use contact_16  contact_16_10
timestamp 1624494425
transform 1 0 1283 0 1 1744
box 0 0 66 58
use contact_16  contact_16_11
timestamp 1624494425
transform 1 0 1203 0 1 1632
box 0 0 66 58
use contact_16  contact_16_6
timestamp 1624494425
transform 1 0 1603 0 1 2058
box 0 0 66 58
use contact_8  contact_8_3
timestamp 1624494425
transform 1 0 2021 0 1 1966
box 0 0 64 64
use contact_9  contact_9_3
timestamp 1624494425
transform 1 0 2020 0 1 1961
box 0 0 66 74
use contact_8  contact_8_13
timestamp 1624494425
transform 1 0 2446 0 1 1966
box 0 0 64 64
use contact_9  contact_9_13
timestamp 1624494425
transform 1 0 2445 0 1 1961
box 0 0 66 74
use contact_8  contact_8_14
timestamp 1624494425
transform 1 0 2878 0 1 1966
box 0 0 64 64
use contact_9  contact_9_14
timestamp 1624494425
transform 1 0 2877 0 1 1961
box 0 0 66 74
use contact_8  contact_8_2
timestamp 1624494425
transform 1 0 3260 0 1 1943
box 0 0 64 64
use contact_9  contact_9_2
timestamp 1624494425
transform 1 0 3259 0 1 1938
box 0 0 66 74
use contact_8  contact_8_12
timestamp 1624494425
transform 1 0 3656 0 1 1943
box 0 0 64 64
use contact_9  contact_9_12
timestamp 1624494425
transform 1 0 3655 0 1 1938
box 0 0 66 74
use and3_dec  and3_dec_2
timestamp 1624494425
transform 1 0 1782 0 -1 2370
box 0 -60 2072 490
use contact_16  contact_16_8
timestamp 1624494425
transform 1 0 1443 0 1 2260
box 0 0 66 58
use contact_16  contact_16_7
timestamp 1624494425
transform 1 0 1283 0 1 2148
box 0 0 66 58
use contact_16  contact_16_5
timestamp 1624494425
transform 1 0 1203 0 1 2422
box 0 0 66 58
use contact_16  contact_16_4
timestamp 1624494425
transform 1 0 1523 0 1 2534
box 0 0 66 58
use contact_16  contact_16_3
timestamp 1624494425
transform 1 0 1603 0 1 2624
box 0 0 66 58
use and3_dec  and3_dec_0
timestamp 1624494425
transform 1 0 1782 0 -1 3160
box 0 -60 2072 490
use and3_dec  and3_dec_1
timestamp 1624494425
transform 1 0 1782 0 1 2370
box 0 -60 2072 490
use contact_7  contact_7_1
timestamp 1624494425
transform 1 0 225 0 1 2844
box 0 0 58 66
use contact_7  contact_7_3
timestamp 1624494425
transform 1 0 145 0 1 2934
box 0 0 58 66
use contact_7  contact_7_5
timestamp 1624494425
transform 1 0 65 0 1 3046
box 0 0 58 66
use contact_16  contact_16_2
timestamp 1624494425
transform 1 0 1443 0 1 3050
box 0 0 66 58
use contact_7  contact_7_4
timestamp 1624494425
transform 1 0 1447 0 1 3046
box 0 0 58 66
use contact_16  contact_16_0
timestamp 1624494425
transform 1 0 1603 0 1 2848
box 0 0 66 58
use contact_16  contact_16_1
timestamp 1624494425
transform 1 0 1523 0 1 2938
box 0 0 66 58
use contact_7  contact_7_0
timestamp 1624494425
transform 1 0 1607 0 1 2844
box 0 0 58 66
use contact_7  contact_7_2
timestamp 1624494425
transform 1 0 1527 0 1 2934
box 0 0 58 66
use contact_9  contact_9_1
timestamp 1624494425
transform 1 0 2020 0 1 2751
box 0 0 66 74
use contact_8  contact_8_1
timestamp 1624494425
transform 1 0 2021 0 1 2756
box 0 0 64 64
use contact_9  contact_9_10
timestamp 1624494425
transform 1 0 2445 0 1 2751
box 0 0 66 74
use contact_8  contact_8_10
timestamp 1624494425
transform 1 0 2446 0 1 2756
box 0 0 64 64
use contact_9  contact_9_11
timestamp 1624494425
transform 1 0 2877 0 1 2751
box 0 0 66 74
use contact_8  contact_8_11
timestamp 1624494425
transform 1 0 2878 0 1 2756
box 0 0 64 64
use contact_9  contact_9_0
timestamp 1624494425
transform 1 0 3259 0 1 2728
box 0 0 66 74
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 3260 0 1 2733
box 0 0 64 64
use contact_9  contact_9_9
timestamp 1624494425
transform 1 0 3655 0 1 2728
box 0 0 66 74
use contact_8  contact_8_9
timestamp 1624494425
transform 1 0 3656 0 1 2733
box 0 0 64 64
<< labels >>
rlabel metal1 s 71 141 117 199 4 in_0
rlabel metal1 s 151 591 197 649 4 in_1
rlabel metal1 s 231 931 277 989 4 in_2
rlabel locali s 3547 120 3547 120 4 out_0
rlabel locali s 3547 670 3547 670 4 out_1
rlabel locali s 3547 910 3547 910 4 out_2
rlabel locali s 3547 1460 3547 1460 4 out_3
rlabel locali s 3547 1700 3547 1700 4 out_4
rlabel locali s 3547 2250 3547 2250 4 out_5
rlabel locali s 3547 2490 3547 2490 4 out_6
rlabel locali s 3547 3040 3547 3040 4 out_7
rlabel metal3 s 2429 1949 2527 2047 4 vdd
rlabel metal3 s 2861 2739 2959 2837 4 vdd
rlabel metal3 s 2861 1949 2959 2047 4 vdd
rlabel metal3 s 2429 1159 2527 1257 4 vdd
rlabel metal3 s 3639 2716 3737 2814 4 vdd
rlabel metal3 s 3639 346 3737 444 4 vdd
rlabel metal3 s 2429 2739 2527 2837 4 vdd
rlabel metal3 s 3639 1136 3737 1234 4 vdd
rlabel metal3 s 2861 369 2959 467 4 vdd
rlabel metal3 s 2429 369 2527 467 4 vdd
rlabel metal3 s 3639 1926 3737 2024 4 vdd
rlabel metal3 s 945 346 1043 444 4 vdd
rlabel metal3 s 2861 1159 2959 1257 4 vdd
rlabel metal3 s 2004 1949 2102 2047 4 gnd
rlabel metal3 s 2004 1159 2102 1257 4 gnd
rlabel metal3 s 2004 369 2102 467 4 gnd
rlabel metal3 s 3243 346 3341 444 4 gnd
rlabel metal3 s 549 346 647 444 4 gnd
rlabel metal3 s 3243 1926 3341 2024 4 gnd
rlabel metal3 s 3243 1136 3341 1234 4 gnd
rlabel metal3 s 2004 2739 2102 2837 4 gnd
rlabel metal3 s 3243 2716 3341 2814 4 gnd
<< properties >>
string FIXED_BBOX 0 0 3836 3160
<< end >>
