magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -2615 -1460 2615 1460
<< nwell >>
rect -1355 -200 1355 200
<< pmos >>
rect -1261 -100 -1061 100
rect -1003 -100 -803 100
rect -745 -100 -545 100
rect -487 -100 -287 100
rect -229 -100 -29 100
rect 29 -100 229 100
rect 287 -100 487 100
rect 545 -100 745 100
rect 803 -100 1003 100
rect 1061 -100 1261 100
<< pdiff >>
rect -1319 85 -1261 100
rect -1319 51 -1307 85
rect -1273 51 -1261 85
rect -1319 17 -1261 51
rect -1319 -17 -1307 17
rect -1273 -17 -1261 17
rect -1319 -51 -1261 -17
rect -1319 -85 -1307 -51
rect -1273 -85 -1261 -51
rect -1319 -100 -1261 -85
rect -1061 85 -1003 100
rect -1061 51 -1049 85
rect -1015 51 -1003 85
rect -1061 17 -1003 51
rect -1061 -17 -1049 17
rect -1015 -17 -1003 17
rect -1061 -51 -1003 -17
rect -1061 -85 -1049 -51
rect -1015 -85 -1003 -51
rect -1061 -100 -1003 -85
rect -803 85 -745 100
rect -803 51 -791 85
rect -757 51 -745 85
rect -803 17 -745 51
rect -803 -17 -791 17
rect -757 -17 -745 17
rect -803 -51 -745 -17
rect -803 -85 -791 -51
rect -757 -85 -745 -51
rect -803 -100 -745 -85
rect -545 85 -487 100
rect -545 51 -533 85
rect -499 51 -487 85
rect -545 17 -487 51
rect -545 -17 -533 17
rect -499 -17 -487 17
rect -545 -51 -487 -17
rect -545 -85 -533 -51
rect -499 -85 -487 -51
rect -545 -100 -487 -85
rect -287 85 -229 100
rect -287 51 -275 85
rect -241 51 -229 85
rect -287 17 -229 51
rect -287 -17 -275 17
rect -241 -17 -229 17
rect -287 -51 -229 -17
rect -287 -85 -275 -51
rect -241 -85 -229 -51
rect -287 -100 -229 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 229 85 287 100
rect 229 51 241 85
rect 275 51 287 85
rect 229 17 287 51
rect 229 -17 241 17
rect 275 -17 287 17
rect 229 -51 287 -17
rect 229 -85 241 -51
rect 275 -85 287 -51
rect 229 -100 287 -85
rect 487 85 545 100
rect 487 51 499 85
rect 533 51 545 85
rect 487 17 545 51
rect 487 -17 499 17
rect 533 -17 545 17
rect 487 -51 545 -17
rect 487 -85 499 -51
rect 533 -85 545 -51
rect 487 -100 545 -85
rect 745 85 803 100
rect 745 51 757 85
rect 791 51 803 85
rect 745 17 803 51
rect 745 -17 757 17
rect 791 -17 803 17
rect 745 -51 803 -17
rect 745 -85 757 -51
rect 791 -85 803 -51
rect 745 -100 803 -85
rect 1003 85 1061 100
rect 1003 51 1015 85
rect 1049 51 1061 85
rect 1003 17 1061 51
rect 1003 -17 1015 17
rect 1049 -17 1061 17
rect 1003 -51 1061 -17
rect 1003 -85 1015 -51
rect 1049 -85 1061 -51
rect 1003 -100 1061 -85
rect 1261 85 1319 100
rect 1261 51 1273 85
rect 1307 51 1319 85
rect 1261 17 1319 51
rect 1261 -17 1273 17
rect 1307 -17 1319 17
rect 1261 -51 1319 -17
rect 1261 -85 1273 -51
rect 1307 -85 1319 -51
rect 1261 -100 1319 -85
<< pdiffc >>
rect -1307 51 -1273 85
rect -1307 -17 -1273 17
rect -1307 -85 -1273 -51
rect -1049 51 -1015 85
rect -1049 -17 -1015 17
rect -1049 -85 -1015 -51
rect -791 51 -757 85
rect -791 -17 -757 17
rect -791 -85 -757 -51
rect -533 51 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -51
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
rect 499 51 533 85
rect 499 -17 533 17
rect 499 -85 533 -51
rect 757 51 791 85
rect 757 -17 791 17
rect 757 -85 791 -51
rect 1015 51 1049 85
rect 1015 -17 1049 17
rect 1015 -85 1049 -51
rect 1273 51 1307 85
rect 1273 -17 1307 17
rect 1273 -85 1307 -51
<< poly >>
rect -1261 181 -1061 197
rect -1261 147 -1212 181
rect -1178 147 -1144 181
rect -1110 147 -1061 181
rect -1261 100 -1061 147
rect -1003 181 -803 197
rect -1003 147 -954 181
rect -920 147 -886 181
rect -852 147 -803 181
rect -1003 100 -803 147
rect -745 181 -545 197
rect -745 147 -696 181
rect -662 147 -628 181
rect -594 147 -545 181
rect -745 100 -545 147
rect -487 181 -287 197
rect -487 147 -438 181
rect -404 147 -370 181
rect -336 147 -287 181
rect -487 100 -287 147
rect -229 181 -29 197
rect -229 147 -180 181
rect -146 147 -112 181
rect -78 147 -29 181
rect -229 100 -29 147
rect 29 181 229 197
rect 29 147 78 181
rect 112 147 146 181
rect 180 147 229 181
rect 29 100 229 147
rect 287 181 487 197
rect 287 147 336 181
rect 370 147 404 181
rect 438 147 487 181
rect 287 100 487 147
rect 545 181 745 197
rect 545 147 594 181
rect 628 147 662 181
rect 696 147 745 181
rect 545 100 745 147
rect 803 181 1003 197
rect 803 147 852 181
rect 886 147 920 181
rect 954 147 1003 181
rect 803 100 1003 147
rect 1061 181 1261 197
rect 1061 147 1110 181
rect 1144 147 1178 181
rect 1212 147 1261 181
rect 1061 100 1261 147
rect -1261 -147 -1061 -100
rect -1261 -181 -1212 -147
rect -1178 -181 -1144 -147
rect -1110 -181 -1061 -147
rect -1261 -197 -1061 -181
rect -1003 -147 -803 -100
rect -1003 -181 -954 -147
rect -920 -181 -886 -147
rect -852 -181 -803 -147
rect -1003 -197 -803 -181
rect -745 -147 -545 -100
rect -745 -181 -696 -147
rect -662 -181 -628 -147
rect -594 -181 -545 -147
rect -745 -197 -545 -181
rect -487 -147 -287 -100
rect -487 -181 -438 -147
rect -404 -181 -370 -147
rect -336 -181 -287 -147
rect -487 -197 -287 -181
rect -229 -147 -29 -100
rect -229 -181 -180 -147
rect -146 -181 -112 -147
rect -78 -181 -29 -147
rect -229 -197 -29 -181
rect 29 -147 229 -100
rect 29 -181 78 -147
rect 112 -181 146 -147
rect 180 -181 229 -147
rect 29 -197 229 -181
rect 287 -147 487 -100
rect 287 -181 336 -147
rect 370 -181 404 -147
rect 438 -181 487 -147
rect 287 -197 487 -181
rect 545 -147 745 -100
rect 545 -181 594 -147
rect 628 -181 662 -147
rect 696 -181 745 -147
rect 545 -197 745 -181
rect 803 -147 1003 -100
rect 803 -181 852 -147
rect 886 -181 920 -147
rect 954 -181 1003 -147
rect 803 -197 1003 -181
rect 1061 -147 1261 -100
rect 1061 -181 1110 -147
rect 1144 -181 1178 -147
rect 1212 -181 1261 -147
rect 1061 -197 1261 -181
<< polycont >>
rect -1212 147 -1178 181
rect -1144 147 -1110 181
rect -954 147 -920 181
rect -886 147 -852 181
rect -696 147 -662 181
rect -628 147 -594 181
rect -438 147 -404 181
rect -370 147 -336 181
rect -180 147 -146 181
rect -112 147 -78 181
rect 78 147 112 181
rect 146 147 180 181
rect 336 147 370 181
rect 404 147 438 181
rect 594 147 628 181
rect 662 147 696 181
rect 852 147 886 181
rect 920 147 954 181
rect 1110 147 1144 181
rect 1178 147 1212 181
rect -1212 -181 -1178 -147
rect -1144 -181 -1110 -147
rect -954 -181 -920 -147
rect -886 -181 -852 -147
rect -696 -181 -662 -147
rect -628 -181 -594 -147
rect -438 -181 -404 -147
rect -370 -181 -336 -147
rect -180 -181 -146 -147
rect -112 -181 -78 -147
rect 78 -181 112 -147
rect 146 -181 180 -147
rect 336 -181 370 -147
rect 404 -181 438 -147
rect 594 -181 628 -147
rect 662 -181 696 -147
rect 852 -181 886 -147
rect 920 -181 954 -147
rect 1110 -181 1144 -147
rect 1178 -181 1212 -147
<< locali >>
rect -1261 147 -1212 181
rect -1110 147 -1061 181
rect -1003 147 -954 181
rect -852 147 -803 181
rect -745 147 -696 181
rect -594 147 -545 181
rect -487 147 -438 181
rect -336 147 -287 181
rect -229 147 -180 181
rect -78 147 -29 181
rect 29 147 78 181
rect 180 147 229 181
rect 287 147 336 181
rect 438 147 487 181
rect 545 147 594 181
rect 696 147 745 181
rect 803 147 852 181
rect 954 147 1003 181
rect 1061 147 1110 181
rect 1212 147 1261 181
rect -1307 85 -1273 104
rect -1307 17 -1273 19
rect -1307 -19 -1273 -17
rect -1307 -104 -1273 -85
rect -1049 85 -1015 104
rect -1049 17 -1015 19
rect -1049 -19 -1015 -17
rect -1049 -104 -1015 -85
rect -791 85 -757 104
rect -791 17 -757 19
rect -791 -19 -757 -17
rect -791 -104 -757 -85
rect -533 85 -499 104
rect -533 17 -499 19
rect -533 -19 -499 -17
rect -533 -104 -499 -85
rect -275 85 -241 104
rect -275 17 -241 19
rect -275 -19 -241 -17
rect -275 -104 -241 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 241 85 275 104
rect 241 17 275 19
rect 241 -19 275 -17
rect 241 -104 275 -85
rect 499 85 533 104
rect 499 17 533 19
rect 499 -19 533 -17
rect 499 -104 533 -85
rect 757 85 791 104
rect 757 17 791 19
rect 757 -19 791 -17
rect 757 -104 791 -85
rect 1015 85 1049 104
rect 1015 17 1049 19
rect 1015 -19 1049 -17
rect 1015 -104 1049 -85
rect 1273 85 1307 104
rect 1273 17 1307 19
rect 1273 -19 1307 -17
rect 1273 -104 1307 -85
rect -1261 -181 -1212 -147
rect -1110 -181 -1061 -147
rect -1003 -181 -954 -147
rect -852 -181 -803 -147
rect -745 -181 -696 -147
rect -594 -181 -545 -147
rect -487 -181 -438 -147
rect -336 -181 -287 -147
rect -229 -181 -180 -147
rect -78 -181 -29 -147
rect 29 -181 78 -147
rect 180 -181 229 -147
rect 287 -181 336 -147
rect 438 -181 487 -147
rect 545 -181 594 -147
rect 696 -181 745 -147
rect 803 -181 852 -147
rect 954 -181 1003 -147
rect 1061 -181 1110 -147
rect 1212 -181 1261 -147
<< viali >>
rect -1178 147 -1144 181
rect -920 147 -886 181
rect -662 147 -628 181
rect -404 147 -370 181
rect -146 147 -112 181
rect 112 147 146 181
rect 370 147 404 181
rect 628 147 662 181
rect 886 147 920 181
rect 1144 147 1178 181
rect -1307 51 -1273 53
rect -1307 19 -1273 51
rect -1307 -51 -1273 -19
rect -1307 -53 -1273 -51
rect -1049 51 -1015 53
rect -1049 19 -1015 51
rect -1049 -51 -1015 -19
rect -1049 -53 -1015 -51
rect -791 51 -757 53
rect -791 19 -757 51
rect -791 -51 -757 -19
rect -791 -53 -757 -51
rect -533 51 -499 53
rect -533 19 -499 51
rect -533 -51 -499 -19
rect -533 -53 -499 -51
rect -275 51 -241 53
rect -275 19 -241 51
rect -275 -51 -241 -19
rect -275 -53 -241 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 241 51 275 53
rect 241 19 275 51
rect 241 -51 275 -19
rect 241 -53 275 -51
rect 499 51 533 53
rect 499 19 533 51
rect 499 -51 533 -19
rect 499 -53 533 -51
rect 757 51 791 53
rect 757 19 791 51
rect 757 -51 791 -19
rect 757 -53 791 -51
rect 1015 51 1049 53
rect 1015 19 1049 51
rect 1015 -51 1049 -19
rect 1015 -53 1049 -51
rect 1273 51 1307 53
rect 1273 19 1307 51
rect 1273 -51 1307 -19
rect 1273 -53 1307 -51
rect -1178 -181 -1144 -147
rect -920 -181 -886 -147
rect -662 -181 -628 -147
rect -404 -181 -370 -147
rect -146 -181 -112 -147
rect 112 -181 146 -147
rect 370 -181 404 -147
rect 628 -181 662 -147
rect 886 -181 920 -147
rect 1144 -181 1178 -147
<< metal1 >>
rect -1215 181 -1107 187
rect -1215 147 -1178 181
rect -1144 147 -1107 181
rect -1215 141 -1107 147
rect -957 181 -849 187
rect -957 147 -920 181
rect -886 147 -849 181
rect -957 141 -849 147
rect -699 181 -591 187
rect -699 147 -662 181
rect -628 147 -591 181
rect -699 141 -591 147
rect -441 181 -333 187
rect -441 147 -404 181
rect -370 147 -333 181
rect -441 141 -333 147
rect -183 181 -75 187
rect -183 147 -146 181
rect -112 147 -75 181
rect -183 141 -75 147
rect 75 181 183 187
rect 75 147 112 181
rect 146 147 183 181
rect 75 141 183 147
rect 333 181 441 187
rect 333 147 370 181
rect 404 147 441 181
rect 333 141 441 147
rect 591 181 699 187
rect 591 147 628 181
rect 662 147 699 181
rect 591 141 699 147
rect 849 181 957 187
rect 849 147 886 181
rect 920 147 957 181
rect 849 141 957 147
rect 1107 181 1215 187
rect 1107 147 1144 181
rect 1178 147 1215 181
rect 1107 141 1215 147
rect -1313 53 -1267 100
rect -1313 19 -1307 53
rect -1273 19 -1267 53
rect -1313 -19 -1267 19
rect -1313 -53 -1307 -19
rect -1273 -53 -1267 -19
rect -1313 -100 -1267 -53
rect -1055 53 -1009 100
rect -1055 19 -1049 53
rect -1015 19 -1009 53
rect -1055 -19 -1009 19
rect -1055 -53 -1049 -19
rect -1015 -53 -1009 -19
rect -1055 -100 -1009 -53
rect -797 53 -751 100
rect -797 19 -791 53
rect -757 19 -751 53
rect -797 -19 -751 19
rect -797 -53 -791 -19
rect -757 -53 -751 -19
rect -797 -100 -751 -53
rect -539 53 -493 100
rect -539 19 -533 53
rect -499 19 -493 53
rect -539 -19 -493 19
rect -539 -53 -533 -19
rect -499 -53 -493 -19
rect -539 -100 -493 -53
rect -281 53 -235 100
rect -281 19 -275 53
rect -241 19 -235 53
rect -281 -19 -235 19
rect -281 -53 -275 -19
rect -241 -53 -235 -19
rect -281 -100 -235 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 235 53 281 100
rect 235 19 241 53
rect 275 19 281 53
rect 235 -19 281 19
rect 235 -53 241 -19
rect 275 -53 281 -19
rect 235 -100 281 -53
rect 493 53 539 100
rect 493 19 499 53
rect 533 19 539 53
rect 493 -19 539 19
rect 493 -53 499 -19
rect 533 -53 539 -19
rect 493 -100 539 -53
rect 751 53 797 100
rect 751 19 757 53
rect 791 19 797 53
rect 751 -19 797 19
rect 751 -53 757 -19
rect 791 -53 797 -19
rect 751 -100 797 -53
rect 1009 53 1055 100
rect 1009 19 1015 53
rect 1049 19 1055 53
rect 1009 -19 1055 19
rect 1009 -53 1015 -19
rect 1049 -53 1055 -19
rect 1009 -100 1055 -53
rect 1267 53 1313 100
rect 1267 19 1273 53
rect 1307 19 1313 53
rect 1267 -19 1313 19
rect 1267 -53 1273 -19
rect 1307 -53 1313 -19
rect 1267 -100 1313 -53
rect -1215 -147 -1107 -141
rect -1215 -181 -1178 -147
rect -1144 -181 -1107 -147
rect -1215 -187 -1107 -181
rect -957 -147 -849 -141
rect -957 -181 -920 -147
rect -886 -181 -849 -147
rect -957 -187 -849 -181
rect -699 -147 -591 -141
rect -699 -181 -662 -147
rect -628 -181 -591 -147
rect -699 -187 -591 -181
rect -441 -147 -333 -141
rect -441 -181 -404 -147
rect -370 -181 -333 -147
rect -441 -187 -333 -181
rect -183 -147 -75 -141
rect -183 -181 -146 -147
rect -112 -181 -75 -147
rect -183 -187 -75 -181
rect 75 -147 183 -141
rect 75 -181 112 -147
rect 146 -181 183 -147
rect 75 -187 183 -181
rect 333 -147 441 -141
rect 333 -181 370 -147
rect 404 -181 441 -147
rect 333 -187 441 -181
rect 591 -147 699 -141
rect 591 -181 628 -147
rect 662 -181 699 -147
rect 591 -187 699 -181
rect 849 -147 957 -141
rect 849 -181 886 -147
rect 920 -181 957 -147
rect 849 -187 957 -181
rect 1107 -147 1215 -141
rect 1107 -181 1144 -147
rect 1178 -181 1215 -147
rect 1107 -187 1215 -181
<< end >>
