magic
tech sky130A
magscale 1 2
timestamp 1621486730
<< pwell >>
rect -941 -310 941 310
<< nmos >>
rect -745 -100 -545 100
rect -487 -100 -287 100
rect -229 -100 -29 100
rect 29 -100 229 100
rect 287 -100 487 100
rect 545 -100 745 100
<< ndiff >>
rect -803 88 -745 100
rect -803 -88 -791 88
rect -757 -88 -745 88
rect -803 -100 -745 -88
rect -545 88 -487 100
rect -545 -88 -533 88
rect -499 -88 -487 88
rect -545 -100 -487 -88
rect -287 88 -229 100
rect -287 -88 -275 88
rect -241 -88 -229 88
rect -287 -100 -229 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 229 88 287 100
rect 229 -88 241 88
rect 275 -88 287 88
rect 229 -100 287 -88
rect 487 88 545 100
rect 487 -88 499 88
rect 533 -88 545 88
rect 487 -100 545 -88
rect 745 88 803 100
rect 745 -88 757 88
rect 791 -88 803 88
rect 745 -100 803 -88
<< ndiffc >>
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
<< psubdiff >>
rect -905 240 -809 274
rect 809 240 905 274
rect -905 178 -871 240
rect 871 178 905 240
rect -905 -240 -871 -178
rect 871 -240 905 -178
rect -905 -274 -809 -240
rect 809 -274 905 -240
<< psubdiffcont >>
rect -809 240 809 274
rect -905 -178 -871 178
rect 871 -178 905 178
rect -809 -274 809 -240
<< poly >>
rect -703 172 -587 188
rect -703 155 -687 172
rect -745 138 -687 155
rect -603 155 -587 172
rect -445 172 -329 188
rect -445 155 -429 172
rect -603 138 -545 155
rect -745 100 -545 138
rect -487 138 -429 155
rect -345 155 -329 172
rect -187 172 -71 188
rect -187 155 -171 172
rect -345 138 -287 155
rect -487 100 -287 138
rect -229 138 -171 155
rect -87 155 -71 172
rect 71 172 187 188
rect 71 155 87 172
rect -87 138 -29 155
rect -229 100 -29 138
rect 29 138 87 155
rect 171 155 187 172
rect 329 172 445 188
rect 329 155 345 172
rect 171 138 229 155
rect 29 100 229 138
rect 287 138 345 155
rect 429 155 445 172
rect 587 172 703 188
rect 587 155 603 172
rect 429 138 487 155
rect 287 100 487 138
rect 545 138 603 155
rect 687 155 703 172
rect 687 138 745 155
rect 545 100 745 138
rect -745 -138 -545 -100
rect -745 -155 -687 -138
rect -703 -172 -687 -155
rect -603 -155 -545 -138
rect -487 -138 -287 -100
rect -487 -155 -429 -138
rect -603 -172 -587 -155
rect -703 -188 -587 -172
rect -445 -172 -429 -155
rect -345 -155 -287 -138
rect -229 -138 -29 -100
rect -229 -155 -171 -138
rect -345 -172 -329 -155
rect -445 -188 -329 -172
rect -187 -172 -171 -155
rect -87 -155 -29 -138
rect 29 -138 229 -100
rect 29 -155 87 -138
rect -87 -172 -71 -155
rect -187 -188 -71 -172
rect 71 -172 87 -155
rect 171 -155 229 -138
rect 287 -138 487 -100
rect 287 -155 345 -138
rect 171 -172 187 -155
rect 71 -188 187 -172
rect 329 -172 345 -155
rect 429 -155 487 -138
rect 545 -138 745 -100
rect 545 -155 603 -138
rect 429 -172 445 -155
rect 329 -188 445 -172
rect 587 -172 603 -155
rect 687 -155 745 -138
rect 687 -172 703 -155
rect 587 -188 703 -172
<< polycont >>
rect -687 138 -603 172
rect -429 138 -345 172
rect -171 138 -87 172
rect 87 138 171 172
rect 345 138 429 172
rect 603 138 687 172
rect -687 -172 -603 -138
rect -429 -172 -345 -138
rect -171 -172 -87 -138
rect 87 -172 171 -138
rect 345 -172 429 -138
rect 603 -172 687 -138
<< locali >>
rect -905 240 -809 274
rect 809 240 905 274
rect -905 178 -871 240
rect 871 178 905 240
rect -703 138 -687 172
rect -603 138 -587 172
rect -445 138 -429 172
rect -345 138 -329 172
rect -187 138 -171 172
rect -87 138 -71 172
rect 71 138 87 172
rect 171 138 187 172
rect 329 138 345 172
rect 429 138 445 172
rect 587 138 603 172
rect 687 138 703 172
rect -791 88 -757 104
rect -791 -104 -757 -88
rect -533 88 -499 104
rect -533 -104 -499 -88
rect -275 88 -241 104
rect -275 -104 -241 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 241 88 275 104
rect 241 -104 275 -88
rect 499 88 533 104
rect 499 -104 533 -88
rect 757 88 791 104
rect 757 -104 791 -88
rect -703 -172 -687 -138
rect -603 -172 -587 -138
rect -445 -172 -429 -138
rect -345 -172 -329 -138
rect -187 -172 -171 -138
rect -87 -172 -71 -138
rect 71 -172 87 -138
rect 171 -172 187 -138
rect 329 -172 345 -138
rect 429 -172 445 -138
rect 587 -172 603 -138
rect 687 -172 703 -138
rect -905 -240 -871 -178
rect 871 -240 905 -178
rect -905 -274 -809 -240
rect 809 -274 905 -240
<< viali >>
rect -687 138 -603 172
rect -429 138 -345 172
rect -171 138 -87 172
rect 87 138 171 172
rect 345 138 429 172
rect 603 138 687 172
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
rect -687 -172 -603 -138
rect -429 -172 -345 -138
rect -171 -172 -87 -138
rect 87 -172 171 -138
rect 345 -172 429 -138
rect 603 -172 687 -138
<< metal1 >>
rect -699 172 -591 178
rect -699 138 -687 172
rect -603 138 -591 172
rect -699 132 -591 138
rect -441 172 -333 178
rect -441 138 -429 172
rect -345 138 -333 172
rect -441 132 -333 138
rect -183 172 -75 178
rect -183 138 -171 172
rect -87 138 -75 172
rect -183 132 -75 138
rect 75 172 183 178
rect 75 138 87 172
rect 171 138 183 172
rect 75 132 183 138
rect 333 172 441 178
rect 333 138 345 172
rect 429 138 441 172
rect 333 132 441 138
rect 591 172 699 178
rect 591 138 603 172
rect 687 138 699 172
rect 591 132 699 138
rect -797 88 -751 100
rect -797 -88 -791 88
rect -757 -88 -751 88
rect -797 -100 -751 -88
rect -539 88 -493 100
rect -539 -88 -533 88
rect -499 -88 -493 88
rect -539 -100 -493 -88
rect -281 88 -235 100
rect -281 -88 -275 88
rect -241 -88 -235 88
rect -281 -100 -235 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 235 88 281 100
rect 235 -88 241 88
rect 275 -88 281 88
rect 235 -100 281 -88
rect 493 88 539 100
rect 493 -88 499 88
rect 533 -88 539 88
rect 493 -100 539 -88
rect 751 88 797 100
rect 751 -88 757 88
rect 791 -88 797 88
rect 751 -100 797 -88
rect -699 -138 -591 -132
rect -699 -172 -687 -138
rect -603 -172 -591 -138
rect -699 -178 -591 -172
rect -441 -138 -333 -132
rect -441 -172 -429 -138
rect -345 -172 -333 -138
rect -441 -178 -333 -172
rect -183 -138 -75 -132
rect -183 -172 -171 -138
rect -87 -172 -75 -138
rect -183 -178 -75 -172
rect 75 -138 183 -132
rect 75 -172 87 -138
rect 171 -172 183 -138
rect 75 -178 183 -172
rect 333 -138 441 -132
rect 333 -172 345 -138
rect 429 -172 441 -138
rect 333 -178 441 -172
rect 591 -138 699 -132
rect 591 -172 603 -138
rect 687 -172 699 -138
rect 591 -178 699 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -888 -257 888 257
string parameters w 1 l 1 m 1 nf 6 diffcov 100 polycov 50 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
